magic
tech gf180mcuB
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 453 4006 1094
<< pwell >>
rect -86 -86 4006 453
<< mvnmos >>
rect 150 175 270 333
rect 374 175 494 333
rect 742 159 862 277
rect 966 159 1086 277
rect 1190 159 1310 277
rect 1358 159 1478 277
rect 1658 215 1778 333
rect 1882 215 2002 333
rect 2106 215 2226 333
rect 2412 69 2532 333
rect 2636 69 2756 333
rect 3004 69 3124 333
rect 3228 69 3348 333
rect 3452 69 3572 333
rect 3676 69 3796 333
<< mvpmos >>
rect 170 573 270 849
rect 374 573 474 849
rect 762 573 862 773
rect 986 573 1086 773
rect 1190 573 1290 773
rect 1378 573 1478 773
rect 1658 573 1758 773
rect 1881 573 1981 773
rect 2192 573 2292 773
rect 2432 573 2532 939
rect 2636 573 2736 939
rect 3024 573 3124 939
rect 3228 573 3328 939
rect 3432 573 3532 939
rect 3636 573 3736 939
<< mvndiff >>
rect 62 320 150 333
rect 62 274 75 320
rect 121 274 150 320
rect 62 175 150 274
rect 270 234 374 333
rect 270 188 299 234
rect 345 188 374 234
rect 270 175 374 188
rect 494 320 582 333
rect 494 274 523 320
rect 569 274 582 320
rect 1578 277 1658 333
rect 494 175 582 274
rect 654 218 742 277
rect 654 172 667 218
rect 713 172 742 218
rect 654 159 742 172
rect 862 264 966 277
rect 862 218 891 264
rect 937 218 966 264
rect 862 159 966 218
rect 1086 264 1190 277
rect 1086 218 1115 264
rect 1161 218 1190 264
rect 1086 159 1190 218
rect 1310 159 1358 277
rect 1478 215 1658 277
rect 1778 320 1882 333
rect 1778 274 1807 320
rect 1853 274 1882 320
rect 1778 215 1882 274
rect 2002 320 2106 333
rect 2002 274 2031 320
rect 2077 274 2106 320
rect 2002 215 2106 274
rect 2226 287 2412 333
rect 2226 215 2337 287
rect 1478 159 1598 215
rect 1538 127 1598 159
rect 1538 114 1610 127
rect 2324 147 2337 215
rect 2383 147 2412 287
rect 1538 68 1551 114
rect 1597 68 1610 114
rect 2324 69 2412 147
rect 2532 128 2636 333
rect 2532 82 2561 128
rect 2607 82 2636 128
rect 2532 69 2636 82
rect 2756 320 2844 333
rect 2756 274 2785 320
rect 2831 274 2844 320
rect 2756 69 2844 274
rect 2916 128 3004 333
rect 2916 82 2929 128
rect 2975 82 3004 128
rect 2916 69 3004 82
rect 3124 320 3228 333
rect 3124 274 3153 320
rect 3199 274 3228 320
rect 3124 69 3228 274
rect 3348 128 3452 333
rect 3348 82 3377 128
rect 3423 82 3452 128
rect 3348 69 3452 82
rect 3572 320 3676 333
rect 3572 274 3601 320
rect 3647 274 3676 320
rect 3572 69 3676 274
rect 3796 222 3884 333
rect 3796 82 3825 222
rect 3871 82 3884 222
rect 3796 69 3884 82
rect 1538 55 1610 68
<< mvpdiff >>
rect 82 739 170 849
rect 82 599 95 739
rect 141 599 170 739
rect 82 573 170 599
rect 270 836 374 849
rect 270 696 299 836
rect 345 696 374 836
rect 270 573 374 696
rect 474 632 562 849
rect 2352 773 2432 939
rect 474 586 503 632
rect 549 586 562 632
rect 474 573 562 586
rect 674 760 762 773
rect 674 714 687 760
rect 733 714 762 760
rect 674 573 762 714
rect 862 726 986 773
rect 862 586 911 726
rect 957 586 986 726
rect 862 573 986 586
rect 1086 726 1190 773
rect 1086 586 1115 726
rect 1161 586 1190 726
rect 1086 573 1190 586
rect 1290 573 1378 773
rect 1478 760 1658 773
rect 1478 620 1507 760
rect 1553 620 1658 760
rect 1478 573 1658 620
rect 1758 726 1881 773
rect 1758 586 1806 726
rect 1852 586 1881 726
rect 1758 573 1881 586
rect 1981 726 2192 773
rect 1981 586 2031 726
rect 2077 586 2192 726
rect 1981 573 2192 586
rect 2292 746 2432 773
rect 2292 700 2357 746
rect 2403 700 2432 746
rect 2292 573 2432 700
rect 2532 926 2636 939
rect 2532 880 2561 926
rect 2607 880 2636 926
rect 2532 573 2636 880
rect 2736 632 2824 939
rect 2736 586 2765 632
rect 2811 586 2824 632
rect 2736 573 2824 586
rect 2936 926 3024 939
rect 2936 880 2949 926
rect 2995 880 3024 926
rect 2936 573 3024 880
rect 3124 635 3228 939
rect 3124 589 3153 635
rect 3199 589 3228 635
rect 3124 573 3228 589
rect 3328 926 3432 939
rect 3328 880 3357 926
rect 3403 880 3432 926
rect 3328 573 3432 880
rect 3532 635 3636 939
rect 3532 589 3561 635
rect 3607 589 3636 635
rect 3532 573 3636 589
rect 3736 926 3824 939
rect 3736 880 3765 926
rect 3811 880 3824 926
rect 3736 573 3824 880
<< mvndiffc >>
rect 75 274 121 320
rect 299 188 345 234
rect 523 274 569 320
rect 667 172 713 218
rect 891 218 937 264
rect 1115 218 1161 264
rect 1807 274 1853 320
rect 2031 274 2077 320
rect 2337 147 2383 287
rect 1551 68 1597 114
rect 2561 82 2607 128
rect 2785 274 2831 320
rect 2929 82 2975 128
rect 3153 274 3199 320
rect 3377 82 3423 128
rect 3601 274 3647 320
rect 3825 82 3871 222
<< mvpdiffc >>
rect 95 599 141 739
rect 299 696 345 836
rect 503 586 549 632
rect 687 714 733 760
rect 911 586 957 726
rect 1115 586 1161 726
rect 1507 620 1553 760
rect 1806 586 1852 726
rect 2031 586 2077 726
rect 2357 700 2403 746
rect 2561 880 2607 926
rect 2765 586 2811 632
rect 2949 880 2995 926
rect 3153 589 3199 635
rect 3357 880 3403 926
rect 3561 589 3607 635
rect 3765 880 3811 926
<< polysilicon >>
rect 374 909 1086 949
rect 2432 939 2532 983
rect 2636 939 2736 983
rect 3024 939 3124 983
rect 3228 939 3328 983
rect 3432 939 3532 983
rect 3636 939 3736 983
rect 170 849 270 893
rect 374 849 474 909
rect 762 773 862 817
rect 986 773 1086 909
rect 1190 865 1981 905
rect 1190 852 1290 865
rect 1190 806 1203 852
rect 1249 806 1290 852
rect 1190 773 1290 806
rect 1378 773 1478 817
rect 1658 773 1758 817
rect 1881 773 1981 865
rect 2192 773 2292 817
rect 170 523 270 573
rect 170 477 183 523
rect 229 477 270 523
rect 170 377 270 477
rect 150 333 270 377
rect 374 412 474 573
rect 374 366 387 412
rect 433 377 474 412
rect 762 512 862 573
rect 986 529 1086 573
rect 762 466 801 512
rect 847 466 862 512
rect 1190 481 1290 573
rect 433 366 494 377
rect 374 333 494 366
rect 762 321 862 466
rect 742 277 862 321
rect 966 441 1290 481
rect 1378 540 1478 573
rect 1378 494 1419 540
rect 1465 494 1478 540
rect 966 277 1086 441
rect 1190 356 1310 369
rect 1190 310 1251 356
rect 1297 310 1310 356
rect 1378 321 1478 494
rect 1658 437 1758 573
rect 1881 513 1981 573
rect 2192 540 2292 573
rect 2192 529 2233 540
rect 1881 473 2146 513
rect 2220 494 2233 529
rect 2279 494 2292 540
rect 2220 481 2292 494
rect 1658 391 1671 437
rect 1717 391 1758 437
rect 1658 377 1758 391
rect 2106 377 2146 473
rect 2432 430 2532 573
rect 2432 384 2473 430
rect 2519 384 2532 430
rect 2432 377 2532 384
rect 1658 333 1778 377
rect 1882 333 2002 377
rect 2106 333 2226 377
rect 2412 333 2532 377
rect 2636 540 2736 573
rect 2636 494 2649 540
rect 2695 494 2736 540
rect 2636 377 2736 494
rect 3024 465 3124 573
rect 3228 465 3328 573
rect 3432 465 3532 573
rect 3636 465 3736 573
rect 3024 431 3736 465
rect 3024 385 3037 431
rect 3083 393 3260 431
rect 3083 385 3124 393
rect 3024 377 3124 385
rect 2636 333 2756 377
rect 3004 333 3124 377
rect 3228 385 3260 393
rect 3306 393 3465 431
rect 3306 385 3348 393
rect 3228 333 3348 385
rect 3452 385 3465 393
rect 3511 393 3736 431
rect 3511 385 3572 393
rect 3452 333 3572 385
rect 3676 377 3736 393
rect 3676 333 3796 377
rect 1190 277 1310 310
rect 1358 277 1478 321
rect 150 131 270 175
rect 374 67 494 175
rect 1658 171 1778 215
rect 1882 182 2002 215
rect 742 115 862 159
rect 966 115 1086 159
rect 1190 67 1310 159
rect 1358 115 1478 159
rect 1882 136 1895 182
rect 1941 136 2002 182
rect 2106 171 2226 215
rect 374 27 1310 67
rect 1882 123 2002 136
rect 2412 25 2532 69
rect 2636 25 2756 69
rect 3004 25 3124 69
rect 3228 25 3348 69
rect 3452 25 3572 69
rect 3676 25 3796 69
<< polycontact >>
rect 1203 806 1249 852
rect 183 477 229 523
rect 387 366 433 412
rect 801 466 847 512
rect 1419 494 1465 540
rect 1251 310 1297 356
rect 2233 494 2279 540
rect 1671 391 1717 437
rect 2473 384 2519 430
rect 2649 494 2695 540
rect 3037 385 3083 431
rect 3260 385 3306 431
rect 3465 385 3511 431
rect 1895 136 1941 182
<< metal1 >>
rect 0 926 3920 1098
rect 0 918 2561 926
rect 299 836 345 918
rect 95 739 141 750
rect 687 760 733 918
rect 687 703 733 714
rect 779 806 1203 852
rect 1249 806 1260 852
rect 299 685 345 696
rect 779 643 825 806
rect 1507 760 1553 918
rect 2607 918 2949 926
rect 2561 869 2607 880
rect 2995 918 3357 926
rect 2949 869 2995 880
rect 3403 918 3765 926
rect 3357 869 3403 880
rect 3811 918 3920 926
rect 3765 869 3811 880
rect 141 599 433 634
rect 95 588 433 599
rect 142 523 341 542
rect 142 477 183 523
rect 229 477 341 523
rect 142 466 341 477
rect 387 412 433 588
rect 75 366 387 401
rect 75 355 433 366
rect 503 632 825 643
rect 549 597 825 632
rect 911 726 958 737
rect 549 586 569 597
rect 75 320 121 355
rect 75 263 121 274
rect 503 320 569 586
rect 957 586 958 726
rect 911 575 958 586
rect 686 512 866 542
rect 686 466 801 512
rect 847 466 866 512
rect 503 274 523 320
rect 912 275 958 575
rect 503 263 569 274
rect 891 264 958 275
rect 299 234 345 245
rect 299 90 345 188
rect 667 218 713 229
rect 937 218 958 264
rect 891 207 958 218
rect 1115 726 1161 737
rect 1507 609 1553 620
rect 1806 726 1853 737
rect 1115 448 1161 586
rect 1852 586 1853 726
rect 1806 540 1853 586
rect 1408 494 1419 540
rect 1465 494 1853 540
rect 1115 437 1717 448
rect 1115 402 1671 437
rect 1115 264 1161 402
rect 1671 380 1717 391
rect 1115 207 1161 218
rect 1240 310 1251 356
rect 1297 310 1308 356
rect 1240 217 1308 310
rect 1807 320 1853 494
rect 1807 263 1853 274
rect 2031 726 2077 737
rect 2346 700 2357 746
rect 2403 700 3750 746
rect 2077 597 2371 643
rect 2031 320 2077 586
rect 2031 263 2077 274
rect 2233 540 2279 551
rect 2325 540 2371 597
rect 2765 632 2811 643
rect 2325 494 2649 540
rect 2695 494 2706 540
rect 2233 217 2279 494
rect 2765 442 2811 586
rect 3142 635 3658 646
rect 3142 589 3153 635
rect 3199 589 3561 635
rect 3607 589 3658 635
rect 3142 578 3658 589
rect 2765 431 3511 442
rect 2765 430 3037 431
rect 2462 384 2473 430
rect 2519 385 3037 430
rect 3083 385 3260 431
rect 3306 385 3465 431
rect 2519 384 3511 385
rect 2774 374 3511 384
rect 2774 320 2842 374
rect 3557 328 3658 578
rect 667 90 713 172
rect 1240 182 2279 217
rect 1240 171 1895 182
rect 1884 136 1895 171
rect 1941 136 2279 182
rect 2337 287 2383 298
rect 2774 274 2785 320
rect 2831 274 2842 320
rect 3142 320 3658 328
rect 3142 274 3153 320
rect 3199 274 3601 320
rect 3647 274 3658 320
rect 3704 228 3750 700
rect 2383 182 3750 228
rect 3825 222 3871 233
rect 2337 136 2383 147
rect 1551 114 1597 125
rect 0 68 1551 90
rect 2550 90 2561 128
rect 1597 82 2561 90
rect 2607 90 2618 128
rect 2918 90 2929 128
rect 2607 82 2929 90
rect 2975 90 2986 128
rect 3366 90 3377 128
rect 2975 82 3377 90
rect 3423 90 3434 128
rect 3423 82 3825 90
rect 3871 82 3920 90
rect 1597 68 3920 82
rect 0 -90 3920 68
<< labels >>
flabel metal1 s 142 466 341 542 0 FreeSans 200 0 0 0 CLKN
port 2 nsew clock input
flabel metal1 s 686 466 866 542 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 3142 578 3658 646 0 FreeSans 200 0 0 0 Q
port 3 nsew default output
flabel metal1 s 0 918 3920 1098 0 FreeSans 200 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 299 233 345 245 0 FreeSans 200 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 5 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 6 nsew ground bidirectional
rlabel metal1 s 3557 328 3658 578 1 Q
port 3 nsew default output
rlabel metal1 s 3142 274 3658 328 1 Q
port 3 nsew default output
rlabel metal1 s 3765 869 3811 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3357 869 3403 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2949 869 2995 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2561 869 2607 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1507 869 1553 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 687 869 733 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 299 869 345 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1507 703 1553 869 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 687 703 733 869 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 299 703 345 869 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1507 685 1553 703 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 299 685 345 703 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1507 609 1553 685 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3825 229 3871 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 299 229 345 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3825 128 3871 229 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 667 128 713 229 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 299 128 345 229 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3825 125 3871 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3366 125 3434 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2918 125 2986 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2550 125 2618 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 667 125 713 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 299 125 345 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3825 90 3871 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3366 90 3434 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2918 90 2986 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2550 90 2618 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1551 90 1597 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 667 90 713 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 299 90 345 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 3920 90 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3920 1008
string GDS_END 1509848
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1501426
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
