magic
tech gf180mcuD
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 352 310 870
<< pwell >>
rect -86 -86 310 352
<< mvpsubdiff >>
rect 56 226 168 256
rect 56 79 89 226
rect 135 79 168 226
rect 56 56 168 79
<< mvnsubdiff >>
rect 72 699 152 712
rect 72 653 89 699
rect 135 653 152 699
rect 72 571 152 653
rect 72 525 89 571
rect 135 525 152 571
rect 72 443 152 525
rect 72 397 89 443
rect 135 397 152 443
rect 72 384 152 397
<< mvpsubdiffcont >>
rect 89 79 135 226
<< mvnsubdiffcont >>
rect 89 653 135 699
rect 89 525 135 571
rect 89 397 135 443
<< metal1 >>
rect 0 724 224 844
rect 78 699 146 724
rect 78 653 89 699
rect 135 653 146 699
rect 78 571 146 653
rect 78 525 89 571
rect 135 525 146 571
rect 78 443 146 525
rect 78 397 89 443
rect 135 397 146 443
rect 78 386 146 397
rect 78 226 146 237
rect 78 79 89 226
rect 135 79 146 226
rect 78 60 146 79
rect 0 -60 224 60
<< labels >>
flabel metal1 s 0 724 224 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 78 60 146 237 0 FreeSans 400 0 0 0 VSS
port 2 nsew ground bidirectional abutment
rlabel metal1 s 78 386 146 724 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 0 -60 224 60 1 VSS
port 2 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 224 784
string GDS_END 423770
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 422058
string LEFclass core WELLTAP
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
