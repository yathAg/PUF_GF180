magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
use M3_M2$$43368492_256x8m81_0  M3_M2$$43368492_256x8m81_0_0
timestamp 1698431365
transform 1 0 5251 0 1 11281
box 0 0 1 1
use M3_M2$$43368492_256x8m81_0  M3_M2$$43368492_256x8m81_0_1
timestamp 1698431365
transform 1 0 12629 0 1 11281
box 0 0 1 1
use M3_M2$$43368492_256x8m81_0  M3_M2$$43368492_256x8m81_0_2
timestamp 1698431365
transform 1 0 23115 0 1 11281
box 0 0 1 1
use M3_M2$$47115308_256x8m81  M3_M2$$47115308_256x8m81_0
timestamp 1698431365
transform 1 0 4256 0 1 12090
box 0 0 1 1
use M3_M2$$47115308_256x8m81  M3_M2$$47115308_256x8m81_1
timestamp 1698431365
transform 1 0 22120 0 1 12090
box 0 0 1 1
use M3_M2$$201412652_256x8m81  M3_M2$$201412652_256x8m81_0
timestamp 1698431365
transform 1 0 15172 0 1 12090
box 0 0 1 1
use xpredec0_256x8m81  xpredec0_256x8m81_0
timestamp 1698431365
transform 1 0 7704 0 1 0
box 0 -1 7186 11377
use xpredec0_256x8m81  xpredec0_256x8m81_1
timestamp 1698431365
transform 1 0 325 0 1 0
box 0 -1 7186 11377
use xpredec1_256x8m81  xpredec1_256x8m81_0
timestamp 1698431365
transform 1 0 15082 0 1 0
box 287 -1 11984 10577
<< properties >>
string GDS_END 1831090
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 1827360
<< end >>
