magic
tech gf180mcuA
magscale 1 10
timestamp 1698431365
<< nwell >>
rect 29138 51874 56005 52390
rect 29138 50321 32850 51874
rect 35260 50809 39818 51874
rect 35260 50633 39436 50809
rect 45169 50633 49764 51874
rect 52285 50633 56005 51874
<< pwell >>
rect 1774 51482 24710 51514
rect 1774 35138 24710 35170
<< mvpsubdiff >>
rect 27479 52963 28511 53046
rect 27479 1117 27498 52963
rect 27744 52942 28511 52963
rect 27744 35996 27846 52942
rect 28492 51528 28511 52942
rect 56613 52963 57645 53046
rect 56613 52942 57380 52963
rect 56613 51528 56632 52942
rect 28492 35996 28911 51528
rect 27744 35977 28911 35996
rect 56256 35996 56632 51528
rect 57278 35996 57380 52942
rect 56256 35977 57380 35996
rect 27744 34621 27763 35977
rect 57361 34621 57380 35977
rect 27744 34602 57380 34621
rect 27744 34256 27846 34602
rect 57292 34256 57380 34602
rect 27744 34237 57380 34256
rect 27744 1117 27763 34237
rect 28620 3906 40188 3925
rect 28620 3860 28639 3906
rect 28685 3860 28755 3906
rect 28801 3860 28871 3906
rect 28917 3860 28987 3906
rect 29033 3860 29103 3906
rect 29149 3860 29219 3906
rect 29265 3860 29335 3906
rect 29381 3860 29451 3906
rect 29497 3860 29567 3906
rect 29613 3860 29683 3906
rect 29729 3860 29799 3906
rect 29845 3860 29915 3906
rect 29961 3860 30031 3906
rect 30077 3860 30147 3906
rect 30193 3860 30263 3906
rect 30309 3860 30379 3906
rect 30425 3860 30495 3906
rect 30541 3860 30611 3906
rect 30657 3860 30727 3906
rect 30773 3860 30843 3906
rect 30889 3860 30959 3906
rect 31005 3860 31075 3906
rect 31121 3860 31191 3906
rect 31237 3860 31307 3906
rect 31353 3860 31423 3906
rect 31469 3860 31539 3906
rect 31585 3860 31655 3906
rect 31701 3860 31771 3906
rect 31817 3860 31887 3906
rect 31933 3860 32003 3906
rect 32049 3860 32119 3906
rect 32165 3860 32235 3906
rect 32281 3860 32351 3906
rect 32397 3860 32467 3906
rect 32513 3860 32583 3906
rect 32629 3860 32699 3906
rect 32745 3860 32815 3906
rect 32861 3860 32931 3906
rect 32977 3860 33047 3906
rect 33093 3860 33163 3906
rect 33209 3860 33279 3906
rect 33325 3860 33395 3906
rect 33441 3860 33511 3906
rect 33557 3860 33627 3906
rect 33673 3860 33743 3906
rect 33789 3860 33859 3906
rect 33905 3860 33975 3906
rect 34021 3860 34091 3906
rect 34137 3860 34207 3906
rect 34253 3860 34323 3906
rect 34369 3860 34439 3906
rect 34485 3860 34555 3906
rect 34601 3860 34671 3906
rect 34717 3860 34787 3906
rect 34833 3860 34903 3906
rect 34949 3860 35019 3906
rect 35065 3860 35135 3906
rect 35181 3860 35251 3906
rect 35297 3860 35367 3906
rect 35413 3860 35483 3906
rect 35529 3860 35599 3906
rect 35645 3860 35715 3906
rect 35761 3860 35831 3906
rect 35877 3860 35947 3906
rect 35993 3860 36063 3906
rect 36109 3860 36179 3906
rect 36225 3860 36295 3906
rect 36341 3860 36411 3906
rect 36457 3860 36527 3906
rect 36573 3860 36643 3906
rect 36689 3860 36759 3906
rect 36805 3860 36875 3906
rect 36921 3860 36991 3906
rect 37037 3860 37107 3906
rect 37153 3860 37223 3906
rect 37269 3860 37339 3906
rect 37385 3860 37455 3906
rect 37501 3860 37571 3906
rect 37617 3860 37687 3906
rect 37733 3860 37803 3906
rect 37849 3860 37919 3906
rect 37965 3860 38035 3906
rect 38081 3860 38151 3906
rect 38197 3860 38267 3906
rect 38313 3860 38383 3906
rect 38429 3860 38499 3906
rect 38545 3860 38615 3906
rect 38661 3860 38731 3906
rect 38777 3860 38847 3906
rect 38893 3860 38963 3906
rect 39009 3860 39079 3906
rect 39125 3860 39195 3906
rect 39241 3860 39311 3906
rect 39357 3860 39427 3906
rect 39473 3860 39543 3906
rect 39589 3860 39659 3906
rect 39705 3860 39775 3906
rect 39821 3860 39891 3906
rect 39937 3860 40007 3906
rect 40053 3860 40123 3906
rect 40169 3860 40188 3906
rect 28620 3790 40188 3860
rect 28620 3744 28639 3790
rect 28685 3744 28755 3790
rect 28801 3744 28871 3790
rect 28917 3744 28987 3790
rect 29033 3744 29103 3790
rect 29149 3744 29219 3790
rect 29265 3744 29335 3790
rect 29381 3744 29451 3790
rect 29497 3744 29567 3790
rect 29613 3744 29683 3790
rect 29729 3744 29799 3790
rect 29845 3744 29915 3790
rect 29961 3744 30031 3790
rect 30077 3744 30147 3790
rect 30193 3744 30263 3790
rect 30309 3744 30379 3790
rect 30425 3744 30495 3790
rect 30541 3744 30611 3790
rect 30657 3744 30727 3790
rect 30773 3744 30843 3790
rect 30889 3744 30959 3790
rect 31005 3744 31075 3790
rect 31121 3744 31191 3790
rect 31237 3744 31307 3790
rect 31353 3744 31423 3790
rect 31469 3744 31539 3790
rect 31585 3744 31655 3790
rect 31701 3744 31771 3790
rect 31817 3744 31887 3790
rect 31933 3744 32003 3790
rect 32049 3744 32119 3790
rect 32165 3744 32235 3790
rect 32281 3744 32351 3790
rect 32397 3744 32467 3790
rect 32513 3744 32583 3790
rect 32629 3744 32699 3790
rect 32745 3744 32815 3790
rect 32861 3744 32931 3790
rect 32977 3744 33047 3790
rect 33093 3744 33163 3790
rect 33209 3744 33279 3790
rect 33325 3744 33395 3790
rect 33441 3744 33511 3790
rect 33557 3744 33627 3790
rect 33673 3744 33743 3790
rect 33789 3744 33859 3790
rect 33905 3744 33975 3790
rect 34021 3744 34091 3790
rect 34137 3744 34207 3790
rect 34253 3744 34323 3790
rect 34369 3744 34439 3790
rect 34485 3744 34555 3790
rect 34601 3744 34671 3790
rect 34717 3744 34787 3790
rect 34833 3744 34903 3790
rect 34949 3744 35019 3790
rect 35065 3744 35135 3790
rect 35181 3744 35251 3790
rect 35297 3744 35367 3790
rect 35413 3744 35483 3790
rect 35529 3744 35599 3790
rect 35645 3744 35715 3790
rect 35761 3744 35831 3790
rect 35877 3744 35947 3790
rect 35993 3744 36063 3790
rect 36109 3744 36179 3790
rect 36225 3744 36295 3790
rect 36341 3744 36411 3790
rect 36457 3744 36527 3790
rect 36573 3744 36643 3790
rect 36689 3744 36759 3790
rect 36805 3744 36875 3790
rect 36921 3744 36991 3790
rect 37037 3744 37107 3790
rect 37153 3744 37223 3790
rect 37269 3744 37339 3790
rect 37385 3744 37455 3790
rect 37501 3744 37571 3790
rect 37617 3744 37687 3790
rect 37733 3744 37803 3790
rect 37849 3744 37919 3790
rect 37965 3744 38035 3790
rect 38081 3744 38151 3790
rect 38197 3744 38267 3790
rect 38313 3744 38383 3790
rect 38429 3744 38499 3790
rect 38545 3744 38615 3790
rect 38661 3744 38731 3790
rect 38777 3744 38847 3790
rect 38893 3744 38963 3790
rect 39009 3744 39079 3790
rect 39125 3744 39195 3790
rect 39241 3744 39311 3790
rect 39357 3744 39427 3790
rect 39473 3744 39543 3790
rect 39589 3744 39659 3790
rect 39705 3744 39775 3790
rect 39821 3744 39891 3790
rect 39937 3744 40007 3790
rect 40053 3744 40123 3790
rect 40169 3744 40188 3790
rect 28620 3674 40188 3744
rect 28620 3628 28639 3674
rect 28685 3628 28755 3674
rect 28801 3628 28871 3674
rect 28917 3628 28987 3674
rect 29033 3628 29103 3674
rect 29149 3628 29219 3674
rect 29265 3628 29335 3674
rect 29381 3628 29451 3674
rect 29497 3628 29567 3674
rect 29613 3628 29683 3674
rect 29729 3628 29799 3674
rect 29845 3628 29915 3674
rect 29961 3628 30031 3674
rect 30077 3628 30147 3674
rect 30193 3628 30263 3674
rect 30309 3628 30379 3674
rect 30425 3628 30495 3674
rect 30541 3628 30611 3674
rect 30657 3628 30727 3674
rect 30773 3628 30843 3674
rect 30889 3628 30959 3674
rect 31005 3628 31075 3674
rect 31121 3628 31191 3674
rect 31237 3628 31307 3674
rect 31353 3628 31423 3674
rect 31469 3628 31539 3674
rect 31585 3628 31655 3674
rect 31701 3628 31771 3674
rect 31817 3628 31887 3674
rect 31933 3628 32003 3674
rect 32049 3628 32119 3674
rect 32165 3628 32235 3674
rect 32281 3628 32351 3674
rect 32397 3628 32467 3674
rect 32513 3628 32583 3674
rect 32629 3628 32699 3674
rect 32745 3628 32815 3674
rect 32861 3628 32931 3674
rect 32977 3628 33047 3674
rect 33093 3628 33163 3674
rect 33209 3628 33279 3674
rect 33325 3628 33395 3674
rect 33441 3628 33511 3674
rect 33557 3628 33627 3674
rect 33673 3628 33743 3674
rect 33789 3628 33859 3674
rect 33905 3628 33975 3674
rect 34021 3628 34091 3674
rect 34137 3628 34207 3674
rect 34253 3628 34323 3674
rect 34369 3628 34439 3674
rect 34485 3628 34555 3674
rect 34601 3628 34671 3674
rect 34717 3628 34787 3674
rect 34833 3628 34903 3674
rect 34949 3628 35019 3674
rect 35065 3628 35135 3674
rect 35181 3628 35251 3674
rect 35297 3628 35367 3674
rect 35413 3628 35483 3674
rect 35529 3628 35599 3674
rect 35645 3628 35715 3674
rect 35761 3628 35831 3674
rect 35877 3628 35947 3674
rect 35993 3628 36063 3674
rect 36109 3628 36179 3674
rect 36225 3628 36295 3674
rect 36341 3628 36411 3674
rect 36457 3628 36527 3674
rect 36573 3628 36643 3674
rect 36689 3628 36759 3674
rect 36805 3628 36875 3674
rect 36921 3628 36991 3674
rect 37037 3628 37107 3674
rect 37153 3628 37223 3674
rect 37269 3628 37339 3674
rect 37385 3628 37455 3674
rect 37501 3628 37571 3674
rect 37617 3628 37687 3674
rect 37733 3628 37803 3674
rect 37849 3628 37919 3674
rect 37965 3628 38035 3674
rect 38081 3628 38151 3674
rect 38197 3628 38267 3674
rect 38313 3628 38383 3674
rect 38429 3628 38499 3674
rect 38545 3628 38615 3674
rect 38661 3628 38731 3674
rect 38777 3628 38847 3674
rect 38893 3628 38963 3674
rect 39009 3628 39079 3674
rect 39125 3628 39195 3674
rect 39241 3628 39311 3674
rect 39357 3628 39427 3674
rect 39473 3628 39543 3674
rect 39589 3628 39659 3674
rect 39705 3628 39775 3674
rect 39821 3628 39891 3674
rect 39937 3628 40007 3674
rect 40053 3628 40123 3674
rect 40169 3628 40188 3674
rect 28620 3558 40188 3628
rect 28620 3512 28639 3558
rect 28685 3512 28755 3558
rect 28801 3512 28871 3558
rect 28917 3512 28987 3558
rect 29033 3512 29103 3558
rect 29149 3512 29219 3558
rect 29265 3512 29335 3558
rect 29381 3512 29451 3558
rect 29497 3512 29567 3558
rect 29613 3512 29683 3558
rect 29729 3512 29799 3558
rect 29845 3512 29915 3558
rect 29961 3512 30031 3558
rect 30077 3512 30147 3558
rect 30193 3512 30263 3558
rect 30309 3512 30379 3558
rect 30425 3512 30495 3558
rect 30541 3512 30611 3558
rect 30657 3512 30727 3558
rect 30773 3512 30843 3558
rect 30889 3512 30959 3558
rect 31005 3512 31075 3558
rect 31121 3512 31191 3558
rect 31237 3512 31307 3558
rect 31353 3512 31423 3558
rect 31469 3512 31539 3558
rect 31585 3512 31655 3558
rect 31701 3512 31771 3558
rect 31817 3512 31887 3558
rect 31933 3512 32003 3558
rect 32049 3512 32119 3558
rect 32165 3512 32235 3558
rect 32281 3512 32351 3558
rect 32397 3512 32467 3558
rect 32513 3512 32583 3558
rect 32629 3512 32699 3558
rect 32745 3512 32815 3558
rect 32861 3512 32931 3558
rect 32977 3512 33047 3558
rect 33093 3512 33163 3558
rect 33209 3512 33279 3558
rect 33325 3512 33395 3558
rect 33441 3512 33511 3558
rect 33557 3512 33627 3558
rect 33673 3512 33743 3558
rect 33789 3512 33859 3558
rect 33905 3512 33975 3558
rect 34021 3512 34091 3558
rect 34137 3512 34207 3558
rect 34253 3512 34323 3558
rect 34369 3512 34439 3558
rect 34485 3512 34555 3558
rect 34601 3512 34671 3558
rect 34717 3512 34787 3558
rect 34833 3512 34903 3558
rect 34949 3512 35019 3558
rect 35065 3512 35135 3558
rect 35181 3512 35251 3558
rect 35297 3512 35367 3558
rect 35413 3512 35483 3558
rect 35529 3512 35599 3558
rect 35645 3512 35715 3558
rect 35761 3512 35831 3558
rect 35877 3512 35947 3558
rect 35993 3512 36063 3558
rect 36109 3512 36179 3558
rect 36225 3512 36295 3558
rect 36341 3512 36411 3558
rect 36457 3512 36527 3558
rect 36573 3512 36643 3558
rect 36689 3512 36759 3558
rect 36805 3512 36875 3558
rect 36921 3512 36991 3558
rect 37037 3512 37107 3558
rect 37153 3512 37223 3558
rect 37269 3512 37339 3558
rect 37385 3512 37455 3558
rect 37501 3512 37571 3558
rect 37617 3512 37687 3558
rect 37733 3512 37803 3558
rect 37849 3512 37919 3558
rect 37965 3512 38035 3558
rect 38081 3512 38151 3558
rect 38197 3512 38267 3558
rect 38313 3512 38383 3558
rect 38429 3512 38499 3558
rect 38545 3512 38615 3558
rect 38661 3512 38731 3558
rect 38777 3512 38847 3558
rect 38893 3512 38963 3558
rect 39009 3512 39079 3558
rect 39125 3512 39195 3558
rect 39241 3512 39311 3558
rect 39357 3512 39427 3558
rect 39473 3512 39543 3558
rect 39589 3512 39659 3558
rect 39705 3512 39775 3558
rect 39821 3512 39891 3558
rect 39937 3512 40007 3558
rect 40053 3512 40123 3558
rect 40169 3512 40188 3558
rect 28620 3442 40188 3512
rect 28620 3396 28639 3442
rect 28685 3396 28755 3442
rect 28801 3396 28871 3442
rect 28917 3396 28987 3442
rect 29033 3396 29103 3442
rect 29149 3396 29219 3442
rect 29265 3396 29335 3442
rect 29381 3396 29451 3442
rect 29497 3396 29567 3442
rect 29613 3396 29683 3442
rect 29729 3396 29799 3442
rect 29845 3396 29915 3442
rect 29961 3396 30031 3442
rect 30077 3396 30147 3442
rect 30193 3396 30263 3442
rect 30309 3396 30379 3442
rect 30425 3396 30495 3442
rect 30541 3396 30611 3442
rect 30657 3396 30727 3442
rect 30773 3396 30843 3442
rect 30889 3396 30959 3442
rect 31005 3396 31075 3442
rect 31121 3396 31191 3442
rect 31237 3396 31307 3442
rect 31353 3396 31423 3442
rect 31469 3396 31539 3442
rect 31585 3396 31655 3442
rect 31701 3396 31771 3442
rect 31817 3396 31887 3442
rect 31933 3396 32003 3442
rect 32049 3396 32119 3442
rect 32165 3396 32235 3442
rect 32281 3396 32351 3442
rect 32397 3396 32467 3442
rect 32513 3396 32583 3442
rect 32629 3396 32699 3442
rect 32745 3396 32815 3442
rect 32861 3396 32931 3442
rect 32977 3396 33047 3442
rect 33093 3396 33163 3442
rect 33209 3396 33279 3442
rect 33325 3396 33395 3442
rect 33441 3396 33511 3442
rect 33557 3396 33627 3442
rect 33673 3396 33743 3442
rect 33789 3396 33859 3442
rect 33905 3396 33975 3442
rect 34021 3396 34091 3442
rect 34137 3396 34207 3442
rect 34253 3396 34323 3442
rect 34369 3396 34439 3442
rect 34485 3396 34555 3442
rect 34601 3396 34671 3442
rect 34717 3396 34787 3442
rect 34833 3396 34903 3442
rect 34949 3396 35019 3442
rect 35065 3396 35135 3442
rect 35181 3396 35251 3442
rect 35297 3396 35367 3442
rect 35413 3396 35483 3442
rect 35529 3396 35599 3442
rect 35645 3396 35715 3442
rect 35761 3396 35831 3442
rect 35877 3396 35947 3442
rect 35993 3396 36063 3442
rect 36109 3396 36179 3442
rect 36225 3396 36295 3442
rect 36341 3396 36411 3442
rect 36457 3396 36527 3442
rect 36573 3396 36643 3442
rect 36689 3396 36759 3442
rect 36805 3396 36875 3442
rect 36921 3396 36991 3442
rect 37037 3396 37107 3442
rect 37153 3396 37223 3442
rect 37269 3396 37339 3442
rect 37385 3396 37455 3442
rect 37501 3396 37571 3442
rect 37617 3396 37687 3442
rect 37733 3396 37803 3442
rect 37849 3396 37919 3442
rect 37965 3396 38035 3442
rect 38081 3396 38151 3442
rect 38197 3396 38267 3442
rect 38313 3396 38383 3442
rect 38429 3396 38499 3442
rect 38545 3396 38615 3442
rect 38661 3396 38731 3442
rect 38777 3396 38847 3442
rect 38893 3396 38963 3442
rect 39009 3396 39079 3442
rect 39125 3396 39195 3442
rect 39241 3396 39311 3442
rect 39357 3396 39427 3442
rect 39473 3396 39543 3442
rect 39589 3396 39659 3442
rect 39705 3396 39775 3442
rect 39821 3396 39891 3442
rect 39937 3396 40007 3442
rect 40053 3396 40123 3442
rect 40169 3396 40188 3442
rect 28620 3326 40188 3396
rect 28620 3280 28639 3326
rect 28685 3280 28755 3326
rect 28801 3280 28871 3326
rect 28917 3280 28987 3326
rect 29033 3280 29103 3326
rect 29149 3280 29219 3326
rect 29265 3280 29335 3326
rect 29381 3280 29451 3326
rect 29497 3280 29567 3326
rect 29613 3280 29683 3326
rect 29729 3280 29799 3326
rect 29845 3280 29915 3326
rect 29961 3280 30031 3326
rect 30077 3280 30147 3326
rect 30193 3280 30263 3326
rect 30309 3280 30379 3326
rect 30425 3280 30495 3326
rect 30541 3280 30611 3326
rect 30657 3280 30727 3326
rect 30773 3280 30843 3326
rect 30889 3280 30959 3326
rect 31005 3280 31075 3326
rect 31121 3280 31191 3326
rect 31237 3280 31307 3326
rect 31353 3280 31423 3326
rect 31469 3280 31539 3326
rect 31585 3280 31655 3326
rect 31701 3280 31771 3326
rect 31817 3280 31887 3326
rect 31933 3280 32003 3326
rect 32049 3280 32119 3326
rect 32165 3280 32235 3326
rect 32281 3280 32351 3326
rect 32397 3280 32467 3326
rect 32513 3280 32583 3326
rect 32629 3280 32699 3326
rect 32745 3280 32815 3326
rect 32861 3280 32931 3326
rect 32977 3280 33047 3326
rect 33093 3280 33163 3326
rect 33209 3280 33279 3326
rect 33325 3280 33395 3326
rect 33441 3280 33511 3326
rect 33557 3280 33627 3326
rect 33673 3280 33743 3326
rect 33789 3280 33859 3326
rect 33905 3280 33975 3326
rect 34021 3280 34091 3326
rect 34137 3280 34207 3326
rect 34253 3280 34323 3326
rect 34369 3280 34439 3326
rect 34485 3280 34555 3326
rect 34601 3280 34671 3326
rect 34717 3280 34787 3326
rect 34833 3280 34903 3326
rect 34949 3280 35019 3326
rect 35065 3280 35135 3326
rect 35181 3280 35251 3326
rect 35297 3280 35367 3326
rect 35413 3280 35483 3326
rect 35529 3280 35599 3326
rect 35645 3280 35715 3326
rect 35761 3280 35831 3326
rect 35877 3280 35947 3326
rect 35993 3280 36063 3326
rect 36109 3280 36179 3326
rect 36225 3280 36295 3326
rect 36341 3280 36411 3326
rect 36457 3280 36527 3326
rect 36573 3280 36643 3326
rect 36689 3280 36759 3326
rect 36805 3280 36875 3326
rect 36921 3280 36991 3326
rect 37037 3280 37107 3326
rect 37153 3280 37223 3326
rect 37269 3280 37339 3326
rect 37385 3280 37455 3326
rect 37501 3280 37571 3326
rect 37617 3280 37687 3326
rect 37733 3280 37803 3326
rect 37849 3280 37919 3326
rect 37965 3280 38035 3326
rect 38081 3280 38151 3326
rect 38197 3280 38267 3326
rect 38313 3280 38383 3326
rect 38429 3280 38499 3326
rect 38545 3280 38615 3326
rect 38661 3280 38731 3326
rect 38777 3280 38847 3326
rect 38893 3280 38963 3326
rect 39009 3280 39079 3326
rect 39125 3280 39195 3326
rect 39241 3280 39311 3326
rect 39357 3280 39427 3326
rect 39473 3280 39543 3326
rect 39589 3280 39659 3326
rect 39705 3280 39775 3326
rect 39821 3280 39891 3326
rect 39937 3280 40007 3326
rect 40053 3280 40123 3326
rect 40169 3280 40188 3326
rect 28620 3210 40188 3280
rect 28620 3164 28639 3210
rect 28685 3164 28755 3210
rect 28801 3164 28871 3210
rect 28917 3164 28987 3210
rect 29033 3164 29103 3210
rect 29149 3164 29219 3210
rect 29265 3164 29335 3210
rect 29381 3164 29451 3210
rect 29497 3164 29567 3210
rect 29613 3164 29683 3210
rect 29729 3164 29799 3210
rect 29845 3164 29915 3210
rect 29961 3164 30031 3210
rect 30077 3164 30147 3210
rect 30193 3164 30263 3210
rect 30309 3164 30379 3210
rect 30425 3164 30495 3210
rect 30541 3164 30611 3210
rect 30657 3164 30727 3210
rect 30773 3164 30843 3210
rect 30889 3164 30959 3210
rect 31005 3164 31075 3210
rect 31121 3164 31191 3210
rect 31237 3164 31307 3210
rect 31353 3164 31423 3210
rect 31469 3164 31539 3210
rect 31585 3164 31655 3210
rect 31701 3164 31771 3210
rect 31817 3164 31887 3210
rect 31933 3164 32003 3210
rect 32049 3164 32119 3210
rect 32165 3164 32235 3210
rect 32281 3164 32351 3210
rect 32397 3164 32467 3210
rect 32513 3164 32583 3210
rect 32629 3164 32699 3210
rect 32745 3164 32815 3210
rect 32861 3164 32931 3210
rect 32977 3164 33047 3210
rect 33093 3164 33163 3210
rect 33209 3164 33279 3210
rect 33325 3164 33395 3210
rect 33441 3164 33511 3210
rect 33557 3164 33627 3210
rect 33673 3164 33743 3210
rect 33789 3164 33859 3210
rect 33905 3164 33975 3210
rect 34021 3164 34091 3210
rect 34137 3164 34207 3210
rect 34253 3164 34323 3210
rect 34369 3164 34439 3210
rect 34485 3164 34555 3210
rect 34601 3164 34671 3210
rect 34717 3164 34787 3210
rect 34833 3164 34903 3210
rect 34949 3164 35019 3210
rect 35065 3164 35135 3210
rect 35181 3164 35251 3210
rect 35297 3164 35367 3210
rect 35413 3164 35483 3210
rect 35529 3164 35599 3210
rect 35645 3164 35715 3210
rect 35761 3164 35831 3210
rect 35877 3164 35947 3210
rect 35993 3164 36063 3210
rect 36109 3164 36179 3210
rect 36225 3164 36295 3210
rect 36341 3164 36411 3210
rect 36457 3164 36527 3210
rect 36573 3164 36643 3210
rect 36689 3164 36759 3210
rect 36805 3164 36875 3210
rect 36921 3164 36991 3210
rect 37037 3164 37107 3210
rect 37153 3164 37223 3210
rect 37269 3164 37339 3210
rect 37385 3164 37455 3210
rect 37501 3164 37571 3210
rect 37617 3164 37687 3210
rect 37733 3164 37803 3210
rect 37849 3164 37919 3210
rect 37965 3164 38035 3210
rect 38081 3164 38151 3210
rect 38197 3164 38267 3210
rect 38313 3164 38383 3210
rect 38429 3164 38499 3210
rect 38545 3164 38615 3210
rect 38661 3164 38731 3210
rect 38777 3164 38847 3210
rect 38893 3164 38963 3210
rect 39009 3164 39079 3210
rect 39125 3164 39195 3210
rect 39241 3164 39311 3210
rect 39357 3164 39427 3210
rect 39473 3164 39543 3210
rect 39589 3164 39659 3210
rect 39705 3164 39775 3210
rect 39821 3164 39891 3210
rect 39937 3164 40007 3210
rect 40053 3164 40123 3210
rect 40169 3164 40188 3210
rect 28620 3094 40188 3164
rect 28620 3048 28639 3094
rect 28685 3048 28755 3094
rect 28801 3048 28871 3094
rect 28917 3048 28987 3094
rect 29033 3048 29103 3094
rect 29149 3048 29219 3094
rect 29265 3048 29335 3094
rect 29381 3048 29451 3094
rect 29497 3048 29567 3094
rect 29613 3048 29683 3094
rect 29729 3048 29799 3094
rect 29845 3048 29915 3094
rect 29961 3048 30031 3094
rect 30077 3048 30147 3094
rect 30193 3048 30263 3094
rect 30309 3048 30379 3094
rect 30425 3048 30495 3094
rect 30541 3048 30611 3094
rect 30657 3048 30727 3094
rect 30773 3048 30843 3094
rect 30889 3048 30959 3094
rect 31005 3048 31075 3094
rect 31121 3048 31191 3094
rect 31237 3048 31307 3094
rect 31353 3048 31423 3094
rect 31469 3048 31539 3094
rect 31585 3048 31655 3094
rect 31701 3048 31771 3094
rect 31817 3048 31887 3094
rect 31933 3048 32003 3094
rect 32049 3048 32119 3094
rect 32165 3048 32235 3094
rect 32281 3048 32351 3094
rect 32397 3048 32467 3094
rect 32513 3048 32583 3094
rect 32629 3048 32699 3094
rect 32745 3048 32815 3094
rect 32861 3048 32931 3094
rect 32977 3048 33047 3094
rect 33093 3048 33163 3094
rect 33209 3048 33279 3094
rect 33325 3048 33395 3094
rect 33441 3048 33511 3094
rect 33557 3048 33627 3094
rect 33673 3048 33743 3094
rect 33789 3048 33859 3094
rect 33905 3048 33975 3094
rect 34021 3048 34091 3094
rect 34137 3048 34207 3094
rect 34253 3048 34323 3094
rect 34369 3048 34439 3094
rect 34485 3048 34555 3094
rect 34601 3048 34671 3094
rect 34717 3048 34787 3094
rect 34833 3048 34903 3094
rect 34949 3048 35019 3094
rect 35065 3048 35135 3094
rect 35181 3048 35251 3094
rect 35297 3048 35367 3094
rect 35413 3048 35483 3094
rect 35529 3048 35599 3094
rect 35645 3048 35715 3094
rect 35761 3048 35831 3094
rect 35877 3048 35947 3094
rect 35993 3048 36063 3094
rect 36109 3048 36179 3094
rect 36225 3048 36295 3094
rect 36341 3048 36411 3094
rect 36457 3048 36527 3094
rect 36573 3048 36643 3094
rect 36689 3048 36759 3094
rect 36805 3048 36875 3094
rect 36921 3048 36991 3094
rect 37037 3048 37107 3094
rect 37153 3048 37223 3094
rect 37269 3048 37339 3094
rect 37385 3048 37455 3094
rect 37501 3048 37571 3094
rect 37617 3048 37687 3094
rect 37733 3048 37803 3094
rect 37849 3048 37919 3094
rect 37965 3048 38035 3094
rect 38081 3048 38151 3094
rect 38197 3048 38267 3094
rect 38313 3048 38383 3094
rect 38429 3048 38499 3094
rect 38545 3048 38615 3094
rect 38661 3048 38731 3094
rect 38777 3048 38847 3094
rect 38893 3048 38963 3094
rect 39009 3048 39079 3094
rect 39125 3048 39195 3094
rect 39241 3048 39311 3094
rect 39357 3048 39427 3094
rect 39473 3048 39543 3094
rect 39589 3048 39659 3094
rect 39705 3048 39775 3094
rect 39821 3048 39891 3094
rect 39937 3048 40007 3094
rect 40053 3048 40123 3094
rect 40169 3048 40188 3094
rect 28620 2978 40188 3048
rect 28620 2932 28639 2978
rect 28685 2932 28755 2978
rect 28801 2932 28871 2978
rect 28917 2932 28987 2978
rect 29033 2932 29103 2978
rect 29149 2932 29219 2978
rect 29265 2932 29335 2978
rect 29381 2932 29451 2978
rect 29497 2932 29567 2978
rect 29613 2932 29683 2978
rect 29729 2932 29799 2978
rect 29845 2932 29915 2978
rect 29961 2932 30031 2978
rect 30077 2932 30147 2978
rect 30193 2932 30263 2978
rect 30309 2932 30379 2978
rect 30425 2932 30495 2978
rect 30541 2932 30611 2978
rect 30657 2932 30727 2978
rect 30773 2932 30843 2978
rect 30889 2932 30959 2978
rect 31005 2932 31075 2978
rect 31121 2932 31191 2978
rect 31237 2932 31307 2978
rect 31353 2932 31423 2978
rect 31469 2932 31539 2978
rect 31585 2932 31655 2978
rect 31701 2932 31771 2978
rect 31817 2932 31887 2978
rect 31933 2932 32003 2978
rect 32049 2932 32119 2978
rect 32165 2932 32235 2978
rect 32281 2932 32351 2978
rect 32397 2932 32467 2978
rect 32513 2932 32583 2978
rect 32629 2932 32699 2978
rect 32745 2932 32815 2978
rect 32861 2932 32931 2978
rect 32977 2932 33047 2978
rect 33093 2932 33163 2978
rect 33209 2932 33279 2978
rect 33325 2932 33395 2978
rect 33441 2932 33511 2978
rect 33557 2932 33627 2978
rect 33673 2932 33743 2978
rect 33789 2932 33859 2978
rect 33905 2932 33975 2978
rect 34021 2932 34091 2978
rect 34137 2932 34207 2978
rect 34253 2932 34323 2978
rect 34369 2932 34439 2978
rect 34485 2932 34555 2978
rect 34601 2932 34671 2978
rect 34717 2932 34787 2978
rect 34833 2932 34903 2978
rect 34949 2932 35019 2978
rect 35065 2932 35135 2978
rect 35181 2932 35251 2978
rect 35297 2932 35367 2978
rect 35413 2932 35483 2978
rect 35529 2932 35599 2978
rect 35645 2932 35715 2978
rect 35761 2932 35831 2978
rect 35877 2932 35947 2978
rect 35993 2932 36063 2978
rect 36109 2932 36179 2978
rect 36225 2932 36295 2978
rect 36341 2932 36411 2978
rect 36457 2932 36527 2978
rect 36573 2932 36643 2978
rect 36689 2932 36759 2978
rect 36805 2932 36875 2978
rect 36921 2932 36991 2978
rect 37037 2932 37107 2978
rect 37153 2932 37223 2978
rect 37269 2932 37339 2978
rect 37385 2932 37455 2978
rect 37501 2932 37571 2978
rect 37617 2932 37687 2978
rect 37733 2932 37803 2978
rect 37849 2932 37919 2978
rect 37965 2932 38035 2978
rect 38081 2932 38151 2978
rect 38197 2932 38267 2978
rect 38313 2932 38383 2978
rect 38429 2932 38499 2978
rect 38545 2932 38615 2978
rect 38661 2932 38731 2978
rect 38777 2932 38847 2978
rect 38893 2932 38963 2978
rect 39009 2932 39079 2978
rect 39125 2932 39195 2978
rect 39241 2932 39311 2978
rect 39357 2932 39427 2978
rect 39473 2932 39543 2978
rect 39589 2932 39659 2978
rect 39705 2932 39775 2978
rect 39821 2932 39891 2978
rect 39937 2932 40007 2978
rect 40053 2932 40123 2978
rect 40169 2932 40188 2978
rect 28620 2862 40188 2932
rect 28620 2816 28639 2862
rect 28685 2816 28755 2862
rect 28801 2816 28871 2862
rect 28917 2816 28987 2862
rect 29033 2816 29103 2862
rect 29149 2816 29219 2862
rect 29265 2816 29335 2862
rect 29381 2816 29451 2862
rect 29497 2816 29567 2862
rect 29613 2816 29683 2862
rect 29729 2816 29799 2862
rect 29845 2816 29915 2862
rect 29961 2816 30031 2862
rect 30077 2816 30147 2862
rect 30193 2816 30263 2862
rect 30309 2816 30379 2862
rect 30425 2816 30495 2862
rect 30541 2816 30611 2862
rect 30657 2816 30727 2862
rect 30773 2816 30843 2862
rect 30889 2816 30959 2862
rect 31005 2816 31075 2862
rect 31121 2816 31191 2862
rect 31237 2816 31307 2862
rect 31353 2816 31423 2862
rect 31469 2816 31539 2862
rect 31585 2816 31655 2862
rect 31701 2816 31771 2862
rect 31817 2816 31887 2862
rect 31933 2816 32003 2862
rect 32049 2816 32119 2862
rect 32165 2816 32235 2862
rect 32281 2816 32351 2862
rect 32397 2816 32467 2862
rect 32513 2816 32583 2862
rect 32629 2816 32699 2862
rect 32745 2816 32815 2862
rect 32861 2816 32931 2862
rect 32977 2816 33047 2862
rect 33093 2816 33163 2862
rect 33209 2816 33279 2862
rect 33325 2816 33395 2862
rect 33441 2816 33511 2862
rect 33557 2816 33627 2862
rect 33673 2816 33743 2862
rect 33789 2816 33859 2862
rect 33905 2816 33975 2862
rect 34021 2816 34091 2862
rect 34137 2816 34207 2862
rect 34253 2816 34323 2862
rect 34369 2816 34439 2862
rect 34485 2816 34555 2862
rect 34601 2816 34671 2862
rect 34717 2816 34787 2862
rect 34833 2816 34903 2862
rect 34949 2816 35019 2862
rect 35065 2816 35135 2862
rect 35181 2816 35251 2862
rect 35297 2816 35367 2862
rect 35413 2816 35483 2862
rect 35529 2816 35599 2862
rect 35645 2816 35715 2862
rect 35761 2816 35831 2862
rect 35877 2816 35947 2862
rect 35993 2816 36063 2862
rect 36109 2816 36179 2862
rect 36225 2816 36295 2862
rect 36341 2816 36411 2862
rect 36457 2816 36527 2862
rect 36573 2816 36643 2862
rect 36689 2816 36759 2862
rect 36805 2816 36875 2862
rect 36921 2816 36991 2862
rect 37037 2816 37107 2862
rect 37153 2816 37223 2862
rect 37269 2816 37339 2862
rect 37385 2816 37455 2862
rect 37501 2816 37571 2862
rect 37617 2816 37687 2862
rect 37733 2816 37803 2862
rect 37849 2816 37919 2862
rect 37965 2816 38035 2862
rect 38081 2816 38151 2862
rect 38197 2816 38267 2862
rect 38313 2816 38383 2862
rect 38429 2816 38499 2862
rect 38545 2816 38615 2862
rect 38661 2816 38731 2862
rect 38777 2816 38847 2862
rect 38893 2816 38963 2862
rect 39009 2816 39079 2862
rect 39125 2816 39195 2862
rect 39241 2816 39311 2862
rect 39357 2816 39427 2862
rect 39473 2816 39543 2862
rect 39589 2816 39659 2862
rect 39705 2816 39775 2862
rect 39821 2816 39891 2862
rect 39937 2816 40007 2862
rect 40053 2816 40123 2862
rect 40169 2816 40188 2862
rect 28620 2746 40188 2816
rect 28620 2700 28639 2746
rect 28685 2700 28755 2746
rect 28801 2700 28871 2746
rect 28917 2700 28987 2746
rect 29033 2700 29103 2746
rect 29149 2700 29219 2746
rect 29265 2700 29335 2746
rect 29381 2700 29451 2746
rect 29497 2700 29567 2746
rect 29613 2700 29683 2746
rect 29729 2700 29799 2746
rect 29845 2700 29915 2746
rect 29961 2700 30031 2746
rect 30077 2700 30147 2746
rect 30193 2700 30263 2746
rect 30309 2700 30379 2746
rect 30425 2700 30495 2746
rect 30541 2700 30611 2746
rect 30657 2700 30727 2746
rect 30773 2700 30843 2746
rect 30889 2700 30959 2746
rect 31005 2700 31075 2746
rect 31121 2700 31191 2746
rect 31237 2700 31307 2746
rect 31353 2700 31423 2746
rect 31469 2700 31539 2746
rect 31585 2700 31655 2746
rect 31701 2700 31771 2746
rect 31817 2700 31887 2746
rect 31933 2700 32003 2746
rect 32049 2700 32119 2746
rect 32165 2700 32235 2746
rect 32281 2700 32351 2746
rect 32397 2700 32467 2746
rect 32513 2700 32583 2746
rect 32629 2700 32699 2746
rect 32745 2700 32815 2746
rect 32861 2700 32931 2746
rect 32977 2700 33047 2746
rect 33093 2700 33163 2746
rect 33209 2700 33279 2746
rect 33325 2700 33395 2746
rect 33441 2700 33511 2746
rect 33557 2700 33627 2746
rect 33673 2700 33743 2746
rect 33789 2700 33859 2746
rect 33905 2700 33975 2746
rect 34021 2700 34091 2746
rect 34137 2700 34207 2746
rect 34253 2700 34323 2746
rect 34369 2700 34439 2746
rect 34485 2700 34555 2746
rect 34601 2700 34671 2746
rect 34717 2700 34787 2746
rect 34833 2700 34903 2746
rect 34949 2700 35019 2746
rect 35065 2700 35135 2746
rect 35181 2700 35251 2746
rect 35297 2700 35367 2746
rect 35413 2700 35483 2746
rect 35529 2700 35599 2746
rect 35645 2700 35715 2746
rect 35761 2700 35831 2746
rect 35877 2700 35947 2746
rect 35993 2700 36063 2746
rect 36109 2700 36179 2746
rect 36225 2700 36295 2746
rect 36341 2700 36411 2746
rect 36457 2700 36527 2746
rect 36573 2700 36643 2746
rect 36689 2700 36759 2746
rect 36805 2700 36875 2746
rect 36921 2700 36991 2746
rect 37037 2700 37107 2746
rect 37153 2700 37223 2746
rect 37269 2700 37339 2746
rect 37385 2700 37455 2746
rect 37501 2700 37571 2746
rect 37617 2700 37687 2746
rect 37733 2700 37803 2746
rect 37849 2700 37919 2746
rect 37965 2700 38035 2746
rect 38081 2700 38151 2746
rect 38197 2700 38267 2746
rect 38313 2700 38383 2746
rect 38429 2700 38499 2746
rect 38545 2700 38615 2746
rect 38661 2700 38731 2746
rect 38777 2700 38847 2746
rect 38893 2700 38963 2746
rect 39009 2700 39079 2746
rect 39125 2700 39195 2746
rect 39241 2700 39311 2746
rect 39357 2700 39427 2746
rect 39473 2700 39543 2746
rect 39589 2700 39659 2746
rect 39705 2700 39775 2746
rect 39821 2700 39891 2746
rect 39937 2700 40007 2746
rect 40053 2700 40123 2746
rect 40169 2700 40188 2746
rect 28620 2630 40188 2700
rect 28620 2584 28639 2630
rect 28685 2584 28755 2630
rect 28801 2584 28871 2630
rect 28917 2584 28987 2630
rect 29033 2584 29103 2630
rect 29149 2584 29219 2630
rect 29265 2584 29335 2630
rect 29381 2584 29451 2630
rect 29497 2584 29567 2630
rect 29613 2584 29683 2630
rect 29729 2584 29799 2630
rect 29845 2584 29915 2630
rect 29961 2584 30031 2630
rect 30077 2584 30147 2630
rect 30193 2584 30263 2630
rect 30309 2584 30379 2630
rect 30425 2584 30495 2630
rect 30541 2584 30611 2630
rect 30657 2584 30727 2630
rect 30773 2584 30843 2630
rect 30889 2584 30959 2630
rect 31005 2584 31075 2630
rect 31121 2584 31191 2630
rect 31237 2584 31307 2630
rect 31353 2584 31423 2630
rect 31469 2584 31539 2630
rect 31585 2584 31655 2630
rect 31701 2584 31771 2630
rect 31817 2584 31887 2630
rect 31933 2584 32003 2630
rect 32049 2584 32119 2630
rect 32165 2584 32235 2630
rect 32281 2584 32351 2630
rect 32397 2584 32467 2630
rect 32513 2584 32583 2630
rect 32629 2584 32699 2630
rect 32745 2584 32815 2630
rect 32861 2584 32931 2630
rect 32977 2584 33047 2630
rect 33093 2584 33163 2630
rect 33209 2584 33279 2630
rect 33325 2584 33395 2630
rect 33441 2584 33511 2630
rect 33557 2584 33627 2630
rect 33673 2584 33743 2630
rect 33789 2584 33859 2630
rect 33905 2584 33975 2630
rect 34021 2584 34091 2630
rect 34137 2584 34207 2630
rect 34253 2584 34323 2630
rect 34369 2584 34439 2630
rect 34485 2584 34555 2630
rect 34601 2584 34671 2630
rect 34717 2584 34787 2630
rect 34833 2584 34903 2630
rect 34949 2584 35019 2630
rect 35065 2584 35135 2630
rect 35181 2584 35251 2630
rect 35297 2584 35367 2630
rect 35413 2584 35483 2630
rect 35529 2584 35599 2630
rect 35645 2584 35715 2630
rect 35761 2584 35831 2630
rect 35877 2584 35947 2630
rect 35993 2584 36063 2630
rect 36109 2584 36179 2630
rect 36225 2584 36295 2630
rect 36341 2584 36411 2630
rect 36457 2584 36527 2630
rect 36573 2584 36643 2630
rect 36689 2584 36759 2630
rect 36805 2584 36875 2630
rect 36921 2584 36991 2630
rect 37037 2584 37107 2630
rect 37153 2584 37223 2630
rect 37269 2584 37339 2630
rect 37385 2584 37455 2630
rect 37501 2584 37571 2630
rect 37617 2584 37687 2630
rect 37733 2584 37803 2630
rect 37849 2584 37919 2630
rect 37965 2584 38035 2630
rect 38081 2584 38151 2630
rect 38197 2584 38267 2630
rect 38313 2584 38383 2630
rect 38429 2584 38499 2630
rect 38545 2584 38615 2630
rect 38661 2584 38731 2630
rect 38777 2584 38847 2630
rect 38893 2584 38963 2630
rect 39009 2584 39079 2630
rect 39125 2584 39195 2630
rect 39241 2584 39311 2630
rect 39357 2584 39427 2630
rect 39473 2584 39543 2630
rect 39589 2584 39659 2630
rect 39705 2584 39775 2630
rect 39821 2584 39891 2630
rect 39937 2584 40007 2630
rect 40053 2584 40123 2630
rect 40169 2584 40188 2630
rect 28620 2514 40188 2584
rect 28620 2468 28639 2514
rect 28685 2468 28755 2514
rect 28801 2468 28871 2514
rect 28917 2468 28987 2514
rect 29033 2468 29103 2514
rect 29149 2468 29219 2514
rect 29265 2468 29335 2514
rect 29381 2468 29451 2514
rect 29497 2468 29567 2514
rect 29613 2468 29683 2514
rect 29729 2468 29799 2514
rect 29845 2468 29915 2514
rect 29961 2468 30031 2514
rect 30077 2468 30147 2514
rect 30193 2468 30263 2514
rect 30309 2468 30379 2514
rect 30425 2468 30495 2514
rect 30541 2468 30611 2514
rect 30657 2468 30727 2514
rect 30773 2468 30843 2514
rect 30889 2468 30959 2514
rect 31005 2468 31075 2514
rect 31121 2468 31191 2514
rect 31237 2468 31307 2514
rect 31353 2468 31423 2514
rect 31469 2468 31539 2514
rect 31585 2468 31655 2514
rect 31701 2468 31771 2514
rect 31817 2468 31887 2514
rect 31933 2468 32003 2514
rect 32049 2468 32119 2514
rect 32165 2468 32235 2514
rect 32281 2468 32351 2514
rect 32397 2468 32467 2514
rect 32513 2468 32583 2514
rect 32629 2468 32699 2514
rect 32745 2468 32815 2514
rect 32861 2468 32931 2514
rect 32977 2468 33047 2514
rect 33093 2468 33163 2514
rect 33209 2468 33279 2514
rect 33325 2468 33395 2514
rect 33441 2468 33511 2514
rect 33557 2468 33627 2514
rect 33673 2468 33743 2514
rect 33789 2468 33859 2514
rect 33905 2468 33975 2514
rect 34021 2468 34091 2514
rect 34137 2468 34207 2514
rect 34253 2468 34323 2514
rect 34369 2468 34439 2514
rect 34485 2468 34555 2514
rect 34601 2468 34671 2514
rect 34717 2468 34787 2514
rect 34833 2468 34903 2514
rect 34949 2468 35019 2514
rect 35065 2468 35135 2514
rect 35181 2468 35251 2514
rect 35297 2468 35367 2514
rect 35413 2468 35483 2514
rect 35529 2468 35599 2514
rect 35645 2468 35715 2514
rect 35761 2468 35831 2514
rect 35877 2468 35947 2514
rect 35993 2468 36063 2514
rect 36109 2468 36179 2514
rect 36225 2468 36295 2514
rect 36341 2468 36411 2514
rect 36457 2468 36527 2514
rect 36573 2468 36643 2514
rect 36689 2468 36759 2514
rect 36805 2468 36875 2514
rect 36921 2468 36991 2514
rect 37037 2468 37107 2514
rect 37153 2468 37223 2514
rect 37269 2468 37339 2514
rect 37385 2468 37455 2514
rect 37501 2468 37571 2514
rect 37617 2468 37687 2514
rect 37733 2468 37803 2514
rect 37849 2468 37919 2514
rect 37965 2468 38035 2514
rect 38081 2468 38151 2514
rect 38197 2468 38267 2514
rect 38313 2468 38383 2514
rect 38429 2468 38499 2514
rect 38545 2468 38615 2514
rect 38661 2468 38731 2514
rect 38777 2468 38847 2514
rect 38893 2468 38963 2514
rect 39009 2468 39079 2514
rect 39125 2468 39195 2514
rect 39241 2468 39311 2514
rect 39357 2468 39427 2514
rect 39473 2468 39543 2514
rect 39589 2468 39659 2514
rect 39705 2468 39775 2514
rect 39821 2468 39891 2514
rect 39937 2468 40007 2514
rect 40053 2468 40123 2514
rect 40169 2468 40188 2514
rect 28620 2398 40188 2468
rect 28620 2352 28639 2398
rect 28685 2352 28755 2398
rect 28801 2352 28871 2398
rect 28917 2352 28987 2398
rect 29033 2352 29103 2398
rect 29149 2352 29219 2398
rect 29265 2352 29335 2398
rect 29381 2352 29451 2398
rect 29497 2352 29567 2398
rect 29613 2352 29683 2398
rect 29729 2352 29799 2398
rect 29845 2352 29915 2398
rect 29961 2352 30031 2398
rect 30077 2352 30147 2398
rect 30193 2352 30263 2398
rect 30309 2352 30379 2398
rect 30425 2352 30495 2398
rect 30541 2352 30611 2398
rect 30657 2352 30727 2398
rect 30773 2352 30843 2398
rect 30889 2352 30959 2398
rect 31005 2352 31075 2398
rect 31121 2352 31191 2398
rect 31237 2352 31307 2398
rect 31353 2352 31423 2398
rect 31469 2352 31539 2398
rect 31585 2352 31655 2398
rect 31701 2352 31771 2398
rect 31817 2352 31887 2398
rect 31933 2352 32003 2398
rect 32049 2352 32119 2398
rect 32165 2352 32235 2398
rect 32281 2352 32351 2398
rect 32397 2352 32467 2398
rect 32513 2352 32583 2398
rect 32629 2352 32699 2398
rect 32745 2352 32815 2398
rect 32861 2352 32931 2398
rect 32977 2352 33047 2398
rect 33093 2352 33163 2398
rect 33209 2352 33279 2398
rect 33325 2352 33395 2398
rect 33441 2352 33511 2398
rect 33557 2352 33627 2398
rect 33673 2352 33743 2398
rect 33789 2352 33859 2398
rect 33905 2352 33975 2398
rect 34021 2352 34091 2398
rect 34137 2352 34207 2398
rect 34253 2352 34323 2398
rect 34369 2352 34439 2398
rect 34485 2352 34555 2398
rect 34601 2352 34671 2398
rect 34717 2352 34787 2398
rect 34833 2352 34903 2398
rect 34949 2352 35019 2398
rect 35065 2352 35135 2398
rect 35181 2352 35251 2398
rect 35297 2352 35367 2398
rect 35413 2352 35483 2398
rect 35529 2352 35599 2398
rect 35645 2352 35715 2398
rect 35761 2352 35831 2398
rect 35877 2352 35947 2398
rect 35993 2352 36063 2398
rect 36109 2352 36179 2398
rect 36225 2352 36295 2398
rect 36341 2352 36411 2398
rect 36457 2352 36527 2398
rect 36573 2352 36643 2398
rect 36689 2352 36759 2398
rect 36805 2352 36875 2398
rect 36921 2352 36991 2398
rect 37037 2352 37107 2398
rect 37153 2352 37223 2398
rect 37269 2352 37339 2398
rect 37385 2352 37455 2398
rect 37501 2352 37571 2398
rect 37617 2352 37687 2398
rect 37733 2352 37803 2398
rect 37849 2352 37919 2398
rect 37965 2352 38035 2398
rect 38081 2352 38151 2398
rect 38197 2352 38267 2398
rect 38313 2352 38383 2398
rect 38429 2352 38499 2398
rect 38545 2352 38615 2398
rect 38661 2352 38731 2398
rect 38777 2352 38847 2398
rect 38893 2352 38963 2398
rect 39009 2352 39079 2398
rect 39125 2352 39195 2398
rect 39241 2352 39311 2398
rect 39357 2352 39427 2398
rect 39473 2352 39543 2398
rect 39589 2352 39659 2398
rect 39705 2352 39775 2398
rect 39821 2352 39891 2398
rect 39937 2352 40007 2398
rect 40053 2352 40123 2398
rect 40169 2352 40188 2398
rect 28620 2282 40188 2352
rect 28620 2236 28639 2282
rect 28685 2236 28755 2282
rect 28801 2236 28871 2282
rect 28917 2236 28987 2282
rect 29033 2236 29103 2282
rect 29149 2236 29219 2282
rect 29265 2236 29335 2282
rect 29381 2236 29451 2282
rect 29497 2236 29567 2282
rect 29613 2236 29683 2282
rect 29729 2236 29799 2282
rect 29845 2236 29915 2282
rect 29961 2236 30031 2282
rect 30077 2236 30147 2282
rect 30193 2236 30263 2282
rect 30309 2236 30379 2282
rect 30425 2236 30495 2282
rect 30541 2236 30611 2282
rect 30657 2236 30727 2282
rect 30773 2236 30843 2282
rect 30889 2236 30959 2282
rect 31005 2236 31075 2282
rect 31121 2236 31191 2282
rect 31237 2236 31307 2282
rect 31353 2236 31423 2282
rect 31469 2236 31539 2282
rect 31585 2236 31655 2282
rect 31701 2236 31771 2282
rect 31817 2236 31887 2282
rect 31933 2236 32003 2282
rect 32049 2236 32119 2282
rect 32165 2236 32235 2282
rect 32281 2236 32351 2282
rect 32397 2236 32467 2282
rect 32513 2236 32583 2282
rect 32629 2236 32699 2282
rect 32745 2236 32815 2282
rect 32861 2236 32931 2282
rect 32977 2236 33047 2282
rect 33093 2236 33163 2282
rect 33209 2236 33279 2282
rect 33325 2236 33395 2282
rect 33441 2236 33511 2282
rect 33557 2236 33627 2282
rect 33673 2236 33743 2282
rect 33789 2236 33859 2282
rect 33905 2236 33975 2282
rect 34021 2236 34091 2282
rect 34137 2236 34207 2282
rect 34253 2236 34323 2282
rect 34369 2236 34439 2282
rect 34485 2236 34555 2282
rect 34601 2236 34671 2282
rect 34717 2236 34787 2282
rect 34833 2236 34903 2282
rect 34949 2236 35019 2282
rect 35065 2236 35135 2282
rect 35181 2236 35251 2282
rect 35297 2236 35367 2282
rect 35413 2236 35483 2282
rect 35529 2236 35599 2282
rect 35645 2236 35715 2282
rect 35761 2236 35831 2282
rect 35877 2236 35947 2282
rect 35993 2236 36063 2282
rect 36109 2236 36179 2282
rect 36225 2236 36295 2282
rect 36341 2236 36411 2282
rect 36457 2236 36527 2282
rect 36573 2236 36643 2282
rect 36689 2236 36759 2282
rect 36805 2236 36875 2282
rect 36921 2236 36991 2282
rect 37037 2236 37107 2282
rect 37153 2236 37223 2282
rect 37269 2236 37339 2282
rect 37385 2236 37455 2282
rect 37501 2236 37571 2282
rect 37617 2236 37687 2282
rect 37733 2236 37803 2282
rect 37849 2236 37919 2282
rect 37965 2236 38035 2282
rect 38081 2236 38151 2282
rect 38197 2236 38267 2282
rect 38313 2236 38383 2282
rect 38429 2236 38499 2282
rect 38545 2236 38615 2282
rect 38661 2236 38731 2282
rect 38777 2236 38847 2282
rect 38893 2236 38963 2282
rect 39009 2236 39079 2282
rect 39125 2236 39195 2282
rect 39241 2236 39311 2282
rect 39357 2236 39427 2282
rect 39473 2236 39543 2282
rect 39589 2236 39659 2282
rect 39705 2236 39775 2282
rect 39821 2236 39891 2282
rect 39937 2236 40007 2282
rect 40053 2236 40123 2282
rect 40169 2236 40188 2282
rect 28620 2166 40188 2236
rect 28620 2120 28639 2166
rect 28685 2120 28755 2166
rect 28801 2120 28871 2166
rect 28917 2120 28987 2166
rect 29033 2120 29103 2166
rect 29149 2120 29219 2166
rect 29265 2120 29335 2166
rect 29381 2120 29451 2166
rect 29497 2120 29567 2166
rect 29613 2120 29683 2166
rect 29729 2120 29799 2166
rect 29845 2120 29915 2166
rect 29961 2120 30031 2166
rect 30077 2120 30147 2166
rect 30193 2120 30263 2166
rect 30309 2120 30379 2166
rect 30425 2120 30495 2166
rect 30541 2120 30611 2166
rect 30657 2120 30727 2166
rect 30773 2120 30843 2166
rect 30889 2120 30959 2166
rect 31005 2120 31075 2166
rect 31121 2120 31191 2166
rect 31237 2120 31307 2166
rect 31353 2120 31423 2166
rect 31469 2120 31539 2166
rect 31585 2120 31655 2166
rect 31701 2120 31771 2166
rect 31817 2120 31887 2166
rect 31933 2120 32003 2166
rect 32049 2120 32119 2166
rect 32165 2120 32235 2166
rect 32281 2120 32351 2166
rect 32397 2120 32467 2166
rect 32513 2120 32583 2166
rect 32629 2120 32699 2166
rect 32745 2120 32815 2166
rect 32861 2120 32931 2166
rect 32977 2120 33047 2166
rect 33093 2120 33163 2166
rect 33209 2120 33279 2166
rect 33325 2120 33395 2166
rect 33441 2120 33511 2166
rect 33557 2120 33627 2166
rect 33673 2120 33743 2166
rect 33789 2120 33859 2166
rect 33905 2120 33975 2166
rect 34021 2120 34091 2166
rect 34137 2120 34207 2166
rect 34253 2120 34323 2166
rect 34369 2120 34439 2166
rect 34485 2120 34555 2166
rect 34601 2120 34671 2166
rect 34717 2120 34787 2166
rect 34833 2120 34903 2166
rect 34949 2120 35019 2166
rect 35065 2120 35135 2166
rect 35181 2120 35251 2166
rect 35297 2120 35367 2166
rect 35413 2120 35483 2166
rect 35529 2120 35599 2166
rect 35645 2120 35715 2166
rect 35761 2120 35831 2166
rect 35877 2120 35947 2166
rect 35993 2120 36063 2166
rect 36109 2120 36179 2166
rect 36225 2120 36295 2166
rect 36341 2120 36411 2166
rect 36457 2120 36527 2166
rect 36573 2120 36643 2166
rect 36689 2120 36759 2166
rect 36805 2120 36875 2166
rect 36921 2120 36991 2166
rect 37037 2120 37107 2166
rect 37153 2120 37223 2166
rect 37269 2120 37339 2166
rect 37385 2120 37455 2166
rect 37501 2120 37571 2166
rect 37617 2120 37687 2166
rect 37733 2120 37803 2166
rect 37849 2120 37919 2166
rect 37965 2120 38035 2166
rect 38081 2120 38151 2166
rect 38197 2120 38267 2166
rect 38313 2120 38383 2166
rect 38429 2120 38499 2166
rect 38545 2120 38615 2166
rect 38661 2120 38731 2166
rect 38777 2120 38847 2166
rect 38893 2120 38963 2166
rect 39009 2120 39079 2166
rect 39125 2120 39195 2166
rect 39241 2120 39311 2166
rect 39357 2120 39427 2166
rect 39473 2120 39543 2166
rect 39589 2120 39659 2166
rect 39705 2120 39775 2166
rect 39821 2120 39891 2166
rect 39937 2120 40007 2166
rect 40053 2120 40123 2166
rect 40169 2120 40188 2166
rect 28620 2050 40188 2120
rect 28620 2004 28639 2050
rect 28685 2004 28755 2050
rect 28801 2004 28871 2050
rect 28917 2004 28987 2050
rect 29033 2004 29103 2050
rect 29149 2004 29219 2050
rect 29265 2004 29335 2050
rect 29381 2004 29451 2050
rect 29497 2004 29567 2050
rect 29613 2004 29683 2050
rect 29729 2004 29799 2050
rect 29845 2004 29915 2050
rect 29961 2004 30031 2050
rect 30077 2004 30147 2050
rect 30193 2004 30263 2050
rect 30309 2004 30379 2050
rect 30425 2004 30495 2050
rect 30541 2004 30611 2050
rect 30657 2004 30727 2050
rect 30773 2004 30843 2050
rect 30889 2004 30959 2050
rect 31005 2004 31075 2050
rect 31121 2004 31191 2050
rect 31237 2004 31307 2050
rect 31353 2004 31423 2050
rect 31469 2004 31539 2050
rect 31585 2004 31655 2050
rect 31701 2004 31771 2050
rect 31817 2004 31887 2050
rect 31933 2004 32003 2050
rect 32049 2004 32119 2050
rect 32165 2004 32235 2050
rect 32281 2004 32351 2050
rect 32397 2004 32467 2050
rect 32513 2004 32583 2050
rect 32629 2004 32699 2050
rect 32745 2004 32815 2050
rect 32861 2004 32931 2050
rect 32977 2004 33047 2050
rect 33093 2004 33163 2050
rect 33209 2004 33279 2050
rect 33325 2004 33395 2050
rect 33441 2004 33511 2050
rect 33557 2004 33627 2050
rect 33673 2004 33743 2050
rect 33789 2004 33859 2050
rect 33905 2004 33975 2050
rect 34021 2004 34091 2050
rect 34137 2004 34207 2050
rect 34253 2004 34323 2050
rect 34369 2004 34439 2050
rect 34485 2004 34555 2050
rect 34601 2004 34671 2050
rect 34717 2004 34787 2050
rect 34833 2004 34903 2050
rect 34949 2004 35019 2050
rect 35065 2004 35135 2050
rect 35181 2004 35251 2050
rect 35297 2004 35367 2050
rect 35413 2004 35483 2050
rect 35529 2004 35599 2050
rect 35645 2004 35715 2050
rect 35761 2004 35831 2050
rect 35877 2004 35947 2050
rect 35993 2004 36063 2050
rect 36109 2004 36179 2050
rect 36225 2004 36295 2050
rect 36341 2004 36411 2050
rect 36457 2004 36527 2050
rect 36573 2004 36643 2050
rect 36689 2004 36759 2050
rect 36805 2004 36875 2050
rect 36921 2004 36991 2050
rect 37037 2004 37107 2050
rect 37153 2004 37223 2050
rect 37269 2004 37339 2050
rect 37385 2004 37455 2050
rect 37501 2004 37571 2050
rect 37617 2004 37687 2050
rect 37733 2004 37803 2050
rect 37849 2004 37919 2050
rect 37965 2004 38035 2050
rect 38081 2004 38151 2050
rect 38197 2004 38267 2050
rect 38313 2004 38383 2050
rect 38429 2004 38499 2050
rect 38545 2004 38615 2050
rect 38661 2004 38731 2050
rect 38777 2004 38847 2050
rect 38893 2004 38963 2050
rect 39009 2004 39079 2050
rect 39125 2004 39195 2050
rect 39241 2004 39311 2050
rect 39357 2004 39427 2050
rect 39473 2004 39543 2050
rect 39589 2004 39659 2050
rect 39705 2004 39775 2050
rect 39821 2004 39891 2050
rect 39937 2004 40007 2050
rect 40053 2004 40123 2050
rect 40169 2004 40188 2050
rect 28620 1934 40188 2004
rect 28620 1888 28639 1934
rect 28685 1888 28755 1934
rect 28801 1888 28871 1934
rect 28917 1888 28987 1934
rect 29033 1888 29103 1934
rect 29149 1888 29219 1934
rect 29265 1888 29335 1934
rect 29381 1888 29451 1934
rect 29497 1888 29567 1934
rect 29613 1888 29683 1934
rect 29729 1888 29799 1934
rect 29845 1888 29915 1934
rect 29961 1888 30031 1934
rect 30077 1888 30147 1934
rect 30193 1888 30263 1934
rect 30309 1888 30379 1934
rect 30425 1888 30495 1934
rect 30541 1888 30611 1934
rect 30657 1888 30727 1934
rect 30773 1888 30843 1934
rect 30889 1888 30959 1934
rect 31005 1888 31075 1934
rect 31121 1888 31191 1934
rect 31237 1888 31307 1934
rect 31353 1888 31423 1934
rect 31469 1888 31539 1934
rect 31585 1888 31655 1934
rect 31701 1888 31771 1934
rect 31817 1888 31887 1934
rect 31933 1888 32003 1934
rect 32049 1888 32119 1934
rect 32165 1888 32235 1934
rect 32281 1888 32351 1934
rect 32397 1888 32467 1934
rect 32513 1888 32583 1934
rect 32629 1888 32699 1934
rect 32745 1888 32815 1934
rect 32861 1888 32931 1934
rect 32977 1888 33047 1934
rect 33093 1888 33163 1934
rect 33209 1888 33279 1934
rect 33325 1888 33395 1934
rect 33441 1888 33511 1934
rect 33557 1888 33627 1934
rect 33673 1888 33743 1934
rect 33789 1888 33859 1934
rect 33905 1888 33975 1934
rect 34021 1888 34091 1934
rect 34137 1888 34207 1934
rect 34253 1888 34323 1934
rect 34369 1888 34439 1934
rect 34485 1888 34555 1934
rect 34601 1888 34671 1934
rect 34717 1888 34787 1934
rect 34833 1888 34903 1934
rect 34949 1888 35019 1934
rect 35065 1888 35135 1934
rect 35181 1888 35251 1934
rect 35297 1888 35367 1934
rect 35413 1888 35483 1934
rect 35529 1888 35599 1934
rect 35645 1888 35715 1934
rect 35761 1888 35831 1934
rect 35877 1888 35947 1934
rect 35993 1888 36063 1934
rect 36109 1888 36179 1934
rect 36225 1888 36295 1934
rect 36341 1888 36411 1934
rect 36457 1888 36527 1934
rect 36573 1888 36643 1934
rect 36689 1888 36759 1934
rect 36805 1888 36875 1934
rect 36921 1888 36991 1934
rect 37037 1888 37107 1934
rect 37153 1888 37223 1934
rect 37269 1888 37339 1934
rect 37385 1888 37455 1934
rect 37501 1888 37571 1934
rect 37617 1888 37687 1934
rect 37733 1888 37803 1934
rect 37849 1888 37919 1934
rect 37965 1888 38035 1934
rect 38081 1888 38151 1934
rect 38197 1888 38267 1934
rect 38313 1888 38383 1934
rect 38429 1888 38499 1934
rect 38545 1888 38615 1934
rect 38661 1888 38731 1934
rect 38777 1888 38847 1934
rect 38893 1888 38963 1934
rect 39009 1888 39079 1934
rect 39125 1888 39195 1934
rect 39241 1888 39311 1934
rect 39357 1888 39427 1934
rect 39473 1888 39543 1934
rect 39589 1888 39659 1934
rect 39705 1888 39775 1934
rect 39821 1888 39891 1934
rect 39937 1888 40007 1934
rect 40053 1888 40123 1934
rect 40169 1888 40188 1934
rect 28620 1818 40188 1888
rect 28620 1772 28639 1818
rect 28685 1772 28755 1818
rect 28801 1772 28871 1818
rect 28917 1772 28987 1818
rect 29033 1772 29103 1818
rect 29149 1772 29219 1818
rect 29265 1772 29335 1818
rect 29381 1772 29451 1818
rect 29497 1772 29567 1818
rect 29613 1772 29683 1818
rect 29729 1772 29799 1818
rect 29845 1772 29915 1818
rect 29961 1772 30031 1818
rect 30077 1772 30147 1818
rect 30193 1772 30263 1818
rect 30309 1772 30379 1818
rect 30425 1772 30495 1818
rect 30541 1772 30611 1818
rect 30657 1772 30727 1818
rect 30773 1772 30843 1818
rect 30889 1772 30959 1818
rect 31005 1772 31075 1818
rect 31121 1772 31191 1818
rect 31237 1772 31307 1818
rect 31353 1772 31423 1818
rect 31469 1772 31539 1818
rect 31585 1772 31655 1818
rect 31701 1772 31771 1818
rect 31817 1772 31887 1818
rect 31933 1772 32003 1818
rect 32049 1772 32119 1818
rect 32165 1772 32235 1818
rect 32281 1772 32351 1818
rect 32397 1772 32467 1818
rect 32513 1772 32583 1818
rect 32629 1772 32699 1818
rect 32745 1772 32815 1818
rect 32861 1772 32931 1818
rect 32977 1772 33047 1818
rect 33093 1772 33163 1818
rect 33209 1772 33279 1818
rect 33325 1772 33395 1818
rect 33441 1772 33511 1818
rect 33557 1772 33627 1818
rect 33673 1772 33743 1818
rect 33789 1772 33859 1818
rect 33905 1772 33975 1818
rect 34021 1772 34091 1818
rect 34137 1772 34207 1818
rect 34253 1772 34323 1818
rect 34369 1772 34439 1818
rect 34485 1772 34555 1818
rect 34601 1772 34671 1818
rect 34717 1772 34787 1818
rect 34833 1772 34903 1818
rect 34949 1772 35019 1818
rect 35065 1772 35135 1818
rect 35181 1772 35251 1818
rect 35297 1772 35367 1818
rect 35413 1772 35483 1818
rect 35529 1772 35599 1818
rect 35645 1772 35715 1818
rect 35761 1772 35831 1818
rect 35877 1772 35947 1818
rect 35993 1772 36063 1818
rect 36109 1772 36179 1818
rect 36225 1772 36295 1818
rect 36341 1772 36411 1818
rect 36457 1772 36527 1818
rect 36573 1772 36643 1818
rect 36689 1772 36759 1818
rect 36805 1772 36875 1818
rect 36921 1772 36991 1818
rect 37037 1772 37107 1818
rect 37153 1772 37223 1818
rect 37269 1772 37339 1818
rect 37385 1772 37455 1818
rect 37501 1772 37571 1818
rect 37617 1772 37687 1818
rect 37733 1772 37803 1818
rect 37849 1772 37919 1818
rect 37965 1772 38035 1818
rect 38081 1772 38151 1818
rect 38197 1772 38267 1818
rect 38313 1772 38383 1818
rect 38429 1772 38499 1818
rect 38545 1772 38615 1818
rect 38661 1772 38731 1818
rect 38777 1772 38847 1818
rect 38893 1772 38963 1818
rect 39009 1772 39079 1818
rect 39125 1772 39195 1818
rect 39241 1772 39311 1818
rect 39357 1772 39427 1818
rect 39473 1772 39543 1818
rect 39589 1772 39659 1818
rect 39705 1772 39775 1818
rect 39821 1772 39891 1818
rect 39937 1772 40007 1818
rect 40053 1772 40123 1818
rect 40169 1772 40188 1818
rect 28620 1702 40188 1772
rect 28620 1656 28639 1702
rect 28685 1656 28755 1702
rect 28801 1656 28871 1702
rect 28917 1656 28987 1702
rect 29033 1656 29103 1702
rect 29149 1656 29219 1702
rect 29265 1656 29335 1702
rect 29381 1656 29451 1702
rect 29497 1656 29567 1702
rect 29613 1656 29683 1702
rect 29729 1656 29799 1702
rect 29845 1656 29915 1702
rect 29961 1656 30031 1702
rect 30077 1656 30147 1702
rect 30193 1656 30263 1702
rect 30309 1656 30379 1702
rect 30425 1656 30495 1702
rect 30541 1656 30611 1702
rect 30657 1656 30727 1702
rect 30773 1656 30843 1702
rect 30889 1656 30959 1702
rect 31005 1656 31075 1702
rect 31121 1656 31191 1702
rect 31237 1656 31307 1702
rect 31353 1656 31423 1702
rect 31469 1656 31539 1702
rect 31585 1656 31655 1702
rect 31701 1656 31771 1702
rect 31817 1656 31887 1702
rect 31933 1656 32003 1702
rect 32049 1656 32119 1702
rect 32165 1656 32235 1702
rect 32281 1656 32351 1702
rect 32397 1656 32467 1702
rect 32513 1656 32583 1702
rect 32629 1656 32699 1702
rect 32745 1656 32815 1702
rect 32861 1656 32931 1702
rect 32977 1656 33047 1702
rect 33093 1656 33163 1702
rect 33209 1656 33279 1702
rect 33325 1656 33395 1702
rect 33441 1656 33511 1702
rect 33557 1656 33627 1702
rect 33673 1656 33743 1702
rect 33789 1656 33859 1702
rect 33905 1656 33975 1702
rect 34021 1656 34091 1702
rect 34137 1656 34207 1702
rect 34253 1656 34323 1702
rect 34369 1656 34439 1702
rect 34485 1656 34555 1702
rect 34601 1656 34671 1702
rect 34717 1656 34787 1702
rect 34833 1656 34903 1702
rect 34949 1656 35019 1702
rect 35065 1656 35135 1702
rect 35181 1656 35251 1702
rect 35297 1656 35367 1702
rect 35413 1656 35483 1702
rect 35529 1656 35599 1702
rect 35645 1656 35715 1702
rect 35761 1656 35831 1702
rect 35877 1656 35947 1702
rect 35993 1656 36063 1702
rect 36109 1656 36179 1702
rect 36225 1656 36295 1702
rect 36341 1656 36411 1702
rect 36457 1656 36527 1702
rect 36573 1656 36643 1702
rect 36689 1656 36759 1702
rect 36805 1656 36875 1702
rect 36921 1656 36991 1702
rect 37037 1656 37107 1702
rect 37153 1656 37223 1702
rect 37269 1656 37339 1702
rect 37385 1656 37455 1702
rect 37501 1656 37571 1702
rect 37617 1656 37687 1702
rect 37733 1656 37803 1702
rect 37849 1656 37919 1702
rect 37965 1656 38035 1702
rect 38081 1656 38151 1702
rect 38197 1656 38267 1702
rect 38313 1656 38383 1702
rect 38429 1656 38499 1702
rect 38545 1656 38615 1702
rect 38661 1656 38731 1702
rect 38777 1656 38847 1702
rect 38893 1656 38963 1702
rect 39009 1656 39079 1702
rect 39125 1656 39195 1702
rect 39241 1656 39311 1702
rect 39357 1656 39427 1702
rect 39473 1656 39543 1702
rect 39589 1656 39659 1702
rect 39705 1656 39775 1702
rect 39821 1656 39891 1702
rect 39937 1656 40007 1702
rect 40053 1656 40123 1702
rect 40169 1656 40188 1702
rect 28620 1637 40188 1656
rect 50826 3906 56594 3925
rect 50826 3860 50845 3906
rect 50891 3860 50961 3906
rect 51007 3860 51077 3906
rect 51123 3860 51193 3906
rect 51239 3860 51309 3906
rect 51355 3860 51425 3906
rect 51471 3860 51541 3906
rect 51587 3860 51657 3906
rect 51703 3860 51773 3906
rect 51819 3860 51889 3906
rect 51935 3860 52005 3906
rect 52051 3860 52121 3906
rect 52167 3860 52237 3906
rect 52283 3860 52353 3906
rect 52399 3860 52469 3906
rect 52515 3860 52585 3906
rect 52631 3860 52701 3906
rect 52747 3860 52817 3906
rect 52863 3860 52933 3906
rect 52979 3860 53049 3906
rect 53095 3860 53165 3906
rect 53211 3860 53281 3906
rect 53327 3860 53397 3906
rect 53443 3860 53513 3906
rect 53559 3860 53629 3906
rect 53675 3860 53745 3906
rect 53791 3860 53861 3906
rect 53907 3860 53977 3906
rect 54023 3860 54093 3906
rect 54139 3860 54209 3906
rect 54255 3860 54325 3906
rect 54371 3860 54441 3906
rect 54487 3860 54557 3906
rect 54603 3860 54673 3906
rect 54719 3860 54789 3906
rect 54835 3860 54905 3906
rect 54951 3860 55021 3906
rect 55067 3860 55137 3906
rect 55183 3860 55253 3906
rect 55299 3860 55369 3906
rect 55415 3860 55485 3906
rect 55531 3860 55601 3906
rect 55647 3860 55717 3906
rect 55763 3860 55833 3906
rect 55879 3860 55949 3906
rect 55995 3860 56065 3906
rect 56111 3860 56181 3906
rect 56227 3860 56297 3906
rect 56343 3860 56413 3906
rect 56459 3860 56529 3906
rect 56575 3860 56594 3906
rect 50826 3790 56594 3860
rect 50826 3744 50845 3790
rect 50891 3744 50961 3790
rect 51007 3744 51077 3790
rect 51123 3744 51193 3790
rect 51239 3744 51309 3790
rect 51355 3744 51425 3790
rect 51471 3744 51541 3790
rect 51587 3744 51657 3790
rect 51703 3744 51773 3790
rect 51819 3744 51889 3790
rect 51935 3744 52005 3790
rect 52051 3744 52121 3790
rect 52167 3744 52237 3790
rect 52283 3744 52353 3790
rect 52399 3744 52469 3790
rect 52515 3744 52585 3790
rect 52631 3744 52701 3790
rect 52747 3744 52817 3790
rect 52863 3744 52933 3790
rect 52979 3744 53049 3790
rect 53095 3744 53165 3790
rect 53211 3744 53281 3790
rect 53327 3744 53397 3790
rect 53443 3744 53513 3790
rect 53559 3744 53629 3790
rect 53675 3744 53745 3790
rect 53791 3744 53861 3790
rect 53907 3744 53977 3790
rect 54023 3744 54093 3790
rect 54139 3744 54209 3790
rect 54255 3744 54325 3790
rect 54371 3744 54441 3790
rect 54487 3744 54557 3790
rect 54603 3744 54673 3790
rect 54719 3744 54789 3790
rect 54835 3744 54905 3790
rect 54951 3744 55021 3790
rect 55067 3744 55137 3790
rect 55183 3744 55253 3790
rect 55299 3744 55369 3790
rect 55415 3744 55485 3790
rect 55531 3744 55601 3790
rect 55647 3744 55717 3790
rect 55763 3744 55833 3790
rect 55879 3744 55949 3790
rect 55995 3744 56065 3790
rect 56111 3744 56181 3790
rect 56227 3744 56297 3790
rect 56343 3744 56413 3790
rect 56459 3744 56529 3790
rect 56575 3744 56594 3790
rect 50826 3674 56594 3744
rect 50826 3628 50845 3674
rect 50891 3628 50961 3674
rect 51007 3628 51077 3674
rect 51123 3628 51193 3674
rect 51239 3628 51309 3674
rect 51355 3628 51425 3674
rect 51471 3628 51541 3674
rect 51587 3628 51657 3674
rect 51703 3628 51773 3674
rect 51819 3628 51889 3674
rect 51935 3628 52005 3674
rect 52051 3628 52121 3674
rect 52167 3628 52237 3674
rect 52283 3628 52353 3674
rect 52399 3628 52469 3674
rect 52515 3628 52585 3674
rect 52631 3628 52701 3674
rect 52747 3628 52817 3674
rect 52863 3628 52933 3674
rect 52979 3628 53049 3674
rect 53095 3628 53165 3674
rect 53211 3628 53281 3674
rect 53327 3628 53397 3674
rect 53443 3628 53513 3674
rect 53559 3628 53629 3674
rect 53675 3628 53745 3674
rect 53791 3628 53861 3674
rect 53907 3628 53977 3674
rect 54023 3628 54093 3674
rect 54139 3628 54209 3674
rect 54255 3628 54325 3674
rect 54371 3628 54441 3674
rect 54487 3628 54557 3674
rect 54603 3628 54673 3674
rect 54719 3628 54789 3674
rect 54835 3628 54905 3674
rect 54951 3628 55021 3674
rect 55067 3628 55137 3674
rect 55183 3628 55253 3674
rect 55299 3628 55369 3674
rect 55415 3628 55485 3674
rect 55531 3628 55601 3674
rect 55647 3628 55717 3674
rect 55763 3628 55833 3674
rect 55879 3628 55949 3674
rect 55995 3628 56065 3674
rect 56111 3628 56181 3674
rect 56227 3628 56297 3674
rect 56343 3628 56413 3674
rect 56459 3628 56529 3674
rect 56575 3628 56594 3674
rect 50826 3558 56594 3628
rect 50826 3512 50845 3558
rect 50891 3512 50961 3558
rect 51007 3512 51077 3558
rect 51123 3512 51193 3558
rect 51239 3512 51309 3558
rect 51355 3512 51425 3558
rect 51471 3512 51541 3558
rect 51587 3512 51657 3558
rect 51703 3512 51773 3558
rect 51819 3512 51889 3558
rect 51935 3512 52005 3558
rect 52051 3512 52121 3558
rect 52167 3512 52237 3558
rect 52283 3512 52353 3558
rect 52399 3512 52469 3558
rect 52515 3512 52585 3558
rect 52631 3512 52701 3558
rect 52747 3512 52817 3558
rect 52863 3512 52933 3558
rect 52979 3512 53049 3558
rect 53095 3512 53165 3558
rect 53211 3512 53281 3558
rect 53327 3512 53397 3558
rect 53443 3512 53513 3558
rect 53559 3512 53629 3558
rect 53675 3512 53745 3558
rect 53791 3512 53861 3558
rect 53907 3512 53977 3558
rect 54023 3512 54093 3558
rect 54139 3512 54209 3558
rect 54255 3512 54325 3558
rect 54371 3512 54441 3558
rect 54487 3512 54557 3558
rect 54603 3512 54673 3558
rect 54719 3512 54789 3558
rect 54835 3512 54905 3558
rect 54951 3512 55021 3558
rect 55067 3512 55137 3558
rect 55183 3512 55253 3558
rect 55299 3512 55369 3558
rect 55415 3512 55485 3558
rect 55531 3512 55601 3558
rect 55647 3512 55717 3558
rect 55763 3512 55833 3558
rect 55879 3512 55949 3558
rect 55995 3512 56065 3558
rect 56111 3512 56181 3558
rect 56227 3512 56297 3558
rect 56343 3512 56413 3558
rect 56459 3512 56529 3558
rect 56575 3512 56594 3558
rect 50826 3442 56594 3512
rect 50826 3396 50845 3442
rect 50891 3396 50961 3442
rect 51007 3396 51077 3442
rect 51123 3396 51193 3442
rect 51239 3396 51309 3442
rect 51355 3396 51425 3442
rect 51471 3396 51541 3442
rect 51587 3396 51657 3442
rect 51703 3396 51773 3442
rect 51819 3396 51889 3442
rect 51935 3396 52005 3442
rect 52051 3396 52121 3442
rect 52167 3396 52237 3442
rect 52283 3396 52353 3442
rect 52399 3396 52469 3442
rect 52515 3396 52585 3442
rect 52631 3396 52701 3442
rect 52747 3396 52817 3442
rect 52863 3396 52933 3442
rect 52979 3396 53049 3442
rect 53095 3396 53165 3442
rect 53211 3396 53281 3442
rect 53327 3396 53397 3442
rect 53443 3396 53513 3442
rect 53559 3396 53629 3442
rect 53675 3396 53745 3442
rect 53791 3396 53861 3442
rect 53907 3396 53977 3442
rect 54023 3396 54093 3442
rect 54139 3396 54209 3442
rect 54255 3396 54325 3442
rect 54371 3396 54441 3442
rect 54487 3396 54557 3442
rect 54603 3396 54673 3442
rect 54719 3396 54789 3442
rect 54835 3396 54905 3442
rect 54951 3396 55021 3442
rect 55067 3396 55137 3442
rect 55183 3396 55253 3442
rect 55299 3396 55369 3442
rect 55415 3396 55485 3442
rect 55531 3396 55601 3442
rect 55647 3396 55717 3442
rect 55763 3396 55833 3442
rect 55879 3396 55949 3442
rect 55995 3396 56065 3442
rect 56111 3396 56181 3442
rect 56227 3396 56297 3442
rect 56343 3396 56413 3442
rect 56459 3396 56529 3442
rect 56575 3396 56594 3442
rect 50826 3326 56594 3396
rect 50826 3280 50845 3326
rect 50891 3280 50961 3326
rect 51007 3280 51077 3326
rect 51123 3280 51193 3326
rect 51239 3280 51309 3326
rect 51355 3280 51425 3326
rect 51471 3280 51541 3326
rect 51587 3280 51657 3326
rect 51703 3280 51773 3326
rect 51819 3280 51889 3326
rect 51935 3280 52005 3326
rect 52051 3280 52121 3326
rect 52167 3280 52237 3326
rect 52283 3280 52353 3326
rect 52399 3280 52469 3326
rect 52515 3280 52585 3326
rect 52631 3280 52701 3326
rect 52747 3280 52817 3326
rect 52863 3280 52933 3326
rect 52979 3280 53049 3326
rect 53095 3280 53165 3326
rect 53211 3280 53281 3326
rect 53327 3280 53397 3326
rect 53443 3280 53513 3326
rect 53559 3280 53629 3326
rect 53675 3280 53745 3326
rect 53791 3280 53861 3326
rect 53907 3280 53977 3326
rect 54023 3280 54093 3326
rect 54139 3280 54209 3326
rect 54255 3280 54325 3326
rect 54371 3280 54441 3326
rect 54487 3280 54557 3326
rect 54603 3280 54673 3326
rect 54719 3280 54789 3326
rect 54835 3280 54905 3326
rect 54951 3280 55021 3326
rect 55067 3280 55137 3326
rect 55183 3280 55253 3326
rect 55299 3280 55369 3326
rect 55415 3280 55485 3326
rect 55531 3280 55601 3326
rect 55647 3280 55717 3326
rect 55763 3280 55833 3326
rect 55879 3280 55949 3326
rect 55995 3280 56065 3326
rect 56111 3280 56181 3326
rect 56227 3280 56297 3326
rect 56343 3280 56413 3326
rect 56459 3280 56529 3326
rect 56575 3280 56594 3326
rect 50826 3210 56594 3280
rect 50826 3164 50845 3210
rect 50891 3164 50961 3210
rect 51007 3164 51077 3210
rect 51123 3164 51193 3210
rect 51239 3164 51309 3210
rect 51355 3164 51425 3210
rect 51471 3164 51541 3210
rect 51587 3164 51657 3210
rect 51703 3164 51773 3210
rect 51819 3164 51889 3210
rect 51935 3164 52005 3210
rect 52051 3164 52121 3210
rect 52167 3164 52237 3210
rect 52283 3164 52353 3210
rect 52399 3164 52469 3210
rect 52515 3164 52585 3210
rect 52631 3164 52701 3210
rect 52747 3164 52817 3210
rect 52863 3164 52933 3210
rect 52979 3164 53049 3210
rect 53095 3164 53165 3210
rect 53211 3164 53281 3210
rect 53327 3164 53397 3210
rect 53443 3164 53513 3210
rect 53559 3164 53629 3210
rect 53675 3164 53745 3210
rect 53791 3164 53861 3210
rect 53907 3164 53977 3210
rect 54023 3164 54093 3210
rect 54139 3164 54209 3210
rect 54255 3164 54325 3210
rect 54371 3164 54441 3210
rect 54487 3164 54557 3210
rect 54603 3164 54673 3210
rect 54719 3164 54789 3210
rect 54835 3164 54905 3210
rect 54951 3164 55021 3210
rect 55067 3164 55137 3210
rect 55183 3164 55253 3210
rect 55299 3164 55369 3210
rect 55415 3164 55485 3210
rect 55531 3164 55601 3210
rect 55647 3164 55717 3210
rect 55763 3164 55833 3210
rect 55879 3164 55949 3210
rect 55995 3164 56065 3210
rect 56111 3164 56181 3210
rect 56227 3164 56297 3210
rect 56343 3164 56413 3210
rect 56459 3164 56529 3210
rect 56575 3164 56594 3210
rect 50826 3094 56594 3164
rect 50826 3048 50845 3094
rect 50891 3048 50961 3094
rect 51007 3048 51077 3094
rect 51123 3048 51193 3094
rect 51239 3048 51309 3094
rect 51355 3048 51425 3094
rect 51471 3048 51541 3094
rect 51587 3048 51657 3094
rect 51703 3048 51773 3094
rect 51819 3048 51889 3094
rect 51935 3048 52005 3094
rect 52051 3048 52121 3094
rect 52167 3048 52237 3094
rect 52283 3048 52353 3094
rect 52399 3048 52469 3094
rect 52515 3048 52585 3094
rect 52631 3048 52701 3094
rect 52747 3048 52817 3094
rect 52863 3048 52933 3094
rect 52979 3048 53049 3094
rect 53095 3048 53165 3094
rect 53211 3048 53281 3094
rect 53327 3048 53397 3094
rect 53443 3048 53513 3094
rect 53559 3048 53629 3094
rect 53675 3048 53745 3094
rect 53791 3048 53861 3094
rect 53907 3048 53977 3094
rect 54023 3048 54093 3094
rect 54139 3048 54209 3094
rect 54255 3048 54325 3094
rect 54371 3048 54441 3094
rect 54487 3048 54557 3094
rect 54603 3048 54673 3094
rect 54719 3048 54789 3094
rect 54835 3048 54905 3094
rect 54951 3048 55021 3094
rect 55067 3048 55137 3094
rect 55183 3048 55253 3094
rect 55299 3048 55369 3094
rect 55415 3048 55485 3094
rect 55531 3048 55601 3094
rect 55647 3048 55717 3094
rect 55763 3048 55833 3094
rect 55879 3048 55949 3094
rect 55995 3048 56065 3094
rect 56111 3048 56181 3094
rect 56227 3048 56297 3094
rect 56343 3048 56413 3094
rect 56459 3048 56529 3094
rect 56575 3048 56594 3094
rect 50826 2978 56594 3048
rect 50826 2932 50845 2978
rect 50891 2932 50961 2978
rect 51007 2932 51077 2978
rect 51123 2932 51193 2978
rect 51239 2932 51309 2978
rect 51355 2932 51425 2978
rect 51471 2932 51541 2978
rect 51587 2932 51657 2978
rect 51703 2932 51773 2978
rect 51819 2932 51889 2978
rect 51935 2932 52005 2978
rect 52051 2932 52121 2978
rect 52167 2932 52237 2978
rect 52283 2932 52353 2978
rect 52399 2932 52469 2978
rect 52515 2932 52585 2978
rect 52631 2932 52701 2978
rect 52747 2932 52817 2978
rect 52863 2932 52933 2978
rect 52979 2932 53049 2978
rect 53095 2932 53165 2978
rect 53211 2932 53281 2978
rect 53327 2932 53397 2978
rect 53443 2932 53513 2978
rect 53559 2932 53629 2978
rect 53675 2932 53745 2978
rect 53791 2932 53861 2978
rect 53907 2932 53977 2978
rect 54023 2932 54093 2978
rect 54139 2932 54209 2978
rect 54255 2932 54325 2978
rect 54371 2932 54441 2978
rect 54487 2932 54557 2978
rect 54603 2932 54673 2978
rect 54719 2932 54789 2978
rect 54835 2932 54905 2978
rect 54951 2932 55021 2978
rect 55067 2932 55137 2978
rect 55183 2932 55253 2978
rect 55299 2932 55369 2978
rect 55415 2932 55485 2978
rect 55531 2932 55601 2978
rect 55647 2932 55717 2978
rect 55763 2932 55833 2978
rect 55879 2932 55949 2978
rect 55995 2932 56065 2978
rect 56111 2932 56181 2978
rect 56227 2932 56297 2978
rect 56343 2932 56413 2978
rect 56459 2932 56529 2978
rect 56575 2932 56594 2978
rect 50826 2862 56594 2932
rect 50826 2816 50845 2862
rect 50891 2816 50961 2862
rect 51007 2816 51077 2862
rect 51123 2816 51193 2862
rect 51239 2816 51309 2862
rect 51355 2816 51425 2862
rect 51471 2816 51541 2862
rect 51587 2816 51657 2862
rect 51703 2816 51773 2862
rect 51819 2816 51889 2862
rect 51935 2816 52005 2862
rect 52051 2816 52121 2862
rect 52167 2816 52237 2862
rect 52283 2816 52353 2862
rect 52399 2816 52469 2862
rect 52515 2816 52585 2862
rect 52631 2816 52701 2862
rect 52747 2816 52817 2862
rect 52863 2816 52933 2862
rect 52979 2816 53049 2862
rect 53095 2816 53165 2862
rect 53211 2816 53281 2862
rect 53327 2816 53397 2862
rect 53443 2816 53513 2862
rect 53559 2816 53629 2862
rect 53675 2816 53745 2862
rect 53791 2816 53861 2862
rect 53907 2816 53977 2862
rect 54023 2816 54093 2862
rect 54139 2816 54209 2862
rect 54255 2816 54325 2862
rect 54371 2816 54441 2862
rect 54487 2816 54557 2862
rect 54603 2816 54673 2862
rect 54719 2816 54789 2862
rect 54835 2816 54905 2862
rect 54951 2816 55021 2862
rect 55067 2816 55137 2862
rect 55183 2816 55253 2862
rect 55299 2816 55369 2862
rect 55415 2816 55485 2862
rect 55531 2816 55601 2862
rect 55647 2816 55717 2862
rect 55763 2816 55833 2862
rect 55879 2816 55949 2862
rect 55995 2816 56065 2862
rect 56111 2816 56181 2862
rect 56227 2816 56297 2862
rect 56343 2816 56413 2862
rect 56459 2816 56529 2862
rect 56575 2816 56594 2862
rect 50826 2746 56594 2816
rect 50826 2700 50845 2746
rect 50891 2700 50961 2746
rect 51007 2700 51077 2746
rect 51123 2700 51193 2746
rect 51239 2700 51309 2746
rect 51355 2700 51425 2746
rect 51471 2700 51541 2746
rect 51587 2700 51657 2746
rect 51703 2700 51773 2746
rect 51819 2700 51889 2746
rect 51935 2700 52005 2746
rect 52051 2700 52121 2746
rect 52167 2700 52237 2746
rect 52283 2700 52353 2746
rect 52399 2700 52469 2746
rect 52515 2700 52585 2746
rect 52631 2700 52701 2746
rect 52747 2700 52817 2746
rect 52863 2700 52933 2746
rect 52979 2700 53049 2746
rect 53095 2700 53165 2746
rect 53211 2700 53281 2746
rect 53327 2700 53397 2746
rect 53443 2700 53513 2746
rect 53559 2700 53629 2746
rect 53675 2700 53745 2746
rect 53791 2700 53861 2746
rect 53907 2700 53977 2746
rect 54023 2700 54093 2746
rect 54139 2700 54209 2746
rect 54255 2700 54325 2746
rect 54371 2700 54441 2746
rect 54487 2700 54557 2746
rect 54603 2700 54673 2746
rect 54719 2700 54789 2746
rect 54835 2700 54905 2746
rect 54951 2700 55021 2746
rect 55067 2700 55137 2746
rect 55183 2700 55253 2746
rect 55299 2700 55369 2746
rect 55415 2700 55485 2746
rect 55531 2700 55601 2746
rect 55647 2700 55717 2746
rect 55763 2700 55833 2746
rect 55879 2700 55949 2746
rect 55995 2700 56065 2746
rect 56111 2700 56181 2746
rect 56227 2700 56297 2746
rect 56343 2700 56413 2746
rect 56459 2700 56529 2746
rect 56575 2700 56594 2746
rect 50826 2630 56594 2700
rect 50826 2584 50845 2630
rect 50891 2584 50961 2630
rect 51007 2584 51077 2630
rect 51123 2584 51193 2630
rect 51239 2584 51309 2630
rect 51355 2584 51425 2630
rect 51471 2584 51541 2630
rect 51587 2584 51657 2630
rect 51703 2584 51773 2630
rect 51819 2584 51889 2630
rect 51935 2584 52005 2630
rect 52051 2584 52121 2630
rect 52167 2584 52237 2630
rect 52283 2584 52353 2630
rect 52399 2584 52469 2630
rect 52515 2584 52585 2630
rect 52631 2584 52701 2630
rect 52747 2584 52817 2630
rect 52863 2584 52933 2630
rect 52979 2584 53049 2630
rect 53095 2584 53165 2630
rect 53211 2584 53281 2630
rect 53327 2584 53397 2630
rect 53443 2584 53513 2630
rect 53559 2584 53629 2630
rect 53675 2584 53745 2630
rect 53791 2584 53861 2630
rect 53907 2584 53977 2630
rect 54023 2584 54093 2630
rect 54139 2584 54209 2630
rect 54255 2584 54325 2630
rect 54371 2584 54441 2630
rect 54487 2584 54557 2630
rect 54603 2584 54673 2630
rect 54719 2584 54789 2630
rect 54835 2584 54905 2630
rect 54951 2584 55021 2630
rect 55067 2584 55137 2630
rect 55183 2584 55253 2630
rect 55299 2584 55369 2630
rect 55415 2584 55485 2630
rect 55531 2584 55601 2630
rect 55647 2584 55717 2630
rect 55763 2584 55833 2630
rect 55879 2584 55949 2630
rect 55995 2584 56065 2630
rect 56111 2584 56181 2630
rect 56227 2584 56297 2630
rect 56343 2584 56413 2630
rect 56459 2584 56529 2630
rect 56575 2584 56594 2630
rect 50826 2514 56594 2584
rect 50826 2468 50845 2514
rect 50891 2468 50961 2514
rect 51007 2468 51077 2514
rect 51123 2468 51193 2514
rect 51239 2468 51309 2514
rect 51355 2468 51425 2514
rect 51471 2468 51541 2514
rect 51587 2468 51657 2514
rect 51703 2468 51773 2514
rect 51819 2468 51889 2514
rect 51935 2468 52005 2514
rect 52051 2468 52121 2514
rect 52167 2468 52237 2514
rect 52283 2468 52353 2514
rect 52399 2468 52469 2514
rect 52515 2468 52585 2514
rect 52631 2468 52701 2514
rect 52747 2468 52817 2514
rect 52863 2468 52933 2514
rect 52979 2468 53049 2514
rect 53095 2468 53165 2514
rect 53211 2468 53281 2514
rect 53327 2468 53397 2514
rect 53443 2468 53513 2514
rect 53559 2468 53629 2514
rect 53675 2468 53745 2514
rect 53791 2468 53861 2514
rect 53907 2468 53977 2514
rect 54023 2468 54093 2514
rect 54139 2468 54209 2514
rect 54255 2468 54325 2514
rect 54371 2468 54441 2514
rect 54487 2468 54557 2514
rect 54603 2468 54673 2514
rect 54719 2468 54789 2514
rect 54835 2468 54905 2514
rect 54951 2468 55021 2514
rect 55067 2468 55137 2514
rect 55183 2468 55253 2514
rect 55299 2468 55369 2514
rect 55415 2468 55485 2514
rect 55531 2468 55601 2514
rect 55647 2468 55717 2514
rect 55763 2468 55833 2514
rect 55879 2468 55949 2514
rect 55995 2468 56065 2514
rect 56111 2468 56181 2514
rect 56227 2468 56297 2514
rect 56343 2468 56413 2514
rect 56459 2468 56529 2514
rect 56575 2468 56594 2514
rect 50826 2398 56594 2468
rect 50826 2352 50845 2398
rect 50891 2352 50961 2398
rect 51007 2352 51077 2398
rect 51123 2352 51193 2398
rect 51239 2352 51309 2398
rect 51355 2352 51425 2398
rect 51471 2352 51541 2398
rect 51587 2352 51657 2398
rect 51703 2352 51773 2398
rect 51819 2352 51889 2398
rect 51935 2352 52005 2398
rect 52051 2352 52121 2398
rect 52167 2352 52237 2398
rect 52283 2352 52353 2398
rect 52399 2352 52469 2398
rect 52515 2352 52585 2398
rect 52631 2352 52701 2398
rect 52747 2352 52817 2398
rect 52863 2352 52933 2398
rect 52979 2352 53049 2398
rect 53095 2352 53165 2398
rect 53211 2352 53281 2398
rect 53327 2352 53397 2398
rect 53443 2352 53513 2398
rect 53559 2352 53629 2398
rect 53675 2352 53745 2398
rect 53791 2352 53861 2398
rect 53907 2352 53977 2398
rect 54023 2352 54093 2398
rect 54139 2352 54209 2398
rect 54255 2352 54325 2398
rect 54371 2352 54441 2398
rect 54487 2352 54557 2398
rect 54603 2352 54673 2398
rect 54719 2352 54789 2398
rect 54835 2352 54905 2398
rect 54951 2352 55021 2398
rect 55067 2352 55137 2398
rect 55183 2352 55253 2398
rect 55299 2352 55369 2398
rect 55415 2352 55485 2398
rect 55531 2352 55601 2398
rect 55647 2352 55717 2398
rect 55763 2352 55833 2398
rect 55879 2352 55949 2398
rect 55995 2352 56065 2398
rect 56111 2352 56181 2398
rect 56227 2352 56297 2398
rect 56343 2352 56413 2398
rect 56459 2352 56529 2398
rect 56575 2352 56594 2398
rect 50826 2282 56594 2352
rect 50826 2236 50845 2282
rect 50891 2236 50961 2282
rect 51007 2236 51077 2282
rect 51123 2236 51193 2282
rect 51239 2236 51309 2282
rect 51355 2236 51425 2282
rect 51471 2236 51541 2282
rect 51587 2236 51657 2282
rect 51703 2236 51773 2282
rect 51819 2236 51889 2282
rect 51935 2236 52005 2282
rect 52051 2236 52121 2282
rect 52167 2236 52237 2282
rect 52283 2236 52353 2282
rect 52399 2236 52469 2282
rect 52515 2236 52585 2282
rect 52631 2236 52701 2282
rect 52747 2236 52817 2282
rect 52863 2236 52933 2282
rect 52979 2236 53049 2282
rect 53095 2236 53165 2282
rect 53211 2236 53281 2282
rect 53327 2236 53397 2282
rect 53443 2236 53513 2282
rect 53559 2236 53629 2282
rect 53675 2236 53745 2282
rect 53791 2236 53861 2282
rect 53907 2236 53977 2282
rect 54023 2236 54093 2282
rect 54139 2236 54209 2282
rect 54255 2236 54325 2282
rect 54371 2236 54441 2282
rect 54487 2236 54557 2282
rect 54603 2236 54673 2282
rect 54719 2236 54789 2282
rect 54835 2236 54905 2282
rect 54951 2236 55021 2282
rect 55067 2236 55137 2282
rect 55183 2236 55253 2282
rect 55299 2236 55369 2282
rect 55415 2236 55485 2282
rect 55531 2236 55601 2282
rect 55647 2236 55717 2282
rect 55763 2236 55833 2282
rect 55879 2236 55949 2282
rect 55995 2236 56065 2282
rect 56111 2236 56181 2282
rect 56227 2236 56297 2282
rect 56343 2236 56413 2282
rect 56459 2236 56529 2282
rect 56575 2236 56594 2282
rect 50826 2166 56594 2236
rect 50826 2120 50845 2166
rect 50891 2120 50961 2166
rect 51007 2120 51077 2166
rect 51123 2120 51193 2166
rect 51239 2120 51309 2166
rect 51355 2120 51425 2166
rect 51471 2120 51541 2166
rect 51587 2120 51657 2166
rect 51703 2120 51773 2166
rect 51819 2120 51889 2166
rect 51935 2120 52005 2166
rect 52051 2120 52121 2166
rect 52167 2120 52237 2166
rect 52283 2120 52353 2166
rect 52399 2120 52469 2166
rect 52515 2120 52585 2166
rect 52631 2120 52701 2166
rect 52747 2120 52817 2166
rect 52863 2120 52933 2166
rect 52979 2120 53049 2166
rect 53095 2120 53165 2166
rect 53211 2120 53281 2166
rect 53327 2120 53397 2166
rect 53443 2120 53513 2166
rect 53559 2120 53629 2166
rect 53675 2120 53745 2166
rect 53791 2120 53861 2166
rect 53907 2120 53977 2166
rect 54023 2120 54093 2166
rect 54139 2120 54209 2166
rect 54255 2120 54325 2166
rect 54371 2120 54441 2166
rect 54487 2120 54557 2166
rect 54603 2120 54673 2166
rect 54719 2120 54789 2166
rect 54835 2120 54905 2166
rect 54951 2120 55021 2166
rect 55067 2120 55137 2166
rect 55183 2120 55253 2166
rect 55299 2120 55369 2166
rect 55415 2120 55485 2166
rect 55531 2120 55601 2166
rect 55647 2120 55717 2166
rect 55763 2120 55833 2166
rect 55879 2120 55949 2166
rect 55995 2120 56065 2166
rect 56111 2120 56181 2166
rect 56227 2120 56297 2166
rect 56343 2120 56413 2166
rect 56459 2120 56529 2166
rect 56575 2120 56594 2166
rect 50826 2050 56594 2120
rect 50826 2004 50845 2050
rect 50891 2004 50961 2050
rect 51007 2004 51077 2050
rect 51123 2004 51193 2050
rect 51239 2004 51309 2050
rect 51355 2004 51425 2050
rect 51471 2004 51541 2050
rect 51587 2004 51657 2050
rect 51703 2004 51773 2050
rect 51819 2004 51889 2050
rect 51935 2004 52005 2050
rect 52051 2004 52121 2050
rect 52167 2004 52237 2050
rect 52283 2004 52353 2050
rect 52399 2004 52469 2050
rect 52515 2004 52585 2050
rect 52631 2004 52701 2050
rect 52747 2004 52817 2050
rect 52863 2004 52933 2050
rect 52979 2004 53049 2050
rect 53095 2004 53165 2050
rect 53211 2004 53281 2050
rect 53327 2004 53397 2050
rect 53443 2004 53513 2050
rect 53559 2004 53629 2050
rect 53675 2004 53745 2050
rect 53791 2004 53861 2050
rect 53907 2004 53977 2050
rect 54023 2004 54093 2050
rect 54139 2004 54209 2050
rect 54255 2004 54325 2050
rect 54371 2004 54441 2050
rect 54487 2004 54557 2050
rect 54603 2004 54673 2050
rect 54719 2004 54789 2050
rect 54835 2004 54905 2050
rect 54951 2004 55021 2050
rect 55067 2004 55137 2050
rect 55183 2004 55253 2050
rect 55299 2004 55369 2050
rect 55415 2004 55485 2050
rect 55531 2004 55601 2050
rect 55647 2004 55717 2050
rect 55763 2004 55833 2050
rect 55879 2004 55949 2050
rect 55995 2004 56065 2050
rect 56111 2004 56181 2050
rect 56227 2004 56297 2050
rect 56343 2004 56413 2050
rect 56459 2004 56529 2050
rect 56575 2004 56594 2050
rect 50826 1934 56594 2004
rect 50826 1888 50845 1934
rect 50891 1888 50961 1934
rect 51007 1888 51077 1934
rect 51123 1888 51193 1934
rect 51239 1888 51309 1934
rect 51355 1888 51425 1934
rect 51471 1888 51541 1934
rect 51587 1888 51657 1934
rect 51703 1888 51773 1934
rect 51819 1888 51889 1934
rect 51935 1888 52005 1934
rect 52051 1888 52121 1934
rect 52167 1888 52237 1934
rect 52283 1888 52353 1934
rect 52399 1888 52469 1934
rect 52515 1888 52585 1934
rect 52631 1888 52701 1934
rect 52747 1888 52817 1934
rect 52863 1888 52933 1934
rect 52979 1888 53049 1934
rect 53095 1888 53165 1934
rect 53211 1888 53281 1934
rect 53327 1888 53397 1934
rect 53443 1888 53513 1934
rect 53559 1888 53629 1934
rect 53675 1888 53745 1934
rect 53791 1888 53861 1934
rect 53907 1888 53977 1934
rect 54023 1888 54093 1934
rect 54139 1888 54209 1934
rect 54255 1888 54325 1934
rect 54371 1888 54441 1934
rect 54487 1888 54557 1934
rect 54603 1888 54673 1934
rect 54719 1888 54789 1934
rect 54835 1888 54905 1934
rect 54951 1888 55021 1934
rect 55067 1888 55137 1934
rect 55183 1888 55253 1934
rect 55299 1888 55369 1934
rect 55415 1888 55485 1934
rect 55531 1888 55601 1934
rect 55647 1888 55717 1934
rect 55763 1888 55833 1934
rect 55879 1888 55949 1934
rect 55995 1888 56065 1934
rect 56111 1888 56181 1934
rect 56227 1888 56297 1934
rect 56343 1888 56413 1934
rect 56459 1888 56529 1934
rect 56575 1888 56594 1934
rect 50826 1818 56594 1888
rect 50826 1772 50845 1818
rect 50891 1772 50961 1818
rect 51007 1772 51077 1818
rect 51123 1772 51193 1818
rect 51239 1772 51309 1818
rect 51355 1772 51425 1818
rect 51471 1772 51541 1818
rect 51587 1772 51657 1818
rect 51703 1772 51773 1818
rect 51819 1772 51889 1818
rect 51935 1772 52005 1818
rect 52051 1772 52121 1818
rect 52167 1772 52237 1818
rect 52283 1772 52353 1818
rect 52399 1772 52469 1818
rect 52515 1772 52585 1818
rect 52631 1772 52701 1818
rect 52747 1772 52817 1818
rect 52863 1772 52933 1818
rect 52979 1772 53049 1818
rect 53095 1772 53165 1818
rect 53211 1772 53281 1818
rect 53327 1772 53397 1818
rect 53443 1772 53513 1818
rect 53559 1772 53629 1818
rect 53675 1772 53745 1818
rect 53791 1772 53861 1818
rect 53907 1772 53977 1818
rect 54023 1772 54093 1818
rect 54139 1772 54209 1818
rect 54255 1772 54325 1818
rect 54371 1772 54441 1818
rect 54487 1772 54557 1818
rect 54603 1772 54673 1818
rect 54719 1772 54789 1818
rect 54835 1772 54905 1818
rect 54951 1772 55021 1818
rect 55067 1772 55137 1818
rect 55183 1772 55253 1818
rect 55299 1772 55369 1818
rect 55415 1772 55485 1818
rect 55531 1772 55601 1818
rect 55647 1772 55717 1818
rect 55763 1772 55833 1818
rect 55879 1772 55949 1818
rect 55995 1772 56065 1818
rect 56111 1772 56181 1818
rect 56227 1772 56297 1818
rect 56343 1772 56413 1818
rect 56459 1772 56529 1818
rect 56575 1772 56594 1818
rect 50826 1702 56594 1772
rect 50826 1656 50845 1702
rect 50891 1656 50961 1702
rect 51007 1656 51077 1702
rect 51123 1656 51193 1702
rect 51239 1656 51309 1702
rect 51355 1656 51425 1702
rect 51471 1656 51541 1702
rect 51587 1656 51657 1702
rect 51703 1656 51773 1702
rect 51819 1656 51889 1702
rect 51935 1656 52005 1702
rect 52051 1656 52121 1702
rect 52167 1656 52237 1702
rect 52283 1656 52353 1702
rect 52399 1656 52469 1702
rect 52515 1656 52585 1702
rect 52631 1656 52701 1702
rect 52747 1656 52817 1702
rect 52863 1656 52933 1702
rect 52979 1656 53049 1702
rect 53095 1656 53165 1702
rect 53211 1656 53281 1702
rect 53327 1656 53397 1702
rect 53443 1656 53513 1702
rect 53559 1656 53629 1702
rect 53675 1656 53745 1702
rect 53791 1656 53861 1702
rect 53907 1656 53977 1702
rect 54023 1656 54093 1702
rect 54139 1656 54209 1702
rect 54255 1656 54325 1702
rect 54371 1656 54441 1702
rect 54487 1656 54557 1702
rect 54603 1656 54673 1702
rect 54719 1656 54789 1702
rect 54835 1656 54905 1702
rect 54951 1656 55021 1702
rect 55067 1656 55137 1702
rect 55183 1656 55253 1702
rect 55299 1656 55369 1702
rect 55415 1656 55485 1702
rect 55531 1656 55601 1702
rect 55647 1656 55717 1702
rect 55763 1656 55833 1702
rect 55879 1656 55949 1702
rect 55995 1656 56065 1702
rect 56111 1656 56181 1702
rect 56227 1656 56297 1702
rect 56343 1656 56413 1702
rect 56459 1656 56529 1702
rect 56575 1656 56594 1702
rect 50826 1637 56594 1656
rect 27479 1030 27763 1117
rect 57361 1117 57380 34237
rect 57626 1117 57645 52963
rect 57361 1030 57645 1117
<< mvpsubdiffcont >>
rect 27498 1117 27744 52963
rect 27846 35996 28492 52942
rect 56632 35996 57278 52942
rect 27846 34256 57292 34602
rect 28639 3860 28685 3906
rect 28755 3860 28801 3906
rect 28871 3860 28917 3906
rect 28987 3860 29033 3906
rect 29103 3860 29149 3906
rect 29219 3860 29265 3906
rect 29335 3860 29381 3906
rect 29451 3860 29497 3906
rect 29567 3860 29613 3906
rect 29683 3860 29729 3906
rect 29799 3860 29845 3906
rect 29915 3860 29961 3906
rect 30031 3860 30077 3906
rect 30147 3860 30193 3906
rect 30263 3860 30309 3906
rect 30379 3860 30425 3906
rect 30495 3860 30541 3906
rect 30611 3860 30657 3906
rect 30727 3860 30773 3906
rect 30843 3860 30889 3906
rect 30959 3860 31005 3906
rect 31075 3860 31121 3906
rect 31191 3860 31237 3906
rect 31307 3860 31353 3906
rect 31423 3860 31469 3906
rect 31539 3860 31585 3906
rect 31655 3860 31701 3906
rect 31771 3860 31817 3906
rect 31887 3860 31933 3906
rect 32003 3860 32049 3906
rect 32119 3860 32165 3906
rect 32235 3860 32281 3906
rect 32351 3860 32397 3906
rect 32467 3860 32513 3906
rect 32583 3860 32629 3906
rect 32699 3860 32745 3906
rect 32815 3860 32861 3906
rect 32931 3860 32977 3906
rect 33047 3860 33093 3906
rect 33163 3860 33209 3906
rect 33279 3860 33325 3906
rect 33395 3860 33441 3906
rect 33511 3860 33557 3906
rect 33627 3860 33673 3906
rect 33743 3860 33789 3906
rect 33859 3860 33905 3906
rect 33975 3860 34021 3906
rect 34091 3860 34137 3906
rect 34207 3860 34253 3906
rect 34323 3860 34369 3906
rect 34439 3860 34485 3906
rect 34555 3860 34601 3906
rect 34671 3860 34717 3906
rect 34787 3860 34833 3906
rect 34903 3860 34949 3906
rect 35019 3860 35065 3906
rect 35135 3860 35181 3906
rect 35251 3860 35297 3906
rect 35367 3860 35413 3906
rect 35483 3860 35529 3906
rect 35599 3860 35645 3906
rect 35715 3860 35761 3906
rect 35831 3860 35877 3906
rect 35947 3860 35993 3906
rect 36063 3860 36109 3906
rect 36179 3860 36225 3906
rect 36295 3860 36341 3906
rect 36411 3860 36457 3906
rect 36527 3860 36573 3906
rect 36643 3860 36689 3906
rect 36759 3860 36805 3906
rect 36875 3860 36921 3906
rect 36991 3860 37037 3906
rect 37107 3860 37153 3906
rect 37223 3860 37269 3906
rect 37339 3860 37385 3906
rect 37455 3860 37501 3906
rect 37571 3860 37617 3906
rect 37687 3860 37733 3906
rect 37803 3860 37849 3906
rect 37919 3860 37965 3906
rect 38035 3860 38081 3906
rect 38151 3860 38197 3906
rect 38267 3860 38313 3906
rect 38383 3860 38429 3906
rect 38499 3860 38545 3906
rect 38615 3860 38661 3906
rect 38731 3860 38777 3906
rect 38847 3860 38893 3906
rect 38963 3860 39009 3906
rect 39079 3860 39125 3906
rect 39195 3860 39241 3906
rect 39311 3860 39357 3906
rect 39427 3860 39473 3906
rect 39543 3860 39589 3906
rect 39659 3860 39705 3906
rect 39775 3860 39821 3906
rect 39891 3860 39937 3906
rect 40007 3860 40053 3906
rect 40123 3860 40169 3906
rect 28639 3744 28685 3790
rect 28755 3744 28801 3790
rect 28871 3744 28917 3790
rect 28987 3744 29033 3790
rect 29103 3744 29149 3790
rect 29219 3744 29265 3790
rect 29335 3744 29381 3790
rect 29451 3744 29497 3790
rect 29567 3744 29613 3790
rect 29683 3744 29729 3790
rect 29799 3744 29845 3790
rect 29915 3744 29961 3790
rect 30031 3744 30077 3790
rect 30147 3744 30193 3790
rect 30263 3744 30309 3790
rect 30379 3744 30425 3790
rect 30495 3744 30541 3790
rect 30611 3744 30657 3790
rect 30727 3744 30773 3790
rect 30843 3744 30889 3790
rect 30959 3744 31005 3790
rect 31075 3744 31121 3790
rect 31191 3744 31237 3790
rect 31307 3744 31353 3790
rect 31423 3744 31469 3790
rect 31539 3744 31585 3790
rect 31655 3744 31701 3790
rect 31771 3744 31817 3790
rect 31887 3744 31933 3790
rect 32003 3744 32049 3790
rect 32119 3744 32165 3790
rect 32235 3744 32281 3790
rect 32351 3744 32397 3790
rect 32467 3744 32513 3790
rect 32583 3744 32629 3790
rect 32699 3744 32745 3790
rect 32815 3744 32861 3790
rect 32931 3744 32977 3790
rect 33047 3744 33093 3790
rect 33163 3744 33209 3790
rect 33279 3744 33325 3790
rect 33395 3744 33441 3790
rect 33511 3744 33557 3790
rect 33627 3744 33673 3790
rect 33743 3744 33789 3790
rect 33859 3744 33905 3790
rect 33975 3744 34021 3790
rect 34091 3744 34137 3790
rect 34207 3744 34253 3790
rect 34323 3744 34369 3790
rect 34439 3744 34485 3790
rect 34555 3744 34601 3790
rect 34671 3744 34717 3790
rect 34787 3744 34833 3790
rect 34903 3744 34949 3790
rect 35019 3744 35065 3790
rect 35135 3744 35181 3790
rect 35251 3744 35297 3790
rect 35367 3744 35413 3790
rect 35483 3744 35529 3790
rect 35599 3744 35645 3790
rect 35715 3744 35761 3790
rect 35831 3744 35877 3790
rect 35947 3744 35993 3790
rect 36063 3744 36109 3790
rect 36179 3744 36225 3790
rect 36295 3744 36341 3790
rect 36411 3744 36457 3790
rect 36527 3744 36573 3790
rect 36643 3744 36689 3790
rect 36759 3744 36805 3790
rect 36875 3744 36921 3790
rect 36991 3744 37037 3790
rect 37107 3744 37153 3790
rect 37223 3744 37269 3790
rect 37339 3744 37385 3790
rect 37455 3744 37501 3790
rect 37571 3744 37617 3790
rect 37687 3744 37733 3790
rect 37803 3744 37849 3790
rect 37919 3744 37965 3790
rect 38035 3744 38081 3790
rect 38151 3744 38197 3790
rect 38267 3744 38313 3790
rect 38383 3744 38429 3790
rect 38499 3744 38545 3790
rect 38615 3744 38661 3790
rect 38731 3744 38777 3790
rect 38847 3744 38893 3790
rect 38963 3744 39009 3790
rect 39079 3744 39125 3790
rect 39195 3744 39241 3790
rect 39311 3744 39357 3790
rect 39427 3744 39473 3790
rect 39543 3744 39589 3790
rect 39659 3744 39705 3790
rect 39775 3744 39821 3790
rect 39891 3744 39937 3790
rect 40007 3744 40053 3790
rect 40123 3744 40169 3790
rect 28639 3628 28685 3674
rect 28755 3628 28801 3674
rect 28871 3628 28917 3674
rect 28987 3628 29033 3674
rect 29103 3628 29149 3674
rect 29219 3628 29265 3674
rect 29335 3628 29381 3674
rect 29451 3628 29497 3674
rect 29567 3628 29613 3674
rect 29683 3628 29729 3674
rect 29799 3628 29845 3674
rect 29915 3628 29961 3674
rect 30031 3628 30077 3674
rect 30147 3628 30193 3674
rect 30263 3628 30309 3674
rect 30379 3628 30425 3674
rect 30495 3628 30541 3674
rect 30611 3628 30657 3674
rect 30727 3628 30773 3674
rect 30843 3628 30889 3674
rect 30959 3628 31005 3674
rect 31075 3628 31121 3674
rect 31191 3628 31237 3674
rect 31307 3628 31353 3674
rect 31423 3628 31469 3674
rect 31539 3628 31585 3674
rect 31655 3628 31701 3674
rect 31771 3628 31817 3674
rect 31887 3628 31933 3674
rect 32003 3628 32049 3674
rect 32119 3628 32165 3674
rect 32235 3628 32281 3674
rect 32351 3628 32397 3674
rect 32467 3628 32513 3674
rect 32583 3628 32629 3674
rect 32699 3628 32745 3674
rect 32815 3628 32861 3674
rect 32931 3628 32977 3674
rect 33047 3628 33093 3674
rect 33163 3628 33209 3674
rect 33279 3628 33325 3674
rect 33395 3628 33441 3674
rect 33511 3628 33557 3674
rect 33627 3628 33673 3674
rect 33743 3628 33789 3674
rect 33859 3628 33905 3674
rect 33975 3628 34021 3674
rect 34091 3628 34137 3674
rect 34207 3628 34253 3674
rect 34323 3628 34369 3674
rect 34439 3628 34485 3674
rect 34555 3628 34601 3674
rect 34671 3628 34717 3674
rect 34787 3628 34833 3674
rect 34903 3628 34949 3674
rect 35019 3628 35065 3674
rect 35135 3628 35181 3674
rect 35251 3628 35297 3674
rect 35367 3628 35413 3674
rect 35483 3628 35529 3674
rect 35599 3628 35645 3674
rect 35715 3628 35761 3674
rect 35831 3628 35877 3674
rect 35947 3628 35993 3674
rect 36063 3628 36109 3674
rect 36179 3628 36225 3674
rect 36295 3628 36341 3674
rect 36411 3628 36457 3674
rect 36527 3628 36573 3674
rect 36643 3628 36689 3674
rect 36759 3628 36805 3674
rect 36875 3628 36921 3674
rect 36991 3628 37037 3674
rect 37107 3628 37153 3674
rect 37223 3628 37269 3674
rect 37339 3628 37385 3674
rect 37455 3628 37501 3674
rect 37571 3628 37617 3674
rect 37687 3628 37733 3674
rect 37803 3628 37849 3674
rect 37919 3628 37965 3674
rect 38035 3628 38081 3674
rect 38151 3628 38197 3674
rect 38267 3628 38313 3674
rect 38383 3628 38429 3674
rect 38499 3628 38545 3674
rect 38615 3628 38661 3674
rect 38731 3628 38777 3674
rect 38847 3628 38893 3674
rect 38963 3628 39009 3674
rect 39079 3628 39125 3674
rect 39195 3628 39241 3674
rect 39311 3628 39357 3674
rect 39427 3628 39473 3674
rect 39543 3628 39589 3674
rect 39659 3628 39705 3674
rect 39775 3628 39821 3674
rect 39891 3628 39937 3674
rect 40007 3628 40053 3674
rect 40123 3628 40169 3674
rect 28639 3512 28685 3558
rect 28755 3512 28801 3558
rect 28871 3512 28917 3558
rect 28987 3512 29033 3558
rect 29103 3512 29149 3558
rect 29219 3512 29265 3558
rect 29335 3512 29381 3558
rect 29451 3512 29497 3558
rect 29567 3512 29613 3558
rect 29683 3512 29729 3558
rect 29799 3512 29845 3558
rect 29915 3512 29961 3558
rect 30031 3512 30077 3558
rect 30147 3512 30193 3558
rect 30263 3512 30309 3558
rect 30379 3512 30425 3558
rect 30495 3512 30541 3558
rect 30611 3512 30657 3558
rect 30727 3512 30773 3558
rect 30843 3512 30889 3558
rect 30959 3512 31005 3558
rect 31075 3512 31121 3558
rect 31191 3512 31237 3558
rect 31307 3512 31353 3558
rect 31423 3512 31469 3558
rect 31539 3512 31585 3558
rect 31655 3512 31701 3558
rect 31771 3512 31817 3558
rect 31887 3512 31933 3558
rect 32003 3512 32049 3558
rect 32119 3512 32165 3558
rect 32235 3512 32281 3558
rect 32351 3512 32397 3558
rect 32467 3512 32513 3558
rect 32583 3512 32629 3558
rect 32699 3512 32745 3558
rect 32815 3512 32861 3558
rect 32931 3512 32977 3558
rect 33047 3512 33093 3558
rect 33163 3512 33209 3558
rect 33279 3512 33325 3558
rect 33395 3512 33441 3558
rect 33511 3512 33557 3558
rect 33627 3512 33673 3558
rect 33743 3512 33789 3558
rect 33859 3512 33905 3558
rect 33975 3512 34021 3558
rect 34091 3512 34137 3558
rect 34207 3512 34253 3558
rect 34323 3512 34369 3558
rect 34439 3512 34485 3558
rect 34555 3512 34601 3558
rect 34671 3512 34717 3558
rect 34787 3512 34833 3558
rect 34903 3512 34949 3558
rect 35019 3512 35065 3558
rect 35135 3512 35181 3558
rect 35251 3512 35297 3558
rect 35367 3512 35413 3558
rect 35483 3512 35529 3558
rect 35599 3512 35645 3558
rect 35715 3512 35761 3558
rect 35831 3512 35877 3558
rect 35947 3512 35993 3558
rect 36063 3512 36109 3558
rect 36179 3512 36225 3558
rect 36295 3512 36341 3558
rect 36411 3512 36457 3558
rect 36527 3512 36573 3558
rect 36643 3512 36689 3558
rect 36759 3512 36805 3558
rect 36875 3512 36921 3558
rect 36991 3512 37037 3558
rect 37107 3512 37153 3558
rect 37223 3512 37269 3558
rect 37339 3512 37385 3558
rect 37455 3512 37501 3558
rect 37571 3512 37617 3558
rect 37687 3512 37733 3558
rect 37803 3512 37849 3558
rect 37919 3512 37965 3558
rect 38035 3512 38081 3558
rect 38151 3512 38197 3558
rect 38267 3512 38313 3558
rect 38383 3512 38429 3558
rect 38499 3512 38545 3558
rect 38615 3512 38661 3558
rect 38731 3512 38777 3558
rect 38847 3512 38893 3558
rect 38963 3512 39009 3558
rect 39079 3512 39125 3558
rect 39195 3512 39241 3558
rect 39311 3512 39357 3558
rect 39427 3512 39473 3558
rect 39543 3512 39589 3558
rect 39659 3512 39705 3558
rect 39775 3512 39821 3558
rect 39891 3512 39937 3558
rect 40007 3512 40053 3558
rect 40123 3512 40169 3558
rect 28639 3396 28685 3442
rect 28755 3396 28801 3442
rect 28871 3396 28917 3442
rect 28987 3396 29033 3442
rect 29103 3396 29149 3442
rect 29219 3396 29265 3442
rect 29335 3396 29381 3442
rect 29451 3396 29497 3442
rect 29567 3396 29613 3442
rect 29683 3396 29729 3442
rect 29799 3396 29845 3442
rect 29915 3396 29961 3442
rect 30031 3396 30077 3442
rect 30147 3396 30193 3442
rect 30263 3396 30309 3442
rect 30379 3396 30425 3442
rect 30495 3396 30541 3442
rect 30611 3396 30657 3442
rect 30727 3396 30773 3442
rect 30843 3396 30889 3442
rect 30959 3396 31005 3442
rect 31075 3396 31121 3442
rect 31191 3396 31237 3442
rect 31307 3396 31353 3442
rect 31423 3396 31469 3442
rect 31539 3396 31585 3442
rect 31655 3396 31701 3442
rect 31771 3396 31817 3442
rect 31887 3396 31933 3442
rect 32003 3396 32049 3442
rect 32119 3396 32165 3442
rect 32235 3396 32281 3442
rect 32351 3396 32397 3442
rect 32467 3396 32513 3442
rect 32583 3396 32629 3442
rect 32699 3396 32745 3442
rect 32815 3396 32861 3442
rect 32931 3396 32977 3442
rect 33047 3396 33093 3442
rect 33163 3396 33209 3442
rect 33279 3396 33325 3442
rect 33395 3396 33441 3442
rect 33511 3396 33557 3442
rect 33627 3396 33673 3442
rect 33743 3396 33789 3442
rect 33859 3396 33905 3442
rect 33975 3396 34021 3442
rect 34091 3396 34137 3442
rect 34207 3396 34253 3442
rect 34323 3396 34369 3442
rect 34439 3396 34485 3442
rect 34555 3396 34601 3442
rect 34671 3396 34717 3442
rect 34787 3396 34833 3442
rect 34903 3396 34949 3442
rect 35019 3396 35065 3442
rect 35135 3396 35181 3442
rect 35251 3396 35297 3442
rect 35367 3396 35413 3442
rect 35483 3396 35529 3442
rect 35599 3396 35645 3442
rect 35715 3396 35761 3442
rect 35831 3396 35877 3442
rect 35947 3396 35993 3442
rect 36063 3396 36109 3442
rect 36179 3396 36225 3442
rect 36295 3396 36341 3442
rect 36411 3396 36457 3442
rect 36527 3396 36573 3442
rect 36643 3396 36689 3442
rect 36759 3396 36805 3442
rect 36875 3396 36921 3442
rect 36991 3396 37037 3442
rect 37107 3396 37153 3442
rect 37223 3396 37269 3442
rect 37339 3396 37385 3442
rect 37455 3396 37501 3442
rect 37571 3396 37617 3442
rect 37687 3396 37733 3442
rect 37803 3396 37849 3442
rect 37919 3396 37965 3442
rect 38035 3396 38081 3442
rect 38151 3396 38197 3442
rect 38267 3396 38313 3442
rect 38383 3396 38429 3442
rect 38499 3396 38545 3442
rect 38615 3396 38661 3442
rect 38731 3396 38777 3442
rect 38847 3396 38893 3442
rect 38963 3396 39009 3442
rect 39079 3396 39125 3442
rect 39195 3396 39241 3442
rect 39311 3396 39357 3442
rect 39427 3396 39473 3442
rect 39543 3396 39589 3442
rect 39659 3396 39705 3442
rect 39775 3396 39821 3442
rect 39891 3396 39937 3442
rect 40007 3396 40053 3442
rect 40123 3396 40169 3442
rect 28639 3280 28685 3326
rect 28755 3280 28801 3326
rect 28871 3280 28917 3326
rect 28987 3280 29033 3326
rect 29103 3280 29149 3326
rect 29219 3280 29265 3326
rect 29335 3280 29381 3326
rect 29451 3280 29497 3326
rect 29567 3280 29613 3326
rect 29683 3280 29729 3326
rect 29799 3280 29845 3326
rect 29915 3280 29961 3326
rect 30031 3280 30077 3326
rect 30147 3280 30193 3326
rect 30263 3280 30309 3326
rect 30379 3280 30425 3326
rect 30495 3280 30541 3326
rect 30611 3280 30657 3326
rect 30727 3280 30773 3326
rect 30843 3280 30889 3326
rect 30959 3280 31005 3326
rect 31075 3280 31121 3326
rect 31191 3280 31237 3326
rect 31307 3280 31353 3326
rect 31423 3280 31469 3326
rect 31539 3280 31585 3326
rect 31655 3280 31701 3326
rect 31771 3280 31817 3326
rect 31887 3280 31933 3326
rect 32003 3280 32049 3326
rect 32119 3280 32165 3326
rect 32235 3280 32281 3326
rect 32351 3280 32397 3326
rect 32467 3280 32513 3326
rect 32583 3280 32629 3326
rect 32699 3280 32745 3326
rect 32815 3280 32861 3326
rect 32931 3280 32977 3326
rect 33047 3280 33093 3326
rect 33163 3280 33209 3326
rect 33279 3280 33325 3326
rect 33395 3280 33441 3326
rect 33511 3280 33557 3326
rect 33627 3280 33673 3326
rect 33743 3280 33789 3326
rect 33859 3280 33905 3326
rect 33975 3280 34021 3326
rect 34091 3280 34137 3326
rect 34207 3280 34253 3326
rect 34323 3280 34369 3326
rect 34439 3280 34485 3326
rect 34555 3280 34601 3326
rect 34671 3280 34717 3326
rect 34787 3280 34833 3326
rect 34903 3280 34949 3326
rect 35019 3280 35065 3326
rect 35135 3280 35181 3326
rect 35251 3280 35297 3326
rect 35367 3280 35413 3326
rect 35483 3280 35529 3326
rect 35599 3280 35645 3326
rect 35715 3280 35761 3326
rect 35831 3280 35877 3326
rect 35947 3280 35993 3326
rect 36063 3280 36109 3326
rect 36179 3280 36225 3326
rect 36295 3280 36341 3326
rect 36411 3280 36457 3326
rect 36527 3280 36573 3326
rect 36643 3280 36689 3326
rect 36759 3280 36805 3326
rect 36875 3280 36921 3326
rect 36991 3280 37037 3326
rect 37107 3280 37153 3326
rect 37223 3280 37269 3326
rect 37339 3280 37385 3326
rect 37455 3280 37501 3326
rect 37571 3280 37617 3326
rect 37687 3280 37733 3326
rect 37803 3280 37849 3326
rect 37919 3280 37965 3326
rect 38035 3280 38081 3326
rect 38151 3280 38197 3326
rect 38267 3280 38313 3326
rect 38383 3280 38429 3326
rect 38499 3280 38545 3326
rect 38615 3280 38661 3326
rect 38731 3280 38777 3326
rect 38847 3280 38893 3326
rect 38963 3280 39009 3326
rect 39079 3280 39125 3326
rect 39195 3280 39241 3326
rect 39311 3280 39357 3326
rect 39427 3280 39473 3326
rect 39543 3280 39589 3326
rect 39659 3280 39705 3326
rect 39775 3280 39821 3326
rect 39891 3280 39937 3326
rect 40007 3280 40053 3326
rect 40123 3280 40169 3326
rect 28639 3164 28685 3210
rect 28755 3164 28801 3210
rect 28871 3164 28917 3210
rect 28987 3164 29033 3210
rect 29103 3164 29149 3210
rect 29219 3164 29265 3210
rect 29335 3164 29381 3210
rect 29451 3164 29497 3210
rect 29567 3164 29613 3210
rect 29683 3164 29729 3210
rect 29799 3164 29845 3210
rect 29915 3164 29961 3210
rect 30031 3164 30077 3210
rect 30147 3164 30193 3210
rect 30263 3164 30309 3210
rect 30379 3164 30425 3210
rect 30495 3164 30541 3210
rect 30611 3164 30657 3210
rect 30727 3164 30773 3210
rect 30843 3164 30889 3210
rect 30959 3164 31005 3210
rect 31075 3164 31121 3210
rect 31191 3164 31237 3210
rect 31307 3164 31353 3210
rect 31423 3164 31469 3210
rect 31539 3164 31585 3210
rect 31655 3164 31701 3210
rect 31771 3164 31817 3210
rect 31887 3164 31933 3210
rect 32003 3164 32049 3210
rect 32119 3164 32165 3210
rect 32235 3164 32281 3210
rect 32351 3164 32397 3210
rect 32467 3164 32513 3210
rect 32583 3164 32629 3210
rect 32699 3164 32745 3210
rect 32815 3164 32861 3210
rect 32931 3164 32977 3210
rect 33047 3164 33093 3210
rect 33163 3164 33209 3210
rect 33279 3164 33325 3210
rect 33395 3164 33441 3210
rect 33511 3164 33557 3210
rect 33627 3164 33673 3210
rect 33743 3164 33789 3210
rect 33859 3164 33905 3210
rect 33975 3164 34021 3210
rect 34091 3164 34137 3210
rect 34207 3164 34253 3210
rect 34323 3164 34369 3210
rect 34439 3164 34485 3210
rect 34555 3164 34601 3210
rect 34671 3164 34717 3210
rect 34787 3164 34833 3210
rect 34903 3164 34949 3210
rect 35019 3164 35065 3210
rect 35135 3164 35181 3210
rect 35251 3164 35297 3210
rect 35367 3164 35413 3210
rect 35483 3164 35529 3210
rect 35599 3164 35645 3210
rect 35715 3164 35761 3210
rect 35831 3164 35877 3210
rect 35947 3164 35993 3210
rect 36063 3164 36109 3210
rect 36179 3164 36225 3210
rect 36295 3164 36341 3210
rect 36411 3164 36457 3210
rect 36527 3164 36573 3210
rect 36643 3164 36689 3210
rect 36759 3164 36805 3210
rect 36875 3164 36921 3210
rect 36991 3164 37037 3210
rect 37107 3164 37153 3210
rect 37223 3164 37269 3210
rect 37339 3164 37385 3210
rect 37455 3164 37501 3210
rect 37571 3164 37617 3210
rect 37687 3164 37733 3210
rect 37803 3164 37849 3210
rect 37919 3164 37965 3210
rect 38035 3164 38081 3210
rect 38151 3164 38197 3210
rect 38267 3164 38313 3210
rect 38383 3164 38429 3210
rect 38499 3164 38545 3210
rect 38615 3164 38661 3210
rect 38731 3164 38777 3210
rect 38847 3164 38893 3210
rect 38963 3164 39009 3210
rect 39079 3164 39125 3210
rect 39195 3164 39241 3210
rect 39311 3164 39357 3210
rect 39427 3164 39473 3210
rect 39543 3164 39589 3210
rect 39659 3164 39705 3210
rect 39775 3164 39821 3210
rect 39891 3164 39937 3210
rect 40007 3164 40053 3210
rect 40123 3164 40169 3210
rect 28639 3048 28685 3094
rect 28755 3048 28801 3094
rect 28871 3048 28917 3094
rect 28987 3048 29033 3094
rect 29103 3048 29149 3094
rect 29219 3048 29265 3094
rect 29335 3048 29381 3094
rect 29451 3048 29497 3094
rect 29567 3048 29613 3094
rect 29683 3048 29729 3094
rect 29799 3048 29845 3094
rect 29915 3048 29961 3094
rect 30031 3048 30077 3094
rect 30147 3048 30193 3094
rect 30263 3048 30309 3094
rect 30379 3048 30425 3094
rect 30495 3048 30541 3094
rect 30611 3048 30657 3094
rect 30727 3048 30773 3094
rect 30843 3048 30889 3094
rect 30959 3048 31005 3094
rect 31075 3048 31121 3094
rect 31191 3048 31237 3094
rect 31307 3048 31353 3094
rect 31423 3048 31469 3094
rect 31539 3048 31585 3094
rect 31655 3048 31701 3094
rect 31771 3048 31817 3094
rect 31887 3048 31933 3094
rect 32003 3048 32049 3094
rect 32119 3048 32165 3094
rect 32235 3048 32281 3094
rect 32351 3048 32397 3094
rect 32467 3048 32513 3094
rect 32583 3048 32629 3094
rect 32699 3048 32745 3094
rect 32815 3048 32861 3094
rect 32931 3048 32977 3094
rect 33047 3048 33093 3094
rect 33163 3048 33209 3094
rect 33279 3048 33325 3094
rect 33395 3048 33441 3094
rect 33511 3048 33557 3094
rect 33627 3048 33673 3094
rect 33743 3048 33789 3094
rect 33859 3048 33905 3094
rect 33975 3048 34021 3094
rect 34091 3048 34137 3094
rect 34207 3048 34253 3094
rect 34323 3048 34369 3094
rect 34439 3048 34485 3094
rect 34555 3048 34601 3094
rect 34671 3048 34717 3094
rect 34787 3048 34833 3094
rect 34903 3048 34949 3094
rect 35019 3048 35065 3094
rect 35135 3048 35181 3094
rect 35251 3048 35297 3094
rect 35367 3048 35413 3094
rect 35483 3048 35529 3094
rect 35599 3048 35645 3094
rect 35715 3048 35761 3094
rect 35831 3048 35877 3094
rect 35947 3048 35993 3094
rect 36063 3048 36109 3094
rect 36179 3048 36225 3094
rect 36295 3048 36341 3094
rect 36411 3048 36457 3094
rect 36527 3048 36573 3094
rect 36643 3048 36689 3094
rect 36759 3048 36805 3094
rect 36875 3048 36921 3094
rect 36991 3048 37037 3094
rect 37107 3048 37153 3094
rect 37223 3048 37269 3094
rect 37339 3048 37385 3094
rect 37455 3048 37501 3094
rect 37571 3048 37617 3094
rect 37687 3048 37733 3094
rect 37803 3048 37849 3094
rect 37919 3048 37965 3094
rect 38035 3048 38081 3094
rect 38151 3048 38197 3094
rect 38267 3048 38313 3094
rect 38383 3048 38429 3094
rect 38499 3048 38545 3094
rect 38615 3048 38661 3094
rect 38731 3048 38777 3094
rect 38847 3048 38893 3094
rect 38963 3048 39009 3094
rect 39079 3048 39125 3094
rect 39195 3048 39241 3094
rect 39311 3048 39357 3094
rect 39427 3048 39473 3094
rect 39543 3048 39589 3094
rect 39659 3048 39705 3094
rect 39775 3048 39821 3094
rect 39891 3048 39937 3094
rect 40007 3048 40053 3094
rect 40123 3048 40169 3094
rect 28639 2932 28685 2978
rect 28755 2932 28801 2978
rect 28871 2932 28917 2978
rect 28987 2932 29033 2978
rect 29103 2932 29149 2978
rect 29219 2932 29265 2978
rect 29335 2932 29381 2978
rect 29451 2932 29497 2978
rect 29567 2932 29613 2978
rect 29683 2932 29729 2978
rect 29799 2932 29845 2978
rect 29915 2932 29961 2978
rect 30031 2932 30077 2978
rect 30147 2932 30193 2978
rect 30263 2932 30309 2978
rect 30379 2932 30425 2978
rect 30495 2932 30541 2978
rect 30611 2932 30657 2978
rect 30727 2932 30773 2978
rect 30843 2932 30889 2978
rect 30959 2932 31005 2978
rect 31075 2932 31121 2978
rect 31191 2932 31237 2978
rect 31307 2932 31353 2978
rect 31423 2932 31469 2978
rect 31539 2932 31585 2978
rect 31655 2932 31701 2978
rect 31771 2932 31817 2978
rect 31887 2932 31933 2978
rect 32003 2932 32049 2978
rect 32119 2932 32165 2978
rect 32235 2932 32281 2978
rect 32351 2932 32397 2978
rect 32467 2932 32513 2978
rect 32583 2932 32629 2978
rect 32699 2932 32745 2978
rect 32815 2932 32861 2978
rect 32931 2932 32977 2978
rect 33047 2932 33093 2978
rect 33163 2932 33209 2978
rect 33279 2932 33325 2978
rect 33395 2932 33441 2978
rect 33511 2932 33557 2978
rect 33627 2932 33673 2978
rect 33743 2932 33789 2978
rect 33859 2932 33905 2978
rect 33975 2932 34021 2978
rect 34091 2932 34137 2978
rect 34207 2932 34253 2978
rect 34323 2932 34369 2978
rect 34439 2932 34485 2978
rect 34555 2932 34601 2978
rect 34671 2932 34717 2978
rect 34787 2932 34833 2978
rect 34903 2932 34949 2978
rect 35019 2932 35065 2978
rect 35135 2932 35181 2978
rect 35251 2932 35297 2978
rect 35367 2932 35413 2978
rect 35483 2932 35529 2978
rect 35599 2932 35645 2978
rect 35715 2932 35761 2978
rect 35831 2932 35877 2978
rect 35947 2932 35993 2978
rect 36063 2932 36109 2978
rect 36179 2932 36225 2978
rect 36295 2932 36341 2978
rect 36411 2932 36457 2978
rect 36527 2932 36573 2978
rect 36643 2932 36689 2978
rect 36759 2932 36805 2978
rect 36875 2932 36921 2978
rect 36991 2932 37037 2978
rect 37107 2932 37153 2978
rect 37223 2932 37269 2978
rect 37339 2932 37385 2978
rect 37455 2932 37501 2978
rect 37571 2932 37617 2978
rect 37687 2932 37733 2978
rect 37803 2932 37849 2978
rect 37919 2932 37965 2978
rect 38035 2932 38081 2978
rect 38151 2932 38197 2978
rect 38267 2932 38313 2978
rect 38383 2932 38429 2978
rect 38499 2932 38545 2978
rect 38615 2932 38661 2978
rect 38731 2932 38777 2978
rect 38847 2932 38893 2978
rect 38963 2932 39009 2978
rect 39079 2932 39125 2978
rect 39195 2932 39241 2978
rect 39311 2932 39357 2978
rect 39427 2932 39473 2978
rect 39543 2932 39589 2978
rect 39659 2932 39705 2978
rect 39775 2932 39821 2978
rect 39891 2932 39937 2978
rect 40007 2932 40053 2978
rect 40123 2932 40169 2978
rect 28639 2816 28685 2862
rect 28755 2816 28801 2862
rect 28871 2816 28917 2862
rect 28987 2816 29033 2862
rect 29103 2816 29149 2862
rect 29219 2816 29265 2862
rect 29335 2816 29381 2862
rect 29451 2816 29497 2862
rect 29567 2816 29613 2862
rect 29683 2816 29729 2862
rect 29799 2816 29845 2862
rect 29915 2816 29961 2862
rect 30031 2816 30077 2862
rect 30147 2816 30193 2862
rect 30263 2816 30309 2862
rect 30379 2816 30425 2862
rect 30495 2816 30541 2862
rect 30611 2816 30657 2862
rect 30727 2816 30773 2862
rect 30843 2816 30889 2862
rect 30959 2816 31005 2862
rect 31075 2816 31121 2862
rect 31191 2816 31237 2862
rect 31307 2816 31353 2862
rect 31423 2816 31469 2862
rect 31539 2816 31585 2862
rect 31655 2816 31701 2862
rect 31771 2816 31817 2862
rect 31887 2816 31933 2862
rect 32003 2816 32049 2862
rect 32119 2816 32165 2862
rect 32235 2816 32281 2862
rect 32351 2816 32397 2862
rect 32467 2816 32513 2862
rect 32583 2816 32629 2862
rect 32699 2816 32745 2862
rect 32815 2816 32861 2862
rect 32931 2816 32977 2862
rect 33047 2816 33093 2862
rect 33163 2816 33209 2862
rect 33279 2816 33325 2862
rect 33395 2816 33441 2862
rect 33511 2816 33557 2862
rect 33627 2816 33673 2862
rect 33743 2816 33789 2862
rect 33859 2816 33905 2862
rect 33975 2816 34021 2862
rect 34091 2816 34137 2862
rect 34207 2816 34253 2862
rect 34323 2816 34369 2862
rect 34439 2816 34485 2862
rect 34555 2816 34601 2862
rect 34671 2816 34717 2862
rect 34787 2816 34833 2862
rect 34903 2816 34949 2862
rect 35019 2816 35065 2862
rect 35135 2816 35181 2862
rect 35251 2816 35297 2862
rect 35367 2816 35413 2862
rect 35483 2816 35529 2862
rect 35599 2816 35645 2862
rect 35715 2816 35761 2862
rect 35831 2816 35877 2862
rect 35947 2816 35993 2862
rect 36063 2816 36109 2862
rect 36179 2816 36225 2862
rect 36295 2816 36341 2862
rect 36411 2816 36457 2862
rect 36527 2816 36573 2862
rect 36643 2816 36689 2862
rect 36759 2816 36805 2862
rect 36875 2816 36921 2862
rect 36991 2816 37037 2862
rect 37107 2816 37153 2862
rect 37223 2816 37269 2862
rect 37339 2816 37385 2862
rect 37455 2816 37501 2862
rect 37571 2816 37617 2862
rect 37687 2816 37733 2862
rect 37803 2816 37849 2862
rect 37919 2816 37965 2862
rect 38035 2816 38081 2862
rect 38151 2816 38197 2862
rect 38267 2816 38313 2862
rect 38383 2816 38429 2862
rect 38499 2816 38545 2862
rect 38615 2816 38661 2862
rect 38731 2816 38777 2862
rect 38847 2816 38893 2862
rect 38963 2816 39009 2862
rect 39079 2816 39125 2862
rect 39195 2816 39241 2862
rect 39311 2816 39357 2862
rect 39427 2816 39473 2862
rect 39543 2816 39589 2862
rect 39659 2816 39705 2862
rect 39775 2816 39821 2862
rect 39891 2816 39937 2862
rect 40007 2816 40053 2862
rect 40123 2816 40169 2862
rect 28639 2700 28685 2746
rect 28755 2700 28801 2746
rect 28871 2700 28917 2746
rect 28987 2700 29033 2746
rect 29103 2700 29149 2746
rect 29219 2700 29265 2746
rect 29335 2700 29381 2746
rect 29451 2700 29497 2746
rect 29567 2700 29613 2746
rect 29683 2700 29729 2746
rect 29799 2700 29845 2746
rect 29915 2700 29961 2746
rect 30031 2700 30077 2746
rect 30147 2700 30193 2746
rect 30263 2700 30309 2746
rect 30379 2700 30425 2746
rect 30495 2700 30541 2746
rect 30611 2700 30657 2746
rect 30727 2700 30773 2746
rect 30843 2700 30889 2746
rect 30959 2700 31005 2746
rect 31075 2700 31121 2746
rect 31191 2700 31237 2746
rect 31307 2700 31353 2746
rect 31423 2700 31469 2746
rect 31539 2700 31585 2746
rect 31655 2700 31701 2746
rect 31771 2700 31817 2746
rect 31887 2700 31933 2746
rect 32003 2700 32049 2746
rect 32119 2700 32165 2746
rect 32235 2700 32281 2746
rect 32351 2700 32397 2746
rect 32467 2700 32513 2746
rect 32583 2700 32629 2746
rect 32699 2700 32745 2746
rect 32815 2700 32861 2746
rect 32931 2700 32977 2746
rect 33047 2700 33093 2746
rect 33163 2700 33209 2746
rect 33279 2700 33325 2746
rect 33395 2700 33441 2746
rect 33511 2700 33557 2746
rect 33627 2700 33673 2746
rect 33743 2700 33789 2746
rect 33859 2700 33905 2746
rect 33975 2700 34021 2746
rect 34091 2700 34137 2746
rect 34207 2700 34253 2746
rect 34323 2700 34369 2746
rect 34439 2700 34485 2746
rect 34555 2700 34601 2746
rect 34671 2700 34717 2746
rect 34787 2700 34833 2746
rect 34903 2700 34949 2746
rect 35019 2700 35065 2746
rect 35135 2700 35181 2746
rect 35251 2700 35297 2746
rect 35367 2700 35413 2746
rect 35483 2700 35529 2746
rect 35599 2700 35645 2746
rect 35715 2700 35761 2746
rect 35831 2700 35877 2746
rect 35947 2700 35993 2746
rect 36063 2700 36109 2746
rect 36179 2700 36225 2746
rect 36295 2700 36341 2746
rect 36411 2700 36457 2746
rect 36527 2700 36573 2746
rect 36643 2700 36689 2746
rect 36759 2700 36805 2746
rect 36875 2700 36921 2746
rect 36991 2700 37037 2746
rect 37107 2700 37153 2746
rect 37223 2700 37269 2746
rect 37339 2700 37385 2746
rect 37455 2700 37501 2746
rect 37571 2700 37617 2746
rect 37687 2700 37733 2746
rect 37803 2700 37849 2746
rect 37919 2700 37965 2746
rect 38035 2700 38081 2746
rect 38151 2700 38197 2746
rect 38267 2700 38313 2746
rect 38383 2700 38429 2746
rect 38499 2700 38545 2746
rect 38615 2700 38661 2746
rect 38731 2700 38777 2746
rect 38847 2700 38893 2746
rect 38963 2700 39009 2746
rect 39079 2700 39125 2746
rect 39195 2700 39241 2746
rect 39311 2700 39357 2746
rect 39427 2700 39473 2746
rect 39543 2700 39589 2746
rect 39659 2700 39705 2746
rect 39775 2700 39821 2746
rect 39891 2700 39937 2746
rect 40007 2700 40053 2746
rect 40123 2700 40169 2746
rect 28639 2584 28685 2630
rect 28755 2584 28801 2630
rect 28871 2584 28917 2630
rect 28987 2584 29033 2630
rect 29103 2584 29149 2630
rect 29219 2584 29265 2630
rect 29335 2584 29381 2630
rect 29451 2584 29497 2630
rect 29567 2584 29613 2630
rect 29683 2584 29729 2630
rect 29799 2584 29845 2630
rect 29915 2584 29961 2630
rect 30031 2584 30077 2630
rect 30147 2584 30193 2630
rect 30263 2584 30309 2630
rect 30379 2584 30425 2630
rect 30495 2584 30541 2630
rect 30611 2584 30657 2630
rect 30727 2584 30773 2630
rect 30843 2584 30889 2630
rect 30959 2584 31005 2630
rect 31075 2584 31121 2630
rect 31191 2584 31237 2630
rect 31307 2584 31353 2630
rect 31423 2584 31469 2630
rect 31539 2584 31585 2630
rect 31655 2584 31701 2630
rect 31771 2584 31817 2630
rect 31887 2584 31933 2630
rect 32003 2584 32049 2630
rect 32119 2584 32165 2630
rect 32235 2584 32281 2630
rect 32351 2584 32397 2630
rect 32467 2584 32513 2630
rect 32583 2584 32629 2630
rect 32699 2584 32745 2630
rect 32815 2584 32861 2630
rect 32931 2584 32977 2630
rect 33047 2584 33093 2630
rect 33163 2584 33209 2630
rect 33279 2584 33325 2630
rect 33395 2584 33441 2630
rect 33511 2584 33557 2630
rect 33627 2584 33673 2630
rect 33743 2584 33789 2630
rect 33859 2584 33905 2630
rect 33975 2584 34021 2630
rect 34091 2584 34137 2630
rect 34207 2584 34253 2630
rect 34323 2584 34369 2630
rect 34439 2584 34485 2630
rect 34555 2584 34601 2630
rect 34671 2584 34717 2630
rect 34787 2584 34833 2630
rect 34903 2584 34949 2630
rect 35019 2584 35065 2630
rect 35135 2584 35181 2630
rect 35251 2584 35297 2630
rect 35367 2584 35413 2630
rect 35483 2584 35529 2630
rect 35599 2584 35645 2630
rect 35715 2584 35761 2630
rect 35831 2584 35877 2630
rect 35947 2584 35993 2630
rect 36063 2584 36109 2630
rect 36179 2584 36225 2630
rect 36295 2584 36341 2630
rect 36411 2584 36457 2630
rect 36527 2584 36573 2630
rect 36643 2584 36689 2630
rect 36759 2584 36805 2630
rect 36875 2584 36921 2630
rect 36991 2584 37037 2630
rect 37107 2584 37153 2630
rect 37223 2584 37269 2630
rect 37339 2584 37385 2630
rect 37455 2584 37501 2630
rect 37571 2584 37617 2630
rect 37687 2584 37733 2630
rect 37803 2584 37849 2630
rect 37919 2584 37965 2630
rect 38035 2584 38081 2630
rect 38151 2584 38197 2630
rect 38267 2584 38313 2630
rect 38383 2584 38429 2630
rect 38499 2584 38545 2630
rect 38615 2584 38661 2630
rect 38731 2584 38777 2630
rect 38847 2584 38893 2630
rect 38963 2584 39009 2630
rect 39079 2584 39125 2630
rect 39195 2584 39241 2630
rect 39311 2584 39357 2630
rect 39427 2584 39473 2630
rect 39543 2584 39589 2630
rect 39659 2584 39705 2630
rect 39775 2584 39821 2630
rect 39891 2584 39937 2630
rect 40007 2584 40053 2630
rect 40123 2584 40169 2630
rect 28639 2468 28685 2514
rect 28755 2468 28801 2514
rect 28871 2468 28917 2514
rect 28987 2468 29033 2514
rect 29103 2468 29149 2514
rect 29219 2468 29265 2514
rect 29335 2468 29381 2514
rect 29451 2468 29497 2514
rect 29567 2468 29613 2514
rect 29683 2468 29729 2514
rect 29799 2468 29845 2514
rect 29915 2468 29961 2514
rect 30031 2468 30077 2514
rect 30147 2468 30193 2514
rect 30263 2468 30309 2514
rect 30379 2468 30425 2514
rect 30495 2468 30541 2514
rect 30611 2468 30657 2514
rect 30727 2468 30773 2514
rect 30843 2468 30889 2514
rect 30959 2468 31005 2514
rect 31075 2468 31121 2514
rect 31191 2468 31237 2514
rect 31307 2468 31353 2514
rect 31423 2468 31469 2514
rect 31539 2468 31585 2514
rect 31655 2468 31701 2514
rect 31771 2468 31817 2514
rect 31887 2468 31933 2514
rect 32003 2468 32049 2514
rect 32119 2468 32165 2514
rect 32235 2468 32281 2514
rect 32351 2468 32397 2514
rect 32467 2468 32513 2514
rect 32583 2468 32629 2514
rect 32699 2468 32745 2514
rect 32815 2468 32861 2514
rect 32931 2468 32977 2514
rect 33047 2468 33093 2514
rect 33163 2468 33209 2514
rect 33279 2468 33325 2514
rect 33395 2468 33441 2514
rect 33511 2468 33557 2514
rect 33627 2468 33673 2514
rect 33743 2468 33789 2514
rect 33859 2468 33905 2514
rect 33975 2468 34021 2514
rect 34091 2468 34137 2514
rect 34207 2468 34253 2514
rect 34323 2468 34369 2514
rect 34439 2468 34485 2514
rect 34555 2468 34601 2514
rect 34671 2468 34717 2514
rect 34787 2468 34833 2514
rect 34903 2468 34949 2514
rect 35019 2468 35065 2514
rect 35135 2468 35181 2514
rect 35251 2468 35297 2514
rect 35367 2468 35413 2514
rect 35483 2468 35529 2514
rect 35599 2468 35645 2514
rect 35715 2468 35761 2514
rect 35831 2468 35877 2514
rect 35947 2468 35993 2514
rect 36063 2468 36109 2514
rect 36179 2468 36225 2514
rect 36295 2468 36341 2514
rect 36411 2468 36457 2514
rect 36527 2468 36573 2514
rect 36643 2468 36689 2514
rect 36759 2468 36805 2514
rect 36875 2468 36921 2514
rect 36991 2468 37037 2514
rect 37107 2468 37153 2514
rect 37223 2468 37269 2514
rect 37339 2468 37385 2514
rect 37455 2468 37501 2514
rect 37571 2468 37617 2514
rect 37687 2468 37733 2514
rect 37803 2468 37849 2514
rect 37919 2468 37965 2514
rect 38035 2468 38081 2514
rect 38151 2468 38197 2514
rect 38267 2468 38313 2514
rect 38383 2468 38429 2514
rect 38499 2468 38545 2514
rect 38615 2468 38661 2514
rect 38731 2468 38777 2514
rect 38847 2468 38893 2514
rect 38963 2468 39009 2514
rect 39079 2468 39125 2514
rect 39195 2468 39241 2514
rect 39311 2468 39357 2514
rect 39427 2468 39473 2514
rect 39543 2468 39589 2514
rect 39659 2468 39705 2514
rect 39775 2468 39821 2514
rect 39891 2468 39937 2514
rect 40007 2468 40053 2514
rect 40123 2468 40169 2514
rect 28639 2352 28685 2398
rect 28755 2352 28801 2398
rect 28871 2352 28917 2398
rect 28987 2352 29033 2398
rect 29103 2352 29149 2398
rect 29219 2352 29265 2398
rect 29335 2352 29381 2398
rect 29451 2352 29497 2398
rect 29567 2352 29613 2398
rect 29683 2352 29729 2398
rect 29799 2352 29845 2398
rect 29915 2352 29961 2398
rect 30031 2352 30077 2398
rect 30147 2352 30193 2398
rect 30263 2352 30309 2398
rect 30379 2352 30425 2398
rect 30495 2352 30541 2398
rect 30611 2352 30657 2398
rect 30727 2352 30773 2398
rect 30843 2352 30889 2398
rect 30959 2352 31005 2398
rect 31075 2352 31121 2398
rect 31191 2352 31237 2398
rect 31307 2352 31353 2398
rect 31423 2352 31469 2398
rect 31539 2352 31585 2398
rect 31655 2352 31701 2398
rect 31771 2352 31817 2398
rect 31887 2352 31933 2398
rect 32003 2352 32049 2398
rect 32119 2352 32165 2398
rect 32235 2352 32281 2398
rect 32351 2352 32397 2398
rect 32467 2352 32513 2398
rect 32583 2352 32629 2398
rect 32699 2352 32745 2398
rect 32815 2352 32861 2398
rect 32931 2352 32977 2398
rect 33047 2352 33093 2398
rect 33163 2352 33209 2398
rect 33279 2352 33325 2398
rect 33395 2352 33441 2398
rect 33511 2352 33557 2398
rect 33627 2352 33673 2398
rect 33743 2352 33789 2398
rect 33859 2352 33905 2398
rect 33975 2352 34021 2398
rect 34091 2352 34137 2398
rect 34207 2352 34253 2398
rect 34323 2352 34369 2398
rect 34439 2352 34485 2398
rect 34555 2352 34601 2398
rect 34671 2352 34717 2398
rect 34787 2352 34833 2398
rect 34903 2352 34949 2398
rect 35019 2352 35065 2398
rect 35135 2352 35181 2398
rect 35251 2352 35297 2398
rect 35367 2352 35413 2398
rect 35483 2352 35529 2398
rect 35599 2352 35645 2398
rect 35715 2352 35761 2398
rect 35831 2352 35877 2398
rect 35947 2352 35993 2398
rect 36063 2352 36109 2398
rect 36179 2352 36225 2398
rect 36295 2352 36341 2398
rect 36411 2352 36457 2398
rect 36527 2352 36573 2398
rect 36643 2352 36689 2398
rect 36759 2352 36805 2398
rect 36875 2352 36921 2398
rect 36991 2352 37037 2398
rect 37107 2352 37153 2398
rect 37223 2352 37269 2398
rect 37339 2352 37385 2398
rect 37455 2352 37501 2398
rect 37571 2352 37617 2398
rect 37687 2352 37733 2398
rect 37803 2352 37849 2398
rect 37919 2352 37965 2398
rect 38035 2352 38081 2398
rect 38151 2352 38197 2398
rect 38267 2352 38313 2398
rect 38383 2352 38429 2398
rect 38499 2352 38545 2398
rect 38615 2352 38661 2398
rect 38731 2352 38777 2398
rect 38847 2352 38893 2398
rect 38963 2352 39009 2398
rect 39079 2352 39125 2398
rect 39195 2352 39241 2398
rect 39311 2352 39357 2398
rect 39427 2352 39473 2398
rect 39543 2352 39589 2398
rect 39659 2352 39705 2398
rect 39775 2352 39821 2398
rect 39891 2352 39937 2398
rect 40007 2352 40053 2398
rect 40123 2352 40169 2398
rect 28639 2236 28685 2282
rect 28755 2236 28801 2282
rect 28871 2236 28917 2282
rect 28987 2236 29033 2282
rect 29103 2236 29149 2282
rect 29219 2236 29265 2282
rect 29335 2236 29381 2282
rect 29451 2236 29497 2282
rect 29567 2236 29613 2282
rect 29683 2236 29729 2282
rect 29799 2236 29845 2282
rect 29915 2236 29961 2282
rect 30031 2236 30077 2282
rect 30147 2236 30193 2282
rect 30263 2236 30309 2282
rect 30379 2236 30425 2282
rect 30495 2236 30541 2282
rect 30611 2236 30657 2282
rect 30727 2236 30773 2282
rect 30843 2236 30889 2282
rect 30959 2236 31005 2282
rect 31075 2236 31121 2282
rect 31191 2236 31237 2282
rect 31307 2236 31353 2282
rect 31423 2236 31469 2282
rect 31539 2236 31585 2282
rect 31655 2236 31701 2282
rect 31771 2236 31817 2282
rect 31887 2236 31933 2282
rect 32003 2236 32049 2282
rect 32119 2236 32165 2282
rect 32235 2236 32281 2282
rect 32351 2236 32397 2282
rect 32467 2236 32513 2282
rect 32583 2236 32629 2282
rect 32699 2236 32745 2282
rect 32815 2236 32861 2282
rect 32931 2236 32977 2282
rect 33047 2236 33093 2282
rect 33163 2236 33209 2282
rect 33279 2236 33325 2282
rect 33395 2236 33441 2282
rect 33511 2236 33557 2282
rect 33627 2236 33673 2282
rect 33743 2236 33789 2282
rect 33859 2236 33905 2282
rect 33975 2236 34021 2282
rect 34091 2236 34137 2282
rect 34207 2236 34253 2282
rect 34323 2236 34369 2282
rect 34439 2236 34485 2282
rect 34555 2236 34601 2282
rect 34671 2236 34717 2282
rect 34787 2236 34833 2282
rect 34903 2236 34949 2282
rect 35019 2236 35065 2282
rect 35135 2236 35181 2282
rect 35251 2236 35297 2282
rect 35367 2236 35413 2282
rect 35483 2236 35529 2282
rect 35599 2236 35645 2282
rect 35715 2236 35761 2282
rect 35831 2236 35877 2282
rect 35947 2236 35993 2282
rect 36063 2236 36109 2282
rect 36179 2236 36225 2282
rect 36295 2236 36341 2282
rect 36411 2236 36457 2282
rect 36527 2236 36573 2282
rect 36643 2236 36689 2282
rect 36759 2236 36805 2282
rect 36875 2236 36921 2282
rect 36991 2236 37037 2282
rect 37107 2236 37153 2282
rect 37223 2236 37269 2282
rect 37339 2236 37385 2282
rect 37455 2236 37501 2282
rect 37571 2236 37617 2282
rect 37687 2236 37733 2282
rect 37803 2236 37849 2282
rect 37919 2236 37965 2282
rect 38035 2236 38081 2282
rect 38151 2236 38197 2282
rect 38267 2236 38313 2282
rect 38383 2236 38429 2282
rect 38499 2236 38545 2282
rect 38615 2236 38661 2282
rect 38731 2236 38777 2282
rect 38847 2236 38893 2282
rect 38963 2236 39009 2282
rect 39079 2236 39125 2282
rect 39195 2236 39241 2282
rect 39311 2236 39357 2282
rect 39427 2236 39473 2282
rect 39543 2236 39589 2282
rect 39659 2236 39705 2282
rect 39775 2236 39821 2282
rect 39891 2236 39937 2282
rect 40007 2236 40053 2282
rect 40123 2236 40169 2282
rect 28639 2120 28685 2166
rect 28755 2120 28801 2166
rect 28871 2120 28917 2166
rect 28987 2120 29033 2166
rect 29103 2120 29149 2166
rect 29219 2120 29265 2166
rect 29335 2120 29381 2166
rect 29451 2120 29497 2166
rect 29567 2120 29613 2166
rect 29683 2120 29729 2166
rect 29799 2120 29845 2166
rect 29915 2120 29961 2166
rect 30031 2120 30077 2166
rect 30147 2120 30193 2166
rect 30263 2120 30309 2166
rect 30379 2120 30425 2166
rect 30495 2120 30541 2166
rect 30611 2120 30657 2166
rect 30727 2120 30773 2166
rect 30843 2120 30889 2166
rect 30959 2120 31005 2166
rect 31075 2120 31121 2166
rect 31191 2120 31237 2166
rect 31307 2120 31353 2166
rect 31423 2120 31469 2166
rect 31539 2120 31585 2166
rect 31655 2120 31701 2166
rect 31771 2120 31817 2166
rect 31887 2120 31933 2166
rect 32003 2120 32049 2166
rect 32119 2120 32165 2166
rect 32235 2120 32281 2166
rect 32351 2120 32397 2166
rect 32467 2120 32513 2166
rect 32583 2120 32629 2166
rect 32699 2120 32745 2166
rect 32815 2120 32861 2166
rect 32931 2120 32977 2166
rect 33047 2120 33093 2166
rect 33163 2120 33209 2166
rect 33279 2120 33325 2166
rect 33395 2120 33441 2166
rect 33511 2120 33557 2166
rect 33627 2120 33673 2166
rect 33743 2120 33789 2166
rect 33859 2120 33905 2166
rect 33975 2120 34021 2166
rect 34091 2120 34137 2166
rect 34207 2120 34253 2166
rect 34323 2120 34369 2166
rect 34439 2120 34485 2166
rect 34555 2120 34601 2166
rect 34671 2120 34717 2166
rect 34787 2120 34833 2166
rect 34903 2120 34949 2166
rect 35019 2120 35065 2166
rect 35135 2120 35181 2166
rect 35251 2120 35297 2166
rect 35367 2120 35413 2166
rect 35483 2120 35529 2166
rect 35599 2120 35645 2166
rect 35715 2120 35761 2166
rect 35831 2120 35877 2166
rect 35947 2120 35993 2166
rect 36063 2120 36109 2166
rect 36179 2120 36225 2166
rect 36295 2120 36341 2166
rect 36411 2120 36457 2166
rect 36527 2120 36573 2166
rect 36643 2120 36689 2166
rect 36759 2120 36805 2166
rect 36875 2120 36921 2166
rect 36991 2120 37037 2166
rect 37107 2120 37153 2166
rect 37223 2120 37269 2166
rect 37339 2120 37385 2166
rect 37455 2120 37501 2166
rect 37571 2120 37617 2166
rect 37687 2120 37733 2166
rect 37803 2120 37849 2166
rect 37919 2120 37965 2166
rect 38035 2120 38081 2166
rect 38151 2120 38197 2166
rect 38267 2120 38313 2166
rect 38383 2120 38429 2166
rect 38499 2120 38545 2166
rect 38615 2120 38661 2166
rect 38731 2120 38777 2166
rect 38847 2120 38893 2166
rect 38963 2120 39009 2166
rect 39079 2120 39125 2166
rect 39195 2120 39241 2166
rect 39311 2120 39357 2166
rect 39427 2120 39473 2166
rect 39543 2120 39589 2166
rect 39659 2120 39705 2166
rect 39775 2120 39821 2166
rect 39891 2120 39937 2166
rect 40007 2120 40053 2166
rect 40123 2120 40169 2166
rect 28639 2004 28685 2050
rect 28755 2004 28801 2050
rect 28871 2004 28917 2050
rect 28987 2004 29033 2050
rect 29103 2004 29149 2050
rect 29219 2004 29265 2050
rect 29335 2004 29381 2050
rect 29451 2004 29497 2050
rect 29567 2004 29613 2050
rect 29683 2004 29729 2050
rect 29799 2004 29845 2050
rect 29915 2004 29961 2050
rect 30031 2004 30077 2050
rect 30147 2004 30193 2050
rect 30263 2004 30309 2050
rect 30379 2004 30425 2050
rect 30495 2004 30541 2050
rect 30611 2004 30657 2050
rect 30727 2004 30773 2050
rect 30843 2004 30889 2050
rect 30959 2004 31005 2050
rect 31075 2004 31121 2050
rect 31191 2004 31237 2050
rect 31307 2004 31353 2050
rect 31423 2004 31469 2050
rect 31539 2004 31585 2050
rect 31655 2004 31701 2050
rect 31771 2004 31817 2050
rect 31887 2004 31933 2050
rect 32003 2004 32049 2050
rect 32119 2004 32165 2050
rect 32235 2004 32281 2050
rect 32351 2004 32397 2050
rect 32467 2004 32513 2050
rect 32583 2004 32629 2050
rect 32699 2004 32745 2050
rect 32815 2004 32861 2050
rect 32931 2004 32977 2050
rect 33047 2004 33093 2050
rect 33163 2004 33209 2050
rect 33279 2004 33325 2050
rect 33395 2004 33441 2050
rect 33511 2004 33557 2050
rect 33627 2004 33673 2050
rect 33743 2004 33789 2050
rect 33859 2004 33905 2050
rect 33975 2004 34021 2050
rect 34091 2004 34137 2050
rect 34207 2004 34253 2050
rect 34323 2004 34369 2050
rect 34439 2004 34485 2050
rect 34555 2004 34601 2050
rect 34671 2004 34717 2050
rect 34787 2004 34833 2050
rect 34903 2004 34949 2050
rect 35019 2004 35065 2050
rect 35135 2004 35181 2050
rect 35251 2004 35297 2050
rect 35367 2004 35413 2050
rect 35483 2004 35529 2050
rect 35599 2004 35645 2050
rect 35715 2004 35761 2050
rect 35831 2004 35877 2050
rect 35947 2004 35993 2050
rect 36063 2004 36109 2050
rect 36179 2004 36225 2050
rect 36295 2004 36341 2050
rect 36411 2004 36457 2050
rect 36527 2004 36573 2050
rect 36643 2004 36689 2050
rect 36759 2004 36805 2050
rect 36875 2004 36921 2050
rect 36991 2004 37037 2050
rect 37107 2004 37153 2050
rect 37223 2004 37269 2050
rect 37339 2004 37385 2050
rect 37455 2004 37501 2050
rect 37571 2004 37617 2050
rect 37687 2004 37733 2050
rect 37803 2004 37849 2050
rect 37919 2004 37965 2050
rect 38035 2004 38081 2050
rect 38151 2004 38197 2050
rect 38267 2004 38313 2050
rect 38383 2004 38429 2050
rect 38499 2004 38545 2050
rect 38615 2004 38661 2050
rect 38731 2004 38777 2050
rect 38847 2004 38893 2050
rect 38963 2004 39009 2050
rect 39079 2004 39125 2050
rect 39195 2004 39241 2050
rect 39311 2004 39357 2050
rect 39427 2004 39473 2050
rect 39543 2004 39589 2050
rect 39659 2004 39705 2050
rect 39775 2004 39821 2050
rect 39891 2004 39937 2050
rect 40007 2004 40053 2050
rect 40123 2004 40169 2050
rect 28639 1888 28685 1934
rect 28755 1888 28801 1934
rect 28871 1888 28917 1934
rect 28987 1888 29033 1934
rect 29103 1888 29149 1934
rect 29219 1888 29265 1934
rect 29335 1888 29381 1934
rect 29451 1888 29497 1934
rect 29567 1888 29613 1934
rect 29683 1888 29729 1934
rect 29799 1888 29845 1934
rect 29915 1888 29961 1934
rect 30031 1888 30077 1934
rect 30147 1888 30193 1934
rect 30263 1888 30309 1934
rect 30379 1888 30425 1934
rect 30495 1888 30541 1934
rect 30611 1888 30657 1934
rect 30727 1888 30773 1934
rect 30843 1888 30889 1934
rect 30959 1888 31005 1934
rect 31075 1888 31121 1934
rect 31191 1888 31237 1934
rect 31307 1888 31353 1934
rect 31423 1888 31469 1934
rect 31539 1888 31585 1934
rect 31655 1888 31701 1934
rect 31771 1888 31817 1934
rect 31887 1888 31933 1934
rect 32003 1888 32049 1934
rect 32119 1888 32165 1934
rect 32235 1888 32281 1934
rect 32351 1888 32397 1934
rect 32467 1888 32513 1934
rect 32583 1888 32629 1934
rect 32699 1888 32745 1934
rect 32815 1888 32861 1934
rect 32931 1888 32977 1934
rect 33047 1888 33093 1934
rect 33163 1888 33209 1934
rect 33279 1888 33325 1934
rect 33395 1888 33441 1934
rect 33511 1888 33557 1934
rect 33627 1888 33673 1934
rect 33743 1888 33789 1934
rect 33859 1888 33905 1934
rect 33975 1888 34021 1934
rect 34091 1888 34137 1934
rect 34207 1888 34253 1934
rect 34323 1888 34369 1934
rect 34439 1888 34485 1934
rect 34555 1888 34601 1934
rect 34671 1888 34717 1934
rect 34787 1888 34833 1934
rect 34903 1888 34949 1934
rect 35019 1888 35065 1934
rect 35135 1888 35181 1934
rect 35251 1888 35297 1934
rect 35367 1888 35413 1934
rect 35483 1888 35529 1934
rect 35599 1888 35645 1934
rect 35715 1888 35761 1934
rect 35831 1888 35877 1934
rect 35947 1888 35993 1934
rect 36063 1888 36109 1934
rect 36179 1888 36225 1934
rect 36295 1888 36341 1934
rect 36411 1888 36457 1934
rect 36527 1888 36573 1934
rect 36643 1888 36689 1934
rect 36759 1888 36805 1934
rect 36875 1888 36921 1934
rect 36991 1888 37037 1934
rect 37107 1888 37153 1934
rect 37223 1888 37269 1934
rect 37339 1888 37385 1934
rect 37455 1888 37501 1934
rect 37571 1888 37617 1934
rect 37687 1888 37733 1934
rect 37803 1888 37849 1934
rect 37919 1888 37965 1934
rect 38035 1888 38081 1934
rect 38151 1888 38197 1934
rect 38267 1888 38313 1934
rect 38383 1888 38429 1934
rect 38499 1888 38545 1934
rect 38615 1888 38661 1934
rect 38731 1888 38777 1934
rect 38847 1888 38893 1934
rect 38963 1888 39009 1934
rect 39079 1888 39125 1934
rect 39195 1888 39241 1934
rect 39311 1888 39357 1934
rect 39427 1888 39473 1934
rect 39543 1888 39589 1934
rect 39659 1888 39705 1934
rect 39775 1888 39821 1934
rect 39891 1888 39937 1934
rect 40007 1888 40053 1934
rect 40123 1888 40169 1934
rect 28639 1772 28685 1818
rect 28755 1772 28801 1818
rect 28871 1772 28917 1818
rect 28987 1772 29033 1818
rect 29103 1772 29149 1818
rect 29219 1772 29265 1818
rect 29335 1772 29381 1818
rect 29451 1772 29497 1818
rect 29567 1772 29613 1818
rect 29683 1772 29729 1818
rect 29799 1772 29845 1818
rect 29915 1772 29961 1818
rect 30031 1772 30077 1818
rect 30147 1772 30193 1818
rect 30263 1772 30309 1818
rect 30379 1772 30425 1818
rect 30495 1772 30541 1818
rect 30611 1772 30657 1818
rect 30727 1772 30773 1818
rect 30843 1772 30889 1818
rect 30959 1772 31005 1818
rect 31075 1772 31121 1818
rect 31191 1772 31237 1818
rect 31307 1772 31353 1818
rect 31423 1772 31469 1818
rect 31539 1772 31585 1818
rect 31655 1772 31701 1818
rect 31771 1772 31817 1818
rect 31887 1772 31933 1818
rect 32003 1772 32049 1818
rect 32119 1772 32165 1818
rect 32235 1772 32281 1818
rect 32351 1772 32397 1818
rect 32467 1772 32513 1818
rect 32583 1772 32629 1818
rect 32699 1772 32745 1818
rect 32815 1772 32861 1818
rect 32931 1772 32977 1818
rect 33047 1772 33093 1818
rect 33163 1772 33209 1818
rect 33279 1772 33325 1818
rect 33395 1772 33441 1818
rect 33511 1772 33557 1818
rect 33627 1772 33673 1818
rect 33743 1772 33789 1818
rect 33859 1772 33905 1818
rect 33975 1772 34021 1818
rect 34091 1772 34137 1818
rect 34207 1772 34253 1818
rect 34323 1772 34369 1818
rect 34439 1772 34485 1818
rect 34555 1772 34601 1818
rect 34671 1772 34717 1818
rect 34787 1772 34833 1818
rect 34903 1772 34949 1818
rect 35019 1772 35065 1818
rect 35135 1772 35181 1818
rect 35251 1772 35297 1818
rect 35367 1772 35413 1818
rect 35483 1772 35529 1818
rect 35599 1772 35645 1818
rect 35715 1772 35761 1818
rect 35831 1772 35877 1818
rect 35947 1772 35993 1818
rect 36063 1772 36109 1818
rect 36179 1772 36225 1818
rect 36295 1772 36341 1818
rect 36411 1772 36457 1818
rect 36527 1772 36573 1818
rect 36643 1772 36689 1818
rect 36759 1772 36805 1818
rect 36875 1772 36921 1818
rect 36991 1772 37037 1818
rect 37107 1772 37153 1818
rect 37223 1772 37269 1818
rect 37339 1772 37385 1818
rect 37455 1772 37501 1818
rect 37571 1772 37617 1818
rect 37687 1772 37733 1818
rect 37803 1772 37849 1818
rect 37919 1772 37965 1818
rect 38035 1772 38081 1818
rect 38151 1772 38197 1818
rect 38267 1772 38313 1818
rect 38383 1772 38429 1818
rect 38499 1772 38545 1818
rect 38615 1772 38661 1818
rect 38731 1772 38777 1818
rect 38847 1772 38893 1818
rect 38963 1772 39009 1818
rect 39079 1772 39125 1818
rect 39195 1772 39241 1818
rect 39311 1772 39357 1818
rect 39427 1772 39473 1818
rect 39543 1772 39589 1818
rect 39659 1772 39705 1818
rect 39775 1772 39821 1818
rect 39891 1772 39937 1818
rect 40007 1772 40053 1818
rect 40123 1772 40169 1818
rect 28639 1656 28685 1702
rect 28755 1656 28801 1702
rect 28871 1656 28917 1702
rect 28987 1656 29033 1702
rect 29103 1656 29149 1702
rect 29219 1656 29265 1702
rect 29335 1656 29381 1702
rect 29451 1656 29497 1702
rect 29567 1656 29613 1702
rect 29683 1656 29729 1702
rect 29799 1656 29845 1702
rect 29915 1656 29961 1702
rect 30031 1656 30077 1702
rect 30147 1656 30193 1702
rect 30263 1656 30309 1702
rect 30379 1656 30425 1702
rect 30495 1656 30541 1702
rect 30611 1656 30657 1702
rect 30727 1656 30773 1702
rect 30843 1656 30889 1702
rect 30959 1656 31005 1702
rect 31075 1656 31121 1702
rect 31191 1656 31237 1702
rect 31307 1656 31353 1702
rect 31423 1656 31469 1702
rect 31539 1656 31585 1702
rect 31655 1656 31701 1702
rect 31771 1656 31817 1702
rect 31887 1656 31933 1702
rect 32003 1656 32049 1702
rect 32119 1656 32165 1702
rect 32235 1656 32281 1702
rect 32351 1656 32397 1702
rect 32467 1656 32513 1702
rect 32583 1656 32629 1702
rect 32699 1656 32745 1702
rect 32815 1656 32861 1702
rect 32931 1656 32977 1702
rect 33047 1656 33093 1702
rect 33163 1656 33209 1702
rect 33279 1656 33325 1702
rect 33395 1656 33441 1702
rect 33511 1656 33557 1702
rect 33627 1656 33673 1702
rect 33743 1656 33789 1702
rect 33859 1656 33905 1702
rect 33975 1656 34021 1702
rect 34091 1656 34137 1702
rect 34207 1656 34253 1702
rect 34323 1656 34369 1702
rect 34439 1656 34485 1702
rect 34555 1656 34601 1702
rect 34671 1656 34717 1702
rect 34787 1656 34833 1702
rect 34903 1656 34949 1702
rect 35019 1656 35065 1702
rect 35135 1656 35181 1702
rect 35251 1656 35297 1702
rect 35367 1656 35413 1702
rect 35483 1656 35529 1702
rect 35599 1656 35645 1702
rect 35715 1656 35761 1702
rect 35831 1656 35877 1702
rect 35947 1656 35993 1702
rect 36063 1656 36109 1702
rect 36179 1656 36225 1702
rect 36295 1656 36341 1702
rect 36411 1656 36457 1702
rect 36527 1656 36573 1702
rect 36643 1656 36689 1702
rect 36759 1656 36805 1702
rect 36875 1656 36921 1702
rect 36991 1656 37037 1702
rect 37107 1656 37153 1702
rect 37223 1656 37269 1702
rect 37339 1656 37385 1702
rect 37455 1656 37501 1702
rect 37571 1656 37617 1702
rect 37687 1656 37733 1702
rect 37803 1656 37849 1702
rect 37919 1656 37965 1702
rect 38035 1656 38081 1702
rect 38151 1656 38197 1702
rect 38267 1656 38313 1702
rect 38383 1656 38429 1702
rect 38499 1656 38545 1702
rect 38615 1656 38661 1702
rect 38731 1656 38777 1702
rect 38847 1656 38893 1702
rect 38963 1656 39009 1702
rect 39079 1656 39125 1702
rect 39195 1656 39241 1702
rect 39311 1656 39357 1702
rect 39427 1656 39473 1702
rect 39543 1656 39589 1702
rect 39659 1656 39705 1702
rect 39775 1656 39821 1702
rect 39891 1656 39937 1702
rect 40007 1656 40053 1702
rect 40123 1656 40169 1702
rect 50845 3860 50891 3906
rect 50961 3860 51007 3906
rect 51077 3860 51123 3906
rect 51193 3860 51239 3906
rect 51309 3860 51355 3906
rect 51425 3860 51471 3906
rect 51541 3860 51587 3906
rect 51657 3860 51703 3906
rect 51773 3860 51819 3906
rect 51889 3860 51935 3906
rect 52005 3860 52051 3906
rect 52121 3860 52167 3906
rect 52237 3860 52283 3906
rect 52353 3860 52399 3906
rect 52469 3860 52515 3906
rect 52585 3860 52631 3906
rect 52701 3860 52747 3906
rect 52817 3860 52863 3906
rect 52933 3860 52979 3906
rect 53049 3860 53095 3906
rect 53165 3860 53211 3906
rect 53281 3860 53327 3906
rect 53397 3860 53443 3906
rect 53513 3860 53559 3906
rect 53629 3860 53675 3906
rect 53745 3860 53791 3906
rect 53861 3860 53907 3906
rect 53977 3860 54023 3906
rect 54093 3860 54139 3906
rect 54209 3860 54255 3906
rect 54325 3860 54371 3906
rect 54441 3860 54487 3906
rect 54557 3860 54603 3906
rect 54673 3860 54719 3906
rect 54789 3860 54835 3906
rect 54905 3860 54951 3906
rect 55021 3860 55067 3906
rect 55137 3860 55183 3906
rect 55253 3860 55299 3906
rect 55369 3860 55415 3906
rect 55485 3860 55531 3906
rect 55601 3860 55647 3906
rect 55717 3860 55763 3906
rect 55833 3860 55879 3906
rect 55949 3860 55995 3906
rect 56065 3860 56111 3906
rect 56181 3860 56227 3906
rect 56297 3860 56343 3906
rect 56413 3860 56459 3906
rect 56529 3860 56575 3906
rect 50845 3744 50891 3790
rect 50961 3744 51007 3790
rect 51077 3744 51123 3790
rect 51193 3744 51239 3790
rect 51309 3744 51355 3790
rect 51425 3744 51471 3790
rect 51541 3744 51587 3790
rect 51657 3744 51703 3790
rect 51773 3744 51819 3790
rect 51889 3744 51935 3790
rect 52005 3744 52051 3790
rect 52121 3744 52167 3790
rect 52237 3744 52283 3790
rect 52353 3744 52399 3790
rect 52469 3744 52515 3790
rect 52585 3744 52631 3790
rect 52701 3744 52747 3790
rect 52817 3744 52863 3790
rect 52933 3744 52979 3790
rect 53049 3744 53095 3790
rect 53165 3744 53211 3790
rect 53281 3744 53327 3790
rect 53397 3744 53443 3790
rect 53513 3744 53559 3790
rect 53629 3744 53675 3790
rect 53745 3744 53791 3790
rect 53861 3744 53907 3790
rect 53977 3744 54023 3790
rect 54093 3744 54139 3790
rect 54209 3744 54255 3790
rect 54325 3744 54371 3790
rect 54441 3744 54487 3790
rect 54557 3744 54603 3790
rect 54673 3744 54719 3790
rect 54789 3744 54835 3790
rect 54905 3744 54951 3790
rect 55021 3744 55067 3790
rect 55137 3744 55183 3790
rect 55253 3744 55299 3790
rect 55369 3744 55415 3790
rect 55485 3744 55531 3790
rect 55601 3744 55647 3790
rect 55717 3744 55763 3790
rect 55833 3744 55879 3790
rect 55949 3744 55995 3790
rect 56065 3744 56111 3790
rect 56181 3744 56227 3790
rect 56297 3744 56343 3790
rect 56413 3744 56459 3790
rect 56529 3744 56575 3790
rect 50845 3628 50891 3674
rect 50961 3628 51007 3674
rect 51077 3628 51123 3674
rect 51193 3628 51239 3674
rect 51309 3628 51355 3674
rect 51425 3628 51471 3674
rect 51541 3628 51587 3674
rect 51657 3628 51703 3674
rect 51773 3628 51819 3674
rect 51889 3628 51935 3674
rect 52005 3628 52051 3674
rect 52121 3628 52167 3674
rect 52237 3628 52283 3674
rect 52353 3628 52399 3674
rect 52469 3628 52515 3674
rect 52585 3628 52631 3674
rect 52701 3628 52747 3674
rect 52817 3628 52863 3674
rect 52933 3628 52979 3674
rect 53049 3628 53095 3674
rect 53165 3628 53211 3674
rect 53281 3628 53327 3674
rect 53397 3628 53443 3674
rect 53513 3628 53559 3674
rect 53629 3628 53675 3674
rect 53745 3628 53791 3674
rect 53861 3628 53907 3674
rect 53977 3628 54023 3674
rect 54093 3628 54139 3674
rect 54209 3628 54255 3674
rect 54325 3628 54371 3674
rect 54441 3628 54487 3674
rect 54557 3628 54603 3674
rect 54673 3628 54719 3674
rect 54789 3628 54835 3674
rect 54905 3628 54951 3674
rect 55021 3628 55067 3674
rect 55137 3628 55183 3674
rect 55253 3628 55299 3674
rect 55369 3628 55415 3674
rect 55485 3628 55531 3674
rect 55601 3628 55647 3674
rect 55717 3628 55763 3674
rect 55833 3628 55879 3674
rect 55949 3628 55995 3674
rect 56065 3628 56111 3674
rect 56181 3628 56227 3674
rect 56297 3628 56343 3674
rect 56413 3628 56459 3674
rect 56529 3628 56575 3674
rect 50845 3512 50891 3558
rect 50961 3512 51007 3558
rect 51077 3512 51123 3558
rect 51193 3512 51239 3558
rect 51309 3512 51355 3558
rect 51425 3512 51471 3558
rect 51541 3512 51587 3558
rect 51657 3512 51703 3558
rect 51773 3512 51819 3558
rect 51889 3512 51935 3558
rect 52005 3512 52051 3558
rect 52121 3512 52167 3558
rect 52237 3512 52283 3558
rect 52353 3512 52399 3558
rect 52469 3512 52515 3558
rect 52585 3512 52631 3558
rect 52701 3512 52747 3558
rect 52817 3512 52863 3558
rect 52933 3512 52979 3558
rect 53049 3512 53095 3558
rect 53165 3512 53211 3558
rect 53281 3512 53327 3558
rect 53397 3512 53443 3558
rect 53513 3512 53559 3558
rect 53629 3512 53675 3558
rect 53745 3512 53791 3558
rect 53861 3512 53907 3558
rect 53977 3512 54023 3558
rect 54093 3512 54139 3558
rect 54209 3512 54255 3558
rect 54325 3512 54371 3558
rect 54441 3512 54487 3558
rect 54557 3512 54603 3558
rect 54673 3512 54719 3558
rect 54789 3512 54835 3558
rect 54905 3512 54951 3558
rect 55021 3512 55067 3558
rect 55137 3512 55183 3558
rect 55253 3512 55299 3558
rect 55369 3512 55415 3558
rect 55485 3512 55531 3558
rect 55601 3512 55647 3558
rect 55717 3512 55763 3558
rect 55833 3512 55879 3558
rect 55949 3512 55995 3558
rect 56065 3512 56111 3558
rect 56181 3512 56227 3558
rect 56297 3512 56343 3558
rect 56413 3512 56459 3558
rect 56529 3512 56575 3558
rect 50845 3396 50891 3442
rect 50961 3396 51007 3442
rect 51077 3396 51123 3442
rect 51193 3396 51239 3442
rect 51309 3396 51355 3442
rect 51425 3396 51471 3442
rect 51541 3396 51587 3442
rect 51657 3396 51703 3442
rect 51773 3396 51819 3442
rect 51889 3396 51935 3442
rect 52005 3396 52051 3442
rect 52121 3396 52167 3442
rect 52237 3396 52283 3442
rect 52353 3396 52399 3442
rect 52469 3396 52515 3442
rect 52585 3396 52631 3442
rect 52701 3396 52747 3442
rect 52817 3396 52863 3442
rect 52933 3396 52979 3442
rect 53049 3396 53095 3442
rect 53165 3396 53211 3442
rect 53281 3396 53327 3442
rect 53397 3396 53443 3442
rect 53513 3396 53559 3442
rect 53629 3396 53675 3442
rect 53745 3396 53791 3442
rect 53861 3396 53907 3442
rect 53977 3396 54023 3442
rect 54093 3396 54139 3442
rect 54209 3396 54255 3442
rect 54325 3396 54371 3442
rect 54441 3396 54487 3442
rect 54557 3396 54603 3442
rect 54673 3396 54719 3442
rect 54789 3396 54835 3442
rect 54905 3396 54951 3442
rect 55021 3396 55067 3442
rect 55137 3396 55183 3442
rect 55253 3396 55299 3442
rect 55369 3396 55415 3442
rect 55485 3396 55531 3442
rect 55601 3396 55647 3442
rect 55717 3396 55763 3442
rect 55833 3396 55879 3442
rect 55949 3396 55995 3442
rect 56065 3396 56111 3442
rect 56181 3396 56227 3442
rect 56297 3396 56343 3442
rect 56413 3396 56459 3442
rect 56529 3396 56575 3442
rect 50845 3280 50891 3326
rect 50961 3280 51007 3326
rect 51077 3280 51123 3326
rect 51193 3280 51239 3326
rect 51309 3280 51355 3326
rect 51425 3280 51471 3326
rect 51541 3280 51587 3326
rect 51657 3280 51703 3326
rect 51773 3280 51819 3326
rect 51889 3280 51935 3326
rect 52005 3280 52051 3326
rect 52121 3280 52167 3326
rect 52237 3280 52283 3326
rect 52353 3280 52399 3326
rect 52469 3280 52515 3326
rect 52585 3280 52631 3326
rect 52701 3280 52747 3326
rect 52817 3280 52863 3326
rect 52933 3280 52979 3326
rect 53049 3280 53095 3326
rect 53165 3280 53211 3326
rect 53281 3280 53327 3326
rect 53397 3280 53443 3326
rect 53513 3280 53559 3326
rect 53629 3280 53675 3326
rect 53745 3280 53791 3326
rect 53861 3280 53907 3326
rect 53977 3280 54023 3326
rect 54093 3280 54139 3326
rect 54209 3280 54255 3326
rect 54325 3280 54371 3326
rect 54441 3280 54487 3326
rect 54557 3280 54603 3326
rect 54673 3280 54719 3326
rect 54789 3280 54835 3326
rect 54905 3280 54951 3326
rect 55021 3280 55067 3326
rect 55137 3280 55183 3326
rect 55253 3280 55299 3326
rect 55369 3280 55415 3326
rect 55485 3280 55531 3326
rect 55601 3280 55647 3326
rect 55717 3280 55763 3326
rect 55833 3280 55879 3326
rect 55949 3280 55995 3326
rect 56065 3280 56111 3326
rect 56181 3280 56227 3326
rect 56297 3280 56343 3326
rect 56413 3280 56459 3326
rect 56529 3280 56575 3326
rect 50845 3164 50891 3210
rect 50961 3164 51007 3210
rect 51077 3164 51123 3210
rect 51193 3164 51239 3210
rect 51309 3164 51355 3210
rect 51425 3164 51471 3210
rect 51541 3164 51587 3210
rect 51657 3164 51703 3210
rect 51773 3164 51819 3210
rect 51889 3164 51935 3210
rect 52005 3164 52051 3210
rect 52121 3164 52167 3210
rect 52237 3164 52283 3210
rect 52353 3164 52399 3210
rect 52469 3164 52515 3210
rect 52585 3164 52631 3210
rect 52701 3164 52747 3210
rect 52817 3164 52863 3210
rect 52933 3164 52979 3210
rect 53049 3164 53095 3210
rect 53165 3164 53211 3210
rect 53281 3164 53327 3210
rect 53397 3164 53443 3210
rect 53513 3164 53559 3210
rect 53629 3164 53675 3210
rect 53745 3164 53791 3210
rect 53861 3164 53907 3210
rect 53977 3164 54023 3210
rect 54093 3164 54139 3210
rect 54209 3164 54255 3210
rect 54325 3164 54371 3210
rect 54441 3164 54487 3210
rect 54557 3164 54603 3210
rect 54673 3164 54719 3210
rect 54789 3164 54835 3210
rect 54905 3164 54951 3210
rect 55021 3164 55067 3210
rect 55137 3164 55183 3210
rect 55253 3164 55299 3210
rect 55369 3164 55415 3210
rect 55485 3164 55531 3210
rect 55601 3164 55647 3210
rect 55717 3164 55763 3210
rect 55833 3164 55879 3210
rect 55949 3164 55995 3210
rect 56065 3164 56111 3210
rect 56181 3164 56227 3210
rect 56297 3164 56343 3210
rect 56413 3164 56459 3210
rect 56529 3164 56575 3210
rect 50845 3048 50891 3094
rect 50961 3048 51007 3094
rect 51077 3048 51123 3094
rect 51193 3048 51239 3094
rect 51309 3048 51355 3094
rect 51425 3048 51471 3094
rect 51541 3048 51587 3094
rect 51657 3048 51703 3094
rect 51773 3048 51819 3094
rect 51889 3048 51935 3094
rect 52005 3048 52051 3094
rect 52121 3048 52167 3094
rect 52237 3048 52283 3094
rect 52353 3048 52399 3094
rect 52469 3048 52515 3094
rect 52585 3048 52631 3094
rect 52701 3048 52747 3094
rect 52817 3048 52863 3094
rect 52933 3048 52979 3094
rect 53049 3048 53095 3094
rect 53165 3048 53211 3094
rect 53281 3048 53327 3094
rect 53397 3048 53443 3094
rect 53513 3048 53559 3094
rect 53629 3048 53675 3094
rect 53745 3048 53791 3094
rect 53861 3048 53907 3094
rect 53977 3048 54023 3094
rect 54093 3048 54139 3094
rect 54209 3048 54255 3094
rect 54325 3048 54371 3094
rect 54441 3048 54487 3094
rect 54557 3048 54603 3094
rect 54673 3048 54719 3094
rect 54789 3048 54835 3094
rect 54905 3048 54951 3094
rect 55021 3048 55067 3094
rect 55137 3048 55183 3094
rect 55253 3048 55299 3094
rect 55369 3048 55415 3094
rect 55485 3048 55531 3094
rect 55601 3048 55647 3094
rect 55717 3048 55763 3094
rect 55833 3048 55879 3094
rect 55949 3048 55995 3094
rect 56065 3048 56111 3094
rect 56181 3048 56227 3094
rect 56297 3048 56343 3094
rect 56413 3048 56459 3094
rect 56529 3048 56575 3094
rect 50845 2932 50891 2978
rect 50961 2932 51007 2978
rect 51077 2932 51123 2978
rect 51193 2932 51239 2978
rect 51309 2932 51355 2978
rect 51425 2932 51471 2978
rect 51541 2932 51587 2978
rect 51657 2932 51703 2978
rect 51773 2932 51819 2978
rect 51889 2932 51935 2978
rect 52005 2932 52051 2978
rect 52121 2932 52167 2978
rect 52237 2932 52283 2978
rect 52353 2932 52399 2978
rect 52469 2932 52515 2978
rect 52585 2932 52631 2978
rect 52701 2932 52747 2978
rect 52817 2932 52863 2978
rect 52933 2932 52979 2978
rect 53049 2932 53095 2978
rect 53165 2932 53211 2978
rect 53281 2932 53327 2978
rect 53397 2932 53443 2978
rect 53513 2932 53559 2978
rect 53629 2932 53675 2978
rect 53745 2932 53791 2978
rect 53861 2932 53907 2978
rect 53977 2932 54023 2978
rect 54093 2932 54139 2978
rect 54209 2932 54255 2978
rect 54325 2932 54371 2978
rect 54441 2932 54487 2978
rect 54557 2932 54603 2978
rect 54673 2932 54719 2978
rect 54789 2932 54835 2978
rect 54905 2932 54951 2978
rect 55021 2932 55067 2978
rect 55137 2932 55183 2978
rect 55253 2932 55299 2978
rect 55369 2932 55415 2978
rect 55485 2932 55531 2978
rect 55601 2932 55647 2978
rect 55717 2932 55763 2978
rect 55833 2932 55879 2978
rect 55949 2932 55995 2978
rect 56065 2932 56111 2978
rect 56181 2932 56227 2978
rect 56297 2932 56343 2978
rect 56413 2932 56459 2978
rect 56529 2932 56575 2978
rect 50845 2816 50891 2862
rect 50961 2816 51007 2862
rect 51077 2816 51123 2862
rect 51193 2816 51239 2862
rect 51309 2816 51355 2862
rect 51425 2816 51471 2862
rect 51541 2816 51587 2862
rect 51657 2816 51703 2862
rect 51773 2816 51819 2862
rect 51889 2816 51935 2862
rect 52005 2816 52051 2862
rect 52121 2816 52167 2862
rect 52237 2816 52283 2862
rect 52353 2816 52399 2862
rect 52469 2816 52515 2862
rect 52585 2816 52631 2862
rect 52701 2816 52747 2862
rect 52817 2816 52863 2862
rect 52933 2816 52979 2862
rect 53049 2816 53095 2862
rect 53165 2816 53211 2862
rect 53281 2816 53327 2862
rect 53397 2816 53443 2862
rect 53513 2816 53559 2862
rect 53629 2816 53675 2862
rect 53745 2816 53791 2862
rect 53861 2816 53907 2862
rect 53977 2816 54023 2862
rect 54093 2816 54139 2862
rect 54209 2816 54255 2862
rect 54325 2816 54371 2862
rect 54441 2816 54487 2862
rect 54557 2816 54603 2862
rect 54673 2816 54719 2862
rect 54789 2816 54835 2862
rect 54905 2816 54951 2862
rect 55021 2816 55067 2862
rect 55137 2816 55183 2862
rect 55253 2816 55299 2862
rect 55369 2816 55415 2862
rect 55485 2816 55531 2862
rect 55601 2816 55647 2862
rect 55717 2816 55763 2862
rect 55833 2816 55879 2862
rect 55949 2816 55995 2862
rect 56065 2816 56111 2862
rect 56181 2816 56227 2862
rect 56297 2816 56343 2862
rect 56413 2816 56459 2862
rect 56529 2816 56575 2862
rect 50845 2700 50891 2746
rect 50961 2700 51007 2746
rect 51077 2700 51123 2746
rect 51193 2700 51239 2746
rect 51309 2700 51355 2746
rect 51425 2700 51471 2746
rect 51541 2700 51587 2746
rect 51657 2700 51703 2746
rect 51773 2700 51819 2746
rect 51889 2700 51935 2746
rect 52005 2700 52051 2746
rect 52121 2700 52167 2746
rect 52237 2700 52283 2746
rect 52353 2700 52399 2746
rect 52469 2700 52515 2746
rect 52585 2700 52631 2746
rect 52701 2700 52747 2746
rect 52817 2700 52863 2746
rect 52933 2700 52979 2746
rect 53049 2700 53095 2746
rect 53165 2700 53211 2746
rect 53281 2700 53327 2746
rect 53397 2700 53443 2746
rect 53513 2700 53559 2746
rect 53629 2700 53675 2746
rect 53745 2700 53791 2746
rect 53861 2700 53907 2746
rect 53977 2700 54023 2746
rect 54093 2700 54139 2746
rect 54209 2700 54255 2746
rect 54325 2700 54371 2746
rect 54441 2700 54487 2746
rect 54557 2700 54603 2746
rect 54673 2700 54719 2746
rect 54789 2700 54835 2746
rect 54905 2700 54951 2746
rect 55021 2700 55067 2746
rect 55137 2700 55183 2746
rect 55253 2700 55299 2746
rect 55369 2700 55415 2746
rect 55485 2700 55531 2746
rect 55601 2700 55647 2746
rect 55717 2700 55763 2746
rect 55833 2700 55879 2746
rect 55949 2700 55995 2746
rect 56065 2700 56111 2746
rect 56181 2700 56227 2746
rect 56297 2700 56343 2746
rect 56413 2700 56459 2746
rect 56529 2700 56575 2746
rect 50845 2584 50891 2630
rect 50961 2584 51007 2630
rect 51077 2584 51123 2630
rect 51193 2584 51239 2630
rect 51309 2584 51355 2630
rect 51425 2584 51471 2630
rect 51541 2584 51587 2630
rect 51657 2584 51703 2630
rect 51773 2584 51819 2630
rect 51889 2584 51935 2630
rect 52005 2584 52051 2630
rect 52121 2584 52167 2630
rect 52237 2584 52283 2630
rect 52353 2584 52399 2630
rect 52469 2584 52515 2630
rect 52585 2584 52631 2630
rect 52701 2584 52747 2630
rect 52817 2584 52863 2630
rect 52933 2584 52979 2630
rect 53049 2584 53095 2630
rect 53165 2584 53211 2630
rect 53281 2584 53327 2630
rect 53397 2584 53443 2630
rect 53513 2584 53559 2630
rect 53629 2584 53675 2630
rect 53745 2584 53791 2630
rect 53861 2584 53907 2630
rect 53977 2584 54023 2630
rect 54093 2584 54139 2630
rect 54209 2584 54255 2630
rect 54325 2584 54371 2630
rect 54441 2584 54487 2630
rect 54557 2584 54603 2630
rect 54673 2584 54719 2630
rect 54789 2584 54835 2630
rect 54905 2584 54951 2630
rect 55021 2584 55067 2630
rect 55137 2584 55183 2630
rect 55253 2584 55299 2630
rect 55369 2584 55415 2630
rect 55485 2584 55531 2630
rect 55601 2584 55647 2630
rect 55717 2584 55763 2630
rect 55833 2584 55879 2630
rect 55949 2584 55995 2630
rect 56065 2584 56111 2630
rect 56181 2584 56227 2630
rect 56297 2584 56343 2630
rect 56413 2584 56459 2630
rect 56529 2584 56575 2630
rect 50845 2468 50891 2514
rect 50961 2468 51007 2514
rect 51077 2468 51123 2514
rect 51193 2468 51239 2514
rect 51309 2468 51355 2514
rect 51425 2468 51471 2514
rect 51541 2468 51587 2514
rect 51657 2468 51703 2514
rect 51773 2468 51819 2514
rect 51889 2468 51935 2514
rect 52005 2468 52051 2514
rect 52121 2468 52167 2514
rect 52237 2468 52283 2514
rect 52353 2468 52399 2514
rect 52469 2468 52515 2514
rect 52585 2468 52631 2514
rect 52701 2468 52747 2514
rect 52817 2468 52863 2514
rect 52933 2468 52979 2514
rect 53049 2468 53095 2514
rect 53165 2468 53211 2514
rect 53281 2468 53327 2514
rect 53397 2468 53443 2514
rect 53513 2468 53559 2514
rect 53629 2468 53675 2514
rect 53745 2468 53791 2514
rect 53861 2468 53907 2514
rect 53977 2468 54023 2514
rect 54093 2468 54139 2514
rect 54209 2468 54255 2514
rect 54325 2468 54371 2514
rect 54441 2468 54487 2514
rect 54557 2468 54603 2514
rect 54673 2468 54719 2514
rect 54789 2468 54835 2514
rect 54905 2468 54951 2514
rect 55021 2468 55067 2514
rect 55137 2468 55183 2514
rect 55253 2468 55299 2514
rect 55369 2468 55415 2514
rect 55485 2468 55531 2514
rect 55601 2468 55647 2514
rect 55717 2468 55763 2514
rect 55833 2468 55879 2514
rect 55949 2468 55995 2514
rect 56065 2468 56111 2514
rect 56181 2468 56227 2514
rect 56297 2468 56343 2514
rect 56413 2468 56459 2514
rect 56529 2468 56575 2514
rect 50845 2352 50891 2398
rect 50961 2352 51007 2398
rect 51077 2352 51123 2398
rect 51193 2352 51239 2398
rect 51309 2352 51355 2398
rect 51425 2352 51471 2398
rect 51541 2352 51587 2398
rect 51657 2352 51703 2398
rect 51773 2352 51819 2398
rect 51889 2352 51935 2398
rect 52005 2352 52051 2398
rect 52121 2352 52167 2398
rect 52237 2352 52283 2398
rect 52353 2352 52399 2398
rect 52469 2352 52515 2398
rect 52585 2352 52631 2398
rect 52701 2352 52747 2398
rect 52817 2352 52863 2398
rect 52933 2352 52979 2398
rect 53049 2352 53095 2398
rect 53165 2352 53211 2398
rect 53281 2352 53327 2398
rect 53397 2352 53443 2398
rect 53513 2352 53559 2398
rect 53629 2352 53675 2398
rect 53745 2352 53791 2398
rect 53861 2352 53907 2398
rect 53977 2352 54023 2398
rect 54093 2352 54139 2398
rect 54209 2352 54255 2398
rect 54325 2352 54371 2398
rect 54441 2352 54487 2398
rect 54557 2352 54603 2398
rect 54673 2352 54719 2398
rect 54789 2352 54835 2398
rect 54905 2352 54951 2398
rect 55021 2352 55067 2398
rect 55137 2352 55183 2398
rect 55253 2352 55299 2398
rect 55369 2352 55415 2398
rect 55485 2352 55531 2398
rect 55601 2352 55647 2398
rect 55717 2352 55763 2398
rect 55833 2352 55879 2398
rect 55949 2352 55995 2398
rect 56065 2352 56111 2398
rect 56181 2352 56227 2398
rect 56297 2352 56343 2398
rect 56413 2352 56459 2398
rect 56529 2352 56575 2398
rect 50845 2236 50891 2282
rect 50961 2236 51007 2282
rect 51077 2236 51123 2282
rect 51193 2236 51239 2282
rect 51309 2236 51355 2282
rect 51425 2236 51471 2282
rect 51541 2236 51587 2282
rect 51657 2236 51703 2282
rect 51773 2236 51819 2282
rect 51889 2236 51935 2282
rect 52005 2236 52051 2282
rect 52121 2236 52167 2282
rect 52237 2236 52283 2282
rect 52353 2236 52399 2282
rect 52469 2236 52515 2282
rect 52585 2236 52631 2282
rect 52701 2236 52747 2282
rect 52817 2236 52863 2282
rect 52933 2236 52979 2282
rect 53049 2236 53095 2282
rect 53165 2236 53211 2282
rect 53281 2236 53327 2282
rect 53397 2236 53443 2282
rect 53513 2236 53559 2282
rect 53629 2236 53675 2282
rect 53745 2236 53791 2282
rect 53861 2236 53907 2282
rect 53977 2236 54023 2282
rect 54093 2236 54139 2282
rect 54209 2236 54255 2282
rect 54325 2236 54371 2282
rect 54441 2236 54487 2282
rect 54557 2236 54603 2282
rect 54673 2236 54719 2282
rect 54789 2236 54835 2282
rect 54905 2236 54951 2282
rect 55021 2236 55067 2282
rect 55137 2236 55183 2282
rect 55253 2236 55299 2282
rect 55369 2236 55415 2282
rect 55485 2236 55531 2282
rect 55601 2236 55647 2282
rect 55717 2236 55763 2282
rect 55833 2236 55879 2282
rect 55949 2236 55995 2282
rect 56065 2236 56111 2282
rect 56181 2236 56227 2282
rect 56297 2236 56343 2282
rect 56413 2236 56459 2282
rect 56529 2236 56575 2282
rect 50845 2120 50891 2166
rect 50961 2120 51007 2166
rect 51077 2120 51123 2166
rect 51193 2120 51239 2166
rect 51309 2120 51355 2166
rect 51425 2120 51471 2166
rect 51541 2120 51587 2166
rect 51657 2120 51703 2166
rect 51773 2120 51819 2166
rect 51889 2120 51935 2166
rect 52005 2120 52051 2166
rect 52121 2120 52167 2166
rect 52237 2120 52283 2166
rect 52353 2120 52399 2166
rect 52469 2120 52515 2166
rect 52585 2120 52631 2166
rect 52701 2120 52747 2166
rect 52817 2120 52863 2166
rect 52933 2120 52979 2166
rect 53049 2120 53095 2166
rect 53165 2120 53211 2166
rect 53281 2120 53327 2166
rect 53397 2120 53443 2166
rect 53513 2120 53559 2166
rect 53629 2120 53675 2166
rect 53745 2120 53791 2166
rect 53861 2120 53907 2166
rect 53977 2120 54023 2166
rect 54093 2120 54139 2166
rect 54209 2120 54255 2166
rect 54325 2120 54371 2166
rect 54441 2120 54487 2166
rect 54557 2120 54603 2166
rect 54673 2120 54719 2166
rect 54789 2120 54835 2166
rect 54905 2120 54951 2166
rect 55021 2120 55067 2166
rect 55137 2120 55183 2166
rect 55253 2120 55299 2166
rect 55369 2120 55415 2166
rect 55485 2120 55531 2166
rect 55601 2120 55647 2166
rect 55717 2120 55763 2166
rect 55833 2120 55879 2166
rect 55949 2120 55995 2166
rect 56065 2120 56111 2166
rect 56181 2120 56227 2166
rect 56297 2120 56343 2166
rect 56413 2120 56459 2166
rect 56529 2120 56575 2166
rect 50845 2004 50891 2050
rect 50961 2004 51007 2050
rect 51077 2004 51123 2050
rect 51193 2004 51239 2050
rect 51309 2004 51355 2050
rect 51425 2004 51471 2050
rect 51541 2004 51587 2050
rect 51657 2004 51703 2050
rect 51773 2004 51819 2050
rect 51889 2004 51935 2050
rect 52005 2004 52051 2050
rect 52121 2004 52167 2050
rect 52237 2004 52283 2050
rect 52353 2004 52399 2050
rect 52469 2004 52515 2050
rect 52585 2004 52631 2050
rect 52701 2004 52747 2050
rect 52817 2004 52863 2050
rect 52933 2004 52979 2050
rect 53049 2004 53095 2050
rect 53165 2004 53211 2050
rect 53281 2004 53327 2050
rect 53397 2004 53443 2050
rect 53513 2004 53559 2050
rect 53629 2004 53675 2050
rect 53745 2004 53791 2050
rect 53861 2004 53907 2050
rect 53977 2004 54023 2050
rect 54093 2004 54139 2050
rect 54209 2004 54255 2050
rect 54325 2004 54371 2050
rect 54441 2004 54487 2050
rect 54557 2004 54603 2050
rect 54673 2004 54719 2050
rect 54789 2004 54835 2050
rect 54905 2004 54951 2050
rect 55021 2004 55067 2050
rect 55137 2004 55183 2050
rect 55253 2004 55299 2050
rect 55369 2004 55415 2050
rect 55485 2004 55531 2050
rect 55601 2004 55647 2050
rect 55717 2004 55763 2050
rect 55833 2004 55879 2050
rect 55949 2004 55995 2050
rect 56065 2004 56111 2050
rect 56181 2004 56227 2050
rect 56297 2004 56343 2050
rect 56413 2004 56459 2050
rect 56529 2004 56575 2050
rect 50845 1888 50891 1934
rect 50961 1888 51007 1934
rect 51077 1888 51123 1934
rect 51193 1888 51239 1934
rect 51309 1888 51355 1934
rect 51425 1888 51471 1934
rect 51541 1888 51587 1934
rect 51657 1888 51703 1934
rect 51773 1888 51819 1934
rect 51889 1888 51935 1934
rect 52005 1888 52051 1934
rect 52121 1888 52167 1934
rect 52237 1888 52283 1934
rect 52353 1888 52399 1934
rect 52469 1888 52515 1934
rect 52585 1888 52631 1934
rect 52701 1888 52747 1934
rect 52817 1888 52863 1934
rect 52933 1888 52979 1934
rect 53049 1888 53095 1934
rect 53165 1888 53211 1934
rect 53281 1888 53327 1934
rect 53397 1888 53443 1934
rect 53513 1888 53559 1934
rect 53629 1888 53675 1934
rect 53745 1888 53791 1934
rect 53861 1888 53907 1934
rect 53977 1888 54023 1934
rect 54093 1888 54139 1934
rect 54209 1888 54255 1934
rect 54325 1888 54371 1934
rect 54441 1888 54487 1934
rect 54557 1888 54603 1934
rect 54673 1888 54719 1934
rect 54789 1888 54835 1934
rect 54905 1888 54951 1934
rect 55021 1888 55067 1934
rect 55137 1888 55183 1934
rect 55253 1888 55299 1934
rect 55369 1888 55415 1934
rect 55485 1888 55531 1934
rect 55601 1888 55647 1934
rect 55717 1888 55763 1934
rect 55833 1888 55879 1934
rect 55949 1888 55995 1934
rect 56065 1888 56111 1934
rect 56181 1888 56227 1934
rect 56297 1888 56343 1934
rect 56413 1888 56459 1934
rect 56529 1888 56575 1934
rect 50845 1772 50891 1818
rect 50961 1772 51007 1818
rect 51077 1772 51123 1818
rect 51193 1772 51239 1818
rect 51309 1772 51355 1818
rect 51425 1772 51471 1818
rect 51541 1772 51587 1818
rect 51657 1772 51703 1818
rect 51773 1772 51819 1818
rect 51889 1772 51935 1818
rect 52005 1772 52051 1818
rect 52121 1772 52167 1818
rect 52237 1772 52283 1818
rect 52353 1772 52399 1818
rect 52469 1772 52515 1818
rect 52585 1772 52631 1818
rect 52701 1772 52747 1818
rect 52817 1772 52863 1818
rect 52933 1772 52979 1818
rect 53049 1772 53095 1818
rect 53165 1772 53211 1818
rect 53281 1772 53327 1818
rect 53397 1772 53443 1818
rect 53513 1772 53559 1818
rect 53629 1772 53675 1818
rect 53745 1772 53791 1818
rect 53861 1772 53907 1818
rect 53977 1772 54023 1818
rect 54093 1772 54139 1818
rect 54209 1772 54255 1818
rect 54325 1772 54371 1818
rect 54441 1772 54487 1818
rect 54557 1772 54603 1818
rect 54673 1772 54719 1818
rect 54789 1772 54835 1818
rect 54905 1772 54951 1818
rect 55021 1772 55067 1818
rect 55137 1772 55183 1818
rect 55253 1772 55299 1818
rect 55369 1772 55415 1818
rect 55485 1772 55531 1818
rect 55601 1772 55647 1818
rect 55717 1772 55763 1818
rect 55833 1772 55879 1818
rect 55949 1772 55995 1818
rect 56065 1772 56111 1818
rect 56181 1772 56227 1818
rect 56297 1772 56343 1818
rect 56413 1772 56459 1818
rect 56529 1772 56575 1818
rect 50845 1656 50891 1702
rect 50961 1656 51007 1702
rect 51077 1656 51123 1702
rect 51193 1656 51239 1702
rect 51309 1656 51355 1702
rect 51425 1656 51471 1702
rect 51541 1656 51587 1702
rect 51657 1656 51703 1702
rect 51773 1656 51819 1702
rect 51889 1656 51935 1702
rect 52005 1656 52051 1702
rect 52121 1656 52167 1702
rect 52237 1656 52283 1702
rect 52353 1656 52399 1702
rect 52469 1656 52515 1702
rect 52585 1656 52631 1702
rect 52701 1656 52747 1702
rect 52817 1656 52863 1702
rect 52933 1656 52979 1702
rect 53049 1656 53095 1702
rect 53165 1656 53211 1702
rect 53281 1656 53327 1702
rect 53397 1656 53443 1702
rect 53513 1656 53559 1702
rect 53629 1656 53675 1702
rect 53745 1656 53791 1702
rect 53861 1656 53907 1702
rect 53977 1656 54023 1702
rect 54093 1656 54139 1702
rect 54209 1656 54255 1702
rect 54325 1656 54371 1702
rect 54441 1656 54487 1702
rect 54557 1656 54603 1702
rect 54673 1656 54719 1702
rect 54789 1656 54835 1702
rect 54905 1656 54951 1702
rect 55021 1656 55067 1702
rect 55137 1656 55183 1702
rect 55253 1656 55299 1702
rect 55369 1656 55415 1702
rect 55485 1656 55531 1702
rect 55601 1656 55647 1702
rect 55717 1656 55763 1702
rect 55833 1656 55879 1702
rect 55949 1656 55995 1702
rect 56065 1656 56111 1702
rect 56181 1656 56227 1702
rect 56297 1656 56343 1702
rect 56413 1656 56459 1702
rect 56529 1656 56575 1702
rect 57380 1117 57626 52963
<< metal1 >>
rect 27387 52963 28911 53137
rect 25313 51579 26039 52644
rect 25313 51527 25400 51579
rect 25452 51527 25524 51579
rect 25576 51527 25648 51579
rect 25700 51527 25772 51579
rect 25824 51527 25896 51579
rect 25948 51527 26039 51579
rect 25313 51455 26039 51527
rect 25313 51403 25400 51455
rect 25452 51403 25524 51455
rect 25576 51403 25648 51455
rect 25700 51403 25772 51455
rect 25824 51403 25896 51455
rect 25948 51403 26039 51455
rect 25313 51331 26039 51403
rect 25313 51279 25400 51331
rect 25452 51279 25524 51331
rect 25576 51279 25648 51331
rect 25700 51279 25772 51331
rect 25824 51279 25896 51331
rect 25948 51279 26039 51331
rect 25313 51195 26039 51279
rect 27387 35273 27498 52963
rect 27744 52942 28911 52963
rect 27744 51453 27846 52942
rect 28492 51526 28911 52942
rect 28492 51494 28757 51526
rect 28492 51453 29146 51494
rect 27744 51401 27790 51453
rect 27842 51401 27846 51453
rect 28492 51401 28634 51453
rect 28686 51401 28845 51453
rect 28897 51401 29056 51453
rect 29108 51401 29146 51453
rect 27744 49653 27846 51401
rect 28492 51360 29146 51401
rect 28492 49694 28757 51360
rect 50636 51285 51451 52995
rect 55927 52974 57369 53223
rect 55927 52963 57637 52974
rect 55927 52942 57380 52963
rect 55927 51453 56632 52942
rect 57278 51453 57380 52942
rect 55927 51401 56015 51453
rect 56067 51401 56226 51453
rect 56278 51401 56437 51453
rect 56489 51401 56632 51453
rect 57278 51401 57281 51453
rect 57333 51401 57380 51453
rect 28492 49653 29146 49694
rect 27744 49601 27790 49653
rect 27842 49601 27846 49653
rect 28492 49601 28634 49653
rect 28686 49601 28845 49653
rect 28897 49601 29056 49653
rect 29108 49601 29146 49653
rect 27744 47853 27846 49601
rect 28492 49560 29146 49601
rect 55927 49653 56632 51401
rect 57278 49653 57380 51401
rect 55927 49601 56015 49653
rect 56067 49601 56226 49653
rect 56278 49601 56437 49653
rect 56489 49601 56632 49653
rect 57278 49601 57281 49653
rect 57333 49601 57380 49653
rect 28492 47894 28757 49560
rect 28492 47853 29146 47894
rect 27744 47801 27790 47853
rect 27842 47801 27846 47853
rect 28492 47801 28634 47853
rect 28686 47801 28845 47853
rect 28897 47801 29056 47853
rect 29108 47801 29146 47853
rect 27744 46053 27846 47801
rect 28492 47760 29146 47801
rect 55927 47853 56632 49601
rect 57278 47853 57380 49601
rect 55927 47801 56015 47853
rect 56067 47801 56226 47853
rect 56278 47801 56437 47853
rect 56489 47801 56632 47853
rect 57278 47801 57281 47853
rect 57333 47801 57380 47853
rect 28492 46094 28757 47760
rect 28492 46053 29146 46094
rect 27744 46001 27790 46053
rect 27842 46001 27846 46053
rect 28492 46001 28634 46053
rect 28686 46001 28845 46053
rect 28897 46001 29056 46053
rect 29108 46001 29146 46053
rect 27744 44253 27846 46001
rect 28492 45960 29146 46001
rect 55927 46053 56632 47801
rect 57278 46053 57380 47801
rect 55927 46001 56015 46053
rect 56067 46001 56226 46053
rect 56278 46001 56437 46053
rect 56489 46001 56632 46053
rect 57278 46001 57281 46053
rect 57333 46001 57380 46053
rect 28492 44294 28757 45960
rect 28492 44253 29146 44294
rect 27744 44201 27790 44253
rect 27842 44201 27846 44253
rect 28492 44201 28634 44253
rect 28686 44201 28845 44253
rect 28897 44201 29056 44253
rect 29108 44201 29146 44253
rect 27744 42453 27846 44201
rect 28492 44160 29146 44201
rect 55927 44253 56632 46001
rect 57278 44253 57380 46001
rect 55927 44201 56015 44253
rect 56067 44201 56226 44253
rect 56278 44201 56437 44253
rect 56489 44201 56632 44253
rect 57278 44201 57281 44253
rect 57333 44201 57380 44253
rect 28492 42494 28757 44160
rect 28492 42453 29146 42494
rect 27744 42401 27790 42453
rect 27842 42401 27846 42453
rect 28492 42401 28634 42453
rect 28686 42401 28845 42453
rect 28897 42401 29056 42453
rect 29108 42401 29146 42453
rect 27744 40653 27846 42401
rect 28492 42360 29146 42401
rect 55927 42453 56632 44201
rect 57278 42453 57380 44201
rect 55927 42401 56015 42453
rect 56067 42401 56226 42453
rect 56278 42401 56437 42453
rect 56489 42401 56632 42453
rect 57278 42401 57281 42453
rect 57333 42401 57380 42453
rect 28492 40694 28757 42360
rect 28492 40653 29146 40694
rect 27744 40601 27790 40653
rect 27842 40601 27846 40653
rect 28492 40601 28634 40653
rect 28686 40601 28845 40653
rect 28897 40601 29056 40653
rect 29108 40601 29146 40653
rect 27744 38853 27846 40601
rect 28492 40560 29146 40601
rect 55927 40653 56632 42401
rect 57278 40653 57380 42401
rect 55927 40601 56015 40653
rect 56067 40601 56226 40653
rect 56278 40601 56437 40653
rect 56489 40601 56632 40653
rect 57278 40601 57281 40653
rect 57333 40601 57380 40653
rect 28492 38894 28757 40560
rect 28492 38853 29146 38894
rect 27744 38801 27790 38853
rect 27842 38801 27846 38853
rect 28492 38801 28634 38853
rect 28686 38801 28845 38853
rect 28897 38801 29056 38853
rect 29108 38801 29146 38853
rect 27744 37053 27846 38801
rect 28492 38760 29146 38801
rect 55927 38853 56632 40601
rect 57278 38853 57380 40601
rect 55927 38801 56015 38853
rect 56067 38801 56226 38853
rect 56278 38801 56437 38853
rect 56489 38801 56632 38853
rect 57278 38801 57281 38853
rect 57333 38801 57380 38853
rect 28492 37094 28757 38760
rect 28492 37053 29146 37094
rect 27744 37001 27790 37053
rect 27842 37001 27846 37053
rect 28492 37001 28634 37053
rect 28686 37001 28845 37053
rect 28897 37001 29056 37053
rect 29108 37001 29146 37053
rect 27744 35996 27846 37001
rect 28492 36960 29146 37001
rect 55927 37053 56632 38801
rect 57278 37053 57380 38801
rect 55927 37001 56015 37053
rect 56067 37001 56226 37053
rect 56278 37001 56437 37053
rect 56489 37001 56632 37053
rect 57278 37001 57281 37053
rect 57333 37001 57380 37053
rect 28492 35996 28757 36960
rect 27744 35985 28757 35996
rect 55927 35996 56632 37001
rect 57278 35996 57380 37001
rect 55927 35985 57380 35996
rect 27387 35221 27440 35273
rect 27492 35221 27498 35273
rect 27387 35149 27498 35221
rect 27387 35097 27440 35149
rect 27492 35097 27498 35149
rect 27387 35025 27498 35097
rect 27387 34973 27440 35025
rect 27492 34973 27498 35025
rect 27387 34901 27498 34973
rect 27387 34849 27440 34901
rect 27492 34849 27498 34901
rect 27387 34777 27498 34849
rect 27387 34725 27440 34777
rect 27492 34725 27498 34777
rect 27387 34653 27498 34725
rect 27387 34601 27440 34653
rect 27492 34601 27498 34653
rect 27744 34613 27828 35985
rect 27744 34602 57303 34613
rect 26772 33432 27214 33519
rect 26772 33380 26861 33432
rect 26913 33380 27073 33432
rect 27125 33380 27214 33432
rect 26772 33215 27214 33380
rect 26772 33163 26861 33215
rect 26913 33163 27073 33215
rect 27125 33163 27214 33215
rect 26772 32997 27214 33163
rect 26772 32945 26861 32997
rect 26913 32945 27073 32997
rect 27125 32945 27214 32997
rect 26772 32779 27214 32945
rect 26772 32727 26861 32779
rect 26913 32727 27073 32779
rect 27125 32727 27214 32779
rect 26772 32562 27214 32727
rect 26772 32510 26861 32562
rect 26913 32510 27073 32562
rect 27125 32510 27214 32562
rect 26772 32344 27214 32510
rect 26772 32292 26861 32344
rect 26913 32292 27073 32344
rect 27125 32292 27214 32344
rect 26772 32127 27214 32292
rect 26772 32075 26861 32127
rect 26913 32075 27073 32127
rect 27125 32075 27214 32127
rect 26772 31909 27214 32075
rect 26772 31857 26861 31909
rect 26913 31857 27073 31909
rect 27125 31857 27214 31909
rect 26772 31691 27214 31857
rect 26772 31639 26861 31691
rect 26913 31639 27073 31691
rect 27125 31639 27214 31691
rect 26772 31474 27214 31639
rect 26772 31422 26861 31474
rect 26913 31422 27073 31474
rect 27125 31422 27214 31474
rect 26772 31256 27214 31422
rect 26772 31204 26861 31256
rect 26913 31204 27073 31256
rect 27125 31204 27214 31256
rect 26772 31038 27214 31204
rect 26772 30986 26861 31038
rect 26913 30986 27073 31038
rect 27125 30986 27214 31038
rect 26772 30821 27214 30986
rect 26772 30769 26861 30821
rect 26913 30769 27073 30821
rect 27125 30769 27214 30821
rect 26772 30603 27214 30769
rect 26772 30551 26861 30603
rect 26913 30551 27073 30603
rect 27125 30551 27214 30603
rect 26772 30386 27214 30551
rect 26772 30334 26861 30386
rect 26913 30334 27073 30386
rect 27125 30334 27214 30386
rect 26772 30168 27214 30334
rect 26772 30116 26861 30168
rect 26913 30116 27073 30168
rect 27125 30116 27214 30168
rect 26772 29950 27214 30116
rect 26772 29898 26861 29950
rect 26913 29898 27073 29950
rect 27125 29898 27214 29950
rect 26772 29733 27214 29898
rect 26772 29681 26861 29733
rect 26913 29681 27073 29733
rect 27125 29681 27214 29733
rect 26772 29515 27214 29681
rect 26772 29463 26861 29515
rect 26913 29463 27073 29515
rect 27125 29463 27214 29515
rect 26772 29297 27214 29463
rect 26772 29245 26861 29297
rect 26913 29245 27073 29297
rect 27125 29245 27214 29297
rect 26772 29080 27214 29245
rect 26772 29028 26861 29080
rect 26913 29028 27073 29080
rect 27125 29028 27214 29080
rect 26772 28862 27214 29028
rect 26772 28810 26861 28862
rect 26913 28810 27073 28862
rect 27125 28810 27214 28862
rect 26772 28644 27214 28810
rect 26772 28592 26861 28644
rect 26913 28592 27073 28644
rect 27125 28592 27214 28644
rect 26772 28427 27214 28592
rect 26772 28375 26861 28427
rect 26913 28375 27073 28427
rect 27125 28375 27214 28427
rect 26772 28209 27214 28375
rect 26772 28157 26861 28209
rect 26913 28157 27073 28209
rect 27125 28157 27214 28209
rect 26772 27992 27214 28157
rect 26772 27940 26861 27992
rect 26913 27940 27073 27992
rect 27125 27940 27214 27992
rect 26772 27774 27214 27940
rect 26772 27722 26861 27774
rect 26913 27722 27073 27774
rect 27125 27722 27214 27774
rect 26772 27556 27214 27722
rect 26772 27504 26861 27556
rect 26913 27504 27073 27556
rect 27125 27504 27214 27556
rect 26772 27339 27214 27504
rect 26772 27287 26861 27339
rect 26913 27287 27073 27339
rect 27125 27287 27214 27339
rect 26772 27121 27214 27287
rect 26772 27069 26861 27121
rect 26913 27069 27073 27121
rect 27125 27069 27214 27121
rect 26772 26903 27214 27069
rect 26772 26851 26861 26903
rect 26913 26851 27073 26903
rect 27125 26851 27214 26903
rect 26772 26686 27214 26851
rect 26772 26634 26861 26686
rect 26913 26634 27073 26686
rect 27125 26634 27214 26686
rect 26772 26468 27214 26634
rect 26772 26416 26861 26468
rect 26913 26416 27073 26468
rect 27125 26416 27214 26468
rect 26772 26250 27214 26416
rect 26772 26198 26861 26250
rect 26913 26198 27073 26250
rect 27125 26198 27214 26250
rect 26772 26033 27214 26198
rect 26772 25981 26861 26033
rect 26913 25981 27073 26033
rect 27125 25981 27214 26033
rect 26772 25815 27214 25981
rect 26772 25763 26861 25815
rect 26913 25763 27073 25815
rect 27125 25763 27214 25815
rect 26772 25598 27214 25763
rect 26772 25546 26861 25598
rect 26913 25546 27073 25598
rect 27125 25546 27214 25598
rect 26772 25380 27214 25546
rect 26772 25328 26861 25380
rect 26913 25328 27073 25380
rect 27125 25328 27214 25380
rect 26772 25162 27214 25328
rect 26772 25110 26861 25162
rect 26913 25110 27073 25162
rect 27125 25110 27214 25162
rect 26772 24945 27214 25110
rect 26772 24893 26861 24945
rect 26913 24893 27073 24945
rect 27125 24893 27214 24945
rect 26772 24727 27214 24893
rect 26772 24675 26861 24727
rect 26913 24675 27073 24727
rect 27125 24675 27214 24727
rect 26772 24509 27214 24675
rect 26772 24457 26861 24509
rect 26913 24457 27073 24509
rect 27125 24457 27214 24509
rect 26772 24292 27214 24457
rect 26772 24240 26861 24292
rect 26913 24240 27073 24292
rect 27125 24240 27214 24292
rect 26772 24074 27214 24240
rect 26772 24022 26861 24074
rect 26913 24022 27073 24074
rect 27125 24022 27214 24074
rect 26772 23857 27214 24022
rect 26772 23805 26861 23857
rect 26913 23805 27073 23857
rect 27125 23805 27214 23857
rect 26772 23639 27214 23805
rect 26772 23587 26861 23639
rect 26913 23587 27073 23639
rect 27125 23587 27214 23639
rect 26772 23421 27214 23587
rect 26772 23369 26861 23421
rect 26913 23369 27073 23421
rect 27125 23369 27214 23421
rect 26772 23204 27214 23369
rect 26772 23152 26861 23204
rect 26913 23152 27073 23204
rect 27125 23152 27214 23204
rect 26772 22986 27214 23152
rect 26772 22934 26861 22986
rect 26913 22934 27073 22986
rect 27125 22934 27214 22986
rect 26772 22768 27214 22934
rect 26772 22716 26861 22768
rect 26913 22716 27073 22768
rect 27125 22716 27214 22768
rect 26772 22551 27214 22716
rect 26772 22499 26861 22551
rect 26913 22499 27073 22551
rect 27125 22499 27214 22551
rect 26772 22333 27214 22499
rect 26772 22281 26861 22333
rect 26913 22281 27073 22333
rect 27125 22281 27214 22333
rect 26772 22115 27214 22281
rect 26772 22063 26861 22115
rect 26913 22063 27073 22115
rect 27125 22063 27214 22115
rect 26772 21898 27214 22063
rect 26772 21846 26861 21898
rect 26913 21846 27073 21898
rect 27125 21846 27214 21898
rect 26772 21680 27214 21846
rect 26772 21628 26861 21680
rect 26913 21628 27073 21680
rect 27125 21628 27214 21680
rect 26772 21463 27214 21628
rect 26772 21411 26861 21463
rect 26913 21411 27073 21463
rect 27125 21411 27214 21463
rect 26772 21245 27214 21411
rect 26772 21193 26861 21245
rect 26913 21193 27073 21245
rect 27125 21193 27214 21245
rect 26772 21027 27214 21193
rect 26772 20975 26861 21027
rect 26913 20975 27073 21027
rect 27125 20975 27214 21027
rect 26772 20810 27214 20975
rect 26772 20758 26861 20810
rect 26913 20758 27073 20810
rect 27125 20758 27214 20810
rect 26772 20592 27214 20758
rect 26772 20540 26861 20592
rect 26913 20540 27073 20592
rect 27125 20540 27214 20592
rect 26772 20374 27214 20540
rect 26772 20322 26861 20374
rect 26913 20322 27073 20374
rect 27125 20322 27214 20374
rect 26772 20157 27214 20322
rect 26772 20105 26861 20157
rect 26913 20105 27073 20157
rect 27125 20105 27214 20157
rect 26772 19939 27214 20105
rect 26772 19887 26861 19939
rect 26913 19887 27073 19939
rect 27125 19887 27214 19939
rect 26772 19722 27214 19887
rect 26772 19670 26861 19722
rect 26913 19670 27073 19722
rect 27125 19670 27214 19722
rect 26772 19504 27214 19670
rect 26772 19452 26861 19504
rect 26913 19452 27073 19504
rect 27125 19452 27214 19504
rect 26772 19286 27214 19452
rect 26772 19234 26861 19286
rect 26913 19234 27073 19286
rect 27125 19234 27214 19286
rect 26772 19068 27214 19234
rect 26772 19016 26861 19068
rect 26913 19016 27073 19068
rect 27125 19016 27214 19068
rect 26772 18851 27214 19016
rect 26772 18799 26861 18851
rect 26913 18799 27073 18851
rect 27125 18799 27214 18851
rect 26772 18633 27214 18799
rect 26772 18581 26861 18633
rect 26913 18581 27073 18633
rect 27125 18581 27214 18633
rect 26772 18416 27214 18581
rect 26772 18364 26861 18416
rect 26913 18364 27073 18416
rect 27125 18364 27214 18416
rect 26772 18198 27214 18364
rect 26772 18146 26861 18198
rect 26913 18146 27073 18198
rect 27125 18146 27214 18198
rect 26772 17980 27214 18146
rect 26772 17928 26861 17980
rect 26913 17928 27073 17980
rect 27125 17928 27214 17980
rect 26772 17763 27214 17928
rect 26772 17711 26861 17763
rect 26913 17711 27073 17763
rect 27125 17711 27214 17763
rect 26772 17545 27214 17711
rect 26772 17493 26861 17545
rect 26913 17493 27073 17545
rect 27125 17493 27214 17545
rect 26772 17327 27214 17493
rect 26772 17275 26861 17327
rect 26913 17275 27073 17327
rect 27125 17275 27214 17327
rect 26772 17110 27214 17275
rect 26772 17058 26861 17110
rect 26913 17058 27073 17110
rect 27125 17058 27214 17110
rect 26772 16892 27214 17058
rect 26772 16840 26861 16892
rect 26913 16840 27073 16892
rect 27125 16840 27214 16892
rect 26772 16675 27214 16840
rect 26772 16623 26861 16675
rect 26913 16623 27073 16675
rect 27125 16623 27214 16675
rect 26772 16457 27214 16623
rect 26772 16405 26861 16457
rect 26913 16405 27073 16457
rect 27125 16405 27214 16457
rect 26772 16239 27214 16405
rect 26772 16187 26861 16239
rect 26913 16187 27073 16239
rect 27125 16187 27214 16239
rect 26772 16022 27214 16187
rect 26772 15970 26861 16022
rect 26913 15970 27073 16022
rect 27125 15970 27214 16022
rect 26772 15804 27214 15970
rect 26772 15752 26861 15804
rect 26913 15752 27073 15804
rect 27125 15752 27214 15804
rect 26772 15586 27214 15752
rect 26772 15534 26861 15586
rect 26913 15534 27073 15586
rect 27125 15534 27214 15586
rect 26772 15369 27214 15534
rect 26772 15317 26861 15369
rect 26913 15317 27073 15369
rect 27125 15317 27214 15369
rect 26772 15151 27214 15317
rect 26772 15099 26861 15151
rect 26913 15099 27073 15151
rect 27125 15099 27214 15151
rect 26772 14933 27214 15099
rect 26772 14881 26861 14933
rect 26913 14881 27073 14933
rect 27125 14881 27214 14933
rect 26772 14716 27214 14881
rect 26772 14664 26861 14716
rect 26913 14664 27073 14716
rect 27125 14664 27214 14716
rect 26772 14498 27214 14664
rect 26772 14446 26861 14498
rect 26913 14446 27073 14498
rect 27125 14446 27214 14498
rect 26772 14281 27214 14446
rect 26772 14229 26861 14281
rect 26913 14229 27073 14281
rect 27125 14229 27214 14281
rect 26772 14063 27214 14229
rect 26772 14011 26861 14063
rect 26913 14011 27073 14063
rect 27125 14011 27214 14063
rect 26772 13845 27214 14011
rect 26772 13793 26861 13845
rect 26913 13793 27073 13845
rect 27125 13793 27214 13845
rect 26772 13628 27214 13793
rect 26772 13576 26861 13628
rect 26913 13576 27073 13628
rect 27125 13576 27214 13628
rect 26772 13410 27214 13576
rect 26772 13358 26861 13410
rect 26913 13358 27073 13410
rect 27125 13358 27214 13410
rect 26772 13192 27214 13358
rect 26772 13140 26861 13192
rect 26913 13140 27073 13192
rect 27125 13140 27214 13192
rect 26772 12975 27214 13140
rect 26772 12923 26861 12975
rect 26913 12923 27073 12975
rect 27125 12923 27214 12975
rect 26772 12757 27214 12923
rect 26772 12705 26861 12757
rect 26913 12705 27073 12757
rect 27125 12705 27214 12757
rect 26772 12540 27214 12705
rect 26772 12488 26861 12540
rect 26913 12488 27073 12540
rect 27125 12488 27214 12540
rect 26772 12322 27214 12488
rect 26772 12270 26861 12322
rect 26913 12270 27073 12322
rect 27125 12270 27214 12322
rect 26772 12104 27214 12270
rect 26772 12052 26861 12104
rect 26913 12052 27073 12104
rect 27125 12052 27214 12104
rect 26772 11887 27214 12052
rect 26772 11835 26861 11887
rect 26913 11835 27073 11887
rect 27125 11835 27214 11887
rect 26772 11669 27214 11835
rect 26772 11617 26861 11669
rect 26913 11617 27073 11669
rect 27125 11617 27214 11669
rect 26772 11451 27214 11617
rect 26772 11399 26861 11451
rect 26913 11399 27073 11451
rect 27125 11399 27214 11451
rect 26772 11234 27214 11399
rect 26772 11182 26861 11234
rect 26913 11182 27073 11234
rect 27125 11182 27214 11234
rect 26772 11016 27214 11182
rect 26772 10964 26861 11016
rect 26913 10964 27073 11016
rect 27125 10964 27214 11016
rect 26772 10798 27214 10964
rect 26772 10746 26861 10798
rect 26913 10746 27073 10798
rect 27125 10746 27214 10798
rect 26772 10581 27214 10746
rect 26772 10529 26861 10581
rect 26913 10529 27073 10581
rect 27125 10529 27214 10581
rect 26772 10363 27214 10529
rect 26772 10311 26861 10363
rect 26913 10311 27073 10363
rect 27125 10311 27214 10363
rect 26772 10146 27214 10311
rect 26772 10094 26861 10146
rect 26913 10094 27073 10146
rect 27125 10094 27214 10146
rect 26772 9928 27214 10094
rect 26772 9876 26861 9928
rect 26913 9876 27073 9928
rect 27125 9876 27214 9928
rect 26772 9710 27214 9876
rect 26772 9658 26861 9710
rect 26913 9658 27073 9710
rect 27125 9658 27214 9710
rect 26772 9493 27214 9658
rect 26772 9441 26861 9493
rect 26913 9441 27073 9493
rect 27125 9441 27214 9493
rect 26772 9275 27214 9441
rect 26772 9223 26861 9275
rect 26913 9223 27073 9275
rect 27125 9223 27214 9275
rect 26772 9057 27214 9223
rect 26772 9005 26861 9057
rect 26913 9005 27073 9057
rect 27125 9005 27214 9057
rect 26772 8840 27214 9005
rect 26772 8788 26861 8840
rect 26913 8788 27073 8840
rect 27125 8788 27214 8840
rect 26772 8622 27214 8788
rect 26772 8570 26861 8622
rect 26913 8570 27073 8622
rect 27125 8570 27214 8622
rect 26772 8404 27214 8570
rect 26772 8352 26861 8404
rect 26913 8352 27073 8404
rect 27125 8352 27214 8404
rect 26772 8187 27214 8352
rect 26772 8135 26861 8187
rect 26913 8135 27073 8187
rect 27125 8135 27214 8187
rect 26772 7969 27214 8135
rect 26772 7917 26861 7969
rect 26913 7917 27073 7969
rect 27125 7917 27214 7969
rect 26772 7752 27214 7917
rect 26772 7700 26861 7752
rect 26913 7700 27073 7752
rect 27125 7700 27214 7752
rect 26772 7534 27214 7700
rect 26772 7482 26861 7534
rect 26913 7482 27073 7534
rect 27125 7482 27214 7534
rect 26772 7316 27214 7482
rect 26772 7264 26861 7316
rect 26913 7264 27073 7316
rect 27125 7264 27214 7316
rect 26772 7099 27214 7264
rect 26772 7047 26861 7099
rect 26913 7047 27073 7099
rect 27125 7047 27214 7099
rect 26772 6881 27214 7047
rect 26772 6829 26861 6881
rect 26913 6829 27073 6881
rect 27125 6829 27214 6881
rect 26772 6663 27214 6829
rect 26772 6611 26861 6663
rect 26913 6611 27073 6663
rect 27125 6611 27214 6663
rect 26772 6446 27214 6611
rect 26772 6394 26861 6446
rect 26913 6394 27073 6446
rect 27125 6394 27214 6446
rect 26772 6228 27214 6394
rect 26772 6176 26861 6228
rect 26913 6176 27073 6228
rect 27125 6176 27214 6228
rect 26772 6011 27214 6176
rect 26772 5959 26861 6011
rect 26913 5959 27073 6011
rect 27125 5959 27214 6011
rect 26772 5793 27214 5959
rect 26772 5741 26861 5793
rect 26913 5741 27073 5793
rect 27125 5741 27214 5793
rect 26772 5575 27214 5741
rect 26772 5523 26861 5575
rect 26913 5523 27073 5575
rect 27125 5523 27214 5575
rect 26772 5358 27214 5523
rect 26772 5306 26861 5358
rect 26913 5306 27073 5358
rect 27125 5306 27214 5358
rect 26772 4587 27214 5306
rect 26772 4535 26861 4587
rect 26913 4535 27073 4587
rect 27125 4535 27214 4587
rect 26772 4370 27214 4535
rect 26772 4318 26861 4370
rect 26913 4318 27073 4370
rect 27125 4318 27214 4370
rect 26772 4152 27214 4318
rect 26772 4100 26861 4152
rect 26913 4100 27073 4152
rect 27125 4100 27214 4152
rect 26772 3934 27214 4100
rect 26772 3882 26861 3934
rect 26913 3882 27073 3934
rect 27125 3882 27214 3934
rect 26772 3717 27214 3882
rect 26772 3665 26861 3717
rect 26913 3665 27073 3717
rect 27125 3665 27214 3717
rect 26772 1777 27214 3665
rect 27387 33432 27498 34601
rect 27744 34256 27846 34602
rect 57292 34256 57303 34602
rect 27744 34245 57303 34256
rect 27387 33380 27476 33432
rect 27387 33215 27498 33380
rect 27387 33163 27476 33215
rect 27387 32997 27498 33163
rect 27387 32945 27476 32997
rect 27387 32779 27498 32945
rect 27387 32727 27476 32779
rect 27387 32562 27498 32727
rect 27387 32510 27476 32562
rect 27387 32344 27498 32510
rect 27387 32292 27476 32344
rect 27387 32127 27498 32292
rect 27387 32075 27476 32127
rect 27387 31909 27498 32075
rect 27387 31857 27476 31909
rect 27387 31691 27498 31857
rect 27387 31639 27476 31691
rect 27387 31474 27498 31639
rect 27387 31422 27476 31474
rect 27387 31256 27498 31422
rect 27387 31204 27476 31256
rect 27387 31038 27498 31204
rect 27387 30986 27476 31038
rect 27387 30821 27498 30986
rect 27387 30769 27476 30821
rect 27387 30603 27498 30769
rect 27387 30551 27476 30603
rect 27387 30386 27498 30551
rect 27387 30334 27476 30386
rect 27387 30168 27498 30334
rect 27387 30116 27476 30168
rect 27387 29950 27498 30116
rect 27387 29898 27476 29950
rect 27387 29733 27498 29898
rect 27387 29681 27476 29733
rect 27387 29515 27498 29681
rect 27387 29463 27476 29515
rect 27387 29297 27498 29463
rect 27387 29245 27476 29297
rect 27387 29080 27498 29245
rect 27387 29028 27476 29080
rect 27387 28862 27498 29028
rect 27387 28810 27476 28862
rect 27387 28644 27498 28810
rect 27387 28592 27476 28644
rect 27387 28427 27498 28592
rect 27387 28375 27476 28427
rect 27387 28209 27498 28375
rect 27387 28157 27476 28209
rect 27387 27992 27498 28157
rect 27387 27940 27476 27992
rect 27387 27774 27498 27940
rect 27387 27722 27476 27774
rect 27387 27556 27498 27722
rect 27387 27504 27476 27556
rect 27387 27339 27498 27504
rect 27387 27287 27476 27339
rect 27387 27121 27498 27287
rect 27387 27069 27476 27121
rect 27387 26903 27498 27069
rect 27387 26851 27476 26903
rect 27387 26686 27498 26851
rect 27387 26634 27476 26686
rect 27387 26468 27498 26634
rect 27387 26416 27476 26468
rect 27387 26250 27498 26416
rect 27387 26198 27476 26250
rect 27387 26033 27498 26198
rect 27387 25981 27476 26033
rect 27387 25815 27498 25981
rect 27387 25763 27476 25815
rect 27387 25598 27498 25763
rect 27387 25546 27476 25598
rect 27387 25380 27498 25546
rect 27387 25328 27476 25380
rect 27387 25162 27498 25328
rect 27387 25110 27476 25162
rect 27387 24945 27498 25110
rect 27387 24893 27476 24945
rect 27387 24727 27498 24893
rect 27387 24675 27476 24727
rect 27387 24509 27498 24675
rect 27387 24457 27476 24509
rect 27387 24292 27498 24457
rect 27387 24240 27476 24292
rect 27387 24074 27498 24240
rect 27387 24022 27476 24074
rect 27387 23857 27498 24022
rect 27387 23805 27476 23857
rect 27387 23639 27498 23805
rect 27387 23587 27476 23639
rect 27387 23421 27498 23587
rect 27387 23369 27476 23421
rect 27387 23204 27498 23369
rect 27387 23152 27476 23204
rect 27387 22986 27498 23152
rect 27387 22934 27476 22986
rect 27387 22768 27498 22934
rect 27387 22716 27476 22768
rect 27387 22551 27498 22716
rect 27387 22499 27476 22551
rect 27387 22333 27498 22499
rect 27387 22281 27476 22333
rect 27387 22115 27498 22281
rect 27387 22063 27476 22115
rect 27387 21898 27498 22063
rect 27387 21846 27476 21898
rect 27387 21680 27498 21846
rect 27387 21628 27476 21680
rect 27387 21463 27498 21628
rect 27387 21411 27476 21463
rect 27387 21245 27498 21411
rect 27387 21193 27476 21245
rect 27387 21027 27498 21193
rect 27387 20975 27476 21027
rect 27387 20810 27498 20975
rect 27387 20758 27476 20810
rect 27387 20592 27498 20758
rect 27387 20540 27476 20592
rect 27387 20374 27498 20540
rect 27387 20322 27476 20374
rect 27387 20157 27498 20322
rect 27387 20105 27476 20157
rect 27387 19939 27498 20105
rect 27387 19887 27476 19939
rect 27387 19722 27498 19887
rect 27387 19670 27476 19722
rect 27387 19504 27498 19670
rect 27387 19452 27476 19504
rect 27387 19286 27498 19452
rect 27387 19234 27476 19286
rect 27387 19068 27498 19234
rect 27387 19016 27476 19068
rect 27387 18851 27498 19016
rect 27387 18799 27476 18851
rect 27387 18633 27498 18799
rect 27387 18581 27476 18633
rect 27387 18416 27498 18581
rect 27387 18364 27476 18416
rect 27387 18198 27498 18364
rect 27387 18146 27476 18198
rect 27387 17980 27498 18146
rect 27387 17928 27476 17980
rect 27387 17763 27498 17928
rect 27387 17711 27476 17763
rect 27387 17545 27498 17711
rect 27387 17493 27476 17545
rect 27387 17327 27498 17493
rect 27387 17275 27476 17327
rect 27387 17110 27498 17275
rect 27387 17058 27476 17110
rect 27387 16892 27498 17058
rect 27387 16840 27476 16892
rect 27387 16675 27498 16840
rect 27387 16623 27476 16675
rect 27387 16457 27498 16623
rect 27387 16405 27476 16457
rect 27387 16239 27498 16405
rect 27387 16187 27476 16239
rect 27387 16022 27498 16187
rect 27387 15970 27476 16022
rect 27387 15804 27498 15970
rect 27387 15752 27476 15804
rect 27387 15586 27498 15752
rect 27387 15534 27476 15586
rect 27387 15369 27498 15534
rect 27387 15317 27476 15369
rect 27387 15151 27498 15317
rect 27387 15099 27476 15151
rect 27387 14933 27498 15099
rect 27387 14881 27476 14933
rect 27387 14716 27498 14881
rect 27387 14664 27476 14716
rect 27387 14498 27498 14664
rect 27387 14446 27476 14498
rect 27387 14281 27498 14446
rect 27387 14229 27476 14281
rect 27387 14063 27498 14229
rect 27387 14011 27476 14063
rect 27387 13845 27498 14011
rect 27387 13793 27476 13845
rect 27387 13628 27498 13793
rect 27387 13576 27476 13628
rect 27387 13410 27498 13576
rect 27387 13358 27476 13410
rect 27387 13192 27498 13358
rect 27387 13140 27476 13192
rect 27387 12975 27498 13140
rect 27387 12923 27476 12975
rect 27387 12757 27498 12923
rect 27387 12705 27476 12757
rect 27387 12540 27498 12705
rect 27387 12488 27476 12540
rect 27387 12322 27498 12488
rect 27387 12270 27476 12322
rect 27387 12104 27498 12270
rect 27387 12052 27476 12104
rect 27387 11887 27498 12052
rect 27387 11835 27476 11887
rect 27387 11669 27498 11835
rect 27387 11617 27476 11669
rect 27387 11451 27498 11617
rect 27387 11399 27476 11451
rect 27387 11234 27498 11399
rect 27387 11182 27476 11234
rect 27387 11016 27498 11182
rect 27387 10964 27476 11016
rect 27387 10798 27498 10964
rect 27387 10746 27476 10798
rect 27387 10581 27498 10746
rect 27387 10529 27476 10581
rect 27387 10363 27498 10529
rect 27387 10311 27476 10363
rect 27387 10146 27498 10311
rect 27387 10094 27476 10146
rect 27387 9928 27498 10094
rect 27387 9876 27476 9928
rect 27387 9710 27498 9876
rect 27387 9658 27476 9710
rect 27387 9493 27498 9658
rect 27387 9441 27476 9493
rect 27387 9275 27498 9441
rect 27387 9223 27476 9275
rect 27387 9057 27498 9223
rect 27387 9005 27476 9057
rect 27387 8840 27498 9005
rect 27387 8788 27476 8840
rect 27387 8622 27498 8788
rect 27387 8570 27476 8622
rect 27387 8404 27498 8570
rect 27387 8352 27476 8404
rect 27387 8187 27498 8352
rect 27387 8135 27476 8187
rect 27387 7969 27498 8135
rect 27387 7917 27476 7969
rect 27387 7752 27498 7917
rect 27387 7700 27476 7752
rect 27387 7534 27498 7700
rect 27387 7482 27476 7534
rect 27387 7316 27498 7482
rect 27387 7264 27476 7316
rect 27387 7099 27498 7264
rect 27387 7047 27476 7099
rect 27387 6881 27498 7047
rect 27387 6829 27476 6881
rect 27387 6663 27498 6829
rect 27387 6611 27476 6663
rect 27387 6446 27498 6611
rect 27387 6394 27476 6446
rect 27387 6228 27498 6394
rect 27387 6176 27476 6228
rect 27387 6011 27498 6176
rect 27387 5959 27476 6011
rect 27387 5793 27498 5959
rect 27387 5741 27476 5793
rect 27387 5575 27498 5741
rect 27387 5523 27476 5575
rect 27387 5358 27498 5523
rect 27387 5306 27476 5358
rect 27387 4587 27498 5306
rect 27387 4535 27476 4587
rect 27387 4370 27498 4535
rect 27387 4318 27476 4370
rect 27387 4152 27498 4318
rect 27387 4100 27476 4152
rect 27387 3934 27498 4100
rect 27387 3882 27476 3934
rect 27387 3717 27498 3882
rect 27387 3665 27476 3717
rect 2562 1689 2742 1701
rect 2562 1637 2574 1689
rect 2730 1637 2742 1689
rect 2562 1625 2742 1637
rect 12627 1689 12807 1701
rect 12627 1637 12639 1689
rect 12795 1637 12807 1689
rect 12627 1625 12807 1637
rect 13077 1689 13257 1701
rect 13077 1637 13089 1689
rect 13245 1637 13257 1689
rect 13077 1625 13257 1637
rect 23427 1689 23607 1701
rect 23427 1637 23439 1689
rect 23595 1637 23607 1689
rect 23427 1625 23607 1637
rect 27387 1282 27498 3665
rect 282 1117 27498 1282
rect 27744 1282 27828 34245
rect 57369 33519 57380 35985
rect 49896 6349 50076 6361
rect 49896 6347 49908 6349
rect 49728 6301 49908 6347
rect 49896 6297 49908 6301
rect 50064 6297 50076 6349
rect 49896 6285 50076 6297
rect 57295 5220 57380 33519
rect 57626 33519 57637 52963
rect 58791 51579 59517 52644
rect 58791 51527 58878 51579
rect 58930 51527 59002 51579
rect 59054 51527 59126 51579
rect 59178 51527 59250 51579
rect 59302 51527 59374 51579
rect 59426 51527 59517 51579
rect 58791 51455 59517 51527
rect 58791 51403 58878 51455
rect 58930 51403 59002 51455
rect 59054 51403 59126 51455
rect 59178 51403 59250 51455
rect 59302 51403 59374 51455
rect 59426 51403 59517 51455
rect 58791 51331 59517 51403
rect 58791 51279 58878 51331
rect 58930 51279 59002 51331
rect 59054 51279 59126 51331
rect 59178 51279 59250 51331
rect 59302 51279 59374 51331
rect 59426 51279 59517 51331
rect 58791 51258 59517 51279
rect 60563 35494 60639 35506
rect 60563 35338 60575 35494
rect 60627 35338 60639 35494
rect 60563 35326 60639 35338
rect 84369 35126 85931 35326
rect 85090 34536 85931 35126
rect 57626 33432 57736 33519
rect 57647 33380 57736 33432
rect 57626 33215 57736 33380
rect 57647 33163 57736 33215
rect 57626 32997 57736 33163
rect 57647 32945 57736 32997
rect 57626 32779 57736 32945
rect 57647 32727 57736 32779
rect 57626 32562 57736 32727
rect 57647 32510 57736 32562
rect 57626 32344 57736 32510
rect 57647 32292 57736 32344
rect 57626 32127 57736 32292
rect 57647 32075 57736 32127
rect 57626 31909 57736 32075
rect 57647 31857 57736 31909
rect 57626 31691 57736 31857
rect 57647 31639 57736 31691
rect 57626 31474 57736 31639
rect 57647 31422 57736 31474
rect 57626 31256 57736 31422
rect 57647 31204 57736 31256
rect 57626 31038 57736 31204
rect 57647 30986 57736 31038
rect 57626 30821 57736 30986
rect 57647 30769 57736 30821
rect 57626 30603 57736 30769
rect 57647 30551 57736 30603
rect 57626 30386 57736 30551
rect 57647 30334 57736 30386
rect 57626 30168 57736 30334
rect 57647 30116 57736 30168
rect 57626 29950 57736 30116
rect 57647 29898 57736 29950
rect 57626 29733 57736 29898
rect 57647 29681 57736 29733
rect 57626 29515 57736 29681
rect 57647 29463 57736 29515
rect 57626 29297 57736 29463
rect 57647 29245 57736 29297
rect 57626 29080 57736 29245
rect 57647 29028 57736 29080
rect 57626 28862 57736 29028
rect 57647 28810 57736 28862
rect 57626 28644 57736 28810
rect 57647 28592 57736 28644
rect 57626 28427 57736 28592
rect 57647 28375 57736 28427
rect 57626 28209 57736 28375
rect 57647 28157 57736 28209
rect 57626 27992 57736 28157
rect 57647 27940 57736 27992
rect 57626 27774 57736 27940
rect 57647 27722 57736 27774
rect 57626 27556 57736 27722
rect 57647 27504 57736 27556
rect 57626 27339 57736 27504
rect 57647 27287 57736 27339
rect 57626 27121 57736 27287
rect 57647 27069 57736 27121
rect 57626 26903 57736 27069
rect 57647 26851 57736 26903
rect 57626 26686 57736 26851
rect 57647 26634 57736 26686
rect 57626 26468 57736 26634
rect 57647 26416 57736 26468
rect 57626 26250 57736 26416
rect 57647 26198 57736 26250
rect 57626 26033 57736 26198
rect 57647 25981 57736 26033
rect 57626 25815 57736 25981
rect 57647 25763 57736 25815
rect 57626 25598 57736 25763
rect 57647 25546 57736 25598
rect 57626 25380 57736 25546
rect 57647 25328 57736 25380
rect 57626 25162 57736 25328
rect 57647 25110 57736 25162
rect 57626 24945 57736 25110
rect 57647 24893 57736 24945
rect 57626 24727 57736 24893
rect 57647 24675 57736 24727
rect 57626 24509 57736 24675
rect 57647 24457 57736 24509
rect 57626 24292 57736 24457
rect 57647 24240 57736 24292
rect 57626 24074 57736 24240
rect 57647 24022 57736 24074
rect 57626 23857 57736 24022
rect 57647 23805 57736 23857
rect 57626 23639 57736 23805
rect 57647 23587 57736 23639
rect 57626 23421 57736 23587
rect 57647 23369 57736 23421
rect 57626 23204 57736 23369
rect 57647 23152 57736 23204
rect 57626 22986 57736 23152
rect 57647 22934 57736 22986
rect 57626 22768 57736 22934
rect 57647 22716 57736 22768
rect 57626 22551 57736 22716
rect 57647 22499 57736 22551
rect 57626 22333 57736 22499
rect 57647 22281 57736 22333
rect 57626 22115 57736 22281
rect 57647 22063 57736 22115
rect 57626 21898 57736 22063
rect 57647 21846 57736 21898
rect 57626 21680 57736 21846
rect 57647 21628 57736 21680
rect 57626 21463 57736 21628
rect 57647 21411 57736 21463
rect 57626 21245 57736 21411
rect 57647 21193 57736 21245
rect 57626 21027 57736 21193
rect 57647 20975 57736 21027
rect 57626 20810 57736 20975
rect 57647 20758 57736 20810
rect 57626 20592 57736 20758
rect 57647 20540 57736 20592
rect 57626 20374 57736 20540
rect 57647 20322 57736 20374
rect 57626 20157 57736 20322
rect 57647 20105 57736 20157
rect 57626 19939 57736 20105
rect 57647 19887 57736 19939
rect 57626 19722 57736 19887
rect 57647 19670 57736 19722
rect 57626 19504 57736 19670
rect 57647 19452 57736 19504
rect 57626 19286 57736 19452
rect 57647 19234 57736 19286
rect 57626 19068 57736 19234
rect 57647 19016 57736 19068
rect 57626 18851 57736 19016
rect 57647 18799 57736 18851
rect 57626 18633 57736 18799
rect 57647 18581 57736 18633
rect 57626 18416 57736 18581
rect 57647 18364 57736 18416
rect 57626 18198 57736 18364
rect 57647 18146 57736 18198
rect 57626 17980 57736 18146
rect 57647 17928 57736 17980
rect 57626 17763 57736 17928
rect 57647 17711 57736 17763
rect 57626 17545 57736 17711
rect 57647 17493 57736 17545
rect 57626 17327 57736 17493
rect 57647 17275 57736 17327
rect 57626 17110 57736 17275
rect 57647 17058 57736 17110
rect 57626 16892 57736 17058
rect 57647 16840 57736 16892
rect 57626 16675 57736 16840
rect 57647 16623 57736 16675
rect 57626 16457 57736 16623
rect 57647 16405 57736 16457
rect 57626 16239 57736 16405
rect 57647 16187 57736 16239
rect 57626 16022 57736 16187
rect 57647 15970 57736 16022
rect 57626 15804 57736 15970
rect 57647 15752 57736 15804
rect 57626 15586 57736 15752
rect 57647 15534 57736 15586
rect 57626 15369 57736 15534
rect 57647 15317 57736 15369
rect 57626 15151 57736 15317
rect 57647 15099 57736 15151
rect 57626 14933 57736 15099
rect 57647 14881 57736 14933
rect 57626 14716 57736 14881
rect 57647 14664 57736 14716
rect 57626 14498 57736 14664
rect 57647 14446 57736 14498
rect 57626 14281 57736 14446
rect 57647 14229 57736 14281
rect 57626 14063 57736 14229
rect 57647 14011 57736 14063
rect 57626 13845 57736 14011
rect 57647 13793 57736 13845
rect 57626 13628 57736 13793
rect 57647 13576 57736 13628
rect 57626 13410 57736 13576
rect 57647 13358 57736 13410
rect 57626 13192 57736 13358
rect 57647 13140 57736 13192
rect 57626 12975 57736 13140
rect 57647 12923 57736 12975
rect 57626 12757 57736 12923
rect 57647 12705 57736 12757
rect 57626 12540 57736 12705
rect 57647 12488 57736 12540
rect 57626 12322 57736 12488
rect 57647 12270 57736 12322
rect 57626 12104 57736 12270
rect 57647 12052 57736 12104
rect 57626 11887 57736 12052
rect 57647 11835 57736 11887
rect 57626 11669 57736 11835
rect 57647 11617 57736 11669
rect 57626 11451 57736 11617
rect 57647 11399 57736 11451
rect 57626 11234 57736 11399
rect 57647 11182 57736 11234
rect 57626 11016 57736 11182
rect 57647 10964 57736 11016
rect 57626 10798 57736 10964
rect 57647 10746 57736 10798
rect 57626 10581 57736 10746
rect 57647 10529 57736 10581
rect 57626 10363 57736 10529
rect 57647 10311 57736 10363
rect 57626 10146 57736 10311
rect 57647 10094 57736 10146
rect 57626 9928 57736 10094
rect 57647 9876 57736 9928
rect 57626 9710 57736 9876
rect 57647 9658 57736 9710
rect 57626 9493 57736 9658
rect 57647 9441 57736 9493
rect 57626 9275 57736 9441
rect 57647 9223 57736 9275
rect 57626 9057 57736 9223
rect 57647 9005 57736 9057
rect 57626 8840 57736 9005
rect 57647 8788 57736 8840
rect 57626 8622 57736 8788
rect 57647 8570 57736 8622
rect 57626 8404 57736 8570
rect 57647 8352 57736 8404
rect 57626 8187 57736 8352
rect 57647 8135 57736 8187
rect 57626 7969 57736 8135
rect 57647 7917 57736 7969
rect 57626 7752 57736 7917
rect 57647 7700 57736 7752
rect 57626 7534 57736 7700
rect 57647 7482 57736 7534
rect 57626 7316 57736 7482
rect 57647 7264 57736 7316
rect 57626 7099 57736 7264
rect 57647 7047 57736 7099
rect 57626 6881 57736 7047
rect 57647 6829 57736 6881
rect 57626 6663 57736 6829
rect 57647 6611 57736 6663
rect 57626 6446 57736 6611
rect 57647 6394 57736 6446
rect 57626 6228 57736 6394
rect 57647 6176 57736 6228
rect 57626 6011 57736 6176
rect 57647 5959 57736 6011
rect 57626 5793 57736 5959
rect 57647 5741 57736 5793
rect 57626 5575 57736 5741
rect 57647 5523 57736 5575
rect 57626 5358 57736 5523
rect 57647 5306 57736 5358
rect 51642 5199 51822 5211
rect 51642 5196 51654 5199
rect 49963 5150 51654 5196
rect 51642 5147 51654 5150
rect 51810 5147 51822 5199
rect 51642 5135 51822 5147
rect 40610 4904 40790 4916
rect 40610 4852 40622 4904
rect 40778 4852 40790 4904
rect 40610 4840 40790 4852
rect 57369 4728 57380 5220
rect 28628 3906 40180 3917
rect 28628 3860 28639 3906
rect 28685 3860 28755 3906
rect 28801 3860 28871 3906
rect 28917 3860 28987 3906
rect 29033 3860 29103 3906
rect 29149 3860 29219 3906
rect 29265 3860 29335 3906
rect 29381 3860 29451 3906
rect 29497 3860 29567 3906
rect 29613 3860 29683 3906
rect 29729 3860 29799 3906
rect 29845 3860 29915 3906
rect 29961 3860 30031 3906
rect 30077 3860 30147 3906
rect 30193 3860 30263 3906
rect 30309 3860 30379 3906
rect 30425 3860 30495 3906
rect 30541 3860 30611 3906
rect 30657 3860 30727 3906
rect 30773 3860 30843 3906
rect 30889 3860 30959 3906
rect 31005 3860 31075 3906
rect 31121 3860 31191 3906
rect 31237 3860 31307 3906
rect 31353 3860 31423 3906
rect 31469 3860 31539 3906
rect 31585 3860 31655 3906
rect 31701 3860 31771 3906
rect 31817 3860 31887 3906
rect 31933 3860 32003 3906
rect 32049 3860 32119 3906
rect 32165 3860 32235 3906
rect 32281 3860 32351 3906
rect 32397 3860 32467 3906
rect 32513 3860 32583 3906
rect 32629 3860 32699 3906
rect 32745 3860 32815 3906
rect 32861 3860 32931 3906
rect 32977 3860 33047 3906
rect 33093 3860 33163 3906
rect 33209 3860 33279 3906
rect 33325 3860 33395 3906
rect 33441 3860 33511 3906
rect 33557 3860 33627 3906
rect 33673 3860 33743 3906
rect 33789 3860 33859 3906
rect 33905 3860 33975 3906
rect 34021 3860 34091 3906
rect 34137 3860 34207 3906
rect 34253 3860 34323 3906
rect 34369 3860 34439 3906
rect 34485 3860 34555 3906
rect 34601 3860 34671 3906
rect 34717 3860 34787 3906
rect 34833 3860 34903 3906
rect 34949 3860 35019 3906
rect 35065 3860 35135 3906
rect 35181 3860 35251 3906
rect 35297 3860 35367 3906
rect 35413 3860 35483 3906
rect 35529 3860 35599 3906
rect 35645 3860 35715 3906
rect 35761 3860 35831 3906
rect 35877 3860 35947 3906
rect 35993 3860 36063 3906
rect 36109 3860 36179 3906
rect 36225 3860 36295 3906
rect 36341 3860 36411 3906
rect 36457 3860 36527 3906
rect 36573 3860 36643 3906
rect 36689 3860 36759 3906
rect 36805 3860 36875 3906
rect 36921 3860 36991 3906
rect 37037 3860 37107 3906
rect 37153 3860 37223 3906
rect 37269 3860 37339 3906
rect 37385 3860 37455 3906
rect 37501 3860 37571 3906
rect 37617 3860 37687 3906
rect 37733 3860 37803 3906
rect 37849 3860 37919 3906
rect 37965 3860 38035 3906
rect 38081 3860 38151 3906
rect 38197 3860 38267 3906
rect 38313 3860 38383 3906
rect 38429 3860 38499 3906
rect 38545 3860 38615 3906
rect 38661 3860 38731 3906
rect 38777 3860 38847 3906
rect 38893 3860 38963 3906
rect 39009 3860 39079 3906
rect 39125 3860 39195 3906
rect 39241 3860 39311 3906
rect 39357 3860 39427 3906
rect 39473 3860 39543 3906
rect 39589 3860 39659 3906
rect 39705 3860 39775 3906
rect 39821 3860 39891 3906
rect 39937 3860 40007 3906
rect 40053 3860 40123 3906
rect 40169 3860 40180 3906
rect 28628 3790 40180 3860
rect 28628 3744 28639 3790
rect 28685 3744 28755 3790
rect 28801 3744 28871 3790
rect 28917 3744 28987 3790
rect 29033 3744 29103 3790
rect 29149 3744 29219 3790
rect 29265 3744 29335 3790
rect 29381 3744 29451 3790
rect 29497 3744 29567 3790
rect 29613 3744 29683 3790
rect 29729 3744 29799 3790
rect 29845 3744 29915 3790
rect 29961 3744 30031 3790
rect 30077 3744 30147 3790
rect 30193 3744 30263 3790
rect 30309 3744 30379 3790
rect 30425 3744 30495 3790
rect 30541 3744 30611 3790
rect 30657 3744 30727 3790
rect 30773 3744 30843 3790
rect 30889 3744 30959 3790
rect 31005 3744 31075 3790
rect 31121 3744 31191 3790
rect 31237 3744 31307 3790
rect 31353 3744 31423 3790
rect 31469 3744 31539 3790
rect 31585 3744 31655 3790
rect 31701 3744 31771 3790
rect 31817 3744 31887 3790
rect 31933 3744 32003 3790
rect 32049 3744 32119 3790
rect 32165 3744 32235 3790
rect 32281 3744 32351 3790
rect 32397 3744 32467 3790
rect 32513 3744 32583 3790
rect 32629 3744 32699 3790
rect 32745 3744 32815 3790
rect 32861 3744 32931 3790
rect 32977 3744 33047 3790
rect 33093 3744 33163 3790
rect 33209 3744 33279 3790
rect 33325 3744 33395 3790
rect 33441 3744 33511 3790
rect 33557 3744 33627 3790
rect 33673 3744 33743 3790
rect 33789 3744 33859 3790
rect 33905 3744 33975 3790
rect 34021 3744 34091 3790
rect 34137 3744 34207 3790
rect 34253 3744 34323 3790
rect 34369 3744 34439 3790
rect 34485 3744 34555 3790
rect 34601 3744 34671 3790
rect 34717 3744 34787 3790
rect 34833 3744 34903 3790
rect 34949 3744 35019 3790
rect 35065 3744 35135 3790
rect 35181 3744 35251 3790
rect 35297 3744 35367 3790
rect 35413 3744 35483 3790
rect 35529 3744 35599 3790
rect 35645 3744 35715 3790
rect 35761 3744 35831 3790
rect 35877 3744 35947 3790
rect 35993 3744 36063 3790
rect 36109 3744 36179 3790
rect 36225 3744 36295 3790
rect 36341 3744 36411 3790
rect 36457 3744 36527 3790
rect 36573 3744 36643 3790
rect 36689 3744 36759 3790
rect 36805 3744 36875 3790
rect 36921 3744 36991 3790
rect 37037 3744 37107 3790
rect 37153 3744 37223 3790
rect 37269 3744 37339 3790
rect 37385 3744 37455 3790
rect 37501 3744 37571 3790
rect 37617 3744 37687 3790
rect 37733 3744 37803 3790
rect 37849 3744 37919 3790
rect 37965 3744 38035 3790
rect 38081 3744 38151 3790
rect 38197 3744 38267 3790
rect 38313 3744 38383 3790
rect 38429 3744 38499 3790
rect 38545 3744 38615 3790
rect 38661 3744 38731 3790
rect 38777 3744 38847 3790
rect 38893 3744 38963 3790
rect 39009 3744 39079 3790
rect 39125 3744 39195 3790
rect 39241 3744 39311 3790
rect 39357 3744 39427 3790
rect 39473 3744 39543 3790
rect 39589 3744 39659 3790
rect 39705 3744 39775 3790
rect 39821 3744 39891 3790
rect 39937 3744 40007 3790
rect 40053 3744 40123 3790
rect 40169 3744 40180 3790
rect 28628 3674 40180 3744
rect 28628 3628 28639 3674
rect 28685 3628 28755 3674
rect 28801 3628 28871 3674
rect 28917 3628 28987 3674
rect 29033 3628 29103 3674
rect 29149 3628 29219 3674
rect 29265 3628 29335 3674
rect 29381 3628 29451 3674
rect 29497 3628 29567 3674
rect 29613 3628 29683 3674
rect 29729 3628 29799 3674
rect 29845 3628 29915 3674
rect 29961 3628 30031 3674
rect 30077 3628 30147 3674
rect 30193 3628 30263 3674
rect 30309 3628 30379 3674
rect 30425 3628 30495 3674
rect 30541 3628 30611 3674
rect 30657 3628 30727 3674
rect 30773 3628 30843 3674
rect 30889 3628 30959 3674
rect 31005 3628 31075 3674
rect 31121 3628 31191 3674
rect 31237 3628 31307 3674
rect 31353 3628 31423 3674
rect 31469 3628 31539 3674
rect 31585 3628 31655 3674
rect 31701 3628 31771 3674
rect 31817 3628 31887 3674
rect 31933 3628 32003 3674
rect 32049 3628 32119 3674
rect 32165 3628 32235 3674
rect 32281 3628 32351 3674
rect 32397 3628 32467 3674
rect 32513 3628 32583 3674
rect 32629 3628 32699 3674
rect 32745 3628 32815 3674
rect 32861 3628 32931 3674
rect 32977 3628 33047 3674
rect 33093 3628 33163 3674
rect 33209 3628 33279 3674
rect 33325 3628 33395 3674
rect 33441 3628 33511 3674
rect 33557 3628 33627 3674
rect 33673 3628 33743 3674
rect 33789 3628 33859 3674
rect 33905 3628 33975 3674
rect 34021 3628 34091 3674
rect 34137 3628 34207 3674
rect 34253 3628 34323 3674
rect 34369 3628 34439 3674
rect 34485 3628 34555 3674
rect 34601 3628 34671 3674
rect 34717 3628 34787 3674
rect 34833 3628 34903 3674
rect 34949 3628 35019 3674
rect 35065 3628 35135 3674
rect 35181 3628 35251 3674
rect 35297 3628 35367 3674
rect 35413 3628 35483 3674
rect 35529 3628 35599 3674
rect 35645 3628 35715 3674
rect 35761 3628 35831 3674
rect 35877 3628 35947 3674
rect 35993 3628 36063 3674
rect 36109 3628 36179 3674
rect 36225 3628 36295 3674
rect 36341 3628 36411 3674
rect 36457 3628 36527 3674
rect 36573 3628 36643 3674
rect 36689 3628 36759 3674
rect 36805 3628 36875 3674
rect 36921 3628 36991 3674
rect 37037 3628 37107 3674
rect 37153 3628 37223 3674
rect 37269 3628 37339 3674
rect 37385 3628 37455 3674
rect 37501 3628 37571 3674
rect 37617 3628 37687 3674
rect 37733 3628 37803 3674
rect 37849 3628 37919 3674
rect 37965 3628 38035 3674
rect 38081 3628 38151 3674
rect 38197 3628 38267 3674
rect 38313 3628 38383 3674
rect 38429 3628 38499 3674
rect 38545 3628 38615 3674
rect 38661 3628 38731 3674
rect 38777 3628 38847 3674
rect 38893 3628 38963 3674
rect 39009 3628 39079 3674
rect 39125 3628 39195 3674
rect 39241 3628 39311 3674
rect 39357 3628 39427 3674
rect 39473 3628 39543 3674
rect 39589 3628 39659 3674
rect 39705 3628 39775 3674
rect 39821 3628 39891 3674
rect 39937 3628 40007 3674
rect 40053 3628 40123 3674
rect 40169 3628 40180 3674
rect 28628 3558 40180 3628
rect 28628 3512 28639 3558
rect 28685 3512 28755 3558
rect 28801 3512 28871 3558
rect 28917 3512 28987 3558
rect 29033 3512 29103 3558
rect 29149 3512 29219 3558
rect 29265 3512 29335 3558
rect 29381 3512 29451 3558
rect 29497 3512 29567 3558
rect 29613 3512 29683 3558
rect 29729 3512 29799 3558
rect 29845 3512 29915 3558
rect 29961 3512 30031 3558
rect 30077 3512 30147 3558
rect 30193 3512 30263 3558
rect 30309 3512 30379 3558
rect 30425 3512 30495 3558
rect 30541 3512 30611 3558
rect 30657 3512 30727 3558
rect 30773 3512 30843 3558
rect 30889 3512 30959 3558
rect 31005 3512 31075 3558
rect 31121 3512 31191 3558
rect 31237 3512 31307 3558
rect 31353 3512 31423 3558
rect 31469 3512 31539 3558
rect 31585 3512 31655 3558
rect 31701 3512 31771 3558
rect 31817 3512 31887 3558
rect 31933 3512 32003 3558
rect 32049 3512 32119 3558
rect 32165 3512 32235 3558
rect 32281 3512 32351 3558
rect 32397 3512 32467 3558
rect 32513 3512 32583 3558
rect 32629 3512 32699 3558
rect 32745 3512 32815 3558
rect 32861 3512 32931 3558
rect 32977 3512 33047 3558
rect 33093 3512 33163 3558
rect 33209 3512 33279 3558
rect 33325 3512 33395 3558
rect 33441 3512 33511 3558
rect 33557 3512 33627 3558
rect 33673 3512 33743 3558
rect 33789 3512 33859 3558
rect 33905 3512 33975 3558
rect 34021 3512 34091 3558
rect 34137 3512 34207 3558
rect 34253 3512 34323 3558
rect 34369 3512 34439 3558
rect 34485 3512 34555 3558
rect 34601 3512 34671 3558
rect 34717 3512 34787 3558
rect 34833 3512 34903 3558
rect 34949 3512 35019 3558
rect 35065 3512 35135 3558
rect 35181 3512 35251 3558
rect 35297 3512 35367 3558
rect 35413 3512 35483 3558
rect 35529 3512 35599 3558
rect 35645 3512 35715 3558
rect 35761 3512 35831 3558
rect 35877 3512 35947 3558
rect 35993 3512 36063 3558
rect 36109 3512 36179 3558
rect 36225 3512 36295 3558
rect 36341 3512 36411 3558
rect 36457 3512 36527 3558
rect 36573 3512 36643 3558
rect 36689 3512 36759 3558
rect 36805 3512 36875 3558
rect 36921 3512 36991 3558
rect 37037 3512 37107 3558
rect 37153 3512 37223 3558
rect 37269 3512 37339 3558
rect 37385 3512 37455 3558
rect 37501 3512 37571 3558
rect 37617 3512 37687 3558
rect 37733 3512 37803 3558
rect 37849 3512 37919 3558
rect 37965 3512 38035 3558
rect 38081 3512 38151 3558
rect 38197 3512 38267 3558
rect 38313 3512 38383 3558
rect 38429 3512 38499 3558
rect 38545 3512 38615 3558
rect 38661 3512 38731 3558
rect 38777 3512 38847 3558
rect 38893 3512 38963 3558
rect 39009 3512 39079 3558
rect 39125 3512 39195 3558
rect 39241 3512 39311 3558
rect 39357 3512 39427 3558
rect 39473 3512 39543 3558
rect 39589 3512 39659 3558
rect 39705 3512 39775 3558
rect 39821 3512 39891 3558
rect 39937 3512 40007 3558
rect 40053 3512 40123 3558
rect 40169 3512 40180 3558
rect 28628 3442 40180 3512
rect 28628 3396 28639 3442
rect 28685 3396 28755 3442
rect 28801 3396 28871 3442
rect 28917 3396 28987 3442
rect 29033 3396 29103 3442
rect 29149 3396 29219 3442
rect 29265 3396 29335 3442
rect 29381 3396 29451 3442
rect 29497 3396 29567 3442
rect 29613 3396 29683 3442
rect 29729 3396 29799 3442
rect 29845 3396 29915 3442
rect 29961 3396 30031 3442
rect 30077 3396 30147 3442
rect 30193 3396 30263 3442
rect 30309 3396 30379 3442
rect 30425 3396 30495 3442
rect 30541 3396 30611 3442
rect 30657 3396 30727 3442
rect 30773 3396 30843 3442
rect 30889 3396 30959 3442
rect 31005 3396 31075 3442
rect 31121 3396 31191 3442
rect 31237 3396 31307 3442
rect 31353 3396 31423 3442
rect 31469 3396 31539 3442
rect 31585 3396 31655 3442
rect 31701 3396 31771 3442
rect 31817 3396 31887 3442
rect 31933 3396 32003 3442
rect 32049 3396 32119 3442
rect 32165 3396 32235 3442
rect 32281 3396 32351 3442
rect 32397 3396 32467 3442
rect 32513 3396 32583 3442
rect 32629 3396 32699 3442
rect 32745 3396 32815 3442
rect 32861 3396 32931 3442
rect 32977 3396 33047 3442
rect 33093 3396 33163 3442
rect 33209 3396 33279 3442
rect 33325 3396 33395 3442
rect 33441 3396 33511 3442
rect 33557 3396 33627 3442
rect 33673 3396 33743 3442
rect 33789 3396 33859 3442
rect 33905 3396 33975 3442
rect 34021 3396 34091 3442
rect 34137 3396 34207 3442
rect 34253 3396 34323 3442
rect 34369 3396 34439 3442
rect 34485 3396 34555 3442
rect 34601 3396 34671 3442
rect 34717 3396 34787 3442
rect 34833 3396 34903 3442
rect 34949 3396 35019 3442
rect 35065 3396 35135 3442
rect 35181 3396 35251 3442
rect 35297 3396 35367 3442
rect 35413 3396 35483 3442
rect 35529 3396 35599 3442
rect 35645 3396 35715 3442
rect 35761 3396 35831 3442
rect 35877 3396 35947 3442
rect 35993 3396 36063 3442
rect 36109 3396 36179 3442
rect 36225 3396 36295 3442
rect 36341 3396 36411 3442
rect 36457 3396 36527 3442
rect 36573 3396 36643 3442
rect 36689 3396 36759 3442
rect 36805 3396 36875 3442
rect 36921 3396 36991 3442
rect 37037 3396 37107 3442
rect 37153 3396 37223 3442
rect 37269 3396 37339 3442
rect 37385 3396 37455 3442
rect 37501 3396 37571 3442
rect 37617 3396 37687 3442
rect 37733 3396 37803 3442
rect 37849 3396 37919 3442
rect 37965 3396 38035 3442
rect 38081 3396 38151 3442
rect 38197 3396 38267 3442
rect 38313 3396 38383 3442
rect 38429 3396 38499 3442
rect 38545 3396 38615 3442
rect 38661 3396 38731 3442
rect 38777 3396 38847 3442
rect 38893 3396 38963 3442
rect 39009 3396 39079 3442
rect 39125 3396 39195 3442
rect 39241 3396 39311 3442
rect 39357 3396 39427 3442
rect 39473 3396 39543 3442
rect 39589 3396 39659 3442
rect 39705 3396 39775 3442
rect 39821 3396 39891 3442
rect 39937 3396 40007 3442
rect 40053 3396 40123 3442
rect 40169 3396 40180 3442
rect 28628 3326 40180 3396
rect 28628 3280 28639 3326
rect 28685 3280 28755 3326
rect 28801 3280 28871 3326
rect 28917 3280 28987 3326
rect 29033 3280 29103 3326
rect 29149 3280 29219 3326
rect 29265 3280 29335 3326
rect 29381 3280 29451 3326
rect 29497 3280 29567 3326
rect 29613 3280 29683 3326
rect 29729 3280 29799 3326
rect 29845 3280 29915 3326
rect 29961 3280 30031 3326
rect 30077 3280 30147 3326
rect 30193 3280 30263 3326
rect 30309 3280 30379 3326
rect 30425 3280 30495 3326
rect 30541 3280 30611 3326
rect 30657 3280 30727 3326
rect 30773 3280 30843 3326
rect 30889 3280 30959 3326
rect 31005 3280 31075 3326
rect 31121 3280 31191 3326
rect 31237 3280 31307 3326
rect 31353 3280 31423 3326
rect 31469 3280 31539 3326
rect 31585 3280 31655 3326
rect 31701 3280 31771 3326
rect 31817 3280 31887 3326
rect 31933 3280 32003 3326
rect 32049 3280 32119 3326
rect 32165 3280 32235 3326
rect 32281 3280 32351 3326
rect 32397 3280 32467 3326
rect 32513 3280 32583 3326
rect 32629 3280 32699 3326
rect 32745 3280 32815 3326
rect 32861 3280 32931 3326
rect 32977 3280 33047 3326
rect 33093 3280 33163 3326
rect 33209 3280 33279 3326
rect 33325 3280 33395 3326
rect 33441 3280 33511 3326
rect 33557 3280 33627 3326
rect 33673 3280 33743 3326
rect 33789 3280 33859 3326
rect 33905 3280 33975 3326
rect 34021 3280 34091 3326
rect 34137 3280 34207 3326
rect 34253 3280 34323 3326
rect 34369 3280 34439 3326
rect 34485 3280 34555 3326
rect 34601 3280 34671 3326
rect 34717 3280 34787 3326
rect 34833 3280 34903 3326
rect 34949 3280 35019 3326
rect 35065 3280 35135 3326
rect 35181 3280 35251 3326
rect 35297 3280 35367 3326
rect 35413 3280 35483 3326
rect 35529 3280 35599 3326
rect 35645 3280 35715 3326
rect 35761 3280 35831 3326
rect 35877 3280 35947 3326
rect 35993 3280 36063 3326
rect 36109 3280 36179 3326
rect 36225 3280 36295 3326
rect 36341 3280 36411 3326
rect 36457 3280 36527 3326
rect 36573 3280 36643 3326
rect 36689 3280 36759 3326
rect 36805 3280 36875 3326
rect 36921 3280 36991 3326
rect 37037 3280 37107 3326
rect 37153 3280 37223 3326
rect 37269 3280 37339 3326
rect 37385 3280 37455 3326
rect 37501 3280 37571 3326
rect 37617 3280 37687 3326
rect 37733 3280 37803 3326
rect 37849 3280 37919 3326
rect 37965 3280 38035 3326
rect 38081 3280 38151 3326
rect 38197 3280 38267 3326
rect 38313 3280 38383 3326
rect 38429 3280 38499 3326
rect 38545 3280 38615 3326
rect 38661 3280 38731 3326
rect 38777 3280 38847 3326
rect 38893 3280 38963 3326
rect 39009 3280 39079 3326
rect 39125 3280 39195 3326
rect 39241 3280 39311 3326
rect 39357 3280 39427 3326
rect 39473 3280 39543 3326
rect 39589 3280 39659 3326
rect 39705 3280 39775 3326
rect 39821 3280 39891 3326
rect 39937 3280 40007 3326
rect 40053 3280 40123 3326
rect 40169 3280 40180 3326
rect 28628 3210 40180 3280
rect 28628 3164 28639 3210
rect 28685 3164 28755 3210
rect 28801 3164 28871 3210
rect 28917 3164 28987 3210
rect 29033 3164 29103 3210
rect 29149 3164 29219 3210
rect 29265 3164 29335 3210
rect 29381 3164 29451 3210
rect 29497 3164 29567 3210
rect 29613 3164 29683 3210
rect 29729 3164 29799 3210
rect 29845 3164 29915 3210
rect 29961 3164 30031 3210
rect 30077 3164 30147 3210
rect 30193 3164 30263 3210
rect 30309 3164 30379 3210
rect 30425 3164 30495 3210
rect 30541 3164 30611 3210
rect 30657 3164 30727 3210
rect 30773 3164 30843 3210
rect 30889 3164 30959 3210
rect 31005 3164 31075 3210
rect 31121 3164 31191 3210
rect 31237 3164 31307 3210
rect 31353 3164 31423 3210
rect 31469 3164 31539 3210
rect 31585 3164 31655 3210
rect 31701 3164 31771 3210
rect 31817 3164 31887 3210
rect 31933 3164 32003 3210
rect 32049 3164 32119 3210
rect 32165 3164 32235 3210
rect 32281 3164 32351 3210
rect 32397 3164 32467 3210
rect 32513 3164 32583 3210
rect 32629 3164 32699 3210
rect 32745 3164 32815 3210
rect 32861 3164 32931 3210
rect 32977 3164 33047 3210
rect 33093 3164 33163 3210
rect 33209 3164 33279 3210
rect 33325 3164 33395 3210
rect 33441 3164 33511 3210
rect 33557 3164 33627 3210
rect 33673 3164 33743 3210
rect 33789 3164 33859 3210
rect 33905 3164 33975 3210
rect 34021 3164 34091 3210
rect 34137 3164 34207 3210
rect 34253 3164 34323 3210
rect 34369 3164 34439 3210
rect 34485 3164 34555 3210
rect 34601 3164 34671 3210
rect 34717 3164 34787 3210
rect 34833 3164 34903 3210
rect 34949 3164 35019 3210
rect 35065 3164 35135 3210
rect 35181 3164 35251 3210
rect 35297 3164 35367 3210
rect 35413 3164 35483 3210
rect 35529 3164 35599 3210
rect 35645 3164 35715 3210
rect 35761 3164 35831 3210
rect 35877 3164 35947 3210
rect 35993 3164 36063 3210
rect 36109 3164 36179 3210
rect 36225 3164 36295 3210
rect 36341 3164 36411 3210
rect 36457 3164 36527 3210
rect 36573 3164 36643 3210
rect 36689 3164 36759 3210
rect 36805 3164 36875 3210
rect 36921 3164 36991 3210
rect 37037 3164 37107 3210
rect 37153 3164 37223 3210
rect 37269 3164 37339 3210
rect 37385 3164 37455 3210
rect 37501 3164 37571 3210
rect 37617 3164 37687 3210
rect 37733 3164 37803 3210
rect 37849 3164 37919 3210
rect 37965 3164 38035 3210
rect 38081 3164 38151 3210
rect 38197 3164 38267 3210
rect 38313 3164 38383 3210
rect 38429 3164 38499 3210
rect 38545 3164 38615 3210
rect 38661 3164 38731 3210
rect 38777 3164 38847 3210
rect 38893 3164 38963 3210
rect 39009 3164 39079 3210
rect 39125 3164 39195 3210
rect 39241 3164 39311 3210
rect 39357 3164 39427 3210
rect 39473 3164 39543 3210
rect 39589 3164 39659 3210
rect 39705 3164 39775 3210
rect 39821 3164 39891 3210
rect 39937 3164 40007 3210
rect 40053 3164 40123 3210
rect 40169 3164 40180 3210
rect 28628 3094 40180 3164
rect 28628 3048 28639 3094
rect 28685 3048 28755 3094
rect 28801 3048 28871 3094
rect 28917 3048 28987 3094
rect 29033 3048 29103 3094
rect 29149 3048 29219 3094
rect 29265 3048 29335 3094
rect 29381 3048 29451 3094
rect 29497 3048 29567 3094
rect 29613 3048 29683 3094
rect 29729 3048 29799 3094
rect 29845 3048 29915 3094
rect 29961 3048 30031 3094
rect 30077 3048 30147 3094
rect 30193 3048 30263 3094
rect 30309 3048 30379 3094
rect 30425 3048 30495 3094
rect 30541 3048 30611 3094
rect 30657 3048 30727 3094
rect 30773 3048 30843 3094
rect 30889 3048 30959 3094
rect 31005 3048 31075 3094
rect 31121 3048 31191 3094
rect 31237 3048 31307 3094
rect 31353 3048 31423 3094
rect 31469 3048 31539 3094
rect 31585 3048 31655 3094
rect 31701 3048 31771 3094
rect 31817 3048 31887 3094
rect 31933 3048 32003 3094
rect 32049 3048 32119 3094
rect 32165 3048 32235 3094
rect 32281 3048 32351 3094
rect 32397 3048 32467 3094
rect 32513 3048 32583 3094
rect 32629 3048 32699 3094
rect 32745 3048 32815 3094
rect 32861 3048 32931 3094
rect 32977 3048 33047 3094
rect 33093 3048 33163 3094
rect 33209 3048 33279 3094
rect 33325 3048 33395 3094
rect 33441 3048 33511 3094
rect 33557 3048 33627 3094
rect 33673 3048 33743 3094
rect 33789 3048 33859 3094
rect 33905 3048 33975 3094
rect 34021 3048 34091 3094
rect 34137 3048 34207 3094
rect 34253 3048 34323 3094
rect 34369 3048 34439 3094
rect 34485 3048 34555 3094
rect 34601 3048 34671 3094
rect 34717 3048 34787 3094
rect 34833 3048 34903 3094
rect 34949 3048 35019 3094
rect 35065 3048 35135 3094
rect 35181 3048 35251 3094
rect 35297 3048 35367 3094
rect 35413 3048 35483 3094
rect 35529 3048 35599 3094
rect 35645 3048 35715 3094
rect 35761 3048 35831 3094
rect 35877 3048 35947 3094
rect 35993 3048 36063 3094
rect 36109 3048 36179 3094
rect 36225 3048 36295 3094
rect 36341 3048 36411 3094
rect 36457 3048 36527 3094
rect 36573 3048 36643 3094
rect 36689 3048 36759 3094
rect 36805 3048 36875 3094
rect 36921 3048 36991 3094
rect 37037 3048 37107 3094
rect 37153 3048 37223 3094
rect 37269 3048 37339 3094
rect 37385 3048 37455 3094
rect 37501 3048 37571 3094
rect 37617 3048 37687 3094
rect 37733 3048 37803 3094
rect 37849 3048 37919 3094
rect 37965 3048 38035 3094
rect 38081 3048 38151 3094
rect 38197 3048 38267 3094
rect 38313 3048 38383 3094
rect 38429 3048 38499 3094
rect 38545 3048 38615 3094
rect 38661 3048 38731 3094
rect 38777 3048 38847 3094
rect 38893 3048 38963 3094
rect 39009 3048 39079 3094
rect 39125 3048 39195 3094
rect 39241 3048 39311 3094
rect 39357 3048 39427 3094
rect 39473 3048 39543 3094
rect 39589 3048 39659 3094
rect 39705 3048 39775 3094
rect 39821 3048 39891 3094
rect 39937 3048 40007 3094
rect 40053 3048 40123 3094
rect 40169 3048 40180 3094
rect 28628 2978 40180 3048
rect 28628 2932 28639 2978
rect 28685 2932 28755 2978
rect 28801 2932 28871 2978
rect 28917 2932 28987 2978
rect 29033 2932 29103 2978
rect 29149 2932 29219 2978
rect 29265 2932 29335 2978
rect 29381 2932 29451 2978
rect 29497 2932 29567 2978
rect 29613 2932 29683 2978
rect 29729 2932 29799 2978
rect 29845 2932 29915 2978
rect 29961 2932 30031 2978
rect 30077 2932 30147 2978
rect 30193 2932 30263 2978
rect 30309 2932 30379 2978
rect 30425 2932 30495 2978
rect 30541 2932 30611 2978
rect 30657 2932 30727 2978
rect 30773 2932 30843 2978
rect 30889 2932 30959 2978
rect 31005 2932 31075 2978
rect 31121 2932 31191 2978
rect 31237 2932 31307 2978
rect 31353 2932 31423 2978
rect 31469 2932 31539 2978
rect 31585 2932 31655 2978
rect 31701 2932 31771 2978
rect 31817 2932 31887 2978
rect 31933 2932 32003 2978
rect 32049 2932 32119 2978
rect 32165 2932 32235 2978
rect 32281 2932 32351 2978
rect 32397 2932 32467 2978
rect 32513 2932 32583 2978
rect 32629 2932 32699 2978
rect 32745 2932 32815 2978
rect 32861 2932 32931 2978
rect 32977 2932 33047 2978
rect 33093 2932 33163 2978
rect 33209 2932 33279 2978
rect 33325 2932 33395 2978
rect 33441 2932 33511 2978
rect 33557 2932 33627 2978
rect 33673 2932 33743 2978
rect 33789 2932 33859 2978
rect 33905 2932 33975 2978
rect 34021 2932 34091 2978
rect 34137 2932 34207 2978
rect 34253 2932 34323 2978
rect 34369 2932 34439 2978
rect 34485 2932 34555 2978
rect 34601 2932 34671 2978
rect 34717 2932 34787 2978
rect 34833 2932 34903 2978
rect 34949 2932 35019 2978
rect 35065 2932 35135 2978
rect 35181 2932 35251 2978
rect 35297 2932 35367 2978
rect 35413 2932 35483 2978
rect 35529 2932 35599 2978
rect 35645 2932 35715 2978
rect 35761 2932 35831 2978
rect 35877 2932 35947 2978
rect 35993 2932 36063 2978
rect 36109 2932 36179 2978
rect 36225 2932 36295 2978
rect 36341 2932 36411 2978
rect 36457 2932 36527 2978
rect 36573 2932 36643 2978
rect 36689 2932 36759 2978
rect 36805 2932 36875 2978
rect 36921 2932 36991 2978
rect 37037 2932 37107 2978
rect 37153 2932 37223 2978
rect 37269 2932 37339 2978
rect 37385 2932 37455 2978
rect 37501 2932 37571 2978
rect 37617 2932 37687 2978
rect 37733 2932 37803 2978
rect 37849 2932 37919 2978
rect 37965 2932 38035 2978
rect 38081 2932 38151 2978
rect 38197 2932 38267 2978
rect 38313 2932 38383 2978
rect 38429 2932 38499 2978
rect 38545 2932 38615 2978
rect 38661 2932 38731 2978
rect 38777 2932 38847 2978
rect 38893 2932 38963 2978
rect 39009 2932 39079 2978
rect 39125 2932 39195 2978
rect 39241 2932 39311 2978
rect 39357 2932 39427 2978
rect 39473 2932 39543 2978
rect 39589 2932 39659 2978
rect 39705 2932 39775 2978
rect 39821 2932 39891 2978
rect 39937 2932 40007 2978
rect 40053 2932 40123 2978
rect 40169 2932 40180 2978
rect 28628 2862 40180 2932
rect 28628 2816 28639 2862
rect 28685 2816 28755 2862
rect 28801 2816 28871 2862
rect 28917 2816 28987 2862
rect 29033 2816 29103 2862
rect 29149 2816 29219 2862
rect 29265 2816 29335 2862
rect 29381 2816 29451 2862
rect 29497 2816 29567 2862
rect 29613 2816 29683 2862
rect 29729 2816 29799 2862
rect 29845 2816 29915 2862
rect 29961 2816 30031 2862
rect 30077 2816 30147 2862
rect 30193 2816 30263 2862
rect 30309 2816 30379 2862
rect 30425 2816 30495 2862
rect 30541 2816 30611 2862
rect 30657 2816 30727 2862
rect 30773 2816 30843 2862
rect 30889 2816 30959 2862
rect 31005 2816 31075 2862
rect 31121 2816 31191 2862
rect 31237 2816 31307 2862
rect 31353 2816 31423 2862
rect 31469 2816 31539 2862
rect 31585 2816 31655 2862
rect 31701 2816 31771 2862
rect 31817 2816 31887 2862
rect 31933 2816 32003 2862
rect 32049 2816 32119 2862
rect 32165 2816 32235 2862
rect 32281 2816 32351 2862
rect 32397 2816 32467 2862
rect 32513 2816 32583 2862
rect 32629 2816 32699 2862
rect 32745 2816 32815 2862
rect 32861 2816 32931 2862
rect 32977 2816 33047 2862
rect 33093 2816 33163 2862
rect 33209 2816 33279 2862
rect 33325 2816 33395 2862
rect 33441 2816 33511 2862
rect 33557 2816 33627 2862
rect 33673 2816 33743 2862
rect 33789 2816 33859 2862
rect 33905 2816 33975 2862
rect 34021 2816 34091 2862
rect 34137 2816 34207 2862
rect 34253 2816 34323 2862
rect 34369 2816 34439 2862
rect 34485 2816 34555 2862
rect 34601 2816 34671 2862
rect 34717 2816 34787 2862
rect 34833 2816 34903 2862
rect 34949 2816 35019 2862
rect 35065 2816 35135 2862
rect 35181 2816 35251 2862
rect 35297 2816 35367 2862
rect 35413 2816 35483 2862
rect 35529 2816 35599 2862
rect 35645 2816 35715 2862
rect 35761 2816 35831 2862
rect 35877 2816 35947 2862
rect 35993 2816 36063 2862
rect 36109 2816 36179 2862
rect 36225 2816 36295 2862
rect 36341 2816 36411 2862
rect 36457 2816 36527 2862
rect 36573 2816 36643 2862
rect 36689 2816 36759 2862
rect 36805 2816 36875 2862
rect 36921 2816 36991 2862
rect 37037 2816 37107 2862
rect 37153 2816 37223 2862
rect 37269 2816 37339 2862
rect 37385 2816 37455 2862
rect 37501 2816 37571 2862
rect 37617 2816 37687 2862
rect 37733 2816 37803 2862
rect 37849 2816 37919 2862
rect 37965 2816 38035 2862
rect 38081 2816 38151 2862
rect 38197 2816 38267 2862
rect 38313 2816 38383 2862
rect 38429 2816 38499 2862
rect 38545 2816 38615 2862
rect 38661 2816 38731 2862
rect 38777 2816 38847 2862
rect 38893 2816 38963 2862
rect 39009 2816 39079 2862
rect 39125 2816 39195 2862
rect 39241 2816 39311 2862
rect 39357 2816 39427 2862
rect 39473 2816 39543 2862
rect 39589 2816 39659 2862
rect 39705 2816 39775 2862
rect 39821 2816 39891 2862
rect 39937 2816 40007 2862
rect 40053 2816 40123 2862
rect 40169 2816 40180 2862
rect 28628 2746 40180 2816
rect 28628 2700 28639 2746
rect 28685 2700 28755 2746
rect 28801 2700 28871 2746
rect 28917 2700 28987 2746
rect 29033 2700 29103 2746
rect 29149 2700 29219 2746
rect 29265 2700 29335 2746
rect 29381 2700 29451 2746
rect 29497 2700 29567 2746
rect 29613 2700 29683 2746
rect 29729 2700 29799 2746
rect 29845 2700 29915 2746
rect 29961 2700 30031 2746
rect 30077 2700 30147 2746
rect 30193 2700 30263 2746
rect 30309 2700 30379 2746
rect 30425 2700 30495 2746
rect 30541 2700 30611 2746
rect 30657 2700 30727 2746
rect 30773 2700 30843 2746
rect 30889 2700 30959 2746
rect 31005 2700 31075 2746
rect 31121 2700 31191 2746
rect 31237 2700 31307 2746
rect 31353 2700 31423 2746
rect 31469 2700 31539 2746
rect 31585 2700 31655 2746
rect 31701 2700 31771 2746
rect 31817 2700 31887 2746
rect 31933 2700 32003 2746
rect 32049 2700 32119 2746
rect 32165 2700 32235 2746
rect 32281 2700 32351 2746
rect 32397 2700 32467 2746
rect 32513 2700 32583 2746
rect 32629 2700 32699 2746
rect 32745 2700 32815 2746
rect 32861 2700 32931 2746
rect 32977 2700 33047 2746
rect 33093 2700 33163 2746
rect 33209 2700 33279 2746
rect 33325 2700 33395 2746
rect 33441 2700 33511 2746
rect 33557 2700 33627 2746
rect 33673 2700 33743 2746
rect 33789 2700 33859 2746
rect 33905 2700 33975 2746
rect 34021 2700 34091 2746
rect 34137 2700 34207 2746
rect 34253 2700 34323 2746
rect 34369 2700 34439 2746
rect 34485 2700 34555 2746
rect 34601 2700 34671 2746
rect 34717 2700 34787 2746
rect 34833 2700 34903 2746
rect 34949 2700 35019 2746
rect 35065 2700 35135 2746
rect 35181 2700 35251 2746
rect 35297 2700 35367 2746
rect 35413 2700 35483 2746
rect 35529 2700 35599 2746
rect 35645 2700 35715 2746
rect 35761 2700 35831 2746
rect 35877 2700 35947 2746
rect 35993 2700 36063 2746
rect 36109 2700 36179 2746
rect 36225 2700 36295 2746
rect 36341 2700 36411 2746
rect 36457 2700 36527 2746
rect 36573 2700 36643 2746
rect 36689 2700 36759 2746
rect 36805 2700 36875 2746
rect 36921 2700 36991 2746
rect 37037 2700 37107 2746
rect 37153 2700 37223 2746
rect 37269 2700 37339 2746
rect 37385 2700 37455 2746
rect 37501 2700 37571 2746
rect 37617 2700 37687 2746
rect 37733 2700 37803 2746
rect 37849 2700 37919 2746
rect 37965 2700 38035 2746
rect 38081 2700 38151 2746
rect 38197 2700 38267 2746
rect 38313 2700 38383 2746
rect 38429 2700 38499 2746
rect 38545 2700 38615 2746
rect 38661 2700 38731 2746
rect 38777 2700 38847 2746
rect 38893 2700 38963 2746
rect 39009 2700 39079 2746
rect 39125 2700 39195 2746
rect 39241 2700 39311 2746
rect 39357 2700 39427 2746
rect 39473 2700 39543 2746
rect 39589 2700 39659 2746
rect 39705 2700 39775 2746
rect 39821 2700 39891 2746
rect 39937 2700 40007 2746
rect 40053 2700 40123 2746
rect 40169 2700 40180 2746
rect 28628 2630 40180 2700
rect 28628 2584 28639 2630
rect 28685 2584 28755 2630
rect 28801 2584 28871 2630
rect 28917 2584 28987 2630
rect 29033 2584 29103 2630
rect 29149 2584 29219 2630
rect 29265 2584 29335 2630
rect 29381 2584 29451 2630
rect 29497 2584 29567 2630
rect 29613 2584 29683 2630
rect 29729 2584 29799 2630
rect 29845 2584 29915 2630
rect 29961 2584 30031 2630
rect 30077 2584 30147 2630
rect 30193 2584 30263 2630
rect 30309 2584 30379 2630
rect 30425 2584 30495 2630
rect 30541 2584 30611 2630
rect 30657 2584 30727 2630
rect 30773 2584 30843 2630
rect 30889 2584 30959 2630
rect 31005 2584 31075 2630
rect 31121 2584 31191 2630
rect 31237 2584 31307 2630
rect 31353 2584 31423 2630
rect 31469 2584 31539 2630
rect 31585 2584 31655 2630
rect 31701 2584 31771 2630
rect 31817 2584 31887 2630
rect 31933 2584 32003 2630
rect 32049 2584 32119 2630
rect 32165 2584 32235 2630
rect 32281 2584 32351 2630
rect 32397 2584 32467 2630
rect 32513 2584 32583 2630
rect 32629 2584 32699 2630
rect 32745 2584 32815 2630
rect 32861 2584 32931 2630
rect 32977 2584 33047 2630
rect 33093 2584 33163 2630
rect 33209 2584 33279 2630
rect 33325 2584 33395 2630
rect 33441 2584 33511 2630
rect 33557 2584 33627 2630
rect 33673 2584 33743 2630
rect 33789 2584 33859 2630
rect 33905 2584 33975 2630
rect 34021 2584 34091 2630
rect 34137 2584 34207 2630
rect 34253 2584 34323 2630
rect 34369 2584 34439 2630
rect 34485 2584 34555 2630
rect 34601 2584 34671 2630
rect 34717 2584 34787 2630
rect 34833 2584 34903 2630
rect 34949 2584 35019 2630
rect 35065 2584 35135 2630
rect 35181 2584 35251 2630
rect 35297 2584 35367 2630
rect 35413 2584 35483 2630
rect 35529 2584 35599 2630
rect 35645 2584 35715 2630
rect 35761 2584 35831 2630
rect 35877 2584 35947 2630
rect 35993 2584 36063 2630
rect 36109 2584 36179 2630
rect 36225 2584 36295 2630
rect 36341 2584 36411 2630
rect 36457 2584 36527 2630
rect 36573 2584 36643 2630
rect 36689 2584 36759 2630
rect 36805 2584 36875 2630
rect 36921 2584 36991 2630
rect 37037 2584 37107 2630
rect 37153 2584 37223 2630
rect 37269 2584 37339 2630
rect 37385 2584 37455 2630
rect 37501 2584 37571 2630
rect 37617 2584 37687 2630
rect 37733 2584 37803 2630
rect 37849 2584 37919 2630
rect 37965 2584 38035 2630
rect 38081 2584 38151 2630
rect 38197 2584 38267 2630
rect 38313 2584 38383 2630
rect 38429 2584 38499 2630
rect 38545 2584 38615 2630
rect 38661 2584 38731 2630
rect 38777 2584 38847 2630
rect 38893 2584 38963 2630
rect 39009 2584 39079 2630
rect 39125 2584 39195 2630
rect 39241 2584 39311 2630
rect 39357 2584 39427 2630
rect 39473 2584 39543 2630
rect 39589 2584 39659 2630
rect 39705 2584 39775 2630
rect 39821 2584 39891 2630
rect 39937 2584 40007 2630
rect 40053 2584 40123 2630
rect 40169 2584 40180 2630
rect 28628 2514 40180 2584
rect 28628 2468 28639 2514
rect 28685 2468 28755 2514
rect 28801 2468 28871 2514
rect 28917 2468 28987 2514
rect 29033 2468 29103 2514
rect 29149 2468 29219 2514
rect 29265 2468 29335 2514
rect 29381 2468 29451 2514
rect 29497 2468 29567 2514
rect 29613 2468 29683 2514
rect 29729 2468 29799 2514
rect 29845 2468 29915 2514
rect 29961 2468 30031 2514
rect 30077 2468 30147 2514
rect 30193 2468 30263 2514
rect 30309 2468 30379 2514
rect 30425 2468 30495 2514
rect 30541 2468 30611 2514
rect 30657 2468 30727 2514
rect 30773 2468 30843 2514
rect 30889 2468 30959 2514
rect 31005 2468 31075 2514
rect 31121 2468 31191 2514
rect 31237 2468 31307 2514
rect 31353 2468 31423 2514
rect 31469 2468 31539 2514
rect 31585 2468 31655 2514
rect 31701 2468 31771 2514
rect 31817 2468 31887 2514
rect 31933 2468 32003 2514
rect 32049 2468 32119 2514
rect 32165 2468 32235 2514
rect 32281 2468 32351 2514
rect 32397 2468 32467 2514
rect 32513 2468 32583 2514
rect 32629 2468 32699 2514
rect 32745 2468 32815 2514
rect 32861 2468 32931 2514
rect 32977 2468 33047 2514
rect 33093 2468 33163 2514
rect 33209 2468 33279 2514
rect 33325 2468 33395 2514
rect 33441 2468 33511 2514
rect 33557 2468 33627 2514
rect 33673 2468 33743 2514
rect 33789 2468 33859 2514
rect 33905 2468 33975 2514
rect 34021 2468 34091 2514
rect 34137 2468 34207 2514
rect 34253 2468 34323 2514
rect 34369 2468 34439 2514
rect 34485 2468 34555 2514
rect 34601 2468 34671 2514
rect 34717 2468 34787 2514
rect 34833 2468 34903 2514
rect 34949 2468 35019 2514
rect 35065 2468 35135 2514
rect 35181 2468 35251 2514
rect 35297 2468 35367 2514
rect 35413 2468 35483 2514
rect 35529 2468 35599 2514
rect 35645 2468 35715 2514
rect 35761 2468 35831 2514
rect 35877 2468 35947 2514
rect 35993 2468 36063 2514
rect 36109 2468 36179 2514
rect 36225 2468 36295 2514
rect 36341 2468 36411 2514
rect 36457 2468 36527 2514
rect 36573 2468 36643 2514
rect 36689 2468 36759 2514
rect 36805 2468 36875 2514
rect 36921 2468 36991 2514
rect 37037 2468 37107 2514
rect 37153 2468 37223 2514
rect 37269 2468 37339 2514
rect 37385 2468 37455 2514
rect 37501 2468 37571 2514
rect 37617 2468 37687 2514
rect 37733 2468 37803 2514
rect 37849 2468 37919 2514
rect 37965 2468 38035 2514
rect 38081 2468 38151 2514
rect 38197 2468 38267 2514
rect 38313 2468 38383 2514
rect 38429 2468 38499 2514
rect 38545 2468 38615 2514
rect 38661 2468 38731 2514
rect 38777 2468 38847 2514
rect 38893 2468 38963 2514
rect 39009 2468 39079 2514
rect 39125 2468 39195 2514
rect 39241 2468 39311 2514
rect 39357 2468 39427 2514
rect 39473 2468 39543 2514
rect 39589 2468 39659 2514
rect 39705 2468 39775 2514
rect 39821 2468 39891 2514
rect 39937 2468 40007 2514
rect 40053 2468 40123 2514
rect 40169 2468 40180 2514
rect 28628 2398 40180 2468
rect 28628 2352 28639 2398
rect 28685 2352 28755 2398
rect 28801 2352 28871 2398
rect 28917 2352 28987 2398
rect 29033 2352 29103 2398
rect 29149 2352 29219 2398
rect 29265 2352 29335 2398
rect 29381 2352 29451 2398
rect 29497 2352 29567 2398
rect 29613 2352 29683 2398
rect 29729 2352 29799 2398
rect 29845 2352 29915 2398
rect 29961 2352 30031 2398
rect 30077 2352 30147 2398
rect 30193 2352 30263 2398
rect 30309 2352 30379 2398
rect 30425 2352 30495 2398
rect 30541 2352 30611 2398
rect 30657 2352 30727 2398
rect 30773 2352 30843 2398
rect 30889 2352 30959 2398
rect 31005 2352 31075 2398
rect 31121 2352 31191 2398
rect 31237 2352 31307 2398
rect 31353 2352 31423 2398
rect 31469 2352 31539 2398
rect 31585 2352 31655 2398
rect 31701 2352 31771 2398
rect 31817 2352 31887 2398
rect 31933 2352 32003 2398
rect 32049 2352 32119 2398
rect 32165 2352 32235 2398
rect 32281 2352 32351 2398
rect 32397 2352 32467 2398
rect 32513 2352 32583 2398
rect 32629 2352 32699 2398
rect 32745 2352 32815 2398
rect 32861 2352 32931 2398
rect 32977 2352 33047 2398
rect 33093 2352 33163 2398
rect 33209 2352 33279 2398
rect 33325 2352 33395 2398
rect 33441 2352 33511 2398
rect 33557 2352 33627 2398
rect 33673 2352 33743 2398
rect 33789 2352 33859 2398
rect 33905 2352 33975 2398
rect 34021 2352 34091 2398
rect 34137 2352 34207 2398
rect 34253 2352 34323 2398
rect 34369 2352 34439 2398
rect 34485 2352 34555 2398
rect 34601 2352 34671 2398
rect 34717 2352 34787 2398
rect 34833 2352 34903 2398
rect 34949 2352 35019 2398
rect 35065 2352 35135 2398
rect 35181 2352 35251 2398
rect 35297 2352 35367 2398
rect 35413 2352 35483 2398
rect 35529 2352 35599 2398
rect 35645 2352 35715 2398
rect 35761 2352 35831 2398
rect 35877 2352 35947 2398
rect 35993 2352 36063 2398
rect 36109 2352 36179 2398
rect 36225 2352 36295 2398
rect 36341 2352 36411 2398
rect 36457 2352 36527 2398
rect 36573 2352 36643 2398
rect 36689 2352 36759 2398
rect 36805 2352 36875 2398
rect 36921 2352 36991 2398
rect 37037 2352 37107 2398
rect 37153 2352 37223 2398
rect 37269 2352 37339 2398
rect 37385 2352 37455 2398
rect 37501 2352 37571 2398
rect 37617 2352 37687 2398
rect 37733 2352 37803 2398
rect 37849 2352 37919 2398
rect 37965 2352 38035 2398
rect 38081 2352 38151 2398
rect 38197 2352 38267 2398
rect 38313 2352 38383 2398
rect 38429 2352 38499 2398
rect 38545 2352 38615 2398
rect 38661 2352 38731 2398
rect 38777 2352 38847 2398
rect 38893 2352 38963 2398
rect 39009 2352 39079 2398
rect 39125 2352 39195 2398
rect 39241 2352 39311 2398
rect 39357 2352 39427 2398
rect 39473 2352 39543 2398
rect 39589 2352 39659 2398
rect 39705 2352 39775 2398
rect 39821 2352 39891 2398
rect 39937 2352 40007 2398
rect 40053 2352 40123 2398
rect 40169 2352 40180 2398
rect 28628 2282 40180 2352
rect 28628 2236 28639 2282
rect 28685 2236 28755 2282
rect 28801 2236 28871 2282
rect 28917 2236 28987 2282
rect 29033 2236 29103 2282
rect 29149 2236 29219 2282
rect 29265 2236 29335 2282
rect 29381 2236 29451 2282
rect 29497 2236 29567 2282
rect 29613 2236 29683 2282
rect 29729 2236 29799 2282
rect 29845 2236 29915 2282
rect 29961 2236 30031 2282
rect 30077 2236 30147 2282
rect 30193 2236 30263 2282
rect 30309 2236 30379 2282
rect 30425 2236 30495 2282
rect 30541 2236 30611 2282
rect 30657 2236 30727 2282
rect 30773 2236 30843 2282
rect 30889 2236 30959 2282
rect 31005 2236 31075 2282
rect 31121 2236 31191 2282
rect 31237 2236 31307 2282
rect 31353 2236 31423 2282
rect 31469 2236 31539 2282
rect 31585 2236 31655 2282
rect 31701 2236 31771 2282
rect 31817 2236 31887 2282
rect 31933 2236 32003 2282
rect 32049 2236 32119 2282
rect 32165 2236 32235 2282
rect 32281 2236 32351 2282
rect 32397 2236 32467 2282
rect 32513 2236 32583 2282
rect 32629 2236 32699 2282
rect 32745 2236 32815 2282
rect 32861 2236 32931 2282
rect 32977 2236 33047 2282
rect 33093 2236 33163 2282
rect 33209 2236 33279 2282
rect 33325 2236 33395 2282
rect 33441 2236 33511 2282
rect 33557 2236 33627 2282
rect 33673 2236 33743 2282
rect 33789 2236 33859 2282
rect 33905 2236 33975 2282
rect 34021 2236 34091 2282
rect 34137 2236 34207 2282
rect 34253 2236 34323 2282
rect 34369 2236 34439 2282
rect 34485 2236 34555 2282
rect 34601 2236 34671 2282
rect 34717 2236 34787 2282
rect 34833 2236 34903 2282
rect 34949 2236 35019 2282
rect 35065 2236 35135 2282
rect 35181 2236 35251 2282
rect 35297 2236 35367 2282
rect 35413 2236 35483 2282
rect 35529 2236 35599 2282
rect 35645 2236 35715 2282
rect 35761 2236 35831 2282
rect 35877 2236 35947 2282
rect 35993 2236 36063 2282
rect 36109 2236 36179 2282
rect 36225 2236 36295 2282
rect 36341 2236 36411 2282
rect 36457 2236 36527 2282
rect 36573 2236 36643 2282
rect 36689 2236 36759 2282
rect 36805 2236 36875 2282
rect 36921 2236 36991 2282
rect 37037 2236 37107 2282
rect 37153 2236 37223 2282
rect 37269 2236 37339 2282
rect 37385 2236 37455 2282
rect 37501 2236 37571 2282
rect 37617 2236 37687 2282
rect 37733 2236 37803 2282
rect 37849 2236 37919 2282
rect 37965 2236 38035 2282
rect 38081 2236 38151 2282
rect 38197 2236 38267 2282
rect 38313 2236 38383 2282
rect 38429 2236 38499 2282
rect 38545 2236 38615 2282
rect 38661 2236 38731 2282
rect 38777 2236 38847 2282
rect 38893 2236 38963 2282
rect 39009 2236 39079 2282
rect 39125 2236 39195 2282
rect 39241 2236 39311 2282
rect 39357 2236 39427 2282
rect 39473 2236 39543 2282
rect 39589 2236 39659 2282
rect 39705 2236 39775 2282
rect 39821 2236 39891 2282
rect 39937 2236 40007 2282
rect 40053 2236 40123 2282
rect 40169 2236 40180 2282
rect 28628 2166 40180 2236
rect 28628 2120 28639 2166
rect 28685 2120 28755 2166
rect 28801 2120 28871 2166
rect 28917 2120 28987 2166
rect 29033 2120 29103 2166
rect 29149 2120 29219 2166
rect 29265 2120 29335 2166
rect 29381 2120 29451 2166
rect 29497 2120 29567 2166
rect 29613 2120 29683 2166
rect 29729 2120 29799 2166
rect 29845 2120 29915 2166
rect 29961 2120 30031 2166
rect 30077 2120 30147 2166
rect 30193 2120 30263 2166
rect 30309 2120 30379 2166
rect 30425 2120 30495 2166
rect 30541 2120 30611 2166
rect 30657 2120 30727 2166
rect 30773 2120 30843 2166
rect 30889 2120 30959 2166
rect 31005 2120 31075 2166
rect 31121 2120 31191 2166
rect 31237 2120 31307 2166
rect 31353 2120 31423 2166
rect 31469 2120 31539 2166
rect 31585 2120 31655 2166
rect 31701 2120 31771 2166
rect 31817 2120 31887 2166
rect 31933 2120 32003 2166
rect 32049 2120 32119 2166
rect 32165 2120 32235 2166
rect 32281 2120 32351 2166
rect 32397 2120 32467 2166
rect 32513 2120 32583 2166
rect 32629 2120 32699 2166
rect 32745 2120 32815 2166
rect 32861 2120 32931 2166
rect 32977 2120 33047 2166
rect 33093 2120 33163 2166
rect 33209 2120 33279 2166
rect 33325 2120 33395 2166
rect 33441 2120 33511 2166
rect 33557 2120 33627 2166
rect 33673 2120 33743 2166
rect 33789 2120 33859 2166
rect 33905 2120 33975 2166
rect 34021 2120 34091 2166
rect 34137 2120 34207 2166
rect 34253 2120 34323 2166
rect 34369 2120 34439 2166
rect 34485 2120 34555 2166
rect 34601 2120 34671 2166
rect 34717 2120 34787 2166
rect 34833 2120 34903 2166
rect 34949 2120 35019 2166
rect 35065 2120 35135 2166
rect 35181 2120 35251 2166
rect 35297 2120 35367 2166
rect 35413 2120 35483 2166
rect 35529 2120 35599 2166
rect 35645 2120 35715 2166
rect 35761 2120 35831 2166
rect 35877 2120 35947 2166
rect 35993 2120 36063 2166
rect 36109 2120 36179 2166
rect 36225 2120 36295 2166
rect 36341 2120 36411 2166
rect 36457 2120 36527 2166
rect 36573 2120 36643 2166
rect 36689 2120 36759 2166
rect 36805 2120 36875 2166
rect 36921 2120 36991 2166
rect 37037 2120 37107 2166
rect 37153 2120 37223 2166
rect 37269 2120 37339 2166
rect 37385 2120 37455 2166
rect 37501 2120 37571 2166
rect 37617 2120 37687 2166
rect 37733 2120 37803 2166
rect 37849 2120 37919 2166
rect 37965 2120 38035 2166
rect 38081 2120 38151 2166
rect 38197 2120 38267 2166
rect 38313 2120 38383 2166
rect 38429 2120 38499 2166
rect 38545 2120 38615 2166
rect 38661 2120 38731 2166
rect 38777 2120 38847 2166
rect 38893 2120 38963 2166
rect 39009 2120 39079 2166
rect 39125 2120 39195 2166
rect 39241 2120 39311 2166
rect 39357 2120 39427 2166
rect 39473 2120 39543 2166
rect 39589 2120 39659 2166
rect 39705 2120 39775 2166
rect 39821 2120 39891 2166
rect 39937 2120 40007 2166
rect 40053 2120 40123 2166
rect 40169 2120 40180 2166
rect 28628 2050 40180 2120
rect 28628 2004 28639 2050
rect 28685 2004 28755 2050
rect 28801 2004 28871 2050
rect 28917 2004 28987 2050
rect 29033 2004 29103 2050
rect 29149 2004 29219 2050
rect 29265 2004 29335 2050
rect 29381 2004 29451 2050
rect 29497 2004 29567 2050
rect 29613 2004 29683 2050
rect 29729 2004 29799 2050
rect 29845 2004 29915 2050
rect 29961 2004 30031 2050
rect 30077 2004 30147 2050
rect 30193 2004 30263 2050
rect 30309 2004 30379 2050
rect 30425 2004 30495 2050
rect 30541 2004 30611 2050
rect 30657 2004 30727 2050
rect 30773 2004 30843 2050
rect 30889 2004 30959 2050
rect 31005 2004 31075 2050
rect 31121 2004 31191 2050
rect 31237 2004 31307 2050
rect 31353 2004 31423 2050
rect 31469 2004 31539 2050
rect 31585 2004 31655 2050
rect 31701 2004 31771 2050
rect 31817 2004 31887 2050
rect 31933 2004 32003 2050
rect 32049 2004 32119 2050
rect 32165 2004 32235 2050
rect 32281 2004 32351 2050
rect 32397 2004 32467 2050
rect 32513 2004 32583 2050
rect 32629 2004 32699 2050
rect 32745 2004 32815 2050
rect 32861 2004 32931 2050
rect 32977 2004 33047 2050
rect 33093 2004 33163 2050
rect 33209 2004 33279 2050
rect 33325 2004 33395 2050
rect 33441 2004 33511 2050
rect 33557 2004 33627 2050
rect 33673 2004 33743 2050
rect 33789 2004 33859 2050
rect 33905 2004 33975 2050
rect 34021 2004 34091 2050
rect 34137 2004 34207 2050
rect 34253 2004 34323 2050
rect 34369 2004 34439 2050
rect 34485 2004 34555 2050
rect 34601 2004 34671 2050
rect 34717 2004 34787 2050
rect 34833 2004 34903 2050
rect 34949 2004 35019 2050
rect 35065 2004 35135 2050
rect 35181 2004 35251 2050
rect 35297 2004 35367 2050
rect 35413 2004 35483 2050
rect 35529 2004 35599 2050
rect 35645 2004 35715 2050
rect 35761 2004 35831 2050
rect 35877 2004 35947 2050
rect 35993 2004 36063 2050
rect 36109 2004 36179 2050
rect 36225 2004 36295 2050
rect 36341 2004 36411 2050
rect 36457 2004 36527 2050
rect 36573 2004 36643 2050
rect 36689 2004 36759 2050
rect 36805 2004 36875 2050
rect 36921 2004 36991 2050
rect 37037 2004 37107 2050
rect 37153 2004 37223 2050
rect 37269 2004 37339 2050
rect 37385 2004 37455 2050
rect 37501 2004 37571 2050
rect 37617 2004 37687 2050
rect 37733 2004 37803 2050
rect 37849 2004 37919 2050
rect 37965 2004 38035 2050
rect 38081 2004 38151 2050
rect 38197 2004 38267 2050
rect 38313 2004 38383 2050
rect 38429 2004 38499 2050
rect 38545 2004 38615 2050
rect 38661 2004 38731 2050
rect 38777 2004 38847 2050
rect 38893 2004 38963 2050
rect 39009 2004 39079 2050
rect 39125 2004 39195 2050
rect 39241 2004 39311 2050
rect 39357 2004 39427 2050
rect 39473 2004 39543 2050
rect 39589 2004 39659 2050
rect 39705 2004 39775 2050
rect 39821 2004 39891 2050
rect 39937 2004 40007 2050
rect 40053 2004 40123 2050
rect 40169 2004 40180 2050
rect 28628 1934 40180 2004
rect 28628 1888 28639 1934
rect 28685 1888 28755 1934
rect 28801 1888 28871 1934
rect 28917 1888 28987 1934
rect 29033 1888 29103 1934
rect 29149 1888 29219 1934
rect 29265 1888 29335 1934
rect 29381 1888 29451 1934
rect 29497 1888 29567 1934
rect 29613 1888 29683 1934
rect 29729 1888 29799 1934
rect 29845 1888 29915 1934
rect 29961 1888 30031 1934
rect 30077 1888 30147 1934
rect 30193 1888 30263 1934
rect 30309 1888 30379 1934
rect 30425 1888 30495 1934
rect 30541 1888 30611 1934
rect 30657 1888 30727 1934
rect 30773 1888 30843 1934
rect 30889 1888 30959 1934
rect 31005 1888 31075 1934
rect 31121 1888 31191 1934
rect 31237 1888 31307 1934
rect 31353 1888 31423 1934
rect 31469 1888 31539 1934
rect 31585 1888 31655 1934
rect 31701 1888 31771 1934
rect 31817 1888 31887 1934
rect 31933 1888 32003 1934
rect 32049 1888 32119 1934
rect 32165 1888 32235 1934
rect 32281 1888 32351 1934
rect 32397 1888 32467 1934
rect 32513 1888 32583 1934
rect 32629 1888 32699 1934
rect 32745 1888 32815 1934
rect 32861 1888 32931 1934
rect 32977 1888 33047 1934
rect 33093 1888 33163 1934
rect 33209 1888 33279 1934
rect 33325 1888 33395 1934
rect 33441 1888 33511 1934
rect 33557 1888 33627 1934
rect 33673 1888 33743 1934
rect 33789 1888 33859 1934
rect 33905 1888 33975 1934
rect 34021 1888 34091 1934
rect 34137 1888 34207 1934
rect 34253 1888 34323 1934
rect 34369 1888 34439 1934
rect 34485 1888 34555 1934
rect 34601 1888 34671 1934
rect 34717 1888 34787 1934
rect 34833 1888 34903 1934
rect 34949 1888 35019 1934
rect 35065 1888 35135 1934
rect 35181 1888 35251 1934
rect 35297 1888 35367 1934
rect 35413 1888 35483 1934
rect 35529 1888 35599 1934
rect 35645 1888 35715 1934
rect 35761 1888 35831 1934
rect 35877 1888 35947 1934
rect 35993 1888 36063 1934
rect 36109 1888 36179 1934
rect 36225 1888 36295 1934
rect 36341 1888 36411 1934
rect 36457 1888 36527 1934
rect 36573 1888 36643 1934
rect 36689 1888 36759 1934
rect 36805 1888 36875 1934
rect 36921 1888 36991 1934
rect 37037 1888 37107 1934
rect 37153 1888 37223 1934
rect 37269 1888 37339 1934
rect 37385 1888 37455 1934
rect 37501 1888 37571 1934
rect 37617 1888 37687 1934
rect 37733 1888 37803 1934
rect 37849 1888 37919 1934
rect 37965 1888 38035 1934
rect 38081 1888 38151 1934
rect 38197 1888 38267 1934
rect 38313 1888 38383 1934
rect 38429 1888 38499 1934
rect 38545 1888 38615 1934
rect 38661 1888 38731 1934
rect 38777 1888 38847 1934
rect 38893 1888 38963 1934
rect 39009 1888 39079 1934
rect 39125 1888 39195 1934
rect 39241 1888 39311 1934
rect 39357 1888 39427 1934
rect 39473 1888 39543 1934
rect 39589 1888 39659 1934
rect 39705 1888 39775 1934
rect 39821 1888 39891 1934
rect 39937 1888 40007 1934
rect 40053 1888 40123 1934
rect 40169 1888 40180 1934
rect 28628 1818 40180 1888
rect 28628 1772 28639 1818
rect 28685 1772 28755 1818
rect 28801 1772 28871 1818
rect 28917 1772 28987 1818
rect 29033 1772 29103 1818
rect 29149 1772 29219 1818
rect 29265 1772 29335 1818
rect 29381 1772 29451 1818
rect 29497 1772 29567 1818
rect 29613 1772 29683 1818
rect 29729 1772 29799 1818
rect 29845 1772 29915 1818
rect 29961 1772 30031 1818
rect 30077 1772 30147 1818
rect 30193 1772 30263 1818
rect 30309 1772 30379 1818
rect 30425 1772 30495 1818
rect 30541 1772 30611 1818
rect 30657 1772 30727 1818
rect 30773 1772 30843 1818
rect 30889 1772 30959 1818
rect 31005 1772 31075 1818
rect 31121 1772 31191 1818
rect 31237 1772 31307 1818
rect 31353 1772 31423 1818
rect 31469 1772 31539 1818
rect 31585 1772 31655 1818
rect 31701 1772 31771 1818
rect 31817 1772 31887 1818
rect 31933 1772 32003 1818
rect 32049 1772 32119 1818
rect 32165 1772 32235 1818
rect 32281 1772 32351 1818
rect 32397 1772 32467 1818
rect 32513 1772 32583 1818
rect 32629 1772 32699 1818
rect 32745 1772 32815 1818
rect 32861 1772 32931 1818
rect 32977 1772 33047 1818
rect 33093 1772 33163 1818
rect 33209 1772 33279 1818
rect 33325 1772 33395 1818
rect 33441 1772 33511 1818
rect 33557 1772 33627 1818
rect 33673 1772 33743 1818
rect 33789 1772 33859 1818
rect 33905 1772 33975 1818
rect 34021 1772 34091 1818
rect 34137 1772 34207 1818
rect 34253 1772 34323 1818
rect 34369 1772 34439 1818
rect 34485 1772 34555 1818
rect 34601 1772 34671 1818
rect 34717 1772 34787 1818
rect 34833 1772 34903 1818
rect 34949 1772 35019 1818
rect 35065 1772 35135 1818
rect 35181 1772 35251 1818
rect 35297 1772 35367 1818
rect 35413 1772 35483 1818
rect 35529 1772 35599 1818
rect 35645 1772 35715 1818
rect 35761 1772 35831 1818
rect 35877 1772 35947 1818
rect 35993 1772 36063 1818
rect 36109 1772 36179 1818
rect 36225 1772 36295 1818
rect 36341 1772 36411 1818
rect 36457 1772 36527 1818
rect 36573 1772 36643 1818
rect 36689 1772 36759 1818
rect 36805 1772 36875 1818
rect 36921 1772 36991 1818
rect 37037 1772 37107 1818
rect 37153 1772 37223 1818
rect 37269 1772 37339 1818
rect 37385 1772 37455 1818
rect 37501 1772 37571 1818
rect 37617 1772 37687 1818
rect 37733 1772 37803 1818
rect 37849 1772 37919 1818
rect 37965 1772 38035 1818
rect 38081 1772 38151 1818
rect 38197 1772 38267 1818
rect 38313 1772 38383 1818
rect 38429 1772 38499 1818
rect 38545 1772 38615 1818
rect 38661 1772 38731 1818
rect 38777 1772 38847 1818
rect 38893 1772 38963 1818
rect 39009 1772 39079 1818
rect 39125 1772 39195 1818
rect 39241 1772 39311 1818
rect 39357 1772 39427 1818
rect 39473 1772 39543 1818
rect 39589 1772 39659 1818
rect 39705 1772 39775 1818
rect 39821 1772 39891 1818
rect 39937 1772 40007 1818
rect 40053 1772 40123 1818
rect 40169 1772 40180 1818
rect 28628 1702 40180 1772
rect 28628 1656 28639 1702
rect 28685 1656 28755 1702
rect 28801 1656 28871 1702
rect 28917 1656 28987 1702
rect 29033 1656 29103 1702
rect 29149 1656 29219 1702
rect 29265 1656 29335 1702
rect 29381 1656 29451 1702
rect 29497 1656 29567 1702
rect 29613 1656 29683 1702
rect 29729 1656 29799 1702
rect 29845 1656 29915 1702
rect 29961 1656 30031 1702
rect 30077 1656 30147 1702
rect 30193 1656 30263 1702
rect 30309 1656 30379 1702
rect 30425 1656 30495 1702
rect 30541 1656 30611 1702
rect 30657 1656 30727 1702
rect 30773 1656 30843 1702
rect 30889 1656 30959 1702
rect 31005 1656 31075 1702
rect 31121 1656 31191 1702
rect 31237 1656 31307 1702
rect 31353 1656 31423 1702
rect 31469 1656 31539 1702
rect 31585 1656 31655 1702
rect 31701 1656 31771 1702
rect 31817 1656 31887 1702
rect 31933 1656 32003 1702
rect 32049 1656 32119 1702
rect 32165 1656 32235 1702
rect 32281 1656 32351 1702
rect 32397 1656 32467 1702
rect 32513 1656 32583 1702
rect 32629 1656 32699 1702
rect 32745 1656 32815 1702
rect 32861 1656 32931 1702
rect 32977 1656 33047 1702
rect 33093 1656 33163 1702
rect 33209 1656 33279 1702
rect 33325 1656 33395 1702
rect 33441 1656 33511 1702
rect 33557 1656 33627 1702
rect 33673 1656 33743 1702
rect 33789 1656 33859 1702
rect 33905 1656 33975 1702
rect 34021 1656 34091 1702
rect 34137 1656 34207 1702
rect 34253 1656 34323 1702
rect 34369 1656 34439 1702
rect 34485 1656 34555 1702
rect 34601 1656 34671 1702
rect 34717 1656 34787 1702
rect 34833 1656 34903 1702
rect 34949 1656 35019 1702
rect 35065 1656 35135 1702
rect 35181 1656 35251 1702
rect 35297 1656 35367 1702
rect 35413 1656 35483 1702
rect 35529 1656 35599 1702
rect 35645 1656 35715 1702
rect 35761 1656 35831 1702
rect 35877 1656 35947 1702
rect 35993 1656 36063 1702
rect 36109 1656 36179 1702
rect 36225 1656 36295 1702
rect 36341 1656 36411 1702
rect 36457 1656 36527 1702
rect 36573 1656 36643 1702
rect 36689 1656 36759 1702
rect 36805 1656 36875 1702
rect 36921 1656 36991 1702
rect 37037 1656 37107 1702
rect 37153 1656 37223 1702
rect 37269 1656 37339 1702
rect 37385 1656 37455 1702
rect 37501 1656 37571 1702
rect 37617 1656 37687 1702
rect 37733 1656 37803 1702
rect 37849 1656 37919 1702
rect 37965 1656 38035 1702
rect 38081 1656 38151 1702
rect 38197 1656 38267 1702
rect 38313 1656 38383 1702
rect 38429 1656 38499 1702
rect 38545 1656 38615 1702
rect 38661 1656 38731 1702
rect 38777 1656 38847 1702
rect 38893 1656 38963 1702
rect 39009 1656 39079 1702
rect 39125 1656 39195 1702
rect 39241 1656 39311 1702
rect 39357 1656 39427 1702
rect 39473 1656 39543 1702
rect 39589 1656 39659 1702
rect 39705 1656 39775 1702
rect 39821 1656 39891 1702
rect 39937 1656 40007 1702
rect 40053 1656 40123 1702
rect 40169 1656 40180 1702
rect 28628 1282 40180 1656
rect 50834 3906 56586 3917
rect 50834 3860 50845 3906
rect 50891 3860 50961 3906
rect 51007 3860 51077 3906
rect 51123 3860 51193 3906
rect 51239 3860 51309 3906
rect 51355 3860 51425 3906
rect 51471 3860 51541 3906
rect 51587 3860 51657 3906
rect 51703 3860 51773 3906
rect 51819 3860 51889 3906
rect 51935 3860 52005 3906
rect 52051 3860 52121 3906
rect 52167 3860 52237 3906
rect 52283 3860 52353 3906
rect 52399 3860 52469 3906
rect 52515 3860 52585 3906
rect 52631 3860 52701 3906
rect 52747 3860 52817 3906
rect 52863 3860 52933 3906
rect 52979 3860 53049 3906
rect 53095 3860 53165 3906
rect 53211 3860 53281 3906
rect 53327 3860 53397 3906
rect 53443 3860 53513 3906
rect 53559 3860 53629 3906
rect 53675 3860 53745 3906
rect 53791 3860 53861 3906
rect 53907 3860 53977 3906
rect 54023 3860 54093 3906
rect 54139 3860 54209 3906
rect 54255 3860 54325 3906
rect 54371 3860 54441 3906
rect 54487 3860 54557 3906
rect 54603 3860 54673 3906
rect 54719 3860 54789 3906
rect 54835 3860 54905 3906
rect 54951 3860 55021 3906
rect 55067 3860 55137 3906
rect 55183 3860 55253 3906
rect 55299 3860 55369 3906
rect 55415 3860 55485 3906
rect 55531 3860 55601 3906
rect 55647 3860 55717 3906
rect 55763 3860 55833 3906
rect 55879 3860 55949 3906
rect 55995 3860 56065 3906
rect 56111 3860 56181 3906
rect 56227 3860 56297 3906
rect 56343 3860 56413 3906
rect 56459 3860 56529 3906
rect 56575 3860 56586 3906
rect 50834 3790 56586 3860
rect 50834 3744 50845 3790
rect 50891 3744 50961 3790
rect 51007 3744 51077 3790
rect 51123 3744 51193 3790
rect 51239 3744 51309 3790
rect 51355 3744 51425 3790
rect 51471 3744 51541 3790
rect 51587 3744 51657 3790
rect 51703 3744 51773 3790
rect 51819 3744 51889 3790
rect 51935 3744 52005 3790
rect 52051 3744 52121 3790
rect 52167 3744 52237 3790
rect 52283 3744 52353 3790
rect 52399 3744 52469 3790
rect 52515 3744 52585 3790
rect 52631 3744 52701 3790
rect 52747 3744 52817 3790
rect 52863 3744 52933 3790
rect 52979 3744 53049 3790
rect 53095 3744 53165 3790
rect 53211 3744 53281 3790
rect 53327 3744 53397 3790
rect 53443 3744 53513 3790
rect 53559 3744 53629 3790
rect 53675 3744 53745 3790
rect 53791 3744 53861 3790
rect 53907 3744 53977 3790
rect 54023 3744 54093 3790
rect 54139 3744 54209 3790
rect 54255 3744 54325 3790
rect 54371 3744 54441 3790
rect 54487 3744 54557 3790
rect 54603 3744 54673 3790
rect 54719 3744 54789 3790
rect 54835 3744 54905 3790
rect 54951 3744 55021 3790
rect 55067 3744 55137 3790
rect 55183 3744 55253 3790
rect 55299 3744 55369 3790
rect 55415 3744 55485 3790
rect 55531 3744 55601 3790
rect 55647 3744 55717 3790
rect 55763 3744 55833 3790
rect 55879 3744 55949 3790
rect 55995 3744 56065 3790
rect 56111 3744 56181 3790
rect 56227 3744 56297 3790
rect 56343 3744 56413 3790
rect 56459 3744 56529 3790
rect 56575 3744 56586 3790
rect 50834 3674 56586 3744
rect 50834 3628 50845 3674
rect 50891 3628 50961 3674
rect 51007 3628 51077 3674
rect 51123 3628 51193 3674
rect 51239 3628 51309 3674
rect 51355 3628 51425 3674
rect 51471 3628 51541 3674
rect 51587 3628 51657 3674
rect 51703 3628 51773 3674
rect 51819 3628 51889 3674
rect 51935 3628 52005 3674
rect 52051 3628 52121 3674
rect 52167 3628 52237 3674
rect 52283 3628 52353 3674
rect 52399 3628 52469 3674
rect 52515 3628 52585 3674
rect 52631 3628 52701 3674
rect 52747 3628 52817 3674
rect 52863 3628 52933 3674
rect 52979 3628 53049 3674
rect 53095 3628 53165 3674
rect 53211 3628 53281 3674
rect 53327 3628 53397 3674
rect 53443 3628 53513 3674
rect 53559 3628 53629 3674
rect 53675 3628 53745 3674
rect 53791 3628 53861 3674
rect 53907 3628 53977 3674
rect 54023 3628 54093 3674
rect 54139 3628 54209 3674
rect 54255 3628 54325 3674
rect 54371 3628 54441 3674
rect 54487 3628 54557 3674
rect 54603 3628 54673 3674
rect 54719 3628 54789 3674
rect 54835 3628 54905 3674
rect 54951 3628 55021 3674
rect 55067 3628 55137 3674
rect 55183 3628 55253 3674
rect 55299 3628 55369 3674
rect 55415 3628 55485 3674
rect 55531 3628 55601 3674
rect 55647 3628 55717 3674
rect 55763 3628 55833 3674
rect 55879 3628 55949 3674
rect 55995 3628 56065 3674
rect 56111 3628 56181 3674
rect 56227 3628 56297 3674
rect 56343 3628 56413 3674
rect 56459 3628 56529 3674
rect 56575 3628 56586 3674
rect 50834 3558 56586 3628
rect 50834 3512 50845 3558
rect 50891 3512 50961 3558
rect 51007 3512 51077 3558
rect 51123 3512 51193 3558
rect 51239 3512 51309 3558
rect 51355 3512 51425 3558
rect 51471 3512 51541 3558
rect 51587 3512 51657 3558
rect 51703 3512 51773 3558
rect 51819 3512 51889 3558
rect 51935 3512 52005 3558
rect 52051 3512 52121 3558
rect 52167 3512 52237 3558
rect 52283 3512 52353 3558
rect 52399 3512 52469 3558
rect 52515 3512 52585 3558
rect 52631 3512 52701 3558
rect 52747 3512 52817 3558
rect 52863 3512 52933 3558
rect 52979 3512 53049 3558
rect 53095 3512 53165 3558
rect 53211 3512 53281 3558
rect 53327 3512 53397 3558
rect 53443 3512 53513 3558
rect 53559 3512 53629 3558
rect 53675 3512 53745 3558
rect 53791 3512 53861 3558
rect 53907 3512 53977 3558
rect 54023 3512 54093 3558
rect 54139 3512 54209 3558
rect 54255 3512 54325 3558
rect 54371 3512 54441 3558
rect 54487 3512 54557 3558
rect 54603 3512 54673 3558
rect 54719 3512 54789 3558
rect 54835 3512 54905 3558
rect 54951 3512 55021 3558
rect 55067 3512 55137 3558
rect 55183 3512 55253 3558
rect 55299 3512 55369 3558
rect 55415 3512 55485 3558
rect 55531 3512 55601 3558
rect 55647 3512 55717 3558
rect 55763 3512 55833 3558
rect 55879 3512 55949 3558
rect 55995 3512 56065 3558
rect 56111 3512 56181 3558
rect 56227 3512 56297 3558
rect 56343 3512 56413 3558
rect 56459 3512 56529 3558
rect 56575 3512 56586 3558
rect 50834 3442 56586 3512
rect 50834 3396 50845 3442
rect 50891 3396 50961 3442
rect 51007 3396 51077 3442
rect 51123 3396 51193 3442
rect 51239 3396 51309 3442
rect 51355 3396 51425 3442
rect 51471 3396 51541 3442
rect 51587 3396 51657 3442
rect 51703 3396 51773 3442
rect 51819 3396 51889 3442
rect 51935 3396 52005 3442
rect 52051 3396 52121 3442
rect 52167 3396 52237 3442
rect 52283 3396 52353 3442
rect 52399 3396 52469 3442
rect 52515 3396 52585 3442
rect 52631 3396 52701 3442
rect 52747 3396 52817 3442
rect 52863 3396 52933 3442
rect 52979 3396 53049 3442
rect 53095 3396 53165 3442
rect 53211 3396 53281 3442
rect 53327 3396 53397 3442
rect 53443 3396 53513 3442
rect 53559 3396 53629 3442
rect 53675 3396 53745 3442
rect 53791 3396 53861 3442
rect 53907 3396 53977 3442
rect 54023 3396 54093 3442
rect 54139 3396 54209 3442
rect 54255 3396 54325 3442
rect 54371 3396 54441 3442
rect 54487 3396 54557 3442
rect 54603 3396 54673 3442
rect 54719 3396 54789 3442
rect 54835 3396 54905 3442
rect 54951 3396 55021 3442
rect 55067 3396 55137 3442
rect 55183 3396 55253 3442
rect 55299 3396 55369 3442
rect 55415 3396 55485 3442
rect 55531 3396 55601 3442
rect 55647 3396 55717 3442
rect 55763 3396 55833 3442
rect 55879 3396 55949 3442
rect 55995 3396 56065 3442
rect 56111 3396 56181 3442
rect 56227 3396 56297 3442
rect 56343 3396 56413 3442
rect 56459 3396 56529 3442
rect 56575 3396 56586 3442
rect 50834 3326 56586 3396
rect 50834 3280 50845 3326
rect 50891 3280 50961 3326
rect 51007 3280 51077 3326
rect 51123 3280 51193 3326
rect 51239 3280 51309 3326
rect 51355 3280 51425 3326
rect 51471 3280 51541 3326
rect 51587 3280 51657 3326
rect 51703 3280 51773 3326
rect 51819 3280 51889 3326
rect 51935 3280 52005 3326
rect 52051 3280 52121 3326
rect 52167 3280 52237 3326
rect 52283 3280 52353 3326
rect 52399 3280 52469 3326
rect 52515 3280 52585 3326
rect 52631 3280 52701 3326
rect 52747 3280 52817 3326
rect 52863 3280 52933 3326
rect 52979 3280 53049 3326
rect 53095 3280 53165 3326
rect 53211 3280 53281 3326
rect 53327 3280 53397 3326
rect 53443 3280 53513 3326
rect 53559 3280 53629 3326
rect 53675 3280 53745 3326
rect 53791 3280 53861 3326
rect 53907 3280 53977 3326
rect 54023 3280 54093 3326
rect 54139 3280 54209 3326
rect 54255 3280 54325 3326
rect 54371 3280 54441 3326
rect 54487 3280 54557 3326
rect 54603 3280 54673 3326
rect 54719 3280 54789 3326
rect 54835 3280 54905 3326
rect 54951 3280 55021 3326
rect 55067 3280 55137 3326
rect 55183 3280 55253 3326
rect 55299 3280 55369 3326
rect 55415 3280 55485 3326
rect 55531 3280 55601 3326
rect 55647 3280 55717 3326
rect 55763 3280 55833 3326
rect 55879 3280 55949 3326
rect 55995 3280 56065 3326
rect 56111 3280 56181 3326
rect 56227 3280 56297 3326
rect 56343 3280 56413 3326
rect 56459 3280 56529 3326
rect 56575 3280 56586 3326
rect 50834 3210 56586 3280
rect 50834 3164 50845 3210
rect 50891 3164 50961 3210
rect 51007 3164 51077 3210
rect 51123 3164 51193 3210
rect 51239 3164 51309 3210
rect 51355 3164 51425 3210
rect 51471 3164 51541 3210
rect 51587 3164 51657 3210
rect 51703 3164 51773 3210
rect 51819 3164 51889 3210
rect 51935 3164 52005 3210
rect 52051 3164 52121 3210
rect 52167 3164 52237 3210
rect 52283 3164 52353 3210
rect 52399 3164 52469 3210
rect 52515 3164 52585 3210
rect 52631 3164 52701 3210
rect 52747 3164 52817 3210
rect 52863 3164 52933 3210
rect 52979 3164 53049 3210
rect 53095 3164 53165 3210
rect 53211 3164 53281 3210
rect 53327 3164 53397 3210
rect 53443 3164 53513 3210
rect 53559 3164 53629 3210
rect 53675 3164 53745 3210
rect 53791 3164 53861 3210
rect 53907 3164 53977 3210
rect 54023 3164 54093 3210
rect 54139 3164 54209 3210
rect 54255 3164 54325 3210
rect 54371 3164 54441 3210
rect 54487 3164 54557 3210
rect 54603 3164 54673 3210
rect 54719 3164 54789 3210
rect 54835 3164 54905 3210
rect 54951 3164 55021 3210
rect 55067 3164 55137 3210
rect 55183 3164 55253 3210
rect 55299 3164 55369 3210
rect 55415 3164 55485 3210
rect 55531 3164 55601 3210
rect 55647 3164 55717 3210
rect 55763 3164 55833 3210
rect 55879 3164 55949 3210
rect 55995 3164 56065 3210
rect 56111 3164 56181 3210
rect 56227 3164 56297 3210
rect 56343 3164 56413 3210
rect 56459 3164 56529 3210
rect 56575 3164 56586 3210
rect 50834 3094 56586 3164
rect 50834 3048 50845 3094
rect 50891 3048 50961 3094
rect 51007 3048 51077 3094
rect 51123 3048 51193 3094
rect 51239 3048 51309 3094
rect 51355 3048 51425 3094
rect 51471 3048 51541 3094
rect 51587 3048 51657 3094
rect 51703 3048 51773 3094
rect 51819 3048 51889 3094
rect 51935 3048 52005 3094
rect 52051 3048 52121 3094
rect 52167 3048 52237 3094
rect 52283 3048 52353 3094
rect 52399 3048 52469 3094
rect 52515 3048 52585 3094
rect 52631 3048 52701 3094
rect 52747 3048 52817 3094
rect 52863 3048 52933 3094
rect 52979 3048 53049 3094
rect 53095 3048 53165 3094
rect 53211 3048 53281 3094
rect 53327 3048 53397 3094
rect 53443 3048 53513 3094
rect 53559 3048 53629 3094
rect 53675 3048 53745 3094
rect 53791 3048 53861 3094
rect 53907 3048 53977 3094
rect 54023 3048 54093 3094
rect 54139 3048 54209 3094
rect 54255 3048 54325 3094
rect 54371 3048 54441 3094
rect 54487 3048 54557 3094
rect 54603 3048 54673 3094
rect 54719 3048 54789 3094
rect 54835 3048 54905 3094
rect 54951 3048 55021 3094
rect 55067 3048 55137 3094
rect 55183 3048 55253 3094
rect 55299 3048 55369 3094
rect 55415 3048 55485 3094
rect 55531 3048 55601 3094
rect 55647 3048 55717 3094
rect 55763 3048 55833 3094
rect 55879 3048 55949 3094
rect 55995 3048 56065 3094
rect 56111 3048 56181 3094
rect 56227 3048 56297 3094
rect 56343 3048 56413 3094
rect 56459 3048 56529 3094
rect 56575 3048 56586 3094
rect 50834 2978 56586 3048
rect 50834 2932 50845 2978
rect 50891 2932 50961 2978
rect 51007 2932 51077 2978
rect 51123 2932 51193 2978
rect 51239 2932 51309 2978
rect 51355 2932 51425 2978
rect 51471 2932 51541 2978
rect 51587 2932 51657 2978
rect 51703 2932 51773 2978
rect 51819 2932 51889 2978
rect 51935 2932 52005 2978
rect 52051 2932 52121 2978
rect 52167 2932 52237 2978
rect 52283 2932 52353 2978
rect 52399 2932 52469 2978
rect 52515 2932 52585 2978
rect 52631 2932 52701 2978
rect 52747 2932 52817 2978
rect 52863 2932 52933 2978
rect 52979 2932 53049 2978
rect 53095 2932 53165 2978
rect 53211 2932 53281 2978
rect 53327 2932 53397 2978
rect 53443 2932 53513 2978
rect 53559 2932 53629 2978
rect 53675 2932 53745 2978
rect 53791 2932 53861 2978
rect 53907 2932 53977 2978
rect 54023 2932 54093 2978
rect 54139 2932 54209 2978
rect 54255 2932 54325 2978
rect 54371 2932 54441 2978
rect 54487 2932 54557 2978
rect 54603 2932 54673 2978
rect 54719 2932 54789 2978
rect 54835 2932 54905 2978
rect 54951 2932 55021 2978
rect 55067 2932 55137 2978
rect 55183 2932 55253 2978
rect 55299 2932 55369 2978
rect 55415 2932 55485 2978
rect 55531 2932 55601 2978
rect 55647 2932 55717 2978
rect 55763 2932 55833 2978
rect 55879 2932 55949 2978
rect 55995 2932 56065 2978
rect 56111 2932 56181 2978
rect 56227 2932 56297 2978
rect 56343 2932 56413 2978
rect 56459 2932 56529 2978
rect 56575 2932 56586 2978
rect 50834 2862 56586 2932
rect 50834 2816 50845 2862
rect 50891 2816 50961 2862
rect 51007 2816 51077 2862
rect 51123 2816 51193 2862
rect 51239 2816 51309 2862
rect 51355 2816 51425 2862
rect 51471 2816 51541 2862
rect 51587 2816 51657 2862
rect 51703 2816 51773 2862
rect 51819 2816 51889 2862
rect 51935 2816 52005 2862
rect 52051 2816 52121 2862
rect 52167 2816 52237 2862
rect 52283 2816 52353 2862
rect 52399 2816 52469 2862
rect 52515 2816 52585 2862
rect 52631 2816 52701 2862
rect 52747 2816 52817 2862
rect 52863 2816 52933 2862
rect 52979 2816 53049 2862
rect 53095 2816 53165 2862
rect 53211 2816 53281 2862
rect 53327 2816 53397 2862
rect 53443 2816 53513 2862
rect 53559 2816 53629 2862
rect 53675 2816 53745 2862
rect 53791 2816 53861 2862
rect 53907 2816 53977 2862
rect 54023 2816 54093 2862
rect 54139 2816 54209 2862
rect 54255 2816 54325 2862
rect 54371 2816 54441 2862
rect 54487 2816 54557 2862
rect 54603 2816 54673 2862
rect 54719 2816 54789 2862
rect 54835 2816 54905 2862
rect 54951 2816 55021 2862
rect 55067 2816 55137 2862
rect 55183 2816 55253 2862
rect 55299 2816 55369 2862
rect 55415 2816 55485 2862
rect 55531 2816 55601 2862
rect 55647 2816 55717 2862
rect 55763 2816 55833 2862
rect 55879 2816 55949 2862
rect 55995 2816 56065 2862
rect 56111 2816 56181 2862
rect 56227 2816 56297 2862
rect 56343 2816 56413 2862
rect 56459 2816 56529 2862
rect 56575 2816 56586 2862
rect 50834 2746 56586 2816
rect 50834 2700 50845 2746
rect 50891 2700 50961 2746
rect 51007 2700 51077 2746
rect 51123 2700 51193 2746
rect 51239 2700 51309 2746
rect 51355 2700 51425 2746
rect 51471 2700 51541 2746
rect 51587 2700 51657 2746
rect 51703 2700 51773 2746
rect 51819 2700 51889 2746
rect 51935 2700 52005 2746
rect 52051 2700 52121 2746
rect 52167 2700 52237 2746
rect 52283 2700 52353 2746
rect 52399 2700 52469 2746
rect 52515 2700 52585 2746
rect 52631 2700 52701 2746
rect 52747 2700 52817 2746
rect 52863 2700 52933 2746
rect 52979 2700 53049 2746
rect 53095 2700 53165 2746
rect 53211 2700 53281 2746
rect 53327 2700 53397 2746
rect 53443 2700 53513 2746
rect 53559 2700 53629 2746
rect 53675 2700 53745 2746
rect 53791 2700 53861 2746
rect 53907 2700 53977 2746
rect 54023 2700 54093 2746
rect 54139 2700 54209 2746
rect 54255 2700 54325 2746
rect 54371 2700 54441 2746
rect 54487 2700 54557 2746
rect 54603 2700 54673 2746
rect 54719 2700 54789 2746
rect 54835 2700 54905 2746
rect 54951 2700 55021 2746
rect 55067 2700 55137 2746
rect 55183 2700 55253 2746
rect 55299 2700 55369 2746
rect 55415 2700 55485 2746
rect 55531 2700 55601 2746
rect 55647 2700 55717 2746
rect 55763 2700 55833 2746
rect 55879 2700 55949 2746
rect 55995 2700 56065 2746
rect 56111 2700 56181 2746
rect 56227 2700 56297 2746
rect 56343 2700 56413 2746
rect 56459 2700 56529 2746
rect 56575 2700 56586 2746
rect 50834 2630 56586 2700
rect 50834 2584 50845 2630
rect 50891 2584 50961 2630
rect 51007 2584 51077 2630
rect 51123 2584 51193 2630
rect 51239 2584 51309 2630
rect 51355 2584 51425 2630
rect 51471 2584 51541 2630
rect 51587 2584 51657 2630
rect 51703 2584 51773 2630
rect 51819 2584 51889 2630
rect 51935 2584 52005 2630
rect 52051 2584 52121 2630
rect 52167 2584 52237 2630
rect 52283 2584 52353 2630
rect 52399 2584 52469 2630
rect 52515 2584 52585 2630
rect 52631 2584 52701 2630
rect 52747 2584 52817 2630
rect 52863 2584 52933 2630
rect 52979 2584 53049 2630
rect 53095 2584 53165 2630
rect 53211 2584 53281 2630
rect 53327 2584 53397 2630
rect 53443 2584 53513 2630
rect 53559 2584 53629 2630
rect 53675 2584 53745 2630
rect 53791 2584 53861 2630
rect 53907 2584 53977 2630
rect 54023 2584 54093 2630
rect 54139 2584 54209 2630
rect 54255 2584 54325 2630
rect 54371 2584 54441 2630
rect 54487 2584 54557 2630
rect 54603 2584 54673 2630
rect 54719 2584 54789 2630
rect 54835 2584 54905 2630
rect 54951 2584 55021 2630
rect 55067 2584 55137 2630
rect 55183 2584 55253 2630
rect 55299 2584 55369 2630
rect 55415 2584 55485 2630
rect 55531 2584 55601 2630
rect 55647 2584 55717 2630
rect 55763 2584 55833 2630
rect 55879 2584 55949 2630
rect 55995 2584 56065 2630
rect 56111 2584 56181 2630
rect 56227 2584 56297 2630
rect 56343 2584 56413 2630
rect 56459 2584 56529 2630
rect 56575 2584 56586 2630
rect 50834 2514 56586 2584
rect 50834 2468 50845 2514
rect 50891 2468 50961 2514
rect 51007 2468 51077 2514
rect 51123 2468 51193 2514
rect 51239 2468 51309 2514
rect 51355 2468 51425 2514
rect 51471 2468 51541 2514
rect 51587 2468 51657 2514
rect 51703 2468 51773 2514
rect 51819 2468 51889 2514
rect 51935 2468 52005 2514
rect 52051 2468 52121 2514
rect 52167 2468 52237 2514
rect 52283 2468 52353 2514
rect 52399 2468 52469 2514
rect 52515 2468 52585 2514
rect 52631 2468 52701 2514
rect 52747 2468 52817 2514
rect 52863 2468 52933 2514
rect 52979 2468 53049 2514
rect 53095 2468 53165 2514
rect 53211 2468 53281 2514
rect 53327 2468 53397 2514
rect 53443 2468 53513 2514
rect 53559 2468 53629 2514
rect 53675 2468 53745 2514
rect 53791 2468 53861 2514
rect 53907 2468 53977 2514
rect 54023 2468 54093 2514
rect 54139 2468 54209 2514
rect 54255 2468 54325 2514
rect 54371 2468 54441 2514
rect 54487 2468 54557 2514
rect 54603 2468 54673 2514
rect 54719 2468 54789 2514
rect 54835 2468 54905 2514
rect 54951 2468 55021 2514
rect 55067 2468 55137 2514
rect 55183 2468 55253 2514
rect 55299 2468 55369 2514
rect 55415 2468 55485 2514
rect 55531 2468 55601 2514
rect 55647 2468 55717 2514
rect 55763 2468 55833 2514
rect 55879 2468 55949 2514
rect 55995 2468 56065 2514
rect 56111 2468 56181 2514
rect 56227 2468 56297 2514
rect 56343 2468 56413 2514
rect 56459 2468 56529 2514
rect 56575 2468 56586 2514
rect 50834 2398 56586 2468
rect 50834 2352 50845 2398
rect 50891 2352 50961 2398
rect 51007 2352 51077 2398
rect 51123 2352 51193 2398
rect 51239 2352 51309 2398
rect 51355 2352 51425 2398
rect 51471 2352 51541 2398
rect 51587 2352 51657 2398
rect 51703 2352 51773 2398
rect 51819 2352 51889 2398
rect 51935 2352 52005 2398
rect 52051 2352 52121 2398
rect 52167 2352 52237 2398
rect 52283 2352 52353 2398
rect 52399 2352 52469 2398
rect 52515 2352 52585 2398
rect 52631 2352 52701 2398
rect 52747 2352 52817 2398
rect 52863 2352 52933 2398
rect 52979 2352 53049 2398
rect 53095 2352 53165 2398
rect 53211 2352 53281 2398
rect 53327 2352 53397 2398
rect 53443 2352 53513 2398
rect 53559 2352 53629 2398
rect 53675 2352 53745 2398
rect 53791 2352 53861 2398
rect 53907 2352 53977 2398
rect 54023 2352 54093 2398
rect 54139 2352 54209 2398
rect 54255 2352 54325 2398
rect 54371 2352 54441 2398
rect 54487 2352 54557 2398
rect 54603 2352 54673 2398
rect 54719 2352 54789 2398
rect 54835 2352 54905 2398
rect 54951 2352 55021 2398
rect 55067 2352 55137 2398
rect 55183 2352 55253 2398
rect 55299 2352 55369 2398
rect 55415 2352 55485 2398
rect 55531 2352 55601 2398
rect 55647 2352 55717 2398
rect 55763 2352 55833 2398
rect 55879 2352 55949 2398
rect 55995 2352 56065 2398
rect 56111 2352 56181 2398
rect 56227 2352 56297 2398
rect 56343 2352 56413 2398
rect 56459 2352 56529 2398
rect 56575 2352 56586 2398
rect 50834 2282 56586 2352
rect 50834 2236 50845 2282
rect 50891 2236 50961 2282
rect 51007 2236 51077 2282
rect 51123 2236 51193 2282
rect 51239 2236 51309 2282
rect 51355 2236 51425 2282
rect 51471 2236 51541 2282
rect 51587 2236 51657 2282
rect 51703 2236 51773 2282
rect 51819 2236 51889 2282
rect 51935 2236 52005 2282
rect 52051 2236 52121 2282
rect 52167 2236 52237 2282
rect 52283 2236 52353 2282
rect 52399 2236 52469 2282
rect 52515 2236 52585 2282
rect 52631 2236 52701 2282
rect 52747 2236 52817 2282
rect 52863 2236 52933 2282
rect 52979 2236 53049 2282
rect 53095 2236 53165 2282
rect 53211 2236 53281 2282
rect 53327 2236 53397 2282
rect 53443 2236 53513 2282
rect 53559 2236 53629 2282
rect 53675 2236 53745 2282
rect 53791 2236 53861 2282
rect 53907 2236 53977 2282
rect 54023 2236 54093 2282
rect 54139 2236 54209 2282
rect 54255 2236 54325 2282
rect 54371 2236 54441 2282
rect 54487 2236 54557 2282
rect 54603 2236 54673 2282
rect 54719 2236 54789 2282
rect 54835 2236 54905 2282
rect 54951 2236 55021 2282
rect 55067 2236 55137 2282
rect 55183 2236 55253 2282
rect 55299 2236 55369 2282
rect 55415 2236 55485 2282
rect 55531 2236 55601 2282
rect 55647 2236 55717 2282
rect 55763 2236 55833 2282
rect 55879 2236 55949 2282
rect 55995 2236 56065 2282
rect 56111 2236 56181 2282
rect 56227 2236 56297 2282
rect 56343 2236 56413 2282
rect 56459 2236 56529 2282
rect 56575 2236 56586 2282
rect 50834 2166 56586 2236
rect 50834 2120 50845 2166
rect 50891 2120 50961 2166
rect 51007 2120 51077 2166
rect 51123 2120 51193 2166
rect 51239 2120 51309 2166
rect 51355 2120 51425 2166
rect 51471 2120 51541 2166
rect 51587 2120 51657 2166
rect 51703 2120 51773 2166
rect 51819 2120 51889 2166
rect 51935 2120 52005 2166
rect 52051 2120 52121 2166
rect 52167 2120 52237 2166
rect 52283 2120 52353 2166
rect 52399 2120 52469 2166
rect 52515 2120 52585 2166
rect 52631 2120 52701 2166
rect 52747 2120 52817 2166
rect 52863 2120 52933 2166
rect 52979 2120 53049 2166
rect 53095 2120 53165 2166
rect 53211 2120 53281 2166
rect 53327 2120 53397 2166
rect 53443 2120 53513 2166
rect 53559 2120 53629 2166
rect 53675 2120 53745 2166
rect 53791 2120 53861 2166
rect 53907 2120 53977 2166
rect 54023 2120 54093 2166
rect 54139 2120 54209 2166
rect 54255 2120 54325 2166
rect 54371 2120 54441 2166
rect 54487 2120 54557 2166
rect 54603 2120 54673 2166
rect 54719 2120 54789 2166
rect 54835 2120 54905 2166
rect 54951 2120 55021 2166
rect 55067 2120 55137 2166
rect 55183 2120 55253 2166
rect 55299 2120 55369 2166
rect 55415 2120 55485 2166
rect 55531 2120 55601 2166
rect 55647 2120 55717 2166
rect 55763 2120 55833 2166
rect 55879 2120 55949 2166
rect 55995 2120 56065 2166
rect 56111 2120 56181 2166
rect 56227 2120 56297 2166
rect 56343 2120 56413 2166
rect 56459 2120 56529 2166
rect 56575 2120 56586 2166
rect 50834 2050 56586 2120
rect 50834 2004 50845 2050
rect 50891 2004 50961 2050
rect 51007 2004 51077 2050
rect 51123 2004 51193 2050
rect 51239 2004 51309 2050
rect 51355 2004 51425 2050
rect 51471 2004 51541 2050
rect 51587 2004 51657 2050
rect 51703 2004 51773 2050
rect 51819 2004 51889 2050
rect 51935 2004 52005 2050
rect 52051 2004 52121 2050
rect 52167 2004 52237 2050
rect 52283 2004 52353 2050
rect 52399 2004 52469 2050
rect 52515 2004 52585 2050
rect 52631 2004 52701 2050
rect 52747 2004 52817 2050
rect 52863 2004 52933 2050
rect 52979 2004 53049 2050
rect 53095 2004 53165 2050
rect 53211 2004 53281 2050
rect 53327 2004 53397 2050
rect 53443 2004 53513 2050
rect 53559 2004 53629 2050
rect 53675 2004 53745 2050
rect 53791 2004 53861 2050
rect 53907 2004 53977 2050
rect 54023 2004 54093 2050
rect 54139 2004 54209 2050
rect 54255 2004 54325 2050
rect 54371 2004 54441 2050
rect 54487 2004 54557 2050
rect 54603 2004 54673 2050
rect 54719 2004 54789 2050
rect 54835 2004 54905 2050
rect 54951 2004 55021 2050
rect 55067 2004 55137 2050
rect 55183 2004 55253 2050
rect 55299 2004 55369 2050
rect 55415 2004 55485 2050
rect 55531 2004 55601 2050
rect 55647 2004 55717 2050
rect 55763 2004 55833 2050
rect 55879 2004 55949 2050
rect 55995 2004 56065 2050
rect 56111 2004 56181 2050
rect 56227 2004 56297 2050
rect 56343 2004 56413 2050
rect 56459 2004 56529 2050
rect 56575 2004 56586 2050
rect 50834 1934 56586 2004
rect 50834 1888 50845 1934
rect 50891 1888 50961 1934
rect 51007 1888 51077 1934
rect 51123 1888 51193 1934
rect 51239 1888 51309 1934
rect 51355 1888 51425 1934
rect 51471 1888 51541 1934
rect 51587 1888 51657 1934
rect 51703 1888 51773 1934
rect 51819 1888 51889 1934
rect 51935 1888 52005 1934
rect 52051 1888 52121 1934
rect 52167 1888 52237 1934
rect 52283 1888 52353 1934
rect 52399 1888 52469 1934
rect 52515 1888 52585 1934
rect 52631 1888 52701 1934
rect 52747 1888 52817 1934
rect 52863 1888 52933 1934
rect 52979 1888 53049 1934
rect 53095 1888 53165 1934
rect 53211 1888 53281 1934
rect 53327 1888 53397 1934
rect 53443 1888 53513 1934
rect 53559 1888 53629 1934
rect 53675 1888 53745 1934
rect 53791 1888 53861 1934
rect 53907 1888 53977 1934
rect 54023 1888 54093 1934
rect 54139 1888 54209 1934
rect 54255 1888 54325 1934
rect 54371 1888 54441 1934
rect 54487 1888 54557 1934
rect 54603 1888 54673 1934
rect 54719 1888 54789 1934
rect 54835 1888 54905 1934
rect 54951 1888 55021 1934
rect 55067 1888 55137 1934
rect 55183 1888 55253 1934
rect 55299 1888 55369 1934
rect 55415 1888 55485 1934
rect 55531 1888 55601 1934
rect 55647 1888 55717 1934
rect 55763 1888 55833 1934
rect 55879 1888 55949 1934
rect 55995 1888 56065 1934
rect 56111 1888 56181 1934
rect 56227 1888 56297 1934
rect 56343 1888 56413 1934
rect 56459 1888 56529 1934
rect 56575 1888 56586 1934
rect 50834 1818 56586 1888
rect 50834 1772 50845 1818
rect 50891 1772 50961 1818
rect 51007 1772 51077 1818
rect 51123 1772 51193 1818
rect 51239 1772 51309 1818
rect 51355 1772 51425 1818
rect 51471 1772 51541 1818
rect 51587 1772 51657 1818
rect 51703 1772 51773 1818
rect 51819 1772 51889 1818
rect 51935 1772 52005 1818
rect 52051 1772 52121 1818
rect 52167 1772 52237 1818
rect 52283 1772 52353 1818
rect 52399 1772 52469 1818
rect 52515 1772 52585 1818
rect 52631 1772 52701 1818
rect 52747 1772 52817 1818
rect 52863 1772 52933 1818
rect 52979 1772 53049 1818
rect 53095 1772 53165 1818
rect 53211 1772 53281 1818
rect 53327 1772 53397 1818
rect 53443 1772 53513 1818
rect 53559 1772 53629 1818
rect 53675 1772 53745 1818
rect 53791 1772 53861 1818
rect 53907 1772 53977 1818
rect 54023 1772 54093 1818
rect 54139 1772 54209 1818
rect 54255 1772 54325 1818
rect 54371 1772 54441 1818
rect 54487 1772 54557 1818
rect 54603 1772 54673 1818
rect 54719 1772 54789 1818
rect 54835 1772 54905 1818
rect 54951 1772 55021 1818
rect 55067 1772 55137 1818
rect 55183 1772 55253 1818
rect 55299 1772 55369 1818
rect 55415 1772 55485 1818
rect 55531 1772 55601 1818
rect 55647 1772 55717 1818
rect 55763 1772 55833 1818
rect 55879 1772 55949 1818
rect 55995 1772 56065 1818
rect 56111 1772 56181 1818
rect 56227 1772 56297 1818
rect 56343 1772 56413 1818
rect 56459 1772 56529 1818
rect 56575 1772 56586 1818
rect 50834 1702 56586 1772
rect 50834 1656 50845 1702
rect 50891 1656 50961 1702
rect 51007 1656 51077 1702
rect 51123 1656 51193 1702
rect 51239 1656 51309 1702
rect 51355 1656 51425 1702
rect 51471 1656 51541 1702
rect 51587 1656 51657 1702
rect 51703 1656 51773 1702
rect 51819 1656 51889 1702
rect 51935 1656 52005 1702
rect 52051 1656 52121 1702
rect 52167 1656 52237 1702
rect 52283 1656 52353 1702
rect 52399 1656 52469 1702
rect 52515 1656 52585 1702
rect 52631 1656 52701 1702
rect 52747 1656 52817 1702
rect 52863 1656 52933 1702
rect 52979 1656 53049 1702
rect 53095 1656 53165 1702
rect 53211 1656 53281 1702
rect 53327 1656 53397 1702
rect 53443 1656 53513 1702
rect 53559 1656 53629 1702
rect 53675 1656 53745 1702
rect 53791 1656 53861 1702
rect 53907 1656 53977 1702
rect 54023 1656 54093 1702
rect 54139 1656 54209 1702
rect 54255 1656 54325 1702
rect 54371 1656 54441 1702
rect 54487 1656 54557 1702
rect 54603 1656 54673 1702
rect 54719 1656 54789 1702
rect 54835 1656 54905 1702
rect 54951 1656 55021 1702
rect 55067 1656 55137 1702
rect 55183 1656 55253 1702
rect 55299 1656 55369 1702
rect 55415 1656 55485 1702
rect 55531 1656 55601 1702
rect 55647 1656 55717 1702
rect 55763 1656 55833 1702
rect 55879 1656 55949 1702
rect 55995 1656 56065 1702
rect 56111 1656 56181 1702
rect 56227 1656 56297 1702
rect 56343 1656 56413 1702
rect 56459 1656 56529 1702
rect 56575 1656 56586 1702
rect 50834 1282 56586 1656
rect 57295 1282 57380 4728
rect 57626 5220 57736 5306
rect 57909 33432 58351 33519
rect 57909 33380 57998 33432
rect 58050 33380 58210 33432
rect 58262 33380 58351 33432
rect 57909 33215 58351 33380
rect 57909 33163 57998 33215
rect 58050 33163 58210 33215
rect 58262 33163 58351 33215
rect 57909 32997 58351 33163
rect 57909 32945 57998 32997
rect 58050 32945 58210 32997
rect 58262 32945 58351 32997
rect 57909 32779 58351 32945
rect 57909 32727 57998 32779
rect 58050 32727 58210 32779
rect 58262 32727 58351 32779
rect 57909 32562 58351 32727
rect 57909 32510 57998 32562
rect 58050 32510 58210 32562
rect 58262 32510 58351 32562
rect 57909 32344 58351 32510
rect 57909 32292 57998 32344
rect 58050 32292 58210 32344
rect 58262 32292 58351 32344
rect 57909 32127 58351 32292
rect 57909 32075 57998 32127
rect 58050 32075 58210 32127
rect 58262 32075 58351 32127
rect 57909 31909 58351 32075
rect 83398 32048 83834 32122
rect 57909 31857 57998 31909
rect 58050 31857 58210 31909
rect 58262 31857 58351 31909
rect 57909 31691 58351 31857
rect 57909 31639 57998 31691
rect 58050 31639 58210 31691
rect 58262 31639 58351 31691
rect 57909 31474 58351 31639
rect 57909 31422 57998 31474
rect 58050 31422 58210 31474
rect 58262 31422 58351 31474
rect 57909 31256 58351 31422
rect 57909 31204 57998 31256
rect 58050 31204 58210 31256
rect 58262 31204 58351 31256
rect 57909 31038 58351 31204
rect 57909 30986 57998 31038
rect 58050 30986 58210 31038
rect 58262 30986 58351 31038
rect 57909 30821 58351 30986
rect 57909 30769 57998 30821
rect 58050 30769 58210 30821
rect 58262 30769 58351 30821
rect 57909 30603 58351 30769
rect 57909 30551 57998 30603
rect 58050 30551 58210 30603
rect 58262 30551 58351 30603
rect 57909 30386 58351 30551
rect 57909 30334 57998 30386
rect 58050 30334 58210 30386
rect 58262 30334 58351 30386
rect 57909 30168 58351 30334
rect 57909 30116 57998 30168
rect 58050 30116 58210 30168
rect 58262 30116 58351 30168
rect 57909 29950 58351 30116
rect 57909 29898 57998 29950
rect 58050 29898 58210 29950
rect 58262 29898 58351 29950
rect 57909 29733 58351 29898
rect 57909 29681 57998 29733
rect 58050 29681 58210 29733
rect 58262 29681 58351 29733
rect 57909 29515 58351 29681
rect 57909 29463 57998 29515
rect 58050 29463 58210 29515
rect 58262 29463 58351 29515
rect 57909 29297 58351 29463
rect 57909 29245 57998 29297
rect 58050 29245 58210 29297
rect 58262 29245 58351 29297
rect 57909 29080 58351 29245
rect 57909 29028 57998 29080
rect 58050 29028 58210 29080
rect 58262 29028 58351 29080
rect 57909 28862 58351 29028
rect 57909 28810 57998 28862
rect 58050 28810 58210 28862
rect 58262 28810 58351 28862
rect 57909 28644 58351 28810
rect 57909 28592 57998 28644
rect 58050 28592 58210 28644
rect 58262 28592 58351 28644
rect 57909 28427 58351 28592
rect 57909 28375 57998 28427
rect 58050 28375 58210 28427
rect 58262 28375 58351 28427
rect 57909 28209 58351 28375
rect 57909 28157 57998 28209
rect 58050 28157 58210 28209
rect 58262 28157 58351 28209
rect 57909 27992 58351 28157
rect 57909 27940 57998 27992
rect 58050 27940 58210 27992
rect 58262 27940 58351 27992
rect 57909 27774 58351 27940
rect 57909 27722 57998 27774
rect 58050 27722 58210 27774
rect 58262 27722 58351 27774
rect 57909 27556 58351 27722
rect 57909 27504 57998 27556
rect 58050 27504 58210 27556
rect 58262 27504 58351 27556
rect 57909 27339 58351 27504
rect 57909 27287 57998 27339
rect 58050 27287 58210 27339
rect 58262 27287 58351 27339
rect 57909 27121 58351 27287
rect 57909 27069 57998 27121
rect 58050 27069 58210 27121
rect 58262 27069 58351 27121
rect 57909 26903 58351 27069
rect 57909 26851 57998 26903
rect 58050 26851 58210 26903
rect 58262 26851 58351 26903
rect 57909 26686 58351 26851
rect 57909 26634 57998 26686
rect 58050 26634 58210 26686
rect 58262 26634 58351 26686
rect 57909 26468 58351 26634
rect 57909 26416 57998 26468
rect 58050 26416 58210 26468
rect 58262 26416 58351 26468
rect 57909 26250 58351 26416
rect 57909 26198 57998 26250
rect 58050 26198 58210 26250
rect 58262 26198 58351 26250
rect 57909 26033 58351 26198
rect 57909 25981 57998 26033
rect 58050 25981 58210 26033
rect 58262 25981 58351 26033
rect 57909 25815 58351 25981
rect 57909 25763 57998 25815
rect 58050 25763 58210 25815
rect 58262 25763 58351 25815
rect 57909 25598 58351 25763
rect 57909 25546 57998 25598
rect 58050 25546 58210 25598
rect 58262 25546 58351 25598
rect 57909 25380 58351 25546
rect 57909 25328 57998 25380
rect 58050 25328 58210 25380
rect 58262 25328 58351 25380
rect 57909 25162 58351 25328
rect 57909 25110 57998 25162
rect 58050 25110 58210 25162
rect 58262 25110 58351 25162
rect 57909 24945 58351 25110
rect 57909 24893 57998 24945
rect 58050 24893 58210 24945
rect 58262 24893 58351 24945
rect 57909 24727 58351 24893
rect 57909 24675 57998 24727
rect 58050 24675 58210 24727
rect 58262 24675 58351 24727
rect 57909 24509 58351 24675
rect 57909 24457 57998 24509
rect 58050 24457 58210 24509
rect 58262 24457 58351 24509
rect 57909 24292 58351 24457
rect 57909 24240 57998 24292
rect 58050 24240 58210 24292
rect 58262 24240 58351 24292
rect 57909 24074 58351 24240
rect 57909 24022 57998 24074
rect 58050 24022 58210 24074
rect 58262 24022 58351 24074
rect 57909 23857 58351 24022
rect 57909 23805 57998 23857
rect 58050 23805 58210 23857
rect 58262 23805 58351 23857
rect 57909 23639 58351 23805
rect 57909 23587 57998 23639
rect 58050 23587 58210 23639
rect 58262 23587 58351 23639
rect 57909 23421 58351 23587
rect 57909 23369 57998 23421
rect 58050 23369 58210 23421
rect 58262 23369 58351 23421
rect 57909 23204 58351 23369
rect 57909 23152 57998 23204
rect 58050 23152 58210 23204
rect 58262 23152 58351 23204
rect 57909 22986 58351 23152
rect 57909 22934 57998 22986
rect 58050 22934 58210 22986
rect 58262 22934 58351 22986
rect 57909 22768 58351 22934
rect 57909 22716 57998 22768
rect 58050 22716 58210 22768
rect 58262 22716 58351 22768
rect 57909 22551 58351 22716
rect 57909 22499 57998 22551
rect 58050 22499 58210 22551
rect 58262 22499 58351 22551
rect 57909 22333 58351 22499
rect 57909 22281 57998 22333
rect 58050 22281 58210 22333
rect 58262 22281 58351 22333
rect 57909 22115 58351 22281
rect 57909 22063 57998 22115
rect 58050 22063 58210 22115
rect 58262 22063 58351 22115
rect 57909 21898 58351 22063
rect 57909 21846 57998 21898
rect 58050 21846 58210 21898
rect 58262 21846 58351 21898
rect 57909 21680 58351 21846
rect 57909 21628 57998 21680
rect 58050 21628 58210 21680
rect 58262 21628 58351 21680
rect 57909 21463 58351 21628
rect 57909 21411 57998 21463
rect 58050 21411 58210 21463
rect 58262 21411 58351 21463
rect 57909 21245 58351 21411
rect 57909 21193 57998 21245
rect 58050 21193 58210 21245
rect 58262 21193 58351 21245
rect 57909 21027 58351 21193
rect 57909 20975 57998 21027
rect 58050 20975 58210 21027
rect 58262 20975 58351 21027
rect 57909 20810 58351 20975
rect 57909 20758 57998 20810
rect 58050 20758 58210 20810
rect 58262 20758 58351 20810
rect 57909 20592 58351 20758
rect 57909 20540 57998 20592
rect 58050 20540 58210 20592
rect 58262 20540 58351 20592
rect 57909 20374 58351 20540
rect 57909 20322 57998 20374
rect 58050 20322 58210 20374
rect 58262 20322 58351 20374
rect 57909 20157 58351 20322
rect 57909 20105 57998 20157
rect 58050 20105 58210 20157
rect 58262 20105 58351 20157
rect 57909 19939 58351 20105
rect 57909 19887 57998 19939
rect 58050 19887 58210 19939
rect 58262 19887 58351 19939
rect 57909 19722 58351 19887
rect 57909 19670 57998 19722
rect 58050 19670 58210 19722
rect 58262 19670 58351 19722
rect 57909 19504 58351 19670
rect 57909 19452 57998 19504
rect 58050 19452 58210 19504
rect 58262 19452 58351 19504
rect 57909 19286 58351 19452
rect 57909 19234 57998 19286
rect 58050 19234 58210 19286
rect 58262 19234 58351 19286
rect 57909 19068 58351 19234
rect 57909 19016 57998 19068
rect 58050 19016 58210 19068
rect 58262 19016 58351 19068
rect 57909 18851 58351 19016
rect 57909 18799 57998 18851
rect 58050 18799 58210 18851
rect 58262 18799 58351 18851
rect 57909 18633 58351 18799
rect 57909 18581 57998 18633
rect 58050 18581 58210 18633
rect 58262 18581 58351 18633
rect 57909 18416 58351 18581
rect 57909 18364 57998 18416
rect 58050 18364 58210 18416
rect 58262 18364 58351 18416
rect 57909 18198 58351 18364
rect 57909 18146 57998 18198
rect 58050 18146 58210 18198
rect 58262 18146 58351 18198
rect 57909 17980 58351 18146
rect 57909 17928 57998 17980
rect 58050 17928 58210 17980
rect 58262 17928 58351 17980
rect 57909 17763 58351 17928
rect 57909 17711 57998 17763
rect 58050 17711 58210 17763
rect 58262 17711 58351 17763
rect 57909 17545 58351 17711
rect 57909 17493 57998 17545
rect 58050 17493 58210 17545
rect 58262 17493 58351 17545
rect 57909 17327 58351 17493
rect 57909 17275 57998 17327
rect 58050 17275 58210 17327
rect 58262 17275 58351 17327
rect 57909 17110 58351 17275
rect 57909 17058 57998 17110
rect 58050 17058 58210 17110
rect 58262 17058 58351 17110
rect 57909 16892 58351 17058
rect 57909 16840 57998 16892
rect 58050 16840 58210 16892
rect 58262 16840 58351 16892
rect 57909 16675 58351 16840
rect 57909 16623 57998 16675
rect 58050 16623 58210 16675
rect 58262 16623 58351 16675
rect 57909 16457 58351 16623
rect 57909 16405 57998 16457
rect 58050 16405 58210 16457
rect 58262 16405 58351 16457
rect 57909 16239 58351 16405
rect 57909 16187 57998 16239
rect 58050 16187 58210 16239
rect 58262 16187 58351 16239
rect 57909 16022 58351 16187
rect 57909 15970 57998 16022
rect 58050 15970 58210 16022
rect 58262 15970 58351 16022
rect 57909 15804 58351 15970
rect 57909 15752 57998 15804
rect 58050 15752 58210 15804
rect 58262 15752 58351 15804
rect 57909 15586 58351 15752
rect 57909 15534 57998 15586
rect 58050 15534 58210 15586
rect 58262 15534 58351 15586
rect 57909 15369 58351 15534
rect 57909 15317 57998 15369
rect 58050 15317 58210 15369
rect 58262 15317 58351 15369
rect 57909 15151 58351 15317
rect 57909 15099 57998 15151
rect 58050 15099 58210 15151
rect 58262 15099 58351 15151
rect 57909 14933 58351 15099
rect 57909 14881 57998 14933
rect 58050 14881 58210 14933
rect 58262 14881 58351 14933
rect 57909 14716 58351 14881
rect 57909 14664 57998 14716
rect 58050 14664 58210 14716
rect 58262 14664 58351 14716
rect 57909 14498 58351 14664
rect 57909 14446 57998 14498
rect 58050 14446 58210 14498
rect 58262 14446 58351 14498
rect 57909 14281 58351 14446
rect 57909 14229 57998 14281
rect 58050 14229 58210 14281
rect 58262 14229 58351 14281
rect 57909 14063 58351 14229
rect 57909 14011 57998 14063
rect 58050 14011 58210 14063
rect 58262 14011 58351 14063
rect 57909 13845 58351 14011
rect 57909 13793 57998 13845
rect 58050 13793 58210 13845
rect 58262 13793 58351 13845
rect 57909 13628 58351 13793
rect 57909 13576 57998 13628
rect 58050 13576 58210 13628
rect 58262 13576 58351 13628
rect 57909 13410 58351 13576
rect 57909 13358 57998 13410
rect 58050 13358 58210 13410
rect 58262 13358 58351 13410
rect 57909 13192 58351 13358
rect 57909 13140 57998 13192
rect 58050 13140 58210 13192
rect 58262 13140 58351 13192
rect 57909 12975 58351 13140
rect 57909 12923 57998 12975
rect 58050 12923 58210 12975
rect 58262 12923 58351 12975
rect 57909 12757 58351 12923
rect 57909 12705 57998 12757
rect 58050 12705 58210 12757
rect 58262 12705 58351 12757
rect 57909 12540 58351 12705
rect 57909 12488 57998 12540
rect 58050 12488 58210 12540
rect 58262 12488 58351 12540
rect 57909 12322 58351 12488
rect 57909 12270 57998 12322
rect 58050 12270 58210 12322
rect 58262 12270 58351 12322
rect 57909 12104 58351 12270
rect 57909 12052 57998 12104
rect 58050 12052 58210 12104
rect 58262 12052 58351 12104
rect 57909 11887 58351 12052
rect 57909 11835 57998 11887
rect 58050 11835 58210 11887
rect 58262 11835 58351 11887
rect 57909 11669 58351 11835
rect 57909 11617 57998 11669
rect 58050 11617 58210 11669
rect 58262 11617 58351 11669
rect 57909 11451 58351 11617
rect 57909 11399 57998 11451
rect 58050 11399 58210 11451
rect 58262 11399 58351 11451
rect 57909 11234 58351 11399
rect 57909 11182 57998 11234
rect 58050 11182 58210 11234
rect 58262 11182 58351 11234
rect 57909 11016 58351 11182
rect 57909 10964 57998 11016
rect 58050 10964 58210 11016
rect 58262 10964 58351 11016
rect 57909 10798 58351 10964
rect 57909 10746 57998 10798
rect 58050 10746 58210 10798
rect 58262 10746 58351 10798
rect 57909 10581 58351 10746
rect 57909 10529 57998 10581
rect 58050 10529 58210 10581
rect 58262 10529 58351 10581
rect 57909 10363 58351 10529
rect 57909 10311 57998 10363
rect 58050 10311 58210 10363
rect 58262 10311 58351 10363
rect 57909 10146 58351 10311
rect 57909 10094 57998 10146
rect 58050 10094 58210 10146
rect 58262 10094 58351 10146
rect 57909 9928 58351 10094
rect 57909 9876 57998 9928
rect 58050 9876 58210 9928
rect 58262 9876 58351 9928
rect 57909 9710 58351 9876
rect 57909 9658 57998 9710
rect 58050 9658 58210 9710
rect 58262 9658 58351 9710
rect 57909 9493 58351 9658
rect 57909 9441 57998 9493
rect 58050 9441 58210 9493
rect 58262 9441 58351 9493
rect 57909 9275 58351 9441
rect 57909 9223 57998 9275
rect 58050 9223 58210 9275
rect 58262 9223 58351 9275
rect 57909 9057 58351 9223
rect 57909 9005 57998 9057
rect 58050 9005 58210 9057
rect 58262 9005 58351 9057
rect 57909 8840 58351 9005
rect 57909 8788 57998 8840
rect 58050 8788 58210 8840
rect 58262 8788 58351 8840
rect 57909 8622 58351 8788
rect 57909 8570 57998 8622
rect 58050 8570 58210 8622
rect 58262 8570 58351 8622
rect 57909 8404 58351 8570
rect 57909 8352 57998 8404
rect 58050 8352 58210 8404
rect 58262 8352 58351 8404
rect 57909 8187 58351 8352
rect 57909 8135 57998 8187
rect 58050 8135 58210 8187
rect 58262 8135 58351 8187
rect 57909 7969 58351 8135
rect 57909 7917 57998 7969
rect 58050 7917 58210 7969
rect 58262 7917 58351 7969
rect 57909 7752 58351 7917
rect 57909 7700 57998 7752
rect 58050 7700 58210 7752
rect 58262 7700 58351 7752
rect 57909 7534 58351 7700
rect 57909 7482 57998 7534
rect 58050 7482 58210 7534
rect 58262 7482 58351 7534
rect 57909 7316 58351 7482
rect 57909 7264 57998 7316
rect 58050 7264 58210 7316
rect 58262 7264 58351 7316
rect 57909 7099 58351 7264
rect 57909 7047 57998 7099
rect 58050 7047 58210 7099
rect 58262 7047 58351 7099
rect 57909 6881 58351 7047
rect 57909 6829 57998 6881
rect 58050 6829 58210 6881
rect 58262 6829 58351 6881
rect 57909 6663 58351 6829
rect 57909 6611 57998 6663
rect 58050 6611 58210 6663
rect 58262 6611 58351 6663
rect 57909 6446 58351 6611
rect 57909 6394 57998 6446
rect 58050 6394 58210 6446
rect 58262 6394 58351 6446
rect 57909 6228 58351 6394
rect 57909 6176 57998 6228
rect 58050 6176 58210 6228
rect 58262 6176 58351 6228
rect 57909 6011 58351 6176
rect 57909 5959 57998 6011
rect 58050 5959 58210 6011
rect 58262 5959 58351 6011
rect 57909 5793 58351 5959
rect 57909 5741 57998 5793
rect 58050 5741 58210 5793
rect 58262 5741 58351 5793
rect 57909 5575 58351 5741
rect 57909 5523 57998 5575
rect 58050 5523 58210 5575
rect 58262 5523 58351 5575
rect 57909 5358 58351 5523
rect 57909 5306 57998 5358
rect 58050 5306 58210 5358
rect 58262 5306 58351 5358
rect 57909 5220 58351 5306
rect 57626 4728 57637 5220
rect 57626 4587 57736 4728
rect 57647 4535 57736 4587
rect 57626 4370 57736 4535
rect 57647 4318 57736 4370
rect 57626 4152 57736 4318
rect 57647 4100 57736 4152
rect 57626 3934 57736 4100
rect 57647 3882 57736 3934
rect 57626 3717 57736 3882
rect 57647 3665 57736 3717
rect 27744 1224 57380 1282
rect 27744 1172 48668 1224
rect 48720 1172 48792 1224
rect 48844 1172 48916 1224
rect 48968 1172 57380 1224
rect 27744 1117 57380 1172
rect 57626 3584 57736 3665
rect 57909 4587 58351 4728
rect 57909 4535 57998 4587
rect 58050 4535 58210 4587
rect 58262 4535 58351 4587
rect 57909 4370 58351 4535
rect 57909 4318 57998 4370
rect 58050 4318 58210 4370
rect 58262 4318 58351 4370
rect 57909 4152 58351 4318
rect 57909 4100 57998 4152
rect 58050 4100 58210 4152
rect 58262 4100 58351 4152
rect 57909 3934 58351 4100
rect 57909 3882 57998 3934
rect 58050 3882 58210 3934
rect 58262 3882 58351 3934
rect 57909 3717 58351 3882
rect 57909 3665 57998 3717
rect 58050 3665 58210 3717
rect 58262 3665 58351 3717
rect 57626 1282 57737 3584
rect 57909 1777 58351 3665
rect 62138 1689 62318 1701
rect 62138 1637 62150 1689
rect 62306 1637 62318 1689
rect 62138 1625 62318 1637
rect 72203 1689 72383 1701
rect 72203 1637 72215 1689
rect 72371 1637 72383 1689
rect 72203 1625 72383 1637
rect 72653 1689 72833 1701
rect 72653 1637 72665 1689
rect 72821 1637 72833 1689
rect 72653 1625 72833 1637
rect 82718 1689 82898 1701
rect 82718 1637 82730 1689
rect 82886 1637 82898 1689
rect 82718 1625 82898 1637
rect 57626 1117 86090 1282
rect 282 1100 86090 1117
rect 282 1048 48668 1100
rect 48720 1048 48792 1100
rect 48844 1048 48916 1100
rect 48968 1048 86090 1100
rect 282 976 86090 1048
rect 282 924 48668 976
rect 48720 924 48792 976
rect 48844 924 48916 976
rect 48968 924 86090 976
rect 282 915 86090 924
rect 282 655 29090 915
rect 29142 655 29792 915
rect 29844 852 86090 915
rect 29844 800 48668 852
rect 48720 800 48792 852
rect 48844 800 48916 852
rect 48968 800 86090 852
rect 29844 728 86090 800
rect 29844 676 48668 728
rect 48720 676 48792 728
rect 48844 676 48916 728
rect 48968 676 86090 728
rect 29844 655 86090 676
rect 282 604 86090 655
rect 282 552 48668 604
rect 48720 552 48792 604
rect 48844 552 48916 604
rect 48968 552 86090 604
rect 282 480 86090 552
rect 282 428 48668 480
rect 48720 428 48792 480
rect 48844 428 48916 480
rect 48968 428 86090 480
rect 282 356 86090 428
rect 282 304 48668 356
rect 48720 304 48792 356
rect 48844 304 48916 356
rect 48968 304 86090 356
rect 282 282 86090 304
<< via1 >>
rect 25400 51527 25452 51579
rect 25524 51527 25576 51579
rect 25648 51527 25700 51579
rect 25772 51527 25824 51579
rect 25896 51527 25948 51579
rect 25400 51403 25452 51455
rect 25524 51403 25576 51455
rect 25648 51403 25700 51455
rect 25772 51403 25824 51455
rect 25896 51403 25948 51455
rect 25400 51279 25452 51331
rect 25524 51279 25576 51331
rect 25648 51279 25700 51331
rect 25772 51279 25824 51331
rect 25896 51279 25948 51331
rect 27790 51401 27842 51453
rect 28001 51401 28053 51453
rect 28212 51401 28264 51453
rect 28423 51401 28475 51453
rect 28634 51401 28686 51453
rect 28845 51401 28897 51453
rect 29056 51401 29108 51453
rect 56015 51401 56067 51453
rect 56226 51401 56278 51453
rect 56437 51401 56489 51453
rect 56648 51401 56700 51453
rect 56859 51401 56911 51453
rect 57070 51401 57122 51453
rect 57281 51401 57333 51453
rect 27790 49601 27842 49653
rect 28001 49601 28053 49653
rect 28212 49601 28264 49653
rect 28423 49601 28475 49653
rect 28634 49601 28686 49653
rect 28845 49601 28897 49653
rect 29056 49601 29108 49653
rect 56015 49601 56067 49653
rect 56226 49601 56278 49653
rect 56437 49601 56489 49653
rect 56648 49601 56700 49653
rect 56859 49601 56911 49653
rect 57070 49601 57122 49653
rect 57281 49601 57333 49653
rect 27790 47801 27842 47853
rect 28001 47801 28053 47853
rect 28212 47801 28264 47853
rect 28423 47801 28475 47853
rect 28634 47801 28686 47853
rect 28845 47801 28897 47853
rect 29056 47801 29108 47853
rect 56015 47801 56067 47853
rect 56226 47801 56278 47853
rect 56437 47801 56489 47853
rect 56648 47801 56700 47853
rect 56859 47801 56911 47853
rect 57070 47801 57122 47853
rect 57281 47801 57333 47853
rect 27790 46001 27842 46053
rect 28001 46001 28053 46053
rect 28212 46001 28264 46053
rect 28423 46001 28475 46053
rect 28634 46001 28686 46053
rect 28845 46001 28897 46053
rect 29056 46001 29108 46053
rect 56015 46001 56067 46053
rect 56226 46001 56278 46053
rect 56437 46001 56489 46053
rect 56648 46001 56700 46053
rect 56859 46001 56911 46053
rect 57070 46001 57122 46053
rect 57281 46001 57333 46053
rect 27790 44201 27842 44253
rect 28001 44201 28053 44253
rect 28212 44201 28264 44253
rect 28423 44201 28475 44253
rect 28634 44201 28686 44253
rect 28845 44201 28897 44253
rect 29056 44201 29108 44253
rect 56015 44201 56067 44253
rect 56226 44201 56278 44253
rect 56437 44201 56489 44253
rect 56648 44201 56700 44253
rect 56859 44201 56911 44253
rect 57070 44201 57122 44253
rect 57281 44201 57333 44253
rect 27790 42401 27842 42453
rect 28001 42401 28053 42453
rect 28212 42401 28264 42453
rect 28423 42401 28475 42453
rect 28634 42401 28686 42453
rect 28845 42401 28897 42453
rect 29056 42401 29108 42453
rect 56015 42401 56067 42453
rect 56226 42401 56278 42453
rect 56437 42401 56489 42453
rect 56648 42401 56700 42453
rect 56859 42401 56911 42453
rect 57070 42401 57122 42453
rect 57281 42401 57333 42453
rect 27790 40601 27842 40653
rect 28001 40601 28053 40653
rect 28212 40601 28264 40653
rect 28423 40601 28475 40653
rect 28634 40601 28686 40653
rect 28845 40601 28897 40653
rect 29056 40601 29108 40653
rect 56015 40601 56067 40653
rect 56226 40601 56278 40653
rect 56437 40601 56489 40653
rect 56648 40601 56700 40653
rect 56859 40601 56911 40653
rect 57070 40601 57122 40653
rect 57281 40601 57333 40653
rect 27790 38801 27842 38853
rect 28001 38801 28053 38853
rect 28212 38801 28264 38853
rect 28423 38801 28475 38853
rect 28634 38801 28686 38853
rect 28845 38801 28897 38853
rect 29056 38801 29108 38853
rect 56015 38801 56067 38853
rect 56226 38801 56278 38853
rect 56437 38801 56489 38853
rect 56648 38801 56700 38853
rect 56859 38801 56911 38853
rect 57070 38801 57122 38853
rect 57281 38801 57333 38853
rect 27790 37001 27842 37053
rect 28001 37001 28053 37053
rect 28212 37001 28264 37053
rect 28423 37001 28475 37053
rect 28634 37001 28686 37053
rect 28845 37001 28897 37053
rect 29056 37001 29108 37053
rect 56015 37001 56067 37053
rect 56226 37001 56278 37053
rect 56437 37001 56489 37053
rect 56648 37001 56700 37053
rect 56859 37001 56911 37053
rect 57070 37001 57122 37053
rect 57281 37001 57333 37053
rect 27440 35221 27492 35273
rect 27564 35221 27616 35273
rect 27688 35221 27740 35273
rect 27440 35097 27492 35149
rect 27564 35097 27616 35149
rect 27688 35097 27740 35149
rect 27440 34973 27492 35025
rect 27564 34973 27616 35025
rect 27688 34973 27740 35025
rect 27440 34849 27492 34901
rect 27564 34849 27616 34901
rect 27688 34849 27740 34901
rect 27440 34725 27492 34777
rect 27564 34725 27616 34777
rect 27688 34725 27740 34777
rect 27440 34601 27492 34653
rect 27564 34601 27616 34653
rect 27688 34601 27740 34653
rect 26861 33380 26913 33432
rect 27073 33380 27125 33432
rect 26861 33163 26913 33215
rect 27073 33163 27125 33215
rect 26861 32945 26913 32997
rect 27073 32945 27125 32997
rect 26861 32727 26913 32779
rect 27073 32727 27125 32779
rect 26861 32510 26913 32562
rect 27073 32510 27125 32562
rect 26861 32292 26913 32344
rect 27073 32292 27125 32344
rect 26861 32075 26913 32127
rect 27073 32075 27125 32127
rect 26861 31857 26913 31909
rect 27073 31857 27125 31909
rect 26861 31639 26913 31691
rect 27073 31639 27125 31691
rect 26861 31422 26913 31474
rect 27073 31422 27125 31474
rect 26861 31204 26913 31256
rect 27073 31204 27125 31256
rect 26861 30986 26913 31038
rect 27073 30986 27125 31038
rect 26861 30769 26913 30821
rect 27073 30769 27125 30821
rect 26861 30551 26913 30603
rect 27073 30551 27125 30603
rect 26861 30334 26913 30386
rect 27073 30334 27125 30386
rect 26861 30116 26913 30168
rect 27073 30116 27125 30168
rect 26861 29898 26913 29950
rect 27073 29898 27125 29950
rect 26861 29681 26913 29733
rect 27073 29681 27125 29733
rect 26861 29463 26913 29515
rect 27073 29463 27125 29515
rect 26861 29245 26913 29297
rect 27073 29245 27125 29297
rect 26861 29028 26913 29080
rect 27073 29028 27125 29080
rect 26861 28810 26913 28862
rect 27073 28810 27125 28862
rect 26861 28592 26913 28644
rect 27073 28592 27125 28644
rect 26861 28375 26913 28427
rect 27073 28375 27125 28427
rect 26861 28157 26913 28209
rect 27073 28157 27125 28209
rect 26861 27940 26913 27992
rect 27073 27940 27125 27992
rect 26861 27722 26913 27774
rect 27073 27722 27125 27774
rect 26861 27504 26913 27556
rect 27073 27504 27125 27556
rect 26861 27287 26913 27339
rect 27073 27287 27125 27339
rect 26861 27069 26913 27121
rect 27073 27069 27125 27121
rect 26861 26851 26913 26903
rect 27073 26851 27125 26903
rect 26861 26634 26913 26686
rect 27073 26634 27125 26686
rect 26861 26416 26913 26468
rect 27073 26416 27125 26468
rect 26861 26198 26913 26250
rect 27073 26198 27125 26250
rect 26861 25981 26913 26033
rect 27073 25981 27125 26033
rect 26861 25763 26913 25815
rect 27073 25763 27125 25815
rect 26861 25546 26913 25598
rect 27073 25546 27125 25598
rect 26861 25328 26913 25380
rect 27073 25328 27125 25380
rect 26861 25110 26913 25162
rect 27073 25110 27125 25162
rect 26861 24893 26913 24945
rect 27073 24893 27125 24945
rect 26861 24675 26913 24727
rect 27073 24675 27125 24727
rect 26861 24457 26913 24509
rect 27073 24457 27125 24509
rect 26861 24240 26913 24292
rect 27073 24240 27125 24292
rect 26861 24022 26913 24074
rect 27073 24022 27125 24074
rect 26861 23805 26913 23857
rect 27073 23805 27125 23857
rect 26861 23587 26913 23639
rect 27073 23587 27125 23639
rect 26861 23369 26913 23421
rect 27073 23369 27125 23421
rect 26861 23152 26913 23204
rect 27073 23152 27125 23204
rect 26861 22934 26913 22986
rect 27073 22934 27125 22986
rect 26861 22716 26913 22768
rect 27073 22716 27125 22768
rect 26861 22499 26913 22551
rect 27073 22499 27125 22551
rect 26861 22281 26913 22333
rect 27073 22281 27125 22333
rect 26861 22063 26913 22115
rect 27073 22063 27125 22115
rect 26861 21846 26913 21898
rect 27073 21846 27125 21898
rect 26861 21628 26913 21680
rect 27073 21628 27125 21680
rect 26861 21411 26913 21463
rect 27073 21411 27125 21463
rect 26861 21193 26913 21245
rect 27073 21193 27125 21245
rect 26861 20975 26913 21027
rect 27073 20975 27125 21027
rect 26861 20758 26913 20810
rect 27073 20758 27125 20810
rect 26861 20540 26913 20592
rect 27073 20540 27125 20592
rect 26861 20322 26913 20374
rect 27073 20322 27125 20374
rect 26861 20105 26913 20157
rect 27073 20105 27125 20157
rect 26861 19887 26913 19939
rect 27073 19887 27125 19939
rect 26861 19670 26913 19722
rect 27073 19670 27125 19722
rect 26861 19452 26913 19504
rect 27073 19452 27125 19504
rect 26861 19234 26913 19286
rect 27073 19234 27125 19286
rect 26861 19016 26913 19068
rect 27073 19016 27125 19068
rect 26861 18799 26913 18851
rect 27073 18799 27125 18851
rect 26861 18581 26913 18633
rect 27073 18581 27125 18633
rect 26861 18364 26913 18416
rect 27073 18364 27125 18416
rect 26861 18146 26913 18198
rect 27073 18146 27125 18198
rect 26861 17928 26913 17980
rect 27073 17928 27125 17980
rect 26861 17711 26913 17763
rect 27073 17711 27125 17763
rect 26861 17493 26913 17545
rect 27073 17493 27125 17545
rect 26861 17275 26913 17327
rect 27073 17275 27125 17327
rect 26861 17058 26913 17110
rect 27073 17058 27125 17110
rect 26861 16840 26913 16892
rect 27073 16840 27125 16892
rect 26861 16623 26913 16675
rect 27073 16623 27125 16675
rect 26861 16405 26913 16457
rect 27073 16405 27125 16457
rect 26861 16187 26913 16239
rect 27073 16187 27125 16239
rect 26861 15970 26913 16022
rect 27073 15970 27125 16022
rect 26861 15752 26913 15804
rect 27073 15752 27125 15804
rect 26861 15534 26913 15586
rect 27073 15534 27125 15586
rect 26861 15317 26913 15369
rect 27073 15317 27125 15369
rect 26861 15099 26913 15151
rect 27073 15099 27125 15151
rect 26861 14881 26913 14933
rect 27073 14881 27125 14933
rect 26861 14664 26913 14716
rect 27073 14664 27125 14716
rect 26861 14446 26913 14498
rect 27073 14446 27125 14498
rect 26861 14229 26913 14281
rect 27073 14229 27125 14281
rect 26861 14011 26913 14063
rect 27073 14011 27125 14063
rect 26861 13793 26913 13845
rect 27073 13793 27125 13845
rect 26861 13576 26913 13628
rect 27073 13576 27125 13628
rect 26861 13358 26913 13410
rect 27073 13358 27125 13410
rect 26861 13140 26913 13192
rect 27073 13140 27125 13192
rect 26861 12923 26913 12975
rect 27073 12923 27125 12975
rect 26861 12705 26913 12757
rect 27073 12705 27125 12757
rect 26861 12488 26913 12540
rect 27073 12488 27125 12540
rect 26861 12270 26913 12322
rect 27073 12270 27125 12322
rect 26861 12052 26913 12104
rect 27073 12052 27125 12104
rect 26861 11835 26913 11887
rect 27073 11835 27125 11887
rect 26861 11617 26913 11669
rect 27073 11617 27125 11669
rect 26861 11399 26913 11451
rect 27073 11399 27125 11451
rect 26861 11182 26913 11234
rect 27073 11182 27125 11234
rect 26861 10964 26913 11016
rect 27073 10964 27125 11016
rect 26861 10746 26913 10798
rect 27073 10746 27125 10798
rect 26861 10529 26913 10581
rect 27073 10529 27125 10581
rect 26861 10311 26913 10363
rect 27073 10311 27125 10363
rect 26861 10094 26913 10146
rect 27073 10094 27125 10146
rect 26861 9876 26913 9928
rect 27073 9876 27125 9928
rect 26861 9658 26913 9710
rect 27073 9658 27125 9710
rect 26861 9441 26913 9493
rect 27073 9441 27125 9493
rect 26861 9223 26913 9275
rect 27073 9223 27125 9275
rect 26861 9005 26913 9057
rect 27073 9005 27125 9057
rect 26861 8788 26913 8840
rect 27073 8788 27125 8840
rect 26861 8570 26913 8622
rect 27073 8570 27125 8622
rect 26861 8352 26913 8404
rect 27073 8352 27125 8404
rect 26861 8135 26913 8187
rect 27073 8135 27125 8187
rect 26861 7917 26913 7969
rect 27073 7917 27125 7969
rect 26861 7700 26913 7752
rect 27073 7700 27125 7752
rect 26861 7482 26913 7534
rect 27073 7482 27125 7534
rect 26861 7264 26913 7316
rect 27073 7264 27125 7316
rect 26861 7047 26913 7099
rect 27073 7047 27125 7099
rect 26861 6829 26913 6881
rect 27073 6829 27125 6881
rect 26861 6611 26913 6663
rect 27073 6611 27125 6663
rect 26861 6394 26913 6446
rect 27073 6394 27125 6446
rect 26861 6176 26913 6228
rect 27073 6176 27125 6228
rect 26861 5959 26913 6011
rect 27073 5959 27125 6011
rect 26861 5741 26913 5793
rect 27073 5741 27125 5793
rect 26861 5523 26913 5575
rect 27073 5523 27125 5575
rect 26861 5306 26913 5358
rect 27073 5306 27125 5358
rect 26861 4535 26913 4587
rect 27073 4535 27125 4587
rect 26861 4318 26913 4370
rect 27073 4318 27125 4370
rect 26861 4100 26913 4152
rect 27073 4100 27125 4152
rect 26861 3882 26913 3934
rect 27073 3882 27125 3934
rect 26861 3665 26913 3717
rect 27073 3665 27125 3717
rect 27476 33380 27498 33432
rect 27498 33380 27528 33432
rect 27688 33380 27740 33432
rect 27476 33163 27498 33215
rect 27498 33163 27528 33215
rect 27688 33163 27740 33215
rect 27476 32945 27498 32997
rect 27498 32945 27528 32997
rect 27688 32945 27740 32997
rect 27476 32727 27498 32779
rect 27498 32727 27528 32779
rect 27688 32727 27740 32779
rect 27476 32510 27498 32562
rect 27498 32510 27528 32562
rect 27688 32510 27740 32562
rect 27476 32292 27498 32344
rect 27498 32292 27528 32344
rect 27688 32292 27740 32344
rect 27476 32075 27498 32127
rect 27498 32075 27528 32127
rect 27688 32075 27740 32127
rect 27476 31857 27498 31909
rect 27498 31857 27528 31909
rect 27688 31857 27740 31909
rect 27476 31639 27498 31691
rect 27498 31639 27528 31691
rect 27688 31639 27740 31691
rect 27476 31422 27498 31474
rect 27498 31422 27528 31474
rect 27688 31422 27740 31474
rect 27476 31204 27498 31256
rect 27498 31204 27528 31256
rect 27688 31204 27740 31256
rect 27476 30986 27498 31038
rect 27498 30986 27528 31038
rect 27688 30986 27740 31038
rect 27476 30769 27498 30821
rect 27498 30769 27528 30821
rect 27688 30769 27740 30821
rect 27476 30551 27498 30603
rect 27498 30551 27528 30603
rect 27688 30551 27740 30603
rect 27476 30334 27498 30386
rect 27498 30334 27528 30386
rect 27688 30334 27740 30386
rect 27476 30116 27498 30168
rect 27498 30116 27528 30168
rect 27688 30116 27740 30168
rect 27476 29898 27498 29950
rect 27498 29898 27528 29950
rect 27688 29898 27740 29950
rect 27476 29681 27498 29733
rect 27498 29681 27528 29733
rect 27688 29681 27740 29733
rect 27476 29463 27498 29515
rect 27498 29463 27528 29515
rect 27688 29463 27740 29515
rect 27476 29245 27498 29297
rect 27498 29245 27528 29297
rect 27688 29245 27740 29297
rect 27476 29028 27498 29080
rect 27498 29028 27528 29080
rect 27688 29028 27740 29080
rect 27476 28810 27498 28862
rect 27498 28810 27528 28862
rect 27688 28810 27740 28862
rect 27476 28592 27498 28644
rect 27498 28592 27528 28644
rect 27688 28592 27740 28644
rect 27476 28375 27498 28427
rect 27498 28375 27528 28427
rect 27688 28375 27740 28427
rect 27476 28157 27498 28209
rect 27498 28157 27528 28209
rect 27688 28157 27740 28209
rect 27476 27940 27498 27992
rect 27498 27940 27528 27992
rect 27688 27940 27740 27992
rect 27476 27722 27498 27774
rect 27498 27722 27528 27774
rect 27688 27722 27740 27774
rect 27476 27504 27498 27556
rect 27498 27504 27528 27556
rect 27688 27504 27740 27556
rect 27476 27287 27498 27339
rect 27498 27287 27528 27339
rect 27688 27287 27740 27339
rect 27476 27069 27498 27121
rect 27498 27069 27528 27121
rect 27688 27069 27740 27121
rect 27476 26851 27498 26903
rect 27498 26851 27528 26903
rect 27688 26851 27740 26903
rect 27476 26634 27498 26686
rect 27498 26634 27528 26686
rect 27688 26634 27740 26686
rect 27476 26416 27498 26468
rect 27498 26416 27528 26468
rect 27688 26416 27740 26468
rect 27476 26198 27498 26250
rect 27498 26198 27528 26250
rect 27688 26198 27740 26250
rect 27476 25981 27498 26033
rect 27498 25981 27528 26033
rect 27688 25981 27740 26033
rect 27476 25763 27498 25815
rect 27498 25763 27528 25815
rect 27688 25763 27740 25815
rect 27476 25546 27498 25598
rect 27498 25546 27528 25598
rect 27688 25546 27740 25598
rect 27476 25328 27498 25380
rect 27498 25328 27528 25380
rect 27688 25328 27740 25380
rect 27476 25110 27498 25162
rect 27498 25110 27528 25162
rect 27688 25110 27740 25162
rect 27476 24893 27498 24945
rect 27498 24893 27528 24945
rect 27688 24893 27740 24945
rect 27476 24675 27498 24727
rect 27498 24675 27528 24727
rect 27688 24675 27740 24727
rect 27476 24457 27498 24509
rect 27498 24457 27528 24509
rect 27688 24457 27740 24509
rect 27476 24240 27498 24292
rect 27498 24240 27528 24292
rect 27688 24240 27740 24292
rect 27476 24022 27498 24074
rect 27498 24022 27528 24074
rect 27688 24022 27740 24074
rect 27476 23805 27498 23857
rect 27498 23805 27528 23857
rect 27688 23805 27740 23857
rect 27476 23587 27498 23639
rect 27498 23587 27528 23639
rect 27688 23587 27740 23639
rect 27476 23369 27498 23421
rect 27498 23369 27528 23421
rect 27688 23369 27740 23421
rect 27476 23152 27498 23204
rect 27498 23152 27528 23204
rect 27688 23152 27740 23204
rect 27476 22934 27498 22986
rect 27498 22934 27528 22986
rect 27688 22934 27740 22986
rect 27476 22716 27498 22768
rect 27498 22716 27528 22768
rect 27688 22716 27740 22768
rect 27476 22499 27498 22551
rect 27498 22499 27528 22551
rect 27688 22499 27740 22551
rect 27476 22281 27498 22333
rect 27498 22281 27528 22333
rect 27688 22281 27740 22333
rect 27476 22063 27498 22115
rect 27498 22063 27528 22115
rect 27688 22063 27740 22115
rect 27476 21846 27498 21898
rect 27498 21846 27528 21898
rect 27688 21846 27740 21898
rect 27476 21628 27498 21680
rect 27498 21628 27528 21680
rect 27688 21628 27740 21680
rect 27476 21411 27498 21463
rect 27498 21411 27528 21463
rect 27688 21411 27740 21463
rect 27476 21193 27498 21245
rect 27498 21193 27528 21245
rect 27688 21193 27740 21245
rect 27476 20975 27498 21027
rect 27498 20975 27528 21027
rect 27688 20975 27740 21027
rect 27476 20758 27498 20810
rect 27498 20758 27528 20810
rect 27688 20758 27740 20810
rect 27476 20540 27498 20592
rect 27498 20540 27528 20592
rect 27688 20540 27740 20592
rect 27476 20322 27498 20374
rect 27498 20322 27528 20374
rect 27688 20322 27740 20374
rect 27476 20105 27498 20157
rect 27498 20105 27528 20157
rect 27688 20105 27740 20157
rect 27476 19887 27498 19939
rect 27498 19887 27528 19939
rect 27688 19887 27740 19939
rect 27476 19670 27498 19722
rect 27498 19670 27528 19722
rect 27688 19670 27740 19722
rect 27476 19452 27498 19504
rect 27498 19452 27528 19504
rect 27688 19452 27740 19504
rect 27476 19234 27498 19286
rect 27498 19234 27528 19286
rect 27688 19234 27740 19286
rect 27476 19016 27498 19068
rect 27498 19016 27528 19068
rect 27688 19016 27740 19068
rect 27476 18799 27498 18851
rect 27498 18799 27528 18851
rect 27688 18799 27740 18851
rect 27476 18581 27498 18633
rect 27498 18581 27528 18633
rect 27688 18581 27740 18633
rect 27476 18364 27498 18416
rect 27498 18364 27528 18416
rect 27688 18364 27740 18416
rect 27476 18146 27498 18198
rect 27498 18146 27528 18198
rect 27688 18146 27740 18198
rect 27476 17928 27498 17980
rect 27498 17928 27528 17980
rect 27688 17928 27740 17980
rect 27476 17711 27498 17763
rect 27498 17711 27528 17763
rect 27688 17711 27740 17763
rect 27476 17493 27498 17545
rect 27498 17493 27528 17545
rect 27688 17493 27740 17545
rect 27476 17275 27498 17327
rect 27498 17275 27528 17327
rect 27688 17275 27740 17327
rect 27476 17058 27498 17110
rect 27498 17058 27528 17110
rect 27688 17058 27740 17110
rect 27476 16840 27498 16892
rect 27498 16840 27528 16892
rect 27688 16840 27740 16892
rect 27476 16623 27498 16675
rect 27498 16623 27528 16675
rect 27688 16623 27740 16675
rect 27476 16405 27498 16457
rect 27498 16405 27528 16457
rect 27688 16405 27740 16457
rect 27476 16187 27498 16239
rect 27498 16187 27528 16239
rect 27688 16187 27740 16239
rect 27476 15970 27498 16022
rect 27498 15970 27528 16022
rect 27688 15970 27740 16022
rect 27476 15752 27498 15804
rect 27498 15752 27528 15804
rect 27688 15752 27740 15804
rect 27476 15534 27498 15586
rect 27498 15534 27528 15586
rect 27688 15534 27740 15586
rect 27476 15317 27498 15369
rect 27498 15317 27528 15369
rect 27688 15317 27740 15369
rect 27476 15099 27498 15151
rect 27498 15099 27528 15151
rect 27688 15099 27740 15151
rect 27476 14881 27498 14933
rect 27498 14881 27528 14933
rect 27688 14881 27740 14933
rect 27476 14664 27498 14716
rect 27498 14664 27528 14716
rect 27688 14664 27740 14716
rect 27476 14446 27498 14498
rect 27498 14446 27528 14498
rect 27688 14446 27740 14498
rect 27476 14229 27498 14281
rect 27498 14229 27528 14281
rect 27688 14229 27740 14281
rect 27476 14011 27498 14063
rect 27498 14011 27528 14063
rect 27688 14011 27740 14063
rect 27476 13793 27498 13845
rect 27498 13793 27528 13845
rect 27688 13793 27740 13845
rect 27476 13576 27498 13628
rect 27498 13576 27528 13628
rect 27688 13576 27740 13628
rect 27476 13358 27498 13410
rect 27498 13358 27528 13410
rect 27688 13358 27740 13410
rect 27476 13140 27498 13192
rect 27498 13140 27528 13192
rect 27688 13140 27740 13192
rect 27476 12923 27498 12975
rect 27498 12923 27528 12975
rect 27688 12923 27740 12975
rect 27476 12705 27498 12757
rect 27498 12705 27528 12757
rect 27688 12705 27740 12757
rect 27476 12488 27498 12540
rect 27498 12488 27528 12540
rect 27688 12488 27740 12540
rect 27476 12270 27498 12322
rect 27498 12270 27528 12322
rect 27688 12270 27740 12322
rect 27476 12052 27498 12104
rect 27498 12052 27528 12104
rect 27688 12052 27740 12104
rect 27476 11835 27498 11887
rect 27498 11835 27528 11887
rect 27688 11835 27740 11887
rect 27476 11617 27498 11669
rect 27498 11617 27528 11669
rect 27688 11617 27740 11669
rect 27476 11399 27498 11451
rect 27498 11399 27528 11451
rect 27688 11399 27740 11451
rect 27476 11182 27498 11234
rect 27498 11182 27528 11234
rect 27688 11182 27740 11234
rect 27476 10964 27498 11016
rect 27498 10964 27528 11016
rect 27688 10964 27740 11016
rect 27476 10746 27498 10798
rect 27498 10746 27528 10798
rect 27688 10746 27740 10798
rect 27476 10529 27498 10581
rect 27498 10529 27528 10581
rect 27688 10529 27740 10581
rect 27476 10311 27498 10363
rect 27498 10311 27528 10363
rect 27688 10311 27740 10363
rect 27476 10094 27498 10146
rect 27498 10094 27528 10146
rect 27688 10094 27740 10146
rect 27476 9876 27498 9928
rect 27498 9876 27528 9928
rect 27688 9876 27740 9928
rect 27476 9658 27498 9710
rect 27498 9658 27528 9710
rect 27688 9658 27740 9710
rect 27476 9441 27498 9493
rect 27498 9441 27528 9493
rect 27688 9441 27740 9493
rect 27476 9223 27498 9275
rect 27498 9223 27528 9275
rect 27688 9223 27740 9275
rect 27476 9005 27498 9057
rect 27498 9005 27528 9057
rect 27688 9005 27740 9057
rect 27476 8788 27498 8840
rect 27498 8788 27528 8840
rect 27688 8788 27740 8840
rect 27476 8570 27498 8622
rect 27498 8570 27528 8622
rect 27688 8570 27740 8622
rect 27476 8352 27498 8404
rect 27498 8352 27528 8404
rect 27688 8352 27740 8404
rect 27476 8135 27498 8187
rect 27498 8135 27528 8187
rect 27688 8135 27740 8187
rect 27476 7917 27498 7969
rect 27498 7917 27528 7969
rect 27688 7917 27740 7969
rect 27476 7700 27498 7752
rect 27498 7700 27528 7752
rect 27688 7700 27740 7752
rect 27476 7482 27498 7534
rect 27498 7482 27528 7534
rect 27688 7482 27740 7534
rect 27476 7264 27498 7316
rect 27498 7264 27528 7316
rect 27688 7264 27740 7316
rect 27476 7047 27498 7099
rect 27498 7047 27528 7099
rect 27688 7047 27740 7099
rect 27476 6829 27498 6881
rect 27498 6829 27528 6881
rect 27688 6829 27740 6881
rect 27476 6611 27498 6663
rect 27498 6611 27528 6663
rect 27688 6611 27740 6663
rect 27476 6394 27498 6446
rect 27498 6394 27528 6446
rect 27688 6394 27740 6446
rect 27476 6176 27498 6228
rect 27498 6176 27528 6228
rect 27688 6176 27740 6228
rect 27476 5959 27498 6011
rect 27498 5959 27528 6011
rect 27688 5959 27740 6011
rect 27476 5741 27498 5793
rect 27498 5741 27528 5793
rect 27688 5741 27740 5793
rect 27476 5523 27498 5575
rect 27498 5523 27528 5575
rect 27688 5523 27740 5575
rect 27476 5306 27498 5358
rect 27498 5306 27528 5358
rect 27688 5306 27740 5358
rect 27476 4535 27498 4587
rect 27498 4535 27528 4587
rect 27688 4535 27740 4587
rect 27476 4318 27498 4370
rect 27498 4318 27528 4370
rect 27688 4318 27740 4370
rect 27476 4100 27498 4152
rect 27498 4100 27528 4152
rect 27688 4100 27740 4152
rect 27476 3882 27498 3934
rect 27498 3882 27528 3934
rect 27688 3882 27740 3934
rect 27476 3665 27498 3717
rect 27498 3665 27528 3717
rect 27688 3665 27740 3717
rect 2574 1637 2730 1689
rect 12639 1637 12795 1689
rect 13089 1637 13245 1689
rect 23439 1637 23595 1689
rect 57419 35190 57471 35242
rect 57543 35190 57595 35242
rect 57419 35066 57471 35118
rect 57543 35066 57595 35118
rect 57419 34942 57471 34994
rect 57543 34942 57595 34994
rect 57419 34818 57471 34870
rect 57543 34818 57595 34870
rect 57419 34694 57471 34746
rect 57543 34694 57595 34746
rect 57419 34570 57471 34622
rect 57543 34570 57595 34622
rect 49908 6297 50064 6349
rect 58878 51527 58930 51579
rect 59002 51527 59054 51579
rect 59126 51527 59178 51579
rect 59250 51527 59302 51579
rect 59374 51527 59426 51579
rect 58878 51403 58930 51455
rect 59002 51403 59054 51455
rect 59126 51403 59178 51455
rect 59250 51403 59302 51455
rect 59374 51403 59426 51455
rect 58878 51279 58930 51331
rect 59002 51279 59054 51331
rect 59126 51279 59178 51331
rect 59250 51279 59302 51331
rect 59374 51279 59426 51331
rect 60575 35338 60627 35494
rect 57383 33380 57435 33432
rect 57595 33380 57626 33432
rect 57626 33380 57647 33432
rect 57383 33163 57435 33215
rect 57595 33163 57626 33215
rect 57626 33163 57647 33215
rect 57383 32945 57435 32997
rect 57595 32945 57626 32997
rect 57626 32945 57647 32997
rect 57383 32727 57435 32779
rect 57595 32727 57626 32779
rect 57626 32727 57647 32779
rect 57383 32510 57435 32562
rect 57595 32510 57626 32562
rect 57626 32510 57647 32562
rect 57383 32292 57435 32344
rect 57595 32292 57626 32344
rect 57626 32292 57647 32344
rect 57383 32075 57435 32127
rect 57595 32075 57626 32127
rect 57626 32075 57647 32127
rect 57383 31857 57435 31909
rect 57595 31857 57626 31909
rect 57626 31857 57647 31909
rect 57383 31639 57435 31691
rect 57595 31639 57626 31691
rect 57626 31639 57647 31691
rect 57383 31422 57435 31474
rect 57595 31422 57626 31474
rect 57626 31422 57647 31474
rect 57383 31204 57435 31256
rect 57595 31204 57626 31256
rect 57626 31204 57647 31256
rect 57383 30986 57435 31038
rect 57595 30986 57626 31038
rect 57626 30986 57647 31038
rect 57383 30769 57435 30821
rect 57595 30769 57626 30821
rect 57626 30769 57647 30821
rect 57383 30551 57435 30603
rect 57595 30551 57626 30603
rect 57626 30551 57647 30603
rect 57383 30334 57435 30386
rect 57595 30334 57626 30386
rect 57626 30334 57647 30386
rect 57383 30116 57435 30168
rect 57595 30116 57626 30168
rect 57626 30116 57647 30168
rect 57383 29898 57435 29950
rect 57595 29898 57626 29950
rect 57626 29898 57647 29950
rect 57383 29681 57435 29733
rect 57595 29681 57626 29733
rect 57626 29681 57647 29733
rect 57383 29463 57435 29515
rect 57595 29463 57626 29515
rect 57626 29463 57647 29515
rect 57383 29245 57435 29297
rect 57595 29245 57626 29297
rect 57626 29245 57647 29297
rect 57383 29028 57435 29080
rect 57595 29028 57626 29080
rect 57626 29028 57647 29080
rect 57383 28810 57435 28862
rect 57595 28810 57626 28862
rect 57626 28810 57647 28862
rect 57383 28592 57435 28644
rect 57595 28592 57626 28644
rect 57626 28592 57647 28644
rect 57383 28375 57435 28427
rect 57595 28375 57626 28427
rect 57626 28375 57647 28427
rect 57383 28157 57435 28209
rect 57595 28157 57626 28209
rect 57626 28157 57647 28209
rect 57383 27940 57435 27992
rect 57595 27940 57626 27992
rect 57626 27940 57647 27992
rect 57383 27722 57435 27774
rect 57595 27722 57626 27774
rect 57626 27722 57647 27774
rect 57383 27504 57435 27556
rect 57595 27504 57626 27556
rect 57626 27504 57647 27556
rect 57383 27287 57435 27339
rect 57595 27287 57626 27339
rect 57626 27287 57647 27339
rect 57383 27069 57435 27121
rect 57595 27069 57626 27121
rect 57626 27069 57647 27121
rect 57383 26851 57435 26903
rect 57595 26851 57626 26903
rect 57626 26851 57647 26903
rect 57383 26634 57435 26686
rect 57595 26634 57626 26686
rect 57626 26634 57647 26686
rect 57383 26416 57435 26468
rect 57595 26416 57626 26468
rect 57626 26416 57647 26468
rect 57383 26198 57435 26250
rect 57595 26198 57626 26250
rect 57626 26198 57647 26250
rect 57383 25981 57435 26033
rect 57595 25981 57626 26033
rect 57626 25981 57647 26033
rect 57383 25763 57435 25815
rect 57595 25763 57626 25815
rect 57626 25763 57647 25815
rect 57383 25546 57435 25598
rect 57595 25546 57626 25598
rect 57626 25546 57647 25598
rect 57383 25328 57435 25380
rect 57595 25328 57626 25380
rect 57626 25328 57647 25380
rect 57383 25110 57435 25162
rect 57595 25110 57626 25162
rect 57626 25110 57647 25162
rect 57383 24893 57435 24945
rect 57595 24893 57626 24945
rect 57626 24893 57647 24945
rect 57383 24675 57435 24727
rect 57595 24675 57626 24727
rect 57626 24675 57647 24727
rect 57383 24457 57435 24509
rect 57595 24457 57626 24509
rect 57626 24457 57647 24509
rect 57383 24240 57435 24292
rect 57595 24240 57626 24292
rect 57626 24240 57647 24292
rect 57383 24022 57435 24074
rect 57595 24022 57626 24074
rect 57626 24022 57647 24074
rect 57383 23805 57435 23857
rect 57595 23805 57626 23857
rect 57626 23805 57647 23857
rect 57383 23587 57435 23639
rect 57595 23587 57626 23639
rect 57626 23587 57647 23639
rect 57383 23369 57435 23421
rect 57595 23369 57626 23421
rect 57626 23369 57647 23421
rect 57383 23152 57435 23204
rect 57595 23152 57626 23204
rect 57626 23152 57647 23204
rect 57383 22934 57435 22986
rect 57595 22934 57626 22986
rect 57626 22934 57647 22986
rect 57383 22716 57435 22768
rect 57595 22716 57626 22768
rect 57626 22716 57647 22768
rect 57383 22499 57435 22551
rect 57595 22499 57626 22551
rect 57626 22499 57647 22551
rect 57383 22281 57435 22333
rect 57595 22281 57626 22333
rect 57626 22281 57647 22333
rect 57383 22063 57435 22115
rect 57595 22063 57626 22115
rect 57626 22063 57647 22115
rect 57383 21846 57435 21898
rect 57595 21846 57626 21898
rect 57626 21846 57647 21898
rect 57383 21628 57435 21680
rect 57595 21628 57626 21680
rect 57626 21628 57647 21680
rect 57383 21411 57435 21463
rect 57595 21411 57626 21463
rect 57626 21411 57647 21463
rect 57383 21193 57435 21245
rect 57595 21193 57626 21245
rect 57626 21193 57647 21245
rect 57383 20975 57435 21027
rect 57595 20975 57626 21027
rect 57626 20975 57647 21027
rect 57383 20758 57435 20810
rect 57595 20758 57626 20810
rect 57626 20758 57647 20810
rect 57383 20540 57435 20592
rect 57595 20540 57626 20592
rect 57626 20540 57647 20592
rect 57383 20322 57435 20374
rect 57595 20322 57626 20374
rect 57626 20322 57647 20374
rect 57383 20105 57435 20157
rect 57595 20105 57626 20157
rect 57626 20105 57647 20157
rect 57383 19887 57435 19939
rect 57595 19887 57626 19939
rect 57626 19887 57647 19939
rect 57383 19670 57435 19722
rect 57595 19670 57626 19722
rect 57626 19670 57647 19722
rect 57383 19452 57435 19504
rect 57595 19452 57626 19504
rect 57626 19452 57647 19504
rect 57383 19234 57435 19286
rect 57595 19234 57626 19286
rect 57626 19234 57647 19286
rect 57383 19016 57435 19068
rect 57595 19016 57626 19068
rect 57626 19016 57647 19068
rect 57383 18799 57435 18851
rect 57595 18799 57626 18851
rect 57626 18799 57647 18851
rect 57383 18581 57435 18633
rect 57595 18581 57626 18633
rect 57626 18581 57647 18633
rect 57383 18364 57435 18416
rect 57595 18364 57626 18416
rect 57626 18364 57647 18416
rect 57383 18146 57435 18198
rect 57595 18146 57626 18198
rect 57626 18146 57647 18198
rect 57383 17928 57435 17980
rect 57595 17928 57626 17980
rect 57626 17928 57647 17980
rect 57383 17711 57435 17763
rect 57595 17711 57626 17763
rect 57626 17711 57647 17763
rect 57383 17493 57435 17545
rect 57595 17493 57626 17545
rect 57626 17493 57647 17545
rect 57383 17275 57435 17327
rect 57595 17275 57626 17327
rect 57626 17275 57647 17327
rect 57383 17058 57435 17110
rect 57595 17058 57626 17110
rect 57626 17058 57647 17110
rect 57383 16840 57435 16892
rect 57595 16840 57626 16892
rect 57626 16840 57647 16892
rect 57383 16623 57435 16675
rect 57595 16623 57626 16675
rect 57626 16623 57647 16675
rect 57383 16405 57435 16457
rect 57595 16405 57626 16457
rect 57626 16405 57647 16457
rect 57383 16187 57435 16239
rect 57595 16187 57626 16239
rect 57626 16187 57647 16239
rect 57383 15970 57435 16022
rect 57595 15970 57626 16022
rect 57626 15970 57647 16022
rect 57383 15752 57435 15804
rect 57595 15752 57626 15804
rect 57626 15752 57647 15804
rect 57383 15534 57435 15586
rect 57595 15534 57626 15586
rect 57626 15534 57647 15586
rect 57383 15317 57435 15369
rect 57595 15317 57626 15369
rect 57626 15317 57647 15369
rect 57383 15099 57435 15151
rect 57595 15099 57626 15151
rect 57626 15099 57647 15151
rect 57383 14881 57435 14933
rect 57595 14881 57626 14933
rect 57626 14881 57647 14933
rect 57383 14664 57435 14716
rect 57595 14664 57626 14716
rect 57626 14664 57647 14716
rect 57383 14446 57435 14498
rect 57595 14446 57626 14498
rect 57626 14446 57647 14498
rect 57383 14229 57435 14281
rect 57595 14229 57626 14281
rect 57626 14229 57647 14281
rect 57383 14011 57435 14063
rect 57595 14011 57626 14063
rect 57626 14011 57647 14063
rect 57383 13793 57435 13845
rect 57595 13793 57626 13845
rect 57626 13793 57647 13845
rect 57383 13576 57435 13628
rect 57595 13576 57626 13628
rect 57626 13576 57647 13628
rect 57383 13358 57435 13410
rect 57595 13358 57626 13410
rect 57626 13358 57647 13410
rect 57383 13140 57435 13192
rect 57595 13140 57626 13192
rect 57626 13140 57647 13192
rect 57383 12923 57435 12975
rect 57595 12923 57626 12975
rect 57626 12923 57647 12975
rect 57383 12705 57435 12757
rect 57595 12705 57626 12757
rect 57626 12705 57647 12757
rect 57383 12488 57435 12540
rect 57595 12488 57626 12540
rect 57626 12488 57647 12540
rect 57383 12270 57435 12322
rect 57595 12270 57626 12322
rect 57626 12270 57647 12322
rect 57383 12052 57435 12104
rect 57595 12052 57626 12104
rect 57626 12052 57647 12104
rect 57383 11835 57435 11887
rect 57595 11835 57626 11887
rect 57626 11835 57647 11887
rect 57383 11617 57435 11669
rect 57595 11617 57626 11669
rect 57626 11617 57647 11669
rect 57383 11399 57435 11451
rect 57595 11399 57626 11451
rect 57626 11399 57647 11451
rect 57383 11182 57435 11234
rect 57595 11182 57626 11234
rect 57626 11182 57647 11234
rect 57383 10964 57435 11016
rect 57595 10964 57626 11016
rect 57626 10964 57647 11016
rect 57383 10746 57435 10798
rect 57595 10746 57626 10798
rect 57626 10746 57647 10798
rect 57383 10529 57435 10581
rect 57595 10529 57626 10581
rect 57626 10529 57647 10581
rect 57383 10311 57435 10363
rect 57595 10311 57626 10363
rect 57626 10311 57647 10363
rect 57383 10094 57435 10146
rect 57595 10094 57626 10146
rect 57626 10094 57647 10146
rect 57383 9876 57435 9928
rect 57595 9876 57626 9928
rect 57626 9876 57647 9928
rect 57383 9658 57435 9710
rect 57595 9658 57626 9710
rect 57626 9658 57647 9710
rect 57383 9441 57435 9493
rect 57595 9441 57626 9493
rect 57626 9441 57647 9493
rect 57383 9223 57435 9275
rect 57595 9223 57626 9275
rect 57626 9223 57647 9275
rect 57383 9005 57435 9057
rect 57595 9005 57626 9057
rect 57626 9005 57647 9057
rect 57383 8788 57435 8840
rect 57595 8788 57626 8840
rect 57626 8788 57647 8840
rect 57383 8570 57435 8622
rect 57595 8570 57626 8622
rect 57626 8570 57647 8622
rect 57383 8352 57435 8404
rect 57595 8352 57626 8404
rect 57626 8352 57647 8404
rect 57383 8135 57435 8187
rect 57595 8135 57626 8187
rect 57626 8135 57647 8187
rect 57383 7917 57435 7969
rect 57595 7917 57626 7969
rect 57626 7917 57647 7969
rect 57383 7700 57435 7752
rect 57595 7700 57626 7752
rect 57626 7700 57647 7752
rect 57383 7482 57435 7534
rect 57595 7482 57626 7534
rect 57626 7482 57647 7534
rect 57383 7264 57435 7316
rect 57595 7264 57626 7316
rect 57626 7264 57647 7316
rect 57383 7047 57435 7099
rect 57595 7047 57626 7099
rect 57626 7047 57647 7099
rect 57383 6829 57435 6881
rect 57595 6829 57626 6881
rect 57626 6829 57647 6881
rect 57383 6611 57435 6663
rect 57595 6611 57626 6663
rect 57626 6611 57647 6663
rect 57383 6394 57435 6446
rect 57595 6394 57626 6446
rect 57626 6394 57647 6446
rect 57383 6176 57435 6228
rect 57595 6176 57626 6228
rect 57626 6176 57647 6228
rect 57383 5959 57435 6011
rect 57595 5959 57626 6011
rect 57626 5959 57647 6011
rect 57383 5741 57435 5793
rect 57595 5741 57626 5793
rect 57626 5741 57647 5793
rect 57383 5523 57435 5575
rect 57595 5523 57626 5575
rect 57626 5523 57647 5575
rect 57383 5306 57435 5358
rect 57595 5306 57626 5358
rect 57626 5306 57647 5358
rect 51654 5147 51810 5199
rect 40622 4852 40778 4904
rect 57998 33380 58050 33432
rect 58210 33380 58262 33432
rect 57998 33163 58050 33215
rect 58210 33163 58262 33215
rect 57998 32945 58050 32997
rect 58210 32945 58262 32997
rect 57998 32727 58050 32779
rect 58210 32727 58262 32779
rect 57998 32510 58050 32562
rect 58210 32510 58262 32562
rect 57998 32292 58050 32344
rect 58210 32292 58262 32344
rect 57998 32075 58050 32127
rect 58210 32075 58262 32127
rect 57998 31857 58050 31909
rect 58210 31857 58262 31909
rect 57998 31639 58050 31691
rect 58210 31639 58262 31691
rect 57998 31422 58050 31474
rect 58210 31422 58262 31474
rect 57998 31204 58050 31256
rect 58210 31204 58262 31256
rect 57998 30986 58050 31038
rect 58210 30986 58262 31038
rect 57998 30769 58050 30821
rect 58210 30769 58262 30821
rect 57998 30551 58050 30603
rect 58210 30551 58262 30603
rect 57998 30334 58050 30386
rect 58210 30334 58262 30386
rect 57998 30116 58050 30168
rect 58210 30116 58262 30168
rect 57998 29898 58050 29950
rect 58210 29898 58262 29950
rect 57998 29681 58050 29733
rect 58210 29681 58262 29733
rect 57998 29463 58050 29515
rect 58210 29463 58262 29515
rect 57998 29245 58050 29297
rect 58210 29245 58262 29297
rect 57998 29028 58050 29080
rect 58210 29028 58262 29080
rect 57998 28810 58050 28862
rect 58210 28810 58262 28862
rect 57998 28592 58050 28644
rect 58210 28592 58262 28644
rect 57998 28375 58050 28427
rect 58210 28375 58262 28427
rect 57998 28157 58050 28209
rect 58210 28157 58262 28209
rect 57998 27940 58050 27992
rect 58210 27940 58262 27992
rect 57998 27722 58050 27774
rect 58210 27722 58262 27774
rect 57998 27504 58050 27556
rect 58210 27504 58262 27556
rect 57998 27287 58050 27339
rect 58210 27287 58262 27339
rect 57998 27069 58050 27121
rect 58210 27069 58262 27121
rect 57998 26851 58050 26903
rect 58210 26851 58262 26903
rect 57998 26634 58050 26686
rect 58210 26634 58262 26686
rect 57998 26416 58050 26468
rect 58210 26416 58262 26468
rect 57998 26198 58050 26250
rect 58210 26198 58262 26250
rect 57998 25981 58050 26033
rect 58210 25981 58262 26033
rect 57998 25763 58050 25815
rect 58210 25763 58262 25815
rect 57998 25546 58050 25598
rect 58210 25546 58262 25598
rect 57998 25328 58050 25380
rect 58210 25328 58262 25380
rect 57998 25110 58050 25162
rect 58210 25110 58262 25162
rect 57998 24893 58050 24945
rect 58210 24893 58262 24945
rect 57998 24675 58050 24727
rect 58210 24675 58262 24727
rect 57998 24457 58050 24509
rect 58210 24457 58262 24509
rect 57998 24240 58050 24292
rect 58210 24240 58262 24292
rect 57998 24022 58050 24074
rect 58210 24022 58262 24074
rect 57998 23805 58050 23857
rect 58210 23805 58262 23857
rect 57998 23587 58050 23639
rect 58210 23587 58262 23639
rect 57998 23369 58050 23421
rect 58210 23369 58262 23421
rect 57998 23152 58050 23204
rect 58210 23152 58262 23204
rect 57998 22934 58050 22986
rect 58210 22934 58262 22986
rect 57998 22716 58050 22768
rect 58210 22716 58262 22768
rect 57998 22499 58050 22551
rect 58210 22499 58262 22551
rect 57998 22281 58050 22333
rect 58210 22281 58262 22333
rect 57998 22063 58050 22115
rect 58210 22063 58262 22115
rect 57998 21846 58050 21898
rect 58210 21846 58262 21898
rect 57998 21628 58050 21680
rect 58210 21628 58262 21680
rect 57998 21411 58050 21463
rect 58210 21411 58262 21463
rect 57998 21193 58050 21245
rect 58210 21193 58262 21245
rect 57998 20975 58050 21027
rect 58210 20975 58262 21027
rect 57998 20758 58050 20810
rect 58210 20758 58262 20810
rect 57998 20540 58050 20592
rect 58210 20540 58262 20592
rect 57998 20322 58050 20374
rect 58210 20322 58262 20374
rect 57998 20105 58050 20157
rect 58210 20105 58262 20157
rect 57998 19887 58050 19939
rect 58210 19887 58262 19939
rect 57998 19670 58050 19722
rect 58210 19670 58262 19722
rect 57998 19452 58050 19504
rect 58210 19452 58262 19504
rect 57998 19234 58050 19286
rect 58210 19234 58262 19286
rect 57998 19016 58050 19068
rect 58210 19016 58262 19068
rect 57998 18799 58050 18851
rect 58210 18799 58262 18851
rect 57998 18581 58050 18633
rect 58210 18581 58262 18633
rect 57998 18364 58050 18416
rect 58210 18364 58262 18416
rect 57998 18146 58050 18198
rect 58210 18146 58262 18198
rect 57998 17928 58050 17980
rect 58210 17928 58262 17980
rect 57998 17711 58050 17763
rect 58210 17711 58262 17763
rect 57998 17493 58050 17545
rect 58210 17493 58262 17545
rect 57998 17275 58050 17327
rect 58210 17275 58262 17327
rect 57998 17058 58050 17110
rect 58210 17058 58262 17110
rect 57998 16840 58050 16892
rect 58210 16840 58262 16892
rect 57998 16623 58050 16675
rect 58210 16623 58262 16675
rect 57998 16405 58050 16457
rect 58210 16405 58262 16457
rect 57998 16187 58050 16239
rect 58210 16187 58262 16239
rect 57998 15970 58050 16022
rect 58210 15970 58262 16022
rect 57998 15752 58050 15804
rect 58210 15752 58262 15804
rect 57998 15534 58050 15586
rect 58210 15534 58262 15586
rect 57998 15317 58050 15369
rect 58210 15317 58262 15369
rect 57998 15099 58050 15151
rect 58210 15099 58262 15151
rect 57998 14881 58050 14933
rect 58210 14881 58262 14933
rect 57998 14664 58050 14716
rect 58210 14664 58262 14716
rect 57998 14446 58050 14498
rect 58210 14446 58262 14498
rect 57998 14229 58050 14281
rect 58210 14229 58262 14281
rect 57998 14011 58050 14063
rect 58210 14011 58262 14063
rect 57998 13793 58050 13845
rect 58210 13793 58262 13845
rect 57998 13576 58050 13628
rect 58210 13576 58262 13628
rect 57998 13358 58050 13410
rect 58210 13358 58262 13410
rect 57998 13140 58050 13192
rect 58210 13140 58262 13192
rect 57998 12923 58050 12975
rect 58210 12923 58262 12975
rect 57998 12705 58050 12757
rect 58210 12705 58262 12757
rect 57998 12488 58050 12540
rect 58210 12488 58262 12540
rect 57998 12270 58050 12322
rect 58210 12270 58262 12322
rect 57998 12052 58050 12104
rect 58210 12052 58262 12104
rect 57998 11835 58050 11887
rect 58210 11835 58262 11887
rect 57998 11617 58050 11669
rect 58210 11617 58262 11669
rect 57998 11399 58050 11451
rect 58210 11399 58262 11451
rect 57998 11182 58050 11234
rect 58210 11182 58262 11234
rect 57998 10964 58050 11016
rect 58210 10964 58262 11016
rect 57998 10746 58050 10798
rect 58210 10746 58262 10798
rect 57998 10529 58050 10581
rect 58210 10529 58262 10581
rect 57998 10311 58050 10363
rect 58210 10311 58262 10363
rect 57998 10094 58050 10146
rect 58210 10094 58262 10146
rect 57998 9876 58050 9928
rect 58210 9876 58262 9928
rect 57998 9658 58050 9710
rect 58210 9658 58262 9710
rect 57998 9441 58050 9493
rect 58210 9441 58262 9493
rect 57998 9223 58050 9275
rect 58210 9223 58262 9275
rect 57998 9005 58050 9057
rect 58210 9005 58262 9057
rect 57998 8788 58050 8840
rect 58210 8788 58262 8840
rect 57998 8570 58050 8622
rect 58210 8570 58262 8622
rect 57998 8352 58050 8404
rect 58210 8352 58262 8404
rect 57998 8135 58050 8187
rect 58210 8135 58262 8187
rect 57998 7917 58050 7969
rect 58210 7917 58262 7969
rect 57998 7700 58050 7752
rect 58210 7700 58262 7752
rect 57998 7482 58050 7534
rect 58210 7482 58262 7534
rect 57998 7264 58050 7316
rect 58210 7264 58262 7316
rect 57998 7047 58050 7099
rect 58210 7047 58262 7099
rect 57998 6829 58050 6881
rect 58210 6829 58262 6881
rect 57998 6611 58050 6663
rect 58210 6611 58262 6663
rect 57998 6394 58050 6446
rect 58210 6394 58262 6446
rect 57998 6176 58050 6228
rect 58210 6176 58262 6228
rect 57998 5959 58050 6011
rect 58210 5959 58262 6011
rect 57998 5741 58050 5793
rect 58210 5741 58262 5793
rect 57998 5523 58050 5575
rect 58210 5523 58262 5575
rect 57998 5306 58050 5358
rect 58210 5306 58262 5358
rect 57383 4535 57435 4587
rect 57595 4535 57626 4587
rect 57626 4535 57647 4587
rect 57383 4318 57435 4370
rect 57595 4318 57626 4370
rect 57626 4318 57647 4370
rect 57383 4100 57435 4152
rect 57595 4100 57626 4152
rect 57626 4100 57647 4152
rect 57383 3882 57435 3934
rect 57595 3882 57626 3934
rect 57626 3882 57647 3934
rect 57383 3665 57435 3717
rect 57595 3665 57626 3717
rect 57626 3665 57647 3717
rect 48668 1172 48720 1224
rect 48792 1172 48844 1224
rect 48916 1172 48968 1224
rect 57998 4535 58050 4587
rect 58210 4535 58262 4587
rect 57998 4318 58050 4370
rect 58210 4318 58262 4370
rect 57998 4100 58050 4152
rect 58210 4100 58262 4152
rect 57998 3882 58050 3934
rect 58210 3882 58262 3934
rect 57998 3665 58050 3717
rect 58210 3665 58262 3717
rect 62150 1637 62306 1689
rect 72215 1637 72371 1689
rect 72665 1637 72821 1689
rect 82730 1637 82886 1689
rect 48668 1048 48720 1100
rect 48792 1048 48844 1100
rect 48916 1048 48968 1100
rect 48668 924 48720 976
rect 48792 924 48844 976
rect 48916 924 48968 976
rect 29090 655 29142 915
rect 29792 655 29844 915
rect 48668 800 48720 852
rect 48792 800 48844 852
rect 48916 800 48968 852
rect 48668 676 48720 728
rect 48792 676 48844 728
rect 48916 676 48968 728
rect 48668 552 48720 604
rect 48792 552 48844 604
rect 48916 552 48968 604
rect 48668 428 48720 480
rect 48792 428 48844 480
rect 48916 428 48968 480
rect 48668 304 48720 356
rect 48792 304 48844 356
rect 48916 304 48968 356
<< metal2 >>
rect 282 53168 86090 53494
rect 706 51976 85666 52976
rect 25313 51579 26039 51627
rect 25313 51572 25400 51579
rect 25452 51572 25524 51579
rect 25576 51572 25648 51579
rect 25700 51572 25772 51579
rect 25824 51572 25896 51579
rect 25948 51572 26039 51579
rect 25313 51516 25398 51572
rect 25454 51516 25522 51572
rect 25578 51516 25646 51572
rect 25702 51516 25770 51572
rect 25826 51516 25894 51572
rect 25950 51516 26039 51572
rect 25313 51455 26039 51516
rect 25313 51448 25400 51455
rect 25452 51448 25524 51455
rect 25576 51448 25648 51455
rect 25700 51448 25772 51455
rect 25824 51448 25896 51455
rect 25948 51448 26039 51455
rect 25313 51392 25398 51448
rect 25454 51392 25522 51448
rect 25578 51392 25646 51448
rect 25702 51392 25770 51448
rect 25826 51392 25894 51448
rect 25950 51392 26039 51448
rect 25313 51331 26039 51392
rect 25313 51324 25400 51331
rect 25452 51324 25524 51331
rect 25576 51324 25648 51331
rect 25700 51324 25772 51331
rect 25824 51324 25896 51331
rect 25948 51324 26039 51331
rect 25313 51268 25398 51324
rect 25454 51268 25522 51324
rect 25578 51268 25646 51324
rect 25702 51268 25770 51324
rect 25826 51268 25894 51324
rect 25950 51268 26039 51324
rect 25313 35275 26039 51268
rect 25313 35219 25384 35275
rect 25440 35219 25508 35275
rect 25564 35219 25632 35275
rect 25688 35219 25756 35275
rect 25812 35219 25880 35275
rect 25936 35219 26039 35275
rect 25313 35151 26039 35219
rect 25313 35095 25384 35151
rect 25440 35095 25508 35151
rect 25564 35095 25632 35151
rect 25688 35095 25756 35151
rect 25812 35095 25880 35151
rect 25936 35095 26039 35151
rect 25313 35027 26039 35095
rect 25313 34971 25384 35027
rect 25440 34971 25508 35027
rect 25564 34971 25632 35027
rect 25688 34971 25756 35027
rect 25812 34971 25880 35027
rect 25936 34971 26039 35027
rect 25313 34903 26039 34971
rect 25313 34847 25384 34903
rect 25440 34847 25508 34903
rect 25564 34847 25632 34903
rect 25688 34847 25756 34903
rect 25812 34847 25880 34903
rect 25936 34847 26039 34903
rect 25313 34779 26039 34847
rect 25313 34723 25384 34779
rect 25440 34723 25508 34779
rect 25564 34723 25632 34779
rect 25688 34723 25756 34779
rect 25812 34723 25880 34779
rect 25936 34723 26039 34779
rect 25313 34655 26039 34723
rect 25313 34599 25384 34655
rect 25440 34599 25508 34655
rect 25564 34599 25632 34655
rect 25688 34599 25756 34655
rect 25812 34599 25880 34655
rect 25936 34599 26039 34655
rect 25313 31248 26039 34599
rect 25313 31192 25398 31248
rect 25454 31192 25522 31248
rect 25578 31192 25646 31248
rect 25702 31192 25770 31248
rect 25826 31192 25894 31248
rect 25950 31192 26039 31248
rect 25313 31124 26039 31192
rect 25313 31068 25398 31124
rect 25454 31068 25522 31124
rect 25578 31068 25646 31124
rect 25702 31068 25770 31124
rect 25826 31068 25894 31124
rect 25950 31068 26039 31124
rect 25313 31000 26039 31068
rect 25313 30944 25398 31000
rect 25454 30944 25522 31000
rect 25578 30944 25646 31000
rect 25702 30944 25770 31000
rect 25826 30944 25894 31000
rect 25950 30944 26039 31000
rect 25313 30793 26039 30944
rect 25313 30737 25398 30793
rect 25454 30737 25522 30793
rect 25578 30737 25646 30793
rect 25702 30737 25770 30793
rect 25826 30737 25894 30793
rect 25950 30737 26039 30793
rect 25313 30669 26039 30737
rect 25313 30613 25398 30669
rect 25454 30613 25522 30669
rect 25578 30613 25646 30669
rect 25702 30613 25770 30669
rect 25826 30613 25894 30669
rect 25950 30613 26039 30669
rect 25313 30545 26039 30613
rect 25313 30489 25398 30545
rect 25454 30489 25522 30545
rect 25578 30489 25646 30545
rect 25702 30489 25770 30545
rect 25826 30489 25894 30545
rect 25950 30489 26039 30545
rect 25313 28263 26039 30489
rect 25313 28207 25404 28263
rect 25460 28207 25528 28263
rect 25584 28207 25652 28263
rect 25708 28207 25776 28263
rect 25832 28207 25900 28263
rect 25956 28207 26039 28263
rect 25313 28139 26039 28207
rect 25313 28083 25404 28139
rect 25460 28083 25528 28139
rect 25584 28083 25652 28139
rect 25708 28083 25776 28139
rect 25832 28083 25900 28139
rect 25956 28083 26039 28139
rect 25313 28015 26039 28083
rect 25313 27959 25404 28015
rect 25460 27959 25528 28015
rect 25584 27959 25652 28015
rect 25708 27959 25776 28015
rect 25832 27959 25900 28015
rect 25956 27959 26039 28015
rect 25313 27891 26039 27959
rect 25313 27835 25404 27891
rect 25460 27835 25528 27891
rect 25584 27835 25652 27891
rect 25708 27835 25776 27891
rect 25832 27835 25900 27891
rect 25956 27835 26039 27891
rect 25313 27767 26039 27835
rect 25313 27711 25404 27767
rect 25460 27711 25528 27767
rect 25584 27711 25652 27767
rect 25708 27711 25776 27767
rect 25832 27711 25900 27767
rect 25956 27711 26039 27767
rect 25313 27643 26039 27711
rect 25313 27587 25404 27643
rect 25460 27587 25528 27643
rect 25584 27587 25652 27643
rect 25708 27587 25776 27643
rect 25832 27587 25900 27643
rect 25956 27587 26039 27643
rect 25313 27519 26039 27587
rect 25313 27463 25404 27519
rect 25460 27463 25528 27519
rect 25584 27463 25652 27519
rect 25708 27463 25776 27519
rect 25832 27463 25900 27519
rect 25956 27463 26039 27519
rect 25313 27395 26039 27463
rect 25313 27339 25404 27395
rect 25460 27339 25528 27395
rect 25584 27339 25652 27395
rect 25708 27339 25776 27395
rect 25832 27339 25900 27395
rect 25956 27339 26039 27395
rect 25313 27271 26039 27339
rect 25313 27215 25404 27271
rect 25460 27215 25528 27271
rect 25584 27215 25652 27271
rect 25708 27215 25776 27271
rect 25832 27215 25900 27271
rect 25956 27215 26039 27271
rect 25313 27147 26039 27215
rect 25313 27091 25404 27147
rect 25460 27091 25528 27147
rect 25584 27091 25652 27147
rect 25708 27091 25776 27147
rect 25832 27091 25900 27147
rect 25956 27091 26039 27147
rect 25313 27023 26039 27091
rect 25313 26967 25404 27023
rect 25460 26967 25528 27023
rect 25584 26967 25652 27023
rect 25708 26967 25776 27023
rect 25832 26967 25900 27023
rect 25956 26967 26039 27023
rect 25313 26899 26039 26967
rect 25313 26843 25404 26899
rect 25460 26843 25528 26899
rect 25584 26843 25652 26899
rect 25708 26843 25776 26899
rect 25832 26843 25900 26899
rect 25956 26843 26039 26899
rect 25313 26775 26039 26843
rect 25313 26719 25404 26775
rect 25460 26719 25528 26775
rect 25584 26719 25652 26775
rect 25708 26719 25776 26775
rect 25832 26719 25900 26775
rect 25956 26719 26039 26775
rect 25313 26651 26039 26719
rect 25313 26595 25404 26651
rect 25460 26595 25528 26651
rect 25584 26595 25652 26651
rect 25708 26595 25776 26651
rect 25832 26595 25900 26651
rect 25956 26595 26039 26651
rect 25313 26527 26039 26595
rect 25313 26471 25404 26527
rect 25460 26471 25528 26527
rect 25584 26471 25652 26527
rect 25708 26471 25776 26527
rect 25832 26471 25900 26527
rect 25956 26471 26039 26527
rect 25313 26433 26039 26471
rect 26823 34011 27163 51976
rect 26823 33955 26859 34011
rect 26915 33955 27071 34011
rect 27127 33955 27163 34011
rect 26823 33793 27163 33955
rect 26823 33737 26859 33793
rect 26915 33737 27071 33793
rect 27127 33737 27163 33793
rect 26823 33576 27163 33737
rect 26823 33520 26859 33576
rect 26915 33520 27071 33576
rect 27127 33520 27163 33576
rect 26823 33432 27163 33520
rect 26823 33380 26861 33432
rect 26913 33380 27073 33432
rect 27125 33380 27163 33432
rect 26823 33358 27163 33380
rect 26823 33302 26859 33358
rect 26915 33302 27071 33358
rect 27127 33302 27163 33358
rect 26823 33215 27163 33302
rect 26823 33163 26861 33215
rect 26913 33163 27073 33215
rect 27125 33163 27163 33215
rect 26823 33140 27163 33163
rect 26823 33084 26859 33140
rect 26915 33084 27071 33140
rect 27127 33084 27163 33140
rect 26823 32997 27163 33084
rect 26823 32945 26861 32997
rect 26913 32945 27073 32997
rect 27125 32945 27163 32997
rect 26823 32922 27163 32945
rect 26823 32866 26859 32922
rect 26915 32866 27071 32922
rect 27127 32866 27163 32922
rect 26823 32779 27163 32866
rect 26823 32727 26861 32779
rect 26913 32727 27073 32779
rect 27125 32727 27163 32779
rect 26823 32705 27163 32727
rect 26823 32649 26859 32705
rect 26915 32649 27071 32705
rect 27127 32649 27163 32705
rect 26823 32562 27163 32649
rect 26823 32510 26861 32562
rect 26913 32510 27073 32562
rect 27125 32510 27163 32562
rect 26823 32487 27163 32510
rect 26823 32431 26859 32487
rect 26915 32431 27071 32487
rect 27127 32431 27163 32487
rect 26823 32344 27163 32431
rect 26823 32292 26861 32344
rect 26913 32292 27073 32344
rect 27125 32292 27163 32344
rect 26823 32127 27163 32292
rect 26823 32088 26861 32127
rect 26913 32088 27073 32127
rect 27125 32088 27163 32127
rect 26823 32032 26859 32088
rect 26915 32032 27071 32088
rect 27127 32032 27163 32088
rect 26823 31909 27163 32032
rect 26823 31870 26861 31909
rect 26913 31870 27073 31909
rect 27125 31870 27163 31909
rect 26823 31814 26859 31870
rect 26915 31814 27071 31870
rect 27127 31814 27163 31870
rect 26823 31691 27163 31814
rect 26823 31652 26861 31691
rect 26913 31652 27073 31691
rect 27125 31652 27163 31691
rect 26823 31596 26859 31652
rect 26915 31596 27071 31652
rect 27127 31596 27163 31652
rect 26823 31474 27163 31596
rect 26823 31422 26861 31474
rect 26913 31422 27073 31474
rect 27125 31422 27163 31474
rect 26823 31256 27163 31422
rect 26823 31204 26861 31256
rect 26913 31204 27073 31256
rect 27125 31204 27163 31256
rect 26823 31038 27163 31204
rect 26823 30986 26861 31038
rect 26913 30986 27073 31038
rect 27125 30986 27163 31038
rect 26823 30821 27163 30986
rect 26823 30769 26861 30821
rect 26913 30769 27073 30821
rect 27125 30769 27163 30821
rect 26823 30603 27163 30769
rect 26823 30551 26861 30603
rect 26913 30551 27073 30603
rect 27125 30551 27163 30603
rect 26823 30386 27163 30551
rect 26823 30334 26861 30386
rect 26913 30334 27073 30386
rect 27125 30334 27163 30386
rect 26823 30168 27163 30334
rect 26823 30116 26861 30168
rect 26913 30116 27073 30168
rect 27125 30116 27163 30168
rect 26823 29968 27163 30116
rect 26823 29912 26859 29968
rect 26915 29912 27071 29968
rect 27127 29912 27163 29968
rect 26823 29898 26861 29912
rect 26913 29898 27073 29912
rect 27125 29898 27163 29912
rect 26823 29750 27163 29898
rect 26823 29694 26859 29750
rect 26915 29694 27071 29750
rect 27127 29694 27163 29750
rect 26823 29681 26861 29694
rect 26913 29681 27073 29694
rect 27125 29681 27163 29694
rect 26823 29533 27163 29681
rect 26823 29477 26859 29533
rect 26915 29477 27071 29533
rect 27127 29477 27163 29533
rect 26823 29463 26861 29477
rect 26913 29463 27073 29477
rect 27125 29463 27163 29477
rect 26823 29315 27163 29463
rect 26823 29259 26859 29315
rect 26915 29259 27071 29315
rect 27127 29259 27163 29315
rect 26823 29245 26861 29259
rect 26913 29245 27073 29259
rect 27125 29245 27163 29259
rect 26823 29098 27163 29245
rect 26823 29042 26859 29098
rect 26915 29042 27071 29098
rect 27127 29042 27163 29098
rect 26823 29028 26861 29042
rect 26913 29028 27073 29042
rect 27125 29028 27163 29042
rect 26823 28880 27163 29028
rect 26823 28824 26859 28880
rect 26915 28824 27071 28880
rect 27127 28824 27163 28880
rect 26823 28810 26861 28824
rect 26913 28810 27073 28824
rect 27125 28810 27163 28824
rect 26823 28662 27163 28810
rect 26823 28606 26859 28662
rect 26915 28606 27071 28662
rect 27127 28606 27163 28662
rect 26823 28592 26861 28606
rect 26913 28592 27073 28606
rect 27125 28592 27163 28606
rect 26823 28444 27163 28592
rect 26823 28388 26859 28444
rect 26915 28388 27071 28444
rect 27127 28388 27163 28444
rect 26823 28375 26861 28388
rect 26913 28375 27073 28388
rect 27125 28375 27163 28388
rect 26823 28227 27163 28375
rect 26823 28171 26859 28227
rect 26915 28171 27071 28227
rect 27127 28171 27163 28227
rect 26823 28157 26861 28171
rect 26913 28157 27073 28171
rect 27125 28157 27163 28171
rect 26823 28009 27163 28157
rect 26823 27953 26859 28009
rect 26915 27953 27071 28009
rect 27127 27953 27163 28009
rect 26823 27940 26861 27953
rect 26913 27940 27073 27953
rect 27125 27940 27163 27953
rect 26823 27792 27163 27940
rect 26823 27736 26859 27792
rect 26915 27736 27071 27792
rect 27127 27736 27163 27792
rect 26823 27722 26861 27736
rect 26913 27722 27073 27736
rect 27125 27722 27163 27736
rect 26823 27574 27163 27722
rect 26823 27518 26859 27574
rect 26915 27518 27071 27574
rect 27127 27518 27163 27574
rect 26823 27504 26861 27518
rect 26913 27504 27073 27518
rect 27125 27504 27163 27518
rect 26823 27339 27163 27504
rect 26823 27287 26861 27339
rect 26913 27287 27073 27339
rect 27125 27287 27163 27339
rect 26823 27121 27163 27287
rect 26823 27069 26861 27121
rect 26913 27069 27073 27121
rect 27125 27069 27163 27121
rect 26823 26903 27163 27069
rect 26823 26851 26861 26903
rect 26913 26851 27073 26903
rect 27125 26851 27163 26903
rect 26823 26686 27163 26851
rect 26823 26634 26861 26686
rect 26913 26634 27073 26686
rect 27125 26634 27163 26686
rect 26823 26468 27163 26634
rect 26823 26416 26861 26468
rect 26913 26416 27073 26468
rect 27125 26416 27163 26468
rect 26435 26286 26643 26321
rect 26435 26126 26450 26286
rect 26610 26126 26643 26286
rect 26077 25967 26285 26002
rect 26077 25807 26092 25967
rect 26252 25807 26285 25967
rect 25741 25647 25949 25676
rect 25741 25487 25756 25647
rect 25916 25487 25949 25647
rect 25406 25328 25614 25357
rect 25406 25168 25421 25328
rect 25581 25168 25614 25328
rect 25066 24637 25274 24666
rect 25066 24477 25081 24637
rect 25241 24477 25274 24637
rect 24729 24316 24937 24345
rect 24729 24156 24744 24316
rect 24904 24156 24937 24316
rect 24401 23995 24609 24024
rect 24401 23835 24416 23995
rect 24576 23835 24609 23995
rect 24042 23673 24250 23702
rect 24042 23513 24057 23673
rect 24217 23513 24250 23673
rect 24042 17317 24250 23513
rect 24401 17656 24609 23835
rect 24729 17977 24937 24156
rect 25066 18350 25274 24477
rect 25406 18684 25614 25168
rect 25741 19027 25949 25487
rect 26077 19347 26285 25807
rect 26435 19692 26643 26126
rect 26435 19532 26465 19692
rect 26625 19532 26643 19692
rect 26435 19502 26643 19532
rect 26823 26250 27163 26416
rect 26823 26198 26861 26250
rect 26913 26198 27073 26250
rect 27125 26198 27163 26250
rect 26823 26033 27163 26198
rect 26823 25981 26861 26033
rect 26913 25981 27073 26033
rect 27125 25981 27163 26033
rect 26823 25815 27163 25981
rect 26823 25763 26861 25815
rect 26913 25763 27073 25815
rect 27125 25763 27163 25815
rect 26823 25598 27163 25763
rect 26823 25546 26861 25598
rect 26913 25546 27073 25598
rect 27125 25546 27163 25598
rect 26823 25380 27163 25546
rect 26823 25328 26861 25380
rect 26913 25328 27073 25380
rect 27125 25328 27163 25380
rect 26823 25162 27163 25328
rect 26823 25110 26861 25162
rect 26913 25110 27073 25162
rect 27125 25110 27163 25162
rect 26823 24945 27163 25110
rect 26823 24893 26861 24945
rect 26913 24893 27073 24945
rect 27125 24893 27163 24945
rect 26823 24727 27163 24893
rect 26823 24675 26861 24727
rect 26913 24675 27073 24727
rect 27125 24675 27163 24727
rect 26823 24509 27163 24675
rect 26823 24457 26861 24509
rect 26913 24457 27073 24509
rect 27125 24457 27163 24509
rect 26823 24292 27163 24457
rect 26823 24240 26861 24292
rect 26913 24240 27073 24292
rect 27125 24240 27163 24292
rect 26823 24075 27163 24240
rect 26823 23187 26858 24075
rect 27122 24074 27163 24075
rect 27125 24022 27163 24074
rect 27122 23857 27163 24022
rect 27125 23805 27163 23857
rect 27122 23639 27163 23805
rect 27125 23587 27163 23639
rect 27122 23421 27163 23587
rect 27125 23369 27163 23421
rect 27122 23204 27163 23369
rect 26823 23152 26861 23187
rect 26913 23152 27073 23187
rect 27125 23152 27163 23204
rect 26823 22986 27163 23152
rect 26823 22934 26861 22986
rect 26913 22934 27073 22986
rect 27125 22934 27163 22986
rect 26823 22768 27163 22934
rect 26823 22716 26861 22768
rect 26913 22716 27073 22768
rect 27125 22716 27163 22768
rect 26823 22551 27163 22716
rect 26823 22499 26861 22551
rect 26913 22499 27073 22551
rect 27125 22499 27163 22551
rect 26823 22333 27163 22499
rect 26823 22281 26861 22333
rect 26913 22281 27073 22333
rect 27125 22281 27163 22333
rect 26823 22115 27163 22281
rect 26823 22063 26861 22115
rect 26913 22063 27073 22115
rect 27125 22063 27163 22115
rect 26823 21898 27163 22063
rect 26823 21846 26861 21898
rect 26913 21846 27073 21898
rect 27125 21846 27163 21898
rect 26823 21680 27163 21846
rect 26823 21628 26861 21680
rect 26913 21628 27073 21680
rect 27125 21628 27163 21680
rect 26823 21463 27163 21628
rect 26823 21411 26861 21463
rect 26913 21411 27073 21463
rect 27125 21411 27163 21463
rect 26823 21245 27163 21411
rect 26823 21193 26861 21245
rect 26913 21193 27073 21245
rect 27125 21193 27163 21245
rect 26823 21027 27163 21193
rect 26823 20975 26861 21027
rect 26913 20975 27073 21027
rect 27125 20975 27163 21027
rect 26823 20810 27163 20975
rect 26823 20758 26861 20810
rect 26913 20758 27073 20810
rect 27125 20758 27163 20810
rect 26823 20592 27163 20758
rect 26823 20540 26861 20592
rect 26913 20570 27073 20592
rect 26913 20540 26924 20570
rect 27125 20540 27163 20592
rect 26823 20410 26924 20540
rect 27084 20410 27163 20540
rect 26823 20374 27163 20410
rect 26823 20322 26861 20374
rect 26913 20322 27073 20374
rect 27125 20322 27163 20374
rect 26823 20226 27163 20322
rect 26823 20157 26924 20226
rect 27084 20157 27163 20226
rect 26823 20105 26861 20157
rect 26913 20105 26924 20157
rect 27125 20105 27163 20157
rect 26823 20066 26924 20105
rect 27084 20066 27163 20105
rect 26823 19939 27163 20066
rect 26823 19887 26861 19939
rect 26913 19887 27073 19939
rect 27125 19887 27163 19939
rect 26823 19722 27163 19887
rect 26823 19670 26861 19722
rect 26913 19670 27073 19722
rect 27125 19670 27163 19722
rect 26823 19504 27163 19670
rect 26077 19187 26107 19347
rect 26267 19187 26285 19347
rect 26077 19162 26285 19187
rect 26823 19452 26861 19504
rect 26913 19452 27073 19504
rect 27125 19452 27163 19504
rect 26823 19286 27163 19452
rect 26823 19234 26861 19286
rect 26913 19234 27073 19286
rect 27125 19234 27163 19286
rect 25741 18867 25771 19027
rect 25931 18867 25949 19027
rect 25741 18822 25949 18867
rect 26823 19068 27163 19234
rect 26823 19016 26861 19068
rect 26913 19016 27073 19068
rect 27125 19016 27163 19068
rect 26823 18851 27163 19016
rect 25406 18524 25434 18684
rect 25594 18524 25614 18684
rect 25406 18482 25614 18524
rect 26823 18799 26861 18851
rect 26913 18799 27073 18851
rect 27125 18799 27163 18851
rect 26823 18633 27163 18799
rect 26823 18581 26861 18633
rect 26913 18581 27073 18633
rect 27125 18581 27163 18633
rect 25066 18190 25094 18350
rect 25254 18190 25274 18350
rect 25066 18142 25274 18190
rect 26823 18416 27163 18581
rect 26823 18364 26861 18416
rect 26913 18364 27073 18416
rect 27125 18364 27163 18416
rect 26823 18198 27163 18364
rect 26823 18146 26861 18198
rect 26913 18146 27073 18198
rect 27125 18146 27163 18198
rect 24729 17817 24757 17977
rect 24917 17817 24937 17977
rect 24729 17803 24937 17817
rect 26823 17980 27163 18146
rect 26823 17928 26861 17980
rect 26913 17928 27073 17980
rect 27125 17928 27163 17980
rect 24401 17496 24429 17656
rect 24589 17496 24609 17656
rect 24401 17462 24609 17496
rect 26823 17763 27163 17928
rect 26823 17711 26861 17763
rect 26913 17711 27073 17763
rect 27125 17711 27163 17763
rect 26823 17545 27163 17711
rect 26823 17493 26861 17545
rect 26913 17493 27073 17545
rect 27125 17493 27163 17545
rect 24042 17157 24069 17317
rect 24229 17157 24250 17317
rect 24042 17122 24250 17157
rect 26823 17327 27163 17493
rect 26823 17275 26861 17327
rect 26913 17275 27073 17327
rect 27125 17275 27163 17327
rect 26823 17110 27163 17275
rect 26823 17058 26861 17110
rect 26913 17058 27073 17110
rect 27125 17058 27163 17110
rect 26823 16892 27163 17058
rect 26823 16840 26861 16892
rect 26913 16840 27073 16892
rect 27125 16840 27163 16892
rect 26823 16675 27163 16840
rect 26823 16623 26861 16675
rect 26913 16623 27073 16675
rect 27125 16623 27163 16675
rect 26823 16457 27163 16623
rect 26823 16405 26861 16457
rect 26913 16405 27073 16457
rect 27125 16405 27163 16457
rect 26823 16239 27163 16405
rect 26823 16187 26861 16239
rect 26913 16187 27073 16239
rect 27125 16187 27163 16239
rect 26823 16022 27163 16187
rect 26823 15970 26861 16022
rect 26913 15970 27073 16022
rect 27125 15970 27163 16022
rect 26823 15804 27163 15970
rect 26823 15752 26861 15804
rect 26913 15752 27073 15804
rect 27125 15752 27163 15804
rect 26823 15586 27163 15752
rect 26823 15534 26861 15586
rect 26913 15534 27073 15586
rect 27125 15534 27163 15586
rect 26823 15369 27163 15534
rect 26823 15317 26861 15369
rect 26913 15317 27073 15369
rect 27125 15317 27163 15369
rect 26823 15151 27163 15317
rect 26823 15099 26861 15151
rect 26913 15099 27073 15151
rect 27125 15099 27163 15151
rect 26823 14933 27163 15099
rect 26823 14881 26861 14933
rect 26913 14881 27073 14933
rect 27125 14881 27163 14933
rect 26823 14716 27163 14881
rect 26823 14664 26861 14716
rect 26913 14664 27073 14716
rect 27125 14664 27163 14716
rect 26823 14498 27163 14664
rect 26823 14446 26861 14498
rect 26913 14446 27073 14498
rect 27125 14446 27163 14498
rect 26823 14281 27163 14446
rect 26823 14229 26861 14281
rect 26913 14229 27073 14281
rect 27125 14229 27163 14281
rect 26823 14119 27163 14229
rect 26823 14063 26859 14119
rect 26915 14063 27071 14119
rect 27127 14063 27163 14119
rect 26823 14011 26861 14063
rect 26913 14011 27073 14063
rect 27125 14011 27163 14063
rect 26823 13902 27163 14011
rect 26823 13846 26859 13902
rect 26915 13846 27071 13902
rect 27127 13846 27163 13902
rect 26823 13845 27163 13846
rect 26823 13793 26861 13845
rect 26913 13793 27073 13845
rect 27125 13793 27163 13845
rect 26823 13684 27163 13793
rect 26823 13628 26859 13684
rect 26915 13628 27071 13684
rect 27127 13628 27163 13684
rect 26823 13576 26861 13628
rect 26913 13576 27073 13628
rect 27125 13576 27163 13628
rect 26823 13467 27163 13576
rect 26823 13411 26859 13467
rect 26915 13411 27071 13467
rect 27127 13411 27163 13467
rect 26823 13410 27163 13411
rect 26823 13358 26861 13410
rect 26913 13358 27073 13410
rect 27125 13358 27163 13410
rect 26823 13249 27163 13358
rect 26823 13193 26859 13249
rect 26915 13193 27071 13249
rect 27127 13193 27163 13249
rect 26823 13192 27163 13193
rect 26823 13140 26861 13192
rect 26913 13140 27073 13192
rect 27125 13140 27163 13192
rect 26823 13031 27163 13140
rect 26823 12975 26859 13031
rect 26915 12975 27071 13031
rect 27127 12975 27163 13031
rect 26823 12923 26861 12975
rect 26913 12923 27073 12975
rect 27125 12923 27163 12975
rect 26823 12813 27163 12923
rect 26823 12757 26859 12813
rect 26915 12757 27071 12813
rect 27127 12757 27163 12813
rect 26823 12705 26861 12757
rect 26913 12705 27073 12757
rect 27125 12705 27163 12757
rect 26823 12596 27163 12705
rect 26823 12540 26859 12596
rect 26915 12540 27071 12596
rect 27127 12540 27163 12596
rect 26823 12488 26861 12540
rect 26913 12488 27073 12540
rect 27125 12488 27163 12540
rect 26823 12378 27163 12488
rect 26823 12322 26859 12378
rect 26915 12322 27071 12378
rect 27127 12322 27163 12378
rect 26823 12270 26861 12322
rect 26913 12270 27073 12322
rect 27125 12270 27163 12322
rect 26823 12161 27163 12270
rect 26823 12105 26859 12161
rect 26915 12105 27071 12161
rect 27127 12105 27163 12161
rect 26823 12104 27163 12105
rect 26823 12052 26861 12104
rect 26913 12052 27073 12104
rect 27125 12052 27163 12104
rect 26823 11887 27163 12052
rect 26823 11835 26861 11887
rect 26913 11835 27073 11887
rect 27125 11835 27163 11887
rect 26823 11669 27163 11835
rect 26823 11617 26861 11669
rect 26913 11617 27073 11669
rect 27125 11617 27163 11669
rect 26823 11451 27163 11617
rect 26823 11399 26861 11451
rect 26913 11399 27073 11451
rect 27125 11399 27163 11451
rect 26823 11234 27163 11399
rect 26823 11182 26861 11234
rect 26913 11182 27073 11234
rect 27125 11182 27163 11234
rect 26823 11016 27163 11182
rect 26823 10964 26861 11016
rect 26913 10964 27073 11016
rect 27125 10964 27163 11016
rect 26823 10798 27163 10964
rect 26823 10746 26861 10798
rect 26913 10746 27073 10798
rect 27125 10746 27163 10798
rect 26823 10581 27163 10746
rect 26823 10529 26861 10581
rect 26913 10529 27073 10581
rect 27125 10529 27163 10581
rect 26823 10363 27163 10529
rect 26823 10311 26861 10363
rect 26913 10311 27073 10363
rect 27125 10311 27163 10363
rect 26823 10146 27163 10311
rect 26823 10094 26861 10146
rect 26913 10094 27073 10146
rect 27125 10094 27163 10146
rect 26823 9928 27163 10094
rect 26823 9876 26861 9928
rect 26913 9876 27073 9928
rect 27125 9876 27163 9928
rect 26823 9710 27163 9876
rect 26823 9658 26861 9710
rect 26913 9658 27073 9710
rect 27125 9658 27163 9710
rect 26823 9493 27163 9658
rect 26823 9441 26861 9493
rect 26913 9441 27073 9493
rect 27125 9441 27163 9493
rect 26823 9407 27163 9441
rect 26823 9351 26859 9407
rect 26915 9351 27071 9407
rect 27127 9351 27163 9407
rect 26823 9275 27163 9351
rect 26823 9223 26861 9275
rect 26913 9223 27073 9275
rect 27125 9223 27163 9275
rect 26823 9190 27163 9223
rect 26823 9134 26859 9190
rect 26915 9134 27071 9190
rect 27127 9134 27163 9190
rect 26823 9057 27163 9134
rect 26823 9005 26861 9057
rect 26913 9005 27073 9057
rect 27125 9005 27163 9057
rect 26823 8972 27163 9005
rect 26823 8916 26859 8972
rect 26915 8916 27071 8972
rect 27127 8916 27163 8972
rect 26823 8840 27163 8916
rect 26823 8788 26861 8840
rect 26913 8788 27073 8840
rect 27125 8788 27163 8840
rect 26823 8754 27163 8788
rect 26823 8698 26859 8754
rect 26915 8698 27071 8754
rect 27127 8698 27163 8754
rect 26823 8622 27163 8698
rect 26823 8570 26861 8622
rect 26913 8570 27073 8622
rect 27125 8570 27163 8622
rect 26823 8536 27163 8570
rect 26823 8480 26859 8536
rect 26915 8480 27071 8536
rect 27127 8480 27163 8536
rect 26823 8404 27163 8480
rect 26823 8352 26861 8404
rect 26913 8352 27073 8404
rect 27125 8352 27163 8404
rect 26823 8319 27163 8352
rect 26823 8263 26859 8319
rect 26915 8263 27071 8319
rect 27127 8263 27163 8319
rect 26823 8187 27163 8263
rect 26823 8135 26861 8187
rect 26913 8135 27073 8187
rect 27125 8135 27163 8187
rect 26823 7969 27163 8135
rect 26823 7917 26861 7969
rect 26913 7917 27073 7969
rect 27125 7917 27163 7969
rect 26823 7752 27163 7917
rect 26823 7700 26861 7752
rect 26913 7700 27073 7752
rect 27125 7700 27163 7752
rect 26823 7534 27163 7700
rect 26823 7482 26861 7534
rect 26913 7482 27073 7534
rect 27125 7482 27163 7534
rect 26823 7316 27163 7482
rect 26823 7264 26861 7316
rect 26913 7264 27073 7316
rect 27125 7264 27163 7316
rect 26823 7099 27163 7264
rect 26823 7047 26861 7099
rect 26913 7047 27073 7099
rect 27125 7047 27163 7099
rect 26823 6881 27163 7047
rect 26823 6829 26861 6881
rect 26913 6829 27073 6881
rect 27125 6829 27163 6881
rect 26823 6663 27163 6829
rect 26823 6611 26861 6663
rect 26913 6611 27073 6663
rect 27125 6611 27163 6663
rect 26823 6446 27163 6611
rect 26823 6394 26861 6446
rect 26913 6394 27073 6446
rect 27125 6394 27163 6446
rect 26823 6228 27163 6394
rect 26823 6176 26861 6228
rect 26913 6176 27073 6228
rect 27125 6176 27163 6228
rect 26823 6011 27163 6176
rect 26823 5959 26861 6011
rect 26913 5959 27073 6011
rect 27125 5959 27163 6011
rect 26823 5793 27163 5959
rect 26823 5741 26861 5793
rect 26913 5741 27073 5793
rect 27125 5741 27163 5793
rect 26823 5575 27163 5741
rect 26823 5539 26861 5575
rect 26913 5539 27073 5575
rect 27125 5539 27163 5575
rect 26823 5483 26859 5539
rect 26915 5483 27071 5539
rect 27127 5483 27163 5539
rect 26823 5358 27163 5483
rect 26823 5321 26861 5358
rect 26913 5321 27073 5358
rect 27125 5321 27163 5358
rect 26823 5265 26859 5321
rect 26915 5265 27071 5321
rect 27127 5265 27163 5321
rect 26823 5226 27163 5265
rect 27387 51455 29146 51494
rect 27387 51399 27788 51455
rect 27844 51399 27999 51455
rect 28055 51399 28210 51455
rect 28266 51399 28421 51455
rect 28477 51399 28632 51455
rect 28688 51399 28843 51455
rect 28899 51399 29054 51455
rect 29110 51399 29146 51455
rect 27387 51360 29146 51399
rect 27387 49694 27828 51360
rect 29486 51285 30364 51976
rect 30769 51285 32888 51976
rect 35128 51285 36415 51976
rect 38953 51471 39618 51976
rect 48789 51285 49990 51976
rect 52226 51285 54354 51976
rect 54758 51285 55638 51976
rect 55977 51455 57371 51494
rect 55977 51399 56013 51455
rect 56069 51399 56224 51455
rect 56280 51399 56435 51455
rect 56491 51399 56646 51455
rect 56702 51399 56857 51455
rect 56913 51399 57068 51455
rect 57124 51399 57279 51455
rect 57335 51399 57371 51455
rect 55977 51360 57371 51399
rect 41865 50613 42045 50623
rect 41865 50453 41875 50613
rect 42035 50453 42045 50613
rect 41865 50443 42045 50453
rect 27387 49655 29146 49694
rect 27387 49599 27788 49655
rect 27844 49599 27999 49655
rect 28055 49599 28210 49655
rect 28266 49599 28421 49655
rect 28477 49599 28632 49655
rect 28688 49599 28843 49655
rect 28899 49599 29054 49655
rect 29110 49599 29146 49655
rect 27387 49560 29146 49599
rect 55977 49655 57371 49694
rect 55977 49599 56013 49655
rect 56069 49599 56224 49655
rect 56280 49599 56435 49655
rect 56491 49599 56646 49655
rect 56702 49599 56857 49655
rect 56913 49599 57068 49655
rect 57124 49599 57279 49655
rect 57335 49599 57371 49655
rect 55977 49560 57371 49599
rect 27387 47894 27828 49560
rect 27387 47855 29146 47894
rect 27387 47799 27788 47855
rect 27844 47799 27999 47855
rect 28055 47799 28210 47855
rect 28266 47799 28421 47855
rect 28477 47799 28632 47855
rect 28688 47799 28843 47855
rect 28899 47799 29054 47855
rect 29110 47799 29146 47855
rect 27387 47760 29146 47799
rect 55977 47855 57371 47894
rect 55977 47799 56013 47855
rect 56069 47799 56224 47855
rect 56280 47799 56435 47855
rect 56491 47799 56646 47855
rect 56702 47799 56857 47855
rect 56913 47799 57068 47855
rect 57124 47799 57279 47855
rect 57335 47799 57371 47855
rect 55977 47760 57371 47799
rect 27387 46094 27828 47760
rect 27387 46055 29146 46094
rect 27387 45999 27788 46055
rect 27844 45999 27999 46055
rect 28055 45999 28210 46055
rect 28266 45999 28421 46055
rect 28477 45999 28632 46055
rect 28688 45999 28843 46055
rect 28899 45999 29054 46055
rect 29110 45999 29146 46055
rect 27387 45960 29146 45999
rect 55977 46055 57371 46094
rect 55977 45999 56013 46055
rect 56069 45999 56224 46055
rect 56280 45999 56435 46055
rect 56491 45999 56646 46055
rect 56702 45999 56857 46055
rect 56913 45999 57068 46055
rect 57124 45999 57279 46055
rect 57335 45999 57371 46055
rect 55977 45960 57371 45999
rect 27387 44294 27828 45960
rect 27387 44255 29146 44294
rect 27387 44199 27788 44255
rect 27844 44199 27999 44255
rect 28055 44199 28210 44255
rect 28266 44199 28421 44255
rect 28477 44199 28632 44255
rect 28688 44199 28843 44255
rect 28899 44199 29054 44255
rect 29110 44199 29146 44255
rect 27387 44160 29146 44199
rect 55977 44255 57371 44294
rect 55977 44199 56013 44255
rect 56069 44199 56224 44255
rect 56280 44199 56435 44255
rect 56491 44199 56646 44255
rect 56702 44199 56857 44255
rect 56913 44199 57068 44255
rect 57124 44199 57279 44255
rect 57335 44199 57371 44255
rect 55977 44160 57371 44199
rect 27387 42494 27828 44160
rect 27387 42455 29146 42494
rect 27387 42399 27788 42455
rect 27844 42399 27999 42455
rect 28055 42399 28210 42455
rect 28266 42399 28421 42455
rect 28477 42399 28632 42455
rect 28688 42399 28843 42455
rect 28899 42399 29054 42455
rect 29110 42399 29146 42455
rect 27387 42360 29146 42399
rect 55977 42455 57371 42494
rect 55977 42399 56013 42455
rect 56069 42399 56224 42455
rect 56280 42399 56435 42455
rect 56491 42399 56646 42455
rect 56702 42399 56857 42455
rect 56913 42399 57068 42455
rect 57124 42399 57279 42455
rect 57335 42399 57371 42455
rect 55977 42360 57371 42399
rect 27387 40694 27828 42360
rect 27387 40655 29146 40694
rect 27387 40599 27788 40655
rect 27844 40599 27999 40655
rect 28055 40599 28210 40655
rect 28266 40599 28421 40655
rect 28477 40599 28632 40655
rect 28688 40599 28843 40655
rect 28899 40599 29054 40655
rect 29110 40599 29146 40655
rect 27387 40560 29146 40599
rect 55977 40655 57371 40694
rect 55977 40599 56013 40655
rect 56069 40599 56224 40655
rect 56280 40599 56435 40655
rect 56491 40599 56646 40655
rect 56702 40599 56857 40655
rect 56913 40599 57068 40655
rect 57124 40599 57279 40655
rect 57335 40599 57371 40655
rect 55977 40560 57371 40599
rect 27387 38894 27828 40560
rect 27387 38855 29146 38894
rect 27387 38799 27788 38855
rect 27844 38799 27999 38855
rect 28055 38799 28210 38855
rect 28266 38799 28421 38855
rect 28477 38799 28632 38855
rect 28688 38799 28843 38855
rect 28899 38799 29054 38855
rect 29110 38799 29146 38855
rect 27387 38760 29146 38799
rect 55977 38855 57371 38894
rect 55977 38799 56013 38855
rect 56069 38799 56224 38855
rect 56280 38799 56435 38855
rect 56491 38799 56646 38855
rect 56702 38799 56857 38855
rect 56913 38799 57068 38855
rect 57124 38799 57279 38855
rect 57335 38799 57371 38855
rect 55977 38760 57371 38799
rect 27387 37094 27828 38760
rect 27387 37055 29146 37094
rect 27387 36999 27788 37055
rect 27844 36999 27999 37055
rect 28055 36999 28210 37055
rect 28266 36999 28421 37055
rect 28477 36999 28632 37055
rect 28688 36999 28843 37055
rect 28899 36999 29054 37055
rect 29110 36999 29146 37055
rect 27387 36960 29146 36999
rect 55977 37055 57371 37094
rect 55977 36999 56013 37055
rect 56069 36999 56224 37055
rect 56280 36999 56435 37055
rect 56491 36999 56646 37055
rect 56702 36999 56857 37055
rect 56913 36999 57068 37055
rect 57124 36999 57279 37055
rect 57335 36999 57371 37055
rect 55977 36960 57371 36999
rect 27387 35275 27828 36960
rect 36863 35881 37743 36650
rect 36863 35825 36958 35881
rect 37014 35825 37169 35881
rect 37225 35825 37381 35881
rect 37437 35825 37592 35881
rect 37648 35825 37743 35881
rect 36863 35786 37743 35825
rect 41472 35761 41694 36096
rect 38596 35532 41694 35761
rect 38596 35516 38817 35532
rect 27387 35219 27438 35275
rect 27494 35219 27562 35275
rect 27618 35219 27686 35275
rect 27742 35219 27828 35275
rect 27387 35151 27828 35219
rect 27387 35095 27438 35151
rect 27494 35095 27562 35151
rect 27618 35095 27686 35151
rect 27742 35095 27828 35151
rect 27387 35027 27828 35095
rect 27387 34971 27438 35027
rect 27494 34971 27562 35027
rect 27618 34971 27686 35027
rect 27742 34971 27828 35027
rect 27387 34903 27828 34971
rect 27387 34847 27438 34903
rect 27494 34847 27562 34903
rect 27618 34847 27686 34903
rect 27742 34847 27828 34903
rect 27387 34779 27828 34847
rect 27387 34723 27438 34779
rect 27494 34723 27562 34779
rect 27618 34723 27686 34779
rect 27742 34723 27828 34779
rect 27387 34655 27828 34723
rect 27387 34599 27438 34655
rect 27494 34599 27562 34655
rect 27618 34599 27686 34655
rect 27742 34599 27828 34655
rect 27387 33432 27828 34599
rect 27387 33380 27476 33432
rect 27528 33380 27688 33432
rect 27740 33380 27828 33432
rect 27387 33215 27828 33380
rect 31615 35287 38817 35516
rect 41850 35425 42072 35528
rect 31615 33349 31836 35287
rect 39077 35197 42072 35425
rect 39077 35171 39298 35197
rect 31970 34943 39298 35171
rect 42228 35090 42449 36096
rect 31970 33349 32192 34943
rect 39755 34861 42449 35090
rect 39755 34675 39977 34861
rect 42603 34754 42825 36085
rect 38301 34491 39977 34675
rect 37201 34446 39977 34491
rect 40106 34526 42825 34754
rect 37201 34263 38523 34446
rect 40106 34312 40328 34526
rect 42983 34419 43205 36096
rect 37201 33360 37423 34263
rect 38642 34156 40328 34312
rect 37557 34084 40328 34156
rect 40458 34190 43205 34419
rect 37557 33927 38863 34084
rect 40458 33977 40679 34190
rect 43359 34083 43580 36085
rect 45513 35842 45735 36096
rect 37557 33349 37778 33927
rect 38993 33748 40679 33977
rect 40809 33855 43580 34083
rect 44646 35614 45735 35842
rect 38993 33360 39215 33748
rect 40809 33625 41031 33855
rect 39349 33397 41031 33625
rect 44646 33576 44867 35614
rect 45891 35507 46112 36096
rect 44997 35278 46112 35507
rect 46268 35681 46490 36096
rect 46268 35453 46501 35681
rect 44997 33576 45219 35278
rect 46279 33576 46501 35453
rect 46646 35346 46868 36085
rect 46631 35117 46868 35346
rect 46631 33564 46852 35117
rect 47026 34836 47248 36085
rect 47402 35171 47623 36096
rect 47779 35507 48001 36096
rect 48157 35842 48379 36096
rect 48157 35614 50120 35842
rect 47779 35278 49769 35507
rect 47402 34943 48486 35171
rect 47026 34607 48135 34836
rect 47913 33564 48135 34607
rect 48265 33576 48486 34943
rect 49547 33576 49769 35278
rect 49898 33576 50120 35614
rect 57407 35242 57607 35254
rect 57407 35190 57419 35242
rect 57471 35190 57543 35242
rect 57595 35190 57607 35242
rect 57407 35118 57607 35190
rect 57407 35066 57419 35118
rect 57471 35066 57543 35118
rect 57595 35066 57607 35118
rect 57407 34994 57607 35066
rect 57407 34942 57419 34994
rect 57471 34942 57543 34994
rect 57595 34942 57607 34994
rect 57407 34870 57607 34942
rect 57407 34818 57419 34870
rect 57471 34818 57543 34870
rect 57595 34818 57607 34870
rect 57407 34746 57607 34818
rect 57407 34694 57419 34746
rect 57471 34694 57543 34746
rect 57595 34694 57607 34746
rect 57407 34622 57607 34694
rect 57407 34570 57419 34622
rect 57471 34570 57543 34622
rect 57595 34570 57607 34622
rect 57407 34558 57607 34570
rect 57909 34011 58351 51976
rect 57909 33955 57996 34011
rect 58052 33955 58208 34011
rect 58264 33955 58351 34011
rect 57909 33793 58351 33955
rect 57909 33737 57996 33793
rect 58052 33737 58208 33793
rect 58264 33737 58351 33793
rect 57909 33576 58351 33737
rect 57909 33520 57996 33576
rect 58052 33520 58208 33576
rect 58264 33520 58351 33576
rect 57295 33432 57736 33519
rect 57295 33380 57383 33432
rect 57435 33380 57595 33432
rect 57647 33380 57736 33432
rect 27387 33163 27476 33215
rect 27528 33163 27688 33215
rect 27740 33163 27828 33215
rect 27387 33141 27828 33163
rect 27387 33085 27474 33141
rect 27530 33085 27686 33141
rect 27742 33085 27828 33141
rect 27387 32997 27828 33085
rect 27387 32945 27476 32997
rect 27528 32945 27688 32997
rect 27740 32945 27828 32997
rect 27387 32923 27828 32945
rect 27387 32867 27474 32923
rect 27530 32867 27686 32923
rect 27742 32867 27828 32923
rect 27387 32779 27828 32867
rect 27387 32727 27476 32779
rect 27528 32727 27688 32779
rect 27740 32727 27828 32779
rect 27387 32705 27828 32727
rect 27387 32649 27474 32705
rect 27530 32649 27686 32705
rect 27742 32649 27828 32705
rect 27387 32562 27828 32649
rect 27387 32510 27476 32562
rect 27528 32510 27688 32562
rect 27740 32510 27828 32562
rect 27387 32487 27828 32510
rect 27387 32431 27474 32487
rect 27530 32431 27686 32487
rect 27742 32431 27828 32487
rect 27387 32344 27828 32431
rect 27387 32292 27476 32344
rect 27528 32292 27688 32344
rect 27740 32292 27828 32344
rect 27387 32127 27828 32292
rect 27387 32075 27476 32127
rect 27528 32075 27688 32127
rect 27740 32075 27828 32127
rect 27387 31909 27828 32075
rect 27387 31857 27476 31909
rect 27528 31857 27688 31909
rect 27740 31857 27828 31909
rect 27387 31691 27828 31857
rect 27387 31639 27476 31691
rect 27528 31639 27688 31691
rect 27740 31639 27828 31691
rect 27387 31474 27828 31639
rect 27387 31422 27476 31474
rect 27528 31422 27688 31474
rect 27740 31422 27828 31474
rect 27387 31256 27828 31422
rect 27387 31252 27476 31256
rect 27528 31252 27688 31256
rect 27740 31252 27828 31256
rect 27387 31196 27474 31252
rect 27530 31196 27686 31252
rect 27742 31196 27828 31252
rect 27387 31038 27828 31196
rect 27387 31034 27476 31038
rect 27528 31034 27688 31038
rect 27740 31034 27828 31038
rect 27387 30978 27474 31034
rect 27530 30978 27686 31034
rect 27742 30978 27828 31034
rect 27387 30821 27828 30978
rect 27387 30816 27476 30821
rect 27528 30816 27688 30821
rect 27740 30816 27828 30821
rect 27387 30760 27474 30816
rect 27530 30760 27686 30816
rect 27742 30760 27828 30816
rect 27387 30603 27828 30760
rect 27387 30598 27476 30603
rect 27528 30598 27688 30603
rect 27740 30598 27828 30603
rect 27387 30542 27474 30598
rect 27530 30542 27686 30598
rect 27742 30542 27828 30598
rect 27387 30386 27828 30542
rect 27387 30334 27476 30386
rect 27528 30334 27688 30386
rect 27740 30334 27828 30386
rect 27387 30168 27828 30334
rect 27387 30116 27476 30168
rect 27528 30116 27688 30168
rect 27740 30116 27828 30168
rect 27387 29950 27828 30116
rect 27387 29898 27476 29950
rect 27528 29898 27688 29950
rect 27740 29898 27828 29950
rect 27387 29733 27828 29898
rect 27387 29681 27476 29733
rect 27528 29681 27688 29733
rect 27740 29681 27828 29733
rect 27387 29515 27828 29681
rect 27387 29463 27476 29515
rect 27528 29463 27688 29515
rect 27740 29463 27828 29515
rect 27387 29297 27828 29463
rect 27387 29245 27476 29297
rect 27528 29245 27688 29297
rect 27740 29245 27828 29297
rect 27387 29080 27828 29245
rect 27387 29028 27476 29080
rect 27528 29028 27688 29080
rect 27740 29028 27828 29080
rect 27387 28862 27828 29028
rect 27387 28810 27476 28862
rect 27528 28810 27688 28862
rect 27740 28810 27828 28862
rect 27387 28644 27828 28810
rect 27387 28592 27476 28644
rect 27528 28592 27688 28644
rect 27740 28592 27828 28644
rect 27387 28427 27828 28592
rect 27387 28375 27476 28427
rect 27528 28375 27688 28427
rect 27740 28375 27828 28427
rect 27387 28209 27828 28375
rect 27387 28157 27476 28209
rect 27528 28157 27688 28209
rect 27740 28157 27828 28209
rect 27387 27992 27828 28157
rect 27387 27940 27476 27992
rect 27528 27940 27688 27992
rect 27740 27940 27828 27992
rect 27387 27774 27828 27940
rect 27387 27722 27476 27774
rect 27528 27722 27688 27774
rect 27740 27722 27828 27774
rect 27387 27556 27828 27722
rect 27387 27504 27476 27556
rect 27528 27504 27688 27556
rect 27740 27504 27828 27556
rect 27387 27339 27828 27504
rect 27387 27287 27476 27339
rect 27528 27287 27688 27339
rect 27740 27287 27828 27339
rect 27387 27121 27828 27287
rect 27387 27069 27476 27121
rect 27528 27069 27688 27121
rect 27740 27069 27828 27121
rect 27387 26903 27828 27069
rect 27387 26851 27476 26903
rect 27528 26851 27688 26903
rect 27740 26851 27828 26903
rect 27387 26799 27828 26851
rect 27387 26743 27474 26799
rect 27530 26743 27686 26799
rect 27742 26743 27828 26799
rect 27387 26686 27828 26743
rect 27387 26634 27476 26686
rect 27528 26634 27688 26686
rect 27740 26634 27828 26686
rect 27387 26581 27828 26634
rect 27387 26525 27474 26581
rect 27530 26525 27686 26581
rect 27742 26525 27828 26581
rect 27387 26468 27828 26525
rect 27387 26416 27476 26468
rect 27528 26416 27688 26468
rect 27740 26416 27828 26468
rect 27387 26250 27828 26416
rect 27387 26198 27476 26250
rect 27528 26198 27688 26250
rect 27740 26198 27828 26250
rect 27387 26033 27828 26198
rect 27387 25981 27476 26033
rect 27528 25981 27688 26033
rect 27740 25981 27828 26033
rect 27387 25815 27828 25981
rect 27387 25763 27476 25815
rect 27528 25763 27688 25815
rect 27740 25763 27828 25815
rect 27387 25598 27828 25763
rect 27387 25546 27476 25598
rect 27528 25546 27688 25598
rect 27740 25546 27828 25598
rect 27387 25380 27828 25546
rect 27387 25328 27476 25380
rect 27528 25328 27688 25380
rect 27740 25328 27828 25380
rect 27387 25162 27828 25328
rect 27387 25110 27476 25162
rect 27528 25110 27688 25162
rect 27740 25110 27828 25162
rect 27387 25028 27828 25110
rect 27387 24972 27474 25028
rect 27530 24972 27686 25028
rect 27742 24972 27828 25028
rect 27387 24945 27828 24972
rect 27387 24893 27476 24945
rect 27528 24893 27688 24945
rect 27740 24893 27828 24945
rect 27387 24810 27828 24893
rect 27387 24754 27474 24810
rect 27530 24754 27686 24810
rect 27742 24754 27828 24810
rect 27387 24727 27828 24754
rect 27387 24675 27476 24727
rect 27528 24675 27688 24727
rect 27740 24675 27828 24727
rect 27387 24509 27828 24675
rect 27387 24457 27476 24509
rect 27528 24457 27688 24509
rect 27740 24457 27828 24509
rect 27387 24292 27828 24457
rect 27387 24240 27476 24292
rect 27528 24240 27688 24292
rect 27740 24240 27828 24292
rect 27387 24074 27828 24240
rect 27387 24022 27476 24074
rect 27528 24022 27688 24074
rect 27740 24022 27828 24074
rect 27387 23857 27828 24022
rect 27387 23805 27476 23857
rect 27528 23805 27688 23857
rect 27740 23805 27828 23857
rect 27387 23639 27828 23805
rect 27387 23587 27476 23639
rect 27528 23587 27688 23639
rect 27740 23587 27828 23639
rect 27387 23421 27828 23587
rect 27387 23369 27476 23421
rect 27528 23369 27688 23421
rect 27740 23369 27828 23421
rect 27387 23204 27828 23369
rect 27387 23152 27476 23204
rect 27528 23152 27688 23204
rect 27740 23152 27828 23204
rect 27387 22986 27828 23152
rect 27387 22936 27476 22986
rect 27528 22936 27688 22986
rect 27387 22048 27475 22936
rect 27740 22934 27828 22986
rect 27739 22768 27828 22934
rect 27740 22716 27828 22768
rect 27739 22551 27828 22716
rect 27740 22499 27828 22551
rect 27739 22333 27828 22499
rect 27740 22281 27828 22333
rect 27739 22115 27828 22281
rect 27740 22063 27828 22115
rect 27739 22048 27828 22063
rect 27387 21898 27828 22048
rect 27387 21846 27476 21898
rect 27528 21846 27688 21898
rect 27740 21846 27828 21898
rect 27387 21680 27828 21846
rect 27387 21628 27476 21680
rect 27528 21628 27688 21680
rect 27740 21628 27828 21680
rect 27387 21463 27828 21628
rect 27387 21411 27476 21463
rect 27528 21411 27688 21463
rect 27740 21411 27828 21463
rect 27387 21245 27828 21411
rect 27387 21193 27476 21245
rect 27528 21193 27688 21245
rect 27740 21193 27828 21245
rect 27387 21027 27828 21193
rect 27387 20975 27476 21027
rect 27528 20975 27688 21027
rect 27740 20975 27828 21027
rect 27387 20810 27828 20975
rect 27387 20758 27476 20810
rect 27528 20758 27688 20810
rect 27740 20758 27828 20810
rect 27387 20592 27828 20758
rect 27387 20540 27476 20592
rect 27528 20540 27688 20592
rect 27740 20540 27828 20592
rect 27387 20374 27828 20540
rect 27387 20322 27476 20374
rect 27528 20322 27688 20374
rect 27740 20322 27828 20374
rect 27387 20157 27828 20322
rect 27387 20105 27476 20157
rect 27528 20105 27688 20157
rect 27740 20105 27828 20157
rect 27387 19939 27828 20105
rect 27387 19887 27476 19939
rect 27528 19887 27688 19939
rect 27740 19887 27828 19939
rect 27387 19722 27828 19887
rect 27387 19670 27476 19722
rect 27528 19670 27688 19722
rect 27740 19670 27828 19722
rect 27387 19504 27828 19670
rect 27387 19452 27476 19504
rect 27528 19452 27688 19504
rect 27740 19452 27828 19504
rect 27387 19286 27828 19452
rect 27387 19234 27476 19286
rect 27528 19234 27688 19286
rect 27740 19234 27828 19286
rect 27387 19068 27828 19234
rect 27387 19016 27476 19068
rect 27528 19016 27688 19068
rect 27740 19016 27828 19068
rect 27387 18851 27828 19016
rect 27387 18799 27476 18851
rect 27528 18799 27688 18851
rect 27740 18799 27828 18851
rect 27387 18633 27828 18799
rect 27387 18581 27476 18633
rect 27528 18581 27688 18633
rect 27740 18581 27828 18633
rect 27387 18416 27828 18581
rect 27387 18364 27476 18416
rect 27528 18364 27688 18416
rect 27740 18364 27828 18416
rect 27387 18198 27828 18364
rect 27387 18146 27476 18198
rect 27528 18146 27688 18198
rect 27740 18146 27828 18198
rect 27387 17980 27828 18146
rect 27387 17928 27476 17980
rect 27528 17928 27688 17980
rect 27740 17928 27828 17980
rect 27387 17763 27828 17928
rect 27387 17711 27476 17763
rect 27528 17711 27688 17763
rect 27740 17711 27828 17763
rect 27387 17545 27828 17711
rect 27387 17493 27476 17545
rect 27528 17493 27688 17545
rect 27740 17493 27828 17545
rect 27387 17327 27828 17493
rect 27387 17275 27476 17327
rect 27528 17275 27688 17327
rect 27740 17275 27828 17327
rect 27387 17110 27828 17275
rect 27387 17058 27476 17110
rect 27528 17058 27688 17110
rect 27740 17058 27828 17110
rect 27387 16892 27828 17058
rect 27387 16840 27476 16892
rect 27528 16840 27688 16892
rect 27740 16840 27828 16892
rect 27387 16675 27828 16840
rect 27387 16623 27476 16675
rect 27528 16623 27688 16675
rect 27740 16623 27828 16675
rect 27387 16470 27828 16623
rect 27387 16414 27474 16470
rect 27530 16414 27686 16470
rect 27742 16414 27828 16470
rect 27387 16405 27476 16414
rect 27528 16405 27688 16414
rect 27740 16405 27828 16414
rect 27387 16253 27828 16405
rect 27387 16197 27474 16253
rect 27530 16197 27686 16253
rect 27742 16197 27828 16253
rect 27387 16187 27476 16197
rect 27528 16187 27688 16197
rect 27740 16187 27828 16197
rect 27387 16035 27828 16187
rect 27387 15979 27474 16035
rect 27530 15979 27686 16035
rect 27742 15979 27828 16035
rect 27387 15970 27476 15979
rect 27528 15970 27688 15979
rect 27740 15970 27828 15979
rect 27387 15818 27828 15970
rect 27387 15762 27474 15818
rect 27530 15762 27686 15818
rect 27742 15762 27828 15818
rect 27387 15752 27476 15762
rect 27528 15752 27688 15762
rect 27740 15752 27828 15762
rect 27387 15600 27828 15752
rect 27387 15544 27474 15600
rect 27530 15544 27686 15600
rect 27742 15544 27828 15600
rect 27387 15534 27476 15544
rect 27528 15534 27688 15544
rect 27740 15534 27828 15544
rect 27387 15382 27828 15534
rect 27387 15326 27474 15382
rect 27530 15326 27686 15382
rect 27742 15326 27828 15382
rect 27387 15317 27476 15326
rect 27528 15317 27688 15326
rect 27740 15317 27828 15326
rect 27387 15164 27828 15317
rect 27387 15108 27474 15164
rect 27530 15108 27686 15164
rect 27742 15108 27828 15164
rect 27387 15099 27476 15108
rect 27528 15099 27688 15108
rect 27740 15099 27828 15108
rect 27387 14947 27828 15099
rect 27387 14891 27474 14947
rect 27530 14891 27686 14947
rect 27742 14891 27828 14947
rect 27387 14881 27476 14891
rect 27528 14881 27688 14891
rect 27740 14881 27828 14891
rect 27387 14729 27828 14881
rect 27387 14673 27474 14729
rect 27530 14673 27686 14729
rect 27742 14673 27828 14729
rect 27387 14664 27476 14673
rect 27528 14664 27688 14673
rect 27740 14664 27828 14673
rect 27387 14512 27828 14664
rect 27387 14456 27474 14512
rect 27530 14456 27686 14512
rect 27742 14456 27828 14512
rect 27387 14446 27476 14456
rect 27528 14446 27688 14456
rect 27740 14446 27828 14456
rect 27387 14281 27828 14446
rect 27387 14231 27476 14281
rect 27528 14231 27688 14281
rect 27740 14231 27828 14281
rect 27387 14175 27474 14231
rect 27530 14175 27686 14231
rect 27742 14175 27828 14231
rect 27387 14063 27828 14175
rect 27387 14014 27476 14063
rect 27528 14014 27688 14063
rect 27740 14014 27828 14063
rect 27387 13958 27474 14014
rect 27530 13958 27686 14014
rect 27742 13958 27828 14014
rect 27387 13845 27828 13958
rect 27387 13796 27476 13845
rect 27528 13796 27688 13845
rect 27740 13796 27828 13845
rect 27387 13740 27474 13796
rect 27530 13740 27686 13796
rect 27742 13740 27828 13796
rect 27387 13628 27828 13740
rect 27387 13578 27476 13628
rect 27528 13578 27688 13628
rect 27740 13578 27828 13628
rect 27387 13522 27474 13578
rect 27530 13522 27686 13578
rect 27742 13522 27828 13578
rect 27387 13410 27828 13522
rect 27387 13361 27476 13410
rect 27528 13361 27688 13410
rect 27740 13361 27828 13410
rect 27387 13305 27474 13361
rect 27530 13305 27686 13361
rect 27742 13305 27828 13361
rect 27387 13192 27828 13305
rect 27387 13140 27476 13192
rect 27528 13140 27688 13192
rect 27740 13140 27828 13192
rect 27387 12975 27828 13140
rect 27387 12923 27476 12975
rect 27528 12923 27688 12975
rect 27740 12923 27828 12975
rect 27387 12757 27828 12923
rect 27387 12705 27476 12757
rect 27528 12705 27688 12757
rect 27740 12705 27828 12757
rect 27387 12540 27828 12705
rect 27387 12488 27476 12540
rect 27528 12488 27688 12540
rect 27740 12488 27828 12540
rect 27387 12322 27828 12488
rect 27387 12270 27476 12322
rect 27528 12270 27688 12322
rect 27740 12270 27828 12322
rect 27387 12104 27828 12270
rect 27387 12052 27476 12104
rect 27528 12052 27688 12104
rect 27740 12052 27828 12104
rect 27387 11887 27828 12052
rect 27387 11835 27476 11887
rect 27528 11835 27688 11887
rect 27740 11835 27828 11887
rect 27387 11669 27828 11835
rect 27387 11617 27476 11669
rect 27528 11617 27688 11669
rect 27740 11617 27828 11669
rect 27387 11451 27828 11617
rect 27387 11406 27476 11451
rect 27528 11406 27688 11451
rect 27740 11406 27828 11451
rect 27387 11350 27474 11406
rect 27530 11350 27686 11406
rect 27742 11350 27828 11406
rect 27387 11234 27828 11350
rect 27387 11189 27476 11234
rect 27528 11189 27688 11234
rect 27740 11189 27828 11234
rect 27387 11133 27474 11189
rect 27530 11133 27686 11189
rect 27742 11133 27828 11189
rect 27387 11016 27828 11133
rect 27387 10971 27476 11016
rect 27528 10971 27688 11016
rect 27740 10971 27828 11016
rect 27387 10915 27474 10971
rect 27530 10915 27686 10971
rect 27742 10915 27828 10971
rect 27387 10798 27828 10915
rect 27387 10753 27476 10798
rect 27528 10753 27688 10798
rect 27740 10753 27828 10798
rect 27387 10697 27474 10753
rect 27530 10697 27686 10753
rect 27742 10697 27828 10753
rect 27387 10581 27828 10697
rect 27387 10535 27476 10581
rect 27528 10535 27688 10581
rect 27740 10535 27828 10581
rect 27387 10479 27474 10535
rect 27530 10479 27686 10535
rect 27742 10479 27828 10535
rect 27387 10363 27828 10479
rect 27387 10318 27476 10363
rect 27528 10318 27688 10363
rect 27740 10318 27828 10363
rect 27387 10262 27474 10318
rect 27530 10262 27686 10318
rect 27742 10262 27828 10318
rect 27387 10146 27828 10262
rect 27387 10094 27476 10146
rect 27528 10094 27688 10146
rect 27740 10094 27828 10146
rect 27387 9928 27828 10094
rect 57295 33215 57736 33380
rect 57295 33163 57383 33215
rect 57435 33163 57595 33215
rect 57647 33163 57736 33215
rect 57295 33141 57736 33163
rect 57295 33085 57381 33141
rect 57437 33085 57593 33141
rect 57649 33085 57736 33141
rect 57295 32997 57736 33085
rect 57295 32945 57383 32997
rect 57435 32945 57595 32997
rect 57647 32945 57736 32997
rect 57295 32923 57736 32945
rect 57295 32867 57381 32923
rect 57437 32867 57593 32923
rect 57649 32867 57736 32923
rect 57295 32779 57736 32867
rect 57295 32727 57383 32779
rect 57435 32727 57595 32779
rect 57647 32727 57736 32779
rect 57295 32705 57736 32727
rect 57295 32649 57381 32705
rect 57437 32649 57593 32705
rect 57649 32649 57736 32705
rect 57295 32562 57736 32649
rect 57295 32510 57383 32562
rect 57435 32510 57595 32562
rect 57647 32510 57736 32562
rect 57295 32487 57736 32510
rect 57295 32431 57381 32487
rect 57437 32431 57593 32487
rect 57649 32431 57736 32487
rect 57295 32344 57736 32431
rect 57295 32292 57383 32344
rect 57435 32292 57595 32344
rect 57647 32292 57736 32344
rect 57295 32127 57736 32292
rect 57295 32075 57383 32127
rect 57435 32075 57595 32127
rect 57647 32075 57736 32127
rect 57295 31909 57736 32075
rect 57295 31857 57383 31909
rect 57435 31857 57595 31909
rect 57647 31857 57736 31909
rect 57295 31691 57736 31857
rect 57295 31639 57383 31691
rect 57435 31639 57595 31691
rect 57647 31639 57736 31691
rect 57295 31474 57736 31639
rect 57295 31422 57383 31474
rect 57435 31422 57595 31474
rect 57647 31422 57736 31474
rect 57295 31256 57736 31422
rect 57295 31252 57383 31256
rect 57435 31252 57595 31256
rect 57647 31252 57736 31256
rect 57295 31196 57381 31252
rect 57437 31196 57593 31252
rect 57649 31196 57736 31252
rect 57295 31038 57736 31196
rect 57295 31034 57383 31038
rect 57435 31034 57595 31038
rect 57647 31034 57736 31038
rect 57295 30978 57381 31034
rect 57437 30978 57593 31034
rect 57649 30978 57736 31034
rect 57295 30821 57736 30978
rect 57295 30816 57383 30821
rect 57435 30816 57595 30821
rect 57647 30816 57736 30821
rect 57295 30760 57381 30816
rect 57437 30760 57593 30816
rect 57649 30760 57736 30816
rect 57295 30603 57736 30760
rect 57295 30598 57383 30603
rect 57435 30598 57595 30603
rect 57647 30598 57736 30603
rect 57295 30542 57381 30598
rect 57437 30542 57593 30598
rect 57649 30542 57736 30598
rect 57295 30386 57736 30542
rect 57295 30334 57383 30386
rect 57435 30334 57595 30386
rect 57647 30334 57736 30386
rect 57295 30168 57736 30334
rect 57295 30116 57383 30168
rect 57435 30116 57595 30168
rect 57647 30116 57736 30168
rect 57295 29950 57736 30116
rect 57295 29898 57383 29950
rect 57435 29898 57595 29950
rect 57647 29898 57736 29950
rect 57295 29733 57736 29898
rect 57295 29681 57383 29733
rect 57435 29681 57595 29733
rect 57647 29681 57736 29733
rect 57295 29515 57736 29681
rect 57295 29463 57383 29515
rect 57435 29463 57595 29515
rect 57647 29463 57736 29515
rect 57295 29297 57736 29463
rect 57295 29245 57383 29297
rect 57435 29245 57595 29297
rect 57647 29245 57736 29297
rect 57295 29080 57736 29245
rect 57295 29028 57383 29080
rect 57435 29028 57595 29080
rect 57647 29028 57736 29080
rect 57295 28862 57736 29028
rect 57295 28810 57383 28862
rect 57435 28810 57595 28862
rect 57647 28810 57736 28862
rect 57295 28644 57736 28810
rect 57295 28592 57383 28644
rect 57435 28592 57595 28644
rect 57647 28592 57736 28644
rect 57295 28427 57736 28592
rect 57295 28375 57383 28427
rect 57435 28375 57595 28427
rect 57647 28375 57736 28427
rect 57295 28209 57736 28375
rect 57295 28157 57383 28209
rect 57435 28157 57595 28209
rect 57647 28157 57736 28209
rect 57295 27992 57736 28157
rect 57295 27940 57383 27992
rect 57435 27940 57595 27992
rect 57647 27940 57736 27992
rect 57295 27774 57736 27940
rect 57295 27722 57383 27774
rect 57435 27722 57595 27774
rect 57647 27722 57736 27774
rect 57295 27556 57736 27722
rect 57295 27504 57383 27556
rect 57435 27504 57595 27556
rect 57647 27504 57736 27556
rect 57295 27339 57736 27504
rect 57295 27287 57383 27339
rect 57435 27287 57595 27339
rect 57647 27287 57736 27339
rect 57295 27121 57736 27287
rect 57295 27069 57383 27121
rect 57435 27069 57595 27121
rect 57647 27069 57736 27121
rect 57295 26903 57736 27069
rect 57295 26851 57383 26903
rect 57435 26851 57595 26903
rect 57647 26851 57736 26903
rect 57295 26799 57736 26851
rect 57295 26743 57381 26799
rect 57437 26743 57593 26799
rect 57649 26743 57736 26799
rect 57295 26686 57736 26743
rect 57295 26634 57383 26686
rect 57435 26634 57595 26686
rect 57647 26634 57736 26686
rect 57295 26581 57736 26634
rect 57295 26525 57381 26581
rect 57437 26525 57593 26581
rect 57649 26525 57736 26581
rect 57295 26468 57736 26525
rect 57295 26416 57383 26468
rect 57435 26416 57595 26468
rect 57647 26416 57736 26468
rect 57295 26250 57736 26416
rect 57295 26198 57383 26250
rect 57435 26198 57595 26250
rect 57647 26198 57736 26250
rect 57295 26033 57736 26198
rect 57295 25981 57383 26033
rect 57435 25981 57595 26033
rect 57647 25981 57736 26033
rect 57295 25815 57736 25981
rect 57295 25763 57383 25815
rect 57435 25763 57595 25815
rect 57647 25763 57736 25815
rect 57295 25598 57736 25763
rect 57295 25546 57383 25598
rect 57435 25546 57595 25598
rect 57647 25546 57736 25598
rect 57295 25380 57736 25546
rect 57295 25328 57383 25380
rect 57435 25328 57595 25380
rect 57647 25328 57736 25380
rect 57295 25162 57736 25328
rect 57295 25110 57383 25162
rect 57435 25110 57595 25162
rect 57647 25110 57736 25162
rect 57295 24945 57736 25110
rect 57295 24893 57383 24945
rect 57435 24893 57595 24945
rect 57647 24893 57736 24945
rect 57295 24727 57736 24893
rect 57295 24675 57383 24727
rect 57435 24675 57595 24727
rect 57647 24675 57736 24727
rect 57295 24509 57736 24675
rect 57295 24457 57383 24509
rect 57435 24457 57595 24509
rect 57647 24457 57736 24509
rect 57295 24292 57736 24457
rect 57295 24240 57383 24292
rect 57435 24240 57595 24292
rect 57647 24240 57736 24292
rect 57295 24074 57736 24240
rect 57295 24022 57383 24074
rect 57435 24022 57595 24074
rect 57647 24022 57736 24074
rect 57295 23857 57736 24022
rect 57295 23805 57383 23857
rect 57435 23805 57595 23857
rect 57647 23805 57736 23857
rect 57295 23639 57736 23805
rect 57295 23587 57383 23639
rect 57435 23587 57595 23639
rect 57647 23587 57736 23639
rect 57295 23421 57736 23587
rect 57295 23369 57383 23421
rect 57435 23369 57595 23421
rect 57647 23369 57736 23421
rect 57295 23204 57736 23369
rect 57295 23152 57383 23204
rect 57435 23152 57595 23204
rect 57647 23152 57736 23204
rect 57295 22986 57736 23152
rect 57295 22934 57383 22986
rect 57435 22934 57595 22986
rect 57647 22934 57736 22986
rect 57295 22923 57736 22934
rect 57295 22035 57363 22923
rect 57627 22768 57736 22923
rect 57647 22716 57736 22768
rect 57627 22551 57736 22716
rect 57647 22499 57736 22551
rect 57627 22333 57736 22499
rect 57647 22281 57736 22333
rect 57627 22115 57736 22281
rect 57647 22063 57736 22115
rect 57627 22035 57736 22063
rect 57295 21898 57736 22035
rect 57295 21846 57383 21898
rect 57435 21846 57595 21898
rect 57647 21846 57736 21898
rect 57295 21680 57736 21846
rect 57295 21628 57383 21680
rect 57435 21628 57595 21680
rect 57647 21628 57736 21680
rect 57295 21463 57736 21628
rect 57295 21411 57383 21463
rect 57435 21411 57595 21463
rect 57647 21411 57736 21463
rect 57295 21245 57736 21411
rect 57295 21193 57383 21245
rect 57435 21193 57595 21245
rect 57647 21193 57736 21245
rect 57295 21027 57736 21193
rect 57295 20975 57383 21027
rect 57435 20975 57595 21027
rect 57647 20975 57736 21027
rect 57295 20810 57736 20975
rect 57295 20758 57383 20810
rect 57435 20758 57595 20810
rect 57647 20758 57736 20810
rect 57295 20592 57736 20758
rect 57295 20540 57383 20592
rect 57435 20540 57595 20592
rect 57647 20540 57736 20592
rect 57295 20374 57736 20540
rect 57295 20322 57383 20374
rect 57435 20322 57595 20374
rect 57647 20322 57736 20374
rect 57295 20157 57736 20322
rect 57295 20105 57383 20157
rect 57435 20105 57595 20157
rect 57647 20105 57736 20157
rect 57295 19939 57736 20105
rect 57295 19887 57383 19939
rect 57435 19887 57595 19939
rect 57647 19887 57736 19939
rect 57295 19722 57736 19887
rect 57295 19670 57383 19722
rect 57435 19670 57595 19722
rect 57647 19670 57736 19722
rect 57295 19504 57736 19670
rect 57295 19452 57383 19504
rect 57435 19452 57595 19504
rect 57647 19452 57736 19504
rect 57295 19286 57736 19452
rect 57295 19234 57383 19286
rect 57435 19234 57595 19286
rect 57647 19234 57736 19286
rect 57295 19068 57736 19234
rect 57295 19016 57383 19068
rect 57435 19016 57595 19068
rect 57647 19016 57736 19068
rect 57295 18851 57736 19016
rect 57295 18799 57383 18851
rect 57435 18799 57595 18851
rect 57647 18799 57736 18851
rect 57295 18633 57736 18799
rect 57295 18581 57383 18633
rect 57435 18581 57595 18633
rect 57647 18581 57736 18633
rect 57295 18416 57736 18581
rect 57295 18364 57383 18416
rect 57435 18364 57595 18416
rect 57647 18364 57736 18416
rect 57295 18198 57736 18364
rect 57295 18146 57383 18198
rect 57435 18146 57595 18198
rect 57647 18146 57736 18198
rect 57295 17980 57736 18146
rect 57295 17928 57383 17980
rect 57435 17928 57595 17980
rect 57647 17928 57736 17980
rect 57295 17763 57736 17928
rect 57295 17711 57383 17763
rect 57435 17711 57595 17763
rect 57647 17711 57736 17763
rect 57295 17545 57736 17711
rect 57295 17493 57383 17545
rect 57435 17493 57595 17545
rect 57647 17493 57736 17545
rect 57295 17327 57736 17493
rect 57295 17275 57383 17327
rect 57435 17275 57595 17327
rect 57647 17275 57736 17327
rect 57295 17110 57736 17275
rect 57295 17058 57383 17110
rect 57435 17058 57595 17110
rect 57647 17058 57736 17110
rect 57295 16892 57736 17058
rect 57295 16840 57383 16892
rect 57435 16840 57595 16892
rect 57647 16840 57736 16892
rect 57295 16678 57736 16840
rect 57295 16622 57381 16678
rect 57437 16622 57593 16678
rect 57649 16622 57736 16678
rect 57295 16461 57736 16622
rect 57295 16405 57381 16461
rect 57437 16405 57593 16461
rect 57649 16405 57736 16461
rect 57295 16243 57736 16405
rect 57295 16187 57381 16243
rect 57437 16187 57593 16243
rect 57649 16187 57736 16243
rect 57295 16026 57736 16187
rect 57295 15970 57381 16026
rect 57437 15970 57593 16026
rect 57649 15970 57736 16026
rect 57295 15808 57736 15970
rect 57295 15752 57381 15808
rect 57437 15752 57593 15808
rect 57649 15752 57736 15808
rect 57295 15590 57736 15752
rect 57295 15534 57381 15590
rect 57437 15534 57593 15590
rect 57649 15534 57736 15590
rect 57295 15372 57736 15534
rect 57295 15316 57381 15372
rect 57437 15316 57593 15372
rect 57649 15316 57736 15372
rect 57295 15155 57736 15316
rect 57295 15099 57381 15155
rect 57437 15099 57593 15155
rect 57649 15099 57736 15155
rect 57295 14937 57736 15099
rect 57295 14881 57381 14937
rect 57437 14881 57593 14937
rect 57649 14881 57736 14937
rect 57295 14720 57736 14881
rect 57295 14664 57381 14720
rect 57437 14664 57593 14720
rect 57649 14664 57736 14720
rect 57295 14498 57736 14664
rect 57295 14446 57383 14498
rect 57435 14446 57595 14498
rect 57647 14446 57736 14498
rect 57295 14281 57736 14446
rect 57295 14229 57383 14281
rect 57435 14229 57595 14281
rect 57647 14229 57736 14281
rect 57295 14063 57736 14229
rect 57295 14011 57383 14063
rect 57435 14011 57595 14063
rect 57647 14011 57736 14063
rect 57295 13845 57736 14011
rect 57295 13793 57383 13845
rect 57435 13793 57595 13845
rect 57647 13793 57736 13845
rect 57295 13628 57736 13793
rect 57295 13576 57383 13628
rect 57435 13576 57595 13628
rect 57647 13576 57736 13628
rect 57295 13410 57736 13576
rect 57295 13358 57383 13410
rect 57435 13358 57595 13410
rect 57647 13358 57736 13410
rect 57295 13192 57736 13358
rect 57295 13140 57383 13192
rect 57435 13140 57595 13192
rect 57647 13140 57736 13192
rect 57295 12975 57736 13140
rect 57295 12923 57383 12975
rect 57435 12923 57595 12975
rect 57647 12923 57736 12975
rect 57295 12757 57736 12923
rect 57295 12705 57383 12757
rect 57435 12705 57595 12757
rect 57647 12705 57736 12757
rect 57295 12540 57736 12705
rect 57295 12488 57383 12540
rect 57435 12488 57595 12540
rect 57647 12488 57736 12540
rect 57295 12322 57736 12488
rect 57295 12270 57383 12322
rect 57435 12270 57595 12322
rect 57647 12270 57736 12322
rect 57295 12104 57736 12270
rect 57295 12052 57383 12104
rect 57435 12052 57595 12104
rect 57647 12052 57736 12104
rect 57295 11887 57736 12052
rect 57295 11835 57383 11887
rect 57435 11835 57595 11887
rect 57647 11835 57736 11887
rect 57295 11669 57736 11835
rect 57295 11617 57383 11669
rect 57435 11617 57595 11669
rect 57647 11617 57736 11669
rect 57295 11451 57736 11617
rect 57295 11406 57383 11451
rect 57435 11406 57595 11451
rect 57647 11406 57736 11451
rect 57295 11350 57381 11406
rect 57437 11350 57593 11406
rect 57649 11350 57736 11406
rect 57295 11234 57736 11350
rect 57295 11189 57383 11234
rect 57435 11189 57595 11234
rect 57647 11189 57736 11234
rect 57295 11133 57381 11189
rect 57437 11133 57593 11189
rect 57649 11133 57736 11189
rect 57295 11016 57736 11133
rect 57295 10971 57383 11016
rect 57435 10971 57595 11016
rect 57647 10971 57736 11016
rect 57295 10915 57381 10971
rect 57437 10915 57593 10971
rect 57649 10915 57736 10971
rect 57295 10798 57736 10915
rect 57295 10753 57383 10798
rect 57435 10753 57595 10798
rect 57647 10753 57736 10798
rect 57295 10697 57381 10753
rect 57437 10697 57593 10753
rect 57649 10697 57736 10753
rect 57295 10581 57736 10697
rect 57295 10535 57383 10581
rect 57435 10535 57595 10581
rect 57647 10535 57736 10581
rect 57295 10479 57381 10535
rect 57437 10479 57593 10535
rect 57649 10479 57736 10535
rect 57295 10363 57736 10479
rect 57295 10318 57383 10363
rect 57435 10318 57595 10363
rect 57647 10318 57736 10363
rect 57295 10262 57381 10318
rect 57437 10262 57593 10318
rect 57649 10262 57736 10318
rect 57295 10146 57736 10262
rect 57295 10094 57383 10146
rect 57435 10094 57595 10146
rect 57647 10094 57736 10146
rect 27387 9876 27476 9928
rect 27528 9876 27688 9928
rect 27740 9876 27828 9928
rect 27387 9710 27828 9876
rect 51756 9971 51832 9981
rect 51756 9811 51766 9971
rect 51822 9811 51832 9971
rect 51756 9801 51832 9811
rect 57295 9928 57736 10094
rect 57295 9876 57383 9928
rect 57435 9876 57595 9928
rect 57647 9876 57736 9928
rect 27387 9658 27476 9710
rect 27528 9658 27688 9710
rect 27740 9658 27828 9710
rect 27387 9493 27828 9658
rect 27387 9441 27476 9493
rect 27528 9441 27688 9493
rect 27740 9441 27828 9493
rect 27387 9275 27828 9441
rect 27387 9223 27476 9275
rect 27528 9223 27688 9275
rect 27740 9223 27828 9275
rect 27387 9057 27828 9223
rect 27387 9005 27476 9057
rect 27528 9005 27688 9057
rect 27740 9005 27828 9057
rect 27387 8840 27828 9005
rect 49896 8956 50076 8966
rect 49896 8900 49906 8956
rect 50066 8900 50076 8956
rect 49896 8890 50076 8900
rect 27387 8788 27476 8840
rect 27528 8788 27688 8840
rect 27740 8788 27828 8840
rect 27387 8622 27828 8788
rect 27387 8570 27476 8622
rect 27528 8570 27688 8622
rect 27740 8570 27828 8622
rect 27387 8404 27828 8570
rect 27387 8352 27476 8404
rect 27528 8352 27688 8404
rect 27740 8352 27828 8404
rect 27387 8187 27828 8352
rect 27387 8135 27476 8187
rect 27528 8135 27688 8187
rect 27740 8135 27828 8187
rect 27387 7969 27828 8135
rect 27387 7917 27476 7969
rect 27528 7917 27688 7969
rect 27740 7917 27828 7969
rect 27387 7752 27828 7917
rect 27387 7700 27476 7752
rect 27528 7700 27688 7752
rect 27740 7700 27828 7752
rect 27387 7535 27828 7700
rect 27387 7479 27474 7535
rect 27530 7479 27686 7535
rect 27742 7479 27828 7535
rect 27387 7317 27828 7479
rect 27387 7261 27474 7317
rect 27530 7261 27686 7317
rect 27742 7261 27828 7317
rect 27387 7099 27828 7261
rect 27387 7043 27474 7099
rect 27530 7043 27686 7099
rect 27742 7043 27828 7099
rect 27387 6881 27828 7043
rect 27387 6829 27476 6881
rect 27528 6829 27688 6881
rect 27740 6829 27828 6881
rect 27387 6663 27828 6829
rect 27387 6611 27476 6663
rect 27528 6611 27688 6663
rect 27740 6611 27828 6663
rect 27387 6446 27828 6611
rect 27387 6394 27476 6446
rect 27528 6394 27688 6446
rect 27740 6394 27828 6446
rect 27387 6228 27828 6394
rect 28237 6836 28999 6874
rect 28237 6780 28273 6836
rect 28329 6780 28484 6836
rect 28540 6780 28696 6836
rect 28752 6780 28907 6836
rect 28963 6780 28999 6836
rect 28237 6618 28999 6780
rect 28237 6562 28273 6618
rect 28329 6562 28484 6618
rect 28540 6562 28696 6618
rect 28752 6562 28907 6618
rect 28963 6562 28999 6618
rect 28237 6400 28999 6562
rect 28237 6344 28273 6400
rect 28329 6344 28484 6400
rect 28540 6344 28696 6400
rect 28752 6344 28907 6400
rect 28963 6344 28999 6400
rect 49958 6361 50014 8890
rect 28237 6306 28999 6344
rect 49896 6349 50076 6361
rect 49896 6297 49908 6349
rect 50064 6297 50076 6349
rect 49896 6285 50076 6297
rect 27387 6176 27476 6228
rect 27528 6176 27688 6228
rect 27740 6176 27828 6228
rect 27387 6120 27828 6176
rect 27387 6064 27474 6120
rect 27530 6064 27686 6120
rect 27742 6064 27828 6120
rect 27387 6011 27828 6064
rect 27387 5959 27476 6011
rect 27528 5959 27688 6011
rect 27740 5959 27828 6011
rect 27387 5902 27828 5959
rect 27387 5846 27474 5902
rect 27530 5846 27686 5902
rect 27742 5846 27828 5902
rect 27387 5793 27828 5846
rect 27387 5741 27476 5793
rect 27528 5741 27688 5793
rect 27740 5741 27828 5793
rect 27387 5575 27828 5741
rect 27387 5523 27476 5575
rect 27528 5523 27688 5575
rect 27740 5523 27828 5575
rect 27387 5358 27828 5523
rect 27387 5306 27476 5358
rect 27528 5306 27688 5358
rect 27740 5306 27828 5358
rect 1864 5024 2509 5135
rect 11727 5073 11783 5140
rect 1864 0 2088 5024
rect 3263 5001 3357 5062
rect 11617 5017 11783 5073
rect 3263 4880 3604 5001
rect 2539 1689 2763 1701
rect 2539 1637 2574 1689
rect 2730 1637 2763 1689
rect 2539 0 2763 1637
rect 3380 0 3604 4880
rect 11617 1701 11673 5017
rect 12575 4740 12631 5185
rect 12290 4684 12631 4740
rect 13253 4740 13309 5185
rect 14101 5073 14157 5140
rect 14101 5017 14267 5073
rect 13253 4684 13594 4740
rect 12290 1701 12346 4684
rect 13538 1701 13594 4684
rect 14211 1701 14267 5017
rect 22527 5001 22621 5062
rect 23375 5024 24019 5135
rect 22279 4880 22621 5001
rect 11533 0 11757 1701
rect 12206 0 12430 1701
rect 12604 1689 12828 1701
rect 12604 1637 12639 1689
rect 12795 1637 12828 1689
rect 12604 0 12828 1637
rect 13054 1689 13278 1701
rect 13054 1637 13089 1689
rect 13245 1637 13278 1689
rect 13054 0 13278 1637
rect 13454 0 13678 1701
rect 14127 0 14351 1701
rect 22279 0 22503 4880
rect 23404 1689 23628 1701
rect 23404 1637 23439 1689
rect 23595 1637 23628 1689
rect 23404 0 23628 1637
rect 23795 0 24019 5024
rect 26823 4587 27163 4628
rect 26823 4535 26861 4587
rect 26913 4535 27073 4587
rect 27125 4535 27163 4587
rect 26823 4528 27163 4535
rect 26823 4472 26859 4528
rect 26915 4472 27071 4528
rect 27127 4472 27163 4528
rect 26823 4370 27163 4472
rect 26823 4318 26861 4370
rect 26913 4318 27073 4370
rect 27125 4318 27163 4370
rect 26823 4310 27163 4318
rect 26823 4254 26859 4310
rect 26915 4254 27071 4310
rect 27127 4254 27163 4310
rect 26823 4152 27163 4254
rect 26823 4100 26861 4152
rect 26913 4100 27073 4152
rect 27125 4100 27163 4152
rect 26823 3934 27163 4100
rect 26823 3882 26861 3934
rect 26913 3882 27073 3934
rect 27125 3882 27163 3934
rect 26823 3717 27163 3882
rect 26823 3665 26861 3717
rect 26913 3665 27073 3717
rect 27125 3665 27163 3717
rect 26823 3624 27163 3665
rect 27387 4587 27828 5306
rect 51766 5211 51822 9801
rect 57295 9710 57736 9876
rect 57295 9658 57383 9710
rect 57435 9658 57595 9710
rect 57647 9658 57736 9710
rect 57295 9493 57736 9658
rect 57295 9441 57383 9493
rect 57435 9441 57595 9493
rect 57647 9441 57736 9493
rect 57295 9275 57736 9441
rect 57295 9223 57383 9275
rect 57435 9223 57595 9275
rect 57647 9223 57736 9275
rect 57295 9057 57736 9223
rect 57295 9005 57383 9057
rect 57435 9005 57595 9057
rect 57647 9005 57736 9057
rect 57295 8840 57736 9005
rect 57295 8837 57383 8840
rect 57435 8837 57595 8840
rect 57647 8837 57736 8840
rect 57295 8781 57381 8837
rect 57437 8781 57593 8837
rect 57649 8781 57736 8837
rect 57295 8622 57736 8781
rect 57295 8619 57383 8622
rect 57435 8619 57595 8622
rect 57647 8619 57736 8622
rect 57295 8563 57381 8619
rect 57437 8563 57593 8619
rect 57649 8563 57736 8619
rect 57295 8404 57736 8563
rect 57295 8402 57383 8404
rect 57435 8402 57595 8404
rect 57647 8402 57736 8404
rect 57295 8346 57381 8402
rect 57437 8346 57593 8402
rect 57649 8346 57736 8402
rect 57295 8187 57736 8346
rect 57295 8184 57383 8187
rect 57435 8184 57595 8187
rect 57647 8184 57736 8187
rect 57295 8128 57381 8184
rect 57437 8128 57593 8184
rect 57649 8128 57736 8184
rect 57295 7969 57736 8128
rect 57295 7966 57383 7969
rect 57435 7966 57595 7969
rect 57647 7966 57736 7969
rect 57295 7910 57381 7966
rect 57437 7910 57593 7966
rect 57649 7910 57736 7966
rect 57295 7752 57736 7910
rect 57295 7749 57383 7752
rect 57435 7749 57595 7752
rect 57647 7749 57736 7752
rect 57295 7693 57381 7749
rect 57437 7693 57593 7749
rect 57649 7693 57736 7749
rect 57295 7534 57736 7693
rect 57295 7531 57383 7534
rect 57435 7531 57595 7534
rect 57647 7531 57736 7534
rect 57295 7475 57381 7531
rect 57437 7475 57593 7531
rect 57649 7475 57736 7531
rect 57295 7316 57736 7475
rect 57295 7313 57383 7316
rect 57435 7313 57595 7316
rect 57647 7313 57736 7316
rect 57295 7257 57381 7313
rect 57437 7257 57593 7313
rect 57649 7257 57736 7313
rect 57295 7099 57736 7257
rect 57295 7096 57383 7099
rect 57435 7096 57595 7099
rect 57647 7096 57736 7099
rect 57295 7040 57381 7096
rect 57437 7040 57593 7096
rect 57649 7040 57736 7096
rect 57295 6881 57736 7040
rect 56124 6836 56886 6874
rect 56124 6780 56160 6836
rect 56216 6780 56371 6836
rect 56427 6780 56583 6836
rect 56639 6780 56794 6836
rect 56850 6780 56886 6836
rect 56124 6618 56886 6780
rect 56124 6562 56160 6618
rect 56216 6562 56371 6618
rect 56427 6562 56583 6618
rect 56639 6562 56794 6618
rect 56850 6562 56886 6618
rect 56124 6400 56886 6562
rect 56124 6344 56160 6400
rect 56216 6344 56371 6400
rect 56427 6344 56583 6400
rect 56639 6344 56794 6400
rect 56850 6344 56886 6400
rect 56124 6306 56886 6344
rect 57295 6829 57383 6881
rect 57435 6829 57595 6881
rect 57647 6829 57736 6881
rect 57295 6663 57736 6829
rect 57295 6611 57383 6663
rect 57435 6611 57595 6663
rect 57647 6611 57736 6663
rect 57295 6446 57736 6611
rect 57295 6394 57383 6446
rect 57435 6394 57595 6446
rect 57647 6394 57736 6446
rect 51642 5199 51822 5211
rect 51642 5147 51654 5199
rect 51810 5147 51822 5199
rect 51642 5135 51822 5147
rect 57295 6228 57736 6394
rect 57295 6176 57383 6228
rect 57435 6176 57595 6228
rect 57647 6176 57736 6228
rect 57295 6120 57736 6176
rect 57295 6064 57381 6120
rect 57437 6064 57593 6120
rect 57649 6064 57736 6120
rect 57295 6011 57736 6064
rect 57295 5959 57383 6011
rect 57435 5959 57595 6011
rect 57647 5959 57736 6011
rect 57295 5902 57736 5959
rect 57295 5846 57381 5902
rect 57437 5846 57593 5902
rect 57649 5846 57736 5902
rect 57295 5793 57736 5846
rect 57295 5741 57383 5793
rect 57435 5741 57595 5793
rect 57647 5741 57736 5793
rect 57295 5575 57736 5741
rect 57295 5523 57383 5575
rect 57435 5523 57595 5575
rect 57647 5523 57736 5575
rect 57295 5358 57736 5523
rect 57295 5306 57383 5358
rect 57435 5306 57595 5358
rect 57647 5306 57736 5358
rect 27387 4535 27476 4587
rect 27528 4535 27688 4587
rect 27740 4535 27828 4587
rect 27387 4370 27828 4535
rect 27387 4318 27476 4370
rect 27528 4318 27688 4370
rect 27740 4318 27828 4370
rect 27387 4152 27828 4318
rect 27387 4100 27476 4152
rect 27528 4100 27688 4152
rect 27740 4100 27828 4152
rect 27387 3934 27828 4100
rect 27387 3882 27476 3934
rect 27528 3882 27688 3934
rect 27740 3882 27828 3934
rect 27387 3837 27828 3882
rect 40588 4904 40812 4928
rect 40588 4852 40622 4904
rect 40778 4852 40812 4904
rect 27387 3781 27474 3837
rect 27530 3781 27686 3837
rect 27742 3781 27828 3837
rect 27387 3717 27828 3781
rect 27387 3665 27476 3717
rect 27528 3665 27688 3717
rect 27740 3665 27828 3717
rect 27387 3619 27828 3665
rect 27387 3563 27474 3619
rect 27530 3563 27686 3619
rect 27742 3563 27828 3619
rect 27387 3524 27828 3563
rect 28764 3837 28894 3876
rect 28764 3781 28801 3837
rect 28857 3781 28894 3837
rect 28764 3619 28894 3781
rect 28764 3563 28801 3619
rect 28857 3563 28894 3619
rect 28764 3525 28894 3563
rect 27936 0 28160 3418
rect 29006 3050 29135 3418
rect 29247 3231 29929 3418
rect 29006 915 29230 3050
rect 29006 655 29090 915
rect 29142 655 29230 915
rect 29006 0 29230 655
rect 29705 915 29929 3231
rect 29705 655 29792 915
rect 29844 655 29929 915
rect 29705 0 29929 655
rect 30859 0 31083 3605
rect 32552 0 32776 3605
rect 34243 0 34467 3605
rect 40588 0 40812 4852
rect 43790 3044 43970 3054
rect 43790 2988 43800 3044
rect 43960 2988 43970 3044
rect 43790 2978 43970 2988
rect 48644 2822 48997 3873
rect 48644 2766 48671 2822
rect 48727 2766 48795 2822
rect 48851 2766 48919 2822
rect 48975 2766 48997 2822
rect 48644 2698 48997 2766
rect 48644 2642 48671 2698
rect 48727 2642 48795 2698
rect 48851 2642 48919 2698
rect 48975 2642 48997 2698
rect 48644 2574 48997 2642
rect 48644 2518 48671 2574
rect 48727 2518 48795 2574
rect 48851 2518 48919 2574
rect 48975 2518 48997 2574
rect 48644 1224 48997 2518
rect 49145 2199 49498 4618
rect 57295 4587 57736 5306
rect 57295 4535 57383 4587
rect 57435 4535 57595 4587
rect 57647 4535 57736 4587
rect 57295 4370 57736 4535
rect 57295 4318 57383 4370
rect 57435 4318 57595 4370
rect 57647 4318 57736 4370
rect 57295 4152 57736 4318
rect 57295 4100 57383 4152
rect 57435 4100 57595 4152
rect 57647 4100 57736 4152
rect 57295 3934 57736 4100
rect 57295 3882 57383 3934
rect 57435 3882 57595 3934
rect 57647 3882 57736 3934
rect 57295 3837 57736 3882
rect 57295 3781 57381 3837
rect 57437 3781 57593 3837
rect 57649 3781 57736 3837
rect 57295 3717 57736 3781
rect 57295 3665 57383 3717
rect 57435 3665 57595 3717
rect 57647 3665 57736 3717
rect 57295 3619 57736 3665
rect 57295 3563 57381 3619
rect 57437 3563 57593 3619
rect 57649 3563 57736 3619
rect 57295 3524 57736 3563
rect 57909 33432 58351 33520
rect 57909 33380 57998 33432
rect 58050 33380 58210 33432
rect 58262 33380 58351 33432
rect 57909 33358 58351 33380
rect 57909 33302 57996 33358
rect 58052 33302 58208 33358
rect 58264 33302 58351 33358
rect 57909 33215 58351 33302
rect 57909 33163 57998 33215
rect 58050 33163 58210 33215
rect 58262 33163 58351 33215
rect 57909 33140 58351 33163
rect 57909 33084 57996 33140
rect 58052 33084 58208 33140
rect 58264 33084 58351 33140
rect 57909 32997 58351 33084
rect 57909 32945 57998 32997
rect 58050 32945 58210 32997
rect 58262 32945 58351 32997
rect 57909 32922 58351 32945
rect 57909 32866 57996 32922
rect 58052 32866 58208 32922
rect 58264 32866 58351 32922
rect 57909 32779 58351 32866
rect 57909 32727 57998 32779
rect 58050 32727 58210 32779
rect 58262 32727 58351 32779
rect 57909 32705 58351 32727
rect 57909 32649 57996 32705
rect 58052 32649 58208 32705
rect 58264 32649 58351 32705
rect 57909 32562 58351 32649
rect 57909 32510 57998 32562
rect 58050 32510 58210 32562
rect 58262 32510 58351 32562
rect 57909 32487 58351 32510
rect 57909 32431 57996 32487
rect 58052 32431 58208 32487
rect 58264 32431 58351 32487
rect 57909 32344 58351 32431
rect 57909 32292 57998 32344
rect 58050 32292 58210 32344
rect 58262 32292 58351 32344
rect 57909 32127 58351 32292
rect 57909 32088 57998 32127
rect 58050 32088 58210 32127
rect 58262 32088 58351 32127
rect 57909 32032 57996 32088
rect 58052 32032 58208 32088
rect 58264 32032 58351 32088
rect 57909 31909 58351 32032
rect 57909 31870 57998 31909
rect 58050 31870 58210 31909
rect 58262 31870 58351 31909
rect 57909 31814 57996 31870
rect 58052 31814 58208 31870
rect 58264 31814 58351 31870
rect 57909 31691 58351 31814
rect 57909 31652 57998 31691
rect 58050 31652 58210 31691
rect 58262 31652 58351 31691
rect 57909 31596 57996 31652
rect 58052 31596 58208 31652
rect 58264 31596 58351 31652
rect 57909 31474 58351 31596
rect 57909 31422 57998 31474
rect 58050 31422 58210 31474
rect 58262 31422 58351 31474
rect 57909 31256 58351 31422
rect 57909 31204 57998 31256
rect 58050 31204 58210 31256
rect 58262 31204 58351 31256
rect 57909 31038 58351 31204
rect 57909 30986 57998 31038
rect 58050 30986 58210 31038
rect 58262 30986 58351 31038
rect 57909 30821 58351 30986
rect 57909 30769 57998 30821
rect 58050 30769 58210 30821
rect 58262 30769 58351 30821
rect 57909 30603 58351 30769
rect 57909 30551 57998 30603
rect 58050 30551 58210 30603
rect 58262 30551 58351 30603
rect 57909 30386 58351 30551
rect 57909 30334 57998 30386
rect 58050 30334 58210 30386
rect 58262 30334 58351 30386
rect 57909 30168 58351 30334
rect 57909 30116 57998 30168
rect 58050 30116 58210 30168
rect 58262 30116 58351 30168
rect 57909 29968 58351 30116
rect 57909 29912 57996 29968
rect 58052 29912 58208 29968
rect 58264 29912 58351 29968
rect 57909 29898 57998 29912
rect 58050 29898 58210 29912
rect 58262 29898 58351 29912
rect 57909 29750 58351 29898
rect 57909 29694 57996 29750
rect 58052 29694 58208 29750
rect 58264 29694 58351 29750
rect 57909 29681 57998 29694
rect 58050 29681 58210 29694
rect 58262 29681 58351 29694
rect 57909 29533 58351 29681
rect 57909 29477 57996 29533
rect 58052 29477 58208 29533
rect 58264 29477 58351 29533
rect 57909 29463 57998 29477
rect 58050 29463 58210 29477
rect 58262 29463 58351 29477
rect 57909 29315 58351 29463
rect 57909 29259 57996 29315
rect 58052 29259 58208 29315
rect 58264 29259 58351 29315
rect 57909 29245 57998 29259
rect 58050 29245 58210 29259
rect 58262 29245 58351 29259
rect 57909 29098 58351 29245
rect 57909 29042 57996 29098
rect 58052 29042 58208 29098
rect 58264 29042 58351 29098
rect 57909 29028 57998 29042
rect 58050 29028 58210 29042
rect 58262 29028 58351 29042
rect 57909 28880 58351 29028
rect 57909 28824 57996 28880
rect 58052 28824 58208 28880
rect 58264 28824 58351 28880
rect 57909 28810 57998 28824
rect 58050 28810 58210 28824
rect 58262 28810 58351 28824
rect 57909 28662 58351 28810
rect 57909 28606 57996 28662
rect 58052 28606 58208 28662
rect 58264 28606 58351 28662
rect 57909 28592 57998 28606
rect 58050 28592 58210 28606
rect 58262 28592 58351 28606
rect 57909 28444 58351 28592
rect 57909 28388 57996 28444
rect 58052 28388 58208 28444
rect 58264 28388 58351 28444
rect 57909 28375 57998 28388
rect 58050 28375 58210 28388
rect 58262 28375 58351 28388
rect 57909 28227 58351 28375
rect 57909 28171 57996 28227
rect 58052 28171 58208 28227
rect 58264 28171 58351 28227
rect 57909 28157 57998 28171
rect 58050 28157 58210 28171
rect 58262 28157 58351 28171
rect 57909 28009 58351 28157
rect 57909 27953 57996 28009
rect 58052 27953 58208 28009
rect 58264 27953 58351 28009
rect 57909 27940 57998 27953
rect 58050 27940 58210 27953
rect 58262 27940 58351 27953
rect 57909 27792 58351 27940
rect 57909 27736 57996 27792
rect 58052 27736 58208 27792
rect 58264 27736 58351 27792
rect 57909 27722 57998 27736
rect 58050 27722 58210 27736
rect 58262 27722 58351 27736
rect 57909 27574 58351 27722
rect 57909 27518 57996 27574
rect 58052 27518 58208 27574
rect 58264 27518 58351 27574
rect 57909 27504 57998 27518
rect 58050 27504 58210 27518
rect 58262 27504 58351 27518
rect 57909 27339 58351 27504
rect 57909 27287 57998 27339
rect 58050 27287 58210 27339
rect 58262 27287 58351 27339
rect 57909 27121 58351 27287
rect 57909 27069 57998 27121
rect 58050 27069 58210 27121
rect 58262 27069 58351 27121
rect 57909 26903 58351 27069
rect 57909 26851 57998 26903
rect 58050 26851 58210 26903
rect 58262 26851 58351 26903
rect 57909 26686 58351 26851
rect 57909 26634 57998 26686
rect 58050 26634 58210 26686
rect 58262 26634 58351 26686
rect 57909 26468 58351 26634
rect 57909 26416 57998 26468
rect 58050 26416 58210 26468
rect 58262 26416 58351 26468
rect 58791 51579 59517 51591
rect 58791 51572 58878 51579
rect 58930 51572 59002 51579
rect 59054 51572 59126 51579
rect 59178 51572 59250 51579
rect 59302 51572 59374 51579
rect 59426 51572 59517 51579
rect 58791 51516 58876 51572
rect 58932 51516 59000 51572
rect 59056 51516 59124 51572
rect 59180 51516 59248 51572
rect 59304 51516 59372 51572
rect 59428 51516 59517 51572
rect 58791 51455 59517 51516
rect 58791 51448 58878 51455
rect 58930 51448 59002 51455
rect 59054 51448 59126 51455
rect 59178 51448 59250 51455
rect 59302 51448 59374 51455
rect 59426 51448 59517 51455
rect 58791 51392 58876 51448
rect 58932 51392 59000 51448
rect 59056 51392 59124 51448
rect 59180 51392 59248 51448
rect 59304 51392 59372 51448
rect 59428 51392 59517 51448
rect 58791 51331 59517 51392
rect 58791 51324 58878 51331
rect 58930 51324 59002 51331
rect 59054 51324 59126 51331
rect 59178 51324 59250 51331
rect 59302 51324 59374 51331
rect 59426 51324 59517 51331
rect 58791 51268 58876 51324
rect 58932 51268 59000 51324
rect 59056 51268 59124 51324
rect 59180 51268 59248 51324
rect 59304 51268 59372 51324
rect 59428 51268 59517 51324
rect 58791 35244 59517 51268
rect 60563 35494 60639 35506
rect 60563 35338 60575 35494
rect 60627 35338 60639 35494
rect 60563 35326 60639 35338
rect 58791 35188 58873 35244
rect 58929 35188 58997 35244
rect 59053 35188 59121 35244
rect 59177 35188 59245 35244
rect 59301 35188 59369 35244
rect 59425 35188 59517 35244
rect 58791 35120 59517 35188
rect 58791 35064 58873 35120
rect 58929 35064 58997 35120
rect 59053 35064 59121 35120
rect 59177 35064 59245 35120
rect 59301 35064 59369 35120
rect 59425 35064 59517 35120
rect 58791 34996 59517 35064
rect 58791 34940 58873 34996
rect 58929 34940 58997 34996
rect 59053 34940 59121 34996
rect 59177 34940 59245 34996
rect 59301 34940 59369 34996
rect 59425 34940 59517 34996
rect 58791 34872 59517 34940
rect 58791 34816 58873 34872
rect 58929 34816 58997 34872
rect 59053 34816 59121 34872
rect 59177 34816 59245 34872
rect 59301 34816 59369 34872
rect 59425 34816 59517 34872
rect 58791 34748 59517 34816
rect 58791 34692 58873 34748
rect 58929 34692 58997 34748
rect 59053 34692 59121 34748
rect 59177 34692 59245 34748
rect 59301 34692 59369 34748
rect 59425 34692 59517 34748
rect 58791 34624 59517 34692
rect 58791 34568 58873 34624
rect 58929 34568 58997 34624
rect 59053 34568 59121 34624
rect 59177 34568 59245 34624
rect 59301 34568 59369 34624
rect 59425 34568 59517 34624
rect 58791 31298 59517 34568
rect 58791 31242 58873 31298
rect 58929 31242 58997 31298
rect 59053 31242 59121 31298
rect 59177 31242 59245 31298
rect 59301 31242 59369 31298
rect 59425 31242 59517 31298
rect 58791 31174 59517 31242
rect 58791 31118 58873 31174
rect 58929 31118 58997 31174
rect 59053 31118 59121 31174
rect 59177 31118 59245 31174
rect 59301 31118 59369 31174
rect 59425 31118 59517 31174
rect 58791 31050 59517 31118
rect 58791 30994 58873 31050
rect 58929 30994 58997 31050
rect 59053 30994 59121 31050
rect 59177 30994 59245 31050
rect 59301 30994 59369 31050
rect 59425 30994 59517 31050
rect 58791 30853 59517 30994
rect 58791 30797 58873 30853
rect 58929 30797 58997 30853
rect 59053 30797 59121 30853
rect 59177 30797 59245 30853
rect 59301 30797 59369 30853
rect 59425 30797 59517 30853
rect 58791 30729 59517 30797
rect 58791 30673 58873 30729
rect 58929 30673 58997 30729
rect 59053 30673 59121 30729
rect 59177 30673 59245 30729
rect 59301 30673 59369 30729
rect 59425 30673 59517 30729
rect 58791 30605 59517 30673
rect 58791 30549 58873 30605
rect 58929 30549 58997 30605
rect 59053 30549 59121 30605
rect 59177 30549 59245 30605
rect 59301 30549 59369 30605
rect 59425 30549 59517 30605
rect 58791 28324 59517 30549
rect 58791 28268 58859 28324
rect 58915 28268 58983 28324
rect 59039 28268 59107 28324
rect 59163 28268 59231 28324
rect 59287 28268 59355 28324
rect 59411 28268 59517 28324
rect 58791 28200 59517 28268
rect 58791 28144 58859 28200
rect 58915 28144 58983 28200
rect 59039 28144 59107 28200
rect 59163 28144 59231 28200
rect 59287 28144 59355 28200
rect 59411 28144 59517 28200
rect 58791 28076 59517 28144
rect 58791 28020 58859 28076
rect 58915 28020 58983 28076
rect 59039 28020 59107 28076
rect 59163 28020 59231 28076
rect 59287 28020 59355 28076
rect 59411 28020 59517 28076
rect 58791 27952 59517 28020
rect 58791 27896 58859 27952
rect 58915 27896 58983 27952
rect 59039 27896 59107 27952
rect 59163 27896 59231 27952
rect 59287 27896 59355 27952
rect 59411 27896 59517 27952
rect 58791 27828 59517 27896
rect 58791 27772 58859 27828
rect 58915 27772 58983 27828
rect 59039 27772 59107 27828
rect 59163 27772 59231 27828
rect 59287 27772 59355 27828
rect 59411 27772 59517 27828
rect 58791 27704 59517 27772
rect 58791 27648 58859 27704
rect 58915 27648 58983 27704
rect 59039 27648 59107 27704
rect 59163 27648 59231 27704
rect 59287 27648 59355 27704
rect 59411 27648 59517 27704
rect 58791 27580 59517 27648
rect 58791 27524 58859 27580
rect 58915 27524 58983 27580
rect 59039 27524 59107 27580
rect 59163 27524 59231 27580
rect 59287 27524 59355 27580
rect 59411 27524 59517 27580
rect 58791 27456 59517 27524
rect 58791 27400 58859 27456
rect 58915 27400 58983 27456
rect 59039 27400 59107 27456
rect 59163 27400 59231 27456
rect 59287 27400 59355 27456
rect 59411 27400 59517 27456
rect 58791 27332 59517 27400
rect 58791 27276 58859 27332
rect 58915 27276 58983 27332
rect 59039 27276 59107 27332
rect 59163 27276 59231 27332
rect 59287 27276 59355 27332
rect 59411 27276 59517 27332
rect 58791 27208 59517 27276
rect 58791 27152 58859 27208
rect 58915 27152 58983 27208
rect 59039 27152 59107 27208
rect 59163 27152 59231 27208
rect 59287 27152 59355 27208
rect 59411 27152 59517 27208
rect 58791 27084 59517 27152
rect 58791 27028 58859 27084
rect 58915 27028 58983 27084
rect 59039 27028 59107 27084
rect 59163 27028 59231 27084
rect 59287 27028 59355 27084
rect 59411 27028 59517 27084
rect 58791 26960 59517 27028
rect 58791 26904 58859 26960
rect 58915 26904 58983 26960
rect 59039 26904 59107 26960
rect 59163 26904 59231 26960
rect 59287 26904 59355 26960
rect 59411 26904 59517 26960
rect 58791 26836 59517 26904
rect 58791 26780 58859 26836
rect 58915 26780 58983 26836
rect 59039 26780 59107 26836
rect 59163 26780 59231 26836
rect 59287 26780 59355 26836
rect 59411 26780 59517 26836
rect 58791 26712 59517 26780
rect 58791 26656 58859 26712
rect 58915 26656 58983 26712
rect 59039 26656 59107 26712
rect 59163 26656 59231 26712
rect 59287 26656 59355 26712
rect 59411 26656 59517 26712
rect 58791 26588 59517 26656
rect 58791 26532 58859 26588
rect 58915 26532 58983 26588
rect 59039 26532 59107 26588
rect 59163 26532 59231 26588
rect 59287 26532 59355 26588
rect 59411 26532 59517 26588
rect 58791 26433 59517 26532
rect 57909 26250 58351 26416
rect 57909 26198 57998 26250
rect 58050 26198 58210 26250
rect 58262 26198 58351 26250
rect 57909 26033 58351 26198
rect 57909 25981 57998 26033
rect 58050 25981 58210 26033
rect 58262 25981 58351 26033
rect 57909 25815 58351 25981
rect 57909 25763 57998 25815
rect 58050 25763 58210 25815
rect 58262 25763 58351 25815
rect 57909 25598 58351 25763
rect 57909 25546 57998 25598
rect 58050 25546 58210 25598
rect 58262 25546 58351 25598
rect 57909 25380 58351 25546
rect 57909 25328 57998 25380
rect 58050 25328 58210 25380
rect 58262 25328 58351 25380
rect 57909 25162 58351 25328
rect 57909 25110 57998 25162
rect 58050 25110 58210 25162
rect 58262 25110 58351 25162
rect 57909 24945 58351 25110
rect 57909 24893 57998 24945
rect 58050 24893 58210 24945
rect 58262 24893 58351 24945
rect 57909 24727 58351 24893
rect 57909 24675 57998 24727
rect 58050 24675 58210 24727
rect 58262 24675 58351 24727
rect 57909 24509 58351 24675
rect 57909 24457 57998 24509
rect 58050 24457 58210 24509
rect 58262 24457 58351 24509
rect 57909 24292 58351 24457
rect 57909 24240 57998 24292
rect 58050 24240 58210 24292
rect 58262 24240 58351 24292
rect 57909 24075 58351 24240
rect 57909 23187 57994 24075
rect 58258 24074 58351 24075
rect 58262 24022 58351 24074
rect 58258 23857 58351 24022
rect 58262 23805 58351 23857
rect 58258 23639 58351 23805
rect 58262 23587 58351 23639
rect 58258 23421 58351 23587
rect 58262 23369 58351 23421
rect 58258 23204 58351 23369
rect 57909 23152 57998 23187
rect 58050 23152 58210 23187
rect 58262 23152 58351 23204
rect 57909 22986 58351 23152
rect 57909 22934 57998 22986
rect 58050 22934 58210 22986
rect 58262 22934 58351 22986
rect 57909 22768 58351 22934
rect 57909 22716 57998 22768
rect 58050 22716 58210 22768
rect 58262 22716 58351 22768
rect 57909 22551 58351 22716
rect 57909 22499 57998 22551
rect 58050 22499 58210 22551
rect 58262 22499 58351 22551
rect 57909 22333 58351 22499
rect 57909 22281 57998 22333
rect 58050 22281 58210 22333
rect 58262 22281 58351 22333
rect 57909 22115 58351 22281
rect 57909 22063 57998 22115
rect 58050 22063 58210 22115
rect 58262 22063 58351 22115
rect 57909 21898 58351 22063
rect 57909 21846 57998 21898
rect 58050 21846 58210 21898
rect 58262 21846 58351 21898
rect 57909 21680 58351 21846
rect 57909 21628 57998 21680
rect 58050 21628 58210 21680
rect 58262 21628 58351 21680
rect 57909 21463 58351 21628
rect 57909 21411 57998 21463
rect 58050 21411 58210 21463
rect 58262 21411 58351 21463
rect 57909 21245 58351 21411
rect 57909 21193 57998 21245
rect 58050 21193 58210 21245
rect 58262 21193 58351 21245
rect 57909 21027 58351 21193
rect 57909 20975 57998 21027
rect 58050 20975 58210 21027
rect 58262 20975 58351 21027
rect 57909 20810 58351 20975
rect 57909 20758 57998 20810
rect 58050 20758 58210 20810
rect 58262 20758 58351 20810
rect 57909 20592 58351 20758
rect 57909 20540 57998 20592
rect 58050 20570 58210 20592
rect 58208 20540 58210 20570
rect 58262 20540 58351 20592
rect 57909 20410 58048 20540
rect 58208 20410 58351 20540
rect 57909 20374 58351 20410
rect 57909 20322 57998 20374
rect 58050 20322 58210 20374
rect 58262 20322 58351 20374
rect 57909 20226 58351 20322
rect 57909 20157 58048 20226
rect 58208 20157 58351 20226
rect 57909 20105 57998 20157
rect 58208 20105 58210 20157
rect 58262 20105 58351 20157
rect 57909 20066 58048 20105
rect 58208 20066 58351 20105
rect 57909 19939 58351 20066
rect 57909 19887 57998 19939
rect 58050 19887 58210 19939
rect 58262 19887 58351 19939
rect 57909 19722 58351 19887
rect 57909 19670 57998 19722
rect 58050 19670 58210 19722
rect 58262 19670 58351 19722
rect 57909 19504 58351 19670
rect 57909 19452 57998 19504
rect 58050 19452 58210 19504
rect 58262 19452 58351 19504
rect 57909 19286 58351 19452
rect 57909 19234 57998 19286
rect 58050 19234 58210 19286
rect 58262 19234 58351 19286
rect 57909 19068 58351 19234
rect 57909 19016 57998 19068
rect 58050 19016 58210 19068
rect 58262 19016 58351 19068
rect 57909 18851 58351 19016
rect 57909 18799 57998 18851
rect 58050 18799 58210 18851
rect 58262 18799 58351 18851
rect 57909 18633 58351 18799
rect 57909 18581 57998 18633
rect 58050 18581 58210 18633
rect 58262 18581 58351 18633
rect 57909 18416 58351 18581
rect 57909 18364 57998 18416
rect 58050 18364 58210 18416
rect 58262 18364 58351 18416
rect 57909 18198 58351 18364
rect 57909 18146 57998 18198
rect 58050 18146 58210 18198
rect 58262 18146 58351 18198
rect 57909 17980 58351 18146
rect 57909 17928 57998 17980
rect 58050 17928 58210 17980
rect 58262 17928 58351 17980
rect 57909 17763 58351 17928
rect 57909 17711 57998 17763
rect 58050 17711 58210 17763
rect 58262 17711 58351 17763
rect 57909 17545 58351 17711
rect 57909 17493 57998 17545
rect 58050 17493 58210 17545
rect 58262 17493 58351 17545
rect 57909 17327 58351 17493
rect 57909 17275 57998 17327
rect 58050 17275 58210 17327
rect 58262 17275 58351 17327
rect 57909 17110 58351 17275
rect 57909 17058 57998 17110
rect 58050 17058 58210 17110
rect 58262 17058 58351 17110
rect 57909 16892 58351 17058
rect 57909 16840 57998 16892
rect 58050 16840 58210 16892
rect 58262 16840 58351 16892
rect 57909 16675 58351 16840
rect 57909 16623 57998 16675
rect 58050 16623 58210 16675
rect 58262 16623 58351 16675
rect 57909 16457 58351 16623
rect 57909 16405 57998 16457
rect 58050 16405 58210 16457
rect 58262 16405 58351 16457
rect 57909 16239 58351 16405
rect 57909 16187 57998 16239
rect 58050 16187 58210 16239
rect 58262 16187 58351 16239
rect 57909 16022 58351 16187
rect 57909 15970 57998 16022
rect 58050 15970 58210 16022
rect 58262 15970 58351 16022
rect 57909 15804 58351 15970
rect 57909 15752 57998 15804
rect 58050 15752 58210 15804
rect 58262 15752 58351 15804
rect 57909 15586 58351 15752
rect 57909 15534 57998 15586
rect 58050 15534 58210 15586
rect 58262 15534 58351 15586
rect 57909 15369 58351 15534
rect 57909 15317 57998 15369
rect 58050 15317 58210 15369
rect 58262 15317 58351 15369
rect 57909 15151 58351 15317
rect 57909 15099 57998 15151
rect 58050 15099 58210 15151
rect 58262 15099 58351 15151
rect 57909 14933 58351 15099
rect 57909 14881 57998 14933
rect 58050 14881 58210 14933
rect 58262 14881 58351 14933
rect 57909 14716 58351 14881
rect 57909 14664 57998 14716
rect 58050 14664 58210 14716
rect 58262 14664 58351 14716
rect 57909 14498 58351 14664
rect 57909 14446 57998 14498
rect 58050 14446 58210 14498
rect 58262 14446 58351 14498
rect 57909 14281 58351 14446
rect 57909 14229 57998 14281
rect 58050 14229 58210 14281
rect 58262 14229 58351 14281
rect 57909 14063 58351 14229
rect 57909 14011 57998 14063
rect 58050 14011 58210 14063
rect 58262 14011 58351 14063
rect 57909 13845 58351 14011
rect 57909 13793 57998 13845
rect 58050 13793 58210 13845
rect 58262 13793 58351 13845
rect 57909 13790 58351 13793
rect 57909 13734 57996 13790
rect 58052 13734 58208 13790
rect 58264 13734 58351 13790
rect 57909 13628 58351 13734
rect 57909 13576 57998 13628
rect 58050 13576 58210 13628
rect 58262 13576 58351 13628
rect 57909 13573 58351 13576
rect 57909 13517 57996 13573
rect 58052 13517 58208 13573
rect 58264 13517 58351 13573
rect 57909 13410 58351 13517
rect 57909 13358 57998 13410
rect 58050 13358 58210 13410
rect 58262 13358 58351 13410
rect 57909 13355 58351 13358
rect 57909 13299 57996 13355
rect 58052 13299 58208 13355
rect 58264 13299 58351 13355
rect 57909 13192 58351 13299
rect 57909 13140 57998 13192
rect 58050 13140 58210 13192
rect 58262 13140 58351 13192
rect 57909 13138 58351 13140
rect 57909 13082 57996 13138
rect 58052 13082 58208 13138
rect 58264 13082 58351 13138
rect 57909 12975 58351 13082
rect 57909 12923 57998 12975
rect 58050 12923 58210 12975
rect 58262 12923 58351 12975
rect 57909 12920 58351 12923
rect 57909 12864 57996 12920
rect 58052 12864 58208 12920
rect 58264 12864 58351 12920
rect 57909 12757 58351 12864
rect 57909 12705 57998 12757
rect 58050 12705 58210 12757
rect 58262 12705 58351 12757
rect 57909 12702 58351 12705
rect 57909 12646 57996 12702
rect 58052 12646 58208 12702
rect 58264 12646 58351 12702
rect 57909 12540 58351 12646
rect 57909 12488 57998 12540
rect 58050 12488 58210 12540
rect 58262 12488 58351 12540
rect 57909 12484 58351 12488
rect 57909 12428 57996 12484
rect 58052 12428 58208 12484
rect 58264 12428 58351 12484
rect 57909 12322 58351 12428
rect 57909 12270 57998 12322
rect 58050 12270 58210 12322
rect 58262 12270 58351 12322
rect 57909 12267 58351 12270
rect 57909 12211 57996 12267
rect 58052 12211 58208 12267
rect 58264 12211 58351 12267
rect 57909 12104 58351 12211
rect 57909 12052 57998 12104
rect 58050 12052 58210 12104
rect 58262 12052 58351 12104
rect 57909 12049 58351 12052
rect 57909 11993 57996 12049
rect 58052 11993 58208 12049
rect 58264 11993 58351 12049
rect 57909 11887 58351 11993
rect 57909 11835 57998 11887
rect 58050 11835 58210 11887
rect 58262 11835 58351 11887
rect 57909 11832 58351 11835
rect 57909 11776 57996 11832
rect 58052 11776 58208 11832
rect 58264 11776 58351 11832
rect 57909 11669 58351 11776
rect 57909 11617 57998 11669
rect 58050 11617 58210 11669
rect 58262 11617 58351 11669
rect 57909 11451 58351 11617
rect 57909 11399 57998 11451
rect 58050 11399 58210 11451
rect 58262 11399 58351 11451
rect 57909 11234 58351 11399
rect 57909 11182 57998 11234
rect 58050 11182 58210 11234
rect 58262 11182 58351 11234
rect 57909 11016 58351 11182
rect 57909 10964 57998 11016
rect 58050 10964 58210 11016
rect 58262 10964 58351 11016
rect 57909 10798 58351 10964
rect 57909 10746 57998 10798
rect 58050 10746 58210 10798
rect 58262 10746 58351 10798
rect 57909 10581 58351 10746
rect 57909 10529 57998 10581
rect 58050 10529 58210 10581
rect 58262 10529 58351 10581
rect 57909 10363 58351 10529
rect 57909 10311 57998 10363
rect 58050 10311 58210 10363
rect 58262 10311 58351 10363
rect 57909 10146 58351 10311
rect 57909 10094 57998 10146
rect 58050 10094 58210 10146
rect 58262 10094 58351 10146
rect 57909 9928 58351 10094
rect 57909 9876 57998 9928
rect 58050 9876 58210 9928
rect 58262 9876 58351 9928
rect 57909 9710 58351 9876
rect 57909 9658 57998 9710
rect 58050 9658 58210 9710
rect 58262 9658 58351 9710
rect 57909 9493 58351 9658
rect 57909 9441 57998 9493
rect 58050 9441 58210 9493
rect 58262 9441 58351 9493
rect 57909 9407 58351 9441
rect 57909 9351 57996 9407
rect 58052 9351 58208 9407
rect 58264 9351 58351 9407
rect 57909 9275 58351 9351
rect 57909 9223 57998 9275
rect 58050 9223 58210 9275
rect 58262 9223 58351 9275
rect 57909 9190 58351 9223
rect 57909 9134 57996 9190
rect 58052 9134 58208 9190
rect 58264 9134 58351 9190
rect 57909 9057 58351 9134
rect 57909 9005 57998 9057
rect 58050 9005 58210 9057
rect 58262 9005 58351 9057
rect 57909 8972 58351 9005
rect 57909 8916 57996 8972
rect 58052 8916 58208 8972
rect 58264 8916 58351 8972
rect 57909 8840 58351 8916
rect 57909 8788 57998 8840
rect 58050 8788 58210 8840
rect 58262 8788 58351 8840
rect 57909 8754 58351 8788
rect 57909 8698 57996 8754
rect 58052 8698 58208 8754
rect 58264 8698 58351 8754
rect 57909 8622 58351 8698
rect 57909 8570 57998 8622
rect 58050 8570 58210 8622
rect 58262 8570 58351 8622
rect 57909 8536 58351 8570
rect 57909 8480 57996 8536
rect 58052 8480 58208 8536
rect 58264 8480 58351 8536
rect 57909 8404 58351 8480
rect 57909 8352 57998 8404
rect 58050 8352 58210 8404
rect 58262 8352 58351 8404
rect 57909 8319 58351 8352
rect 57909 8263 57996 8319
rect 58052 8263 58208 8319
rect 58264 8263 58351 8319
rect 57909 8187 58351 8263
rect 57909 8135 57998 8187
rect 58050 8135 58210 8187
rect 58262 8135 58351 8187
rect 57909 7969 58351 8135
rect 57909 7917 57998 7969
rect 58050 7917 58210 7969
rect 58262 7917 58351 7969
rect 57909 7752 58351 7917
rect 57909 7700 57998 7752
rect 58050 7700 58210 7752
rect 58262 7700 58351 7752
rect 57909 7534 58351 7700
rect 57909 7482 57998 7534
rect 58050 7482 58210 7534
rect 58262 7482 58351 7534
rect 57909 7316 58351 7482
rect 57909 7264 57998 7316
rect 58050 7264 58210 7316
rect 58262 7264 58351 7316
rect 57909 7099 58351 7264
rect 57909 7047 57998 7099
rect 58050 7047 58210 7099
rect 58262 7047 58351 7099
rect 57909 6881 58351 7047
rect 57909 6829 57998 6881
rect 58050 6829 58210 6881
rect 58262 6829 58351 6881
rect 57909 6663 58351 6829
rect 57909 6611 57998 6663
rect 58050 6611 58210 6663
rect 58262 6611 58351 6663
rect 57909 6446 58351 6611
rect 57909 6394 57998 6446
rect 58050 6394 58210 6446
rect 58262 6394 58351 6446
rect 57909 6228 58351 6394
rect 57909 6176 57998 6228
rect 58050 6176 58210 6228
rect 58262 6176 58351 6228
rect 57909 6011 58351 6176
rect 57909 5959 57998 6011
rect 58050 5959 58210 6011
rect 58262 5959 58351 6011
rect 57909 5793 58351 5959
rect 57909 5741 57998 5793
rect 58050 5741 58210 5793
rect 58262 5741 58351 5793
rect 57909 5575 58351 5741
rect 57909 5539 57998 5575
rect 58050 5539 58210 5575
rect 58262 5539 58351 5575
rect 57909 5483 57996 5539
rect 58052 5483 58208 5539
rect 58264 5483 58351 5539
rect 57909 5358 58351 5483
rect 57909 5321 57998 5358
rect 58050 5321 58210 5358
rect 58262 5321 58351 5358
rect 57909 5265 57996 5321
rect 58052 5265 58208 5321
rect 58264 5265 58351 5321
rect 57909 4587 58351 5265
rect 57909 4535 57998 4587
rect 58050 4535 58210 4587
rect 58262 4535 58351 4587
rect 57909 4528 58351 4535
rect 57909 4472 57996 4528
rect 58052 4472 58208 4528
rect 58264 4472 58351 4528
rect 57909 4370 58351 4472
rect 57909 4318 57998 4370
rect 58050 4318 58210 4370
rect 58262 4318 58351 4370
rect 57909 4310 58351 4318
rect 57909 4254 57996 4310
rect 58052 4254 58208 4310
rect 58264 4254 58351 4310
rect 57909 4152 58351 4254
rect 57909 4100 57998 4152
rect 58050 4100 58210 4152
rect 58262 4100 58351 4152
rect 57909 3934 58351 4100
rect 57909 3882 57998 3934
rect 58050 3882 58210 3934
rect 58262 3882 58351 3934
rect 57909 3717 58351 3882
rect 57909 3665 57998 3717
rect 58050 3665 58210 3717
rect 58262 3665 58351 3717
rect 57909 3524 58351 3665
rect 61507 5024 62085 5135
rect 71303 5073 71359 5140
rect 49145 2143 49161 2199
rect 49217 2143 49285 2199
rect 49341 2143 49409 2199
rect 49465 2143 49498 2199
rect 49145 2075 49498 2143
rect 49145 2019 49161 2075
rect 49217 2019 49285 2075
rect 49341 2019 49409 2075
rect 49465 2019 49498 2075
rect 49145 1951 49498 2019
rect 49145 1895 49161 1951
rect 49217 1895 49285 1951
rect 49341 1895 49409 1951
rect 49465 1895 49498 1951
rect 49145 1827 49498 1895
rect 49145 1771 49161 1827
rect 49217 1771 49285 1827
rect 49341 1771 49409 1827
rect 49465 1771 49498 1827
rect 49145 1703 49498 1771
rect 49145 1647 49161 1703
rect 49217 1647 49285 1703
rect 49341 1647 49409 1703
rect 49465 1647 49498 1703
rect 49145 1579 49498 1647
rect 49145 1523 49161 1579
rect 49217 1523 49285 1579
rect 49341 1523 49409 1579
rect 49465 1523 49498 1579
rect 49145 1455 49498 1523
rect 49145 1399 49161 1455
rect 49217 1399 49285 1455
rect 49341 1399 49409 1455
rect 49465 1399 49498 1455
rect 49145 1331 49498 1399
rect 49145 1275 49161 1331
rect 49217 1275 49285 1331
rect 49341 1275 49409 1331
rect 49465 1275 49498 1331
rect 49145 1232 49498 1275
rect 48644 1172 48668 1224
rect 48720 1172 48792 1224
rect 48844 1172 48916 1224
rect 48968 1172 48997 1224
rect 48644 1100 48997 1172
rect 48644 1048 48668 1100
rect 48720 1048 48792 1100
rect 48844 1048 48916 1100
rect 48968 1048 48997 1100
rect 48644 976 48997 1048
rect 48644 924 48668 976
rect 48720 924 48792 976
rect 48844 924 48916 976
rect 48968 924 48997 976
rect 48644 852 48997 924
rect 48644 800 48668 852
rect 48720 800 48792 852
rect 48844 800 48916 852
rect 48968 800 48997 852
rect 48644 728 48997 800
rect 48644 676 48668 728
rect 48720 676 48792 728
rect 48844 676 48916 728
rect 48968 676 48997 728
rect 48644 604 48997 676
rect 48644 552 48668 604
rect 48720 552 48792 604
rect 48844 552 48916 604
rect 48968 552 48997 604
rect 48644 480 48997 552
rect 48644 428 48668 480
rect 48720 428 48792 480
rect 48844 428 48916 480
rect 48968 428 48997 480
rect 48644 356 48997 428
rect 48644 304 48668 356
rect 48720 304 48792 356
rect 48844 304 48916 356
rect 48968 304 48997 356
rect 48644 282 48997 304
rect 50342 0 50566 3517
rect 53772 3255 55669 3418
rect 53772 0 53996 3255
rect 55781 2974 55911 3418
rect 54417 2789 55911 2974
rect 54417 0 54641 2789
rect 56023 2480 56152 3418
rect 55164 2224 56152 2480
rect 55164 0 55388 2224
rect 56265 0 56489 3481
rect 61507 1701 61601 5024
rect 62839 5001 62933 5062
rect 71193 5017 71359 5073
rect 62839 4880 63115 5001
rect 63021 1701 63115 4880
rect 71193 1701 71249 5017
rect 72151 4740 72207 5185
rect 71866 4684 72207 4740
rect 72829 4740 72885 5185
rect 73677 5073 73733 5140
rect 73677 5017 73843 5073
rect 72829 4684 73170 4740
rect 71866 1701 71922 4684
rect 73114 1701 73170 4684
rect 73787 1701 73843 5017
rect 82103 5001 82197 5062
rect 82951 5024 83529 5135
rect 81921 4880 82197 5001
rect 81921 1701 82015 4880
rect 83435 1701 83529 5024
rect 61447 0 61671 1701
rect 62115 1689 62339 1701
rect 62115 1637 62150 1689
rect 62306 1637 62339 1689
rect 62115 0 62339 1637
rect 62958 0 63182 1701
rect 71109 0 71333 1701
rect 71782 0 72006 1701
rect 72180 1689 72404 1701
rect 72180 1637 72215 1689
rect 72371 1637 72404 1689
rect 72180 0 72404 1637
rect 72630 1689 72854 1701
rect 72630 1637 72665 1689
rect 72821 1637 72854 1689
rect 72630 0 72854 1637
rect 73030 0 73254 1701
rect 73703 0 73927 1701
rect 81855 0 82079 1701
rect 82695 1689 82919 1701
rect 82695 1637 82730 1689
rect 82886 1637 82919 1689
rect 82695 0 82919 1637
rect 83372 0 83596 1701
<< via2 >>
rect 25398 51527 25400 51572
rect 25400 51527 25452 51572
rect 25452 51527 25454 51572
rect 25398 51516 25454 51527
rect 25522 51527 25524 51572
rect 25524 51527 25576 51572
rect 25576 51527 25578 51572
rect 25522 51516 25578 51527
rect 25646 51527 25648 51572
rect 25648 51527 25700 51572
rect 25700 51527 25702 51572
rect 25646 51516 25702 51527
rect 25770 51527 25772 51572
rect 25772 51527 25824 51572
rect 25824 51527 25826 51572
rect 25770 51516 25826 51527
rect 25894 51527 25896 51572
rect 25896 51527 25948 51572
rect 25948 51527 25950 51572
rect 25894 51516 25950 51527
rect 25398 51403 25400 51448
rect 25400 51403 25452 51448
rect 25452 51403 25454 51448
rect 25398 51392 25454 51403
rect 25522 51403 25524 51448
rect 25524 51403 25576 51448
rect 25576 51403 25578 51448
rect 25522 51392 25578 51403
rect 25646 51403 25648 51448
rect 25648 51403 25700 51448
rect 25700 51403 25702 51448
rect 25646 51392 25702 51403
rect 25770 51403 25772 51448
rect 25772 51403 25824 51448
rect 25824 51403 25826 51448
rect 25770 51392 25826 51403
rect 25894 51403 25896 51448
rect 25896 51403 25948 51448
rect 25948 51403 25950 51448
rect 25894 51392 25950 51403
rect 25398 51279 25400 51324
rect 25400 51279 25452 51324
rect 25452 51279 25454 51324
rect 25398 51268 25454 51279
rect 25522 51279 25524 51324
rect 25524 51279 25576 51324
rect 25576 51279 25578 51324
rect 25522 51268 25578 51279
rect 25646 51279 25648 51324
rect 25648 51279 25700 51324
rect 25700 51279 25702 51324
rect 25646 51268 25702 51279
rect 25770 51279 25772 51324
rect 25772 51279 25824 51324
rect 25824 51279 25826 51324
rect 25770 51268 25826 51279
rect 25894 51279 25896 51324
rect 25896 51279 25948 51324
rect 25948 51279 25950 51324
rect 25894 51268 25950 51279
rect 25384 35219 25440 35275
rect 25508 35219 25564 35275
rect 25632 35219 25688 35275
rect 25756 35219 25812 35275
rect 25880 35219 25936 35275
rect 25384 35095 25440 35151
rect 25508 35095 25564 35151
rect 25632 35095 25688 35151
rect 25756 35095 25812 35151
rect 25880 35095 25936 35151
rect 25384 34971 25440 35027
rect 25508 34971 25564 35027
rect 25632 34971 25688 35027
rect 25756 34971 25812 35027
rect 25880 34971 25936 35027
rect 25384 34847 25440 34903
rect 25508 34847 25564 34903
rect 25632 34847 25688 34903
rect 25756 34847 25812 34903
rect 25880 34847 25936 34903
rect 25384 34723 25440 34779
rect 25508 34723 25564 34779
rect 25632 34723 25688 34779
rect 25756 34723 25812 34779
rect 25880 34723 25936 34779
rect 25384 34599 25440 34655
rect 25508 34599 25564 34655
rect 25632 34599 25688 34655
rect 25756 34599 25812 34655
rect 25880 34599 25936 34655
rect 25398 31192 25454 31248
rect 25522 31192 25578 31248
rect 25646 31192 25702 31248
rect 25770 31192 25826 31248
rect 25894 31192 25950 31248
rect 25398 31068 25454 31124
rect 25522 31068 25578 31124
rect 25646 31068 25702 31124
rect 25770 31068 25826 31124
rect 25894 31068 25950 31124
rect 25398 30944 25454 31000
rect 25522 30944 25578 31000
rect 25646 30944 25702 31000
rect 25770 30944 25826 31000
rect 25894 30944 25950 31000
rect 25398 30737 25454 30793
rect 25522 30737 25578 30793
rect 25646 30737 25702 30793
rect 25770 30737 25826 30793
rect 25894 30737 25950 30793
rect 25398 30613 25454 30669
rect 25522 30613 25578 30669
rect 25646 30613 25702 30669
rect 25770 30613 25826 30669
rect 25894 30613 25950 30669
rect 25398 30489 25454 30545
rect 25522 30489 25578 30545
rect 25646 30489 25702 30545
rect 25770 30489 25826 30545
rect 25894 30489 25950 30545
rect 25404 28207 25460 28263
rect 25528 28207 25584 28263
rect 25652 28207 25708 28263
rect 25776 28207 25832 28263
rect 25900 28207 25956 28263
rect 25404 28083 25460 28139
rect 25528 28083 25584 28139
rect 25652 28083 25708 28139
rect 25776 28083 25832 28139
rect 25900 28083 25956 28139
rect 25404 27959 25460 28015
rect 25528 27959 25584 28015
rect 25652 27959 25708 28015
rect 25776 27959 25832 28015
rect 25900 27959 25956 28015
rect 25404 27835 25460 27891
rect 25528 27835 25584 27891
rect 25652 27835 25708 27891
rect 25776 27835 25832 27891
rect 25900 27835 25956 27891
rect 25404 27711 25460 27767
rect 25528 27711 25584 27767
rect 25652 27711 25708 27767
rect 25776 27711 25832 27767
rect 25900 27711 25956 27767
rect 25404 27587 25460 27643
rect 25528 27587 25584 27643
rect 25652 27587 25708 27643
rect 25776 27587 25832 27643
rect 25900 27587 25956 27643
rect 25404 27463 25460 27519
rect 25528 27463 25584 27519
rect 25652 27463 25708 27519
rect 25776 27463 25832 27519
rect 25900 27463 25956 27519
rect 25404 27339 25460 27395
rect 25528 27339 25584 27395
rect 25652 27339 25708 27395
rect 25776 27339 25832 27395
rect 25900 27339 25956 27395
rect 25404 27215 25460 27271
rect 25528 27215 25584 27271
rect 25652 27215 25708 27271
rect 25776 27215 25832 27271
rect 25900 27215 25956 27271
rect 25404 27091 25460 27147
rect 25528 27091 25584 27147
rect 25652 27091 25708 27147
rect 25776 27091 25832 27147
rect 25900 27091 25956 27147
rect 25404 26967 25460 27023
rect 25528 26967 25584 27023
rect 25652 26967 25708 27023
rect 25776 26967 25832 27023
rect 25900 26967 25956 27023
rect 25404 26843 25460 26899
rect 25528 26843 25584 26899
rect 25652 26843 25708 26899
rect 25776 26843 25832 26899
rect 25900 26843 25956 26899
rect 25404 26719 25460 26775
rect 25528 26719 25584 26775
rect 25652 26719 25708 26775
rect 25776 26719 25832 26775
rect 25900 26719 25956 26775
rect 25404 26595 25460 26651
rect 25528 26595 25584 26651
rect 25652 26595 25708 26651
rect 25776 26595 25832 26651
rect 25900 26595 25956 26651
rect 25404 26471 25460 26527
rect 25528 26471 25584 26527
rect 25652 26471 25708 26527
rect 25776 26471 25832 26527
rect 25900 26471 25956 26527
rect 26859 33955 26915 34011
rect 27071 33955 27127 34011
rect 26859 33737 26915 33793
rect 27071 33737 27127 33793
rect 26859 33520 26915 33576
rect 27071 33520 27127 33576
rect 26859 33302 26915 33358
rect 27071 33302 27127 33358
rect 26859 33084 26915 33140
rect 27071 33084 27127 33140
rect 26859 32866 26915 32922
rect 27071 32866 27127 32922
rect 26859 32649 26915 32705
rect 27071 32649 27127 32705
rect 26859 32431 26915 32487
rect 27071 32431 27127 32487
rect 26859 32075 26861 32088
rect 26861 32075 26913 32088
rect 26913 32075 26915 32088
rect 26859 32032 26915 32075
rect 27071 32075 27073 32088
rect 27073 32075 27125 32088
rect 27125 32075 27127 32088
rect 27071 32032 27127 32075
rect 26859 31857 26861 31870
rect 26861 31857 26913 31870
rect 26913 31857 26915 31870
rect 26859 31814 26915 31857
rect 27071 31857 27073 31870
rect 27073 31857 27125 31870
rect 27125 31857 27127 31870
rect 27071 31814 27127 31857
rect 26859 31639 26861 31652
rect 26861 31639 26913 31652
rect 26913 31639 26915 31652
rect 26859 31596 26915 31639
rect 27071 31639 27073 31652
rect 27073 31639 27125 31652
rect 27125 31639 27127 31652
rect 27071 31596 27127 31639
rect 26859 29950 26915 29968
rect 26859 29912 26861 29950
rect 26861 29912 26913 29950
rect 26913 29912 26915 29950
rect 27071 29950 27127 29968
rect 27071 29912 27073 29950
rect 27073 29912 27125 29950
rect 27125 29912 27127 29950
rect 26859 29733 26915 29750
rect 26859 29694 26861 29733
rect 26861 29694 26913 29733
rect 26913 29694 26915 29733
rect 27071 29733 27127 29750
rect 27071 29694 27073 29733
rect 27073 29694 27125 29733
rect 27125 29694 27127 29733
rect 26859 29515 26915 29533
rect 26859 29477 26861 29515
rect 26861 29477 26913 29515
rect 26913 29477 26915 29515
rect 27071 29515 27127 29533
rect 27071 29477 27073 29515
rect 27073 29477 27125 29515
rect 27125 29477 27127 29515
rect 26859 29297 26915 29315
rect 26859 29259 26861 29297
rect 26861 29259 26913 29297
rect 26913 29259 26915 29297
rect 27071 29297 27127 29315
rect 27071 29259 27073 29297
rect 27073 29259 27125 29297
rect 27125 29259 27127 29297
rect 26859 29080 26915 29098
rect 26859 29042 26861 29080
rect 26861 29042 26913 29080
rect 26913 29042 26915 29080
rect 27071 29080 27127 29098
rect 27071 29042 27073 29080
rect 27073 29042 27125 29080
rect 27125 29042 27127 29080
rect 26859 28862 26915 28880
rect 26859 28824 26861 28862
rect 26861 28824 26913 28862
rect 26913 28824 26915 28862
rect 27071 28862 27127 28880
rect 27071 28824 27073 28862
rect 27073 28824 27125 28862
rect 27125 28824 27127 28862
rect 26859 28644 26915 28662
rect 26859 28606 26861 28644
rect 26861 28606 26913 28644
rect 26913 28606 26915 28644
rect 27071 28644 27127 28662
rect 27071 28606 27073 28644
rect 27073 28606 27125 28644
rect 27125 28606 27127 28644
rect 26859 28427 26915 28444
rect 26859 28388 26861 28427
rect 26861 28388 26913 28427
rect 26913 28388 26915 28427
rect 27071 28427 27127 28444
rect 27071 28388 27073 28427
rect 27073 28388 27125 28427
rect 27125 28388 27127 28427
rect 26859 28209 26915 28227
rect 26859 28171 26861 28209
rect 26861 28171 26913 28209
rect 26913 28171 26915 28209
rect 27071 28209 27127 28227
rect 27071 28171 27073 28209
rect 27073 28171 27125 28209
rect 27125 28171 27127 28209
rect 26859 27992 26915 28009
rect 26859 27953 26861 27992
rect 26861 27953 26913 27992
rect 26913 27953 26915 27992
rect 27071 27992 27127 28009
rect 27071 27953 27073 27992
rect 27073 27953 27125 27992
rect 27125 27953 27127 27992
rect 26859 27774 26915 27792
rect 26859 27736 26861 27774
rect 26861 27736 26913 27774
rect 26913 27736 26915 27774
rect 27071 27774 27127 27792
rect 27071 27736 27073 27774
rect 27073 27736 27125 27774
rect 27125 27736 27127 27774
rect 26859 27556 26915 27574
rect 26859 27518 26861 27556
rect 26861 27518 26913 27556
rect 26913 27518 26915 27556
rect 27071 27556 27127 27574
rect 27071 27518 27073 27556
rect 27073 27518 27125 27556
rect 27125 27518 27127 27556
rect 26450 26126 26610 26286
rect 26092 25807 26252 25967
rect 25756 25487 25916 25647
rect 25421 25168 25581 25328
rect 25081 24477 25241 24637
rect 24744 24156 24904 24316
rect 24416 23835 24576 23995
rect 24057 23513 24217 23673
rect 26465 19532 26625 19692
rect 26858 24074 27122 24075
rect 26858 24022 26861 24074
rect 26861 24022 26913 24074
rect 26913 24022 27073 24074
rect 27073 24022 27122 24074
rect 26858 23857 27122 24022
rect 26858 23805 26861 23857
rect 26861 23805 26913 23857
rect 26913 23805 27073 23857
rect 27073 23805 27122 23857
rect 26858 23639 27122 23805
rect 26858 23587 26861 23639
rect 26861 23587 26913 23639
rect 26913 23587 27073 23639
rect 27073 23587 27122 23639
rect 26858 23421 27122 23587
rect 26858 23369 26861 23421
rect 26861 23369 26913 23421
rect 26913 23369 27073 23421
rect 27073 23369 27122 23421
rect 26858 23204 27122 23369
rect 26858 23187 26861 23204
rect 26861 23187 26913 23204
rect 26913 23187 27073 23204
rect 27073 23187 27122 23204
rect 26924 20540 27073 20570
rect 27073 20540 27084 20570
rect 26924 20410 27084 20540
rect 26924 20157 27084 20226
rect 26924 20105 27073 20157
rect 27073 20105 27084 20157
rect 26924 20066 27084 20105
rect 26107 19187 26267 19347
rect 25771 18867 25931 19027
rect 25434 18524 25594 18684
rect 25094 18190 25254 18350
rect 24757 17817 24917 17977
rect 24429 17496 24589 17656
rect 24069 17157 24229 17317
rect 26859 14063 26915 14119
rect 27071 14063 27127 14119
rect 26859 13846 26915 13902
rect 27071 13846 27127 13902
rect 26859 13628 26915 13684
rect 27071 13628 27127 13684
rect 26859 13411 26915 13467
rect 27071 13411 27127 13467
rect 26859 13193 26915 13249
rect 27071 13193 27127 13249
rect 26859 12975 26915 13031
rect 27071 12975 27127 13031
rect 26859 12757 26915 12813
rect 27071 12757 27127 12813
rect 26859 12540 26915 12596
rect 27071 12540 27127 12596
rect 26859 12322 26915 12378
rect 27071 12322 27127 12378
rect 26859 12105 26915 12161
rect 27071 12105 27127 12161
rect 26859 9351 26915 9407
rect 27071 9351 27127 9407
rect 26859 9134 26915 9190
rect 27071 9134 27127 9190
rect 26859 8916 26915 8972
rect 27071 8916 27127 8972
rect 26859 8698 26915 8754
rect 27071 8698 27127 8754
rect 26859 8480 26915 8536
rect 27071 8480 27127 8536
rect 26859 8263 26915 8319
rect 27071 8263 27127 8319
rect 26859 5523 26861 5539
rect 26861 5523 26913 5539
rect 26913 5523 26915 5539
rect 26859 5483 26915 5523
rect 27071 5523 27073 5539
rect 27073 5523 27125 5539
rect 27125 5523 27127 5539
rect 27071 5483 27127 5523
rect 26859 5306 26861 5321
rect 26861 5306 26913 5321
rect 26913 5306 26915 5321
rect 26859 5265 26915 5306
rect 27071 5306 27073 5321
rect 27073 5306 27125 5321
rect 27125 5306 27127 5321
rect 27071 5265 27127 5306
rect 27788 51453 27844 51455
rect 27788 51401 27790 51453
rect 27790 51401 27842 51453
rect 27842 51401 27844 51453
rect 27788 51399 27844 51401
rect 27999 51453 28055 51455
rect 27999 51401 28001 51453
rect 28001 51401 28053 51453
rect 28053 51401 28055 51453
rect 27999 51399 28055 51401
rect 28210 51453 28266 51455
rect 28210 51401 28212 51453
rect 28212 51401 28264 51453
rect 28264 51401 28266 51453
rect 28210 51399 28266 51401
rect 28421 51453 28477 51455
rect 28421 51401 28423 51453
rect 28423 51401 28475 51453
rect 28475 51401 28477 51453
rect 28421 51399 28477 51401
rect 28632 51453 28688 51455
rect 28632 51401 28634 51453
rect 28634 51401 28686 51453
rect 28686 51401 28688 51453
rect 28632 51399 28688 51401
rect 28843 51453 28899 51455
rect 28843 51401 28845 51453
rect 28845 51401 28897 51453
rect 28897 51401 28899 51453
rect 28843 51399 28899 51401
rect 29054 51453 29110 51455
rect 29054 51401 29056 51453
rect 29056 51401 29108 51453
rect 29108 51401 29110 51453
rect 29054 51399 29110 51401
rect 56013 51453 56069 51455
rect 56013 51401 56015 51453
rect 56015 51401 56067 51453
rect 56067 51401 56069 51453
rect 56013 51399 56069 51401
rect 56224 51453 56280 51455
rect 56224 51401 56226 51453
rect 56226 51401 56278 51453
rect 56278 51401 56280 51453
rect 56224 51399 56280 51401
rect 56435 51453 56491 51455
rect 56435 51401 56437 51453
rect 56437 51401 56489 51453
rect 56489 51401 56491 51453
rect 56435 51399 56491 51401
rect 56646 51453 56702 51455
rect 56646 51401 56648 51453
rect 56648 51401 56700 51453
rect 56700 51401 56702 51453
rect 56646 51399 56702 51401
rect 56857 51453 56913 51455
rect 56857 51401 56859 51453
rect 56859 51401 56911 51453
rect 56911 51401 56913 51453
rect 56857 51399 56913 51401
rect 57068 51453 57124 51455
rect 57068 51401 57070 51453
rect 57070 51401 57122 51453
rect 57122 51401 57124 51453
rect 57068 51399 57124 51401
rect 57279 51453 57335 51455
rect 57279 51401 57281 51453
rect 57281 51401 57333 51453
rect 57333 51401 57335 51453
rect 57279 51399 57335 51401
rect 41875 50453 42035 50613
rect 27788 49653 27844 49655
rect 27788 49601 27790 49653
rect 27790 49601 27842 49653
rect 27842 49601 27844 49653
rect 27788 49599 27844 49601
rect 27999 49653 28055 49655
rect 27999 49601 28001 49653
rect 28001 49601 28053 49653
rect 28053 49601 28055 49653
rect 27999 49599 28055 49601
rect 28210 49653 28266 49655
rect 28210 49601 28212 49653
rect 28212 49601 28264 49653
rect 28264 49601 28266 49653
rect 28210 49599 28266 49601
rect 28421 49653 28477 49655
rect 28421 49601 28423 49653
rect 28423 49601 28475 49653
rect 28475 49601 28477 49653
rect 28421 49599 28477 49601
rect 28632 49653 28688 49655
rect 28632 49601 28634 49653
rect 28634 49601 28686 49653
rect 28686 49601 28688 49653
rect 28632 49599 28688 49601
rect 28843 49653 28899 49655
rect 28843 49601 28845 49653
rect 28845 49601 28897 49653
rect 28897 49601 28899 49653
rect 28843 49599 28899 49601
rect 29054 49653 29110 49655
rect 29054 49601 29056 49653
rect 29056 49601 29108 49653
rect 29108 49601 29110 49653
rect 29054 49599 29110 49601
rect 56013 49653 56069 49655
rect 56013 49601 56015 49653
rect 56015 49601 56067 49653
rect 56067 49601 56069 49653
rect 56013 49599 56069 49601
rect 56224 49653 56280 49655
rect 56224 49601 56226 49653
rect 56226 49601 56278 49653
rect 56278 49601 56280 49653
rect 56224 49599 56280 49601
rect 56435 49653 56491 49655
rect 56435 49601 56437 49653
rect 56437 49601 56489 49653
rect 56489 49601 56491 49653
rect 56435 49599 56491 49601
rect 56646 49653 56702 49655
rect 56646 49601 56648 49653
rect 56648 49601 56700 49653
rect 56700 49601 56702 49653
rect 56646 49599 56702 49601
rect 56857 49653 56913 49655
rect 56857 49601 56859 49653
rect 56859 49601 56911 49653
rect 56911 49601 56913 49653
rect 56857 49599 56913 49601
rect 57068 49653 57124 49655
rect 57068 49601 57070 49653
rect 57070 49601 57122 49653
rect 57122 49601 57124 49653
rect 57068 49599 57124 49601
rect 57279 49653 57335 49655
rect 57279 49601 57281 49653
rect 57281 49601 57333 49653
rect 57333 49601 57335 49653
rect 57279 49599 57335 49601
rect 27788 47853 27844 47855
rect 27788 47801 27790 47853
rect 27790 47801 27842 47853
rect 27842 47801 27844 47853
rect 27788 47799 27844 47801
rect 27999 47853 28055 47855
rect 27999 47801 28001 47853
rect 28001 47801 28053 47853
rect 28053 47801 28055 47853
rect 27999 47799 28055 47801
rect 28210 47853 28266 47855
rect 28210 47801 28212 47853
rect 28212 47801 28264 47853
rect 28264 47801 28266 47853
rect 28210 47799 28266 47801
rect 28421 47853 28477 47855
rect 28421 47801 28423 47853
rect 28423 47801 28475 47853
rect 28475 47801 28477 47853
rect 28421 47799 28477 47801
rect 28632 47853 28688 47855
rect 28632 47801 28634 47853
rect 28634 47801 28686 47853
rect 28686 47801 28688 47853
rect 28632 47799 28688 47801
rect 28843 47853 28899 47855
rect 28843 47801 28845 47853
rect 28845 47801 28897 47853
rect 28897 47801 28899 47853
rect 28843 47799 28899 47801
rect 29054 47853 29110 47855
rect 29054 47801 29056 47853
rect 29056 47801 29108 47853
rect 29108 47801 29110 47853
rect 29054 47799 29110 47801
rect 56013 47853 56069 47855
rect 56013 47801 56015 47853
rect 56015 47801 56067 47853
rect 56067 47801 56069 47853
rect 56013 47799 56069 47801
rect 56224 47853 56280 47855
rect 56224 47801 56226 47853
rect 56226 47801 56278 47853
rect 56278 47801 56280 47853
rect 56224 47799 56280 47801
rect 56435 47853 56491 47855
rect 56435 47801 56437 47853
rect 56437 47801 56489 47853
rect 56489 47801 56491 47853
rect 56435 47799 56491 47801
rect 56646 47853 56702 47855
rect 56646 47801 56648 47853
rect 56648 47801 56700 47853
rect 56700 47801 56702 47853
rect 56646 47799 56702 47801
rect 56857 47853 56913 47855
rect 56857 47801 56859 47853
rect 56859 47801 56911 47853
rect 56911 47801 56913 47853
rect 56857 47799 56913 47801
rect 57068 47853 57124 47855
rect 57068 47801 57070 47853
rect 57070 47801 57122 47853
rect 57122 47801 57124 47853
rect 57068 47799 57124 47801
rect 57279 47853 57335 47855
rect 57279 47801 57281 47853
rect 57281 47801 57333 47853
rect 57333 47801 57335 47853
rect 57279 47799 57335 47801
rect 27788 46053 27844 46055
rect 27788 46001 27790 46053
rect 27790 46001 27842 46053
rect 27842 46001 27844 46053
rect 27788 45999 27844 46001
rect 27999 46053 28055 46055
rect 27999 46001 28001 46053
rect 28001 46001 28053 46053
rect 28053 46001 28055 46053
rect 27999 45999 28055 46001
rect 28210 46053 28266 46055
rect 28210 46001 28212 46053
rect 28212 46001 28264 46053
rect 28264 46001 28266 46053
rect 28210 45999 28266 46001
rect 28421 46053 28477 46055
rect 28421 46001 28423 46053
rect 28423 46001 28475 46053
rect 28475 46001 28477 46053
rect 28421 45999 28477 46001
rect 28632 46053 28688 46055
rect 28632 46001 28634 46053
rect 28634 46001 28686 46053
rect 28686 46001 28688 46053
rect 28632 45999 28688 46001
rect 28843 46053 28899 46055
rect 28843 46001 28845 46053
rect 28845 46001 28897 46053
rect 28897 46001 28899 46053
rect 28843 45999 28899 46001
rect 29054 46053 29110 46055
rect 29054 46001 29056 46053
rect 29056 46001 29108 46053
rect 29108 46001 29110 46053
rect 29054 45999 29110 46001
rect 56013 46053 56069 46055
rect 56013 46001 56015 46053
rect 56015 46001 56067 46053
rect 56067 46001 56069 46053
rect 56013 45999 56069 46001
rect 56224 46053 56280 46055
rect 56224 46001 56226 46053
rect 56226 46001 56278 46053
rect 56278 46001 56280 46053
rect 56224 45999 56280 46001
rect 56435 46053 56491 46055
rect 56435 46001 56437 46053
rect 56437 46001 56489 46053
rect 56489 46001 56491 46053
rect 56435 45999 56491 46001
rect 56646 46053 56702 46055
rect 56646 46001 56648 46053
rect 56648 46001 56700 46053
rect 56700 46001 56702 46053
rect 56646 45999 56702 46001
rect 56857 46053 56913 46055
rect 56857 46001 56859 46053
rect 56859 46001 56911 46053
rect 56911 46001 56913 46053
rect 56857 45999 56913 46001
rect 57068 46053 57124 46055
rect 57068 46001 57070 46053
rect 57070 46001 57122 46053
rect 57122 46001 57124 46053
rect 57068 45999 57124 46001
rect 57279 46053 57335 46055
rect 57279 46001 57281 46053
rect 57281 46001 57333 46053
rect 57333 46001 57335 46053
rect 57279 45999 57335 46001
rect 27788 44253 27844 44255
rect 27788 44201 27790 44253
rect 27790 44201 27842 44253
rect 27842 44201 27844 44253
rect 27788 44199 27844 44201
rect 27999 44253 28055 44255
rect 27999 44201 28001 44253
rect 28001 44201 28053 44253
rect 28053 44201 28055 44253
rect 27999 44199 28055 44201
rect 28210 44253 28266 44255
rect 28210 44201 28212 44253
rect 28212 44201 28264 44253
rect 28264 44201 28266 44253
rect 28210 44199 28266 44201
rect 28421 44253 28477 44255
rect 28421 44201 28423 44253
rect 28423 44201 28475 44253
rect 28475 44201 28477 44253
rect 28421 44199 28477 44201
rect 28632 44253 28688 44255
rect 28632 44201 28634 44253
rect 28634 44201 28686 44253
rect 28686 44201 28688 44253
rect 28632 44199 28688 44201
rect 28843 44253 28899 44255
rect 28843 44201 28845 44253
rect 28845 44201 28897 44253
rect 28897 44201 28899 44253
rect 28843 44199 28899 44201
rect 29054 44253 29110 44255
rect 29054 44201 29056 44253
rect 29056 44201 29108 44253
rect 29108 44201 29110 44253
rect 29054 44199 29110 44201
rect 56013 44253 56069 44255
rect 56013 44201 56015 44253
rect 56015 44201 56067 44253
rect 56067 44201 56069 44253
rect 56013 44199 56069 44201
rect 56224 44253 56280 44255
rect 56224 44201 56226 44253
rect 56226 44201 56278 44253
rect 56278 44201 56280 44253
rect 56224 44199 56280 44201
rect 56435 44253 56491 44255
rect 56435 44201 56437 44253
rect 56437 44201 56489 44253
rect 56489 44201 56491 44253
rect 56435 44199 56491 44201
rect 56646 44253 56702 44255
rect 56646 44201 56648 44253
rect 56648 44201 56700 44253
rect 56700 44201 56702 44253
rect 56646 44199 56702 44201
rect 56857 44253 56913 44255
rect 56857 44201 56859 44253
rect 56859 44201 56911 44253
rect 56911 44201 56913 44253
rect 56857 44199 56913 44201
rect 57068 44253 57124 44255
rect 57068 44201 57070 44253
rect 57070 44201 57122 44253
rect 57122 44201 57124 44253
rect 57068 44199 57124 44201
rect 57279 44253 57335 44255
rect 57279 44201 57281 44253
rect 57281 44201 57333 44253
rect 57333 44201 57335 44253
rect 57279 44199 57335 44201
rect 27788 42453 27844 42455
rect 27788 42401 27790 42453
rect 27790 42401 27842 42453
rect 27842 42401 27844 42453
rect 27788 42399 27844 42401
rect 27999 42453 28055 42455
rect 27999 42401 28001 42453
rect 28001 42401 28053 42453
rect 28053 42401 28055 42453
rect 27999 42399 28055 42401
rect 28210 42453 28266 42455
rect 28210 42401 28212 42453
rect 28212 42401 28264 42453
rect 28264 42401 28266 42453
rect 28210 42399 28266 42401
rect 28421 42453 28477 42455
rect 28421 42401 28423 42453
rect 28423 42401 28475 42453
rect 28475 42401 28477 42453
rect 28421 42399 28477 42401
rect 28632 42453 28688 42455
rect 28632 42401 28634 42453
rect 28634 42401 28686 42453
rect 28686 42401 28688 42453
rect 28632 42399 28688 42401
rect 28843 42453 28899 42455
rect 28843 42401 28845 42453
rect 28845 42401 28897 42453
rect 28897 42401 28899 42453
rect 28843 42399 28899 42401
rect 29054 42453 29110 42455
rect 29054 42401 29056 42453
rect 29056 42401 29108 42453
rect 29108 42401 29110 42453
rect 29054 42399 29110 42401
rect 56013 42453 56069 42455
rect 56013 42401 56015 42453
rect 56015 42401 56067 42453
rect 56067 42401 56069 42453
rect 56013 42399 56069 42401
rect 56224 42453 56280 42455
rect 56224 42401 56226 42453
rect 56226 42401 56278 42453
rect 56278 42401 56280 42453
rect 56224 42399 56280 42401
rect 56435 42453 56491 42455
rect 56435 42401 56437 42453
rect 56437 42401 56489 42453
rect 56489 42401 56491 42453
rect 56435 42399 56491 42401
rect 56646 42453 56702 42455
rect 56646 42401 56648 42453
rect 56648 42401 56700 42453
rect 56700 42401 56702 42453
rect 56646 42399 56702 42401
rect 56857 42453 56913 42455
rect 56857 42401 56859 42453
rect 56859 42401 56911 42453
rect 56911 42401 56913 42453
rect 56857 42399 56913 42401
rect 57068 42453 57124 42455
rect 57068 42401 57070 42453
rect 57070 42401 57122 42453
rect 57122 42401 57124 42453
rect 57068 42399 57124 42401
rect 57279 42453 57335 42455
rect 57279 42401 57281 42453
rect 57281 42401 57333 42453
rect 57333 42401 57335 42453
rect 57279 42399 57335 42401
rect 27788 40653 27844 40655
rect 27788 40601 27790 40653
rect 27790 40601 27842 40653
rect 27842 40601 27844 40653
rect 27788 40599 27844 40601
rect 27999 40653 28055 40655
rect 27999 40601 28001 40653
rect 28001 40601 28053 40653
rect 28053 40601 28055 40653
rect 27999 40599 28055 40601
rect 28210 40653 28266 40655
rect 28210 40601 28212 40653
rect 28212 40601 28264 40653
rect 28264 40601 28266 40653
rect 28210 40599 28266 40601
rect 28421 40653 28477 40655
rect 28421 40601 28423 40653
rect 28423 40601 28475 40653
rect 28475 40601 28477 40653
rect 28421 40599 28477 40601
rect 28632 40653 28688 40655
rect 28632 40601 28634 40653
rect 28634 40601 28686 40653
rect 28686 40601 28688 40653
rect 28632 40599 28688 40601
rect 28843 40653 28899 40655
rect 28843 40601 28845 40653
rect 28845 40601 28897 40653
rect 28897 40601 28899 40653
rect 28843 40599 28899 40601
rect 29054 40653 29110 40655
rect 29054 40601 29056 40653
rect 29056 40601 29108 40653
rect 29108 40601 29110 40653
rect 29054 40599 29110 40601
rect 56013 40653 56069 40655
rect 56013 40601 56015 40653
rect 56015 40601 56067 40653
rect 56067 40601 56069 40653
rect 56013 40599 56069 40601
rect 56224 40653 56280 40655
rect 56224 40601 56226 40653
rect 56226 40601 56278 40653
rect 56278 40601 56280 40653
rect 56224 40599 56280 40601
rect 56435 40653 56491 40655
rect 56435 40601 56437 40653
rect 56437 40601 56489 40653
rect 56489 40601 56491 40653
rect 56435 40599 56491 40601
rect 56646 40653 56702 40655
rect 56646 40601 56648 40653
rect 56648 40601 56700 40653
rect 56700 40601 56702 40653
rect 56646 40599 56702 40601
rect 56857 40653 56913 40655
rect 56857 40601 56859 40653
rect 56859 40601 56911 40653
rect 56911 40601 56913 40653
rect 56857 40599 56913 40601
rect 57068 40653 57124 40655
rect 57068 40601 57070 40653
rect 57070 40601 57122 40653
rect 57122 40601 57124 40653
rect 57068 40599 57124 40601
rect 57279 40653 57335 40655
rect 57279 40601 57281 40653
rect 57281 40601 57333 40653
rect 57333 40601 57335 40653
rect 57279 40599 57335 40601
rect 27788 38853 27844 38855
rect 27788 38801 27790 38853
rect 27790 38801 27842 38853
rect 27842 38801 27844 38853
rect 27788 38799 27844 38801
rect 27999 38853 28055 38855
rect 27999 38801 28001 38853
rect 28001 38801 28053 38853
rect 28053 38801 28055 38853
rect 27999 38799 28055 38801
rect 28210 38853 28266 38855
rect 28210 38801 28212 38853
rect 28212 38801 28264 38853
rect 28264 38801 28266 38853
rect 28210 38799 28266 38801
rect 28421 38853 28477 38855
rect 28421 38801 28423 38853
rect 28423 38801 28475 38853
rect 28475 38801 28477 38853
rect 28421 38799 28477 38801
rect 28632 38853 28688 38855
rect 28632 38801 28634 38853
rect 28634 38801 28686 38853
rect 28686 38801 28688 38853
rect 28632 38799 28688 38801
rect 28843 38853 28899 38855
rect 28843 38801 28845 38853
rect 28845 38801 28897 38853
rect 28897 38801 28899 38853
rect 28843 38799 28899 38801
rect 29054 38853 29110 38855
rect 29054 38801 29056 38853
rect 29056 38801 29108 38853
rect 29108 38801 29110 38853
rect 29054 38799 29110 38801
rect 56013 38853 56069 38855
rect 56013 38801 56015 38853
rect 56015 38801 56067 38853
rect 56067 38801 56069 38853
rect 56013 38799 56069 38801
rect 56224 38853 56280 38855
rect 56224 38801 56226 38853
rect 56226 38801 56278 38853
rect 56278 38801 56280 38853
rect 56224 38799 56280 38801
rect 56435 38853 56491 38855
rect 56435 38801 56437 38853
rect 56437 38801 56489 38853
rect 56489 38801 56491 38853
rect 56435 38799 56491 38801
rect 56646 38853 56702 38855
rect 56646 38801 56648 38853
rect 56648 38801 56700 38853
rect 56700 38801 56702 38853
rect 56646 38799 56702 38801
rect 56857 38853 56913 38855
rect 56857 38801 56859 38853
rect 56859 38801 56911 38853
rect 56911 38801 56913 38853
rect 56857 38799 56913 38801
rect 57068 38853 57124 38855
rect 57068 38801 57070 38853
rect 57070 38801 57122 38853
rect 57122 38801 57124 38853
rect 57068 38799 57124 38801
rect 57279 38853 57335 38855
rect 57279 38801 57281 38853
rect 57281 38801 57333 38853
rect 57333 38801 57335 38853
rect 57279 38799 57335 38801
rect 27788 37053 27844 37055
rect 27788 37001 27790 37053
rect 27790 37001 27842 37053
rect 27842 37001 27844 37053
rect 27788 36999 27844 37001
rect 27999 37053 28055 37055
rect 27999 37001 28001 37053
rect 28001 37001 28053 37053
rect 28053 37001 28055 37053
rect 27999 36999 28055 37001
rect 28210 37053 28266 37055
rect 28210 37001 28212 37053
rect 28212 37001 28264 37053
rect 28264 37001 28266 37053
rect 28210 36999 28266 37001
rect 28421 37053 28477 37055
rect 28421 37001 28423 37053
rect 28423 37001 28475 37053
rect 28475 37001 28477 37053
rect 28421 36999 28477 37001
rect 28632 37053 28688 37055
rect 28632 37001 28634 37053
rect 28634 37001 28686 37053
rect 28686 37001 28688 37053
rect 28632 36999 28688 37001
rect 28843 37053 28899 37055
rect 28843 37001 28845 37053
rect 28845 37001 28897 37053
rect 28897 37001 28899 37053
rect 28843 36999 28899 37001
rect 29054 37053 29110 37055
rect 29054 37001 29056 37053
rect 29056 37001 29108 37053
rect 29108 37001 29110 37053
rect 29054 36999 29110 37001
rect 56013 37053 56069 37055
rect 56013 37001 56015 37053
rect 56015 37001 56067 37053
rect 56067 37001 56069 37053
rect 56013 36999 56069 37001
rect 56224 37053 56280 37055
rect 56224 37001 56226 37053
rect 56226 37001 56278 37053
rect 56278 37001 56280 37053
rect 56224 36999 56280 37001
rect 56435 37053 56491 37055
rect 56435 37001 56437 37053
rect 56437 37001 56489 37053
rect 56489 37001 56491 37053
rect 56435 36999 56491 37001
rect 56646 37053 56702 37055
rect 56646 37001 56648 37053
rect 56648 37001 56700 37053
rect 56700 37001 56702 37053
rect 56646 36999 56702 37001
rect 56857 37053 56913 37055
rect 56857 37001 56859 37053
rect 56859 37001 56911 37053
rect 56911 37001 56913 37053
rect 56857 36999 56913 37001
rect 57068 37053 57124 37055
rect 57068 37001 57070 37053
rect 57070 37001 57122 37053
rect 57122 37001 57124 37053
rect 57068 36999 57124 37001
rect 57279 37053 57335 37055
rect 57279 37001 57281 37053
rect 57281 37001 57333 37053
rect 57333 37001 57335 37053
rect 57279 36999 57335 37001
rect 36958 35825 37014 35881
rect 37169 35825 37225 35881
rect 37381 35825 37437 35881
rect 37592 35825 37648 35881
rect 27438 35273 27494 35275
rect 27438 35221 27440 35273
rect 27440 35221 27492 35273
rect 27492 35221 27494 35273
rect 27438 35219 27494 35221
rect 27562 35273 27618 35275
rect 27562 35221 27564 35273
rect 27564 35221 27616 35273
rect 27616 35221 27618 35273
rect 27562 35219 27618 35221
rect 27686 35273 27742 35275
rect 27686 35221 27688 35273
rect 27688 35221 27740 35273
rect 27740 35221 27742 35273
rect 27686 35219 27742 35221
rect 27438 35149 27494 35151
rect 27438 35097 27440 35149
rect 27440 35097 27492 35149
rect 27492 35097 27494 35149
rect 27438 35095 27494 35097
rect 27562 35149 27618 35151
rect 27562 35097 27564 35149
rect 27564 35097 27616 35149
rect 27616 35097 27618 35149
rect 27562 35095 27618 35097
rect 27686 35149 27742 35151
rect 27686 35097 27688 35149
rect 27688 35097 27740 35149
rect 27740 35097 27742 35149
rect 27686 35095 27742 35097
rect 27438 35025 27494 35027
rect 27438 34973 27440 35025
rect 27440 34973 27492 35025
rect 27492 34973 27494 35025
rect 27438 34971 27494 34973
rect 27562 35025 27618 35027
rect 27562 34973 27564 35025
rect 27564 34973 27616 35025
rect 27616 34973 27618 35025
rect 27562 34971 27618 34973
rect 27686 35025 27742 35027
rect 27686 34973 27688 35025
rect 27688 34973 27740 35025
rect 27740 34973 27742 35025
rect 27686 34971 27742 34973
rect 27438 34901 27494 34903
rect 27438 34849 27440 34901
rect 27440 34849 27492 34901
rect 27492 34849 27494 34901
rect 27438 34847 27494 34849
rect 27562 34901 27618 34903
rect 27562 34849 27564 34901
rect 27564 34849 27616 34901
rect 27616 34849 27618 34901
rect 27562 34847 27618 34849
rect 27686 34901 27742 34903
rect 27686 34849 27688 34901
rect 27688 34849 27740 34901
rect 27740 34849 27742 34901
rect 27686 34847 27742 34849
rect 27438 34777 27494 34779
rect 27438 34725 27440 34777
rect 27440 34725 27492 34777
rect 27492 34725 27494 34777
rect 27438 34723 27494 34725
rect 27562 34777 27618 34779
rect 27562 34725 27564 34777
rect 27564 34725 27616 34777
rect 27616 34725 27618 34777
rect 27562 34723 27618 34725
rect 27686 34777 27742 34779
rect 27686 34725 27688 34777
rect 27688 34725 27740 34777
rect 27740 34725 27742 34777
rect 27686 34723 27742 34725
rect 27438 34653 27494 34655
rect 27438 34601 27440 34653
rect 27440 34601 27492 34653
rect 27492 34601 27494 34653
rect 27438 34599 27494 34601
rect 27562 34653 27618 34655
rect 27562 34601 27564 34653
rect 27564 34601 27616 34653
rect 27616 34601 27618 34653
rect 27562 34599 27618 34601
rect 27686 34653 27742 34655
rect 27686 34601 27688 34653
rect 27688 34601 27740 34653
rect 27740 34601 27742 34653
rect 27686 34599 27742 34601
rect 57996 33955 58052 34011
rect 58208 33955 58264 34011
rect 57996 33737 58052 33793
rect 58208 33737 58264 33793
rect 57996 33520 58052 33576
rect 58208 33520 58264 33576
rect 27474 33085 27530 33141
rect 27686 33085 27742 33141
rect 27474 32867 27530 32923
rect 27686 32867 27742 32923
rect 27474 32649 27530 32705
rect 27686 32649 27742 32705
rect 27474 32431 27530 32487
rect 27686 32431 27742 32487
rect 27474 31204 27476 31252
rect 27476 31204 27528 31252
rect 27528 31204 27530 31252
rect 27474 31196 27530 31204
rect 27686 31204 27688 31252
rect 27688 31204 27740 31252
rect 27740 31204 27742 31252
rect 27686 31196 27742 31204
rect 27474 30986 27476 31034
rect 27476 30986 27528 31034
rect 27528 30986 27530 31034
rect 27474 30978 27530 30986
rect 27686 30986 27688 31034
rect 27688 30986 27740 31034
rect 27740 30986 27742 31034
rect 27686 30978 27742 30986
rect 27474 30769 27476 30816
rect 27476 30769 27528 30816
rect 27528 30769 27530 30816
rect 27474 30760 27530 30769
rect 27686 30769 27688 30816
rect 27688 30769 27740 30816
rect 27740 30769 27742 30816
rect 27686 30760 27742 30769
rect 27474 30551 27476 30598
rect 27476 30551 27528 30598
rect 27528 30551 27530 30598
rect 27474 30542 27530 30551
rect 27686 30551 27688 30598
rect 27688 30551 27740 30598
rect 27740 30551 27742 30598
rect 27686 30542 27742 30551
rect 27474 26743 27530 26799
rect 27686 26743 27742 26799
rect 27474 26525 27530 26581
rect 27686 26525 27742 26581
rect 27474 24972 27530 25028
rect 27686 24972 27742 25028
rect 27474 24754 27530 24810
rect 27686 24754 27742 24810
rect 27475 22934 27476 22936
rect 27476 22934 27528 22936
rect 27528 22934 27688 22936
rect 27688 22934 27739 22936
rect 27475 22768 27739 22934
rect 27475 22716 27476 22768
rect 27476 22716 27528 22768
rect 27528 22716 27688 22768
rect 27688 22716 27739 22768
rect 27475 22551 27739 22716
rect 27475 22499 27476 22551
rect 27476 22499 27528 22551
rect 27528 22499 27688 22551
rect 27688 22499 27739 22551
rect 27475 22333 27739 22499
rect 27475 22281 27476 22333
rect 27476 22281 27528 22333
rect 27528 22281 27688 22333
rect 27688 22281 27739 22333
rect 27475 22115 27739 22281
rect 27475 22063 27476 22115
rect 27476 22063 27528 22115
rect 27528 22063 27688 22115
rect 27688 22063 27739 22115
rect 27475 22048 27739 22063
rect 27474 16457 27530 16470
rect 27474 16414 27476 16457
rect 27476 16414 27528 16457
rect 27528 16414 27530 16457
rect 27686 16457 27742 16470
rect 27686 16414 27688 16457
rect 27688 16414 27740 16457
rect 27740 16414 27742 16457
rect 27474 16239 27530 16253
rect 27474 16197 27476 16239
rect 27476 16197 27528 16239
rect 27528 16197 27530 16239
rect 27686 16239 27742 16253
rect 27686 16197 27688 16239
rect 27688 16197 27740 16239
rect 27740 16197 27742 16239
rect 27474 16022 27530 16035
rect 27474 15979 27476 16022
rect 27476 15979 27528 16022
rect 27528 15979 27530 16022
rect 27686 16022 27742 16035
rect 27686 15979 27688 16022
rect 27688 15979 27740 16022
rect 27740 15979 27742 16022
rect 27474 15804 27530 15818
rect 27474 15762 27476 15804
rect 27476 15762 27528 15804
rect 27528 15762 27530 15804
rect 27686 15804 27742 15818
rect 27686 15762 27688 15804
rect 27688 15762 27740 15804
rect 27740 15762 27742 15804
rect 27474 15586 27530 15600
rect 27474 15544 27476 15586
rect 27476 15544 27528 15586
rect 27528 15544 27530 15586
rect 27686 15586 27742 15600
rect 27686 15544 27688 15586
rect 27688 15544 27740 15586
rect 27740 15544 27742 15586
rect 27474 15369 27530 15382
rect 27474 15326 27476 15369
rect 27476 15326 27528 15369
rect 27528 15326 27530 15369
rect 27686 15369 27742 15382
rect 27686 15326 27688 15369
rect 27688 15326 27740 15369
rect 27740 15326 27742 15369
rect 27474 15151 27530 15164
rect 27474 15108 27476 15151
rect 27476 15108 27528 15151
rect 27528 15108 27530 15151
rect 27686 15151 27742 15164
rect 27686 15108 27688 15151
rect 27688 15108 27740 15151
rect 27740 15108 27742 15151
rect 27474 14933 27530 14947
rect 27474 14891 27476 14933
rect 27476 14891 27528 14933
rect 27528 14891 27530 14933
rect 27686 14933 27742 14947
rect 27686 14891 27688 14933
rect 27688 14891 27740 14933
rect 27740 14891 27742 14933
rect 27474 14716 27530 14729
rect 27474 14673 27476 14716
rect 27476 14673 27528 14716
rect 27528 14673 27530 14716
rect 27686 14716 27742 14729
rect 27686 14673 27688 14716
rect 27688 14673 27740 14716
rect 27740 14673 27742 14716
rect 27474 14498 27530 14512
rect 27474 14456 27476 14498
rect 27476 14456 27528 14498
rect 27528 14456 27530 14498
rect 27686 14498 27742 14512
rect 27686 14456 27688 14498
rect 27688 14456 27740 14498
rect 27740 14456 27742 14498
rect 27474 14229 27476 14231
rect 27476 14229 27528 14231
rect 27528 14229 27530 14231
rect 27474 14175 27530 14229
rect 27686 14229 27688 14231
rect 27688 14229 27740 14231
rect 27740 14229 27742 14231
rect 27686 14175 27742 14229
rect 27474 14011 27476 14014
rect 27476 14011 27528 14014
rect 27528 14011 27530 14014
rect 27474 13958 27530 14011
rect 27686 14011 27688 14014
rect 27688 14011 27740 14014
rect 27740 14011 27742 14014
rect 27686 13958 27742 14011
rect 27474 13793 27476 13796
rect 27476 13793 27528 13796
rect 27528 13793 27530 13796
rect 27474 13740 27530 13793
rect 27686 13793 27688 13796
rect 27688 13793 27740 13796
rect 27740 13793 27742 13796
rect 27686 13740 27742 13793
rect 27474 13576 27476 13578
rect 27476 13576 27528 13578
rect 27528 13576 27530 13578
rect 27474 13522 27530 13576
rect 27686 13576 27688 13578
rect 27688 13576 27740 13578
rect 27740 13576 27742 13578
rect 27686 13522 27742 13576
rect 27474 13358 27476 13361
rect 27476 13358 27528 13361
rect 27528 13358 27530 13361
rect 27474 13305 27530 13358
rect 27686 13358 27688 13361
rect 27688 13358 27740 13361
rect 27740 13358 27742 13361
rect 27686 13305 27742 13358
rect 27474 11399 27476 11406
rect 27476 11399 27528 11406
rect 27528 11399 27530 11406
rect 27474 11350 27530 11399
rect 27686 11399 27688 11406
rect 27688 11399 27740 11406
rect 27740 11399 27742 11406
rect 27686 11350 27742 11399
rect 27474 11182 27476 11189
rect 27476 11182 27528 11189
rect 27528 11182 27530 11189
rect 27474 11133 27530 11182
rect 27686 11182 27688 11189
rect 27688 11182 27740 11189
rect 27740 11182 27742 11189
rect 27686 11133 27742 11182
rect 27474 10964 27476 10971
rect 27476 10964 27528 10971
rect 27528 10964 27530 10971
rect 27474 10915 27530 10964
rect 27686 10964 27688 10971
rect 27688 10964 27740 10971
rect 27740 10964 27742 10971
rect 27686 10915 27742 10964
rect 27474 10746 27476 10753
rect 27476 10746 27528 10753
rect 27528 10746 27530 10753
rect 27474 10697 27530 10746
rect 27686 10746 27688 10753
rect 27688 10746 27740 10753
rect 27740 10746 27742 10753
rect 27686 10697 27742 10746
rect 27474 10529 27476 10535
rect 27476 10529 27528 10535
rect 27528 10529 27530 10535
rect 27474 10479 27530 10529
rect 27686 10529 27688 10535
rect 27688 10529 27740 10535
rect 27740 10529 27742 10535
rect 27686 10479 27742 10529
rect 27474 10311 27476 10318
rect 27476 10311 27528 10318
rect 27528 10311 27530 10318
rect 27474 10262 27530 10311
rect 27686 10311 27688 10318
rect 27688 10311 27740 10318
rect 27740 10311 27742 10318
rect 27686 10262 27742 10311
rect 57381 33085 57437 33141
rect 57593 33085 57649 33141
rect 57381 32867 57437 32923
rect 57593 32867 57649 32923
rect 57381 32649 57437 32705
rect 57593 32649 57649 32705
rect 57381 32431 57437 32487
rect 57593 32431 57649 32487
rect 57381 31204 57383 31252
rect 57383 31204 57435 31252
rect 57435 31204 57437 31252
rect 57381 31196 57437 31204
rect 57593 31204 57595 31252
rect 57595 31204 57647 31252
rect 57647 31204 57649 31252
rect 57593 31196 57649 31204
rect 57381 30986 57383 31034
rect 57383 30986 57435 31034
rect 57435 30986 57437 31034
rect 57381 30978 57437 30986
rect 57593 30986 57595 31034
rect 57595 30986 57647 31034
rect 57647 30986 57649 31034
rect 57593 30978 57649 30986
rect 57381 30769 57383 30816
rect 57383 30769 57435 30816
rect 57435 30769 57437 30816
rect 57381 30760 57437 30769
rect 57593 30769 57595 30816
rect 57595 30769 57647 30816
rect 57647 30769 57649 30816
rect 57593 30760 57649 30769
rect 57381 30551 57383 30598
rect 57383 30551 57435 30598
rect 57435 30551 57437 30598
rect 57381 30542 57437 30551
rect 57593 30551 57595 30598
rect 57595 30551 57647 30598
rect 57647 30551 57649 30598
rect 57593 30542 57649 30551
rect 57381 26743 57437 26799
rect 57593 26743 57649 26799
rect 57381 26525 57437 26581
rect 57593 26525 57649 26581
rect 57363 22768 57627 22923
rect 57363 22716 57383 22768
rect 57383 22716 57435 22768
rect 57435 22716 57595 22768
rect 57595 22716 57627 22768
rect 57363 22551 57627 22716
rect 57363 22499 57383 22551
rect 57383 22499 57435 22551
rect 57435 22499 57595 22551
rect 57595 22499 57627 22551
rect 57363 22333 57627 22499
rect 57363 22281 57383 22333
rect 57383 22281 57435 22333
rect 57435 22281 57595 22333
rect 57595 22281 57627 22333
rect 57363 22115 57627 22281
rect 57363 22063 57383 22115
rect 57383 22063 57435 22115
rect 57435 22063 57595 22115
rect 57595 22063 57627 22115
rect 57363 22035 57627 22063
rect 57381 16675 57437 16678
rect 57381 16623 57383 16675
rect 57383 16623 57435 16675
rect 57435 16623 57437 16675
rect 57381 16622 57437 16623
rect 57593 16675 57649 16678
rect 57593 16623 57595 16675
rect 57595 16623 57647 16675
rect 57647 16623 57649 16675
rect 57593 16622 57649 16623
rect 57381 16457 57437 16461
rect 57381 16405 57383 16457
rect 57383 16405 57435 16457
rect 57435 16405 57437 16457
rect 57593 16457 57649 16461
rect 57593 16405 57595 16457
rect 57595 16405 57647 16457
rect 57647 16405 57649 16457
rect 57381 16239 57437 16243
rect 57381 16187 57383 16239
rect 57383 16187 57435 16239
rect 57435 16187 57437 16239
rect 57593 16239 57649 16243
rect 57593 16187 57595 16239
rect 57595 16187 57647 16239
rect 57647 16187 57649 16239
rect 57381 16022 57437 16026
rect 57381 15970 57383 16022
rect 57383 15970 57435 16022
rect 57435 15970 57437 16022
rect 57593 16022 57649 16026
rect 57593 15970 57595 16022
rect 57595 15970 57647 16022
rect 57647 15970 57649 16022
rect 57381 15804 57437 15808
rect 57381 15752 57383 15804
rect 57383 15752 57435 15804
rect 57435 15752 57437 15804
rect 57593 15804 57649 15808
rect 57593 15752 57595 15804
rect 57595 15752 57647 15804
rect 57647 15752 57649 15804
rect 57381 15586 57437 15590
rect 57381 15534 57383 15586
rect 57383 15534 57435 15586
rect 57435 15534 57437 15586
rect 57593 15586 57649 15590
rect 57593 15534 57595 15586
rect 57595 15534 57647 15586
rect 57647 15534 57649 15586
rect 57381 15369 57437 15372
rect 57381 15317 57383 15369
rect 57383 15317 57435 15369
rect 57435 15317 57437 15369
rect 57381 15316 57437 15317
rect 57593 15369 57649 15372
rect 57593 15317 57595 15369
rect 57595 15317 57647 15369
rect 57647 15317 57649 15369
rect 57593 15316 57649 15317
rect 57381 15151 57437 15155
rect 57381 15099 57383 15151
rect 57383 15099 57435 15151
rect 57435 15099 57437 15151
rect 57593 15151 57649 15155
rect 57593 15099 57595 15151
rect 57595 15099 57647 15151
rect 57647 15099 57649 15151
rect 57381 14933 57437 14937
rect 57381 14881 57383 14933
rect 57383 14881 57435 14933
rect 57435 14881 57437 14933
rect 57593 14933 57649 14937
rect 57593 14881 57595 14933
rect 57595 14881 57647 14933
rect 57647 14881 57649 14933
rect 57381 14716 57437 14720
rect 57381 14664 57383 14716
rect 57383 14664 57435 14716
rect 57435 14664 57437 14716
rect 57593 14716 57649 14720
rect 57593 14664 57595 14716
rect 57595 14664 57647 14716
rect 57647 14664 57649 14716
rect 57381 11399 57383 11406
rect 57383 11399 57435 11406
rect 57435 11399 57437 11406
rect 57381 11350 57437 11399
rect 57593 11399 57595 11406
rect 57595 11399 57647 11406
rect 57647 11399 57649 11406
rect 57593 11350 57649 11399
rect 57381 11182 57383 11189
rect 57383 11182 57435 11189
rect 57435 11182 57437 11189
rect 57381 11133 57437 11182
rect 57593 11182 57595 11189
rect 57595 11182 57647 11189
rect 57647 11182 57649 11189
rect 57593 11133 57649 11182
rect 57381 10964 57383 10971
rect 57383 10964 57435 10971
rect 57435 10964 57437 10971
rect 57381 10915 57437 10964
rect 57593 10964 57595 10971
rect 57595 10964 57647 10971
rect 57647 10964 57649 10971
rect 57593 10915 57649 10964
rect 57381 10746 57383 10753
rect 57383 10746 57435 10753
rect 57435 10746 57437 10753
rect 57381 10697 57437 10746
rect 57593 10746 57595 10753
rect 57595 10746 57647 10753
rect 57647 10746 57649 10753
rect 57593 10697 57649 10746
rect 57381 10529 57383 10535
rect 57383 10529 57435 10535
rect 57435 10529 57437 10535
rect 57381 10479 57437 10529
rect 57593 10529 57595 10535
rect 57595 10529 57647 10535
rect 57647 10529 57649 10535
rect 57593 10479 57649 10529
rect 57381 10311 57383 10318
rect 57383 10311 57435 10318
rect 57435 10311 57437 10318
rect 57381 10262 57437 10311
rect 57593 10311 57595 10318
rect 57595 10311 57647 10318
rect 57647 10311 57649 10318
rect 57593 10262 57649 10311
rect 51766 9811 51822 9971
rect 49906 8900 50066 8956
rect 27474 7534 27530 7535
rect 27474 7482 27476 7534
rect 27476 7482 27528 7534
rect 27528 7482 27530 7534
rect 27474 7479 27530 7482
rect 27686 7534 27742 7535
rect 27686 7482 27688 7534
rect 27688 7482 27740 7534
rect 27740 7482 27742 7534
rect 27686 7479 27742 7482
rect 27474 7316 27530 7317
rect 27474 7264 27476 7316
rect 27476 7264 27528 7316
rect 27528 7264 27530 7316
rect 27474 7261 27530 7264
rect 27686 7316 27742 7317
rect 27686 7264 27688 7316
rect 27688 7264 27740 7316
rect 27740 7264 27742 7316
rect 27686 7261 27742 7264
rect 27474 7047 27476 7099
rect 27476 7047 27528 7099
rect 27528 7047 27530 7099
rect 27474 7043 27530 7047
rect 27686 7047 27688 7099
rect 27688 7047 27740 7099
rect 27740 7047 27742 7099
rect 27686 7043 27742 7047
rect 28273 6780 28329 6836
rect 28484 6780 28540 6836
rect 28696 6780 28752 6836
rect 28907 6780 28963 6836
rect 28273 6562 28329 6618
rect 28484 6562 28540 6618
rect 28696 6562 28752 6618
rect 28907 6562 28963 6618
rect 28273 6344 28329 6400
rect 28484 6344 28540 6400
rect 28696 6344 28752 6400
rect 28907 6344 28963 6400
rect 27474 6064 27530 6120
rect 27686 6064 27742 6120
rect 27474 5846 27530 5902
rect 27686 5846 27742 5902
rect 26859 4472 26915 4528
rect 27071 4472 27127 4528
rect 26859 4254 26915 4310
rect 27071 4254 27127 4310
rect 57381 8788 57383 8837
rect 57383 8788 57435 8837
rect 57435 8788 57437 8837
rect 57381 8781 57437 8788
rect 57593 8788 57595 8837
rect 57595 8788 57647 8837
rect 57647 8788 57649 8837
rect 57593 8781 57649 8788
rect 57381 8570 57383 8619
rect 57383 8570 57435 8619
rect 57435 8570 57437 8619
rect 57381 8563 57437 8570
rect 57593 8570 57595 8619
rect 57595 8570 57647 8619
rect 57647 8570 57649 8619
rect 57593 8563 57649 8570
rect 57381 8352 57383 8402
rect 57383 8352 57435 8402
rect 57435 8352 57437 8402
rect 57381 8346 57437 8352
rect 57593 8352 57595 8402
rect 57595 8352 57647 8402
rect 57647 8352 57649 8402
rect 57593 8346 57649 8352
rect 57381 8135 57383 8184
rect 57383 8135 57435 8184
rect 57435 8135 57437 8184
rect 57381 8128 57437 8135
rect 57593 8135 57595 8184
rect 57595 8135 57647 8184
rect 57647 8135 57649 8184
rect 57593 8128 57649 8135
rect 57381 7917 57383 7966
rect 57383 7917 57435 7966
rect 57435 7917 57437 7966
rect 57381 7910 57437 7917
rect 57593 7917 57595 7966
rect 57595 7917 57647 7966
rect 57647 7917 57649 7966
rect 57593 7910 57649 7917
rect 57381 7700 57383 7749
rect 57383 7700 57435 7749
rect 57435 7700 57437 7749
rect 57381 7693 57437 7700
rect 57593 7700 57595 7749
rect 57595 7700 57647 7749
rect 57647 7700 57649 7749
rect 57593 7693 57649 7700
rect 57381 7482 57383 7531
rect 57383 7482 57435 7531
rect 57435 7482 57437 7531
rect 57381 7475 57437 7482
rect 57593 7482 57595 7531
rect 57595 7482 57647 7531
rect 57647 7482 57649 7531
rect 57593 7475 57649 7482
rect 57381 7264 57383 7313
rect 57383 7264 57435 7313
rect 57435 7264 57437 7313
rect 57381 7257 57437 7264
rect 57593 7264 57595 7313
rect 57595 7264 57647 7313
rect 57647 7264 57649 7313
rect 57593 7257 57649 7264
rect 57381 7047 57383 7096
rect 57383 7047 57435 7096
rect 57435 7047 57437 7096
rect 57381 7040 57437 7047
rect 57593 7047 57595 7096
rect 57595 7047 57647 7096
rect 57647 7047 57649 7096
rect 57593 7040 57649 7047
rect 56160 6780 56216 6836
rect 56371 6780 56427 6836
rect 56583 6780 56639 6836
rect 56794 6780 56850 6836
rect 56160 6562 56216 6618
rect 56371 6562 56427 6618
rect 56583 6562 56639 6618
rect 56794 6562 56850 6618
rect 56160 6344 56216 6400
rect 56371 6344 56427 6400
rect 56583 6344 56639 6400
rect 56794 6344 56850 6400
rect 57381 6064 57437 6120
rect 57593 6064 57649 6120
rect 57381 5846 57437 5902
rect 57593 5846 57649 5902
rect 27474 3781 27530 3837
rect 27686 3781 27742 3837
rect 27474 3563 27530 3619
rect 27686 3563 27742 3619
rect 28801 3781 28857 3837
rect 28801 3563 28857 3619
rect 43800 2988 43960 3044
rect 48671 2766 48727 2822
rect 48795 2766 48851 2822
rect 48919 2766 48975 2822
rect 48671 2642 48727 2698
rect 48795 2642 48851 2698
rect 48919 2642 48975 2698
rect 48671 2518 48727 2574
rect 48795 2518 48851 2574
rect 48919 2518 48975 2574
rect 57381 3781 57437 3837
rect 57593 3781 57649 3837
rect 57381 3563 57437 3619
rect 57593 3563 57649 3619
rect 57996 33302 58052 33358
rect 58208 33302 58264 33358
rect 57996 33084 58052 33140
rect 58208 33084 58264 33140
rect 57996 32866 58052 32922
rect 58208 32866 58264 32922
rect 57996 32649 58052 32705
rect 58208 32649 58264 32705
rect 57996 32431 58052 32487
rect 58208 32431 58264 32487
rect 57996 32075 57998 32088
rect 57998 32075 58050 32088
rect 58050 32075 58052 32088
rect 57996 32032 58052 32075
rect 58208 32075 58210 32088
rect 58210 32075 58262 32088
rect 58262 32075 58264 32088
rect 58208 32032 58264 32075
rect 57996 31857 57998 31870
rect 57998 31857 58050 31870
rect 58050 31857 58052 31870
rect 57996 31814 58052 31857
rect 58208 31857 58210 31870
rect 58210 31857 58262 31870
rect 58262 31857 58264 31870
rect 58208 31814 58264 31857
rect 57996 31639 57998 31652
rect 57998 31639 58050 31652
rect 58050 31639 58052 31652
rect 57996 31596 58052 31639
rect 58208 31639 58210 31652
rect 58210 31639 58262 31652
rect 58262 31639 58264 31652
rect 58208 31596 58264 31639
rect 57996 29950 58052 29968
rect 57996 29912 57998 29950
rect 57998 29912 58050 29950
rect 58050 29912 58052 29950
rect 58208 29950 58264 29968
rect 58208 29912 58210 29950
rect 58210 29912 58262 29950
rect 58262 29912 58264 29950
rect 57996 29733 58052 29750
rect 57996 29694 57998 29733
rect 57998 29694 58050 29733
rect 58050 29694 58052 29733
rect 58208 29733 58264 29750
rect 58208 29694 58210 29733
rect 58210 29694 58262 29733
rect 58262 29694 58264 29733
rect 57996 29515 58052 29533
rect 57996 29477 57998 29515
rect 57998 29477 58050 29515
rect 58050 29477 58052 29515
rect 58208 29515 58264 29533
rect 58208 29477 58210 29515
rect 58210 29477 58262 29515
rect 58262 29477 58264 29515
rect 57996 29297 58052 29315
rect 57996 29259 57998 29297
rect 57998 29259 58050 29297
rect 58050 29259 58052 29297
rect 58208 29297 58264 29315
rect 58208 29259 58210 29297
rect 58210 29259 58262 29297
rect 58262 29259 58264 29297
rect 57996 29080 58052 29098
rect 57996 29042 57998 29080
rect 57998 29042 58050 29080
rect 58050 29042 58052 29080
rect 58208 29080 58264 29098
rect 58208 29042 58210 29080
rect 58210 29042 58262 29080
rect 58262 29042 58264 29080
rect 57996 28862 58052 28880
rect 57996 28824 57998 28862
rect 57998 28824 58050 28862
rect 58050 28824 58052 28862
rect 58208 28862 58264 28880
rect 58208 28824 58210 28862
rect 58210 28824 58262 28862
rect 58262 28824 58264 28862
rect 57996 28644 58052 28662
rect 57996 28606 57998 28644
rect 57998 28606 58050 28644
rect 58050 28606 58052 28644
rect 58208 28644 58264 28662
rect 58208 28606 58210 28644
rect 58210 28606 58262 28644
rect 58262 28606 58264 28644
rect 57996 28427 58052 28444
rect 57996 28388 57998 28427
rect 57998 28388 58050 28427
rect 58050 28388 58052 28427
rect 58208 28427 58264 28444
rect 58208 28388 58210 28427
rect 58210 28388 58262 28427
rect 58262 28388 58264 28427
rect 57996 28209 58052 28227
rect 57996 28171 57998 28209
rect 57998 28171 58050 28209
rect 58050 28171 58052 28209
rect 58208 28209 58264 28227
rect 58208 28171 58210 28209
rect 58210 28171 58262 28209
rect 58262 28171 58264 28209
rect 57996 27992 58052 28009
rect 57996 27953 57998 27992
rect 57998 27953 58050 27992
rect 58050 27953 58052 27992
rect 58208 27992 58264 28009
rect 58208 27953 58210 27992
rect 58210 27953 58262 27992
rect 58262 27953 58264 27992
rect 57996 27774 58052 27792
rect 57996 27736 57998 27774
rect 57998 27736 58050 27774
rect 58050 27736 58052 27774
rect 58208 27774 58264 27792
rect 58208 27736 58210 27774
rect 58210 27736 58262 27774
rect 58262 27736 58264 27774
rect 57996 27556 58052 27574
rect 57996 27518 57998 27556
rect 57998 27518 58050 27556
rect 58050 27518 58052 27556
rect 58208 27556 58264 27574
rect 58208 27518 58210 27556
rect 58210 27518 58262 27556
rect 58262 27518 58264 27556
rect 58876 51527 58878 51572
rect 58878 51527 58930 51572
rect 58930 51527 58932 51572
rect 58876 51516 58932 51527
rect 59000 51527 59002 51572
rect 59002 51527 59054 51572
rect 59054 51527 59056 51572
rect 59000 51516 59056 51527
rect 59124 51527 59126 51572
rect 59126 51527 59178 51572
rect 59178 51527 59180 51572
rect 59124 51516 59180 51527
rect 59248 51527 59250 51572
rect 59250 51527 59302 51572
rect 59302 51527 59304 51572
rect 59248 51516 59304 51527
rect 59372 51527 59374 51572
rect 59374 51527 59426 51572
rect 59426 51527 59428 51572
rect 59372 51516 59428 51527
rect 58876 51403 58878 51448
rect 58878 51403 58930 51448
rect 58930 51403 58932 51448
rect 58876 51392 58932 51403
rect 59000 51403 59002 51448
rect 59002 51403 59054 51448
rect 59054 51403 59056 51448
rect 59000 51392 59056 51403
rect 59124 51403 59126 51448
rect 59126 51403 59178 51448
rect 59178 51403 59180 51448
rect 59124 51392 59180 51403
rect 59248 51403 59250 51448
rect 59250 51403 59302 51448
rect 59302 51403 59304 51448
rect 59248 51392 59304 51403
rect 59372 51403 59374 51448
rect 59374 51403 59426 51448
rect 59426 51403 59428 51448
rect 59372 51392 59428 51403
rect 58876 51279 58878 51324
rect 58878 51279 58930 51324
rect 58930 51279 58932 51324
rect 58876 51268 58932 51279
rect 59000 51279 59002 51324
rect 59002 51279 59054 51324
rect 59054 51279 59056 51324
rect 59000 51268 59056 51279
rect 59124 51279 59126 51324
rect 59126 51279 59178 51324
rect 59178 51279 59180 51324
rect 59124 51268 59180 51279
rect 59248 51279 59250 51324
rect 59250 51279 59302 51324
rect 59302 51279 59304 51324
rect 59248 51268 59304 51279
rect 59372 51279 59374 51324
rect 59374 51279 59426 51324
rect 59426 51279 59428 51324
rect 59372 51268 59428 51279
rect 58873 35188 58929 35244
rect 58997 35188 59053 35244
rect 59121 35188 59177 35244
rect 59245 35188 59301 35244
rect 59369 35188 59425 35244
rect 58873 35064 58929 35120
rect 58997 35064 59053 35120
rect 59121 35064 59177 35120
rect 59245 35064 59301 35120
rect 59369 35064 59425 35120
rect 58873 34940 58929 34996
rect 58997 34940 59053 34996
rect 59121 34940 59177 34996
rect 59245 34940 59301 34996
rect 59369 34940 59425 34996
rect 58873 34816 58929 34872
rect 58997 34816 59053 34872
rect 59121 34816 59177 34872
rect 59245 34816 59301 34872
rect 59369 34816 59425 34872
rect 58873 34692 58929 34748
rect 58997 34692 59053 34748
rect 59121 34692 59177 34748
rect 59245 34692 59301 34748
rect 59369 34692 59425 34748
rect 58873 34568 58929 34624
rect 58997 34568 59053 34624
rect 59121 34568 59177 34624
rect 59245 34568 59301 34624
rect 59369 34568 59425 34624
rect 58873 31242 58929 31298
rect 58997 31242 59053 31298
rect 59121 31242 59177 31298
rect 59245 31242 59301 31298
rect 59369 31242 59425 31298
rect 58873 31118 58929 31174
rect 58997 31118 59053 31174
rect 59121 31118 59177 31174
rect 59245 31118 59301 31174
rect 59369 31118 59425 31174
rect 58873 30994 58929 31050
rect 58997 30994 59053 31050
rect 59121 30994 59177 31050
rect 59245 30994 59301 31050
rect 59369 30994 59425 31050
rect 58873 30797 58929 30853
rect 58997 30797 59053 30853
rect 59121 30797 59177 30853
rect 59245 30797 59301 30853
rect 59369 30797 59425 30853
rect 58873 30673 58929 30729
rect 58997 30673 59053 30729
rect 59121 30673 59177 30729
rect 59245 30673 59301 30729
rect 59369 30673 59425 30729
rect 58873 30549 58929 30605
rect 58997 30549 59053 30605
rect 59121 30549 59177 30605
rect 59245 30549 59301 30605
rect 59369 30549 59425 30605
rect 58859 28268 58915 28324
rect 58983 28268 59039 28324
rect 59107 28268 59163 28324
rect 59231 28268 59287 28324
rect 59355 28268 59411 28324
rect 58859 28144 58915 28200
rect 58983 28144 59039 28200
rect 59107 28144 59163 28200
rect 59231 28144 59287 28200
rect 59355 28144 59411 28200
rect 58859 28020 58915 28076
rect 58983 28020 59039 28076
rect 59107 28020 59163 28076
rect 59231 28020 59287 28076
rect 59355 28020 59411 28076
rect 58859 27896 58915 27952
rect 58983 27896 59039 27952
rect 59107 27896 59163 27952
rect 59231 27896 59287 27952
rect 59355 27896 59411 27952
rect 58859 27772 58915 27828
rect 58983 27772 59039 27828
rect 59107 27772 59163 27828
rect 59231 27772 59287 27828
rect 59355 27772 59411 27828
rect 58859 27648 58915 27704
rect 58983 27648 59039 27704
rect 59107 27648 59163 27704
rect 59231 27648 59287 27704
rect 59355 27648 59411 27704
rect 58859 27524 58915 27580
rect 58983 27524 59039 27580
rect 59107 27524 59163 27580
rect 59231 27524 59287 27580
rect 59355 27524 59411 27580
rect 58859 27400 58915 27456
rect 58983 27400 59039 27456
rect 59107 27400 59163 27456
rect 59231 27400 59287 27456
rect 59355 27400 59411 27456
rect 58859 27276 58915 27332
rect 58983 27276 59039 27332
rect 59107 27276 59163 27332
rect 59231 27276 59287 27332
rect 59355 27276 59411 27332
rect 58859 27152 58915 27208
rect 58983 27152 59039 27208
rect 59107 27152 59163 27208
rect 59231 27152 59287 27208
rect 59355 27152 59411 27208
rect 58859 27028 58915 27084
rect 58983 27028 59039 27084
rect 59107 27028 59163 27084
rect 59231 27028 59287 27084
rect 59355 27028 59411 27084
rect 58859 26904 58915 26960
rect 58983 26904 59039 26960
rect 59107 26904 59163 26960
rect 59231 26904 59287 26960
rect 59355 26904 59411 26960
rect 58859 26780 58915 26836
rect 58983 26780 59039 26836
rect 59107 26780 59163 26836
rect 59231 26780 59287 26836
rect 59355 26780 59411 26836
rect 58859 26656 58915 26712
rect 58983 26656 59039 26712
rect 59107 26656 59163 26712
rect 59231 26656 59287 26712
rect 59355 26656 59411 26712
rect 58859 26532 58915 26588
rect 58983 26532 59039 26588
rect 59107 26532 59163 26588
rect 59231 26532 59287 26588
rect 59355 26532 59411 26588
rect 57994 24074 58258 24075
rect 57994 24022 57998 24074
rect 57998 24022 58050 24074
rect 58050 24022 58210 24074
rect 58210 24022 58258 24074
rect 57994 23857 58258 24022
rect 57994 23805 57998 23857
rect 57998 23805 58050 23857
rect 58050 23805 58210 23857
rect 58210 23805 58258 23857
rect 57994 23639 58258 23805
rect 57994 23587 57998 23639
rect 57998 23587 58050 23639
rect 58050 23587 58210 23639
rect 58210 23587 58258 23639
rect 57994 23421 58258 23587
rect 57994 23369 57998 23421
rect 57998 23369 58050 23421
rect 58050 23369 58210 23421
rect 58210 23369 58258 23421
rect 57994 23204 58258 23369
rect 57994 23187 57998 23204
rect 57998 23187 58050 23204
rect 58050 23187 58210 23204
rect 58210 23187 58258 23204
rect 58048 20540 58050 20570
rect 58050 20540 58208 20570
rect 58048 20410 58208 20540
rect 58048 20157 58208 20226
rect 58048 20105 58050 20157
rect 58050 20105 58208 20157
rect 58048 20066 58208 20105
rect 57996 13734 58052 13790
rect 58208 13734 58264 13790
rect 57996 13517 58052 13573
rect 58208 13517 58264 13573
rect 57996 13299 58052 13355
rect 58208 13299 58264 13355
rect 57996 13082 58052 13138
rect 58208 13082 58264 13138
rect 57996 12864 58052 12920
rect 58208 12864 58264 12920
rect 57996 12646 58052 12702
rect 58208 12646 58264 12702
rect 57996 12428 58052 12484
rect 58208 12428 58264 12484
rect 57996 12211 58052 12267
rect 58208 12211 58264 12267
rect 57996 11993 58052 12049
rect 58208 11993 58264 12049
rect 57996 11776 58052 11832
rect 58208 11776 58264 11832
rect 57996 9351 58052 9407
rect 58208 9351 58264 9407
rect 57996 9134 58052 9190
rect 58208 9134 58264 9190
rect 57996 8916 58052 8972
rect 58208 8916 58264 8972
rect 57996 8698 58052 8754
rect 58208 8698 58264 8754
rect 57996 8480 58052 8536
rect 58208 8480 58264 8536
rect 57996 8263 58052 8319
rect 58208 8263 58264 8319
rect 57996 5523 57998 5539
rect 57998 5523 58050 5539
rect 58050 5523 58052 5539
rect 57996 5483 58052 5523
rect 58208 5523 58210 5539
rect 58210 5523 58262 5539
rect 58262 5523 58264 5539
rect 58208 5483 58264 5523
rect 57996 5306 57998 5321
rect 57998 5306 58050 5321
rect 58050 5306 58052 5321
rect 57996 5265 58052 5306
rect 58208 5306 58210 5321
rect 58210 5306 58262 5321
rect 58262 5306 58264 5321
rect 58208 5265 58264 5306
rect 57996 4472 58052 4528
rect 58208 4472 58264 4528
rect 57996 4254 58052 4310
rect 58208 4254 58264 4310
rect 49161 2143 49217 2199
rect 49285 2143 49341 2199
rect 49409 2143 49465 2199
rect 49161 2019 49217 2075
rect 49285 2019 49341 2075
rect 49409 2019 49465 2075
rect 49161 1895 49217 1951
rect 49285 1895 49341 1951
rect 49409 1895 49465 1951
rect 49161 1771 49217 1827
rect 49285 1771 49341 1827
rect 49409 1771 49465 1827
rect 49161 1647 49217 1703
rect 49285 1647 49341 1703
rect 49409 1647 49465 1703
rect 49161 1523 49217 1579
rect 49285 1523 49341 1579
rect 49409 1523 49465 1579
rect 49161 1399 49217 1455
rect 49285 1399 49341 1455
rect 49409 1399 49465 1455
rect 49161 1275 49217 1331
rect 49285 1275 49341 1331
rect 49409 1275 49465 1331
<< metal3 >>
rect 1401 52976 2401 53776
rect 2626 53168 3626 53776
rect 4137 52976 5137 53776
rect 5362 53168 6362 53776
rect 6801 52976 7801 53776
rect 8026 53168 9026 53776
rect 9537 52976 10537 53776
rect 10762 53168 11762 53776
rect 12201 52976 13201 53776
rect 13426 53168 14426 53776
rect 14937 52976 15937 53776
rect 16162 53168 17162 53776
rect 17601 52976 18601 53776
rect 18826 53168 19826 53776
rect 20653 52976 21653 53776
rect 22258 53168 23258 53776
rect 23483 52976 24483 53776
rect 25158 53168 26158 53776
rect 26572 52976 27572 53776
rect 27877 53168 28877 53776
rect 29273 53168 30273 53776
rect 30710 52976 31710 53776
rect 32381 53168 33381 53776
rect 34024 53168 35024 53776
rect 35415 52976 36415 53776
rect 36948 53168 37948 53776
rect 38585 52976 39585 53776
rect 39882 53168 40882 53776
rect 41230 52976 42230 53776
rect 42430 53168 43430 53776
rect 43713 53168 44713 53776
rect 45069 52976 46069 53776
rect 46313 52976 47313 53776
rect 47538 53168 48538 53776
rect 48901 52976 49901 53776
rect 50465 53168 51465 53776
rect 52569 52976 53569 53776
rect 54262 52976 55262 53776
rect 55990 53168 56990 53776
rect 57547 52976 58547 53776
rect 58791 53168 59791 53776
rect 60977 52976 61977 53776
rect 62202 53168 63202 53776
rect 63713 52976 64713 53776
rect 64938 53168 65938 53776
rect 66377 52976 67377 53776
rect 67602 53168 68602 53776
rect 69113 52976 70113 53776
rect 70338 53168 71338 53776
rect 71777 52976 72777 53776
rect 73002 53168 74002 53776
rect 74513 52976 75513 53776
rect 75738 53168 76738 53776
rect 77177 52976 78177 53776
rect 78402 53168 79402 53776
rect 80229 52976 81229 53776
rect 81834 53168 82834 53776
rect 83059 52976 84059 53776
rect 84666 52976 85666 53776
rect 0 51976 86372 52976
rect 0 51626 1014 51776
rect 0 51572 27779 51626
rect 0 51516 25398 51572
rect 25454 51516 25522 51572
rect 25578 51516 25646 51572
rect 25702 51516 25770 51572
rect 25826 51516 25894 51572
rect 25950 51528 27779 51572
rect 58791 51576 59517 51591
rect 85358 51576 86372 51776
rect 58791 51572 86372 51576
rect 58791 51528 58876 51572
rect 25950 51516 58876 51528
rect 58932 51516 59000 51572
rect 59056 51516 59124 51572
rect 59180 51516 59248 51572
rect 59304 51516 59372 51572
rect 59428 51516 86372 51572
rect 0 51455 86372 51516
rect 0 51448 27788 51455
rect 0 51392 25398 51448
rect 25454 51392 25522 51448
rect 25578 51392 25646 51448
rect 25702 51392 25770 51448
rect 25826 51392 25894 51448
rect 25950 51399 27788 51448
rect 27844 51399 27999 51455
rect 28055 51399 28210 51455
rect 28266 51399 28421 51455
rect 28477 51399 28632 51455
rect 28688 51399 28843 51455
rect 28899 51399 29054 51455
rect 29110 51399 56013 51455
rect 56069 51399 56224 51455
rect 56280 51399 56435 51455
rect 56491 51399 56646 51455
rect 56702 51399 56857 51455
rect 56913 51399 57068 51455
rect 57124 51399 57279 51455
rect 57335 51448 86372 51455
rect 57335 51399 58876 51448
rect 25950 51392 58876 51399
rect 58932 51392 59000 51448
rect 59056 51392 59124 51448
rect 59180 51392 59248 51448
rect 59304 51392 59372 51448
rect 59428 51392 86372 51448
rect 0 51327 86372 51392
rect 0 51324 27779 51327
rect 30402 51326 54622 51327
rect 0 51268 25398 51324
rect 25454 51268 25522 51324
rect 25578 51268 25646 51324
rect 25702 51268 25770 51324
rect 25826 51268 25894 51324
rect 25950 51268 27779 51324
rect 0 51226 27779 51268
rect 58791 51324 86372 51327
rect 58791 51268 58876 51324
rect 58932 51268 59000 51324
rect 59056 51268 59124 51324
rect 59180 51268 59248 51324
rect 59304 51268 59372 51324
rect 59428 51276 86372 51324
rect 59428 51268 59517 51276
rect 58791 51258 59517 51268
rect 0 51076 1014 51226
rect 85358 51076 86372 51276
rect 0 50176 1706 50876
rect 56271 50866 61644 51068
rect 41865 50613 42045 50623
rect 41865 50453 41875 50613
rect 42035 50453 42045 50613
rect 41865 50443 42045 50453
rect 84666 50176 86372 50876
rect 0 49776 1014 49976
rect 85358 49776 86372 49976
rect 0 49726 27272 49776
rect 30403 49726 54622 49728
rect 59421 49726 86372 49776
rect 0 49655 86372 49726
rect 0 49599 27788 49655
rect 27844 49599 27999 49655
rect 28055 49599 28210 49655
rect 28266 49599 28421 49655
rect 28477 49599 28632 49655
rect 28688 49599 28843 49655
rect 28899 49599 29054 49655
rect 29110 49599 56013 49655
rect 56069 49599 56224 49655
rect 56280 49599 56435 49655
rect 56491 49599 56646 49655
rect 56702 49599 56857 49655
rect 56913 49599 57068 49655
rect 57124 49599 57279 49655
rect 57335 49599 86372 49655
rect 0 49526 86372 49599
rect 0 49476 27272 49526
rect 59421 49476 86372 49526
rect 0 49276 1014 49476
rect 85358 49276 86372 49476
rect 0 48376 1706 49076
rect 84666 48376 86372 49076
rect 0 47976 1014 48176
rect 85358 47976 86372 48176
rect 0 47926 27272 47976
rect 30403 47926 54622 47928
rect 59421 47926 86372 47976
rect 0 47855 86372 47926
rect 0 47799 27788 47855
rect 27844 47799 27999 47855
rect 28055 47799 28210 47855
rect 28266 47799 28421 47855
rect 28477 47799 28632 47855
rect 28688 47799 28843 47855
rect 28899 47799 29054 47855
rect 29110 47799 56013 47855
rect 56069 47799 56224 47855
rect 56280 47799 56435 47855
rect 56491 47799 56646 47855
rect 56702 47799 56857 47855
rect 56913 47799 57068 47855
rect 57124 47799 57279 47855
rect 57335 47799 86372 47855
rect 0 47726 86372 47799
rect 0 47676 27272 47726
rect 59421 47676 86372 47726
rect 0 47476 1014 47676
rect 85358 47476 86372 47676
rect 0 46576 1706 47276
rect 84666 46576 86372 47276
rect 0 46176 1014 46376
rect 85358 46176 86372 46376
rect 0 46126 27272 46176
rect 30403 46126 54622 46128
rect 59421 46126 86372 46176
rect 0 46055 86372 46126
rect 0 45999 27788 46055
rect 27844 45999 27999 46055
rect 28055 45999 28210 46055
rect 28266 45999 28421 46055
rect 28477 45999 28632 46055
rect 28688 45999 28843 46055
rect 28899 45999 29054 46055
rect 29110 45999 56013 46055
rect 56069 45999 56224 46055
rect 56280 45999 56435 46055
rect 56491 45999 56646 46055
rect 56702 45999 56857 46055
rect 56913 45999 57068 46055
rect 57124 45999 57279 46055
rect 57335 45999 86372 46055
rect 0 45926 86372 45999
rect 0 45876 27272 45926
rect 59421 45876 86372 45926
rect 0 45676 1014 45876
rect 85358 45676 86372 45876
rect 0 44776 1706 45476
rect 84666 44776 86372 45476
rect 0 44376 1014 44576
rect 85358 44376 86372 44576
rect 0 44326 27272 44376
rect 30403 44326 54622 44328
rect 59421 44326 86372 44376
rect 0 44255 86372 44326
rect 0 44199 27788 44255
rect 27844 44199 27999 44255
rect 28055 44199 28210 44255
rect 28266 44199 28421 44255
rect 28477 44199 28632 44255
rect 28688 44199 28843 44255
rect 28899 44199 29054 44255
rect 29110 44199 56013 44255
rect 56069 44199 56224 44255
rect 56280 44199 56435 44255
rect 56491 44199 56646 44255
rect 56702 44199 56857 44255
rect 56913 44199 57068 44255
rect 57124 44199 57279 44255
rect 57335 44199 86372 44255
rect 0 44126 86372 44199
rect 0 44076 27272 44126
rect 59421 44076 86372 44126
rect 0 43876 1014 44076
rect 85358 43876 86372 44076
rect 0 42976 1706 43676
rect 84666 42976 86372 43676
rect 0 42576 1014 42776
rect 85358 42576 86372 42776
rect 0 42526 27272 42576
rect 30403 42526 54622 42528
rect 59421 42526 86372 42576
rect 0 42455 86372 42526
rect 0 42399 27788 42455
rect 27844 42399 27999 42455
rect 28055 42399 28210 42455
rect 28266 42399 28421 42455
rect 28477 42399 28632 42455
rect 28688 42399 28843 42455
rect 28899 42399 29054 42455
rect 29110 42399 56013 42455
rect 56069 42399 56224 42455
rect 56280 42399 56435 42455
rect 56491 42399 56646 42455
rect 56702 42399 56857 42455
rect 56913 42399 57068 42455
rect 57124 42399 57279 42455
rect 57335 42399 86372 42455
rect 0 42326 86372 42399
rect 0 42276 27272 42326
rect 59421 42276 86372 42326
rect 0 42076 1014 42276
rect 85358 42076 86372 42276
rect 0 41176 1706 41876
rect 84666 41176 86372 41876
rect 0 40776 1014 40976
rect 85358 40776 86372 40976
rect 0 40726 27272 40776
rect 30403 40726 54622 40728
rect 59421 40726 86372 40776
rect 0 40655 86372 40726
rect 0 40599 27788 40655
rect 27844 40599 27999 40655
rect 28055 40599 28210 40655
rect 28266 40599 28421 40655
rect 28477 40599 28632 40655
rect 28688 40599 28843 40655
rect 28899 40599 29054 40655
rect 29110 40599 56013 40655
rect 56069 40599 56224 40655
rect 56280 40599 56435 40655
rect 56491 40599 56646 40655
rect 56702 40599 56857 40655
rect 56913 40599 57068 40655
rect 57124 40599 57279 40655
rect 57335 40599 86372 40655
rect 0 40526 86372 40599
rect 0 40476 27272 40526
rect 59421 40476 86372 40526
rect 0 40276 1014 40476
rect 85358 40276 86372 40476
rect 0 39376 1706 40076
rect 84666 39376 86372 40076
rect 0 38976 1014 39176
rect 85358 38976 86372 39176
rect 0 38926 27272 38976
rect 30403 38926 54622 38928
rect 59421 38926 86372 38976
rect 0 38855 86372 38926
rect 0 38799 27788 38855
rect 27844 38799 27999 38855
rect 28055 38799 28210 38855
rect 28266 38799 28421 38855
rect 28477 38799 28632 38855
rect 28688 38799 28843 38855
rect 28899 38799 29054 38855
rect 29110 38799 56013 38855
rect 56069 38799 56224 38855
rect 56280 38799 56435 38855
rect 56491 38799 56646 38855
rect 56702 38799 56857 38855
rect 56913 38799 57068 38855
rect 57124 38799 57279 38855
rect 57335 38799 86372 38855
rect 0 38726 86372 38799
rect 0 38676 27272 38726
rect 59421 38676 86372 38726
rect 0 38476 1014 38676
rect 85358 38476 86372 38676
rect 0 37576 1706 38276
rect 84666 37576 86372 38276
rect 0 37176 1014 37376
rect 85358 37176 86372 37376
rect 0 37126 27272 37176
rect 30403 37126 54622 37128
rect 59421 37126 86372 37176
rect 0 37055 86372 37126
rect 0 36999 27788 37055
rect 27844 36999 27999 37055
rect 28055 36999 28210 37055
rect 28266 36999 28421 37055
rect 28477 36999 28632 37055
rect 28688 36999 28843 37055
rect 28899 36999 29054 37055
rect 29110 36999 56013 37055
rect 56069 36999 56224 37055
rect 56280 36999 56435 37055
rect 56491 36999 56646 37055
rect 56702 36999 56857 37055
rect 56913 36999 57068 37055
rect 57124 36999 57279 37055
rect 57335 36999 86372 37055
rect 0 36926 86372 36999
rect 0 36876 27272 36926
rect 59421 36876 86372 36926
rect 0 36676 1014 36876
rect 85358 36676 86372 36876
rect 0 35776 1706 36476
rect 36863 35881 37743 35920
rect 36863 35825 36958 35881
rect 37014 35825 37169 35881
rect 37225 35825 37381 35881
rect 37437 35825 37592 35881
rect 37648 35825 37743 35881
rect 0 35275 27828 35326
rect 0 35219 25384 35275
rect 25440 35219 25508 35275
rect 25564 35219 25632 35275
rect 25688 35219 25756 35275
rect 25812 35219 25880 35275
rect 25936 35219 27438 35275
rect 27494 35219 27562 35275
rect 27618 35219 27686 35275
rect 27742 35219 27828 35275
rect 0 35151 27828 35219
rect 0 35095 25384 35151
rect 25440 35095 25508 35151
rect 25564 35095 25632 35151
rect 25688 35095 25756 35151
rect 25812 35095 25880 35151
rect 25936 35095 27438 35151
rect 27494 35095 27562 35151
rect 27618 35095 27686 35151
rect 27742 35095 27828 35151
rect 0 35027 27828 35095
rect 0 34971 25384 35027
rect 25440 34971 25508 35027
rect 25564 34971 25632 35027
rect 25688 34971 25756 35027
rect 25812 34971 25880 35027
rect 25936 34971 27438 35027
rect 27494 34971 27562 35027
rect 27618 34971 27686 35027
rect 27742 34971 27828 35027
rect 0 34903 27828 34971
rect 0 34847 25384 34903
rect 25440 34847 25508 34903
rect 25564 34847 25632 34903
rect 25688 34847 25756 34903
rect 25812 34847 25880 34903
rect 25936 34847 27438 34903
rect 27494 34847 27562 34903
rect 27618 34847 27686 34903
rect 27742 34847 27828 34903
rect 0 34779 27828 34847
rect 0 34723 25384 34779
rect 25440 34723 25508 34779
rect 25564 34723 25632 34779
rect 25688 34723 25756 34779
rect 25812 34723 25880 34779
rect 25936 34723 27438 34779
rect 27494 34723 27562 34779
rect 27618 34723 27686 34779
rect 27742 34723 27828 34779
rect 0 34655 27828 34723
rect 0 34599 25384 34655
rect 25440 34599 25508 34655
rect 25564 34599 25632 34655
rect 25688 34599 25756 34655
rect 25812 34599 25880 34655
rect 25936 34599 27438 34655
rect 27494 34599 27562 34655
rect 27618 34599 27686 34655
rect 27742 34599 27828 34655
rect 0 34536 27828 34599
rect 2095 34125 2188 34126
rect 0 34124 25085 34125
rect 0 34011 27214 34124
rect 0 33955 26859 34011
rect 26915 33955 27071 34011
rect 27127 33955 27214 34011
rect 0 33793 27214 33955
rect 36863 33927 37743 35825
rect 84666 35776 86372 36476
rect 57369 35244 86372 35326
rect 57369 35188 58873 35244
rect 58929 35188 58997 35244
rect 59053 35188 59121 35244
rect 59177 35188 59245 35244
rect 59301 35188 59369 35244
rect 59425 35188 86372 35244
rect 57369 35120 86372 35188
rect 57369 35064 58873 35120
rect 58929 35064 58997 35120
rect 59053 35064 59121 35120
rect 59177 35064 59245 35120
rect 59301 35064 59369 35120
rect 59425 35064 86372 35120
rect 57369 34996 86372 35064
rect 57369 34940 58873 34996
rect 58929 34940 58997 34996
rect 59053 34940 59121 34996
rect 59177 34940 59245 34996
rect 59301 34940 59369 34996
rect 59425 34940 86372 34996
rect 57369 34872 86372 34940
rect 57369 34816 58873 34872
rect 58929 34816 58997 34872
rect 59053 34816 59121 34872
rect 59177 34816 59245 34872
rect 59301 34816 59369 34872
rect 59425 34816 86372 34872
rect 57369 34748 86372 34816
rect 57369 34692 58873 34748
rect 58929 34692 58997 34748
rect 59053 34692 59121 34748
rect 59177 34692 59245 34748
rect 59301 34692 59369 34748
rect 59425 34692 86372 34748
rect 57369 34624 86372 34692
rect 57369 34568 58873 34624
rect 58929 34568 58997 34624
rect 59053 34568 59121 34624
rect 59177 34568 59245 34624
rect 59301 34568 59369 34624
rect 59425 34568 86372 34624
rect 57369 34536 86372 34568
rect 61853 34124 72383 34125
rect 72653 34124 86372 34125
rect 57908 34011 86372 34124
rect 57908 33955 57996 34011
rect 58052 33955 58208 34011
rect 58264 33955 86372 34011
rect 0 33737 26859 33793
rect 26915 33737 27071 33793
rect 27127 33737 27214 33793
rect 0 33576 27214 33737
rect 0 33520 26859 33576
rect 26915 33520 27071 33576
rect 27127 33520 27214 33576
rect 0 33358 27214 33520
rect 0 33302 26859 33358
rect 26915 33302 27071 33358
rect 27127 33302 27214 33358
rect 0 33140 27214 33302
rect 57908 33793 86372 33955
rect 57908 33737 57996 33793
rect 58052 33737 58208 33793
rect 58264 33737 86372 33793
rect 57908 33576 86372 33737
rect 57908 33520 57996 33576
rect 58052 33520 58208 33576
rect 58264 33520 86372 33576
rect 57908 33358 86372 33520
rect 57908 33302 57996 33358
rect 58052 33302 58208 33358
rect 58264 33302 86372 33358
rect 0 33084 26859 33140
rect 26915 33084 27071 33140
rect 27127 33084 27214 33140
rect 0 32922 27214 33084
rect 0 32866 26859 32922
rect 26915 32866 27071 32922
rect 27127 32866 27214 32922
rect 0 32705 27214 32866
rect 0 32649 26859 32705
rect 26915 32649 27071 32705
rect 27127 32649 27214 32705
rect 0 32487 27214 32649
rect 0 32431 26859 32487
rect 26915 32431 27071 32487
rect 27127 32431 27214 32487
rect 0 32318 27214 32431
rect 27387 33141 28929 33263
rect 27387 33085 27474 33141
rect 27530 33085 27686 33141
rect 27742 33085 28929 33141
rect 27387 32923 28929 33085
rect 27387 32867 27474 32923
rect 27530 32867 27686 32923
rect 27742 32867 28929 32923
rect 27387 32705 28929 32867
rect 27387 32649 27474 32705
rect 27530 32649 27686 32705
rect 27742 32649 28929 32705
rect 27387 32487 28929 32649
rect 27387 32431 27474 32487
rect 27530 32431 27686 32487
rect 27742 32431 28929 32487
rect 0 32316 25085 32318
rect 0 32315 3011 32316
rect 0 29714 1706 32315
rect 27387 32311 28929 32431
rect 56135 33141 57736 33263
rect 56135 33085 57381 33141
rect 57437 33085 57593 33141
rect 57649 33085 57736 33141
rect 56135 32923 57736 33085
rect 56135 32867 57381 32923
rect 57437 32867 57593 32923
rect 57649 32867 57736 32923
rect 56135 32705 57736 32867
rect 56135 32649 57381 32705
rect 57437 32649 57593 32705
rect 57649 32649 57736 32705
rect 56135 32487 57736 32649
rect 56135 32431 57381 32487
rect 57437 32431 57593 32487
rect 57649 32431 57736 32487
rect 56135 32311 57736 32431
rect 57908 33140 86372 33302
rect 57908 33084 57996 33140
rect 58052 33084 58208 33140
rect 58264 33084 86372 33140
rect 57908 32922 86372 33084
rect 57908 32866 57996 32922
rect 58052 32866 58208 32922
rect 58264 32866 86372 32922
rect 57908 32705 86372 32866
rect 57908 32649 57996 32705
rect 58052 32649 58208 32705
rect 58264 32649 86372 32705
rect 57908 32487 86372 32649
rect 57908 32431 57996 32487
rect 58052 32431 58208 32487
rect 58264 32431 86372 32487
rect 57908 32315 86372 32431
rect 57908 32199 58351 32315
rect 26772 32088 58351 32199
rect 26772 32032 26859 32088
rect 26915 32032 27071 32088
rect 27127 32032 57996 32088
rect 58052 32032 58208 32088
rect 58264 32032 58351 32088
rect 26772 31870 58351 32032
rect 26772 31814 26859 31870
rect 26915 31814 27071 31870
rect 27127 31814 57996 31870
rect 58052 31814 58208 31870
rect 58264 31814 58351 31870
rect 26772 31652 58351 31814
rect 26772 31596 26859 31652
rect 26915 31596 27071 31652
rect 27127 31596 57996 31652
rect 58052 31596 58208 31652
rect 58264 31596 58351 31652
rect 26772 31486 58351 31596
rect 25293 31252 28929 31352
rect 25293 31248 27474 31252
rect 25293 31192 25398 31248
rect 25454 31192 25522 31248
rect 25578 31192 25646 31248
rect 25702 31192 25770 31248
rect 25826 31192 25894 31248
rect 25950 31196 27474 31248
rect 27530 31196 27686 31252
rect 27742 31196 28929 31252
rect 25950 31192 28929 31196
rect 25293 31124 28929 31192
rect 25293 31068 25398 31124
rect 25454 31068 25522 31124
rect 25578 31068 25646 31124
rect 25702 31068 25770 31124
rect 25826 31068 25894 31124
rect 25950 31068 28929 31124
rect 25293 31034 28929 31068
rect 25293 31000 27474 31034
rect 25293 30944 25398 31000
rect 25454 30944 25522 31000
rect 25578 30944 25646 31000
rect 25702 30944 25770 31000
rect 25826 30944 25894 31000
rect 25950 30978 27474 31000
rect 27530 30978 27686 31034
rect 27742 30978 28929 31034
rect 25950 30944 28929 30978
rect 25293 30816 28929 30944
rect 25293 30793 27474 30816
rect 25293 30737 25398 30793
rect 25454 30737 25522 30793
rect 25578 30737 25646 30793
rect 25702 30737 25770 30793
rect 25826 30737 25894 30793
rect 25950 30760 27474 30793
rect 27530 30760 27686 30816
rect 27742 30760 28929 30816
rect 25950 30737 28929 30760
rect 25293 30669 28929 30737
rect 25293 30613 25398 30669
rect 25454 30613 25522 30669
rect 25578 30613 25646 30669
rect 25702 30613 25770 30669
rect 25826 30613 25894 30669
rect 25950 30613 28929 30669
rect 25293 30598 28929 30613
rect 25293 30545 27474 30598
rect 25293 30489 25398 30545
rect 25454 30489 25522 30545
rect 25578 30489 25646 30545
rect 25702 30489 25770 30545
rect 25826 30489 25894 30545
rect 25950 30542 27474 30545
rect 27530 30542 27686 30598
rect 27742 30542 28929 30598
rect 25950 30489 28929 30542
rect 25293 30443 28929 30489
rect 56186 31298 59524 31352
rect 56186 31252 58873 31298
rect 56186 31196 57381 31252
rect 57437 31196 57593 31252
rect 57649 31242 58873 31252
rect 58929 31242 58997 31298
rect 59053 31242 59121 31298
rect 59177 31242 59245 31298
rect 59301 31242 59369 31298
rect 59425 31242 59524 31298
rect 57649 31196 59524 31242
rect 56186 31174 59524 31196
rect 56186 31118 58873 31174
rect 58929 31118 58997 31174
rect 59053 31118 59121 31174
rect 59177 31118 59245 31174
rect 59301 31118 59369 31174
rect 59425 31118 59524 31174
rect 56186 31050 59524 31118
rect 56186 31034 58873 31050
rect 56186 30978 57381 31034
rect 57437 30978 57593 31034
rect 57649 30994 58873 31034
rect 58929 30994 58997 31050
rect 59053 30994 59121 31050
rect 59177 30994 59245 31050
rect 59301 30994 59369 31050
rect 59425 30994 59524 31050
rect 57649 30978 59524 30994
rect 56186 30853 59524 30978
rect 56186 30816 58873 30853
rect 56186 30760 57381 30816
rect 57437 30760 57593 30816
rect 57649 30797 58873 30816
rect 58929 30797 58997 30853
rect 59053 30797 59121 30853
rect 59177 30797 59245 30853
rect 59301 30797 59369 30853
rect 59425 30797 59524 30853
rect 57649 30760 59524 30797
rect 56186 30729 59524 30760
rect 56186 30673 58873 30729
rect 58929 30673 58997 30729
rect 59053 30673 59121 30729
rect 59177 30673 59245 30729
rect 59301 30673 59369 30729
rect 59425 30673 59524 30729
rect 56186 30605 59524 30673
rect 56186 30598 58873 30605
rect 56186 30542 57381 30598
rect 57437 30542 57593 30598
rect 57649 30549 58873 30598
rect 58929 30549 58997 30605
rect 59053 30549 59121 30605
rect 59177 30549 59245 30605
rect 59301 30549 59369 30605
rect 59425 30549 59524 30605
rect 57649 30542 59524 30549
rect 56186 30443 59524 30542
rect 26772 29968 58351 30105
rect 26772 29912 26859 29968
rect 26915 29912 27071 29968
rect 27127 29912 57996 29968
rect 58052 29912 58208 29968
rect 58264 29912 58351 29968
rect 26772 29750 58351 29912
rect 26772 29714 26859 29750
rect 0 29694 26859 29714
rect 26915 29694 27071 29750
rect 27127 29694 57996 29750
rect 58052 29694 58208 29750
rect 58264 29714 58351 29750
rect 84666 29714 86372 32315
rect 58264 29694 86372 29714
rect 0 29533 86372 29694
rect 0 29477 26859 29533
rect 26915 29477 27071 29533
rect 27127 29477 57996 29533
rect 58052 29477 58208 29533
rect 58264 29477 86372 29533
rect 0 29430 86372 29477
rect 26772 29315 58351 29430
rect 26772 29259 26859 29315
rect 26915 29259 27071 29315
rect 27127 29259 57996 29315
rect 58052 29259 58208 29315
rect 58264 29259 58351 29315
rect 26772 29098 58351 29259
rect 26772 29042 26859 29098
rect 26915 29042 27071 29098
rect 27127 29042 57996 29098
rect 58052 29042 58208 29098
rect 58264 29042 58351 29098
rect 26772 28880 58351 29042
rect 26772 28824 26859 28880
rect 26915 28824 27071 28880
rect 27127 28824 57996 28880
rect 58052 28824 58208 28880
rect 58264 28824 58351 28880
rect 26772 28662 58351 28824
rect 26772 28606 26859 28662
rect 26915 28606 27071 28662
rect 27127 28606 57996 28662
rect 58052 28606 58208 28662
rect 58264 28606 58351 28662
rect 26772 28444 58351 28606
rect 0 28263 26070 28416
rect 0 28207 25404 28263
rect 25460 28207 25528 28263
rect 25584 28207 25652 28263
rect 25708 28207 25776 28263
rect 25832 28207 25900 28263
rect 25956 28207 26070 28263
rect 0 28139 26070 28207
rect 0 28083 25404 28139
rect 25460 28083 25528 28139
rect 25584 28083 25652 28139
rect 25708 28083 25776 28139
rect 25832 28083 25900 28139
rect 25956 28083 26070 28139
rect 0 28015 26070 28083
rect 0 27959 25404 28015
rect 25460 27959 25528 28015
rect 25584 27959 25652 28015
rect 25708 27959 25776 28015
rect 25832 27959 25900 28015
rect 25956 27959 26070 28015
rect 0 27891 26070 27959
rect 0 27835 25404 27891
rect 25460 27835 25528 27891
rect 25584 27835 25652 27891
rect 25708 27835 25776 27891
rect 25832 27835 25900 27891
rect 25956 27835 26070 27891
rect 0 27767 26070 27835
rect 0 27711 25404 27767
rect 25460 27711 25528 27767
rect 25584 27711 25652 27767
rect 25708 27711 25776 27767
rect 25832 27711 25900 27767
rect 25956 27711 26070 27767
rect 0 27643 26070 27711
rect 0 27587 25404 27643
rect 25460 27587 25528 27643
rect 25584 27587 25652 27643
rect 25708 27587 25776 27643
rect 25832 27587 25900 27643
rect 25956 27587 26070 27643
rect 0 27519 26070 27587
rect 0 27463 25404 27519
rect 25460 27463 25528 27519
rect 25584 27463 25652 27519
rect 25708 27463 25776 27519
rect 25832 27463 25900 27519
rect 25956 27463 26070 27519
rect 0 27395 26070 27463
rect 0 27339 25404 27395
rect 25460 27339 25528 27395
rect 25584 27339 25652 27395
rect 25708 27339 25776 27395
rect 25832 27339 25900 27395
rect 25956 27339 26070 27395
rect 26772 28388 26859 28444
rect 26915 28388 27071 28444
rect 27127 28388 57996 28444
rect 58052 28388 58208 28444
rect 58264 28388 58351 28444
rect 26772 28227 58351 28388
rect 26772 28171 26859 28227
rect 26915 28171 27071 28227
rect 27127 28171 57996 28227
rect 58052 28171 58208 28227
rect 58264 28171 58351 28227
rect 26772 28009 58351 28171
rect 26772 27953 26859 28009
rect 26915 27953 27071 28009
rect 27127 27953 57996 28009
rect 58052 27953 58208 28009
rect 58264 27953 58351 28009
rect 26772 27792 58351 27953
rect 26772 27736 26859 27792
rect 26915 27736 27071 27792
rect 27127 27736 57996 27792
rect 58052 27736 58208 27792
rect 58264 27736 58351 27792
rect 26772 27574 58351 27736
rect 26772 27518 26859 27574
rect 26915 27518 27071 27574
rect 27127 27518 57996 27574
rect 58052 27518 58208 27574
rect 58264 27518 58351 27574
rect 26772 27382 58351 27518
rect 58785 28324 86372 28416
rect 58785 28268 58859 28324
rect 58915 28268 58983 28324
rect 59039 28268 59107 28324
rect 59163 28268 59231 28324
rect 59287 28268 59355 28324
rect 59411 28268 86372 28324
rect 58785 28200 86372 28268
rect 58785 28144 58859 28200
rect 58915 28144 58983 28200
rect 59039 28144 59107 28200
rect 59163 28144 59231 28200
rect 59287 28144 59355 28200
rect 59411 28144 86372 28200
rect 58785 28076 86372 28144
rect 58785 28020 58859 28076
rect 58915 28020 58983 28076
rect 59039 28020 59107 28076
rect 59163 28020 59231 28076
rect 59287 28020 59355 28076
rect 59411 28020 86372 28076
rect 58785 27952 86372 28020
rect 58785 27896 58859 27952
rect 58915 27896 58983 27952
rect 59039 27896 59107 27952
rect 59163 27896 59231 27952
rect 59287 27896 59355 27952
rect 59411 27896 86372 27952
rect 58785 27828 86372 27896
rect 58785 27772 58859 27828
rect 58915 27772 58983 27828
rect 59039 27772 59107 27828
rect 59163 27772 59231 27828
rect 59287 27772 59355 27828
rect 59411 27772 86372 27828
rect 58785 27704 86372 27772
rect 58785 27648 58859 27704
rect 58915 27648 58983 27704
rect 59039 27648 59107 27704
rect 59163 27648 59231 27704
rect 59287 27648 59355 27704
rect 59411 27648 86372 27704
rect 58785 27580 86372 27648
rect 58785 27524 58859 27580
rect 58915 27524 58983 27580
rect 59039 27524 59107 27580
rect 59163 27524 59231 27580
rect 59287 27524 59355 27580
rect 59411 27524 86372 27580
rect 58785 27456 86372 27524
rect 58785 27400 58859 27456
rect 58915 27400 58983 27456
rect 59039 27400 59107 27456
rect 59163 27400 59231 27456
rect 59287 27400 59355 27456
rect 59411 27400 86372 27456
rect 0 27271 26070 27339
rect 0 27215 25404 27271
rect 25460 27215 25528 27271
rect 25584 27215 25652 27271
rect 25708 27215 25776 27271
rect 25832 27215 25900 27271
rect 25956 27215 26070 27271
rect 0 27147 26070 27215
rect 0 27091 25404 27147
rect 25460 27091 25528 27147
rect 25584 27091 25652 27147
rect 25708 27091 25776 27147
rect 25832 27091 25900 27147
rect 25956 27091 26070 27147
rect 0 27023 26070 27091
rect 0 26967 25404 27023
rect 25460 26967 25528 27023
rect 25584 26967 25652 27023
rect 25708 26967 25776 27023
rect 25832 26967 25900 27023
rect 25956 26967 26070 27023
rect 0 26899 26070 26967
rect 0 26843 25404 26899
rect 25460 26843 25528 26899
rect 25584 26843 25652 26899
rect 25708 26843 25776 26899
rect 25832 26843 25900 26899
rect 25956 26890 26070 26899
rect 58785 27332 86372 27400
rect 58785 27276 58859 27332
rect 58915 27276 58983 27332
rect 59039 27276 59107 27332
rect 59163 27276 59231 27332
rect 59287 27276 59355 27332
rect 59411 27276 86372 27332
rect 58785 27208 86372 27276
rect 58785 27152 58859 27208
rect 58915 27152 58983 27208
rect 59039 27152 59107 27208
rect 59163 27152 59231 27208
rect 59287 27152 59355 27208
rect 59411 27152 86372 27208
rect 58785 27084 86372 27152
rect 58785 27028 58859 27084
rect 58915 27028 58983 27084
rect 59039 27028 59107 27084
rect 59163 27028 59231 27084
rect 59287 27028 59355 27084
rect 59411 27028 86372 27084
rect 58785 26960 86372 27028
rect 58785 26904 58859 26960
rect 58915 26904 58983 26960
rect 59039 26904 59107 26960
rect 59163 26904 59231 26960
rect 59287 26904 59355 26960
rect 59411 26904 86372 26960
rect 58785 26890 86372 26904
rect 25956 26843 27828 26890
rect 0 26799 27828 26843
rect 0 26775 27474 26799
rect 0 26719 25404 26775
rect 25460 26719 25528 26775
rect 25584 26719 25652 26775
rect 25708 26719 25776 26775
rect 25832 26719 25900 26775
rect 25956 26743 27474 26775
rect 27530 26743 27686 26799
rect 27742 26743 27828 26799
rect 25956 26719 27828 26743
rect 0 26651 27828 26719
rect 0 26595 25404 26651
rect 25460 26595 25528 26651
rect 25584 26595 25652 26651
rect 25708 26595 25776 26651
rect 25832 26595 25900 26651
rect 25956 26595 27828 26651
rect 0 26581 27828 26595
rect 0 26527 27474 26581
rect 0 26471 25404 26527
rect 25460 26471 25528 26527
rect 25584 26471 25652 26527
rect 25708 26471 25776 26527
rect 25832 26471 25900 26527
rect 25956 26525 27474 26527
rect 27530 26525 27686 26581
rect 27742 26525 27828 26581
rect 25956 26471 27828 26525
rect 0 26435 27828 26471
rect 57295 26836 86372 26890
rect 57295 26799 58859 26836
rect 57295 26743 57381 26799
rect 57437 26743 57593 26799
rect 57649 26780 58859 26799
rect 58915 26780 58983 26836
rect 59039 26780 59107 26836
rect 59163 26780 59231 26836
rect 59287 26780 59355 26836
rect 59411 26780 86372 26836
rect 57649 26743 86372 26780
rect 57295 26712 86372 26743
rect 57295 26656 58859 26712
rect 58915 26656 58983 26712
rect 59039 26656 59107 26712
rect 59163 26656 59231 26712
rect 59287 26656 59355 26712
rect 59411 26656 86372 26712
rect 57295 26588 86372 26656
rect 57295 26581 58859 26588
rect 57295 26525 57381 26581
rect 57437 26525 57593 26581
rect 57649 26532 58859 26581
rect 58915 26532 58983 26588
rect 59039 26532 59107 26588
rect 59163 26532 59231 26588
rect 59287 26532 59355 26588
rect 59411 26532 86372 26588
rect 57649 26525 86372 26532
rect 57295 26435 86372 26525
rect 6921 26434 8163 26435
rect 17721 26434 18963 26435
rect 66497 26434 67739 26435
rect 77297 26434 78539 26435
rect 23828 26286 26642 26324
rect 23828 26126 26450 26286
rect 26610 26126 26642 26286
rect 23828 26109 26642 26126
rect 23828 25967 26285 26002
rect 23828 25807 26092 25967
rect 26252 25807 26285 25967
rect 23828 25787 26285 25807
rect 23828 25647 25949 25681
rect 23828 25487 25756 25647
rect 25916 25487 25949 25647
rect 23828 25466 25949 25487
rect 23828 25328 25614 25359
rect 23828 25168 25421 25328
rect 25581 25168 25614 25328
rect 23828 25144 25614 25168
rect 27382 25028 29699 25208
rect 27382 24972 27474 25028
rect 27530 24972 27686 25028
rect 27742 24972 29699 25028
rect 27382 24810 29699 24972
rect 27382 24754 27474 24810
rect 27530 24754 27686 24810
rect 27742 24754 29699 24810
rect 23828 24637 25274 24667
rect 23828 24477 25081 24637
rect 25241 24477 25274 24637
rect 27382 24526 29699 24754
rect 23828 24452 25274 24477
rect 23828 24316 24935 24345
rect 23828 24156 24744 24316
rect 24904 24156 24935 24316
rect 23828 24130 24935 24156
rect 26770 24075 58348 24278
rect 23828 23995 24607 24024
rect 0 23380 1706 23938
rect 23828 23835 24416 23995
rect 24576 23835 24607 23995
rect 23828 23809 24607 23835
rect 24047 23673 24227 23683
rect 24047 23513 24057 23673
rect 24217 23513 24227 23673
rect 24047 23503 24227 23513
rect 26770 23380 26858 24075
rect 0 23187 26858 23380
rect 27122 23370 57994 24075
rect 27122 23187 27214 23370
rect 0 22938 27214 23187
rect 27387 22936 57677 23199
rect 57908 23187 57994 23370
rect 58258 23380 58348 24075
rect 84666 23380 86372 23938
rect 58258 23187 86372 23380
rect 57908 22938 86372 23187
rect 57908 22937 83763 22938
rect 27387 22282 27475 22936
rect 0 22048 27475 22282
rect 27739 22923 57677 22936
rect 27739 22291 57363 22923
rect 27739 22048 27826 22291
rect 0 21827 27826 22048
rect 0 21282 1014 21827
rect 24036 21826 27826 21827
rect 56078 22035 57363 22291
rect 57627 22282 57677 22923
rect 57627 22035 86372 22282
rect 56078 21827 86372 22035
rect 56078 21826 83763 21827
rect 44432 21707 55645 21708
rect 29521 21625 55645 21707
rect 29513 20739 55645 21625
rect 85358 21282 86372 21827
rect 0 20570 86372 20739
rect 0 20410 26924 20570
rect 27084 20410 58048 20570
rect 58208 20410 86372 20570
rect 0 20226 86372 20410
rect 0 20066 26924 20226
rect 27084 20066 58048 20226
rect 58208 20066 86372 20226
rect 0 19969 86372 20066
rect 0 18016 24250 19969
rect 26435 19692 29403 19731
rect 26435 19532 26465 19692
rect 26625 19532 29403 19692
rect 26435 19502 29403 19532
rect 55720 19502 58817 19731
rect 26077 19347 29403 19391
rect 26077 19187 26107 19347
rect 26267 19187 29403 19347
rect 26077 19162 29403 19187
rect 55720 19162 59177 19391
rect 25742 19027 29403 19051
rect 25742 18867 25771 19027
rect 25931 18867 29403 19027
rect 25742 18822 29403 18867
rect 55720 18822 59515 19051
rect 25406 18684 29403 18711
rect 25406 18524 25434 18684
rect 25594 18524 29403 18684
rect 25406 18482 29403 18524
rect 55720 18482 59846 18711
rect 25066 18350 29403 18371
rect 25066 18190 25094 18350
rect 25254 18190 29403 18350
rect 25066 18142 29403 18190
rect 55720 18142 60184 18371
rect 24730 17977 29403 18031
rect 24730 17817 24757 17977
rect 24917 17817 29403 17977
rect 24730 17802 29403 17817
rect 55720 17802 60525 18031
rect 61807 18016 86372 19969
rect 61825 18015 83763 18016
rect 0 16597 23678 17730
rect 24401 17656 29403 17691
rect 24401 17496 24429 17656
rect 24589 17496 29403 17656
rect 24401 17462 29403 17496
rect 55720 17462 60855 17691
rect 24042 17317 29403 17351
rect 24042 17157 24069 17317
rect 24229 17157 29403 17317
rect 24042 17122 29403 17157
rect 55720 17122 61205 17351
rect 61807 16784 86372 17730
rect 46982 16678 86372 16784
rect 46982 16622 57381 16678
rect 57437 16622 57593 16678
rect 57649 16622 86372 16678
rect 24111 16597 27828 16598
rect 0 16470 27828 16597
rect 0 16414 27474 16470
rect 27530 16414 27686 16470
rect 27742 16414 27828 16470
rect 0 16253 27828 16414
rect 0 16197 27474 16253
rect 27530 16197 27686 16253
rect 27742 16197 27828 16253
rect 0 16035 27828 16197
rect 0 15979 27474 16035
rect 27530 15979 27686 16035
rect 27742 15979 27828 16035
rect 0 15818 27828 15979
rect 0 15762 27474 15818
rect 27530 15762 27686 15818
rect 27742 15762 27828 15818
rect 0 15600 27828 15762
rect 0 15544 27474 15600
rect 27530 15544 27686 15600
rect 27742 15544 27828 15600
rect 0 15382 27828 15544
rect 0 15326 27474 15382
rect 27530 15326 27686 15382
rect 27742 15326 27828 15382
rect 0 15164 27828 15326
rect 0 15108 27474 15164
rect 27530 15108 27686 15164
rect 27742 15108 27828 15164
rect 0 15015 27828 15108
rect 46982 16461 86372 16622
rect 46982 16405 57381 16461
rect 57437 16405 57593 16461
rect 57649 16405 86372 16461
rect 46982 16243 86372 16405
rect 46982 16187 57381 16243
rect 57437 16187 57593 16243
rect 57649 16187 86372 16243
rect 46982 16026 86372 16187
rect 46982 15970 57381 16026
rect 57437 15970 57593 16026
rect 57649 15970 86372 16026
rect 46982 15808 86372 15970
rect 46982 15752 57381 15808
rect 57437 15752 57593 15808
rect 57649 15752 86372 15808
rect 46982 15590 86372 15752
rect 46982 15534 57381 15590
rect 57437 15534 57593 15590
rect 57649 15534 86372 15590
rect 46982 15372 86372 15534
rect 46982 15316 57381 15372
rect 57437 15316 57593 15372
rect 57649 15316 86372 15372
rect 46982 15155 86372 15316
rect 46982 15099 57381 15155
rect 57437 15099 57593 15155
rect 57649 15099 86372 15155
rect 46982 15015 86372 15099
rect 0 14968 86372 15015
rect 0 14966 55645 14968
rect 0 14947 51760 14966
rect 0 14891 27474 14947
rect 27530 14891 27686 14947
rect 27742 14936 51760 14947
rect 57295 14937 86372 14968
rect 27742 14891 47683 14936
rect 0 14729 47683 14891
rect 0 14673 27474 14729
rect 27530 14673 27686 14729
rect 27742 14673 47683 14729
rect 0 14512 47683 14673
rect 0 14456 27474 14512
rect 27530 14456 27686 14512
rect 27742 14491 47683 14512
rect 57295 14881 57381 14937
rect 57437 14881 57593 14937
rect 57649 14881 86372 14937
rect 57295 14720 86372 14881
rect 57295 14664 57381 14720
rect 57437 14664 57593 14720
rect 57649 14664 86372 14720
rect 27742 14456 45977 14491
rect 0 14329 45977 14456
rect 0 14328 24250 14329
rect 27387 14231 45977 14329
rect 57295 14328 86372 14664
rect 57295 14327 83763 14328
rect 24047 14178 27214 14179
rect 0 14119 27214 14178
rect 0 14063 26859 14119
rect 26915 14063 27071 14119
rect 27127 14063 27214 14119
rect 0 13902 27214 14063
rect 0 13846 26859 13902
rect 26915 13846 27071 13902
rect 27127 13846 27214 13902
rect 0 13684 27214 13846
rect 0 13628 26859 13684
rect 26915 13628 27071 13684
rect 27127 13628 27214 13684
rect 0 13467 27214 13628
rect 0 13461 26859 13467
rect 0 12846 1706 13461
rect 24047 13411 26859 13461
rect 26915 13411 27071 13467
rect 27127 13411 27214 13467
rect 24047 13249 27214 13411
rect 24047 13193 26859 13249
rect 26915 13193 27071 13249
rect 27127 13193 27214 13249
rect 27387 14175 27474 14231
rect 27530 14175 27686 14231
rect 27742 14175 45977 14231
rect 83169 14178 84221 14179
rect 61807 14177 72429 14178
rect 72607 14177 86372 14178
rect 27387 14014 45977 14175
rect 27387 13958 27474 14014
rect 27530 13958 27686 14014
rect 27742 13958 45977 14014
rect 27387 13796 45977 13958
rect 59826 13866 60026 14017
rect 61773 13866 86372 14177
rect 27387 13740 27474 13796
rect 27530 13740 27686 13796
rect 27742 13760 45977 13796
rect 50228 13790 86372 13866
rect 27742 13740 49775 13760
rect 27387 13578 49775 13740
rect 27387 13522 27474 13578
rect 27530 13522 27686 13578
rect 27742 13522 49775 13578
rect 27387 13361 49775 13522
rect 27387 13305 27474 13361
rect 27530 13305 27686 13361
rect 27742 13305 49775 13361
rect 27387 13245 49775 13305
rect 29478 13243 49775 13245
rect 24047 13031 27214 13193
rect 41493 13078 49775 13243
rect 50228 13734 57996 13790
rect 58052 13734 58208 13790
rect 58264 13734 86372 13790
rect 50228 13573 86372 13734
rect 50228 13517 57996 13573
rect 58052 13517 58208 13573
rect 58264 13517 86372 13573
rect 50228 13461 86372 13517
rect 50228 13355 58421 13461
rect 50228 13299 57996 13355
rect 58052 13299 58208 13355
rect 58264 13299 58421 13355
rect 50228 13138 58421 13299
rect 50228 13082 57996 13138
rect 58052 13082 58208 13138
rect 58264 13082 58421 13138
rect 24047 12975 26859 13031
rect 26915 12975 27071 13031
rect 27127 12975 27214 13031
rect 24047 12934 27214 12975
rect 24047 12847 34761 12934
rect 23821 12846 34761 12847
rect 0 12813 34761 12846
rect 0 12757 26859 12813
rect 26915 12757 27071 12813
rect 27127 12757 34761 12813
rect 0 12596 34761 12757
rect 0 12540 26859 12596
rect 26915 12540 27071 12596
rect 27127 12574 34761 12596
rect 50228 12920 58421 13082
rect 50228 12864 57996 12920
rect 58052 12864 58208 12920
rect 58264 12864 58421 12920
rect 50228 12846 58421 12864
rect 59826 12846 60026 13461
rect 83169 12846 84221 12847
rect 84666 12846 86372 13461
rect 50228 12702 86372 12846
rect 50228 12646 57996 12702
rect 58052 12646 58208 12702
rect 58264 12646 86372 12702
rect 50228 12574 86372 12646
rect 27127 12540 86372 12574
rect 0 12484 86372 12540
rect 0 12428 57996 12484
rect 58052 12428 58208 12484
rect 58264 12428 86372 12484
rect 0 12378 86372 12428
rect 0 12322 26859 12378
rect 26915 12322 27071 12378
rect 27127 12322 86372 12378
rect 0 12267 86372 12322
rect 0 12211 57996 12267
rect 58052 12211 58208 12267
rect 58264 12211 86372 12267
rect 0 12161 86372 12211
rect 0 12105 26859 12161
rect 26915 12105 27071 12161
rect 27127 12105 86372 12161
rect 0 12049 86372 12105
rect 0 12046 57996 12049
rect 0 12036 24250 12046
rect 26772 11993 57996 12046
rect 58052 11993 58208 12049
rect 58264 12036 86372 12049
rect 58264 12035 84999 12036
rect 58264 11993 58351 12035
rect 26772 11844 58351 11993
rect 29478 11832 58351 11844
rect 29478 11776 57996 11832
rect 58052 11776 58208 11832
rect 58264 11776 58351 11832
rect 29478 11697 58351 11776
rect 0 11491 3011 11493
rect 24047 11491 27828 11493
rect 0 11406 27828 11491
rect 0 11350 27474 11406
rect 27530 11350 27686 11406
rect 27742 11350 27828 11406
rect 0 11189 27828 11350
rect 0 11133 27474 11189
rect 27530 11133 27686 11189
rect 27742 11133 27828 11189
rect 0 10971 27828 11133
rect 0 10915 27474 10971
rect 27530 10915 27686 10971
rect 27742 10915 27828 10971
rect 0 10753 27828 10915
rect 29478 10756 41516 11697
rect 0 10697 27474 10753
rect 27530 10697 27686 10753
rect 27742 10697 27828 10753
rect 0 10535 27828 10697
rect 0 10479 27474 10535
rect 27530 10479 27686 10535
rect 27742 10479 27828 10535
rect 0 10318 27828 10479
rect 0 10262 27474 10318
rect 27530 10262 27686 10318
rect 27742 10262 27828 10318
rect 0 10176 27828 10262
rect 2229 10175 24250 10176
rect 2249 10174 24250 10175
rect 23612 9942 29221 10030
rect 34741 9972 41516 10756
rect 42261 11491 57736 11527
rect 61825 11491 86372 11493
rect 42261 11406 86372 11491
rect 42261 11350 57381 11406
rect 57437 11350 57593 11406
rect 57649 11350 86372 11406
rect 42261 11189 86372 11350
rect 42261 11133 57381 11189
rect 57437 11133 57593 11189
rect 57649 11133 86372 11189
rect 42261 10971 86372 11133
rect 42261 10915 57381 10971
rect 57437 10915 57593 10971
rect 57649 10915 86372 10971
rect 42261 10753 86372 10915
rect 42261 10740 57381 10753
rect 57295 10697 57381 10740
rect 57437 10697 57593 10753
rect 57649 10697 86372 10753
rect 57295 10535 86372 10697
rect 57295 10479 57381 10535
rect 57437 10479 57593 10535
rect 57649 10479 86372 10535
rect 24047 9515 28729 9516
rect 0 9407 28729 9515
rect 0 9351 26859 9407
rect 26915 9351 27071 9407
rect 27127 9351 28729 9407
rect 0 9190 28729 9351
rect 29133 9302 29221 9942
rect 41857 9502 51430 10420
rect 57295 10318 86372 10479
rect 57295 10262 57381 10318
rect 57437 10262 57593 10318
rect 57649 10262 86372 10318
rect 51750 10097 54952 10185
rect 57295 10176 86372 10262
rect 61805 10175 84482 10176
rect 61825 10173 84482 10175
rect 51750 9971 51838 10097
rect 51750 9811 51766 9971
rect 51822 9811 51838 9971
rect 54864 10028 54952 10097
rect 54864 9940 62145 10028
rect 51750 9801 51838 9811
rect 58688 9681 61743 9777
rect 57909 9514 62278 9516
rect 83361 9514 86372 9515
rect 29133 9214 41656 9302
rect 0 9134 26859 9190
rect 26915 9134 27071 9190
rect 27127 9134 28729 9190
rect 0 8972 28729 9134
rect 0 8916 26859 8972
rect 26915 8916 27071 8972
rect 27127 8916 28729 8972
rect 0 8754 28729 8916
rect 41568 8972 41656 9214
rect 41857 9165 55482 9502
rect 41568 8956 50076 8972
rect 41568 8900 49906 8956
rect 50066 8900 50076 8956
rect 41568 8884 50076 8900
rect 50922 8888 55482 9165
rect 57909 9407 86372 9514
rect 57909 9351 57996 9407
rect 58052 9351 58208 9407
rect 58264 9351 86372 9407
rect 57909 9190 86372 9351
rect 57909 9134 57996 9190
rect 58052 9134 58208 9190
rect 58264 9134 86372 9190
rect 57909 8972 86372 9134
rect 57909 8916 57996 8972
rect 58052 8916 58208 8972
rect 58264 8916 86372 8972
rect 0 8698 26859 8754
rect 26915 8698 27071 8754
rect 27127 8698 28729 8754
rect 0 8536 28729 8698
rect 50922 8837 57736 8888
rect 50922 8781 57381 8837
rect 57437 8781 57593 8837
rect 57649 8781 57736 8837
rect 50922 8619 57736 8781
rect 0 8480 26859 8536
rect 26915 8480 27071 8536
rect 27127 8480 28729 8536
rect 0 8319 28729 8480
rect 0 8263 26859 8319
rect 26915 8263 27071 8319
rect 27127 8263 28729 8319
rect 0 8154 28729 8263
rect 0 8153 24250 8154
rect 0 8152 3011 8153
rect 28178 7652 28729 8154
rect 29513 7900 41397 8582
rect 0 7595 3011 7596
rect 23625 7595 27828 7596
rect 0 7535 27828 7595
rect 0 7479 27474 7535
rect 27530 7479 27686 7535
rect 27742 7479 27828 7535
rect 0 7317 27828 7479
rect 0 7261 27474 7317
rect 27530 7261 27686 7317
rect 27742 7261 27828 7317
rect 0 7099 27828 7261
rect 0 7043 27474 7099
rect 27530 7043 27686 7099
rect 27742 7043 27828 7099
rect 28178 7084 34622 7652
rect 0 6982 27828 7043
rect 0 6199 1014 6982
rect 2226 6981 24250 6982
rect 2249 6980 24250 6981
rect 23625 6836 29058 6875
rect 23625 6780 28273 6836
rect 28329 6780 28484 6836
rect 28540 6780 28696 6836
rect 28752 6780 28907 6836
rect 28963 6780 29058 6836
rect 23625 6618 29058 6780
rect 29537 6744 34622 7084
rect 34860 7392 41397 7900
rect 50922 8563 57381 8619
rect 57437 8563 57593 8619
rect 57649 8563 57736 8619
rect 50922 8402 57736 8563
rect 50922 8346 57381 8402
rect 57437 8346 57593 8402
rect 57649 8346 57736 8402
rect 50922 8184 57736 8346
rect 50922 8128 57381 8184
rect 57437 8128 57593 8184
rect 57649 8128 57736 8184
rect 57909 8754 86372 8916
rect 57909 8698 57996 8754
rect 58052 8698 58208 8754
rect 58264 8698 86372 8754
rect 57909 8536 86372 8698
rect 57909 8480 57996 8536
rect 58052 8480 58208 8536
rect 58264 8480 86372 8536
rect 57909 8319 86372 8480
rect 57909 8263 57996 8319
rect 58052 8263 58208 8319
rect 58264 8263 86372 8319
rect 57909 8154 86372 8263
rect 61802 8153 86372 8154
rect 61825 8152 86372 8153
rect 50922 7966 57736 8128
rect 50922 7910 57381 7966
rect 57437 7910 57593 7966
rect 57649 7910 57736 7966
rect 50922 7749 57736 7910
rect 50922 7693 57381 7749
rect 57437 7693 57593 7749
rect 57649 7693 57736 7749
rect 50922 7596 57736 7693
rect 50922 7595 62747 7596
rect 83361 7595 86372 7596
rect 50922 7531 86372 7595
rect 50922 7475 57381 7531
rect 57437 7475 57593 7531
rect 57649 7475 86372 7531
rect 50922 7392 86372 7475
rect 34860 7313 86372 7392
rect 34860 7257 57381 7313
rect 57437 7257 57593 7313
rect 57649 7257 86372 7313
rect 34860 7096 86372 7257
rect 34860 7040 57381 7096
rect 57437 7040 57593 7096
rect 57649 7040 86372 7096
rect 34860 6984 86372 7040
rect 23625 6562 28273 6618
rect 28329 6562 28484 6618
rect 28540 6562 28696 6618
rect 28752 6562 28907 6618
rect 28963 6562 29058 6618
rect 34860 6592 55482 6984
rect 57295 6982 86372 6984
rect 61802 6981 84787 6982
rect 61825 6980 84787 6981
rect 34860 6573 41397 6592
rect 23625 6400 29058 6562
rect 23625 6344 28273 6400
rect 28329 6344 28484 6400
rect 28540 6344 28696 6400
rect 28752 6344 28907 6400
rect 28963 6344 29058 6400
rect 23625 6306 29058 6344
rect 29458 6199 41397 6573
rect 0 6198 3011 6199
rect 23687 6198 41397 6199
rect 0 6177 41397 6198
rect 50922 6199 55482 6592
rect 56065 6836 62747 6875
rect 56065 6780 56160 6836
rect 56216 6780 56371 6836
rect 56427 6780 56583 6836
rect 56639 6780 56794 6836
rect 56850 6780 62747 6836
rect 56065 6618 62747 6780
rect 56065 6562 56160 6618
rect 56216 6562 56371 6618
rect 56427 6562 56583 6618
rect 56639 6562 56794 6618
rect 56850 6562 62747 6618
rect 56065 6400 62747 6562
rect 56065 6344 56160 6400
rect 56216 6344 56371 6400
rect 56427 6344 56583 6400
rect 56639 6344 56794 6400
rect 56850 6344 62747 6400
rect 56065 6306 62747 6344
rect 85358 6199 86372 6982
rect 50922 6198 62429 6199
rect 83361 6198 86372 6199
rect 0 6120 34622 6177
rect 0 6064 27474 6120
rect 27530 6064 27686 6120
rect 27742 6064 34622 6120
rect 0 5902 34622 6064
rect 0 5846 27474 5902
rect 27530 5846 27686 5902
rect 27742 5846 34622 5902
rect 0 5766 34622 5846
rect 29458 5665 34622 5766
rect 50922 6120 86372 6198
rect 50922 6064 57381 6120
rect 57437 6064 57593 6120
rect 57649 6064 86372 6120
rect 50922 5902 86372 6064
rect 50922 5846 57381 5902
rect 57437 5846 57593 5902
rect 57649 5846 86372 5902
rect 50922 5766 86372 5846
rect 23687 5629 27214 5630
rect 0 5539 27214 5629
rect 50922 5605 55482 5766
rect 57909 5629 62429 5630
rect 0 5483 26859 5539
rect 26915 5483 27071 5539
rect 27127 5483 27214 5539
rect 0 5321 27214 5483
rect 0 5265 26859 5321
rect 26915 5265 27071 5321
rect 27127 5265 27214 5321
rect 0 5175 27214 5265
rect 57909 5539 86372 5629
rect 57909 5483 57996 5539
rect 58052 5483 58208 5539
rect 58264 5483 86372 5539
rect 57909 5321 86372 5483
rect 57909 5265 57996 5321
rect 58052 5265 58208 5321
rect 58264 5265 86372 5321
rect 57909 5175 86372 5265
rect 0 5174 24250 5175
rect 61802 5174 86372 5175
rect 0 5173 3011 5174
rect 83361 5173 86372 5174
rect 0 4515 1712 5173
rect 57909 4619 62429 4621
rect 23909 4528 62429 4619
rect 23909 4515 26859 4528
rect 0 4472 26859 4515
rect 26915 4472 27071 4528
rect 27127 4472 57996 4528
rect 58052 4472 58208 4528
rect 58264 4515 62429 4528
rect 84660 4515 86372 5173
rect 58264 4472 86372 4515
rect 0 4310 86372 4472
rect 0 4254 26859 4310
rect 26915 4254 27071 4310
rect 27127 4254 57996 4310
rect 58052 4254 58208 4310
rect 58264 4254 86372 4310
rect 0 4166 86372 4254
rect 0 4164 59323 4166
rect 0 4060 24341 4164
rect 61788 4060 86372 4166
rect 27438 3875 27778 3876
rect 28764 3875 28894 3876
rect 41774 3875 41904 3876
rect 42299 3875 42429 3876
rect 46873 3875 47003 3876
rect 47321 3875 47451 3876
rect 47769 3875 47899 3876
rect 48217 3875 48347 3876
rect 57345 3875 61215 3876
rect 23909 3837 61215 3875
rect 23909 3781 27474 3837
rect 27530 3781 27686 3837
rect 27742 3781 28801 3837
rect 28857 3781 57381 3837
rect 57437 3781 57593 3837
rect 57649 3781 61215 3837
rect 23909 3772 61215 3781
rect 0 3619 86372 3772
rect 0 3563 27474 3619
rect 27530 3563 27686 3619
rect 27742 3563 28801 3619
rect 28857 3563 57381 3619
rect 57437 3563 57593 3619
rect 57649 3563 86372 3619
rect 0 3524 86372 3563
rect 0 3421 24341 3524
rect 0 3420 3011 3421
rect 60886 3420 86372 3524
rect 0 2854 1000 3420
rect 24169 3044 62588 3066
rect 24169 2988 43800 3044
rect 43960 2988 62588 3044
rect 24169 2978 62588 2988
rect 85358 2854 86372 3420
rect 0 2822 86372 2854
rect 0 2766 48671 2822
rect 48727 2766 48795 2822
rect 48851 2766 48919 2822
rect 48975 2766 86372 2822
rect 0 2698 86372 2766
rect 0 2642 48671 2698
rect 48727 2642 48795 2698
rect 48851 2642 48919 2698
rect 48975 2642 86372 2698
rect 0 2574 86372 2642
rect 0 2518 48671 2574
rect 48727 2518 48795 2574
rect 48851 2518 48919 2574
rect 48975 2518 86372 2574
rect 0 2502 86372 2518
rect 0 2199 86372 2232
rect 0 2143 49161 2199
rect 49217 2143 49285 2199
rect 49341 2143 49409 2199
rect 49465 2143 86372 2199
rect 0 2075 86372 2143
rect 0 2019 49161 2075
rect 49217 2019 49285 2075
rect 49341 2019 49409 2075
rect 49465 2019 86372 2075
rect 0 1951 86372 2019
rect 0 1895 49161 1951
rect 49217 1895 49285 1951
rect 49341 1895 49409 1951
rect 49465 1895 86372 1951
rect 0 1827 86372 1895
rect 0 1771 49161 1827
rect 49217 1771 49285 1827
rect 49341 1771 49409 1827
rect 49465 1771 86372 1827
rect 0 1703 86372 1771
rect 0 1647 49161 1703
rect 49217 1647 49285 1703
rect 49341 1647 49409 1703
rect 49465 1647 86372 1703
rect 0 1579 86372 1647
rect 0 1523 49161 1579
rect 49217 1523 49285 1579
rect 49341 1523 49409 1579
rect 49465 1523 86372 1579
rect 0 1455 86372 1523
rect 0 1399 49161 1455
rect 49217 1399 49285 1455
rect 49341 1399 49409 1455
rect 49465 1399 86372 1455
rect 0 1331 86372 1399
rect 0 1275 49161 1331
rect 49217 1275 49285 1331
rect 49341 1275 49409 1331
rect 49465 1275 86372 1331
rect 0 1232 86372 1275
rect 706 0 1706 1232
rect 2039 0 3039 1232
rect 3442 0 4442 1232
rect 4642 0 5642 932
rect 5842 0 6842 1232
rect 7042 0 8042 1232
rect 8242 0 9242 1232
rect 9442 0 10442 932
rect 10642 0 11642 1232
rect 12443 0 13443 1232
rect 14242 0 15242 1232
rect 15442 0 16442 932
rect 16642 0 17642 1232
rect 17842 0 18842 1232
rect 19042 0 20042 1232
rect 20242 0 21242 932
rect 21910 0 22910 1232
rect 23110 0 24110 1232
rect 24410 0 25410 1232
rect 25710 0 26710 1232
rect 27010 0 28010 1232
rect 28310 0 29310 1232
rect 29610 0 30610 1232
rect 31324 0 32324 932
rect 33022 0 34022 932
rect 34831 0 35831 932
rect 36031 0 37031 1232
rect 38028 0 39028 932
rect 39228 0 40228 1232
rect 41233 0 42233 932
rect 42433 0 43433 1232
rect 43633 0 44633 932
rect 44833 0 45833 1232
rect 46033 0 47033 932
rect 47233 0 48233 1232
rect 48566 0 49566 1232
rect 49876 0 50876 1232
rect 51233 0 52233 932
rect 52478 0 53478 932
rect 54458 0 55458 1232
rect 55758 0 56758 1232
rect 57058 0 58058 1232
rect 58358 0 59358 1232
rect 59658 0 60658 1232
rect 60958 0 61958 1232
rect 62295 0 63295 1232
rect 64218 0 65218 932
rect 65418 0 66418 1232
rect 66618 0 67618 1232
rect 67818 0 68818 1232
rect 69018 0 70018 932
rect 70218 0 71218 1232
rect 72017 0 73017 1232
rect 73818 0 74818 1232
rect 75018 0 76018 932
rect 76218 0 77218 1232
rect 77418 0 78418 1232
rect 78618 0 79618 1232
rect 79818 0 80818 932
rect 81018 0 82018 1232
rect 82419 0 83419 1232
rect 84666 0 85666 1232
use 128x8M8WM1_PWR_128x8m81  128x8M8WM1_PWR_128x8m81_0
timestamp 1698431365
transform 1 0 0 0 1 0
box 1912 6592 83548 35222
use control_512x8_128x8m81  control_512x8_128x8m81_0
timestamp 1698431365
transform 1 0 27533 0 1 4711
box -3624 -1833 31790 30125
use G_ring_128x8m81  G_ring_128x8m81_0
timestamp 1698431365
transform 1 0 282 0 1 0
box 0 0 85816 53502
use GF018_128x8M8WM1_lef_128x8m81  GF018_128x8M8WM1_lef_128x8m81_0
timestamp 1698431365
transform 1 0 0 0 1 0
box 0 0 86372 53776
use lcol4_128_128x8m81  lcol4_128_128x8m81_0
timestamp 1698431365
transform 1 0 2921 0 1 5019
box -1235 -3416 22810 46507
use M1_PSUB431059054877_128x8m81  M1_PSUB431059054877_128x8m81_0
timestamp 1698431365
transform 1 0 53710 0 1 2781
box 0 0 1 1
use M1_PSUB4310590548712_128x8m81  M1_PSUB4310590548712_128x8m81_0
timestamp 1698431365
transform 1 0 34404 0 1 2781
box 0 0 1 1
use M1_PSUB4310590548715_128x8m81  M1_PSUB4310590548715_128x8m81_0
timestamp 1698431365
transform 1 0 57403 0 1 1140
box 0 0 1 1
use M1_PSUB4310590548715_128x8m81  M1_PSUB4310590548715_128x8m81_1
timestamp 1698431365
transform 1 0 27521 0 1 1140
box 0 0 1 1
use M1_PSUB4310590548716_128x8m81  M1_PSUB4310590548716_128x8m81_0
timestamp 1698431365
transform 1 0 27869 0 1 34279
box 0 0 1 1
use M1_PSUB4310590548717_128x8m81  M1_PSUB4310590548717_128x8m81_0
timestamp 1698431365
transform 1 0 27869 0 1 36019
box 0 0 1 1
use M1_PSUB4310590548717_128x8m81  M1_PSUB4310590548717_128x8m81_1
timestamp 1698431365
transform 1 0 56655 0 1 36019
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_0
timestamp 1698431365
transform 1 0 28449 0 1 49627
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_1
timestamp 1698431365
transform 1 0 28449 0 1 47827
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_2
timestamp 1698431365
transform 1 0 28449 0 1 46027
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_3
timestamp 1698431365
transform 1 0 28449 0 1 44227
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_4
timestamp 1698431365
transform 1 0 28449 0 1 42427
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_5
timestamp 1698431365
transform 1 0 28449 0 1 37027
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_6
timestamp 1698431365
transform 1 0 28449 0 1 38827
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_7
timestamp 1698431365
transform 1 0 28449 0 1 40627
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_8
timestamp 1698431365
transform 1 0 28449 0 1 51427
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_9
timestamp 1698431365
transform 1 0 56674 0 1 47827
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_10
timestamp 1698431365
transform 1 0 56674 0 1 49627
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_11
timestamp 1698431365
transform 1 0 56674 0 1 51427
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_12
timestamp 1698431365
transform 1 0 56674 0 1 37027
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_13
timestamp 1698431365
transform 1 0 56674 0 1 38827
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_14
timestamp 1698431365
transform 1 0 56674 0 1 40627
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_15
timestamp 1698431365
transform 1 0 56674 0 1 42427
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_16
timestamp 1698431365
transform 1 0 56674 0 1 44227
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_17
timestamp 1698431365
transform 1 0 56674 0 1 46027
box 0 0 1 1
use M2_M1$$201260076_128x8m81  M2_M1$$201260076_128x8m81_0
timestamp 1698431365
transform -1 0 57515 0 1 19369
box 0 0 1 1
use M2_M1$$201260076_128x8m81  M2_M1$$201260076_128x8m81_1
timestamp 1698431365
transform -1 0 58130 0 1 19369
box 0 0 1 1
use M2_M1$$201260076_128x8m81  M2_M1$$201260076_128x8m81_2
timestamp 1698431365
transform 1 0 27608 0 1 19369
box 0 0 1 1
use M2_M1$$201260076_128x8m81  M2_M1$$201260076_128x8m81_3
timestamp 1698431365
transform 1 0 26993 0 1 19369
box 0 0 1 1
use M2_M1$$201261100_128x8m81  M2_M1$$201261100_128x8m81_0
timestamp 1698431365
transform -1 0 58130 0 1 4126
box 0 0 1 1
use M2_M1$$201261100_128x8m81  M2_M1$$201261100_128x8m81_1
timestamp 1698431365
transform -1 0 57515 0 1 4126
box 0 0 1 1
use M2_M1$$201261100_128x8m81  M2_M1$$201261100_128x8m81_2
timestamp 1698431365
transform 1 0 27608 0 1 4126
box 0 0 1 1
use M2_M1$$201261100_128x8m81  M2_M1$$201261100_128x8m81_3
timestamp 1698431365
transform 1 0 26993 0 1 4126
box 0 0 1 1
use M2_M1431059054870_128x8m81  M2_M1431059054870_128x8m81_0
timestamp 1698431365
transform 1 0 82808 0 1 1663
box 0 0 1 1
use M2_M1431059054870_128x8m81  M2_M1431059054870_128x8m81_1
timestamp 1698431365
transform 1 0 51732 0 1 5173
box 0 0 1 1
use M2_M1431059054870_128x8m81  M2_M1431059054870_128x8m81_2
timestamp 1698431365
transform 1 0 72743 0 1 1663
box 0 0 1 1
use M2_M1431059054870_128x8m81  M2_M1431059054870_128x8m81_3
timestamp 1698431365
transform 1 0 72293 0 1 1663
box 0 0 1 1
use M2_M1431059054870_128x8m81  M2_M1431059054870_128x8m81_4
timestamp 1698431365
transform 1 0 62228 0 1 1663
box 0 0 1 1
use M2_M1431059054870_128x8m81  M2_M1431059054870_128x8m81_5
timestamp 1698431365
transform 1 0 49986 0 1 6323
box 0 0 1 1
use M2_M1431059054870_128x8m81  M2_M1431059054870_128x8m81_6
timestamp 1698431365
transform 1 0 40700 0 1 4878
box 0 0 1 1
use M2_M1431059054870_128x8m81  M2_M1431059054870_128x8m81_7
timestamp 1698431365
transform 1 0 23517 0 1 1663
box 0 0 1 1
use M2_M1431059054870_128x8m81  M2_M1431059054870_128x8m81_8
timestamp 1698431365
transform 1 0 13167 0 1 1663
box 0 0 1 1
use M2_M1431059054870_128x8m81  M2_M1431059054870_128x8m81_9
timestamp 1698431365
transform 1 0 12717 0 1 1663
box 0 0 1 1
use M2_M1431059054870_128x8m81  M2_M1431059054870_128x8m81_10
timestamp 1698431365
transform 1 0 2652 0 1 1663
box 0 0 1 1
use M2_M1431059054873_128x8m81  M2_M1431059054873_128x8m81_0
timestamp 1698431365
transform 1 0 27590 0 1 34937
box 0 0 1 1
use M2_M1431059054875_128x8m81  M2_M1431059054875_128x8m81_0
timestamp 1698431365
transform 1 0 60601 0 1 35416
box 0 0 1 1
use M2_M14310590548711_128x8m81  M2_M14310590548711_128x8m81_0
timestamp 1698431365
transform 1 0 57507 0 1 34906
box 0 0 1 1
use M2_M14310590548713_128x8m81  M2_M14310590548713_128x8m81_0
timestamp 1698431365
transform 1 0 29818 0 1 785
box 0 0 1 1
use M2_M14310590548713_128x8m81  M2_M14310590548713_128x8m81_1
timestamp 1698431365
transform 1 0 29116 0 1 785
box 0 0 1 1
use M2_M14310590548719_128x8m81  M2_M14310590548719_128x8m81_0
timestamp 1698431365
transform 1 0 25674 0 1 51429
box 0 0 1 1
use M2_M14310590548719_128x8m81  M2_M14310590548719_128x8m81_1
timestamp 1698431365
transform 1 0 59152 0 1 51429
box 0 0 1 1
use M2_M14310590548721_128x8m81  M2_M14310590548721_128x8m81_0
timestamp 1698431365
transform 1 0 48818 0 1 764
box 0 0 1 1
use m2m3_128x8m81  m2m3_128x8m81_0
timestamp 1698431365
transform 1 0 58611 0 1 17122
box 0 0 3541 9202
use M3_M2$$201248812_128x8m81  M3_M2$$201248812_128x8m81_0
timestamp 1698431365
transform -1 0 58130 0 1 12783
box 0 0 1 1
use M3_M2$$201248812_128x8m81  M3_M2$$201248812_128x8m81_1
timestamp 1698431365
transform -1 0 57515 0 1 15671
box 0 0 1 1
use M3_M2$$201248812_128x8m81  M3_M2$$201248812_128x8m81_2
timestamp 1698431365
transform 1 0 27608 0 1 15463
box 0 0 1 1
use M3_M2$$201248812_128x8m81  M3_M2$$201248812_128x8m81_3
timestamp 1698431365
transform 1 0 26993 0 1 13112
box 0 0 1 1
use M3_M2$$201249836_128x8m81  M3_M2$$201249836_128x8m81_0
timestamp 1698431365
transform -1 0 57515 0 1 10834
box 0 0 1 1
use M3_M2$$201249836_128x8m81  M3_M2$$201249836_128x8m81_1
timestamp 1698431365
transform -1 0 58130 0 1 8835
box 0 0 1 1
use M3_M2$$201249836_128x8m81  M3_M2$$201249836_128x8m81_2
timestamp 1698431365
transform 1 0 27608 0 1 10834
box 0 0 1 1
use M3_M2$$201249836_128x8m81  M3_M2$$201249836_128x8m81_3
timestamp 1698431365
transform 1 0 26993 0 1 8835
box 0 0 1 1
use M3_M2$$201250860_128x8m81  M3_M2$$201250860_128x8m81_0
timestamp 1698431365
transform -1 0 56505 0 1 6590
box 0 0 1 1
use M3_M2$$201250860_128x8m81  M3_M2$$201250860_128x8m81_1
timestamp 1698431365
transform 1 0 28618 0 1 6590
box 0 0 1 1
use M3_M2$$201251884_128x8m81  M3_M2$$201251884_128x8m81_0
timestamp 1698431365
transform 1 0 37303 0 1 35853
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_0
timestamp 1698431365
transform 1 0 28829 0 1 3700
box 0 0 1 1
use M3_M2$$201253932_128x8m81  M3_M2$$201253932_128x8m81_0
timestamp 1698431365
transform 1 0 57515 0 1 8156
box 0 0 1 1
use M3_M2$$201254956_128x8m81  M3_M2$$201254956_128x8m81_0
timestamp 1698431365
transform 1 0 27608 0 1 13768
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_0
timestamp 1698431365
transform 1 0 28449 0 1 46027
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_1
timestamp 1698431365
transform 1 0 28449 0 1 44227
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_2
timestamp 1698431365
transform 1 0 28449 0 1 42427
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_3
timestamp 1698431365
transform 1 0 28449 0 1 40627
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_4
timestamp 1698431365
transform 1 0 28449 0 1 38827
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_5
timestamp 1698431365
transform 1 0 28449 0 1 37027
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_6
timestamp 1698431365
transform 1 0 28449 0 1 51427
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_7
timestamp 1698431365
transform 1 0 28449 0 1 49627
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_8
timestamp 1698431365
transform 1 0 28449 0 1 47827
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_9
timestamp 1698431365
transform 1 0 56674 0 1 38827
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_10
timestamp 1698431365
transform 1 0 56674 0 1 40627
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_11
timestamp 1698431365
transform 1 0 56674 0 1 42427
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_12
timestamp 1698431365
transform 1 0 56674 0 1 44227
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_13
timestamp 1698431365
transform 1 0 56674 0 1 46027
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_14
timestamp 1698431365
transform 1 0 56674 0 1 47827
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_15
timestamp 1698431365
transform 1 0 56674 0 1 49627
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_16
timestamp 1698431365
transform 1 0 56674 0 1 51427
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_17
timestamp 1698431365
transform 1 0 56674 0 1 37027
box 0 0 1 1
use M3_M2$$201412652_128x8m81  M3_M2$$201412652_128x8m81_0
timestamp 1698431365
transform 1 0 27608 0 1 32786
box 0 0 1 1
use M3_M2$$201412652_128x8m81  M3_M2$$201412652_128x8m81_1
timestamp 1698431365
transform 1 0 27608 0 1 30897
box 0 0 1 1
use M3_M2$$201412652_128x8m81  M3_M2$$201412652_128x8m81_2
timestamp 1698431365
transform -1 0 57515 0 1 30897
box 0 0 1 1
use M3_M2$$201412652_128x8m81  M3_M2$$201412652_128x8m81_3
timestamp 1698431365
transform -1 0 57515 0 1 32786
box 0 0 1 1
use M3_M2$$201413676_128x8m81  M3_M2$$201413676_128x8m81_0
timestamp 1698431365
transform 1 0 27608 0 1 7289
box 0 0 1 1
use M3_M2$$201413676_128x8m81  M3_M2$$201413676_128x8m81_1
timestamp 1698431365
transform 1 0 26993 0 1 31842
box 0 0 1 1
use M3_M2$$201413676_128x8m81  M3_M2$$201413676_128x8m81_2
timestamp 1698431365
transform -1 0 58130 0 1 31842
box 0 0 1 1
use M3_M2$$201414700_128x8m81  M3_M2$$201414700_128x8m81_0
timestamp 1698431365
transform 1 0 26993 0 1 33221
box 0 0 1 1
use M3_M2$$201414700_128x8m81  M3_M2$$201414700_128x8m81_1
timestamp 1698431365
transform -1 0 58130 0 1 33221
box 0 0 1 1
use M3_M2$$201415724_128x8m81  M3_M2$$201415724_128x8m81_0
timestamp 1698431365
transform 1 0 26993 0 1 28743
box 0 0 1 1
use M3_M2$$201415724_128x8m81  M3_M2$$201415724_128x8m81_1
timestamp 1698431365
transform -1 0 58130 0 1 28743
box 0 0 1 1
use M3_M2$$201416748_128x8m81  M3_M2$$201416748_128x8m81_0
timestamp 1698431365
transform -1 0 58130 0 1 4391
box 0 0 1 1
use M3_M2$$201416748_128x8m81  M3_M2$$201416748_128x8m81_1
timestamp 1698431365
transform -1 0 57515 0 1 26662
box 0 0 1 1
use M3_M2$$201416748_128x8m81  M3_M2$$201416748_128x8m81_2
timestamp 1698431365
transform -1 0 57515 0 1 3700
box 0 0 1 1
use M3_M2$$201416748_128x8m81  M3_M2$$201416748_128x8m81_3
timestamp 1698431365
transform -1 0 58130 0 1 5402
box 0 0 1 1
use M3_M2$$201416748_128x8m81  M3_M2$$201416748_128x8m81_4
timestamp 1698431365
transform -1 0 57515 0 1 5983
box 0 0 1 1
use M3_M2$$201416748_128x8m81  M3_M2$$201416748_128x8m81_5
timestamp 1698431365
transform 1 0 27608 0 1 3700
box 0 0 1 1
use M3_M2$$201416748_128x8m81  M3_M2$$201416748_128x8m81_6
timestamp 1698431365
transform 1 0 26993 0 1 4391
box 0 0 1 1
use M3_M2$$201416748_128x8m81  M3_M2$$201416748_128x8m81_7
timestamp 1698431365
transform 1 0 27608 0 1 5983
box 0 0 1 1
use M3_M2$$201416748_128x8m81  M3_M2$$201416748_128x8m81_8
timestamp 1698431365
transform 1 0 26993 0 1 5402
box 0 0 1 1
use M3_M2$$201416748_128x8m81  M3_M2$$201416748_128x8m81_9
timestamp 1698431365
transform 1 0 27608 0 1 26662
box 0 0 1 1
use M3_M2$$201416748_128x8m81  M3_M2$$201416748_128x8m81_10
timestamp 1698431365
transform 1 0 27608 0 1 24891
box 0 0 1 1
use M3_M2431059054871_128x8m81  M3_M2431059054871_128x8m81_0
timestamp 1698431365
transform 0 -1 49986 1 0 8928
box 0 0 1 1
use M3_M2431059054871_128x8m81  M3_M2431059054871_128x8m81_1
timestamp 1698431365
transform 1 0 51794 0 1 9891
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_0
timestamp 1698431365
transform 1 0 58128 0 1 20490
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_1
timestamp 1698431365
transform 1 0 58128 0 1 20146
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_2
timestamp 1698431365
transform 1 0 26187 0 1 19267
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_3
timestamp 1698431365
transform 1 0 26530 0 1 26206
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_4
timestamp 1698431365
transform 1 0 26545 0 1 19612
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_5
timestamp 1698431365
transform 1 0 27004 0 1 20490
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_6
timestamp 1698431365
transform 1 0 27004 0 1 20146
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_7
timestamp 1698431365
transform 1 0 24137 0 1 23593
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_8
timestamp 1698431365
transform 1 0 24149 0 1 17237
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_9
timestamp 1698431365
transform 1 0 24496 0 1 23915
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_10
timestamp 1698431365
transform 1 0 24509 0 1 17576
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_11
timestamp 1698431365
transform 1 0 24824 0 1 24236
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_12
timestamp 1698431365
transform 1 0 24837 0 1 17897
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_13
timestamp 1698431365
transform 1 0 25161 0 1 24557
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_14
timestamp 1698431365
transform 1 0 25174 0 1 18270
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_15
timestamp 1698431365
transform 1 0 25501 0 1 25248
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_16
timestamp 1698431365
transform 1 0 25514 0 1 18604
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_17
timestamp 1698431365
transform 1 0 25836 0 1 25567
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_18
timestamp 1698431365
transform 1 0 25851 0 1 18947
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_19
timestamp 1698431365
transform 1 0 26172 0 1 25887
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_20
timestamp 1698431365
transform 1 0 41955 0 1 50533
box 0 0 1 1
use M3_M2431059054874_128x8m81  M3_M2431059054874_128x8m81_0
timestamp 1698431365
transform 1 0 43880 0 1 3016
box 0 0 1 1
use M3_M2431059054876_128x8m81  M3_M2431059054876_128x8m81_0
timestamp 1698431365
transform 1 0 25674 0 1 51420
box 0 0 1 1
use M3_M2431059054876_128x8m81  M3_M2431059054876_128x8m81_1
timestamp 1698431365
transform 1 0 25674 0 1 31096
box 0 0 1 1
use M3_M2431059054876_128x8m81  M3_M2431059054876_128x8m81_2
timestamp 1698431365
transform 1 0 25674 0 1 30641
box 0 0 1 1
use M3_M2431059054876_128x8m81  M3_M2431059054876_128x8m81_3
timestamp 1698431365
transform 1 0 59149 0 1 31146
box 0 0 1 1
use M3_M2431059054876_128x8m81  M3_M2431059054876_128x8m81_4
timestamp 1698431365
transform 1 0 59149 0 1 30701
box 0 0 1 1
use M3_M2431059054876_128x8m81  M3_M2431059054876_128x8m81_5
timestamp 1698431365
transform 1 0 59152 0 1 51420
box 0 0 1 1
use M3_M2431059054878_128x8m81  M3_M2431059054878_128x8m81_0
timestamp 1698431365
transform 1 0 25660 0 1 34937
box 0 0 1 1
use M3_M2431059054878_128x8m81  M3_M2431059054878_128x8m81_1
timestamp 1698431365
transform 1 0 59149 0 1 34906
box 0 0 1 1
use M3_M2431059054879_128x8m81  M3_M2431059054879_128x8m81_0
timestamp 1698431365
transform 1 0 49313 0 1 1737
box 0 0 1 1
use M3_M24310590548710_128x8m81  M3_M24310590548710_128x8m81_0
timestamp 1698431365
transform 1 0 48823 0 1 2670
box 0 0 1 1
use M3_M24310590548714_128x8m81  M3_M24310590548714_128x8m81_0
timestamp 1698431365
transform 1 0 59135 0 1 27428
box 0 0 1 1
use M3_M24310590548714_128x8m81  M3_M24310590548714_128x8m81_1
timestamp 1698431365
transform 1 0 25680 0 1 27367
box 0 0 1 1
use M3_M24310590548718_128x8m81  M3_M24310590548718_128x8m81_0
timestamp 1698431365
transform 1 0 27590 0 1 34937
box 0 0 1 1
use M3_M24310590548720_128x8m81  M3_M24310590548720_128x8m81_0
timestamp 1698431365
transform 1 0 57495 0 1 22479
box 0 0 1 1
use M3_M24310590548720_128x8m81  M3_M24310590548720_128x8m81_1
timestamp 1698431365
transform 1 0 58126 0 1 23631
box 0 0 1 1
use M3_M24310590548720_128x8m81  M3_M24310590548720_128x8m81_2
timestamp 1698431365
transform 1 0 26990 0 1 23631
box 0 0 1 1
use M3_M24310590548720_128x8m81  M3_M24310590548720_128x8m81_3
timestamp 1698431365
transform 1 0 27607 0 1 22492
box 0 0 1 1
use power_a_128x8m81  power_a_128x8m81_0
timestamp 1698431365
transform -1 0 80818 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_1
timestamp 1698431365
transform 1 0 51233 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_2
timestamp 1698431365
transform 1 0 64218 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_3
timestamp 1698431365
transform 1 0 52478 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_4
timestamp 1698431365
transform 1 0 75018 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_5
timestamp 1698431365
transform 1 0 46033 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_6
timestamp 1698431365
transform 1 0 43633 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_7
timestamp 1698431365
transform -1 0 70018 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_8
timestamp 1698431365
transform -1 0 10442 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_9
timestamp 1698431365
transform -1 0 32324 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_10
timestamp 1698431365
transform -1 0 21242 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_11
timestamp 1698431365
transform -1 0 34022 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_12
timestamp 1698431365
transform 1 0 41233 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_13
timestamp 1698431365
transform 1 0 34831 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_14
timestamp 1698431365
transform 1 0 15442 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_15
timestamp 1698431365
transform 1 0 38028 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_16
timestamp 1698431365
transform 1 0 4642 0 1 282
box 0 -282 1000 1000
use power_route_01_a_128x8m81  power_route_01_a_128x8m81_0
timestamp 1698431365
transform 1 0 15448 0 1 51346
box -511 630 1714 2430
use power_route_01_a_128x8m81  power_route_01_a_128x8m81_1
timestamp 1698431365
transform 1 0 10048 0 1 51346
box -511 630 1714 2430
use power_route_01_a_128x8m81  power_route_01_a_128x8m81_2
timestamp 1698431365
transform 1 0 4648 0 1 51346
box -511 630 1714 2430
use power_route_01_a_128x8m81  power_route_01_a_128x8m81_3
timestamp 1698431365
transform 1 0 64224 0 1 51346
box -511 630 1714 2430
use power_route_01_a_128x8m81  power_route_01_a_128x8m81_4
timestamp 1698431365
transform 1 0 69624 0 1 51346
box -511 630 1714 2430
use power_route_01_a_128x8m81  power_route_01_a_128x8m81_5
timestamp 1698431365
transform 1 0 75024 0 1 51346
box -511 630 1714 2430
use power_route_01_a_128x8m81  power_route_01_a_128x8m81_6
timestamp 1698431365
transform 1 0 46824 0 1 51346
box -511 630 1714 2430
use power_route_01_b_128x8m81  power_route_01_b_128x8m81_0
timestamp 1698431365
transform -1 0 21142 0 1 51346
box -511 630 489 2430
use power_route_01_b_128x8m81  power_route_01_b_128x8m81_1
timestamp 1698431365
transform -1 0 41719 0 1 51346
box -511 630 489 2430
use power_route_01_b_128x8m81  power_route_01_b_128x8m81_2
timestamp 1698431365
transform -1 0 80718 0 1 51346
box -511 630 489 2430
use power_route_01_b_128x8m81  power_route_01_b_128x8m81_3
timestamp 1698431365
transform -1 0 85155 0 1 51346
box -511 630 489 2430
use power_route_01_b_128x8m81  power_route_01_b_128x8m81_4
timestamp 1698431365
transform -1 0 45558 0 1 51346
box -511 630 489 2430
use power_route_01_c_128x8m81  power_route_01_c_128x8m81_0
timestamp 1698431365
transform -1 0 34095 0 1 51346
box 714 1822 1714 2430
use power_route_01_c_128x8m81  power_route_01_c_128x8m81_1
timestamp 1698431365
transform -1 0 38662 0 1 51346
box 714 1822 1714 2430
use power_route_01_c_128x8m81  power_route_01_c_128x8m81_2
timestamp 1698431365
transform -1 0 30987 0 1 51346
box 714 1822 1714 2430
use power_route_01_c_128x8m81  power_route_01_c_128x8m81_3
timestamp 1698431365
transform -1 0 29591 0 1 51346
box 714 1822 1714 2430
use power_route_01_c_128x8m81  power_route_01_c_128x8m81_4
timestamp 1698431365
transform -1 0 44144 0 1 51346
box 714 1822 1714 2430
use power_route_128_128x8m81  power_route_128_128x8m81_0
timestamp 1698431365
transform 1 0 -1921 0 1 -2063
box 1921 2345 88293 55839
use rcol4_128_128x8m81  rcol4_128_128x8m81_0
timestamp 1698431365
transform 1 0 60511 0 1 5019
box -1090 -3398 24602 46517
use xdec16_128_128x8m81  xdec16_128_128x8m81_0
timestamp 1698431365
transform 1 0 28677 0 1 36127
box -3364 -228 31133 15548
<< labels >>
flabel metal3 s 2626 53168 3626 53776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 50176 1706 50876 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 48376 1706 49076 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 4642 0 5642 932 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 5362 53168 6362 53776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 46576 1706 47276 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 44776 1706 45476 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 8026 53168 9026 53776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 42976 1706 43676 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 41176 1706 41876 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 39376 1706 40076 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 37576 1706 38276 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 9442 0 10442 932 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 35776 1706 36476 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 8152 3011 9515 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 10762 53168 11762 53776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 8153 24250 9515 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 13426 53168 14426 53776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 15442 0 16442 932 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 16162 53168 17162 53776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 28178 7084 28729 9516 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 24047 8154 28729 9516 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 29537 6744 34622 7652 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 18826 53168 19826 53776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 20242 0 21242 932 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 28178 7084 34622 7652 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 22258 53168 23258 53776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 25158 53168 26158 53776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 1401 51976 2401 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 4137 51976 5137 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 34536 27828 35326 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 6801 51976 7801 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 6921 26434 8163 28416 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 17721 26434 18963 28416 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 26435 26070 28416 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 9537 51976 10537 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 26435 27828 26890 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 12201 51976 13201 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 14937 51976 15937 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 10176 3011 11493 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 2249 10174 24250 11491 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 17601 51976 18601 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 20653 51976 21653 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 2229 10175 24250 11491 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 24047 10176 27828 11493 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 27877 53168 28877 53776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 29273 53168 30273 53776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 23483 51976 24483 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 31324 0 32324 932 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 26572 51976 27572 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 32381 53168 33381 53776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 30710 51976 31710 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 35415 51976 36415 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 33022 0 34022 932 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 38585 51976 39585 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 34024 53168 35024 53776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 34831 0 35831 932 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 41230 51976 42230 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 45069 51976 46069 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 36948 53168 37948 53776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 38028 0 39028 932 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 39882 53168 40882 53776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 46313 51976 47313 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 41233 0 42233 932 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 42430 53168 43430 53776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 48901 51976 49901 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 52569 51976 53569 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 54262 51976 55262 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 43633 0 44633 932 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 43713 53168 44713 53776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 57547 51976 58547 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 60977 51976 61977 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 46033 0 47033 932 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 47538 53168 48538 53776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 63713 51976 64713 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 50465 53168 51465 53776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 66377 51976 67377 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 51233 0 52233 932 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 69113 51976 70113 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 71777 51976 72777 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 52478 0 53478 932 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 55990 53168 56990 53776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 74513 51976 75513 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 77177 51976 78177 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 80229 51976 81229 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 83059 51976 84059 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 84666 51976 85666 53776 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 51976 86372 52976 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 84666 50176 86372 50876 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 58791 53168 59791 53776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 62202 53168 63202 53776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 64218 0 65218 932 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 84666 48376 86372 49076 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 64938 53168 65938 53776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 67602 53168 68602 53776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 84666 46576 86372 47276 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 69018 0 70018 932 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 70338 53168 71338 53776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 84666 44776 86372 45476 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 84666 42976 86372 43676 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 73002 53168 74002 53776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 75018 0 76018 932 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 75738 53168 76738 53776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 84666 41176 86372 41876 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 78402 53168 79402 53776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 84666 39376 86372 40076 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 79818 0 80818 932 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 84666 37576 86372 38276 0 FreeSans 1600 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 81834 53168 82834 53776 0 FreeSans 1600 180 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 84666 35776 86372 36476 0 FreeSans 1600 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 29430 1706 34125 0 FreeSans 1600 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 2095 32315 2188 34126 0 FreeSans 1600 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 51076 1014 51776 0 FreeSans 1600 180 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 32315 3011 34125 0 FreeSans 1600 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 32316 25085 34125 0 FreeSans 1600 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 51226 27779 51626 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 32318 27214 34124 0 FreeSans 1600 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 26772 31486 58351 32199 0 FreeSans 1600 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 30402 51326 54622 51528 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 26772 27382 58351 30105 0 FreeSans 1600 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 57908 31486 58351 34124 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 61853 32315 72383 34125 0 FreeSans 1600 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 57908 32315 86372 34124 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 51327 86372 51528 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 29430 86372 29714 0 FreeSans 1600 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 84666 29430 86372 34125 0 FreeSans 1600 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 58791 51258 59517 51591 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 72653 32315 86372 34125 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 58791 51276 86372 51576 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 22938 1706 23938 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 85358 51076 86372 51776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 22938 27214 23380 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 49276 1014 49976 0 FreeSans 1600 180 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 26770 23370 58348 24278 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 57908 22937 83763 23380 0 FreeSans 1600 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 57908 22938 86372 23380 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 84666 22938 86372 23938 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 18016 24250 20739 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 49476 27272 49776 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 29513 19969 55645 21625 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 30403 49526 54622 49728 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 49526 86372 49726 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 59421 49476 86372 49776 0 FreeSans 1600 180 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 85358 49276 86372 49976 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 29521 19969 55645 21707 0 FreeSans 1600 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 44432 19969 55645 21708 0 FreeSans 1600 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 61825 18015 83763 20739 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 61807 18016 86372 20739 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 19969 86372 20739 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 47476 1014 48176 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 47676 27272 47976 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 12036 1706 14178 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 23821 12046 34761 12847 0 FreeSans 1600 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 13461 27214 14178 0 FreeSans 1600 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 12036 24250 12846 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 24047 12046 27214 14179 0 FreeSans 1600 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 30403 47726 54622 47928 0 FreeSans 1600 180 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 24047 12046 34761 12934 0 FreeSans 1600 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 34741 9972 41516 12574 0 FreeSans 1600 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 29478 10756 41516 12574 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 29478 11697 58351 12574 0 FreeSans 1600 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 47726 86372 47926 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 59421 47676 86372 47976 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 85358 47476 86372 48176 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 45676 1014 46376 0 FreeSans 1600 180 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 26772 11844 58351 12574 0 FreeSans 1600 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 50228 12035 58421 13866 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 59826 12035 60026 14017 0 FreeSans 1600 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 50228 13461 86372 13866 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 61807 13461 72429 14178 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 61773 13461 86372 14177 0 FreeSans 1600 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 83169 12035 84221 12847 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 45876 27272 46176 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 83169 13461 84221 14179 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 50228 12036 86372 12846 0 FreeSans 1600 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 26772 12035 84999 12574 0 FreeSans 1600 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 84666 12036 86372 14178 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 72607 13461 86372 14178 0 FreeSans 1600 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 61802 8153 86372 9514 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 57909 8154 62278 9516 0 FreeSans 1600 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 61825 8152 86372 9514 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 30403 45926 54622 46128 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 83361 8152 86372 9515 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 45926 86372 46126 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 59421 45876 86372 46176 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 4060 1712 5629 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 85358 45676 86372 46376 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 5173 3011 5629 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 43876 1014 44576 0 FreeSans 1600 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 5174 24250 5629 0 FreeSans 1600 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 4060 24341 4515 0 FreeSans 1600 180 0 0 VDD
port 27 nsew power bidirectional
rlabel metal2 s 27936 0 28160 200 4 CLK
port 9 nsew signal input
rlabel metal2 s 1864 0 2088 200 4 D[0]
port 17 nsew signal input
rlabel metal2 s 30859 0 31083 200 4 A[2]
port 5 nsew signal input
rlabel metal2 s 32552 0 32776 200 4 A[1]
port 6 nsew signal input
rlabel metal2 s 34243 0 34467 200 4 A[0]
port 7 nsew signal input
rlabel metal2 s 14127 0 14351 200 4 Q[2]
port 24 nsew signal output
rlabel metal2 s 22279 0 22503 200 4 Q[3]
port 23 nsew signal output
rlabel metal2 s 50342 0 50566 200 4 CEN
port 8 nsew signal input
rlabel metal2 s 54417 0 54641 200 4 A[5]
port 2 nsew signal input
rlabel metal2 s 53772 0 53996 200 4 A[6]
port 1 nsew signal input
rlabel metal2 s 55164 0 55388 200 4 A[4]
port 3 nsew signal input
rlabel metal2 s 23404 0 23628 200 4 WEN[3]
port 33 nsew signal input
rlabel metal2 s 83372 0 83596 200 4 D[7]
port 10 nsew signal input
rlabel metal2 s 81855 0 82079 200 4 Q[7]
port 19 nsew signal output
rlabel metal2 s 23795 0 24019 200 4 D[3]
port 14 nsew signal input
rlabel metal2 s 12206 0 12430 200 4 D[1]
port 16 nsew signal input
rlabel metal2 s 13454 0 13678 200 4 D[2]
port 15 nsew signal input
rlabel metal2 s 56265 0 56489 200 4 A[3]
port 4 nsew signal input
rlabel metal2 s 11533 0 11757 200 4 Q[1]
port 25 nsew signal output
rlabel metal2 s 73703 0 73927 200 4 Q[6]
port 20 nsew signal output
rlabel metal2 s 71782 0 72006 200 4 D[5]
port 12 nsew signal input
rlabel metal2 s 62958 0 63182 200 4 Q[4]
port 22 nsew signal output
rlabel metal2 s 72180 0 72404 200 4 WEN[5]
port 31 nsew signal input
rlabel metal2 s 13054 0 13278 200 4 WEN[2]
port 34 nsew signal input
rlabel metal2 s 12604 0 12828 200 4 WEN[1]
port 35 nsew signal input
rlabel metal2 s 62115 0 62339 200 4 WEN[4]
port 32 nsew signal input
rlabel metal2 s 82695 0 82919 200 4 WEN[7]
port 29 nsew signal input
rlabel metal2 s 72630 0 72854 200 4 WEN[6]
port 30 nsew signal input
rlabel metal2 s 61447 0 61671 200 4 D[4]
port 13 nsew signal input
rlabel metal2 s 73030 0 73254 200 4 D[6]
port 11 nsew signal input
rlabel metal2 s 71109 0 71333 200 4 Q[5]
port 21 nsew signal output
rlabel metal2 s 3380 0 3604 200 4 Q[0]
port 26 nsew signal output
rlabel metal2 s 40588 0 40812 200 4 GWEN
port 18 nsew signal input
rlabel metal2 s 2539 0 2763 200 4 WEN[0]
port 36 nsew signal input
rlabel metal3 s 23687 5175 27214 5630 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 23909 4166 62429 4619 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 4164 59323 4515 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 57909 4166 62429 4621 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 57909 5175 62429 5630 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 61788 4060 86372 4515 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 83361 5173 86372 5629 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 61802 5174 86372 5629 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 84660 4060 86372 5629 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 706 0 1706 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 2039 0 3039 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 3442 0 4442 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 5842 0 6842 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 7042 0 8042 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 8242 0 9242 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 10642 0 11642 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 12443 0 13443 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 14242 0 15242 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 16642 0 17642 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 17842 0 18842 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 19042 0 20042 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 21910 0 22910 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 23110 0 24110 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 24410 0 25410 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 25710 0 26710 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 27010 0 28010 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 28310 0 29310 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 29610 0 30610 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 36031 0 37031 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 39228 0 40228 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 42433 0 43433 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 44833 0 45833 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 47233 0 48233 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 48566 0 49566 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 49876 0 50876 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 54458 0 55458 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 55758 0 56758 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 57058 0 58058 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 58358 0 59358 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 59658 0 60658 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 60958 0 61958 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 62295 0 63295 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 65418 0 66418 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 66618 0 67618 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 67818 0 68818 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 70218 0 71218 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 72017 0 73017 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 73818 0 74818 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 76218 0 77218 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 77418 0 78418 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 78618 0 79618 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 81018 0 82018 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 82419 0 83419 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 84666 0 85666 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 1232 86372 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 44076 27272 44376 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 30403 44126 54622 44328 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 44126 86372 44326 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 59421 44076 86372 44376 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 85358 43876 86372 44576 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 42076 1014 42776 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 42276 27272 42576 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 30403 42326 54622 42528 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 42326 86372 42526 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 59421 42276 86372 42576 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 85358 42076 86372 42776 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 40276 1014 40976 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 40476 27272 40776 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 30403 40526 54622 40728 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 40526 86372 40726 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 59421 40476 86372 40776 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 85358 40276 86372 40976 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 38476 1014 39176 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 38676 27272 38976 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 30403 38726 54622 38928 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 38726 86372 38926 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 59421 38676 86372 38976 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 85358 38476 86372 39176 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 36676 1014 37376 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 36876 27272 37176 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 30403 36926 54622 37128 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 36926 86372 37126 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 59421 36876 86372 37176 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 85358 36676 86372 37376 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 57369 34536 86372 35326 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 57295 26435 86372 26890 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 66497 26434 67739 28416 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 77297 26434 78539 28416 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 58785 26435 86372 28416 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 21282 1014 22282 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 24036 21826 27826 22282 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 21827 27826 22282 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 27387 21826 27826 23199 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 56078 21826 57677 23199 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 27387 22291 57677 23199 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 56078 21826 83763 22282 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 85358 21282 86372 22282 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 56078 21827 86372 22282 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 14328 23678 17730 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 14328 24250 16597 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 24111 14329 27828 16598 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 29478 13243 45977 15015 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 27387 13245 45977 15015 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 14491 47683 15015 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 41493 13078 49775 13760 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 14936 51760 15015 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 14966 55645 15015 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 46982 14968 86372 16784 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 57295 14327 83763 16784 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 61807 14328 86372 17730 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 42261 10740 57736 11527 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 57295 10176 86372 11491 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 61825 10173 84482 11493 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 61805 10175 84482 11491 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 61825 10176 86372 11493 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 5766 1014 7596 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 5766 3011 6199 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 6982 3011 7596 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 2249 6980 24250 7595 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 2226 6981 24250 7595 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 23625 6982 27828 7596 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 23687 6177 41397 6199 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 29458 5665 34622 6573 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 5766 34622 6198 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 29458 6177 41397 6573 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 34860 6177 41397 8582 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 29513 7900 41397 8582 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 34860 6592 55482 7392 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 41857 9165 51430 10420 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 50922 5605 55482 9502 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 50922 6984 57736 8888 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 57295 6982 86372 7595 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 50922 5766 62429 6199 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 50922 6984 62747 7596 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 50922 5766 86372 6198 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 61825 6980 84787 7595 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 61802 6981 84787 7595 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 83361 5766 86372 6199 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 85358 5766 86372 7596 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 83361 6982 86372 7596 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 2502 1000 3772 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 3420 3011 3772 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 3421 24341 3772 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 27438 3524 27778 3876 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 28764 3524 28894 3876 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 41774 3524 41904 3876 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 42299 3524 42429 3876 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 46873 3524 47003 3876 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 47321 3524 47451 3876 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 47769 3524 47899 3876 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 48217 3524 48347 3876 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 23909 3524 61215 3875 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 57345 3524 61215 3876 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 2502 86372 2854 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 60886 3420 86372 3772 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 85358 2502 86372 3772 1 VSS
port 28 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 86372 53776
string GDS_END 2348274
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 2298700
string LEFclass BLOCK
string LEFsymmetry X Y R90
string path 307.290 11.160 307.290 0.000 
<< end >>
