magic
tech gf180mcuA
magscale 1 10
timestamp 1698431365
<< nwell >>
rect 600 14610 3070 14628
rect 255 -210 3070 14610
rect 4721 -178 7236 14578
rect 600 -228 3070 -210
rect 8461 -228 9061 14628
rect 14259 14577 18306 14627
rect 23622 14609 24064 14610
rect 14259 -177 19597 14577
rect 14259 -227 18306 -177
rect 21249 -209 24064 14609
rect 23622 -210 24064 -209
<< nmos >>
rect 13292 14217 13922 14337
rect 3268 13748 4268 13868
rect 13292 14004 13922 14124
rect 13292 13780 13922 13900
rect 20051 13748 21051 13868
rect 3268 13132 4268 13252
rect 13292 13100 13922 13220
rect 20051 13132 21051 13252
rect 13292 12876 13922 12996
rect 13292 12663 13922 12783
rect 13292 12417 13922 12537
rect 3268 11948 4268 12068
rect 13292 12204 13922 12324
rect 13292 11980 13922 12100
rect 20051 11948 21051 12068
rect 3268 11332 4268 11452
rect 13292 11300 13922 11420
rect 20051 11332 21051 11452
rect 13292 11076 13922 11196
rect 13292 10863 13922 10983
rect 13292 10617 13922 10737
rect 3268 10148 4268 10268
rect 13292 10404 13922 10524
rect 13292 10180 13922 10300
rect 20051 10148 21051 10268
rect 3268 9532 4268 9652
rect 13292 9500 13922 9620
rect 20051 9532 21051 9652
rect 13292 9276 13922 9396
rect 13292 9063 13922 9183
rect 13292 8817 13922 8937
rect 3268 8348 4268 8468
rect 13292 8604 13922 8724
rect 13292 8380 13922 8500
rect 20051 8348 21051 8468
rect 3268 7732 4268 7852
rect 13292 7700 13922 7820
rect 20051 7732 21051 7852
rect 13292 7476 13922 7596
rect 13292 7263 13922 7383
rect 13292 7017 13922 7137
rect 3268 6548 4268 6668
rect 13292 6804 13922 6924
rect 13292 6580 13922 6700
rect 20051 6548 21051 6668
rect 3268 5932 4268 6052
rect 13292 5900 13922 6020
rect 20051 5932 21051 6052
rect 13292 5676 13922 5796
rect 13292 5463 13922 5583
rect 13292 5217 13922 5337
rect 3268 4748 4268 4868
rect 13292 5004 13922 5124
rect 13292 4780 13922 4900
rect 20051 4748 21051 4868
rect 3268 4132 4268 4252
rect 13292 4100 13922 4220
rect 20051 4132 21051 4252
rect 13292 3876 13922 3996
rect 13292 3663 13922 3783
rect 13292 3417 13922 3537
rect 3268 2948 4268 3068
rect 13292 3204 13922 3324
rect 13292 2980 13922 3100
rect 20051 2948 21051 3068
rect 3268 2332 4268 2452
rect 13292 2300 13922 2420
rect 20051 2332 21051 2452
rect 13292 2076 13922 2196
rect 13292 1863 13922 1983
rect 13292 1617 13922 1737
rect 3268 1148 4268 1268
rect 13292 1404 13922 1524
rect 13292 1180 13922 1300
rect 20051 1148 21051 1268
rect 3268 532 4268 652
rect 13292 500 13922 620
rect 20051 532 21051 652
rect 13292 276 13922 396
rect 13292 63 13922 183
<< mvnmos >>
rect 3268 14228 4268 14348
rect 9324 14228 9764 14348
rect 3268 14004 4268 14124
rect 20051 14228 21051 14348
rect 7493 13917 8153 14037
rect 7493 13693 8153 13813
rect 9195 13693 9327 13813
rect 20051 14004 21051 14124
rect 3268 12876 4268 12996
rect 7493 13187 8153 13307
rect 7493 12963 8153 13083
rect 9195 13187 9327 13307
rect 20051 12876 21051 12996
rect 3268 12652 4268 12772
rect 3268 12428 4268 12548
rect 9324 12652 9764 12772
rect 9324 12428 9764 12548
rect 20051 12652 21051 12772
rect 3268 12204 4268 12324
rect 20051 12428 21051 12548
rect 7493 12117 8153 12237
rect 7493 11893 8153 12013
rect 9195 11893 9327 12013
rect 20051 12204 21051 12324
rect 3268 11076 4268 11196
rect 7493 11387 8153 11507
rect 7493 11163 8153 11283
rect 9195 11387 9327 11507
rect 20051 11076 21051 11196
rect 3268 10852 4268 10972
rect 3268 10628 4268 10748
rect 9324 10852 9764 10972
rect 9324 10628 9764 10748
rect 20051 10852 21051 10972
rect 3268 10404 4268 10524
rect 20051 10628 21051 10748
rect 7493 10317 8153 10437
rect 7493 10093 8153 10213
rect 9195 10093 9327 10213
rect 20051 10404 21051 10524
rect 3268 9276 4268 9396
rect 7493 9587 8153 9707
rect 7493 9363 8153 9483
rect 9195 9587 9327 9707
rect 20051 9276 21051 9396
rect 3268 9052 4268 9172
rect 3268 8828 4268 8948
rect 9324 9052 9764 9172
rect 9324 8828 9764 8948
rect 20051 9052 21051 9172
rect 3268 8604 4268 8724
rect 20051 8828 21051 8948
rect 7493 8517 8153 8637
rect 7493 8293 8153 8413
rect 9195 8293 9327 8413
rect 20051 8604 21051 8724
rect 3268 7476 4268 7596
rect 7493 7787 8153 7907
rect 7493 7563 8153 7683
rect 9195 7787 9327 7907
rect 20051 7476 21051 7596
rect 3268 7252 4268 7372
rect 3268 7028 4268 7148
rect 9324 7252 9764 7372
rect 9324 7028 9764 7148
rect 20051 7252 21051 7372
rect 3268 6804 4268 6924
rect 20051 7028 21051 7148
rect 7493 6717 8153 6837
rect 7493 6493 8153 6613
rect 9195 6493 9327 6613
rect 20051 6804 21051 6924
rect 3268 5676 4268 5796
rect 7493 5987 8153 6107
rect 7493 5763 8153 5883
rect 9195 5987 9327 6107
rect 20051 5676 21051 5796
rect 3268 5452 4268 5572
rect 3268 5228 4268 5348
rect 9324 5452 9764 5572
rect 9324 5228 9764 5348
rect 20051 5452 21051 5572
rect 3268 5004 4268 5124
rect 20051 5228 21051 5348
rect 7493 4917 8153 5037
rect 7493 4693 8153 4813
rect 9195 4693 9327 4813
rect 20051 5004 21051 5124
rect 3268 3876 4268 3996
rect 7493 4187 8153 4307
rect 7493 3963 8153 4083
rect 9195 4187 9327 4307
rect 20051 3876 21051 3996
rect 3268 3652 4268 3772
rect 3268 3428 4268 3548
rect 9324 3652 9764 3772
rect 9324 3428 9764 3548
rect 20051 3652 21051 3772
rect 3268 3204 4268 3324
rect 20051 3428 21051 3548
rect 7493 3117 8153 3237
rect 7493 2893 8153 3013
rect 9195 2893 9327 3013
rect 20051 3204 21051 3324
rect 3268 2076 4268 2196
rect 7493 2387 8153 2507
rect 7493 2163 8153 2283
rect 9195 2387 9327 2507
rect 20051 2076 21051 2196
rect 3268 1852 4268 1972
rect 3268 1628 4268 1748
rect 9324 1852 9764 1972
rect 9324 1628 9764 1748
rect 20051 1852 21051 1972
rect 3268 1404 4268 1524
rect 20051 1628 21051 1748
rect 7493 1317 8153 1437
rect 7493 1093 8153 1213
rect 9195 1093 9327 1213
rect 20051 1404 21051 1524
rect 3268 276 4268 396
rect 7493 587 8153 707
rect 7493 363 8153 483
rect 9195 587 9327 707
rect 20051 276 21051 396
rect 3268 52 4268 172
rect 9324 52 9764 172
rect 20051 52 21051 172
<< mvpmos >>
rect 933 14228 2933 14348
rect 933 14004 2933 14124
rect 933 13780 2933 13900
rect 14396 14228 14920 14348
rect 21386 14228 23386 14348
rect 4857 13917 5957 14037
rect 4857 13693 5957 13813
rect 6438 13917 7098 14037
rect 14396 14004 14920 14124
rect 6438 13693 7098 13813
rect 8605 13693 8923 13813
rect 14396 13780 14920 13900
rect 18362 13917 19462 14037
rect 18362 13693 19462 13813
rect 21386 14004 23386 14124
rect 21386 13780 23386 13900
rect 933 13100 2933 13220
rect 933 12876 2933 12996
rect 933 12652 2933 12772
rect 4857 13187 5957 13307
rect 4857 12963 5957 13083
rect 6438 13187 7098 13307
rect 6438 12963 7098 13083
rect 8605 13187 8923 13307
rect 14396 13100 14920 13220
rect 18362 13187 19462 13307
rect 14396 12876 14920 12996
rect 18362 12963 19462 13083
rect 933 12428 2933 12548
rect 933 12204 2933 12324
rect 933 11980 2933 12100
rect 14396 12652 14920 12772
rect 21386 13100 23386 13220
rect 21386 12876 23386 12996
rect 21386 12652 23386 12772
rect 14396 12428 14920 12548
rect 21386 12428 23386 12548
rect 4857 12117 5957 12237
rect 4857 11893 5957 12013
rect 6438 12117 7098 12237
rect 14396 12204 14920 12324
rect 6438 11893 7098 12013
rect 8605 11893 8923 12013
rect 14396 11980 14920 12100
rect 18362 12117 19462 12237
rect 18362 11893 19462 12013
rect 21386 12204 23386 12324
rect 21386 11980 23386 12100
rect 933 11300 2933 11420
rect 933 11076 2933 11196
rect 933 10852 2933 10972
rect 4857 11387 5957 11507
rect 4857 11163 5957 11283
rect 6438 11387 7098 11507
rect 6438 11163 7098 11283
rect 8605 11387 8923 11507
rect 14396 11300 14920 11420
rect 18362 11387 19462 11507
rect 14396 11076 14920 11196
rect 18362 11163 19462 11283
rect 933 10628 2933 10748
rect 933 10404 2933 10524
rect 933 10180 2933 10300
rect 14396 10852 14920 10972
rect 21386 11300 23386 11420
rect 21386 11076 23386 11196
rect 21386 10852 23386 10972
rect 14396 10628 14920 10748
rect 21386 10628 23386 10748
rect 4857 10317 5957 10437
rect 4857 10093 5957 10213
rect 6438 10317 7098 10437
rect 14396 10404 14920 10524
rect 6438 10093 7098 10213
rect 8605 10093 8923 10213
rect 14396 10180 14920 10300
rect 18362 10317 19462 10437
rect 18362 10093 19462 10213
rect 21386 10404 23386 10524
rect 21386 10180 23386 10300
rect 933 9500 2933 9620
rect 933 9276 2933 9396
rect 933 9052 2933 9172
rect 4857 9587 5957 9707
rect 4857 9363 5957 9483
rect 6438 9587 7098 9707
rect 6438 9363 7098 9483
rect 8605 9587 8923 9707
rect 14396 9500 14920 9620
rect 18362 9587 19462 9707
rect 14396 9276 14920 9396
rect 18362 9363 19462 9483
rect 933 8828 2933 8948
rect 933 8604 2933 8724
rect 933 8380 2933 8500
rect 14396 9052 14920 9172
rect 21386 9500 23386 9620
rect 21386 9276 23386 9396
rect 21386 9052 23386 9172
rect 14396 8828 14920 8948
rect 21386 8828 23386 8948
rect 4857 8517 5957 8637
rect 4857 8293 5957 8413
rect 6438 8517 7098 8637
rect 14396 8604 14920 8724
rect 6438 8293 7098 8413
rect 8605 8293 8923 8413
rect 14396 8380 14920 8500
rect 18362 8517 19462 8637
rect 18362 8293 19462 8413
rect 21386 8604 23386 8724
rect 21386 8380 23386 8500
rect 933 7700 2933 7820
rect 933 7476 2933 7596
rect 933 7252 2933 7372
rect 4857 7787 5957 7907
rect 4857 7563 5957 7683
rect 6438 7787 7098 7907
rect 6438 7563 7098 7683
rect 8605 7787 8923 7907
rect 14396 7700 14920 7820
rect 18362 7787 19462 7907
rect 14396 7476 14920 7596
rect 18362 7563 19462 7683
rect 933 7028 2933 7148
rect 933 6804 2933 6924
rect 933 6580 2933 6700
rect 14396 7252 14920 7372
rect 21386 7700 23386 7820
rect 21386 7476 23386 7596
rect 21386 7252 23386 7372
rect 14396 7028 14920 7148
rect 21386 7028 23386 7148
rect 4857 6717 5957 6837
rect 4857 6493 5957 6613
rect 6438 6717 7098 6837
rect 14396 6804 14920 6924
rect 6438 6493 7098 6613
rect 8605 6493 8923 6613
rect 14396 6580 14920 6700
rect 18362 6717 19462 6837
rect 18362 6493 19462 6613
rect 21386 6804 23386 6924
rect 21386 6580 23386 6700
rect 933 5900 2933 6020
rect 933 5676 2933 5796
rect 933 5452 2933 5572
rect 4857 5987 5957 6107
rect 4857 5763 5957 5883
rect 6438 5987 7098 6107
rect 6438 5763 7098 5883
rect 8605 5987 8923 6107
rect 14396 5900 14920 6020
rect 18362 5987 19462 6107
rect 14396 5676 14920 5796
rect 18362 5763 19462 5883
rect 933 5228 2933 5348
rect 933 5004 2933 5124
rect 933 4780 2933 4900
rect 14396 5452 14920 5572
rect 21386 5900 23386 6020
rect 21386 5676 23386 5796
rect 21386 5452 23386 5572
rect 14396 5228 14920 5348
rect 21386 5228 23386 5348
rect 4857 4917 5957 5037
rect 4857 4693 5957 4813
rect 6438 4917 7098 5037
rect 14396 5004 14920 5124
rect 6438 4693 7098 4813
rect 8605 4693 8923 4813
rect 14396 4780 14920 4900
rect 18362 4917 19462 5037
rect 18362 4693 19462 4813
rect 21386 5004 23386 5124
rect 21386 4780 23386 4900
rect 933 4100 2933 4220
rect 933 3876 2933 3996
rect 933 3652 2933 3772
rect 4857 4187 5957 4307
rect 4857 3963 5957 4083
rect 6438 4187 7098 4307
rect 6438 3963 7098 4083
rect 8605 4187 8923 4307
rect 14396 4100 14920 4220
rect 18362 4187 19462 4307
rect 14396 3876 14920 3996
rect 18362 3963 19462 4083
rect 933 3428 2933 3548
rect 933 3204 2933 3324
rect 933 2980 2933 3100
rect 14396 3652 14920 3772
rect 21386 4100 23386 4220
rect 21386 3876 23386 3996
rect 21386 3652 23386 3772
rect 14396 3428 14920 3548
rect 21386 3428 23386 3548
rect 4857 3117 5957 3237
rect 4857 2893 5957 3013
rect 6438 3117 7098 3237
rect 14396 3204 14920 3324
rect 6438 2893 7098 3013
rect 8605 2893 8923 3013
rect 14396 2980 14920 3100
rect 18362 3117 19462 3237
rect 18362 2893 19462 3013
rect 21386 3204 23386 3324
rect 21386 2980 23386 3100
rect 933 2300 2933 2420
rect 933 2076 2933 2196
rect 933 1852 2933 1972
rect 4857 2387 5957 2507
rect 4857 2163 5957 2283
rect 6438 2387 7098 2507
rect 6438 2163 7098 2283
rect 8605 2387 8923 2507
rect 14396 2300 14920 2420
rect 18362 2387 19462 2507
rect 14396 2076 14920 2196
rect 18362 2163 19462 2283
rect 933 1628 2933 1748
rect 933 1404 2933 1524
rect 933 1180 2933 1300
rect 14396 1852 14920 1972
rect 21386 2300 23386 2420
rect 21386 2076 23386 2196
rect 21386 1852 23386 1972
rect 14396 1628 14920 1748
rect 21386 1628 23386 1748
rect 4857 1317 5957 1437
rect 4857 1093 5957 1213
rect 6438 1317 7098 1437
rect 14396 1404 14920 1524
rect 6438 1093 7098 1213
rect 8605 1093 8923 1213
rect 14396 1180 14920 1300
rect 18362 1317 19462 1437
rect 18362 1093 19462 1213
rect 21386 1404 23386 1524
rect 21386 1180 23386 1300
rect 933 500 2933 620
rect 933 276 2933 396
rect 933 52 2933 172
rect 4857 587 5957 707
rect 4857 363 5957 483
rect 6438 587 7098 707
rect 6438 363 7098 483
rect 8605 587 8923 707
rect 14396 500 14920 620
rect 18362 587 19462 707
rect 14396 276 14920 396
rect 18362 363 19462 483
rect 14396 52 14920 172
rect 21386 500 23386 620
rect 21386 276 23386 396
rect 21386 52 23386 172
<< ndiff >>
rect 13292 14423 13922 14469
rect 13292 14377 13336 14423
rect 13382 14377 13503 14423
rect 13549 14377 13668 14423
rect 13714 14377 13833 14423
rect 13879 14377 13922 14423
rect 13292 14337 13922 14377
rect 13292 14124 13922 14217
rect 3268 13716 4268 13748
rect 3268 13670 3413 13716
rect 3459 13670 3599 13716
rect 3645 13670 3786 13716
rect 3832 13670 3973 13716
rect 4019 13670 4159 13716
rect 4205 13670 4268 13716
rect 13292 13900 13922 14004
rect 13292 13730 13922 13780
rect 3268 13624 4268 13670
rect 13292 13684 13336 13730
rect 13382 13684 13503 13730
rect 13549 13684 13668 13730
rect 13714 13684 13833 13730
rect 13879 13684 13922 13730
rect 20051 13716 21051 13748
rect 13292 13637 13922 13684
rect 20051 13670 20113 13716
rect 20159 13670 20300 13716
rect 20346 13670 20487 13716
rect 20533 13670 20673 13716
rect 20719 13670 20860 13716
rect 20906 13670 21051 13716
rect 20051 13624 21051 13670
rect 3268 13330 4268 13376
rect 3268 13284 3413 13330
rect 3459 13284 3599 13330
rect 3645 13284 3786 13330
rect 3832 13284 3973 13330
rect 4019 13284 4159 13330
rect 4205 13284 4268 13330
rect 13292 13316 13922 13363
rect 3268 13252 4268 13284
rect 13292 13270 13336 13316
rect 13382 13270 13503 13316
rect 13549 13270 13668 13316
rect 13714 13270 13833 13316
rect 13879 13270 13922 13316
rect 13292 13220 13922 13270
rect 20051 13330 21051 13376
rect 20051 13284 20113 13330
rect 20159 13284 20300 13330
rect 20346 13284 20487 13330
rect 20533 13284 20673 13330
rect 20719 13284 20860 13330
rect 20906 13284 21051 13330
rect 20051 13252 21051 13284
rect 13292 12996 13922 13100
rect 13292 12783 13922 12876
rect 13292 12623 13922 12663
rect 13292 12577 13336 12623
rect 13382 12577 13503 12623
rect 13549 12577 13668 12623
rect 13714 12577 13833 12623
rect 13879 12577 13922 12623
rect 13292 12537 13922 12577
rect 13292 12324 13922 12417
rect 3268 11916 4268 11948
rect 3268 11870 3413 11916
rect 3459 11870 3599 11916
rect 3645 11870 3786 11916
rect 3832 11870 3973 11916
rect 4019 11870 4159 11916
rect 4205 11870 4268 11916
rect 13292 12100 13922 12204
rect 13292 11930 13922 11980
rect 3268 11824 4268 11870
rect 13292 11884 13336 11930
rect 13382 11884 13503 11930
rect 13549 11884 13668 11930
rect 13714 11884 13833 11930
rect 13879 11884 13922 11930
rect 20051 11916 21051 11948
rect 13292 11837 13922 11884
rect 20051 11870 20113 11916
rect 20159 11870 20300 11916
rect 20346 11870 20487 11916
rect 20533 11870 20673 11916
rect 20719 11870 20860 11916
rect 20906 11870 21051 11916
rect 20051 11824 21051 11870
rect 3268 11530 4268 11576
rect 3268 11484 3413 11530
rect 3459 11484 3599 11530
rect 3645 11484 3786 11530
rect 3832 11484 3973 11530
rect 4019 11484 4159 11530
rect 4205 11484 4268 11530
rect 13292 11516 13922 11563
rect 3268 11452 4268 11484
rect 13292 11470 13336 11516
rect 13382 11470 13503 11516
rect 13549 11470 13668 11516
rect 13714 11470 13833 11516
rect 13879 11470 13922 11516
rect 13292 11420 13922 11470
rect 20051 11530 21051 11576
rect 20051 11484 20113 11530
rect 20159 11484 20300 11530
rect 20346 11484 20487 11530
rect 20533 11484 20673 11530
rect 20719 11484 20860 11530
rect 20906 11484 21051 11530
rect 20051 11452 21051 11484
rect 13292 11196 13922 11300
rect 13292 10983 13922 11076
rect 13292 10823 13922 10863
rect 13292 10777 13336 10823
rect 13382 10777 13503 10823
rect 13549 10777 13668 10823
rect 13714 10777 13833 10823
rect 13879 10777 13922 10823
rect 13292 10737 13922 10777
rect 13292 10524 13922 10617
rect 3268 10116 4268 10148
rect 3268 10070 3413 10116
rect 3459 10070 3599 10116
rect 3645 10070 3786 10116
rect 3832 10070 3973 10116
rect 4019 10070 4159 10116
rect 4205 10070 4268 10116
rect 13292 10300 13922 10404
rect 13292 10130 13922 10180
rect 3268 10024 4268 10070
rect 13292 10084 13336 10130
rect 13382 10084 13503 10130
rect 13549 10084 13668 10130
rect 13714 10084 13833 10130
rect 13879 10084 13922 10130
rect 20051 10116 21051 10148
rect 13292 10037 13922 10084
rect 20051 10070 20113 10116
rect 20159 10070 20300 10116
rect 20346 10070 20487 10116
rect 20533 10070 20673 10116
rect 20719 10070 20860 10116
rect 20906 10070 21051 10116
rect 20051 10024 21051 10070
rect 3268 9730 4268 9776
rect 3268 9684 3413 9730
rect 3459 9684 3599 9730
rect 3645 9684 3786 9730
rect 3832 9684 3973 9730
rect 4019 9684 4159 9730
rect 4205 9684 4268 9730
rect 13292 9716 13922 9763
rect 3268 9652 4268 9684
rect 13292 9670 13336 9716
rect 13382 9670 13503 9716
rect 13549 9670 13668 9716
rect 13714 9670 13833 9716
rect 13879 9670 13922 9716
rect 13292 9620 13922 9670
rect 20051 9730 21051 9776
rect 20051 9684 20113 9730
rect 20159 9684 20300 9730
rect 20346 9684 20487 9730
rect 20533 9684 20673 9730
rect 20719 9684 20860 9730
rect 20906 9684 21051 9730
rect 20051 9652 21051 9684
rect 13292 9396 13922 9500
rect 13292 9183 13922 9276
rect 13292 9023 13922 9063
rect 13292 8977 13336 9023
rect 13382 8977 13503 9023
rect 13549 8977 13668 9023
rect 13714 8977 13833 9023
rect 13879 8977 13922 9023
rect 13292 8937 13922 8977
rect 13292 8724 13922 8817
rect 3268 8316 4268 8348
rect 3268 8270 3413 8316
rect 3459 8270 3599 8316
rect 3645 8270 3786 8316
rect 3832 8270 3973 8316
rect 4019 8270 4159 8316
rect 4205 8270 4268 8316
rect 13292 8500 13922 8604
rect 13292 8330 13922 8380
rect 3268 8224 4268 8270
rect 13292 8284 13336 8330
rect 13382 8284 13503 8330
rect 13549 8284 13668 8330
rect 13714 8284 13833 8330
rect 13879 8284 13922 8330
rect 20051 8316 21051 8348
rect 13292 8237 13922 8284
rect 20051 8270 20113 8316
rect 20159 8270 20300 8316
rect 20346 8270 20487 8316
rect 20533 8270 20673 8316
rect 20719 8270 20860 8316
rect 20906 8270 21051 8316
rect 20051 8224 21051 8270
rect 3268 7930 4268 7976
rect 3268 7884 3413 7930
rect 3459 7884 3599 7930
rect 3645 7884 3786 7930
rect 3832 7884 3973 7930
rect 4019 7884 4159 7930
rect 4205 7884 4268 7930
rect 13292 7916 13922 7963
rect 3268 7852 4268 7884
rect 13292 7870 13336 7916
rect 13382 7870 13503 7916
rect 13549 7870 13668 7916
rect 13714 7870 13833 7916
rect 13879 7870 13922 7916
rect 13292 7820 13922 7870
rect 20051 7930 21051 7976
rect 20051 7884 20113 7930
rect 20159 7884 20300 7930
rect 20346 7884 20487 7930
rect 20533 7884 20673 7930
rect 20719 7884 20860 7930
rect 20906 7884 21051 7930
rect 20051 7852 21051 7884
rect 13292 7596 13922 7700
rect 13292 7383 13922 7476
rect 13292 7223 13922 7263
rect 13292 7177 13336 7223
rect 13382 7177 13503 7223
rect 13549 7177 13668 7223
rect 13714 7177 13833 7223
rect 13879 7177 13922 7223
rect 13292 7137 13922 7177
rect 13292 6924 13922 7017
rect 3268 6516 4268 6548
rect 3268 6470 3413 6516
rect 3459 6470 3599 6516
rect 3645 6470 3786 6516
rect 3832 6470 3973 6516
rect 4019 6470 4159 6516
rect 4205 6470 4268 6516
rect 13292 6700 13922 6804
rect 13292 6530 13922 6580
rect 3268 6424 4268 6470
rect 13292 6484 13336 6530
rect 13382 6484 13503 6530
rect 13549 6484 13668 6530
rect 13714 6484 13833 6530
rect 13879 6484 13922 6530
rect 20051 6516 21051 6548
rect 13292 6437 13922 6484
rect 20051 6470 20113 6516
rect 20159 6470 20300 6516
rect 20346 6470 20487 6516
rect 20533 6470 20673 6516
rect 20719 6470 20860 6516
rect 20906 6470 21051 6516
rect 20051 6424 21051 6470
rect 3268 6130 4268 6176
rect 3268 6084 3413 6130
rect 3459 6084 3599 6130
rect 3645 6084 3786 6130
rect 3832 6084 3973 6130
rect 4019 6084 4159 6130
rect 4205 6084 4268 6130
rect 13292 6116 13922 6163
rect 3268 6052 4268 6084
rect 13292 6070 13336 6116
rect 13382 6070 13503 6116
rect 13549 6070 13668 6116
rect 13714 6070 13833 6116
rect 13879 6070 13922 6116
rect 13292 6020 13922 6070
rect 20051 6130 21051 6176
rect 20051 6084 20113 6130
rect 20159 6084 20300 6130
rect 20346 6084 20487 6130
rect 20533 6084 20673 6130
rect 20719 6084 20860 6130
rect 20906 6084 21051 6130
rect 20051 6052 21051 6084
rect 13292 5796 13922 5900
rect 13292 5583 13922 5676
rect 13292 5423 13922 5463
rect 13292 5377 13336 5423
rect 13382 5377 13503 5423
rect 13549 5377 13668 5423
rect 13714 5377 13833 5423
rect 13879 5377 13922 5423
rect 13292 5337 13922 5377
rect 13292 5124 13922 5217
rect 3268 4716 4268 4748
rect 3268 4670 3413 4716
rect 3459 4670 3599 4716
rect 3645 4670 3786 4716
rect 3832 4670 3973 4716
rect 4019 4670 4159 4716
rect 4205 4670 4268 4716
rect 13292 4900 13922 5004
rect 13292 4730 13922 4780
rect 3268 4624 4268 4670
rect 13292 4684 13336 4730
rect 13382 4684 13503 4730
rect 13549 4684 13668 4730
rect 13714 4684 13833 4730
rect 13879 4684 13922 4730
rect 20051 4716 21051 4748
rect 13292 4637 13922 4684
rect 20051 4670 20113 4716
rect 20159 4670 20300 4716
rect 20346 4670 20487 4716
rect 20533 4670 20673 4716
rect 20719 4670 20860 4716
rect 20906 4670 21051 4716
rect 20051 4624 21051 4670
rect 3268 4330 4268 4376
rect 3268 4284 3413 4330
rect 3459 4284 3599 4330
rect 3645 4284 3786 4330
rect 3832 4284 3973 4330
rect 4019 4284 4159 4330
rect 4205 4284 4268 4330
rect 13292 4316 13922 4363
rect 3268 4252 4268 4284
rect 13292 4270 13336 4316
rect 13382 4270 13503 4316
rect 13549 4270 13668 4316
rect 13714 4270 13833 4316
rect 13879 4270 13922 4316
rect 13292 4220 13922 4270
rect 20051 4330 21051 4376
rect 20051 4284 20113 4330
rect 20159 4284 20300 4330
rect 20346 4284 20487 4330
rect 20533 4284 20673 4330
rect 20719 4284 20860 4330
rect 20906 4284 21051 4330
rect 20051 4252 21051 4284
rect 13292 3996 13922 4100
rect 13292 3783 13922 3876
rect 13292 3623 13922 3663
rect 13292 3577 13336 3623
rect 13382 3577 13503 3623
rect 13549 3577 13668 3623
rect 13714 3577 13833 3623
rect 13879 3577 13922 3623
rect 13292 3537 13922 3577
rect 13292 3324 13922 3417
rect 3268 2916 4268 2948
rect 3268 2870 3413 2916
rect 3459 2870 3599 2916
rect 3645 2870 3786 2916
rect 3832 2870 3973 2916
rect 4019 2870 4159 2916
rect 4205 2870 4268 2916
rect 13292 3100 13922 3204
rect 13292 2930 13922 2980
rect 3268 2824 4268 2870
rect 13292 2884 13336 2930
rect 13382 2884 13503 2930
rect 13549 2884 13668 2930
rect 13714 2884 13833 2930
rect 13879 2884 13922 2930
rect 20051 2916 21051 2948
rect 13292 2837 13922 2884
rect 20051 2870 20113 2916
rect 20159 2870 20300 2916
rect 20346 2870 20487 2916
rect 20533 2870 20673 2916
rect 20719 2870 20860 2916
rect 20906 2870 21051 2916
rect 20051 2824 21051 2870
rect 3268 2530 4268 2576
rect 3268 2484 3413 2530
rect 3459 2484 3599 2530
rect 3645 2484 3786 2530
rect 3832 2484 3973 2530
rect 4019 2484 4159 2530
rect 4205 2484 4268 2530
rect 13292 2516 13922 2563
rect 3268 2452 4268 2484
rect 13292 2470 13336 2516
rect 13382 2470 13503 2516
rect 13549 2470 13668 2516
rect 13714 2470 13833 2516
rect 13879 2470 13922 2516
rect 13292 2420 13922 2470
rect 20051 2530 21051 2576
rect 20051 2484 20113 2530
rect 20159 2484 20300 2530
rect 20346 2484 20487 2530
rect 20533 2484 20673 2530
rect 20719 2484 20860 2530
rect 20906 2484 21051 2530
rect 20051 2452 21051 2484
rect 13292 2196 13922 2300
rect 13292 1983 13922 2076
rect 13292 1823 13922 1863
rect 13292 1777 13336 1823
rect 13382 1777 13503 1823
rect 13549 1777 13668 1823
rect 13714 1777 13833 1823
rect 13879 1777 13922 1823
rect 13292 1737 13922 1777
rect 13292 1524 13922 1617
rect 3268 1116 4268 1148
rect 3268 1070 3413 1116
rect 3459 1070 3599 1116
rect 3645 1070 3786 1116
rect 3832 1070 3973 1116
rect 4019 1070 4159 1116
rect 4205 1070 4268 1116
rect 13292 1300 13922 1404
rect 13292 1130 13922 1180
rect 3268 1024 4268 1070
rect 13292 1084 13336 1130
rect 13382 1084 13503 1130
rect 13549 1084 13668 1130
rect 13714 1084 13833 1130
rect 13879 1084 13922 1130
rect 20051 1116 21051 1148
rect 13292 1037 13922 1084
rect 20051 1070 20113 1116
rect 20159 1070 20300 1116
rect 20346 1070 20487 1116
rect 20533 1070 20673 1116
rect 20719 1070 20860 1116
rect 20906 1070 21051 1116
rect 20051 1024 21051 1070
rect 3268 730 4268 776
rect 3268 684 3413 730
rect 3459 684 3599 730
rect 3645 684 3786 730
rect 3832 684 3973 730
rect 4019 684 4159 730
rect 4205 684 4268 730
rect 13292 716 13922 763
rect 3268 652 4268 684
rect 13292 670 13336 716
rect 13382 670 13503 716
rect 13549 670 13668 716
rect 13714 670 13833 716
rect 13879 670 13922 716
rect 13292 620 13922 670
rect 20051 730 21051 776
rect 20051 684 20113 730
rect 20159 684 20300 730
rect 20346 684 20487 730
rect 20533 684 20673 730
rect 20719 684 20860 730
rect 20906 684 21051 730
rect 20051 652 21051 684
rect 13292 396 13922 500
rect 13292 183 13922 276
rect 13292 23 13922 63
rect 13292 -23 13336 23
rect 13382 -23 13503 23
rect 13549 -23 13668 23
rect 13714 -23 13833 23
rect 13879 -23 13922 23
rect 13292 -69 13922 -23
<< mvndiff >>
rect 3268 14423 4268 14436
rect 3268 14377 3281 14423
rect 3327 14377 3384 14423
rect 3430 14377 3487 14423
rect 3533 14377 3590 14423
rect 3636 14377 3693 14423
rect 3739 14377 3796 14423
rect 3842 14377 3899 14423
rect 3945 14377 4002 14423
rect 4048 14377 4105 14423
rect 4151 14377 4209 14423
rect 4255 14377 4268 14423
rect 3268 14348 4268 14377
rect 9324 14423 9764 14436
rect 9324 14377 9337 14423
rect 9383 14377 9459 14423
rect 9505 14377 9582 14423
rect 9628 14377 9705 14423
rect 9751 14377 9764 14423
rect 9324 14348 9764 14377
rect 3268 14199 4268 14228
rect 3268 14153 3281 14199
rect 3327 14153 3384 14199
rect 3430 14153 3487 14199
rect 3533 14153 3590 14199
rect 3636 14153 3693 14199
rect 3739 14153 3796 14199
rect 3842 14153 3899 14199
rect 3945 14153 4002 14199
rect 4048 14153 4105 14199
rect 4151 14153 4209 14199
rect 4255 14153 4268 14199
rect 3268 14124 4268 14153
rect 9324 14199 9764 14228
rect 9324 14153 9337 14199
rect 9383 14153 9459 14199
rect 9505 14153 9582 14199
rect 9628 14153 9705 14199
rect 9751 14153 9764 14199
rect 9324 14140 9764 14153
rect 20051 14423 21051 14436
rect 20051 14377 20064 14423
rect 20110 14377 20168 14423
rect 20214 14377 20271 14423
rect 20317 14377 20374 14423
rect 20420 14377 20477 14423
rect 20523 14377 20580 14423
rect 20626 14377 20683 14423
rect 20729 14377 20786 14423
rect 20832 14377 20889 14423
rect 20935 14377 20992 14423
rect 21038 14377 21051 14423
rect 20051 14348 21051 14377
rect 7493 14112 8153 14125
rect 20051 14199 21051 14228
rect 20051 14153 20064 14199
rect 20110 14153 20168 14199
rect 20214 14153 20271 14199
rect 20317 14153 20374 14199
rect 20420 14153 20477 14199
rect 20523 14153 20580 14199
rect 20626 14153 20683 14199
rect 20729 14153 20786 14199
rect 20832 14153 20889 14199
rect 20935 14153 20992 14199
rect 21038 14153 21051 14199
rect 7493 14066 7506 14112
rect 7552 14066 7623 14112
rect 7669 14066 7740 14112
rect 7786 14066 7858 14112
rect 7904 14066 7976 14112
rect 8022 14066 8094 14112
rect 8140 14066 8153 14112
rect 7493 14037 8153 14066
rect 3268 13975 4268 14004
rect 3268 13929 3281 13975
rect 3327 13929 3384 13975
rect 3430 13929 3487 13975
rect 3533 13929 3590 13975
rect 3636 13929 3693 13975
rect 3739 13929 3796 13975
rect 3842 13929 3899 13975
rect 3945 13929 4002 13975
rect 4048 13929 4105 13975
rect 4151 13929 4209 13975
rect 4255 13929 4268 13975
rect 3268 13868 4268 13929
rect 20051 14124 21051 14153
rect 7493 13888 8153 13917
rect 7493 13842 7506 13888
rect 7552 13842 7623 13888
rect 7669 13842 7740 13888
rect 7786 13842 7858 13888
rect 7904 13842 7976 13888
rect 8022 13842 8094 13888
rect 8140 13842 8153 13888
rect 7493 13813 8153 13842
rect 9195 13888 9327 13901
rect 9195 13842 9238 13888
rect 9284 13842 9327 13888
rect 9195 13813 9327 13842
rect 20051 13975 21051 14004
rect 20051 13929 20064 13975
rect 20110 13929 20168 13975
rect 20214 13929 20271 13975
rect 20317 13929 20374 13975
rect 20420 13929 20477 13975
rect 20523 13929 20580 13975
rect 20626 13929 20683 13975
rect 20729 13929 20786 13975
rect 20832 13929 20889 13975
rect 20935 13929 20992 13975
rect 21038 13929 21051 13975
rect 20051 13868 21051 13929
rect 7493 13664 8153 13693
rect 7493 13618 7506 13664
rect 7552 13618 7623 13664
rect 7669 13618 7740 13664
rect 7786 13618 7858 13664
rect 7904 13618 7976 13664
rect 8022 13618 8094 13664
rect 8140 13618 8153 13664
rect 7493 13605 8153 13618
rect 9195 13664 9327 13693
rect 9195 13618 9238 13664
rect 9284 13618 9327 13664
rect 9195 13605 9327 13618
rect 7493 13382 8153 13395
rect 7493 13336 7506 13382
rect 7552 13336 7623 13382
rect 7669 13336 7740 13382
rect 7786 13336 7858 13382
rect 7904 13336 7976 13382
rect 8022 13336 8094 13382
rect 8140 13336 8153 13382
rect 7493 13307 8153 13336
rect 9195 13382 9327 13395
rect 9195 13336 9238 13382
rect 9284 13336 9327 13382
rect 9195 13307 9327 13336
rect 3268 13071 4268 13132
rect 3268 13025 3281 13071
rect 3327 13025 3384 13071
rect 3430 13025 3487 13071
rect 3533 13025 3590 13071
rect 3636 13025 3693 13071
rect 3739 13025 3796 13071
rect 3842 13025 3899 13071
rect 3945 13025 4002 13071
rect 4048 13025 4105 13071
rect 4151 13025 4209 13071
rect 4255 13025 4268 13071
rect 3268 12996 4268 13025
rect 7493 13158 8153 13187
rect 7493 13112 7506 13158
rect 7552 13112 7623 13158
rect 7669 13112 7740 13158
rect 7786 13112 7858 13158
rect 7904 13112 7976 13158
rect 8022 13112 8094 13158
rect 8140 13112 8153 13158
rect 7493 13083 8153 13112
rect 9195 13158 9327 13187
rect 9195 13112 9238 13158
rect 9284 13112 9327 13158
rect 9195 13099 9327 13112
rect 3268 12847 4268 12876
rect 7493 12934 8153 12963
rect 7493 12888 7506 12934
rect 7552 12888 7623 12934
rect 7669 12888 7740 12934
rect 7786 12888 7858 12934
rect 7904 12888 7976 12934
rect 8022 12888 8094 12934
rect 8140 12888 8153 12934
rect 7493 12875 8153 12888
rect 20051 13071 21051 13132
rect 20051 13025 20064 13071
rect 20110 13025 20168 13071
rect 20214 13025 20271 13071
rect 20317 13025 20374 13071
rect 20420 13025 20477 13071
rect 20523 13025 20580 13071
rect 20626 13025 20683 13071
rect 20729 13025 20786 13071
rect 20832 13025 20889 13071
rect 20935 13025 20992 13071
rect 21038 13025 21051 13071
rect 20051 12996 21051 13025
rect 3268 12801 3281 12847
rect 3327 12801 3384 12847
rect 3430 12801 3487 12847
rect 3533 12801 3590 12847
rect 3636 12801 3693 12847
rect 3739 12801 3796 12847
rect 3842 12801 3899 12847
rect 3945 12801 4002 12847
rect 4048 12801 4105 12847
rect 4151 12801 4209 12847
rect 4255 12801 4268 12847
rect 3268 12772 4268 12801
rect 9324 12847 9764 12860
rect 9324 12801 9337 12847
rect 9383 12801 9459 12847
rect 9505 12801 9582 12847
rect 9628 12801 9705 12847
rect 9751 12801 9764 12847
rect 9324 12772 9764 12801
rect 20051 12847 21051 12876
rect 3268 12623 4268 12652
rect 3268 12577 3281 12623
rect 3327 12577 3384 12623
rect 3430 12577 3487 12623
rect 3533 12577 3590 12623
rect 3636 12577 3693 12623
rect 3739 12577 3796 12623
rect 3842 12577 3899 12623
rect 3945 12577 4002 12623
rect 4048 12577 4105 12623
rect 4151 12577 4209 12623
rect 4255 12577 4268 12623
rect 3268 12548 4268 12577
rect 9324 12623 9764 12652
rect 9324 12577 9337 12623
rect 9383 12577 9459 12623
rect 9505 12577 9582 12623
rect 9628 12577 9705 12623
rect 9751 12577 9764 12623
rect 9324 12548 9764 12577
rect 20051 12801 20064 12847
rect 20110 12801 20168 12847
rect 20214 12801 20271 12847
rect 20317 12801 20374 12847
rect 20420 12801 20477 12847
rect 20523 12801 20580 12847
rect 20626 12801 20683 12847
rect 20729 12801 20786 12847
rect 20832 12801 20889 12847
rect 20935 12801 20992 12847
rect 21038 12801 21051 12847
rect 20051 12772 21051 12801
rect 3268 12399 4268 12428
rect 3268 12353 3281 12399
rect 3327 12353 3384 12399
rect 3430 12353 3487 12399
rect 3533 12353 3590 12399
rect 3636 12353 3693 12399
rect 3739 12353 3796 12399
rect 3842 12353 3899 12399
rect 3945 12353 4002 12399
rect 4048 12353 4105 12399
rect 4151 12353 4209 12399
rect 4255 12353 4268 12399
rect 3268 12324 4268 12353
rect 9324 12399 9764 12428
rect 9324 12353 9337 12399
rect 9383 12353 9459 12399
rect 9505 12353 9582 12399
rect 9628 12353 9705 12399
rect 9751 12353 9764 12399
rect 9324 12340 9764 12353
rect 20051 12623 21051 12652
rect 20051 12577 20064 12623
rect 20110 12577 20168 12623
rect 20214 12577 20271 12623
rect 20317 12577 20374 12623
rect 20420 12577 20477 12623
rect 20523 12577 20580 12623
rect 20626 12577 20683 12623
rect 20729 12577 20786 12623
rect 20832 12577 20889 12623
rect 20935 12577 20992 12623
rect 21038 12577 21051 12623
rect 20051 12548 21051 12577
rect 7493 12312 8153 12325
rect 20051 12399 21051 12428
rect 20051 12353 20064 12399
rect 20110 12353 20168 12399
rect 20214 12353 20271 12399
rect 20317 12353 20374 12399
rect 20420 12353 20477 12399
rect 20523 12353 20580 12399
rect 20626 12353 20683 12399
rect 20729 12353 20786 12399
rect 20832 12353 20889 12399
rect 20935 12353 20992 12399
rect 21038 12353 21051 12399
rect 7493 12266 7506 12312
rect 7552 12266 7623 12312
rect 7669 12266 7740 12312
rect 7786 12266 7858 12312
rect 7904 12266 7976 12312
rect 8022 12266 8094 12312
rect 8140 12266 8153 12312
rect 7493 12237 8153 12266
rect 3268 12175 4268 12204
rect 3268 12129 3281 12175
rect 3327 12129 3384 12175
rect 3430 12129 3487 12175
rect 3533 12129 3590 12175
rect 3636 12129 3693 12175
rect 3739 12129 3796 12175
rect 3842 12129 3899 12175
rect 3945 12129 4002 12175
rect 4048 12129 4105 12175
rect 4151 12129 4209 12175
rect 4255 12129 4268 12175
rect 3268 12068 4268 12129
rect 20051 12324 21051 12353
rect 7493 12088 8153 12117
rect 7493 12042 7506 12088
rect 7552 12042 7623 12088
rect 7669 12042 7740 12088
rect 7786 12042 7858 12088
rect 7904 12042 7976 12088
rect 8022 12042 8094 12088
rect 8140 12042 8153 12088
rect 7493 12013 8153 12042
rect 9195 12088 9327 12101
rect 9195 12042 9238 12088
rect 9284 12042 9327 12088
rect 9195 12013 9327 12042
rect 20051 12175 21051 12204
rect 20051 12129 20064 12175
rect 20110 12129 20168 12175
rect 20214 12129 20271 12175
rect 20317 12129 20374 12175
rect 20420 12129 20477 12175
rect 20523 12129 20580 12175
rect 20626 12129 20683 12175
rect 20729 12129 20786 12175
rect 20832 12129 20889 12175
rect 20935 12129 20992 12175
rect 21038 12129 21051 12175
rect 20051 12068 21051 12129
rect 7493 11864 8153 11893
rect 7493 11818 7506 11864
rect 7552 11818 7623 11864
rect 7669 11818 7740 11864
rect 7786 11818 7858 11864
rect 7904 11818 7976 11864
rect 8022 11818 8094 11864
rect 8140 11818 8153 11864
rect 7493 11805 8153 11818
rect 9195 11864 9327 11893
rect 9195 11818 9238 11864
rect 9284 11818 9327 11864
rect 9195 11805 9327 11818
rect 7493 11582 8153 11595
rect 7493 11536 7506 11582
rect 7552 11536 7623 11582
rect 7669 11536 7740 11582
rect 7786 11536 7858 11582
rect 7904 11536 7976 11582
rect 8022 11536 8094 11582
rect 8140 11536 8153 11582
rect 7493 11507 8153 11536
rect 9195 11582 9327 11595
rect 9195 11536 9238 11582
rect 9284 11536 9327 11582
rect 9195 11507 9327 11536
rect 3268 11271 4268 11332
rect 3268 11225 3281 11271
rect 3327 11225 3384 11271
rect 3430 11225 3487 11271
rect 3533 11225 3590 11271
rect 3636 11225 3693 11271
rect 3739 11225 3796 11271
rect 3842 11225 3899 11271
rect 3945 11225 4002 11271
rect 4048 11225 4105 11271
rect 4151 11225 4209 11271
rect 4255 11225 4268 11271
rect 3268 11196 4268 11225
rect 7493 11358 8153 11387
rect 7493 11312 7506 11358
rect 7552 11312 7623 11358
rect 7669 11312 7740 11358
rect 7786 11312 7858 11358
rect 7904 11312 7976 11358
rect 8022 11312 8094 11358
rect 8140 11312 8153 11358
rect 7493 11283 8153 11312
rect 9195 11358 9327 11387
rect 9195 11312 9238 11358
rect 9284 11312 9327 11358
rect 9195 11299 9327 11312
rect 3268 11047 4268 11076
rect 7493 11134 8153 11163
rect 7493 11088 7506 11134
rect 7552 11088 7623 11134
rect 7669 11088 7740 11134
rect 7786 11088 7858 11134
rect 7904 11088 7976 11134
rect 8022 11088 8094 11134
rect 8140 11088 8153 11134
rect 7493 11075 8153 11088
rect 20051 11271 21051 11332
rect 20051 11225 20064 11271
rect 20110 11225 20168 11271
rect 20214 11225 20271 11271
rect 20317 11225 20374 11271
rect 20420 11225 20477 11271
rect 20523 11225 20580 11271
rect 20626 11225 20683 11271
rect 20729 11225 20786 11271
rect 20832 11225 20889 11271
rect 20935 11225 20992 11271
rect 21038 11225 21051 11271
rect 20051 11196 21051 11225
rect 3268 11001 3281 11047
rect 3327 11001 3384 11047
rect 3430 11001 3487 11047
rect 3533 11001 3590 11047
rect 3636 11001 3693 11047
rect 3739 11001 3796 11047
rect 3842 11001 3899 11047
rect 3945 11001 4002 11047
rect 4048 11001 4105 11047
rect 4151 11001 4209 11047
rect 4255 11001 4268 11047
rect 3268 10972 4268 11001
rect 9324 11047 9764 11060
rect 9324 11001 9337 11047
rect 9383 11001 9459 11047
rect 9505 11001 9582 11047
rect 9628 11001 9705 11047
rect 9751 11001 9764 11047
rect 9324 10972 9764 11001
rect 20051 11047 21051 11076
rect 3268 10823 4268 10852
rect 3268 10777 3281 10823
rect 3327 10777 3384 10823
rect 3430 10777 3487 10823
rect 3533 10777 3590 10823
rect 3636 10777 3693 10823
rect 3739 10777 3796 10823
rect 3842 10777 3899 10823
rect 3945 10777 4002 10823
rect 4048 10777 4105 10823
rect 4151 10777 4209 10823
rect 4255 10777 4268 10823
rect 3268 10748 4268 10777
rect 9324 10823 9764 10852
rect 9324 10777 9337 10823
rect 9383 10777 9459 10823
rect 9505 10777 9582 10823
rect 9628 10777 9705 10823
rect 9751 10777 9764 10823
rect 9324 10748 9764 10777
rect 20051 11001 20064 11047
rect 20110 11001 20168 11047
rect 20214 11001 20271 11047
rect 20317 11001 20374 11047
rect 20420 11001 20477 11047
rect 20523 11001 20580 11047
rect 20626 11001 20683 11047
rect 20729 11001 20786 11047
rect 20832 11001 20889 11047
rect 20935 11001 20992 11047
rect 21038 11001 21051 11047
rect 20051 10972 21051 11001
rect 3268 10599 4268 10628
rect 3268 10553 3281 10599
rect 3327 10553 3384 10599
rect 3430 10553 3487 10599
rect 3533 10553 3590 10599
rect 3636 10553 3693 10599
rect 3739 10553 3796 10599
rect 3842 10553 3899 10599
rect 3945 10553 4002 10599
rect 4048 10553 4105 10599
rect 4151 10553 4209 10599
rect 4255 10553 4268 10599
rect 3268 10524 4268 10553
rect 9324 10599 9764 10628
rect 9324 10553 9337 10599
rect 9383 10553 9459 10599
rect 9505 10553 9582 10599
rect 9628 10553 9705 10599
rect 9751 10553 9764 10599
rect 9324 10540 9764 10553
rect 20051 10823 21051 10852
rect 20051 10777 20064 10823
rect 20110 10777 20168 10823
rect 20214 10777 20271 10823
rect 20317 10777 20374 10823
rect 20420 10777 20477 10823
rect 20523 10777 20580 10823
rect 20626 10777 20683 10823
rect 20729 10777 20786 10823
rect 20832 10777 20889 10823
rect 20935 10777 20992 10823
rect 21038 10777 21051 10823
rect 20051 10748 21051 10777
rect 7493 10512 8153 10525
rect 20051 10599 21051 10628
rect 20051 10553 20064 10599
rect 20110 10553 20168 10599
rect 20214 10553 20271 10599
rect 20317 10553 20374 10599
rect 20420 10553 20477 10599
rect 20523 10553 20580 10599
rect 20626 10553 20683 10599
rect 20729 10553 20786 10599
rect 20832 10553 20889 10599
rect 20935 10553 20992 10599
rect 21038 10553 21051 10599
rect 7493 10466 7506 10512
rect 7552 10466 7623 10512
rect 7669 10466 7740 10512
rect 7786 10466 7858 10512
rect 7904 10466 7976 10512
rect 8022 10466 8094 10512
rect 8140 10466 8153 10512
rect 7493 10437 8153 10466
rect 3268 10375 4268 10404
rect 3268 10329 3281 10375
rect 3327 10329 3384 10375
rect 3430 10329 3487 10375
rect 3533 10329 3590 10375
rect 3636 10329 3693 10375
rect 3739 10329 3796 10375
rect 3842 10329 3899 10375
rect 3945 10329 4002 10375
rect 4048 10329 4105 10375
rect 4151 10329 4209 10375
rect 4255 10329 4268 10375
rect 3268 10268 4268 10329
rect 20051 10524 21051 10553
rect 7493 10288 8153 10317
rect 7493 10242 7506 10288
rect 7552 10242 7623 10288
rect 7669 10242 7740 10288
rect 7786 10242 7858 10288
rect 7904 10242 7976 10288
rect 8022 10242 8094 10288
rect 8140 10242 8153 10288
rect 7493 10213 8153 10242
rect 9195 10288 9327 10301
rect 9195 10242 9238 10288
rect 9284 10242 9327 10288
rect 9195 10213 9327 10242
rect 20051 10375 21051 10404
rect 20051 10329 20064 10375
rect 20110 10329 20168 10375
rect 20214 10329 20271 10375
rect 20317 10329 20374 10375
rect 20420 10329 20477 10375
rect 20523 10329 20580 10375
rect 20626 10329 20683 10375
rect 20729 10329 20786 10375
rect 20832 10329 20889 10375
rect 20935 10329 20992 10375
rect 21038 10329 21051 10375
rect 20051 10268 21051 10329
rect 7493 10064 8153 10093
rect 7493 10018 7506 10064
rect 7552 10018 7623 10064
rect 7669 10018 7740 10064
rect 7786 10018 7858 10064
rect 7904 10018 7976 10064
rect 8022 10018 8094 10064
rect 8140 10018 8153 10064
rect 7493 10005 8153 10018
rect 9195 10064 9327 10093
rect 9195 10018 9238 10064
rect 9284 10018 9327 10064
rect 9195 10005 9327 10018
rect 7493 9782 8153 9795
rect 7493 9736 7506 9782
rect 7552 9736 7623 9782
rect 7669 9736 7740 9782
rect 7786 9736 7858 9782
rect 7904 9736 7976 9782
rect 8022 9736 8094 9782
rect 8140 9736 8153 9782
rect 7493 9707 8153 9736
rect 9195 9782 9327 9795
rect 9195 9736 9238 9782
rect 9284 9736 9327 9782
rect 9195 9707 9327 9736
rect 3268 9471 4268 9532
rect 3268 9425 3281 9471
rect 3327 9425 3384 9471
rect 3430 9425 3487 9471
rect 3533 9425 3590 9471
rect 3636 9425 3693 9471
rect 3739 9425 3796 9471
rect 3842 9425 3899 9471
rect 3945 9425 4002 9471
rect 4048 9425 4105 9471
rect 4151 9425 4209 9471
rect 4255 9425 4268 9471
rect 3268 9396 4268 9425
rect 7493 9558 8153 9587
rect 7493 9512 7506 9558
rect 7552 9512 7623 9558
rect 7669 9512 7740 9558
rect 7786 9512 7858 9558
rect 7904 9512 7976 9558
rect 8022 9512 8094 9558
rect 8140 9512 8153 9558
rect 7493 9483 8153 9512
rect 9195 9558 9327 9587
rect 9195 9512 9238 9558
rect 9284 9512 9327 9558
rect 9195 9499 9327 9512
rect 3268 9247 4268 9276
rect 7493 9334 8153 9363
rect 7493 9288 7506 9334
rect 7552 9288 7623 9334
rect 7669 9288 7740 9334
rect 7786 9288 7858 9334
rect 7904 9288 7976 9334
rect 8022 9288 8094 9334
rect 8140 9288 8153 9334
rect 7493 9275 8153 9288
rect 20051 9471 21051 9532
rect 20051 9425 20064 9471
rect 20110 9425 20168 9471
rect 20214 9425 20271 9471
rect 20317 9425 20374 9471
rect 20420 9425 20477 9471
rect 20523 9425 20580 9471
rect 20626 9425 20683 9471
rect 20729 9425 20786 9471
rect 20832 9425 20889 9471
rect 20935 9425 20992 9471
rect 21038 9425 21051 9471
rect 20051 9396 21051 9425
rect 3268 9201 3281 9247
rect 3327 9201 3384 9247
rect 3430 9201 3487 9247
rect 3533 9201 3590 9247
rect 3636 9201 3693 9247
rect 3739 9201 3796 9247
rect 3842 9201 3899 9247
rect 3945 9201 4002 9247
rect 4048 9201 4105 9247
rect 4151 9201 4209 9247
rect 4255 9201 4268 9247
rect 3268 9172 4268 9201
rect 9324 9247 9764 9260
rect 9324 9201 9337 9247
rect 9383 9201 9459 9247
rect 9505 9201 9582 9247
rect 9628 9201 9705 9247
rect 9751 9201 9764 9247
rect 9324 9172 9764 9201
rect 20051 9247 21051 9276
rect 3268 9023 4268 9052
rect 3268 8977 3281 9023
rect 3327 8977 3384 9023
rect 3430 8977 3487 9023
rect 3533 8977 3590 9023
rect 3636 8977 3693 9023
rect 3739 8977 3796 9023
rect 3842 8977 3899 9023
rect 3945 8977 4002 9023
rect 4048 8977 4105 9023
rect 4151 8977 4209 9023
rect 4255 8977 4268 9023
rect 3268 8948 4268 8977
rect 9324 9023 9764 9052
rect 9324 8977 9337 9023
rect 9383 8977 9459 9023
rect 9505 8977 9582 9023
rect 9628 8977 9705 9023
rect 9751 8977 9764 9023
rect 9324 8948 9764 8977
rect 20051 9201 20064 9247
rect 20110 9201 20168 9247
rect 20214 9201 20271 9247
rect 20317 9201 20374 9247
rect 20420 9201 20477 9247
rect 20523 9201 20580 9247
rect 20626 9201 20683 9247
rect 20729 9201 20786 9247
rect 20832 9201 20889 9247
rect 20935 9201 20992 9247
rect 21038 9201 21051 9247
rect 20051 9172 21051 9201
rect 3268 8799 4268 8828
rect 3268 8753 3281 8799
rect 3327 8753 3384 8799
rect 3430 8753 3487 8799
rect 3533 8753 3590 8799
rect 3636 8753 3693 8799
rect 3739 8753 3796 8799
rect 3842 8753 3899 8799
rect 3945 8753 4002 8799
rect 4048 8753 4105 8799
rect 4151 8753 4209 8799
rect 4255 8753 4268 8799
rect 3268 8724 4268 8753
rect 9324 8799 9764 8828
rect 9324 8753 9337 8799
rect 9383 8753 9459 8799
rect 9505 8753 9582 8799
rect 9628 8753 9705 8799
rect 9751 8753 9764 8799
rect 9324 8740 9764 8753
rect 20051 9023 21051 9052
rect 20051 8977 20064 9023
rect 20110 8977 20168 9023
rect 20214 8977 20271 9023
rect 20317 8977 20374 9023
rect 20420 8977 20477 9023
rect 20523 8977 20580 9023
rect 20626 8977 20683 9023
rect 20729 8977 20786 9023
rect 20832 8977 20889 9023
rect 20935 8977 20992 9023
rect 21038 8977 21051 9023
rect 20051 8948 21051 8977
rect 7493 8712 8153 8725
rect 20051 8799 21051 8828
rect 20051 8753 20064 8799
rect 20110 8753 20168 8799
rect 20214 8753 20271 8799
rect 20317 8753 20374 8799
rect 20420 8753 20477 8799
rect 20523 8753 20580 8799
rect 20626 8753 20683 8799
rect 20729 8753 20786 8799
rect 20832 8753 20889 8799
rect 20935 8753 20992 8799
rect 21038 8753 21051 8799
rect 7493 8666 7506 8712
rect 7552 8666 7623 8712
rect 7669 8666 7740 8712
rect 7786 8666 7858 8712
rect 7904 8666 7976 8712
rect 8022 8666 8094 8712
rect 8140 8666 8153 8712
rect 7493 8637 8153 8666
rect 3268 8575 4268 8604
rect 3268 8529 3281 8575
rect 3327 8529 3384 8575
rect 3430 8529 3487 8575
rect 3533 8529 3590 8575
rect 3636 8529 3693 8575
rect 3739 8529 3796 8575
rect 3842 8529 3899 8575
rect 3945 8529 4002 8575
rect 4048 8529 4105 8575
rect 4151 8529 4209 8575
rect 4255 8529 4268 8575
rect 3268 8468 4268 8529
rect 20051 8724 21051 8753
rect 7493 8488 8153 8517
rect 7493 8442 7506 8488
rect 7552 8442 7623 8488
rect 7669 8442 7740 8488
rect 7786 8442 7858 8488
rect 7904 8442 7976 8488
rect 8022 8442 8094 8488
rect 8140 8442 8153 8488
rect 7493 8413 8153 8442
rect 9195 8488 9327 8501
rect 9195 8442 9238 8488
rect 9284 8442 9327 8488
rect 9195 8413 9327 8442
rect 20051 8575 21051 8604
rect 20051 8529 20064 8575
rect 20110 8529 20168 8575
rect 20214 8529 20271 8575
rect 20317 8529 20374 8575
rect 20420 8529 20477 8575
rect 20523 8529 20580 8575
rect 20626 8529 20683 8575
rect 20729 8529 20786 8575
rect 20832 8529 20889 8575
rect 20935 8529 20992 8575
rect 21038 8529 21051 8575
rect 20051 8468 21051 8529
rect 7493 8264 8153 8293
rect 7493 8218 7506 8264
rect 7552 8218 7623 8264
rect 7669 8218 7740 8264
rect 7786 8218 7858 8264
rect 7904 8218 7976 8264
rect 8022 8218 8094 8264
rect 8140 8218 8153 8264
rect 7493 8205 8153 8218
rect 9195 8264 9327 8293
rect 9195 8218 9238 8264
rect 9284 8218 9327 8264
rect 9195 8205 9327 8218
rect 7493 7982 8153 7995
rect 7493 7936 7506 7982
rect 7552 7936 7623 7982
rect 7669 7936 7740 7982
rect 7786 7936 7858 7982
rect 7904 7936 7976 7982
rect 8022 7936 8094 7982
rect 8140 7936 8153 7982
rect 7493 7907 8153 7936
rect 9195 7982 9327 7995
rect 9195 7936 9238 7982
rect 9284 7936 9327 7982
rect 9195 7907 9327 7936
rect 3268 7671 4268 7732
rect 3268 7625 3281 7671
rect 3327 7625 3384 7671
rect 3430 7625 3487 7671
rect 3533 7625 3590 7671
rect 3636 7625 3693 7671
rect 3739 7625 3796 7671
rect 3842 7625 3899 7671
rect 3945 7625 4002 7671
rect 4048 7625 4105 7671
rect 4151 7625 4209 7671
rect 4255 7625 4268 7671
rect 3268 7596 4268 7625
rect 7493 7758 8153 7787
rect 7493 7712 7506 7758
rect 7552 7712 7623 7758
rect 7669 7712 7740 7758
rect 7786 7712 7858 7758
rect 7904 7712 7976 7758
rect 8022 7712 8094 7758
rect 8140 7712 8153 7758
rect 7493 7683 8153 7712
rect 9195 7758 9327 7787
rect 9195 7712 9238 7758
rect 9284 7712 9327 7758
rect 9195 7699 9327 7712
rect 3268 7447 4268 7476
rect 7493 7534 8153 7563
rect 7493 7488 7506 7534
rect 7552 7488 7623 7534
rect 7669 7488 7740 7534
rect 7786 7488 7858 7534
rect 7904 7488 7976 7534
rect 8022 7488 8094 7534
rect 8140 7488 8153 7534
rect 7493 7475 8153 7488
rect 20051 7671 21051 7732
rect 20051 7625 20064 7671
rect 20110 7625 20168 7671
rect 20214 7625 20271 7671
rect 20317 7625 20374 7671
rect 20420 7625 20477 7671
rect 20523 7625 20580 7671
rect 20626 7625 20683 7671
rect 20729 7625 20786 7671
rect 20832 7625 20889 7671
rect 20935 7625 20992 7671
rect 21038 7625 21051 7671
rect 20051 7596 21051 7625
rect 3268 7401 3281 7447
rect 3327 7401 3384 7447
rect 3430 7401 3487 7447
rect 3533 7401 3590 7447
rect 3636 7401 3693 7447
rect 3739 7401 3796 7447
rect 3842 7401 3899 7447
rect 3945 7401 4002 7447
rect 4048 7401 4105 7447
rect 4151 7401 4209 7447
rect 4255 7401 4268 7447
rect 3268 7372 4268 7401
rect 9324 7447 9764 7460
rect 9324 7401 9337 7447
rect 9383 7401 9459 7447
rect 9505 7401 9582 7447
rect 9628 7401 9705 7447
rect 9751 7401 9764 7447
rect 9324 7372 9764 7401
rect 20051 7447 21051 7476
rect 3268 7223 4268 7252
rect 3268 7177 3281 7223
rect 3327 7177 3384 7223
rect 3430 7177 3487 7223
rect 3533 7177 3590 7223
rect 3636 7177 3693 7223
rect 3739 7177 3796 7223
rect 3842 7177 3899 7223
rect 3945 7177 4002 7223
rect 4048 7177 4105 7223
rect 4151 7177 4209 7223
rect 4255 7177 4268 7223
rect 3268 7148 4268 7177
rect 9324 7223 9764 7252
rect 9324 7177 9337 7223
rect 9383 7177 9459 7223
rect 9505 7177 9582 7223
rect 9628 7177 9705 7223
rect 9751 7177 9764 7223
rect 9324 7148 9764 7177
rect 20051 7401 20064 7447
rect 20110 7401 20168 7447
rect 20214 7401 20271 7447
rect 20317 7401 20374 7447
rect 20420 7401 20477 7447
rect 20523 7401 20580 7447
rect 20626 7401 20683 7447
rect 20729 7401 20786 7447
rect 20832 7401 20889 7447
rect 20935 7401 20992 7447
rect 21038 7401 21051 7447
rect 20051 7372 21051 7401
rect 3268 6999 4268 7028
rect 3268 6953 3281 6999
rect 3327 6953 3384 6999
rect 3430 6953 3487 6999
rect 3533 6953 3590 6999
rect 3636 6953 3693 6999
rect 3739 6953 3796 6999
rect 3842 6953 3899 6999
rect 3945 6953 4002 6999
rect 4048 6953 4105 6999
rect 4151 6953 4209 6999
rect 4255 6953 4268 6999
rect 3268 6924 4268 6953
rect 9324 6999 9764 7028
rect 9324 6953 9337 6999
rect 9383 6953 9459 6999
rect 9505 6953 9582 6999
rect 9628 6953 9705 6999
rect 9751 6953 9764 6999
rect 9324 6940 9764 6953
rect 20051 7223 21051 7252
rect 20051 7177 20064 7223
rect 20110 7177 20168 7223
rect 20214 7177 20271 7223
rect 20317 7177 20374 7223
rect 20420 7177 20477 7223
rect 20523 7177 20580 7223
rect 20626 7177 20683 7223
rect 20729 7177 20786 7223
rect 20832 7177 20889 7223
rect 20935 7177 20992 7223
rect 21038 7177 21051 7223
rect 20051 7148 21051 7177
rect 7493 6912 8153 6925
rect 20051 6999 21051 7028
rect 20051 6953 20064 6999
rect 20110 6953 20168 6999
rect 20214 6953 20271 6999
rect 20317 6953 20374 6999
rect 20420 6953 20477 6999
rect 20523 6953 20580 6999
rect 20626 6953 20683 6999
rect 20729 6953 20786 6999
rect 20832 6953 20889 6999
rect 20935 6953 20992 6999
rect 21038 6953 21051 6999
rect 7493 6866 7506 6912
rect 7552 6866 7623 6912
rect 7669 6866 7740 6912
rect 7786 6866 7858 6912
rect 7904 6866 7976 6912
rect 8022 6866 8094 6912
rect 8140 6866 8153 6912
rect 7493 6837 8153 6866
rect 3268 6775 4268 6804
rect 3268 6729 3281 6775
rect 3327 6729 3384 6775
rect 3430 6729 3487 6775
rect 3533 6729 3590 6775
rect 3636 6729 3693 6775
rect 3739 6729 3796 6775
rect 3842 6729 3899 6775
rect 3945 6729 4002 6775
rect 4048 6729 4105 6775
rect 4151 6729 4209 6775
rect 4255 6729 4268 6775
rect 3268 6668 4268 6729
rect 20051 6924 21051 6953
rect 7493 6688 8153 6717
rect 7493 6642 7506 6688
rect 7552 6642 7623 6688
rect 7669 6642 7740 6688
rect 7786 6642 7858 6688
rect 7904 6642 7976 6688
rect 8022 6642 8094 6688
rect 8140 6642 8153 6688
rect 7493 6613 8153 6642
rect 9195 6688 9327 6701
rect 9195 6642 9238 6688
rect 9284 6642 9327 6688
rect 9195 6613 9327 6642
rect 20051 6775 21051 6804
rect 20051 6729 20064 6775
rect 20110 6729 20168 6775
rect 20214 6729 20271 6775
rect 20317 6729 20374 6775
rect 20420 6729 20477 6775
rect 20523 6729 20580 6775
rect 20626 6729 20683 6775
rect 20729 6729 20786 6775
rect 20832 6729 20889 6775
rect 20935 6729 20992 6775
rect 21038 6729 21051 6775
rect 20051 6668 21051 6729
rect 7493 6464 8153 6493
rect 7493 6418 7506 6464
rect 7552 6418 7623 6464
rect 7669 6418 7740 6464
rect 7786 6418 7858 6464
rect 7904 6418 7976 6464
rect 8022 6418 8094 6464
rect 8140 6418 8153 6464
rect 7493 6405 8153 6418
rect 9195 6464 9327 6493
rect 9195 6418 9238 6464
rect 9284 6418 9327 6464
rect 9195 6405 9327 6418
rect 7493 6182 8153 6195
rect 7493 6136 7506 6182
rect 7552 6136 7623 6182
rect 7669 6136 7740 6182
rect 7786 6136 7858 6182
rect 7904 6136 7976 6182
rect 8022 6136 8094 6182
rect 8140 6136 8153 6182
rect 7493 6107 8153 6136
rect 9195 6182 9327 6195
rect 9195 6136 9238 6182
rect 9284 6136 9327 6182
rect 9195 6107 9327 6136
rect 3268 5871 4268 5932
rect 3268 5825 3281 5871
rect 3327 5825 3384 5871
rect 3430 5825 3487 5871
rect 3533 5825 3590 5871
rect 3636 5825 3693 5871
rect 3739 5825 3796 5871
rect 3842 5825 3899 5871
rect 3945 5825 4002 5871
rect 4048 5825 4105 5871
rect 4151 5825 4209 5871
rect 4255 5825 4268 5871
rect 3268 5796 4268 5825
rect 7493 5958 8153 5987
rect 7493 5912 7506 5958
rect 7552 5912 7623 5958
rect 7669 5912 7740 5958
rect 7786 5912 7858 5958
rect 7904 5912 7976 5958
rect 8022 5912 8094 5958
rect 8140 5912 8153 5958
rect 7493 5883 8153 5912
rect 9195 5958 9327 5987
rect 9195 5912 9238 5958
rect 9284 5912 9327 5958
rect 9195 5899 9327 5912
rect 3268 5647 4268 5676
rect 7493 5734 8153 5763
rect 7493 5688 7506 5734
rect 7552 5688 7623 5734
rect 7669 5688 7740 5734
rect 7786 5688 7858 5734
rect 7904 5688 7976 5734
rect 8022 5688 8094 5734
rect 8140 5688 8153 5734
rect 7493 5675 8153 5688
rect 20051 5871 21051 5932
rect 20051 5825 20064 5871
rect 20110 5825 20168 5871
rect 20214 5825 20271 5871
rect 20317 5825 20374 5871
rect 20420 5825 20477 5871
rect 20523 5825 20580 5871
rect 20626 5825 20683 5871
rect 20729 5825 20786 5871
rect 20832 5825 20889 5871
rect 20935 5825 20992 5871
rect 21038 5825 21051 5871
rect 20051 5796 21051 5825
rect 3268 5601 3281 5647
rect 3327 5601 3384 5647
rect 3430 5601 3487 5647
rect 3533 5601 3590 5647
rect 3636 5601 3693 5647
rect 3739 5601 3796 5647
rect 3842 5601 3899 5647
rect 3945 5601 4002 5647
rect 4048 5601 4105 5647
rect 4151 5601 4209 5647
rect 4255 5601 4268 5647
rect 3268 5572 4268 5601
rect 9324 5647 9764 5660
rect 9324 5601 9337 5647
rect 9383 5601 9459 5647
rect 9505 5601 9582 5647
rect 9628 5601 9705 5647
rect 9751 5601 9764 5647
rect 9324 5572 9764 5601
rect 20051 5647 21051 5676
rect 3268 5423 4268 5452
rect 3268 5377 3281 5423
rect 3327 5377 3384 5423
rect 3430 5377 3487 5423
rect 3533 5377 3590 5423
rect 3636 5377 3693 5423
rect 3739 5377 3796 5423
rect 3842 5377 3899 5423
rect 3945 5377 4002 5423
rect 4048 5377 4105 5423
rect 4151 5377 4209 5423
rect 4255 5377 4268 5423
rect 3268 5348 4268 5377
rect 9324 5423 9764 5452
rect 9324 5377 9337 5423
rect 9383 5377 9459 5423
rect 9505 5377 9582 5423
rect 9628 5377 9705 5423
rect 9751 5377 9764 5423
rect 9324 5348 9764 5377
rect 20051 5601 20064 5647
rect 20110 5601 20168 5647
rect 20214 5601 20271 5647
rect 20317 5601 20374 5647
rect 20420 5601 20477 5647
rect 20523 5601 20580 5647
rect 20626 5601 20683 5647
rect 20729 5601 20786 5647
rect 20832 5601 20889 5647
rect 20935 5601 20992 5647
rect 21038 5601 21051 5647
rect 20051 5572 21051 5601
rect 3268 5199 4268 5228
rect 3268 5153 3281 5199
rect 3327 5153 3384 5199
rect 3430 5153 3487 5199
rect 3533 5153 3590 5199
rect 3636 5153 3693 5199
rect 3739 5153 3796 5199
rect 3842 5153 3899 5199
rect 3945 5153 4002 5199
rect 4048 5153 4105 5199
rect 4151 5153 4209 5199
rect 4255 5153 4268 5199
rect 3268 5124 4268 5153
rect 9324 5199 9764 5228
rect 9324 5153 9337 5199
rect 9383 5153 9459 5199
rect 9505 5153 9582 5199
rect 9628 5153 9705 5199
rect 9751 5153 9764 5199
rect 9324 5140 9764 5153
rect 20051 5423 21051 5452
rect 20051 5377 20064 5423
rect 20110 5377 20168 5423
rect 20214 5377 20271 5423
rect 20317 5377 20374 5423
rect 20420 5377 20477 5423
rect 20523 5377 20580 5423
rect 20626 5377 20683 5423
rect 20729 5377 20786 5423
rect 20832 5377 20889 5423
rect 20935 5377 20992 5423
rect 21038 5377 21051 5423
rect 20051 5348 21051 5377
rect 7493 5112 8153 5125
rect 20051 5199 21051 5228
rect 20051 5153 20064 5199
rect 20110 5153 20168 5199
rect 20214 5153 20271 5199
rect 20317 5153 20374 5199
rect 20420 5153 20477 5199
rect 20523 5153 20580 5199
rect 20626 5153 20683 5199
rect 20729 5153 20786 5199
rect 20832 5153 20889 5199
rect 20935 5153 20992 5199
rect 21038 5153 21051 5199
rect 7493 5066 7506 5112
rect 7552 5066 7623 5112
rect 7669 5066 7740 5112
rect 7786 5066 7858 5112
rect 7904 5066 7976 5112
rect 8022 5066 8094 5112
rect 8140 5066 8153 5112
rect 7493 5037 8153 5066
rect 3268 4975 4268 5004
rect 3268 4929 3281 4975
rect 3327 4929 3384 4975
rect 3430 4929 3487 4975
rect 3533 4929 3590 4975
rect 3636 4929 3693 4975
rect 3739 4929 3796 4975
rect 3842 4929 3899 4975
rect 3945 4929 4002 4975
rect 4048 4929 4105 4975
rect 4151 4929 4209 4975
rect 4255 4929 4268 4975
rect 3268 4868 4268 4929
rect 20051 5124 21051 5153
rect 7493 4888 8153 4917
rect 7493 4842 7506 4888
rect 7552 4842 7623 4888
rect 7669 4842 7740 4888
rect 7786 4842 7858 4888
rect 7904 4842 7976 4888
rect 8022 4842 8094 4888
rect 8140 4842 8153 4888
rect 7493 4813 8153 4842
rect 9195 4888 9327 4901
rect 9195 4842 9238 4888
rect 9284 4842 9327 4888
rect 9195 4813 9327 4842
rect 20051 4975 21051 5004
rect 20051 4929 20064 4975
rect 20110 4929 20168 4975
rect 20214 4929 20271 4975
rect 20317 4929 20374 4975
rect 20420 4929 20477 4975
rect 20523 4929 20580 4975
rect 20626 4929 20683 4975
rect 20729 4929 20786 4975
rect 20832 4929 20889 4975
rect 20935 4929 20992 4975
rect 21038 4929 21051 4975
rect 20051 4868 21051 4929
rect 7493 4664 8153 4693
rect 7493 4618 7506 4664
rect 7552 4618 7623 4664
rect 7669 4618 7740 4664
rect 7786 4618 7858 4664
rect 7904 4618 7976 4664
rect 8022 4618 8094 4664
rect 8140 4618 8153 4664
rect 7493 4605 8153 4618
rect 9195 4664 9327 4693
rect 9195 4618 9238 4664
rect 9284 4618 9327 4664
rect 9195 4605 9327 4618
rect 7493 4382 8153 4395
rect 7493 4336 7506 4382
rect 7552 4336 7623 4382
rect 7669 4336 7740 4382
rect 7786 4336 7858 4382
rect 7904 4336 7976 4382
rect 8022 4336 8094 4382
rect 8140 4336 8153 4382
rect 7493 4307 8153 4336
rect 9195 4382 9327 4395
rect 9195 4336 9238 4382
rect 9284 4336 9327 4382
rect 9195 4307 9327 4336
rect 3268 4071 4268 4132
rect 3268 4025 3281 4071
rect 3327 4025 3384 4071
rect 3430 4025 3487 4071
rect 3533 4025 3590 4071
rect 3636 4025 3693 4071
rect 3739 4025 3796 4071
rect 3842 4025 3899 4071
rect 3945 4025 4002 4071
rect 4048 4025 4105 4071
rect 4151 4025 4209 4071
rect 4255 4025 4268 4071
rect 3268 3996 4268 4025
rect 7493 4158 8153 4187
rect 7493 4112 7506 4158
rect 7552 4112 7623 4158
rect 7669 4112 7740 4158
rect 7786 4112 7858 4158
rect 7904 4112 7976 4158
rect 8022 4112 8094 4158
rect 8140 4112 8153 4158
rect 7493 4083 8153 4112
rect 9195 4158 9327 4187
rect 9195 4112 9238 4158
rect 9284 4112 9327 4158
rect 9195 4099 9327 4112
rect 3268 3847 4268 3876
rect 7493 3934 8153 3963
rect 7493 3888 7506 3934
rect 7552 3888 7623 3934
rect 7669 3888 7740 3934
rect 7786 3888 7858 3934
rect 7904 3888 7976 3934
rect 8022 3888 8094 3934
rect 8140 3888 8153 3934
rect 7493 3875 8153 3888
rect 20051 4071 21051 4132
rect 20051 4025 20064 4071
rect 20110 4025 20168 4071
rect 20214 4025 20271 4071
rect 20317 4025 20374 4071
rect 20420 4025 20477 4071
rect 20523 4025 20580 4071
rect 20626 4025 20683 4071
rect 20729 4025 20786 4071
rect 20832 4025 20889 4071
rect 20935 4025 20992 4071
rect 21038 4025 21051 4071
rect 20051 3996 21051 4025
rect 3268 3801 3281 3847
rect 3327 3801 3384 3847
rect 3430 3801 3487 3847
rect 3533 3801 3590 3847
rect 3636 3801 3693 3847
rect 3739 3801 3796 3847
rect 3842 3801 3899 3847
rect 3945 3801 4002 3847
rect 4048 3801 4105 3847
rect 4151 3801 4209 3847
rect 4255 3801 4268 3847
rect 3268 3772 4268 3801
rect 9324 3847 9764 3860
rect 9324 3801 9337 3847
rect 9383 3801 9459 3847
rect 9505 3801 9582 3847
rect 9628 3801 9705 3847
rect 9751 3801 9764 3847
rect 9324 3772 9764 3801
rect 20051 3847 21051 3876
rect 3268 3623 4268 3652
rect 3268 3577 3281 3623
rect 3327 3577 3384 3623
rect 3430 3577 3487 3623
rect 3533 3577 3590 3623
rect 3636 3577 3693 3623
rect 3739 3577 3796 3623
rect 3842 3577 3899 3623
rect 3945 3577 4002 3623
rect 4048 3577 4105 3623
rect 4151 3577 4209 3623
rect 4255 3577 4268 3623
rect 3268 3548 4268 3577
rect 9324 3623 9764 3652
rect 9324 3577 9337 3623
rect 9383 3577 9459 3623
rect 9505 3577 9582 3623
rect 9628 3577 9705 3623
rect 9751 3577 9764 3623
rect 9324 3548 9764 3577
rect 20051 3801 20064 3847
rect 20110 3801 20168 3847
rect 20214 3801 20271 3847
rect 20317 3801 20374 3847
rect 20420 3801 20477 3847
rect 20523 3801 20580 3847
rect 20626 3801 20683 3847
rect 20729 3801 20786 3847
rect 20832 3801 20889 3847
rect 20935 3801 20992 3847
rect 21038 3801 21051 3847
rect 20051 3772 21051 3801
rect 3268 3399 4268 3428
rect 3268 3353 3281 3399
rect 3327 3353 3384 3399
rect 3430 3353 3487 3399
rect 3533 3353 3590 3399
rect 3636 3353 3693 3399
rect 3739 3353 3796 3399
rect 3842 3353 3899 3399
rect 3945 3353 4002 3399
rect 4048 3353 4105 3399
rect 4151 3353 4209 3399
rect 4255 3353 4268 3399
rect 3268 3324 4268 3353
rect 9324 3399 9764 3428
rect 9324 3353 9337 3399
rect 9383 3353 9459 3399
rect 9505 3353 9582 3399
rect 9628 3353 9705 3399
rect 9751 3353 9764 3399
rect 9324 3340 9764 3353
rect 20051 3623 21051 3652
rect 20051 3577 20064 3623
rect 20110 3577 20168 3623
rect 20214 3577 20271 3623
rect 20317 3577 20374 3623
rect 20420 3577 20477 3623
rect 20523 3577 20580 3623
rect 20626 3577 20683 3623
rect 20729 3577 20786 3623
rect 20832 3577 20889 3623
rect 20935 3577 20992 3623
rect 21038 3577 21051 3623
rect 20051 3548 21051 3577
rect 7493 3312 8153 3325
rect 20051 3399 21051 3428
rect 20051 3353 20064 3399
rect 20110 3353 20168 3399
rect 20214 3353 20271 3399
rect 20317 3353 20374 3399
rect 20420 3353 20477 3399
rect 20523 3353 20580 3399
rect 20626 3353 20683 3399
rect 20729 3353 20786 3399
rect 20832 3353 20889 3399
rect 20935 3353 20992 3399
rect 21038 3353 21051 3399
rect 7493 3266 7506 3312
rect 7552 3266 7623 3312
rect 7669 3266 7740 3312
rect 7786 3266 7858 3312
rect 7904 3266 7976 3312
rect 8022 3266 8094 3312
rect 8140 3266 8153 3312
rect 7493 3237 8153 3266
rect 3268 3175 4268 3204
rect 3268 3129 3281 3175
rect 3327 3129 3384 3175
rect 3430 3129 3487 3175
rect 3533 3129 3590 3175
rect 3636 3129 3693 3175
rect 3739 3129 3796 3175
rect 3842 3129 3899 3175
rect 3945 3129 4002 3175
rect 4048 3129 4105 3175
rect 4151 3129 4209 3175
rect 4255 3129 4268 3175
rect 3268 3068 4268 3129
rect 20051 3324 21051 3353
rect 7493 3088 8153 3117
rect 7493 3042 7506 3088
rect 7552 3042 7623 3088
rect 7669 3042 7740 3088
rect 7786 3042 7858 3088
rect 7904 3042 7976 3088
rect 8022 3042 8094 3088
rect 8140 3042 8153 3088
rect 7493 3013 8153 3042
rect 9195 3088 9327 3101
rect 9195 3042 9238 3088
rect 9284 3042 9327 3088
rect 9195 3013 9327 3042
rect 20051 3175 21051 3204
rect 20051 3129 20064 3175
rect 20110 3129 20168 3175
rect 20214 3129 20271 3175
rect 20317 3129 20374 3175
rect 20420 3129 20477 3175
rect 20523 3129 20580 3175
rect 20626 3129 20683 3175
rect 20729 3129 20786 3175
rect 20832 3129 20889 3175
rect 20935 3129 20992 3175
rect 21038 3129 21051 3175
rect 20051 3068 21051 3129
rect 7493 2864 8153 2893
rect 7493 2818 7506 2864
rect 7552 2818 7623 2864
rect 7669 2818 7740 2864
rect 7786 2818 7858 2864
rect 7904 2818 7976 2864
rect 8022 2818 8094 2864
rect 8140 2818 8153 2864
rect 7493 2805 8153 2818
rect 9195 2864 9327 2893
rect 9195 2818 9238 2864
rect 9284 2818 9327 2864
rect 9195 2805 9327 2818
rect 7493 2582 8153 2595
rect 7493 2536 7506 2582
rect 7552 2536 7623 2582
rect 7669 2536 7740 2582
rect 7786 2536 7858 2582
rect 7904 2536 7976 2582
rect 8022 2536 8094 2582
rect 8140 2536 8153 2582
rect 7493 2507 8153 2536
rect 9195 2582 9327 2595
rect 9195 2536 9238 2582
rect 9284 2536 9327 2582
rect 9195 2507 9327 2536
rect 3268 2271 4268 2332
rect 3268 2225 3281 2271
rect 3327 2225 3384 2271
rect 3430 2225 3487 2271
rect 3533 2225 3590 2271
rect 3636 2225 3693 2271
rect 3739 2225 3796 2271
rect 3842 2225 3899 2271
rect 3945 2225 4002 2271
rect 4048 2225 4105 2271
rect 4151 2225 4209 2271
rect 4255 2225 4268 2271
rect 3268 2196 4268 2225
rect 7493 2358 8153 2387
rect 7493 2312 7506 2358
rect 7552 2312 7623 2358
rect 7669 2312 7740 2358
rect 7786 2312 7858 2358
rect 7904 2312 7976 2358
rect 8022 2312 8094 2358
rect 8140 2312 8153 2358
rect 7493 2283 8153 2312
rect 9195 2358 9327 2387
rect 9195 2312 9238 2358
rect 9284 2312 9327 2358
rect 9195 2299 9327 2312
rect 3268 2047 4268 2076
rect 7493 2134 8153 2163
rect 7493 2088 7506 2134
rect 7552 2088 7623 2134
rect 7669 2088 7740 2134
rect 7786 2088 7858 2134
rect 7904 2088 7976 2134
rect 8022 2088 8094 2134
rect 8140 2088 8153 2134
rect 7493 2075 8153 2088
rect 20051 2271 21051 2332
rect 20051 2225 20064 2271
rect 20110 2225 20168 2271
rect 20214 2225 20271 2271
rect 20317 2225 20374 2271
rect 20420 2225 20477 2271
rect 20523 2225 20580 2271
rect 20626 2225 20683 2271
rect 20729 2225 20786 2271
rect 20832 2225 20889 2271
rect 20935 2225 20992 2271
rect 21038 2225 21051 2271
rect 20051 2196 21051 2225
rect 3268 2001 3281 2047
rect 3327 2001 3384 2047
rect 3430 2001 3487 2047
rect 3533 2001 3590 2047
rect 3636 2001 3693 2047
rect 3739 2001 3796 2047
rect 3842 2001 3899 2047
rect 3945 2001 4002 2047
rect 4048 2001 4105 2047
rect 4151 2001 4209 2047
rect 4255 2001 4268 2047
rect 3268 1972 4268 2001
rect 9324 2047 9764 2060
rect 9324 2001 9337 2047
rect 9383 2001 9459 2047
rect 9505 2001 9582 2047
rect 9628 2001 9705 2047
rect 9751 2001 9764 2047
rect 9324 1972 9764 2001
rect 20051 2047 21051 2076
rect 3268 1823 4268 1852
rect 3268 1777 3281 1823
rect 3327 1777 3384 1823
rect 3430 1777 3487 1823
rect 3533 1777 3590 1823
rect 3636 1777 3693 1823
rect 3739 1777 3796 1823
rect 3842 1777 3899 1823
rect 3945 1777 4002 1823
rect 4048 1777 4105 1823
rect 4151 1777 4209 1823
rect 4255 1777 4268 1823
rect 3268 1748 4268 1777
rect 9324 1823 9764 1852
rect 9324 1777 9337 1823
rect 9383 1777 9459 1823
rect 9505 1777 9582 1823
rect 9628 1777 9705 1823
rect 9751 1777 9764 1823
rect 9324 1748 9764 1777
rect 20051 2001 20064 2047
rect 20110 2001 20168 2047
rect 20214 2001 20271 2047
rect 20317 2001 20374 2047
rect 20420 2001 20477 2047
rect 20523 2001 20580 2047
rect 20626 2001 20683 2047
rect 20729 2001 20786 2047
rect 20832 2001 20889 2047
rect 20935 2001 20992 2047
rect 21038 2001 21051 2047
rect 20051 1972 21051 2001
rect 3268 1599 4268 1628
rect 3268 1553 3281 1599
rect 3327 1553 3384 1599
rect 3430 1553 3487 1599
rect 3533 1553 3590 1599
rect 3636 1553 3693 1599
rect 3739 1553 3796 1599
rect 3842 1553 3899 1599
rect 3945 1553 4002 1599
rect 4048 1553 4105 1599
rect 4151 1553 4209 1599
rect 4255 1553 4268 1599
rect 3268 1524 4268 1553
rect 9324 1599 9764 1628
rect 9324 1553 9337 1599
rect 9383 1553 9459 1599
rect 9505 1553 9582 1599
rect 9628 1553 9705 1599
rect 9751 1553 9764 1599
rect 9324 1540 9764 1553
rect 20051 1823 21051 1852
rect 20051 1777 20064 1823
rect 20110 1777 20168 1823
rect 20214 1777 20271 1823
rect 20317 1777 20374 1823
rect 20420 1777 20477 1823
rect 20523 1777 20580 1823
rect 20626 1777 20683 1823
rect 20729 1777 20786 1823
rect 20832 1777 20889 1823
rect 20935 1777 20992 1823
rect 21038 1777 21051 1823
rect 20051 1748 21051 1777
rect 7493 1512 8153 1525
rect 20051 1599 21051 1628
rect 20051 1553 20064 1599
rect 20110 1553 20168 1599
rect 20214 1553 20271 1599
rect 20317 1553 20374 1599
rect 20420 1553 20477 1599
rect 20523 1553 20580 1599
rect 20626 1553 20683 1599
rect 20729 1553 20786 1599
rect 20832 1553 20889 1599
rect 20935 1553 20992 1599
rect 21038 1553 21051 1599
rect 7493 1466 7506 1512
rect 7552 1466 7623 1512
rect 7669 1466 7740 1512
rect 7786 1466 7858 1512
rect 7904 1466 7976 1512
rect 8022 1466 8094 1512
rect 8140 1466 8153 1512
rect 7493 1437 8153 1466
rect 3268 1375 4268 1404
rect 3268 1329 3281 1375
rect 3327 1329 3384 1375
rect 3430 1329 3487 1375
rect 3533 1329 3590 1375
rect 3636 1329 3693 1375
rect 3739 1329 3796 1375
rect 3842 1329 3899 1375
rect 3945 1329 4002 1375
rect 4048 1329 4105 1375
rect 4151 1329 4209 1375
rect 4255 1329 4268 1375
rect 3268 1268 4268 1329
rect 20051 1524 21051 1553
rect 7493 1288 8153 1317
rect 7493 1242 7506 1288
rect 7552 1242 7623 1288
rect 7669 1242 7740 1288
rect 7786 1242 7858 1288
rect 7904 1242 7976 1288
rect 8022 1242 8094 1288
rect 8140 1242 8153 1288
rect 7493 1213 8153 1242
rect 9195 1288 9327 1301
rect 9195 1242 9238 1288
rect 9284 1242 9327 1288
rect 9195 1213 9327 1242
rect 20051 1375 21051 1404
rect 20051 1329 20064 1375
rect 20110 1329 20168 1375
rect 20214 1329 20271 1375
rect 20317 1329 20374 1375
rect 20420 1329 20477 1375
rect 20523 1329 20580 1375
rect 20626 1329 20683 1375
rect 20729 1329 20786 1375
rect 20832 1329 20889 1375
rect 20935 1329 20992 1375
rect 21038 1329 21051 1375
rect 20051 1268 21051 1329
rect 7493 1064 8153 1093
rect 7493 1018 7506 1064
rect 7552 1018 7623 1064
rect 7669 1018 7740 1064
rect 7786 1018 7858 1064
rect 7904 1018 7976 1064
rect 8022 1018 8094 1064
rect 8140 1018 8153 1064
rect 7493 1005 8153 1018
rect 9195 1064 9327 1093
rect 9195 1018 9238 1064
rect 9284 1018 9327 1064
rect 9195 1005 9327 1018
rect 7493 782 8153 795
rect 7493 736 7506 782
rect 7552 736 7623 782
rect 7669 736 7740 782
rect 7786 736 7858 782
rect 7904 736 7976 782
rect 8022 736 8094 782
rect 8140 736 8153 782
rect 7493 707 8153 736
rect 9195 782 9327 795
rect 9195 736 9238 782
rect 9284 736 9327 782
rect 9195 707 9327 736
rect 3268 471 4268 532
rect 3268 425 3281 471
rect 3327 425 3384 471
rect 3430 425 3487 471
rect 3533 425 3590 471
rect 3636 425 3693 471
rect 3739 425 3796 471
rect 3842 425 3899 471
rect 3945 425 4002 471
rect 4048 425 4105 471
rect 4151 425 4209 471
rect 4255 425 4268 471
rect 3268 396 4268 425
rect 7493 558 8153 587
rect 7493 512 7506 558
rect 7552 512 7623 558
rect 7669 512 7740 558
rect 7786 512 7858 558
rect 7904 512 7976 558
rect 8022 512 8094 558
rect 8140 512 8153 558
rect 7493 483 8153 512
rect 9195 558 9327 587
rect 9195 512 9238 558
rect 9284 512 9327 558
rect 9195 499 9327 512
rect 3268 247 4268 276
rect 7493 334 8153 363
rect 7493 288 7506 334
rect 7552 288 7623 334
rect 7669 288 7740 334
rect 7786 288 7858 334
rect 7904 288 7976 334
rect 8022 288 8094 334
rect 8140 288 8153 334
rect 7493 275 8153 288
rect 20051 471 21051 532
rect 20051 425 20064 471
rect 20110 425 20168 471
rect 20214 425 20271 471
rect 20317 425 20374 471
rect 20420 425 20477 471
rect 20523 425 20580 471
rect 20626 425 20683 471
rect 20729 425 20786 471
rect 20832 425 20889 471
rect 20935 425 20992 471
rect 21038 425 21051 471
rect 20051 396 21051 425
rect 3268 201 3281 247
rect 3327 201 3384 247
rect 3430 201 3487 247
rect 3533 201 3590 247
rect 3636 201 3693 247
rect 3739 201 3796 247
rect 3842 201 3899 247
rect 3945 201 4002 247
rect 4048 201 4105 247
rect 4151 201 4209 247
rect 4255 201 4268 247
rect 3268 172 4268 201
rect 9324 247 9764 260
rect 9324 201 9337 247
rect 9383 201 9459 247
rect 9505 201 9582 247
rect 9628 201 9705 247
rect 9751 201 9764 247
rect 9324 172 9764 201
rect 20051 247 21051 276
rect 3268 23 4268 52
rect 3268 -23 3281 23
rect 3327 -23 3384 23
rect 3430 -23 3487 23
rect 3533 -23 3590 23
rect 3636 -23 3693 23
rect 3739 -23 3796 23
rect 3842 -23 3899 23
rect 3945 -23 4002 23
rect 4048 -23 4105 23
rect 4151 -23 4209 23
rect 4255 -23 4268 23
rect 3268 -36 4268 -23
rect 9324 23 9764 52
rect 9324 -23 9337 23
rect 9383 -23 9459 23
rect 9505 -23 9582 23
rect 9628 -23 9705 23
rect 9751 -23 9764 23
rect 9324 -36 9764 -23
rect 20051 201 20064 247
rect 20110 201 20168 247
rect 20214 201 20271 247
rect 20317 201 20374 247
rect 20420 201 20477 247
rect 20523 201 20580 247
rect 20626 201 20683 247
rect 20729 201 20786 247
rect 20832 201 20889 247
rect 20935 201 20992 247
rect 21038 201 21051 247
rect 20051 172 21051 201
rect 20051 23 21051 52
rect 20051 -23 20064 23
rect 20110 -23 20168 23
rect 20214 -23 20271 23
rect 20317 -23 20374 23
rect 20420 -23 20477 23
rect 20523 -23 20580 23
rect 20626 -23 20683 23
rect 20729 -23 20786 23
rect 20832 -23 20889 23
rect 20935 -23 20992 23
rect 21038 -23 21051 23
rect 20051 -36 21051 -23
<< mvpdiff >>
rect 933 14423 2933 14436
rect 933 14377 946 14423
rect 2920 14377 2933 14423
rect 933 14348 2933 14377
rect 933 14199 2933 14228
rect 933 14153 946 14199
rect 2920 14153 2933 14199
rect 933 14124 2933 14153
rect 933 13975 2933 14004
rect 933 13929 946 13975
rect 2920 13929 2933 13975
rect 933 13900 2933 13929
rect 14396 14423 14920 14436
rect 14396 14377 14409 14423
rect 14455 14377 14522 14423
rect 14568 14377 14635 14423
rect 14681 14377 14748 14423
rect 14794 14377 14861 14423
rect 14907 14377 14920 14423
rect 14396 14348 14920 14377
rect 21386 14423 23386 14436
rect 21386 14377 21399 14423
rect 23373 14377 23386 14423
rect 21386 14348 23386 14377
rect 4857 14112 5957 14125
rect 4857 14066 4870 14112
rect 5120 14066 5177 14112
rect 5223 14066 5280 14112
rect 5326 14066 5383 14112
rect 5429 14066 5486 14112
rect 5532 14066 5589 14112
rect 5635 14066 5692 14112
rect 5738 14066 5795 14112
rect 5841 14066 5898 14112
rect 5944 14066 5957 14112
rect 4857 14037 5957 14066
rect 6438 14112 7098 14125
rect 6438 14066 6451 14112
rect 6497 14066 6568 14112
rect 6614 14066 6685 14112
rect 6731 14066 6803 14112
rect 6849 14066 6921 14112
rect 6967 14066 7039 14112
rect 7085 14066 7098 14112
rect 6438 14037 7098 14066
rect 14396 14199 14920 14228
rect 14396 14153 14409 14199
rect 14455 14153 14522 14199
rect 14568 14153 14635 14199
rect 14681 14153 14748 14199
rect 14794 14153 14861 14199
rect 14907 14153 14920 14199
rect 14396 14124 14920 14153
rect 933 13751 2933 13780
rect 933 13705 946 13751
rect 2920 13705 2933 13751
rect 4857 13888 5957 13917
rect 4857 13842 4870 13888
rect 5120 13842 5177 13888
rect 5223 13842 5280 13888
rect 5326 13842 5383 13888
rect 5429 13842 5486 13888
rect 5532 13842 5589 13888
rect 5635 13842 5692 13888
rect 5738 13842 5795 13888
rect 5841 13842 5898 13888
rect 5944 13842 5957 13888
rect 4857 13813 5957 13842
rect 933 13692 2933 13705
rect 18362 14112 19462 14125
rect 18362 14066 18375 14112
rect 18421 14066 18478 14112
rect 18524 14066 18581 14112
rect 18627 14066 18684 14112
rect 18730 14066 18787 14112
rect 18833 14066 18890 14112
rect 18936 14066 18993 14112
rect 19039 14066 19096 14112
rect 19142 14066 19199 14112
rect 19449 14066 19462 14112
rect 18362 14037 19462 14066
rect 6438 13888 7098 13917
rect 6438 13842 6451 13888
rect 6497 13842 6568 13888
rect 6614 13842 6685 13888
rect 6731 13842 6803 13888
rect 6849 13842 6921 13888
rect 6967 13842 7039 13888
rect 7085 13842 7098 13888
rect 6438 13813 7098 13842
rect 8605 13888 8923 13901
rect 8605 13842 8618 13888
rect 8664 13842 8741 13888
rect 8787 13842 8864 13888
rect 8910 13842 8923 13888
rect 8605 13813 8923 13842
rect 14396 13975 14920 14004
rect 14396 13929 14409 13975
rect 14455 13929 14522 13975
rect 14568 13929 14635 13975
rect 14681 13929 14748 13975
rect 14794 13929 14861 13975
rect 14907 13929 14920 13975
rect 14396 13900 14920 13929
rect 18362 13888 19462 13917
rect 18362 13842 18375 13888
rect 18421 13842 18478 13888
rect 18524 13842 18581 13888
rect 18627 13842 18684 13888
rect 18730 13842 18787 13888
rect 18833 13842 18890 13888
rect 18936 13842 18993 13888
rect 19039 13842 19096 13888
rect 19142 13842 19199 13888
rect 19449 13842 19462 13888
rect 18362 13813 19462 13842
rect 4857 13664 5957 13693
rect 4857 13618 4870 13664
rect 5120 13618 5177 13664
rect 5223 13618 5280 13664
rect 5326 13618 5383 13664
rect 5429 13618 5486 13664
rect 5532 13618 5589 13664
rect 5635 13618 5692 13664
rect 5738 13618 5795 13664
rect 5841 13618 5898 13664
rect 5944 13618 5957 13664
rect 4857 13605 5957 13618
rect 6438 13664 7098 13693
rect 6438 13618 6451 13664
rect 6497 13618 6568 13664
rect 6614 13618 6685 13664
rect 6731 13618 6803 13664
rect 6849 13618 6921 13664
rect 6967 13618 7039 13664
rect 7085 13618 7098 13664
rect 6438 13605 7098 13618
rect 8605 13664 8923 13693
rect 8605 13618 8618 13664
rect 8664 13618 8741 13664
rect 8787 13618 8864 13664
rect 8910 13618 8923 13664
rect 8605 13605 8923 13618
rect 14396 13751 14920 13780
rect 14396 13705 14409 13751
rect 14455 13705 14522 13751
rect 14568 13705 14635 13751
rect 14681 13705 14748 13751
rect 14794 13705 14861 13751
rect 14907 13705 14920 13751
rect 14396 13692 14920 13705
rect 21386 14199 23386 14228
rect 21386 14153 21399 14199
rect 23373 14153 23386 14199
rect 21386 14124 23386 14153
rect 21386 13975 23386 14004
rect 21386 13929 21399 13975
rect 23373 13929 23386 13975
rect 21386 13900 23386 13929
rect 21386 13751 23386 13780
rect 18362 13664 19462 13693
rect 18362 13618 18375 13664
rect 18421 13618 18478 13664
rect 18524 13618 18581 13664
rect 18627 13618 18684 13664
rect 18730 13618 18787 13664
rect 18833 13618 18890 13664
rect 18936 13618 18993 13664
rect 19039 13618 19096 13664
rect 19142 13618 19199 13664
rect 19449 13618 19462 13664
rect 21386 13705 21399 13751
rect 23373 13705 23386 13751
rect 21386 13692 23386 13705
rect 18362 13605 19462 13618
rect 4857 13382 5957 13395
rect 933 13295 2933 13308
rect 933 13249 946 13295
rect 2920 13249 2933 13295
rect 4857 13336 4870 13382
rect 5120 13336 5177 13382
rect 5223 13336 5280 13382
rect 5326 13336 5383 13382
rect 5429 13336 5486 13382
rect 5532 13336 5589 13382
rect 5635 13336 5692 13382
rect 5738 13336 5795 13382
rect 5841 13336 5898 13382
rect 5944 13336 5957 13382
rect 4857 13307 5957 13336
rect 6438 13382 7098 13395
rect 6438 13336 6451 13382
rect 6497 13336 6568 13382
rect 6614 13336 6685 13382
rect 6731 13336 6803 13382
rect 6849 13336 6921 13382
rect 6967 13336 7039 13382
rect 7085 13336 7098 13382
rect 6438 13307 7098 13336
rect 8605 13382 8923 13395
rect 8605 13336 8618 13382
rect 8664 13336 8741 13382
rect 8787 13336 8864 13382
rect 8910 13336 8923 13382
rect 8605 13307 8923 13336
rect 18362 13382 19462 13395
rect 933 13220 2933 13249
rect 933 13071 2933 13100
rect 933 13025 946 13071
rect 2920 13025 2933 13071
rect 933 12996 2933 13025
rect 933 12847 2933 12876
rect 933 12801 946 12847
rect 2920 12801 2933 12847
rect 933 12772 2933 12801
rect 4857 13158 5957 13187
rect 4857 13112 4870 13158
rect 5120 13112 5177 13158
rect 5223 13112 5280 13158
rect 5326 13112 5383 13158
rect 5429 13112 5486 13158
rect 5532 13112 5589 13158
rect 5635 13112 5692 13158
rect 5738 13112 5795 13158
rect 5841 13112 5898 13158
rect 5944 13112 5957 13158
rect 4857 13083 5957 13112
rect 6438 13158 7098 13187
rect 6438 13112 6451 13158
rect 6497 13112 6568 13158
rect 6614 13112 6685 13158
rect 6731 13112 6803 13158
rect 6849 13112 6921 13158
rect 6967 13112 7039 13158
rect 7085 13112 7098 13158
rect 6438 13083 7098 13112
rect 18362 13336 18375 13382
rect 18421 13336 18478 13382
rect 18524 13336 18581 13382
rect 18627 13336 18684 13382
rect 18730 13336 18787 13382
rect 18833 13336 18890 13382
rect 18936 13336 18993 13382
rect 19039 13336 19096 13382
rect 19142 13336 19199 13382
rect 19449 13336 19462 13382
rect 14396 13295 14920 13308
rect 18362 13307 19462 13336
rect 14396 13249 14409 13295
rect 14455 13249 14522 13295
rect 14568 13249 14635 13295
rect 14681 13249 14748 13295
rect 14794 13249 14861 13295
rect 14907 13249 14920 13295
rect 14396 13220 14920 13249
rect 8605 13158 8923 13187
rect 8605 13112 8618 13158
rect 8664 13112 8741 13158
rect 8787 13112 8864 13158
rect 8910 13112 8923 13158
rect 8605 13099 8923 13112
rect 21386 13295 23386 13308
rect 14396 13071 14920 13100
rect 14396 13025 14409 13071
rect 14455 13025 14522 13071
rect 14568 13025 14635 13071
rect 14681 13025 14748 13071
rect 14794 13025 14861 13071
rect 14907 13025 14920 13071
rect 14396 12996 14920 13025
rect 18362 13158 19462 13187
rect 18362 13112 18375 13158
rect 18421 13112 18478 13158
rect 18524 13112 18581 13158
rect 18627 13112 18684 13158
rect 18730 13112 18787 13158
rect 18833 13112 18890 13158
rect 18936 13112 18993 13158
rect 19039 13112 19096 13158
rect 19142 13112 19199 13158
rect 19449 13112 19462 13158
rect 18362 13083 19462 13112
rect 21386 13249 21399 13295
rect 23373 13249 23386 13295
rect 21386 13220 23386 13249
rect 4857 12934 5957 12963
rect 4857 12888 4870 12934
rect 5120 12888 5177 12934
rect 5223 12888 5280 12934
rect 5326 12888 5383 12934
rect 5429 12888 5486 12934
rect 5532 12888 5589 12934
rect 5635 12888 5692 12934
rect 5738 12888 5795 12934
rect 5841 12888 5898 12934
rect 5944 12888 5957 12934
rect 4857 12875 5957 12888
rect 6438 12934 7098 12963
rect 6438 12888 6451 12934
rect 6497 12888 6568 12934
rect 6614 12888 6685 12934
rect 6731 12888 6803 12934
rect 6849 12888 6921 12934
rect 6967 12888 7039 12934
rect 7085 12888 7098 12934
rect 6438 12875 7098 12888
rect 18362 12934 19462 12963
rect 18362 12888 18375 12934
rect 18421 12888 18478 12934
rect 18524 12888 18581 12934
rect 18627 12888 18684 12934
rect 18730 12888 18787 12934
rect 18833 12888 18890 12934
rect 18936 12888 18993 12934
rect 19039 12888 19096 12934
rect 19142 12888 19199 12934
rect 19449 12888 19462 12934
rect 14396 12847 14920 12876
rect 18362 12875 19462 12888
rect 14396 12801 14409 12847
rect 14455 12801 14522 12847
rect 14568 12801 14635 12847
rect 14681 12801 14748 12847
rect 14794 12801 14861 12847
rect 14907 12801 14920 12847
rect 933 12623 2933 12652
rect 933 12577 946 12623
rect 2920 12577 2933 12623
rect 933 12548 2933 12577
rect 933 12399 2933 12428
rect 933 12353 946 12399
rect 2920 12353 2933 12399
rect 933 12324 2933 12353
rect 933 12175 2933 12204
rect 933 12129 946 12175
rect 2920 12129 2933 12175
rect 933 12100 2933 12129
rect 14396 12772 14920 12801
rect 21386 13071 23386 13100
rect 21386 13025 21399 13071
rect 23373 13025 23386 13071
rect 21386 12996 23386 13025
rect 21386 12847 23386 12876
rect 21386 12801 21399 12847
rect 23373 12801 23386 12847
rect 21386 12772 23386 12801
rect 14396 12623 14920 12652
rect 14396 12577 14409 12623
rect 14455 12577 14522 12623
rect 14568 12577 14635 12623
rect 14681 12577 14748 12623
rect 14794 12577 14861 12623
rect 14907 12577 14920 12623
rect 14396 12548 14920 12577
rect 21386 12623 23386 12652
rect 21386 12577 21399 12623
rect 23373 12577 23386 12623
rect 21386 12548 23386 12577
rect 4857 12312 5957 12325
rect 4857 12266 4870 12312
rect 5120 12266 5177 12312
rect 5223 12266 5280 12312
rect 5326 12266 5383 12312
rect 5429 12266 5486 12312
rect 5532 12266 5589 12312
rect 5635 12266 5692 12312
rect 5738 12266 5795 12312
rect 5841 12266 5898 12312
rect 5944 12266 5957 12312
rect 4857 12237 5957 12266
rect 6438 12312 7098 12325
rect 6438 12266 6451 12312
rect 6497 12266 6568 12312
rect 6614 12266 6685 12312
rect 6731 12266 6803 12312
rect 6849 12266 6921 12312
rect 6967 12266 7039 12312
rect 7085 12266 7098 12312
rect 6438 12237 7098 12266
rect 14396 12399 14920 12428
rect 14396 12353 14409 12399
rect 14455 12353 14522 12399
rect 14568 12353 14635 12399
rect 14681 12353 14748 12399
rect 14794 12353 14861 12399
rect 14907 12353 14920 12399
rect 14396 12324 14920 12353
rect 933 11951 2933 11980
rect 933 11905 946 11951
rect 2920 11905 2933 11951
rect 4857 12088 5957 12117
rect 4857 12042 4870 12088
rect 5120 12042 5177 12088
rect 5223 12042 5280 12088
rect 5326 12042 5383 12088
rect 5429 12042 5486 12088
rect 5532 12042 5589 12088
rect 5635 12042 5692 12088
rect 5738 12042 5795 12088
rect 5841 12042 5898 12088
rect 5944 12042 5957 12088
rect 4857 12013 5957 12042
rect 933 11892 2933 11905
rect 18362 12312 19462 12325
rect 18362 12266 18375 12312
rect 18421 12266 18478 12312
rect 18524 12266 18581 12312
rect 18627 12266 18684 12312
rect 18730 12266 18787 12312
rect 18833 12266 18890 12312
rect 18936 12266 18993 12312
rect 19039 12266 19096 12312
rect 19142 12266 19199 12312
rect 19449 12266 19462 12312
rect 18362 12237 19462 12266
rect 6438 12088 7098 12117
rect 6438 12042 6451 12088
rect 6497 12042 6568 12088
rect 6614 12042 6685 12088
rect 6731 12042 6803 12088
rect 6849 12042 6921 12088
rect 6967 12042 7039 12088
rect 7085 12042 7098 12088
rect 6438 12013 7098 12042
rect 8605 12088 8923 12101
rect 8605 12042 8618 12088
rect 8664 12042 8741 12088
rect 8787 12042 8864 12088
rect 8910 12042 8923 12088
rect 8605 12013 8923 12042
rect 14396 12175 14920 12204
rect 14396 12129 14409 12175
rect 14455 12129 14522 12175
rect 14568 12129 14635 12175
rect 14681 12129 14748 12175
rect 14794 12129 14861 12175
rect 14907 12129 14920 12175
rect 14396 12100 14920 12129
rect 18362 12088 19462 12117
rect 18362 12042 18375 12088
rect 18421 12042 18478 12088
rect 18524 12042 18581 12088
rect 18627 12042 18684 12088
rect 18730 12042 18787 12088
rect 18833 12042 18890 12088
rect 18936 12042 18993 12088
rect 19039 12042 19096 12088
rect 19142 12042 19199 12088
rect 19449 12042 19462 12088
rect 18362 12013 19462 12042
rect 4857 11864 5957 11893
rect 4857 11818 4870 11864
rect 5120 11818 5177 11864
rect 5223 11818 5280 11864
rect 5326 11818 5383 11864
rect 5429 11818 5486 11864
rect 5532 11818 5589 11864
rect 5635 11818 5692 11864
rect 5738 11818 5795 11864
rect 5841 11818 5898 11864
rect 5944 11818 5957 11864
rect 4857 11805 5957 11818
rect 6438 11864 7098 11893
rect 6438 11818 6451 11864
rect 6497 11818 6568 11864
rect 6614 11818 6685 11864
rect 6731 11818 6803 11864
rect 6849 11818 6921 11864
rect 6967 11818 7039 11864
rect 7085 11818 7098 11864
rect 6438 11805 7098 11818
rect 8605 11864 8923 11893
rect 8605 11818 8618 11864
rect 8664 11818 8741 11864
rect 8787 11818 8864 11864
rect 8910 11818 8923 11864
rect 8605 11805 8923 11818
rect 14396 11951 14920 11980
rect 14396 11905 14409 11951
rect 14455 11905 14522 11951
rect 14568 11905 14635 11951
rect 14681 11905 14748 11951
rect 14794 11905 14861 11951
rect 14907 11905 14920 11951
rect 14396 11892 14920 11905
rect 21386 12399 23386 12428
rect 21386 12353 21399 12399
rect 23373 12353 23386 12399
rect 21386 12324 23386 12353
rect 21386 12175 23386 12204
rect 21386 12129 21399 12175
rect 23373 12129 23386 12175
rect 21386 12100 23386 12129
rect 21386 11951 23386 11980
rect 18362 11864 19462 11893
rect 18362 11818 18375 11864
rect 18421 11818 18478 11864
rect 18524 11818 18581 11864
rect 18627 11818 18684 11864
rect 18730 11818 18787 11864
rect 18833 11818 18890 11864
rect 18936 11818 18993 11864
rect 19039 11818 19096 11864
rect 19142 11818 19199 11864
rect 19449 11818 19462 11864
rect 21386 11905 21399 11951
rect 23373 11905 23386 11951
rect 21386 11892 23386 11905
rect 18362 11805 19462 11818
rect 4857 11582 5957 11595
rect 933 11495 2933 11508
rect 933 11449 946 11495
rect 2920 11449 2933 11495
rect 4857 11536 4870 11582
rect 5120 11536 5177 11582
rect 5223 11536 5280 11582
rect 5326 11536 5383 11582
rect 5429 11536 5486 11582
rect 5532 11536 5589 11582
rect 5635 11536 5692 11582
rect 5738 11536 5795 11582
rect 5841 11536 5898 11582
rect 5944 11536 5957 11582
rect 4857 11507 5957 11536
rect 6438 11582 7098 11595
rect 6438 11536 6451 11582
rect 6497 11536 6568 11582
rect 6614 11536 6685 11582
rect 6731 11536 6803 11582
rect 6849 11536 6921 11582
rect 6967 11536 7039 11582
rect 7085 11536 7098 11582
rect 6438 11507 7098 11536
rect 8605 11582 8923 11595
rect 8605 11536 8618 11582
rect 8664 11536 8741 11582
rect 8787 11536 8864 11582
rect 8910 11536 8923 11582
rect 8605 11507 8923 11536
rect 18362 11582 19462 11595
rect 933 11420 2933 11449
rect 933 11271 2933 11300
rect 933 11225 946 11271
rect 2920 11225 2933 11271
rect 933 11196 2933 11225
rect 933 11047 2933 11076
rect 933 11001 946 11047
rect 2920 11001 2933 11047
rect 933 10972 2933 11001
rect 4857 11358 5957 11387
rect 4857 11312 4870 11358
rect 5120 11312 5177 11358
rect 5223 11312 5280 11358
rect 5326 11312 5383 11358
rect 5429 11312 5486 11358
rect 5532 11312 5589 11358
rect 5635 11312 5692 11358
rect 5738 11312 5795 11358
rect 5841 11312 5898 11358
rect 5944 11312 5957 11358
rect 4857 11283 5957 11312
rect 6438 11358 7098 11387
rect 6438 11312 6451 11358
rect 6497 11312 6568 11358
rect 6614 11312 6685 11358
rect 6731 11312 6803 11358
rect 6849 11312 6921 11358
rect 6967 11312 7039 11358
rect 7085 11312 7098 11358
rect 6438 11283 7098 11312
rect 18362 11536 18375 11582
rect 18421 11536 18478 11582
rect 18524 11536 18581 11582
rect 18627 11536 18684 11582
rect 18730 11536 18787 11582
rect 18833 11536 18890 11582
rect 18936 11536 18993 11582
rect 19039 11536 19096 11582
rect 19142 11536 19199 11582
rect 19449 11536 19462 11582
rect 14396 11495 14920 11508
rect 18362 11507 19462 11536
rect 14396 11449 14409 11495
rect 14455 11449 14522 11495
rect 14568 11449 14635 11495
rect 14681 11449 14748 11495
rect 14794 11449 14861 11495
rect 14907 11449 14920 11495
rect 14396 11420 14920 11449
rect 8605 11358 8923 11387
rect 8605 11312 8618 11358
rect 8664 11312 8741 11358
rect 8787 11312 8864 11358
rect 8910 11312 8923 11358
rect 8605 11299 8923 11312
rect 21386 11495 23386 11508
rect 14396 11271 14920 11300
rect 14396 11225 14409 11271
rect 14455 11225 14522 11271
rect 14568 11225 14635 11271
rect 14681 11225 14748 11271
rect 14794 11225 14861 11271
rect 14907 11225 14920 11271
rect 14396 11196 14920 11225
rect 18362 11358 19462 11387
rect 18362 11312 18375 11358
rect 18421 11312 18478 11358
rect 18524 11312 18581 11358
rect 18627 11312 18684 11358
rect 18730 11312 18787 11358
rect 18833 11312 18890 11358
rect 18936 11312 18993 11358
rect 19039 11312 19096 11358
rect 19142 11312 19199 11358
rect 19449 11312 19462 11358
rect 18362 11283 19462 11312
rect 21386 11449 21399 11495
rect 23373 11449 23386 11495
rect 21386 11420 23386 11449
rect 4857 11134 5957 11163
rect 4857 11088 4870 11134
rect 5120 11088 5177 11134
rect 5223 11088 5280 11134
rect 5326 11088 5383 11134
rect 5429 11088 5486 11134
rect 5532 11088 5589 11134
rect 5635 11088 5692 11134
rect 5738 11088 5795 11134
rect 5841 11088 5898 11134
rect 5944 11088 5957 11134
rect 4857 11075 5957 11088
rect 6438 11134 7098 11163
rect 6438 11088 6451 11134
rect 6497 11088 6568 11134
rect 6614 11088 6685 11134
rect 6731 11088 6803 11134
rect 6849 11088 6921 11134
rect 6967 11088 7039 11134
rect 7085 11088 7098 11134
rect 6438 11075 7098 11088
rect 18362 11134 19462 11163
rect 18362 11088 18375 11134
rect 18421 11088 18478 11134
rect 18524 11088 18581 11134
rect 18627 11088 18684 11134
rect 18730 11088 18787 11134
rect 18833 11088 18890 11134
rect 18936 11088 18993 11134
rect 19039 11088 19096 11134
rect 19142 11088 19199 11134
rect 19449 11088 19462 11134
rect 14396 11047 14920 11076
rect 18362 11075 19462 11088
rect 14396 11001 14409 11047
rect 14455 11001 14522 11047
rect 14568 11001 14635 11047
rect 14681 11001 14748 11047
rect 14794 11001 14861 11047
rect 14907 11001 14920 11047
rect 933 10823 2933 10852
rect 933 10777 946 10823
rect 2920 10777 2933 10823
rect 933 10748 2933 10777
rect 933 10599 2933 10628
rect 933 10553 946 10599
rect 2920 10553 2933 10599
rect 933 10524 2933 10553
rect 933 10375 2933 10404
rect 933 10329 946 10375
rect 2920 10329 2933 10375
rect 933 10300 2933 10329
rect 14396 10972 14920 11001
rect 21386 11271 23386 11300
rect 21386 11225 21399 11271
rect 23373 11225 23386 11271
rect 21386 11196 23386 11225
rect 21386 11047 23386 11076
rect 21386 11001 21399 11047
rect 23373 11001 23386 11047
rect 21386 10972 23386 11001
rect 14396 10823 14920 10852
rect 14396 10777 14409 10823
rect 14455 10777 14522 10823
rect 14568 10777 14635 10823
rect 14681 10777 14748 10823
rect 14794 10777 14861 10823
rect 14907 10777 14920 10823
rect 14396 10748 14920 10777
rect 21386 10823 23386 10852
rect 21386 10777 21399 10823
rect 23373 10777 23386 10823
rect 21386 10748 23386 10777
rect 4857 10512 5957 10525
rect 4857 10466 4870 10512
rect 5120 10466 5177 10512
rect 5223 10466 5280 10512
rect 5326 10466 5383 10512
rect 5429 10466 5486 10512
rect 5532 10466 5589 10512
rect 5635 10466 5692 10512
rect 5738 10466 5795 10512
rect 5841 10466 5898 10512
rect 5944 10466 5957 10512
rect 4857 10437 5957 10466
rect 6438 10512 7098 10525
rect 6438 10466 6451 10512
rect 6497 10466 6568 10512
rect 6614 10466 6685 10512
rect 6731 10466 6803 10512
rect 6849 10466 6921 10512
rect 6967 10466 7039 10512
rect 7085 10466 7098 10512
rect 6438 10437 7098 10466
rect 14396 10599 14920 10628
rect 14396 10553 14409 10599
rect 14455 10553 14522 10599
rect 14568 10553 14635 10599
rect 14681 10553 14748 10599
rect 14794 10553 14861 10599
rect 14907 10553 14920 10599
rect 14396 10524 14920 10553
rect 933 10151 2933 10180
rect 933 10105 946 10151
rect 2920 10105 2933 10151
rect 4857 10288 5957 10317
rect 4857 10242 4870 10288
rect 5120 10242 5177 10288
rect 5223 10242 5280 10288
rect 5326 10242 5383 10288
rect 5429 10242 5486 10288
rect 5532 10242 5589 10288
rect 5635 10242 5692 10288
rect 5738 10242 5795 10288
rect 5841 10242 5898 10288
rect 5944 10242 5957 10288
rect 4857 10213 5957 10242
rect 933 10092 2933 10105
rect 18362 10512 19462 10525
rect 18362 10466 18375 10512
rect 18421 10466 18478 10512
rect 18524 10466 18581 10512
rect 18627 10466 18684 10512
rect 18730 10466 18787 10512
rect 18833 10466 18890 10512
rect 18936 10466 18993 10512
rect 19039 10466 19096 10512
rect 19142 10466 19199 10512
rect 19449 10466 19462 10512
rect 18362 10437 19462 10466
rect 6438 10288 7098 10317
rect 6438 10242 6451 10288
rect 6497 10242 6568 10288
rect 6614 10242 6685 10288
rect 6731 10242 6803 10288
rect 6849 10242 6921 10288
rect 6967 10242 7039 10288
rect 7085 10242 7098 10288
rect 6438 10213 7098 10242
rect 8605 10288 8923 10301
rect 8605 10242 8618 10288
rect 8664 10242 8741 10288
rect 8787 10242 8864 10288
rect 8910 10242 8923 10288
rect 8605 10213 8923 10242
rect 14396 10375 14920 10404
rect 14396 10329 14409 10375
rect 14455 10329 14522 10375
rect 14568 10329 14635 10375
rect 14681 10329 14748 10375
rect 14794 10329 14861 10375
rect 14907 10329 14920 10375
rect 14396 10300 14920 10329
rect 18362 10288 19462 10317
rect 18362 10242 18375 10288
rect 18421 10242 18478 10288
rect 18524 10242 18581 10288
rect 18627 10242 18684 10288
rect 18730 10242 18787 10288
rect 18833 10242 18890 10288
rect 18936 10242 18993 10288
rect 19039 10242 19096 10288
rect 19142 10242 19199 10288
rect 19449 10242 19462 10288
rect 18362 10213 19462 10242
rect 4857 10064 5957 10093
rect 4857 10018 4870 10064
rect 5120 10018 5177 10064
rect 5223 10018 5280 10064
rect 5326 10018 5383 10064
rect 5429 10018 5486 10064
rect 5532 10018 5589 10064
rect 5635 10018 5692 10064
rect 5738 10018 5795 10064
rect 5841 10018 5898 10064
rect 5944 10018 5957 10064
rect 4857 10005 5957 10018
rect 6438 10064 7098 10093
rect 6438 10018 6451 10064
rect 6497 10018 6568 10064
rect 6614 10018 6685 10064
rect 6731 10018 6803 10064
rect 6849 10018 6921 10064
rect 6967 10018 7039 10064
rect 7085 10018 7098 10064
rect 6438 10005 7098 10018
rect 8605 10064 8923 10093
rect 8605 10018 8618 10064
rect 8664 10018 8741 10064
rect 8787 10018 8864 10064
rect 8910 10018 8923 10064
rect 8605 10005 8923 10018
rect 14396 10151 14920 10180
rect 14396 10105 14409 10151
rect 14455 10105 14522 10151
rect 14568 10105 14635 10151
rect 14681 10105 14748 10151
rect 14794 10105 14861 10151
rect 14907 10105 14920 10151
rect 14396 10092 14920 10105
rect 21386 10599 23386 10628
rect 21386 10553 21399 10599
rect 23373 10553 23386 10599
rect 21386 10524 23386 10553
rect 21386 10375 23386 10404
rect 21386 10329 21399 10375
rect 23373 10329 23386 10375
rect 21386 10300 23386 10329
rect 21386 10151 23386 10180
rect 18362 10064 19462 10093
rect 18362 10018 18375 10064
rect 18421 10018 18478 10064
rect 18524 10018 18581 10064
rect 18627 10018 18684 10064
rect 18730 10018 18787 10064
rect 18833 10018 18890 10064
rect 18936 10018 18993 10064
rect 19039 10018 19096 10064
rect 19142 10018 19199 10064
rect 19449 10018 19462 10064
rect 21386 10105 21399 10151
rect 23373 10105 23386 10151
rect 21386 10092 23386 10105
rect 18362 10005 19462 10018
rect 4857 9782 5957 9795
rect 933 9695 2933 9708
rect 933 9649 946 9695
rect 2920 9649 2933 9695
rect 4857 9736 4870 9782
rect 5120 9736 5177 9782
rect 5223 9736 5280 9782
rect 5326 9736 5383 9782
rect 5429 9736 5486 9782
rect 5532 9736 5589 9782
rect 5635 9736 5692 9782
rect 5738 9736 5795 9782
rect 5841 9736 5898 9782
rect 5944 9736 5957 9782
rect 4857 9707 5957 9736
rect 6438 9782 7098 9795
rect 6438 9736 6451 9782
rect 6497 9736 6568 9782
rect 6614 9736 6685 9782
rect 6731 9736 6803 9782
rect 6849 9736 6921 9782
rect 6967 9736 7039 9782
rect 7085 9736 7098 9782
rect 6438 9707 7098 9736
rect 8605 9782 8923 9795
rect 8605 9736 8618 9782
rect 8664 9736 8741 9782
rect 8787 9736 8864 9782
rect 8910 9736 8923 9782
rect 8605 9707 8923 9736
rect 18362 9782 19462 9795
rect 933 9620 2933 9649
rect 933 9471 2933 9500
rect 933 9425 946 9471
rect 2920 9425 2933 9471
rect 933 9396 2933 9425
rect 933 9247 2933 9276
rect 933 9201 946 9247
rect 2920 9201 2933 9247
rect 933 9172 2933 9201
rect 4857 9558 5957 9587
rect 4857 9512 4870 9558
rect 5120 9512 5177 9558
rect 5223 9512 5280 9558
rect 5326 9512 5383 9558
rect 5429 9512 5486 9558
rect 5532 9512 5589 9558
rect 5635 9512 5692 9558
rect 5738 9512 5795 9558
rect 5841 9512 5898 9558
rect 5944 9512 5957 9558
rect 4857 9483 5957 9512
rect 6438 9558 7098 9587
rect 6438 9512 6451 9558
rect 6497 9512 6568 9558
rect 6614 9512 6685 9558
rect 6731 9512 6803 9558
rect 6849 9512 6921 9558
rect 6967 9512 7039 9558
rect 7085 9512 7098 9558
rect 6438 9483 7098 9512
rect 18362 9736 18375 9782
rect 18421 9736 18478 9782
rect 18524 9736 18581 9782
rect 18627 9736 18684 9782
rect 18730 9736 18787 9782
rect 18833 9736 18890 9782
rect 18936 9736 18993 9782
rect 19039 9736 19096 9782
rect 19142 9736 19199 9782
rect 19449 9736 19462 9782
rect 14396 9695 14920 9708
rect 18362 9707 19462 9736
rect 14396 9649 14409 9695
rect 14455 9649 14522 9695
rect 14568 9649 14635 9695
rect 14681 9649 14748 9695
rect 14794 9649 14861 9695
rect 14907 9649 14920 9695
rect 14396 9620 14920 9649
rect 8605 9558 8923 9587
rect 8605 9512 8618 9558
rect 8664 9512 8741 9558
rect 8787 9512 8864 9558
rect 8910 9512 8923 9558
rect 8605 9499 8923 9512
rect 21386 9695 23386 9708
rect 14396 9471 14920 9500
rect 14396 9425 14409 9471
rect 14455 9425 14522 9471
rect 14568 9425 14635 9471
rect 14681 9425 14748 9471
rect 14794 9425 14861 9471
rect 14907 9425 14920 9471
rect 14396 9396 14920 9425
rect 18362 9558 19462 9587
rect 18362 9512 18375 9558
rect 18421 9512 18478 9558
rect 18524 9512 18581 9558
rect 18627 9512 18684 9558
rect 18730 9512 18787 9558
rect 18833 9512 18890 9558
rect 18936 9512 18993 9558
rect 19039 9512 19096 9558
rect 19142 9512 19199 9558
rect 19449 9512 19462 9558
rect 18362 9483 19462 9512
rect 21386 9649 21399 9695
rect 23373 9649 23386 9695
rect 21386 9620 23386 9649
rect 4857 9334 5957 9363
rect 4857 9288 4870 9334
rect 5120 9288 5177 9334
rect 5223 9288 5280 9334
rect 5326 9288 5383 9334
rect 5429 9288 5486 9334
rect 5532 9288 5589 9334
rect 5635 9288 5692 9334
rect 5738 9288 5795 9334
rect 5841 9288 5898 9334
rect 5944 9288 5957 9334
rect 4857 9275 5957 9288
rect 6438 9334 7098 9363
rect 6438 9288 6451 9334
rect 6497 9288 6568 9334
rect 6614 9288 6685 9334
rect 6731 9288 6803 9334
rect 6849 9288 6921 9334
rect 6967 9288 7039 9334
rect 7085 9288 7098 9334
rect 6438 9275 7098 9288
rect 18362 9334 19462 9363
rect 18362 9288 18375 9334
rect 18421 9288 18478 9334
rect 18524 9288 18581 9334
rect 18627 9288 18684 9334
rect 18730 9288 18787 9334
rect 18833 9288 18890 9334
rect 18936 9288 18993 9334
rect 19039 9288 19096 9334
rect 19142 9288 19199 9334
rect 19449 9288 19462 9334
rect 14396 9247 14920 9276
rect 18362 9275 19462 9288
rect 14396 9201 14409 9247
rect 14455 9201 14522 9247
rect 14568 9201 14635 9247
rect 14681 9201 14748 9247
rect 14794 9201 14861 9247
rect 14907 9201 14920 9247
rect 933 9023 2933 9052
rect 933 8977 946 9023
rect 2920 8977 2933 9023
rect 933 8948 2933 8977
rect 933 8799 2933 8828
rect 933 8753 946 8799
rect 2920 8753 2933 8799
rect 933 8724 2933 8753
rect 933 8575 2933 8604
rect 933 8529 946 8575
rect 2920 8529 2933 8575
rect 933 8500 2933 8529
rect 14396 9172 14920 9201
rect 21386 9471 23386 9500
rect 21386 9425 21399 9471
rect 23373 9425 23386 9471
rect 21386 9396 23386 9425
rect 21386 9247 23386 9276
rect 21386 9201 21399 9247
rect 23373 9201 23386 9247
rect 21386 9172 23386 9201
rect 14396 9023 14920 9052
rect 14396 8977 14409 9023
rect 14455 8977 14522 9023
rect 14568 8977 14635 9023
rect 14681 8977 14748 9023
rect 14794 8977 14861 9023
rect 14907 8977 14920 9023
rect 14396 8948 14920 8977
rect 21386 9023 23386 9052
rect 21386 8977 21399 9023
rect 23373 8977 23386 9023
rect 21386 8948 23386 8977
rect 4857 8712 5957 8725
rect 4857 8666 4870 8712
rect 5120 8666 5177 8712
rect 5223 8666 5280 8712
rect 5326 8666 5383 8712
rect 5429 8666 5486 8712
rect 5532 8666 5589 8712
rect 5635 8666 5692 8712
rect 5738 8666 5795 8712
rect 5841 8666 5898 8712
rect 5944 8666 5957 8712
rect 4857 8637 5957 8666
rect 6438 8712 7098 8725
rect 6438 8666 6451 8712
rect 6497 8666 6568 8712
rect 6614 8666 6685 8712
rect 6731 8666 6803 8712
rect 6849 8666 6921 8712
rect 6967 8666 7039 8712
rect 7085 8666 7098 8712
rect 6438 8637 7098 8666
rect 14396 8799 14920 8828
rect 14396 8753 14409 8799
rect 14455 8753 14522 8799
rect 14568 8753 14635 8799
rect 14681 8753 14748 8799
rect 14794 8753 14861 8799
rect 14907 8753 14920 8799
rect 14396 8724 14920 8753
rect 933 8351 2933 8380
rect 933 8305 946 8351
rect 2920 8305 2933 8351
rect 4857 8488 5957 8517
rect 4857 8442 4870 8488
rect 5120 8442 5177 8488
rect 5223 8442 5280 8488
rect 5326 8442 5383 8488
rect 5429 8442 5486 8488
rect 5532 8442 5589 8488
rect 5635 8442 5692 8488
rect 5738 8442 5795 8488
rect 5841 8442 5898 8488
rect 5944 8442 5957 8488
rect 4857 8413 5957 8442
rect 933 8292 2933 8305
rect 18362 8712 19462 8725
rect 18362 8666 18375 8712
rect 18421 8666 18478 8712
rect 18524 8666 18581 8712
rect 18627 8666 18684 8712
rect 18730 8666 18787 8712
rect 18833 8666 18890 8712
rect 18936 8666 18993 8712
rect 19039 8666 19096 8712
rect 19142 8666 19199 8712
rect 19449 8666 19462 8712
rect 18362 8637 19462 8666
rect 6438 8488 7098 8517
rect 6438 8442 6451 8488
rect 6497 8442 6568 8488
rect 6614 8442 6685 8488
rect 6731 8442 6803 8488
rect 6849 8442 6921 8488
rect 6967 8442 7039 8488
rect 7085 8442 7098 8488
rect 6438 8413 7098 8442
rect 8605 8488 8923 8501
rect 8605 8442 8618 8488
rect 8664 8442 8741 8488
rect 8787 8442 8864 8488
rect 8910 8442 8923 8488
rect 8605 8413 8923 8442
rect 14396 8575 14920 8604
rect 14396 8529 14409 8575
rect 14455 8529 14522 8575
rect 14568 8529 14635 8575
rect 14681 8529 14748 8575
rect 14794 8529 14861 8575
rect 14907 8529 14920 8575
rect 14396 8500 14920 8529
rect 18362 8488 19462 8517
rect 18362 8442 18375 8488
rect 18421 8442 18478 8488
rect 18524 8442 18581 8488
rect 18627 8442 18684 8488
rect 18730 8442 18787 8488
rect 18833 8442 18890 8488
rect 18936 8442 18993 8488
rect 19039 8442 19096 8488
rect 19142 8442 19199 8488
rect 19449 8442 19462 8488
rect 18362 8413 19462 8442
rect 4857 8264 5957 8293
rect 4857 8218 4870 8264
rect 5120 8218 5177 8264
rect 5223 8218 5280 8264
rect 5326 8218 5383 8264
rect 5429 8218 5486 8264
rect 5532 8218 5589 8264
rect 5635 8218 5692 8264
rect 5738 8218 5795 8264
rect 5841 8218 5898 8264
rect 5944 8218 5957 8264
rect 4857 8205 5957 8218
rect 6438 8264 7098 8293
rect 6438 8218 6451 8264
rect 6497 8218 6568 8264
rect 6614 8218 6685 8264
rect 6731 8218 6803 8264
rect 6849 8218 6921 8264
rect 6967 8218 7039 8264
rect 7085 8218 7098 8264
rect 6438 8205 7098 8218
rect 8605 8264 8923 8293
rect 8605 8218 8618 8264
rect 8664 8218 8741 8264
rect 8787 8218 8864 8264
rect 8910 8218 8923 8264
rect 8605 8205 8923 8218
rect 14396 8351 14920 8380
rect 14396 8305 14409 8351
rect 14455 8305 14522 8351
rect 14568 8305 14635 8351
rect 14681 8305 14748 8351
rect 14794 8305 14861 8351
rect 14907 8305 14920 8351
rect 14396 8292 14920 8305
rect 21386 8799 23386 8828
rect 21386 8753 21399 8799
rect 23373 8753 23386 8799
rect 21386 8724 23386 8753
rect 21386 8575 23386 8604
rect 21386 8529 21399 8575
rect 23373 8529 23386 8575
rect 21386 8500 23386 8529
rect 21386 8351 23386 8380
rect 18362 8264 19462 8293
rect 18362 8218 18375 8264
rect 18421 8218 18478 8264
rect 18524 8218 18581 8264
rect 18627 8218 18684 8264
rect 18730 8218 18787 8264
rect 18833 8218 18890 8264
rect 18936 8218 18993 8264
rect 19039 8218 19096 8264
rect 19142 8218 19199 8264
rect 19449 8218 19462 8264
rect 21386 8305 21399 8351
rect 23373 8305 23386 8351
rect 21386 8292 23386 8305
rect 18362 8205 19462 8218
rect 4857 7982 5957 7995
rect 933 7895 2933 7908
rect 933 7849 946 7895
rect 2920 7849 2933 7895
rect 4857 7936 4870 7982
rect 5120 7936 5177 7982
rect 5223 7936 5280 7982
rect 5326 7936 5383 7982
rect 5429 7936 5486 7982
rect 5532 7936 5589 7982
rect 5635 7936 5692 7982
rect 5738 7936 5795 7982
rect 5841 7936 5898 7982
rect 5944 7936 5957 7982
rect 4857 7907 5957 7936
rect 6438 7982 7098 7995
rect 6438 7936 6451 7982
rect 6497 7936 6568 7982
rect 6614 7936 6685 7982
rect 6731 7936 6803 7982
rect 6849 7936 6921 7982
rect 6967 7936 7039 7982
rect 7085 7936 7098 7982
rect 6438 7907 7098 7936
rect 8605 7982 8923 7995
rect 8605 7936 8618 7982
rect 8664 7936 8741 7982
rect 8787 7936 8864 7982
rect 8910 7936 8923 7982
rect 8605 7907 8923 7936
rect 18362 7982 19462 7995
rect 933 7820 2933 7849
rect 933 7671 2933 7700
rect 933 7625 946 7671
rect 2920 7625 2933 7671
rect 933 7596 2933 7625
rect 933 7447 2933 7476
rect 933 7401 946 7447
rect 2920 7401 2933 7447
rect 933 7372 2933 7401
rect 4857 7758 5957 7787
rect 4857 7712 4870 7758
rect 5120 7712 5177 7758
rect 5223 7712 5280 7758
rect 5326 7712 5383 7758
rect 5429 7712 5486 7758
rect 5532 7712 5589 7758
rect 5635 7712 5692 7758
rect 5738 7712 5795 7758
rect 5841 7712 5898 7758
rect 5944 7712 5957 7758
rect 4857 7683 5957 7712
rect 6438 7758 7098 7787
rect 6438 7712 6451 7758
rect 6497 7712 6568 7758
rect 6614 7712 6685 7758
rect 6731 7712 6803 7758
rect 6849 7712 6921 7758
rect 6967 7712 7039 7758
rect 7085 7712 7098 7758
rect 6438 7683 7098 7712
rect 18362 7936 18375 7982
rect 18421 7936 18478 7982
rect 18524 7936 18581 7982
rect 18627 7936 18684 7982
rect 18730 7936 18787 7982
rect 18833 7936 18890 7982
rect 18936 7936 18993 7982
rect 19039 7936 19096 7982
rect 19142 7936 19199 7982
rect 19449 7936 19462 7982
rect 14396 7895 14920 7908
rect 18362 7907 19462 7936
rect 14396 7849 14409 7895
rect 14455 7849 14522 7895
rect 14568 7849 14635 7895
rect 14681 7849 14748 7895
rect 14794 7849 14861 7895
rect 14907 7849 14920 7895
rect 14396 7820 14920 7849
rect 8605 7758 8923 7787
rect 8605 7712 8618 7758
rect 8664 7712 8741 7758
rect 8787 7712 8864 7758
rect 8910 7712 8923 7758
rect 8605 7699 8923 7712
rect 21386 7895 23386 7908
rect 14396 7671 14920 7700
rect 14396 7625 14409 7671
rect 14455 7625 14522 7671
rect 14568 7625 14635 7671
rect 14681 7625 14748 7671
rect 14794 7625 14861 7671
rect 14907 7625 14920 7671
rect 14396 7596 14920 7625
rect 18362 7758 19462 7787
rect 18362 7712 18375 7758
rect 18421 7712 18478 7758
rect 18524 7712 18581 7758
rect 18627 7712 18684 7758
rect 18730 7712 18787 7758
rect 18833 7712 18890 7758
rect 18936 7712 18993 7758
rect 19039 7712 19096 7758
rect 19142 7712 19199 7758
rect 19449 7712 19462 7758
rect 18362 7683 19462 7712
rect 21386 7849 21399 7895
rect 23373 7849 23386 7895
rect 21386 7820 23386 7849
rect 4857 7534 5957 7563
rect 4857 7488 4870 7534
rect 5120 7488 5177 7534
rect 5223 7488 5280 7534
rect 5326 7488 5383 7534
rect 5429 7488 5486 7534
rect 5532 7488 5589 7534
rect 5635 7488 5692 7534
rect 5738 7488 5795 7534
rect 5841 7488 5898 7534
rect 5944 7488 5957 7534
rect 4857 7475 5957 7488
rect 6438 7534 7098 7563
rect 6438 7488 6451 7534
rect 6497 7488 6568 7534
rect 6614 7488 6685 7534
rect 6731 7488 6803 7534
rect 6849 7488 6921 7534
rect 6967 7488 7039 7534
rect 7085 7488 7098 7534
rect 6438 7475 7098 7488
rect 18362 7534 19462 7563
rect 18362 7488 18375 7534
rect 18421 7488 18478 7534
rect 18524 7488 18581 7534
rect 18627 7488 18684 7534
rect 18730 7488 18787 7534
rect 18833 7488 18890 7534
rect 18936 7488 18993 7534
rect 19039 7488 19096 7534
rect 19142 7488 19199 7534
rect 19449 7488 19462 7534
rect 14396 7447 14920 7476
rect 18362 7475 19462 7488
rect 14396 7401 14409 7447
rect 14455 7401 14522 7447
rect 14568 7401 14635 7447
rect 14681 7401 14748 7447
rect 14794 7401 14861 7447
rect 14907 7401 14920 7447
rect 933 7223 2933 7252
rect 933 7177 946 7223
rect 2920 7177 2933 7223
rect 933 7148 2933 7177
rect 933 6999 2933 7028
rect 933 6953 946 6999
rect 2920 6953 2933 6999
rect 933 6924 2933 6953
rect 933 6775 2933 6804
rect 933 6729 946 6775
rect 2920 6729 2933 6775
rect 933 6700 2933 6729
rect 14396 7372 14920 7401
rect 21386 7671 23386 7700
rect 21386 7625 21399 7671
rect 23373 7625 23386 7671
rect 21386 7596 23386 7625
rect 21386 7447 23386 7476
rect 21386 7401 21399 7447
rect 23373 7401 23386 7447
rect 21386 7372 23386 7401
rect 14396 7223 14920 7252
rect 14396 7177 14409 7223
rect 14455 7177 14522 7223
rect 14568 7177 14635 7223
rect 14681 7177 14748 7223
rect 14794 7177 14861 7223
rect 14907 7177 14920 7223
rect 14396 7148 14920 7177
rect 21386 7223 23386 7252
rect 21386 7177 21399 7223
rect 23373 7177 23386 7223
rect 21386 7148 23386 7177
rect 4857 6912 5957 6925
rect 4857 6866 4870 6912
rect 5120 6866 5177 6912
rect 5223 6866 5280 6912
rect 5326 6866 5383 6912
rect 5429 6866 5486 6912
rect 5532 6866 5589 6912
rect 5635 6866 5692 6912
rect 5738 6866 5795 6912
rect 5841 6866 5898 6912
rect 5944 6866 5957 6912
rect 4857 6837 5957 6866
rect 6438 6912 7098 6925
rect 6438 6866 6451 6912
rect 6497 6866 6568 6912
rect 6614 6866 6685 6912
rect 6731 6866 6803 6912
rect 6849 6866 6921 6912
rect 6967 6866 7039 6912
rect 7085 6866 7098 6912
rect 6438 6837 7098 6866
rect 14396 6999 14920 7028
rect 14396 6953 14409 6999
rect 14455 6953 14522 6999
rect 14568 6953 14635 6999
rect 14681 6953 14748 6999
rect 14794 6953 14861 6999
rect 14907 6953 14920 6999
rect 14396 6924 14920 6953
rect 933 6551 2933 6580
rect 933 6505 946 6551
rect 2920 6505 2933 6551
rect 4857 6688 5957 6717
rect 4857 6642 4870 6688
rect 5120 6642 5177 6688
rect 5223 6642 5280 6688
rect 5326 6642 5383 6688
rect 5429 6642 5486 6688
rect 5532 6642 5589 6688
rect 5635 6642 5692 6688
rect 5738 6642 5795 6688
rect 5841 6642 5898 6688
rect 5944 6642 5957 6688
rect 4857 6613 5957 6642
rect 933 6492 2933 6505
rect 18362 6912 19462 6925
rect 18362 6866 18375 6912
rect 18421 6866 18478 6912
rect 18524 6866 18581 6912
rect 18627 6866 18684 6912
rect 18730 6866 18787 6912
rect 18833 6866 18890 6912
rect 18936 6866 18993 6912
rect 19039 6866 19096 6912
rect 19142 6866 19199 6912
rect 19449 6866 19462 6912
rect 18362 6837 19462 6866
rect 6438 6688 7098 6717
rect 6438 6642 6451 6688
rect 6497 6642 6568 6688
rect 6614 6642 6685 6688
rect 6731 6642 6803 6688
rect 6849 6642 6921 6688
rect 6967 6642 7039 6688
rect 7085 6642 7098 6688
rect 6438 6613 7098 6642
rect 8605 6688 8923 6701
rect 8605 6642 8618 6688
rect 8664 6642 8741 6688
rect 8787 6642 8864 6688
rect 8910 6642 8923 6688
rect 8605 6613 8923 6642
rect 14396 6775 14920 6804
rect 14396 6729 14409 6775
rect 14455 6729 14522 6775
rect 14568 6729 14635 6775
rect 14681 6729 14748 6775
rect 14794 6729 14861 6775
rect 14907 6729 14920 6775
rect 14396 6700 14920 6729
rect 18362 6688 19462 6717
rect 18362 6642 18375 6688
rect 18421 6642 18478 6688
rect 18524 6642 18581 6688
rect 18627 6642 18684 6688
rect 18730 6642 18787 6688
rect 18833 6642 18890 6688
rect 18936 6642 18993 6688
rect 19039 6642 19096 6688
rect 19142 6642 19199 6688
rect 19449 6642 19462 6688
rect 18362 6613 19462 6642
rect 4857 6464 5957 6493
rect 4857 6418 4870 6464
rect 5120 6418 5177 6464
rect 5223 6418 5280 6464
rect 5326 6418 5383 6464
rect 5429 6418 5486 6464
rect 5532 6418 5589 6464
rect 5635 6418 5692 6464
rect 5738 6418 5795 6464
rect 5841 6418 5898 6464
rect 5944 6418 5957 6464
rect 4857 6405 5957 6418
rect 6438 6464 7098 6493
rect 6438 6418 6451 6464
rect 6497 6418 6568 6464
rect 6614 6418 6685 6464
rect 6731 6418 6803 6464
rect 6849 6418 6921 6464
rect 6967 6418 7039 6464
rect 7085 6418 7098 6464
rect 6438 6405 7098 6418
rect 8605 6464 8923 6493
rect 8605 6418 8618 6464
rect 8664 6418 8741 6464
rect 8787 6418 8864 6464
rect 8910 6418 8923 6464
rect 8605 6405 8923 6418
rect 14396 6551 14920 6580
rect 14396 6505 14409 6551
rect 14455 6505 14522 6551
rect 14568 6505 14635 6551
rect 14681 6505 14748 6551
rect 14794 6505 14861 6551
rect 14907 6505 14920 6551
rect 14396 6492 14920 6505
rect 21386 6999 23386 7028
rect 21386 6953 21399 6999
rect 23373 6953 23386 6999
rect 21386 6924 23386 6953
rect 21386 6775 23386 6804
rect 21386 6729 21399 6775
rect 23373 6729 23386 6775
rect 21386 6700 23386 6729
rect 21386 6551 23386 6580
rect 18362 6464 19462 6493
rect 18362 6418 18375 6464
rect 18421 6418 18478 6464
rect 18524 6418 18581 6464
rect 18627 6418 18684 6464
rect 18730 6418 18787 6464
rect 18833 6418 18890 6464
rect 18936 6418 18993 6464
rect 19039 6418 19096 6464
rect 19142 6418 19199 6464
rect 19449 6418 19462 6464
rect 21386 6505 21399 6551
rect 23373 6505 23386 6551
rect 21386 6492 23386 6505
rect 18362 6405 19462 6418
rect 4857 6182 5957 6195
rect 933 6095 2933 6108
rect 933 6049 946 6095
rect 2920 6049 2933 6095
rect 4857 6136 4870 6182
rect 5120 6136 5177 6182
rect 5223 6136 5280 6182
rect 5326 6136 5383 6182
rect 5429 6136 5486 6182
rect 5532 6136 5589 6182
rect 5635 6136 5692 6182
rect 5738 6136 5795 6182
rect 5841 6136 5898 6182
rect 5944 6136 5957 6182
rect 4857 6107 5957 6136
rect 6438 6182 7098 6195
rect 6438 6136 6451 6182
rect 6497 6136 6568 6182
rect 6614 6136 6685 6182
rect 6731 6136 6803 6182
rect 6849 6136 6921 6182
rect 6967 6136 7039 6182
rect 7085 6136 7098 6182
rect 6438 6107 7098 6136
rect 8605 6182 8923 6195
rect 8605 6136 8618 6182
rect 8664 6136 8741 6182
rect 8787 6136 8864 6182
rect 8910 6136 8923 6182
rect 8605 6107 8923 6136
rect 18362 6182 19462 6195
rect 933 6020 2933 6049
rect 933 5871 2933 5900
rect 933 5825 946 5871
rect 2920 5825 2933 5871
rect 933 5796 2933 5825
rect 933 5647 2933 5676
rect 933 5601 946 5647
rect 2920 5601 2933 5647
rect 933 5572 2933 5601
rect 4857 5958 5957 5987
rect 4857 5912 4870 5958
rect 5120 5912 5177 5958
rect 5223 5912 5280 5958
rect 5326 5912 5383 5958
rect 5429 5912 5486 5958
rect 5532 5912 5589 5958
rect 5635 5912 5692 5958
rect 5738 5912 5795 5958
rect 5841 5912 5898 5958
rect 5944 5912 5957 5958
rect 4857 5883 5957 5912
rect 6438 5958 7098 5987
rect 6438 5912 6451 5958
rect 6497 5912 6568 5958
rect 6614 5912 6685 5958
rect 6731 5912 6803 5958
rect 6849 5912 6921 5958
rect 6967 5912 7039 5958
rect 7085 5912 7098 5958
rect 6438 5883 7098 5912
rect 18362 6136 18375 6182
rect 18421 6136 18478 6182
rect 18524 6136 18581 6182
rect 18627 6136 18684 6182
rect 18730 6136 18787 6182
rect 18833 6136 18890 6182
rect 18936 6136 18993 6182
rect 19039 6136 19096 6182
rect 19142 6136 19199 6182
rect 19449 6136 19462 6182
rect 14396 6095 14920 6108
rect 18362 6107 19462 6136
rect 14396 6049 14409 6095
rect 14455 6049 14522 6095
rect 14568 6049 14635 6095
rect 14681 6049 14748 6095
rect 14794 6049 14861 6095
rect 14907 6049 14920 6095
rect 14396 6020 14920 6049
rect 8605 5958 8923 5987
rect 8605 5912 8618 5958
rect 8664 5912 8741 5958
rect 8787 5912 8864 5958
rect 8910 5912 8923 5958
rect 8605 5899 8923 5912
rect 21386 6095 23386 6108
rect 14396 5871 14920 5900
rect 14396 5825 14409 5871
rect 14455 5825 14522 5871
rect 14568 5825 14635 5871
rect 14681 5825 14748 5871
rect 14794 5825 14861 5871
rect 14907 5825 14920 5871
rect 14396 5796 14920 5825
rect 18362 5958 19462 5987
rect 18362 5912 18375 5958
rect 18421 5912 18478 5958
rect 18524 5912 18581 5958
rect 18627 5912 18684 5958
rect 18730 5912 18787 5958
rect 18833 5912 18890 5958
rect 18936 5912 18993 5958
rect 19039 5912 19096 5958
rect 19142 5912 19199 5958
rect 19449 5912 19462 5958
rect 18362 5883 19462 5912
rect 21386 6049 21399 6095
rect 23373 6049 23386 6095
rect 21386 6020 23386 6049
rect 4857 5734 5957 5763
rect 4857 5688 4870 5734
rect 5120 5688 5177 5734
rect 5223 5688 5280 5734
rect 5326 5688 5383 5734
rect 5429 5688 5486 5734
rect 5532 5688 5589 5734
rect 5635 5688 5692 5734
rect 5738 5688 5795 5734
rect 5841 5688 5898 5734
rect 5944 5688 5957 5734
rect 4857 5675 5957 5688
rect 6438 5734 7098 5763
rect 6438 5688 6451 5734
rect 6497 5688 6568 5734
rect 6614 5688 6685 5734
rect 6731 5688 6803 5734
rect 6849 5688 6921 5734
rect 6967 5688 7039 5734
rect 7085 5688 7098 5734
rect 6438 5675 7098 5688
rect 18362 5734 19462 5763
rect 18362 5688 18375 5734
rect 18421 5688 18478 5734
rect 18524 5688 18581 5734
rect 18627 5688 18684 5734
rect 18730 5688 18787 5734
rect 18833 5688 18890 5734
rect 18936 5688 18993 5734
rect 19039 5688 19096 5734
rect 19142 5688 19199 5734
rect 19449 5688 19462 5734
rect 14396 5647 14920 5676
rect 18362 5675 19462 5688
rect 14396 5601 14409 5647
rect 14455 5601 14522 5647
rect 14568 5601 14635 5647
rect 14681 5601 14748 5647
rect 14794 5601 14861 5647
rect 14907 5601 14920 5647
rect 933 5423 2933 5452
rect 933 5377 946 5423
rect 2920 5377 2933 5423
rect 933 5348 2933 5377
rect 933 5199 2933 5228
rect 933 5153 946 5199
rect 2920 5153 2933 5199
rect 933 5124 2933 5153
rect 933 4975 2933 5004
rect 933 4929 946 4975
rect 2920 4929 2933 4975
rect 933 4900 2933 4929
rect 14396 5572 14920 5601
rect 21386 5871 23386 5900
rect 21386 5825 21399 5871
rect 23373 5825 23386 5871
rect 21386 5796 23386 5825
rect 21386 5647 23386 5676
rect 21386 5601 21399 5647
rect 23373 5601 23386 5647
rect 21386 5572 23386 5601
rect 14396 5423 14920 5452
rect 14396 5377 14409 5423
rect 14455 5377 14522 5423
rect 14568 5377 14635 5423
rect 14681 5377 14748 5423
rect 14794 5377 14861 5423
rect 14907 5377 14920 5423
rect 14396 5348 14920 5377
rect 21386 5423 23386 5452
rect 21386 5377 21399 5423
rect 23373 5377 23386 5423
rect 21386 5348 23386 5377
rect 4857 5112 5957 5125
rect 4857 5066 4870 5112
rect 5120 5066 5177 5112
rect 5223 5066 5280 5112
rect 5326 5066 5383 5112
rect 5429 5066 5486 5112
rect 5532 5066 5589 5112
rect 5635 5066 5692 5112
rect 5738 5066 5795 5112
rect 5841 5066 5898 5112
rect 5944 5066 5957 5112
rect 4857 5037 5957 5066
rect 6438 5112 7098 5125
rect 6438 5066 6451 5112
rect 6497 5066 6568 5112
rect 6614 5066 6685 5112
rect 6731 5066 6803 5112
rect 6849 5066 6921 5112
rect 6967 5066 7039 5112
rect 7085 5066 7098 5112
rect 6438 5037 7098 5066
rect 14396 5199 14920 5228
rect 14396 5153 14409 5199
rect 14455 5153 14522 5199
rect 14568 5153 14635 5199
rect 14681 5153 14748 5199
rect 14794 5153 14861 5199
rect 14907 5153 14920 5199
rect 14396 5124 14920 5153
rect 933 4751 2933 4780
rect 933 4705 946 4751
rect 2920 4705 2933 4751
rect 4857 4888 5957 4917
rect 4857 4842 4870 4888
rect 5120 4842 5177 4888
rect 5223 4842 5280 4888
rect 5326 4842 5383 4888
rect 5429 4842 5486 4888
rect 5532 4842 5589 4888
rect 5635 4842 5692 4888
rect 5738 4842 5795 4888
rect 5841 4842 5898 4888
rect 5944 4842 5957 4888
rect 4857 4813 5957 4842
rect 933 4692 2933 4705
rect 18362 5112 19462 5125
rect 18362 5066 18375 5112
rect 18421 5066 18478 5112
rect 18524 5066 18581 5112
rect 18627 5066 18684 5112
rect 18730 5066 18787 5112
rect 18833 5066 18890 5112
rect 18936 5066 18993 5112
rect 19039 5066 19096 5112
rect 19142 5066 19199 5112
rect 19449 5066 19462 5112
rect 18362 5037 19462 5066
rect 6438 4888 7098 4917
rect 6438 4842 6451 4888
rect 6497 4842 6568 4888
rect 6614 4842 6685 4888
rect 6731 4842 6803 4888
rect 6849 4842 6921 4888
rect 6967 4842 7039 4888
rect 7085 4842 7098 4888
rect 6438 4813 7098 4842
rect 8605 4888 8923 4901
rect 8605 4842 8618 4888
rect 8664 4842 8741 4888
rect 8787 4842 8864 4888
rect 8910 4842 8923 4888
rect 8605 4813 8923 4842
rect 14396 4975 14920 5004
rect 14396 4929 14409 4975
rect 14455 4929 14522 4975
rect 14568 4929 14635 4975
rect 14681 4929 14748 4975
rect 14794 4929 14861 4975
rect 14907 4929 14920 4975
rect 14396 4900 14920 4929
rect 18362 4888 19462 4917
rect 18362 4842 18375 4888
rect 18421 4842 18478 4888
rect 18524 4842 18581 4888
rect 18627 4842 18684 4888
rect 18730 4842 18787 4888
rect 18833 4842 18890 4888
rect 18936 4842 18993 4888
rect 19039 4842 19096 4888
rect 19142 4842 19199 4888
rect 19449 4842 19462 4888
rect 18362 4813 19462 4842
rect 4857 4664 5957 4693
rect 4857 4618 4870 4664
rect 5120 4618 5177 4664
rect 5223 4618 5280 4664
rect 5326 4618 5383 4664
rect 5429 4618 5486 4664
rect 5532 4618 5589 4664
rect 5635 4618 5692 4664
rect 5738 4618 5795 4664
rect 5841 4618 5898 4664
rect 5944 4618 5957 4664
rect 4857 4605 5957 4618
rect 6438 4664 7098 4693
rect 6438 4618 6451 4664
rect 6497 4618 6568 4664
rect 6614 4618 6685 4664
rect 6731 4618 6803 4664
rect 6849 4618 6921 4664
rect 6967 4618 7039 4664
rect 7085 4618 7098 4664
rect 6438 4605 7098 4618
rect 8605 4664 8923 4693
rect 8605 4618 8618 4664
rect 8664 4618 8741 4664
rect 8787 4618 8864 4664
rect 8910 4618 8923 4664
rect 8605 4605 8923 4618
rect 14396 4751 14920 4780
rect 14396 4705 14409 4751
rect 14455 4705 14522 4751
rect 14568 4705 14635 4751
rect 14681 4705 14748 4751
rect 14794 4705 14861 4751
rect 14907 4705 14920 4751
rect 14396 4692 14920 4705
rect 21386 5199 23386 5228
rect 21386 5153 21399 5199
rect 23373 5153 23386 5199
rect 21386 5124 23386 5153
rect 21386 4975 23386 5004
rect 21386 4929 21399 4975
rect 23373 4929 23386 4975
rect 21386 4900 23386 4929
rect 21386 4751 23386 4780
rect 18362 4664 19462 4693
rect 18362 4618 18375 4664
rect 18421 4618 18478 4664
rect 18524 4618 18581 4664
rect 18627 4618 18684 4664
rect 18730 4618 18787 4664
rect 18833 4618 18890 4664
rect 18936 4618 18993 4664
rect 19039 4618 19096 4664
rect 19142 4618 19199 4664
rect 19449 4618 19462 4664
rect 21386 4705 21399 4751
rect 23373 4705 23386 4751
rect 21386 4692 23386 4705
rect 18362 4605 19462 4618
rect 4857 4382 5957 4395
rect 933 4295 2933 4308
rect 933 4249 946 4295
rect 2920 4249 2933 4295
rect 4857 4336 4870 4382
rect 5120 4336 5177 4382
rect 5223 4336 5280 4382
rect 5326 4336 5383 4382
rect 5429 4336 5486 4382
rect 5532 4336 5589 4382
rect 5635 4336 5692 4382
rect 5738 4336 5795 4382
rect 5841 4336 5898 4382
rect 5944 4336 5957 4382
rect 4857 4307 5957 4336
rect 6438 4382 7098 4395
rect 6438 4336 6451 4382
rect 6497 4336 6568 4382
rect 6614 4336 6685 4382
rect 6731 4336 6803 4382
rect 6849 4336 6921 4382
rect 6967 4336 7039 4382
rect 7085 4336 7098 4382
rect 6438 4307 7098 4336
rect 8605 4382 8923 4395
rect 8605 4336 8618 4382
rect 8664 4336 8741 4382
rect 8787 4336 8864 4382
rect 8910 4336 8923 4382
rect 8605 4307 8923 4336
rect 18362 4382 19462 4395
rect 933 4220 2933 4249
rect 933 4071 2933 4100
rect 933 4025 946 4071
rect 2920 4025 2933 4071
rect 933 3996 2933 4025
rect 933 3847 2933 3876
rect 933 3801 946 3847
rect 2920 3801 2933 3847
rect 933 3772 2933 3801
rect 4857 4158 5957 4187
rect 4857 4112 4870 4158
rect 5120 4112 5177 4158
rect 5223 4112 5280 4158
rect 5326 4112 5383 4158
rect 5429 4112 5486 4158
rect 5532 4112 5589 4158
rect 5635 4112 5692 4158
rect 5738 4112 5795 4158
rect 5841 4112 5898 4158
rect 5944 4112 5957 4158
rect 4857 4083 5957 4112
rect 6438 4158 7098 4187
rect 6438 4112 6451 4158
rect 6497 4112 6568 4158
rect 6614 4112 6685 4158
rect 6731 4112 6803 4158
rect 6849 4112 6921 4158
rect 6967 4112 7039 4158
rect 7085 4112 7098 4158
rect 6438 4083 7098 4112
rect 18362 4336 18375 4382
rect 18421 4336 18478 4382
rect 18524 4336 18581 4382
rect 18627 4336 18684 4382
rect 18730 4336 18787 4382
rect 18833 4336 18890 4382
rect 18936 4336 18993 4382
rect 19039 4336 19096 4382
rect 19142 4336 19199 4382
rect 19449 4336 19462 4382
rect 14396 4295 14920 4308
rect 18362 4307 19462 4336
rect 14396 4249 14409 4295
rect 14455 4249 14522 4295
rect 14568 4249 14635 4295
rect 14681 4249 14748 4295
rect 14794 4249 14861 4295
rect 14907 4249 14920 4295
rect 14396 4220 14920 4249
rect 8605 4158 8923 4187
rect 8605 4112 8618 4158
rect 8664 4112 8741 4158
rect 8787 4112 8864 4158
rect 8910 4112 8923 4158
rect 8605 4099 8923 4112
rect 21386 4295 23386 4308
rect 14396 4071 14920 4100
rect 14396 4025 14409 4071
rect 14455 4025 14522 4071
rect 14568 4025 14635 4071
rect 14681 4025 14748 4071
rect 14794 4025 14861 4071
rect 14907 4025 14920 4071
rect 14396 3996 14920 4025
rect 18362 4158 19462 4187
rect 18362 4112 18375 4158
rect 18421 4112 18478 4158
rect 18524 4112 18581 4158
rect 18627 4112 18684 4158
rect 18730 4112 18787 4158
rect 18833 4112 18890 4158
rect 18936 4112 18993 4158
rect 19039 4112 19096 4158
rect 19142 4112 19199 4158
rect 19449 4112 19462 4158
rect 18362 4083 19462 4112
rect 21386 4249 21399 4295
rect 23373 4249 23386 4295
rect 21386 4220 23386 4249
rect 4857 3934 5957 3963
rect 4857 3888 4870 3934
rect 5120 3888 5177 3934
rect 5223 3888 5280 3934
rect 5326 3888 5383 3934
rect 5429 3888 5486 3934
rect 5532 3888 5589 3934
rect 5635 3888 5692 3934
rect 5738 3888 5795 3934
rect 5841 3888 5898 3934
rect 5944 3888 5957 3934
rect 4857 3875 5957 3888
rect 6438 3934 7098 3963
rect 6438 3888 6451 3934
rect 6497 3888 6568 3934
rect 6614 3888 6685 3934
rect 6731 3888 6803 3934
rect 6849 3888 6921 3934
rect 6967 3888 7039 3934
rect 7085 3888 7098 3934
rect 6438 3875 7098 3888
rect 18362 3934 19462 3963
rect 18362 3888 18375 3934
rect 18421 3888 18478 3934
rect 18524 3888 18581 3934
rect 18627 3888 18684 3934
rect 18730 3888 18787 3934
rect 18833 3888 18890 3934
rect 18936 3888 18993 3934
rect 19039 3888 19096 3934
rect 19142 3888 19199 3934
rect 19449 3888 19462 3934
rect 14396 3847 14920 3876
rect 18362 3875 19462 3888
rect 14396 3801 14409 3847
rect 14455 3801 14522 3847
rect 14568 3801 14635 3847
rect 14681 3801 14748 3847
rect 14794 3801 14861 3847
rect 14907 3801 14920 3847
rect 933 3623 2933 3652
rect 933 3577 946 3623
rect 2920 3577 2933 3623
rect 933 3548 2933 3577
rect 933 3399 2933 3428
rect 933 3353 946 3399
rect 2920 3353 2933 3399
rect 933 3324 2933 3353
rect 933 3175 2933 3204
rect 933 3129 946 3175
rect 2920 3129 2933 3175
rect 933 3100 2933 3129
rect 14396 3772 14920 3801
rect 21386 4071 23386 4100
rect 21386 4025 21399 4071
rect 23373 4025 23386 4071
rect 21386 3996 23386 4025
rect 21386 3847 23386 3876
rect 21386 3801 21399 3847
rect 23373 3801 23386 3847
rect 21386 3772 23386 3801
rect 14396 3623 14920 3652
rect 14396 3577 14409 3623
rect 14455 3577 14522 3623
rect 14568 3577 14635 3623
rect 14681 3577 14748 3623
rect 14794 3577 14861 3623
rect 14907 3577 14920 3623
rect 14396 3548 14920 3577
rect 21386 3623 23386 3652
rect 21386 3577 21399 3623
rect 23373 3577 23386 3623
rect 21386 3548 23386 3577
rect 4857 3312 5957 3325
rect 4857 3266 4870 3312
rect 5120 3266 5177 3312
rect 5223 3266 5280 3312
rect 5326 3266 5383 3312
rect 5429 3266 5486 3312
rect 5532 3266 5589 3312
rect 5635 3266 5692 3312
rect 5738 3266 5795 3312
rect 5841 3266 5898 3312
rect 5944 3266 5957 3312
rect 4857 3237 5957 3266
rect 6438 3312 7098 3325
rect 6438 3266 6451 3312
rect 6497 3266 6568 3312
rect 6614 3266 6685 3312
rect 6731 3266 6803 3312
rect 6849 3266 6921 3312
rect 6967 3266 7039 3312
rect 7085 3266 7098 3312
rect 6438 3237 7098 3266
rect 14396 3399 14920 3428
rect 14396 3353 14409 3399
rect 14455 3353 14522 3399
rect 14568 3353 14635 3399
rect 14681 3353 14748 3399
rect 14794 3353 14861 3399
rect 14907 3353 14920 3399
rect 14396 3324 14920 3353
rect 933 2951 2933 2980
rect 933 2905 946 2951
rect 2920 2905 2933 2951
rect 4857 3088 5957 3117
rect 4857 3042 4870 3088
rect 5120 3042 5177 3088
rect 5223 3042 5280 3088
rect 5326 3042 5383 3088
rect 5429 3042 5486 3088
rect 5532 3042 5589 3088
rect 5635 3042 5692 3088
rect 5738 3042 5795 3088
rect 5841 3042 5898 3088
rect 5944 3042 5957 3088
rect 4857 3013 5957 3042
rect 933 2892 2933 2905
rect 18362 3312 19462 3325
rect 18362 3266 18375 3312
rect 18421 3266 18478 3312
rect 18524 3266 18581 3312
rect 18627 3266 18684 3312
rect 18730 3266 18787 3312
rect 18833 3266 18890 3312
rect 18936 3266 18993 3312
rect 19039 3266 19096 3312
rect 19142 3266 19199 3312
rect 19449 3266 19462 3312
rect 18362 3237 19462 3266
rect 6438 3088 7098 3117
rect 6438 3042 6451 3088
rect 6497 3042 6568 3088
rect 6614 3042 6685 3088
rect 6731 3042 6803 3088
rect 6849 3042 6921 3088
rect 6967 3042 7039 3088
rect 7085 3042 7098 3088
rect 6438 3013 7098 3042
rect 8605 3088 8923 3101
rect 8605 3042 8618 3088
rect 8664 3042 8741 3088
rect 8787 3042 8864 3088
rect 8910 3042 8923 3088
rect 8605 3013 8923 3042
rect 14396 3175 14920 3204
rect 14396 3129 14409 3175
rect 14455 3129 14522 3175
rect 14568 3129 14635 3175
rect 14681 3129 14748 3175
rect 14794 3129 14861 3175
rect 14907 3129 14920 3175
rect 14396 3100 14920 3129
rect 18362 3088 19462 3117
rect 18362 3042 18375 3088
rect 18421 3042 18478 3088
rect 18524 3042 18581 3088
rect 18627 3042 18684 3088
rect 18730 3042 18787 3088
rect 18833 3042 18890 3088
rect 18936 3042 18993 3088
rect 19039 3042 19096 3088
rect 19142 3042 19199 3088
rect 19449 3042 19462 3088
rect 18362 3013 19462 3042
rect 4857 2864 5957 2893
rect 4857 2818 4870 2864
rect 5120 2818 5177 2864
rect 5223 2818 5280 2864
rect 5326 2818 5383 2864
rect 5429 2818 5486 2864
rect 5532 2818 5589 2864
rect 5635 2818 5692 2864
rect 5738 2818 5795 2864
rect 5841 2818 5898 2864
rect 5944 2818 5957 2864
rect 4857 2805 5957 2818
rect 6438 2864 7098 2893
rect 6438 2818 6451 2864
rect 6497 2818 6568 2864
rect 6614 2818 6685 2864
rect 6731 2818 6803 2864
rect 6849 2818 6921 2864
rect 6967 2818 7039 2864
rect 7085 2818 7098 2864
rect 6438 2805 7098 2818
rect 8605 2864 8923 2893
rect 8605 2818 8618 2864
rect 8664 2818 8741 2864
rect 8787 2818 8864 2864
rect 8910 2818 8923 2864
rect 8605 2805 8923 2818
rect 14396 2951 14920 2980
rect 14396 2905 14409 2951
rect 14455 2905 14522 2951
rect 14568 2905 14635 2951
rect 14681 2905 14748 2951
rect 14794 2905 14861 2951
rect 14907 2905 14920 2951
rect 14396 2892 14920 2905
rect 21386 3399 23386 3428
rect 21386 3353 21399 3399
rect 23373 3353 23386 3399
rect 21386 3324 23386 3353
rect 21386 3175 23386 3204
rect 21386 3129 21399 3175
rect 23373 3129 23386 3175
rect 21386 3100 23386 3129
rect 21386 2951 23386 2980
rect 18362 2864 19462 2893
rect 18362 2818 18375 2864
rect 18421 2818 18478 2864
rect 18524 2818 18581 2864
rect 18627 2818 18684 2864
rect 18730 2818 18787 2864
rect 18833 2818 18890 2864
rect 18936 2818 18993 2864
rect 19039 2818 19096 2864
rect 19142 2818 19199 2864
rect 19449 2818 19462 2864
rect 21386 2905 21399 2951
rect 23373 2905 23386 2951
rect 21386 2892 23386 2905
rect 18362 2805 19462 2818
rect 4857 2582 5957 2595
rect 933 2495 2933 2508
rect 933 2449 946 2495
rect 2920 2449 2933 2495
rect 4857 2536 4870 2582
rect 5120 2536 5177 2582
rect 5223 2536 5280 2582
rect 5326 2536 5383 2582
rect 5429 2536 5486 2582
rect 5532 2536 5589 2582
rect 5635 2536 5692 2582
rect 5738 2536 5795 2582
rect 5841 2536 5898 2582
rect 5944 2536 5957 2582
rect 4857 2507 5957 2536
rect 6438 2582 7098 2595
rect 6438 2536 6451 2582
rect 6497 2536 6568 2582
rect 6614 2536 6685 2582
rect 6731 2536 6803 2582
rect 6849 2536 6921 2582
rect 6967 2536 7039 2582
rect 7085 2536 7098 2582
rect 6438 2507 7098 2536
rect 8605 2582 8923 2595
rect 8605 2536 8618 2582
rect 8664 2536 8741 2582
rect 8787 2536 8864 2582
rect 8910 2536 8923 2582
rect 8605 2507 8923 2536
rect 18362 2582 19462 2595
rect 933 2420 2933 2449
rect 933 2271 2933 2300
rect 933 2225 946 2271
rect 2920 2225 2933 2271
rect 933 2196 2933 2225
rect 933 2047 2933 2076
rect 933 2001 946 2047
rect 2920 2001 2933 2047
rect 933 1972 2933 2001
rect 4857 2358 5957 2387
rect 4857 2312 4870 2358
rect 5120 2312 5177 2358
rect 5223 2312 5280 2358
rect 5326 2312 5383 2358
rect 5429 2312 5486 2358
rect 5532 2312 5589 2358
rect 5635 2312 5692 2358
rect 5738 2312 5795 2358
rect 5841 2312 5898 2358
rect 5944 2312 5957 2358
rect 4857 2283 5957 2312
rect 6438 2358 7098 2387
rect 6438 2312 6451 2358
rect 6497 2312 6568 2358
rect 6614 2312 6685 2358
rect 6731 2312 6803 2358
rect 6849 2312 6921 2358
rect 6967 2312 7039 2358
rect 7085 2312 7098 2358
rect 6438 2283 7098 2312
rect 18362 2536 18375 2582
rect 18421 2536 18478 2582
rect 18524 2536 18581 2582
rect 18627 2536 18684 2582
rect 18730 2536 18787 2582
rect 18833 2536 18890 2582
rect 18936 2536 18993 2582
rect 19039 2536 19096 2582
rect 19142 2536 19199 2582
rect 19449 2536 19462 2582
rect 14396 2495 14920 2508
rect 18362 2507 19462 2536
rect 14396 2449 14409 2495
rect 14455 2449 14522 2495
rect 14568 2449 14635 2495
rect 14681 2449 14748 2495
rect 14794 2449 14861 2495
rect 14907 2449 14920 2495
rect 14396 2420 14920 2449
rect 8605 2358 8923 2387
rect 8605 2312 8618 2358
rect 8664 2312 8741 2358
rect 8787 2312 8864 2358
rect 8910 2312 8923 2358
rect 8605 2299 8923 2312
rect 21386 2495 23386 2508
rect 14396 2271 14920 2300
rect 14396 2225 14409 2271
rect 14455 2225 14522 2271
rect 14568 2225 14635 2271
rect 14681 2225 14748 2271
rect 14794 2225 14861 2271
rect 14907 2225 14920 2271
rect 14396 2196 14920 2225
rect 18362 2358 19462 2387
rect 18362 2312 18375 2358
rect 18421 2312 18478 2358
rect 18524 2312 18581 2358
rect 18627 2312 18684 2358
rect 18730 2312 18787 2358
rect 18833 2312 18890 2358
rect 18936 2312 18993 2358
rect 19039 2312 19096 2358
rect 19142 2312 19199 2358
rect 19449 2312 19462 2358
rect 18362 2283 19462 2312
rect 21386 2449 21399 2495
rect 23373 2449 23386 2495
rect 21386 2420 23386 2449
rect 4857 2134 5957 2163
rect 4857 2088 4870 2134
rect 5120 2088 5177 2134
rect 5223 2088 5280 2134
rect 5326 2088 5383 2134
rect 5429 2088 5486 2134
rect 5532 2088 5589 2134
rect 5635 2088 5692 2134
rect 5738 2088 5795 2134
rect 5841 2088 5898 2134
rect 5944 2088 5957 2134
rect 4857 2075 5957 2088
rect 6438 2134 7098 2163
rect 6438 2088 6451 2134
rect 6497 2088 6568 2134
rect 6614 2088 6685 2134
rect 6731 2088 6803 2134
rect 6849 2088 6921 2134
rect 6967 2088 7039 2134
rect 7085 2088 7098 2134
rect 6438 2075 7098 2088
rect 18362 2134 19462 2163
rect 18362 2088 18375 2134
rect 18421 2088 18478 2134
rect 18524 2088 18581 2134
rect 18627 2088 18684 2134
rect 18730 2088 18787 2134
rect 18833 2088 18890 2134
rect 18936 2088 18993 2134
rect 19039 2088 19096 2134
rect 19142 2088 19199 2134
rect 19449 2088 19462 2134
rect 14396 2047 14920 2076
rect 18362 2075 19462 2088
rect 14396 2001 14409 2047
rect 14455 2001 14522 2047
rect 14568 2001 14635 2047
rect 14681 2001 14748 2047
rect 14794 2001 14861 2047
rect 14907 2001 14920 2047
rect 933 1823 2933 1852
rect 933 1777 946 1823
rect 2920 1777 2933 1823
rect 933 1748 2933 1777
rect 933 1599 2933 1628
rect 933 1553 946 1599
rect 2920 1553 2933 1599
rect 933 1524 2933 1553
rect 933 1375 2933 1404
rect 933 1329 946 1375
rect 2920 1329 2933 1375
rect 933 1300 2933 1329
rect 14396 1972 14920 2001
rect 21386 2271 23386 2300
rect 21386 2225 21399 2271
rect 23373 2225 23386 2271
rect 21386 2196 23386 2225
rect 21386 2047 23386 2076
rect 21386 2001 21399 2047
rect 23373 2001 23386 2047
rect 21386 1972 23386 2001
rect 14396 1823 14920 1852
rect 14396 1777 14409 1823
rect 14455 1777 14522 1823
rect 14568 1777 14635 1823
rect 14681 1777 14748 1823
rect 14794 1777 14861 1823
rect 14907 1777 14920 1823
rect 14396 1748 14920 1777
rect 21386 1823 23386 1852
rect 21386 1777 21399 1823
rect 23373 1777 23386 1823
rect 21386 1748 23386 1777
rect 4857 1512 5957 1525
rect 4857 1466 4870 1512
rect 5120 1466 5177 1512
rect 5223 1466 5280 1512
rect 5326 1466 5383 1512
rect 5429 1466 5486 1512
rect 5532 1466 5589 1512
rect 5635 1466 5692 1512
rect 5738 1466 5795 1512
rect 5841 1466 5898 1512
rect 5944 1466 5957 1512
rect 4857 1437 5957 1466
rect 6438 1512 7098 1525
rect 6438 1466 6451 1512
rect 6497 1466 6568 1512
rect 6614 1466 6685 1512
rect 6731 1466 6803 1512
rect 6849 1466 6921 1512
rect 6967 1466 7039 1512
rect 7085 1466 7098 1512
rect 6438 1437 7098 1466
rect 14396 1599 14920 1628
rect 14396 1553 14409 1599
rect 14455 1553 14522 1599
rect 14568 1553 14635 1599
rect 14681 1553 14748 1599
rect 14794 1553 14861 1599
rect 14907 1553 14920 1599
rect 14396 1524 14920 1553
rect 933 1151 2933 1180
rect 933 1105 946 1151
rect 2920 1105 2933 1151
rect 4857 1288 5957 1317
rect 4857 1242 4870 1288
rect 5120 1242 5177 1288
rect 5223 1242 5280 1288
rect 5326 1242 5383 1288
rect 5429 1242 5486 1288
rect 5532 1242 5589 1288
rect 5635 1242 5692 1288
rect 5738 1242 5795 1288
rect 5841 1242 5898 1288
rect 5944 1242 5957 1288
rect 4857 1213 5957 1242
rect 933 1092 2933 1105
rect 18362 1512 19462 1525
rect 18362 1466 18375 1512
rect 18421 1466 18478 1512
rect 18524 1466 18581 1512
rect 18627 1466 18684 1512
rect 18730 1466 18787 1512
rect 18833 1466 18890 1512
rect 18936 1466 18993 1512
rect 19039 1466 19096 1512
rect 19142 1466 19199 1512
rect 19449 1466 19462 1512
rect 18362 1437 19462 1466
rect 6438 1288 7098 1317
rect 6438 1242 6451 1288
rect 6497 1242 6568 1288
rect 6614 1242 6685 1288
rect 6731 1242 6803 1288
rect 6849 1242 6921 1288
rect 6967 1242 7039 1288
rect 7085 1242 7098 1288
rect 6438 1213 7098 1242
rect 8605 1288 8923 1301
rect 8605 1242 8618 1288
rect 8664 1242 8741 1288
rect 8787 1242 8864 1288
rect 8910 1242 8923 1288
rect 8605 1213 8923 1242
rect 14396 1375 14920 1404
rect 14396 1329 14409 1375
rect 14455 1329 14522 1375
rect 14568 1329 14635 1375
rect 14681 1329 14748 1375
rect 14794 1329 14861 1375
rect 14907 1329 14920 1375
rect 14396 1300 14920 1329
rect 18362 1288 19462 1317
rect 18362 1242 18375 1288
rect 18421 1242 18478 1288
rect 18524 1242 18581 1288
rect 18627 1242 18684 1288
rect 18730 1242 18787 1288
rect 18833 1242 18890 1288
rect 18936 1242 18993 1288
rect 19039 1242 19096 1288
rect 19142 1242 19199 1288
rect 19449 1242 19462 1288
rect 18362 1213 19462 1242
rect 4857 1064 5957 1093
rect 4857 1018 4870 1064
rect 5120 1018 5177 1064
rect 5223 1018 5280 1064
rect 5326 1018 5383 1064
rect 5429 1018 5486 1064
rect 5532 1018 5589 1064
rect 5635 1018 5692 1064
rect 5738 1018 5795 1064
rect 5841 1018 5898 1064
rect 5944 1018 5957 1064
rect 4857 1005 5957 1018
rect 6438 1064 7098 1093
rect 6438 1018 6451 1064
rect 6497 1018 6568 1064
rect 6614 1018 6685 1064
rect 6731 1018 6803 1064
rect 6849 1018 6921 1064
rect 6967 1018 7039 1064
rect 7085 1018 7098 1064
rect 6438 1005 7098 1018
rect 8605 1064 8923 1093
rect 8605 1018 8618 1064
rect 8664 1018 8741 1064
rect 8787 1018 8864 1064
rect 8910 1018 8923 1064
rect 8605 1005 8923 1018
rect 14396 1151 14920 1180
rect 14396 1105 14409 1151
rect 14455 1105 14522 1151
rect 14568 1105 14635 1151
rect 14681 1105 14748 1151
rect 14794 1105 14861 1151
rect 14907 1105 14920 1151
rect 14396 1092 14920 1105
rect 21386 1599 23386 1628
rect 21386 1553 21399 1599
rect 23373 1553 23386 1599
rect 21386 1524 23386 1553
rect 21386 1375 23386 1404
rect 21386 1329 21399 1375
rect 23373 1329 23386 1375
rect 21386 1300 23386 1329
rect 21386 1151 23386 1180
rect 18362 1064 19462 1093
rect 18362 1018 18375 1064
rect 18421 1018 18478 1064
rect 18524 1018 18581 1064
rect 18627 1018 18684 1064
rect 18730 1018 18787 1064
rect 18833 1018 18890 1064
rect 18936 1018 18993 1064
rect 19039 1018 19096 1064
rect 19142 1018 19199 1064
rect 19449 1018 19462 1064
rect 21386 1105 21399 1151
rect 23373 1105 23386 1151
rect 21386 1092 23386 1105
rect 18362 1005 19462 1018
rect 4857 782 5957 795
rect 933 695 2933 708
rect 933 649 946 695
rect 2920 649 2933 695
rect 4857 736 4870 782
rect 5120 736 5177 782
rect 5223 736 5280 782
rect 5326 736 5383 782
rect 5429 736 5486 782
rect 5532 736 5589 782
rect 5635 736 5692 782
rect 5738 736 5795 782
rect 5841 736 5898 782
rect 5944 736 5957 782
rect 4857 707 5957 736
rect 6438 782 7098 795
rect 6438 736 6451 782
rect 6497 736 6568 782
rect 6614 736 6685 782
rect 6731 736 6803 782
rect 6849 736 6921 782
rect 6967 736 7039 782
rect 7085 736 7098 782
rect 6438 707 7098 736
rect 8605 782 8923 795
rect 8605 736 8618 782
rect 8664 736 8741 782
rect 8787 736 8864 782
rect 8910 736 8923 782
rect 8605 707 8923 736
rect 18362 782 19462 795
rect 933 620 2933 649
rect 933 471 2933 500
rect 933 425 946 471
rect 2920 425 2933 471
rect 933 396 2933 425
rect 933 247 2933 276
rect 933 201 946 247
rect 2920 201 2933 247
rect 933 172 2933 201
rect 4857 558 5957 587
rect 4857 512 4870 558
rect 5120 512 5177 558
rect 5223 512 5280 558
rect 5326 512 5383 558
rect 5429 512 5486 558
rect 5532 512 5589 558
rect 5635 512 5692 558
rect 5738 512 5795 558
rect 5841 512 5898 558
rect 5944 512 5957 558
rect 4857 483 5957 512
rect 6438 558 7098 587
rect 6438 512 6451 558
rect 6497 512 6568 558
rect 6614 512 6685 558
rect 6731 512 6803 558
rect 6849 512 6921 558
rect 6967 512 7039 558
rect 7085 512 7098 558
rect 6438 483 7098 512
rect 18362 736 18375 782
rect 18421 736 18478 782
rect 18524 736 18581 782
rect 18627 736 18684 782
rect 18730 736 18787 782
rect 18833 736 18890 782
rect 18936 736 18993 782
rect 19039 736 19096 782
rect 19142 736 19199 782
rect 19449 736 19462 782
rect 14396 695 14920 708
rect 18362 707 19462 736
rect 14396 649 14409 695
rect 14455 649 14522 695
rect 14568 649 14635 695
rect 14681 649 14748 695
rect 14794 649 14861 695
rect 14907 649 14920 695
rect 14396 620 14920 649
rect 8605 558 8923 587
rect 8605 512 8618 558
rect 8664 512 8741 558
rect 8787 512 8864 558
rect 8910 512 8923 558
rect 8605 499 8923 512
rect 21386 695 23386 708
rect 14396 471 14920 500
rect 14396 425 14409 471
rect 14455 425 14522 471
rect 14568 425 14635 471
rect 14681 425 14748 471
rect 14794 425 14861 471
rect 14907 425 14920 471
rect 14396 396 14920 425
rect 18362 558 19462 587
rect 18362 512 18375 558
rect 18421 512 18478 558
rect 18524 512 18581 558
rect 18627 512 18684 558
rect 18730 512 18787 558
rect 18833 512 18890 558
rect 18936 512 18993 558
rect 19039 512 19096 558
rect 19142 512 19199 558
rect 19449 512 19462 558
rect 18362 483 19462 512
rect 21386 649 21399 695
rect 23373 649 23386 695
rect 21386 620 23386 649
rect 4857 334 5957 363
rect 4857 288 4870 334
rect 5120 288 5177 334
rect 5223 288 5280 334
rect 5326 288 5383 334
rect 5429 288 5486 334
rect 5532 288 5589 334
rect 5635 288 5692 334
rect 5738 288 5795 334
rect 5841 288 5898 334
rect 5944 288 5957 334
rect 4857 275 5957 288
rect 6438 334 7098 363
rect 6438 288 6451 334
rect 6497 288 6568 334
rect 6614 288 6685 334
rect 6731 288 6803 334
rect 6849 288 6921 334
rect 6967 288 7039 334
rect 7085 288 7098 334
rect 6438 275 7098 288
rect 18362 334 19462 363
rect 18362 288 18375 334
rect 18421 288 18478 334
rect 18524 288 18581 334
rect 18627 288 18684 334
rect 18730 288 18787 334
rect 18833 288 18890 334
rect 18936 288 18993 334
rect 19039 288 19096 334
rect 19142 288 19199 334
rect 19449 288 19462 334
rect 14396 247 14920 276
rect 18362 275 19462 288
rect 14396 201 14409 247
rect 14455 201 14522 247
rect 14568 201 14635 247
rect 14681 201 14748 247
rect 14794 201 14861 247
rect 14907 201 14920 247
rect 933 23 2933 52
rect 933 -23 946 23
rect 2920 -23 2933 23
rect 933 -36 2933 -23
rect 14396 172 14920 201
rect 21386 471 23386 500
rect 21386 425 21399 471
rect 23373 425 23386 471
rect 21386 396 23386 425
rect 21386 247 23386 276
rect 21386 201 21399 247
rect 23373 201 23386 247
rect 21386 172 23386 201
rect 14396 23 14920 52
rect 14396 -23 14409 23
rect 14455 -23 14522 23
rect 14568 -23 14635 23
rect 14681 -23 14748 23
rect 14794 -23 14861 23
rect 14907 -23 14920 23
rect 14396 -36 14920 -23
rect 21386 23 23386 52
rect 21386 -23 21399 23
rect 23373 -23 23386 23
rect 21386 -36 23386 -23
<< ndiffc >>
rect 13336 14377 13382 14423
rect 13503 14377 13549 14423
rect 13668 14377 13714 14423
rect 13833 14377 13879 14423
rect 3413 13670 3459 13716
rect 3599 13670 3645 13716
rect 3786 13670 3832 13716
rect 3973 13670 4019 13716
rect 4159 13670 4205 13716
rect 13336 13684 13382 13730
rect 13503 13684 13549 13730
rect 13668 13684 13714 13730
rect 13833 13684 13879 13730
rect 20113 13670 20159 13716
rect 20300 13670 20346 13716
rect 20487 13670 20533 13716
rect 20673 13670 20719 13716
rect 20860 13670 20906 13716
rect 3413 13284 3459 13330
rect 3599 13284 3645 13330
rect 3786 13284 3832 13330
rect 3973 13284 4019 13330
rect 4159 13284 4205 13330
rect 13336 13270 13382 13316
rect 13503 13270 13549 13316
rect 13668 13270 13714 13316
rect 13833 13270 13879 13316
rect 20113 13284 20159 13330
rect 20300 13284 20346 13330
rect 20487 13284 20533 13330
rect 20673 13284 20719 13330
rect 20860 13284 20906 13330
rect 13336 12577 13382 12623
rect 13503 12577 13549 12623
rect 13668 12577 13714 12623
rect 13833 12577 13879 12623
rect 3413 11870 3459 11916
rect 3599 11870 3645 11916
rect 3786 11870 3832 11916
rect 3973 11870 4019 11916
rect 4159 11870 4205 11916
rect 13336 11884 13382 11930
rect 13503 11884 13549 11930
rect 13668 11884 13714 11930
rect 13833 11884 13879 11930
rect 20113 11870 20159 11916
rect 20300 11870 20346 11916
rect 20487 11870 20533 11916
rect 20673 11870 20719 11916
rect 20860 11870 20906 11916
rect 3413 11484 3459 11530
rect 3599 11484 3645 11530
rect 3786 11484 3832 11530
rect 3973 11484 4019 11530
rect 4159 11484 4205 11530
rect 13336 11470 13382 11516
rect 13503 11470 13549 11516
rect 13668 11470 13714 11516
rect 13833 11470 13879 11516
rect 20113 11484 20159 11530
rect 20300 11484 20346 11530
rect 20487 11484 20533 11530
rect 20673 11484 20719 11530
rect 20860 11484 20906 11530
rect 13336 10777 13382 10823
rect 13503 10777 13549 10823
rect 13668 10777 13714 10823
rect 13833 10777 13879 10823
rect 3413 10070 3459 10116
rect 3599 10070 3645 10116
rect 3786 10070 3832 10116
rect 3973 10070 4019 10116
rect 4159 10070 4205 10116
rect 13336 10084 13382 10130
rect 13503 10084 13549 10130
rect 13668 10084 13714 10130
rect 13833 10084 13879 10130
rect 20113 10070 20159 10116
rect 20300 10070 20346 10116
rect 20487 10070 20533 10116
rect 20673 10070 20719 10116
rect 20860 10070 20906 10116
rect 3413 9684 3459 9730
rect 3599 9684 3645 9730
rect 3786 9684 3832 9730
rect 3973 9684 4019 9730
rect 4159 9684 4205 9730
rect 13336 9670 13382 9716
rect 13503 9670 13549 9716
rect 13668 9670 13714 9716
rect 13833 9670 13879 9716
rect 20113 9684 20159 9730
rect 20300 9684 20346 9730
rect 20487 9684 20533 9730
rect 20673 9684 20719 9730
rect 20860 9684 20906 9730
rect 13336 8977 13382 9023
rect 13503 8977 13549 9023
rect 13668 8977 13714 9023
rect 13833 8977 13879 9023
rect 3413 8270 3459 8316
rect 3599 8270 3645 8316
rect 3786 8270 3832 8316
rect 3973 8270 4019 8316
rect 4159 8270 4205 8316
rect 13336 8284 13382 8330
rect 13503 8284 13549 8330
rect 13668 8284 13714 8330
rect 13833 8284 13879 8330
rect 20113 8270 20159 8316
rect 20300 8270 20346 8316
rect 20487 8270 20533 8316
rect 20673 8270 20719 8316
rect 20860 8270 20906 8316
rect 3413 7884 3459 7930
rect 3599 7884 3645 7930
rect 3786 7884 3832 7930
rect 3973 7884 4019 7930
rect 4159 7884 4205 7930
rect 13336 7870 13382 7916
rect 13503 7870 13549 7916
rect 13668 7870 13714 7916
rect 13833 7870 13879 7916
rect 20113 7884 20159 7930
rect 20300 7884 20346 7930
rect 20487 7884 20533 7930
rect 20673 7884 20719 7930
rect 20860 7884 20906 7930
rect 13336 7177 13382 7223
rect 13503 7177 13549 7223
rect 13668 7177 13714 7223
rect 13833 7177 13879 7223
rect 3413 6470 3459 6516
rect 3599 6470 3645 6516
rect 3786 6470 3832 6516
rect 3973 6470 4019 6516
rect 4159 6470 4205 6516
rect 13336 6484 13382 6530
rect 13503 6484 13549 6530
rect 13668 6484 13714 6530
rect 13833 6484 13879 6530
rect 20113 6470 20159 6516
rect 20300 6470 20346 6516
rect 20487 6470 20533 6516
rect 20673 6470 20719 6516
rect 20860 6470 20906 6516
rect 3413 6084 3459 6130
rect 3599 6084 3645 6130
rect 3786 6084 3832 6130
rect 3973 6084 4019 6130
rect 4159 6084 4205 6130
rect 13336 6070 13382 6116
rect 13503 6070 13549 6116
rect 13668 6070 13714 6116
rect 13833 6070 13879 6116
rect 20113 6084 20159 6130
rect 20300 6084 20346 6130
rect 20487 6084 20533 6130
rect 20673 6084 20719 6130
rect 20860 6084 20906 6130
rect 13336 5377 13382 5423
rect 13503 5377 13549 5423
rect 13668 5377 13714 5423
rect 13833 5377 13879 5423
rect 3413 4670 3459 4716
rect 3599 4670 3645 4716
rect 3786 4670 3832 4716
rect 3973 4670 4019 4716
rect 4159 4670 4205 4716
rect 13336 4684 13382 4730
rect 13503 4684 13549 4730
rect 13668 4684 13714 4730
rect 13833 4684 13879 4730
rect 20113 4670 20159 4716
rect 20300 4670 20346 4716
rect 20487 4670 20533 4716
rect 20673 4670 20719 4716
rect 20860 4670 20906 4716
rect 3413 4284 3459 4330
rect 3599 4284 3645 4330
rect 3786 4284 3832 4330
rect 3973 4284 4019 4330
rect 4159 4284 4205 4330
rect 13336 4270 13382 4316
rect 13503 4270 13549 4316
rect 13668 4270 13714 4316
rect 13833 4270 13879 4316
rect 20113 4284 20159 4330
rect 20300 4284 20346 4330
rect 20487 4284 20533 4330
rect 20673 4284 20719 4330
rect 20860 4284 20906 4330
rect 13336 3577 13382 3623
rect 13503 3577 13549 3623
rect 13668 3577 13714 3623
rect 13833 3577 13879 3623
rect 3413 2870 3459 2916
rect 3599 2870 3645 2916
rect 3786 2870 3832 2916
rect 3973 2870 4019 2916
rect 4159 2870 4205 2916
rect 13336 2884 13382 2930
rect 13503 2884 13549 2930
rect 13668 2884 13714 2930
rect 13833 2884 13879 2930
rect 20113 2870 20159 2916
rect 20300 2870 20346 2916
rect 20487 2870 20533 2916
rect 20673 2870 20719 2916
rect 20860 2870 20906 2916
rect 3413 2484 3459 2530
rect 3599 2484 3645 2530
rect 3786 2484 3832 2530
rect 3973 2484 4019 2530
rect 4159 2484 4205 2530
rect 13336 2470 13382 2516
rect 13503 2470 13549 2516
rect 13668 2470 13714 2516
rect 13833 2470 13879 2516
rect 20113 2484 20159 2530
rect 20300 2484 20346 2530
rect 20487 2484 20533 2530
rect 20673 2484 20719 2530
rect 20860 2484 20906 2530
rect 13336 1777 13382 1823
rect 13503 1777 13549 1823
rect 13668 1777 13714 1823
rect 13833 1777 13879 1823
rect 3413 1070 3459 1116
rect 3599 1070 3645 1116
rect 3786 1070 3832 1116
rect 3973 1070 4019 1116
rect 4159 1070 4205 1116
rect 13336 1084 13382 1130
rect 13503 1084 13549 1130
rect 13668 1084 13714 1130
rect 13833 1084 13879 1130
rect 20113 1070 20159 1116
rect 20300 1070 20346 1116
rect 20487 1070 20533 1116
rect 20673 1070 20719 1116
rect 20860 1070 20906 1116
rect 3413 684 3459 730
rect 3599 684 3645 730
rect 3786 684 3832 730
rect 3973 684 4019 730
rect 4159 684 4205 730
rect 13336 670 13382 716
rect 13503 670 13549 716
rect 13668 670 13714 716
rect 13833 670 13879 716
rect 20113 684 20159 730
rect 20300 684 20346 730
rect 20487 684 20533 730
rect 20673 684 20719 730
rect 20860 684 20906 730
rect 13336 -23 13382 23
rect 13503 -23 13549 23
rect 13668 -23 13714 23
rect 13833 -23 13879 23
<< mvndiffc >>
rect 3281 14377 3327 14423
rect 3384 14377 3430 14423
rect 3487 14377 3533 14423
rect 3590 14377 3636 14423
rect 3693 14377 3739 14423
rect 3796 14377 3842 14423
rect 3899 14377 3945 14423
rect 4002 14377 4048 14423
rect 4105 14377 4151 14423
rect 4209 14377 4255 14423
rect 9337 14377 9383 14423
rect 9459 14377 9505 14423
rect 9582 14377 9628 14423
rect 9705 14377 9751 14423
rect 3281 14153 3327 14199
rect 3384 14153 3430 14199
rect 3487 14153 3533 14199
rect 3590 14153 3636 14199
rect 3693 14153 3739 14199
rect 3796 14153 3842 14199
rect 3899 14153 3945 14199
rect 4002 14153 4048 14199
rect 4105 14153 4151 14199
rect 4209 14153 4255 14199
rect 9337 14153 9383 14199
rect 9459 14153 9505 14199
rect 9582 14153 9628 14199
rect 9705 14153 9751 14199
rect 20064 14377 20110 14423
rect 20168 14377 20214 14423
rect 20271 14377 20317 14423
rect 20374 14377 20420 14423
rect 20477 14377 20523 14423
rect 20580 14377 20626 14423
rect 20683 14377 20729 14423
rect 20786 14377 20832 14423
rect 20889 14377 20935 14423
rect 20992 14377 21038 14423
rect 20064 14153 20110 14199
rect 20168 14153 20214 14199
rect 20271 14153 20317 14199
rect 20374 14153 20420 14199
rect 20477 14153 20523 14199
rect 20580 14153 20626 14199
rect 20683 14153 20729 14199
rect 20786 14153 20832 14199
rect 20889 14153 20935 14199
rect 20992 14153 21038 14199
rect 7506 14066 7552 14112
rect 7623 14066 7669 14112
rect 7740 14066 7786 14112
rect 7858 14066 7904 14112
rect 7976 14066 8022 14112
rect 8094 14066 8140 14112
rect 3281 13929 3327 13975
rect 3384 13929 3430 13975
rect 3487 13929 3533 13975
rect 3590 13929 3636 13975
rect 3693 13929 3739 13975
rect 3796 13929 3842 13975
rect 3899 13929 3945 13975
rect 4002 13929 4048 13975
rect 4105 13929 4151 13975
rect 4209 13929 4255 13975
rect 7506 13842 7552 13888
rect 7623 13842 7669 13888
rect 7740 13842 7786 13888
rect 7858 13842 7904 13888
rect 7976 13842 8022 13888
rect 8094 13842 8140 13888
rect 9238 13842 9284 13888
rect 20064 13929 20110 13975
rect 20168 13929 20214 13975
rect 20271 13929 20317 13975
rect 20374 13929 20420 13975
rect 20477 13929 20523 13975
rect 20580 13929 20626 13975
rect 20683 13929 20729 13975
rect 20786 13929 20832 13975
rect 20889 13929 20935 13975
rect 20992 13929 21038 13975
rect 7506 13618 7552 13664
rect 7623 13618 7669 13664
rect 7740 13618 7786 13664
rect 7858 13618 7904 13664
rect 7976 13618 8022 13664
rect 8094 13618 8140 13664
rect 9238 13618 9284 13664
rect 7506 13336 7552 13382
rect 7623 13336 7669 13382
rect 7740 13336 7786 13382
rect 7858 13336 7904 13382
rect 7976 13336 8022 13382
rect 8094 13336 8140 13382
rect 9238 13336 9284 13382
rect 3281 13025 3327 13071
rect 3384 13025 3430 13071
rect 3487 13025 3533 13071
rect 3590 13025 3636 13071
rect 3693 13025 3739 13071
rect 3796 13025 3842 13071
rect 3899 13025 3945 13071
rect 4002 13025 4048 13071
rect 4105 13025 4151 13071
rect 4209 13025 4255 13071
rect 7506 13112 7552 13158
rect 7623 13112 7669 13158
rect 7740 13112 7786 13158
rect 7858 13112 7904 13158
rect 7976 13112 8022 13158
rect 8094 13112 8140 13158
rect 9238 13112 9284 13158
rect 7506 12888 7552 12934
rect 7623 12888 7669 12934
rect 7740 12888 7786 12934
rect 7858 12888 7904 12934
rect 7976 12888 8022 12934
rect 8094 12888 8140 12934
rect 20064 13025 20110 13071
rect 20168 13025 20214 13071
rect 20271 13025 20317 13071
rect 20374 13025 20420 13071
rect 20477 13025 20523 13071
rect 20580 13025 20626 13071
rect 20683 13025 20729 13071
rect 20786 13025 20832 13071
rect 20889 13025 20935 13071
rect 20992 13025 21038 13071
rect 3281 12801 3327 12847
rect 3384 12801 3430 12847
rect 3487 12801 3533 12847
rect 3590 12801 3636 12847
rect 3693 12801 3739 12847
rect 3796 12801 3842 12847
rect 3899 12801 3945 12847
rect 4002 12801 4048 12847
rect 4105 12801 4151 12847
rect 4209 12801 4255 12847
rect 9337 12801 9383 12847
rect 9459 12801 9505 12847
rect 9582 12801 9628 12847
rect 9705 12801 9751 12847
rect 3281 12577 3327 12623
rect 3384 12577 3430 12623
rect 3487 12577 3533 12623
rect 3590 12577 3636 12623
rect 3693 12577 3739 12623
rect 3796 12577 3842 12623
rect 3899 12577 3945 12623
rect 4002 12577 4048 12623
rect 4105 12577 4151 12623
rect 4209 12577 4255 12623
rect 9337 12577 9383 12623
rect 9459 12577 9505 12623
rect 9582 12577 9628 12623
rect 9705 12577 9751 12623
rect 20064 12801 20110 12847
rect 20168 12801 20214 12847
rect 20271 12801 20317 12847
rect 20374 12801 20420 12847
rect 20477 12801 20523 12847
rect 20580 12801 20626 12847
rect 20683 12801 20729 12847
rect 20786 12801 20832 12847
rect 20889 12801 20935 12847
rect 20992 12801 21038 12847
rect 3281 12353 3327 12399
rect 3384 12353 3430 12399
rect 3487 12353 3533 12399
rect 3590 12353 3636 12399
rect 3693 12353 3739 12399
rect 3796 12353 3842 12399
rect 3899 12353 3945 12399
rect 4002 12353 4048 12399
rect 4105 12353 4151 12399
rect 4209 12353 4255 12399
rect 9337 12353 9383 12399
rect 9459 12353 9505 12399
rect 9582 12353 9628 12399
rect 9705 12353 9751 12399
rect 20064 12577 20110 12623
rect 20168 12577 20214 12623
rect 20271 12577 20317 12623
rect 20374 12577 20420 12623
rect 20477 12577 20523 12623
rect 20580 12577 20626 12623
rect 20683 12577 20729 12623
rect 20786 12577 20832 12623
rect 20889 12577 20935 12623
rect 20992 12577 21038 12623
rect 20064 12353 20110 12399
rect 20168 12353 20214 12399
rect 20271 12353 20317 12399
rect 20374 12353 20420 12399
rect 20477 12353 20523 12399
rect 20580 12353 20626 12399
rect 20683 12353 20729 12399
rect 20786 12353 20832 12399
rect 20889 12353 20935 12399
rect 20992 12353 21038 12399
rect 7506 12266 7552 12312
rect 7623 12266 7669 12312
rect 7740 12266 7786 12312
rect 7858 12266 7904 12312
rect 7976 12266 8022 12312
rect 8094 12266 8140 12312
rect 3281 12129 3327 12175
rect 3384 12129 3430 12175
rect 3487 12129 3533 12175
rect 3590 12129 3636 12175
rect 3693 12129 3739 12175
rect 3796 12129 3842 12175
rect 3899 12129 3945 12175
rect 4002 12129 4048 12175
rect 4105 12129 4151 12175
rect 4209 12129 4255 12175
rect 7506 12042 7552 12088
rect 7623 12042 7669 12088
rect 7740 12042 7786 12088
rect 7858 12042 7904 12088
rect 7976 12042 8022 12088
rect 8094 12042 8140 12088
rect 9238 12042 9284 12088
rect 20064 12129 20110 12175
rect 20168 12129 20214 12175
rect 20271 12129 20317 12175
rect 20374 12129 20420 12175
rect 20477 12129 20523 12175
rect 20580 12129 20626 12175
rect 20683 12129 20729 12175
rect 20786 12129 20832 12175
rect 20889 12129 20935 12175
rect 20992 12129 21038 12175
rect 7506 11818 7552 11864
rect 7623 11818 7669 11864
rect 7740 11818 7786 11864
rect 7858 11818 7904 11864
rect 7976 11818 8022 11864
rect 8094 11818 8140 11864
rect 9238 11818 9284 11864
rect 7506 11536 7552 11582
rect 7623 11536 7669 11582
rect 7740 11536 7786 11582
rect 7858 11536 7904 11582
rect 7976 11536 8022 11582
rect 8094 11536 8140 11582
rect 9238 11536 9284 11582
rect 3281 11225 3327 11271
rect 3384 11225 3430 11271
rect 3487 11225 3533 11271
rect 3590 11225 3636 11271
rect 3693 11225 3739 11271
rect 3796 11225 3842 11271
rect 3899 11225 3945 11271
rect 4002 11225 4048 11271
rect 4105 11225 4151 11271
rect 4209 11225 4255 11271
rect 7506 11312 7552 11358
rect 7623 11312 7669 11358
rect 7740 11312 7786 11358
rect 7858 11312 7904 11358
rect 7976 11312 8022 11358
rect 8094 11312 8140 11358
rect 9238 11312 9284 11358
rect 7506 11088 7552 11134
rect 7623 11088 7669 11134
rect 7740 11088 7786 11134
rect 7858 11088 7904 11134
rect 7976 11088 8022 11134
rect 8094 11088 8140 11134
rect 20064 11225 20110 11271
rect 20168 11225 20214 11271
rect 20271 11225 20317 11271
rect 20374 11225 20420 11271
rect 20477 11225 20523 11271
rect 20580 11225 20626 11271
rect 20683 11225 20729 11271
rect 20786 11225 20832 11271
rect 20889 11225 20935 11271
rect 20992 11225 21038 11271
rect 3281 11001 3327 11047
rect 3384 11001 3430 11047
rect 3487 11001 3533 11047
rect 3590 11001 3636 11047
rect 3693 11001 3739 11047
rect 3796 11001 3842 11047
rect 3899 11001 3945 11047
rect 4002 11001 4048 11047
rect 4105 11001 4151 11047
rect 4209 11001 4255 11047
rect 9337 11001 9383 11047
rect 9459 11001 9505 11047
rect 9582 11001 9628 11047
rect 9705 11001 9751 11047
rect 3281 10777 3327 10823
rect 3384 10777 3430 10823
rect 3487 10777 3533 10823
rect 3590 10777 3636 10823
rect 3693 10777 3739 10823
rect 3796 10777 3842 10823
rect 3899 10777 3945 10823
rect 4002 10777 4048 10823
rect 4105 10777 4151 10823
rect 4209 10777 4255 10823
rect 9337 10777 9383 10823
rect 9459 10777 9505 10823
rect 9582 10777 9628 10823
rect 9705 10777 9751 10823
rect 20064 11001 20110 11047
rect 20168 11001 20214 11047
rect 20271 11001 20317 11047
rect 20374 11001 20420 11047
rect 20477 11001 20523 11047
rect 20580 11001 20626 11047
rect 20683 11001 20729 11047
rect 20786 11001 20832 11047
rect 20889 11001 20935 11047
rect 20992 11001 21038 11047
rect 3281 10553 3327 10599
rect 3384 10553 3430 10599
rect 3487 10553 3533 10599
rect 3590 10553 3636 10599
rect 3693 10553 3739 10599
rect 3796 10553 3842 10599
rect 3899 10553 3945 10599
rect 4002 10553 4048 10599
rect 4105 10553 4151 10599
rect 4209 10553 4255 10599
rect 9337 10553 9383 10599
rect 9459 10553 9505 10599
rect 9582 10553 9628 10599
rect 9705 10553 9751 10599
rect 20064 10777 20110 10823
rect 20168 10777 20214 10823
rect 20271 10777 20317 10823
rect 20374 10777 20420 10823
rect 20477 10777 20523 10823
rect 20580 10777 20626 10823
rect 20683 10777 20729 10823
rect 20786 10777 20832 10823
rect 20889 10777 20935 10823
rect 20992 10777 21038 10823
rect 20064 10553 20110 10599
rect 20168 10553 20214 10599
rect 20271 10553 20317 10599
rect 20374 10553 20420 10599
rect 20477 10553 20523 10599
rect 20580 10553 20626 10599
rect 20683 10553 20729 10599
rect 20786 10553 20832 10599
rect 20889 10553 20935 10599
rect 20992 10553 21038 10599
rect 7506 10466 7552 10512
rect 7623 10466 7669 10512
rect 7740 10466 7786 10512
rect 7858 10466 7904 10512
rect 7976 10466 8022 10512
rect 8094 10466 8140 10512
rect 3281 10329 3327 10375
rect 3384 10329 3430 10375
rect 3487 10329 3533 10375
rect 3590 10329 3636 10375
rect 3693 10329 3739 10375
rect 3796 10329 3842 10375
rect 3899 10329 3945 10375
rect 4002 10329 4048 10375
rect 4105 10329 4151 10375
rect 4209 10329 4255 10375
rect 7506 10242 7552 10288
rect 7623 10242 7669 10288
rect 7740 10242 7786 10288
rect 7858 10242 7904 10288
rect 7976 10242 8022 10288
rect 8094 10242 8140 10288
rect 9238 10242 9284 10288
rect 20064 10329 20110 10375
rect 20168 10329 20214 10375
rect 20271 10329 20317 10375
rect 20374 10329 20420 10375
rect 20477 10329 20523 10375
rect 20580 10329 20626 10375
rect 20683 10329 20729 10375
rect 20786 10329 20832 10375
rect 20889 10329 20935 10375
rect 20992 10329 21038 10375
rect 7506 10018 7552 10064
rect 7623 10018 7669 10064
rect 7740 10018 7786 10064
rect 7858 10018 7904 10064
rect 7976 10018 8022 10064
rect 8094 10018 8140 10064
rect 9238 10018 9284 10064
rect 7506 9736 7552 9782
rect 7623 9736 7669 9782
rect 7740 9736 7786 9782
rect 7858 9736 7904 9782
rect 7976 9736 8022 9782
rect 8094 9736 8140 9782
rect 9238 9736 9284 9782
rect 3281 9425 3327 9471
rect 3384 9425 3430 9471
rect 3487 9425 3533 9471
rect 3590 9425 3636 9471
rect 3693 9425 3739 9471
rect 3796 9425 3842 9471
rect 3899 9425 3945 9471
rect 4002 9425 4048 9471
rect 4105 9425 4151 9471
rect 4209 9425 4255 9471
rect 7506 9512 7552 9558
rect 7623 9512 7669 9558
rect 7740 9512 7786 9558
rect 7858 9512 7904 9558
rect 7976 9512 8022 9558
rect 8094 9512 8140 9558
rect 9238 9512 9284 9558
rect 7506 9288 7552 9334
rect 7623 9288 7669 9334
rect 7740 9288 7786 9334
rect 7858 9288 7904 9334
rect 7976 9288 8022 9334
rect 8094 9288 8140 9334
rect 20064 9425 20110 9471
rect 20168 9425 20214 9471
rect 20271 9425 20317 9471
rect 20374 9425 20420 9471
rect 20477 9425 20523 9471
rect 20580 9425 20626 9471
rect 20683 9425 20729 9471
rect 20786 9425 20832 9471
rect 20889 9425 20935 9471
rect 20992 9425 21038 9471
rect 3281 9201 3327 9247
rect 3384 9201 3430 9247
rect 3487 9201 3533 9247
rect 3590 9201 3636 9247
rect 3693 9201 3739 9247
rect 3796 9201 3842 9247
rect 3899 9201 3945 9247
rect 4002 9201 4048 9247
rect 4105 9201 4151 9247
rect 4209 9201 4255 9247
rect 9337 9201 9383 9247
rect 9459 9201 9505 9247
rect 9582 9201 9628 9247
rect 9705 9201 9751 9247
rect 3281 8977 3327 9023
rect 3384 8977 3430 9023
rect 3487 8977 3533 9023
rect 3590 8977 3636 9023
rect 3693 8977 3739 9023
rect 3796 8977 3842 9023
rect 3899 8977 3945 9023
rect 4002 8977 4048 9023
rect 4105 8977 4151 9023
rect 4209 8977 4255 9023
rect 9337 8977 9383 9023
rect 9459 8977 9505 9023
rect 9582 8977 9628 9023
rect 9705 8977 9751 9023
rect 20064 9201 20110 9247
rect 20168 9201 20214 9247
rect 20271 9201 20317 9247
rect 20374 9201 20420 9247
rect 20477 9201 20523 9247
rect 20580 9201 20626 9247
rect 20683 9201 20729 9247
rect 20786 9201 20832 9247
rect 20889 9201 20935 9247
rect 20992 9201 21038 9247
rect 3281 8753 3327 8799
rect 3384 8753 3430 8799
rect 3487 8753 3533 8799
rect 3590 8753 3636 8799
rect 3693 8753 3739 8799
rect 3796 8753 3842 8799
rect 3899 8753 3945 8799
rect 4002 8753 4048 8799
rect 4105 8753 4151 8799
rect 4209 8753 4255 8799
rect 9337 8753 9383 8799
rect 9459 8753 9505 8799
rect 9582 8753 9628 8799
rect 9705 8753 9751 8799
rect 20064 8977 20110 9023
rect 20168 8977 20214 9023
rect 20271 8977 20317 9023
rect 20374 8977 20420 9023
rect 20477 8977 20523 9023
rect 20580 8977 20626 9023
rect 20683 8977 20729 9023
rect 20786 8977 20832 9023
rect 20889 8977 20935 9023
rect 20992 8977 21038 9023
rect 20064 8753 20110 8799
rect 20168 8753 20214 8799
rect 20271 8753 20317 8799
rect 20374 8753 20420 8799
rect 20477 8753 20523 8799
rect 20580 8753 20626 8799
rect 20683 8753 20729 8799
rect 20786 8753 20832 8799
rect 20889 8753 20935 8799
rect 20992 8753 21038 8799
rect 7506 8666 7552 8712
rect 7623 8666 7669 8712
rect 7740 8666 7786 8712
rect 7858 8666 7904 8712
rect 7976 8666 8022 8712
rect 8094 8666 8140 8712
rect 3281 8529 3327 8575
rect 3384 8529 3430 8575
rect 3487 8529 3533 8575
rect 3590 8529 3636 8575
rect 3693 8529 3739 8575
rect 3796 8529 3842 8575
rect 3899 8529 3945 8575
rect 4002 8529 4048 8575
rect 4105 8529 4151 8575
rect 4209 8529 4255 8575
rect 7506 8442 7552 8488
rect 7623 8442 7669 8488
rect 7740 8442 7786 8488
rect 7858 8442 7904 8488
rect 7976 8442 8022 8488
rect 8094 8442 8140 8488
rect 9238 8442 9284 8488
rect 20064 8529 20110 8575
rect 20168 8529 20214 8575
rect 20271 8529 20317 8575
rect 20374 8529 20420 8575
rect 20477 8529 20523 8575
rect 20580 8529 20626 8575
rect 20683 8529 20729 8575
rect 20786 8529 20832 8575
rect 20889 8529 20935 8575
rect 20992 8529 21038 8575
rect 7506 8218 7552 8264
rect 7623 8218 7669 8264
rect 7740 8218 7786 8264
rect 7858 8218 7904 8264
rect 7976 8218 8022 8264
rect 8094 8218 8140 8264
rect 9238 8218 9284 8264
rect 7506 7936 7552 7982
rect 7623 7936 7669 7982
rect 7740 7936 7786 7982
rect 7858 7936 7904 7982
rect 7976 7936 8022 7982
rect 8094 7936 8140 7982
rect 9238 7936 9284 7982
rect 3281 7625 3327 7671
rect 3384 7625 3430 7671
rect 3487 7625 3533 7671
rect 3590 7625 3636 7671
rect 3693 7625 3739 7671
rect 3796 7625 3842 7671
rect 3899 7625 3945 7671
rect 4002 7625 4048 7671
rect 4105 7625 4151 7671
rect 4209 7625 4255 7671
rect 7506 7712 7552 7758
rect 7623 7712 7669 7758
rect 7740 7712 7786 7758
rect 7858 7712 7904 7758
rect 7976 7712 8022 7758
rect 8094 7712 8140 7758
rect 9238 7712 9284 7758
rect 7506 7488 7552 7534
rect 7623 7488 7669 7534
rect 7740 7488 7786 7534
rect 7858 7488 7904 7534
rect 7976 7488 8022 7534
rect 8094 7488 8140 7534
rect 20064 7625 20110 7671
rect 20168 7625 20214 7671
rect 20271 7625 20317 7671
rect 20374 7625 20420 7671
rect 20477 7625 20523 7671
rect 20580 7625 20626 7671
rect 20683 7625 20729 7671
rect 20786 7625 20832 7671
rect 20889 7625 20935 7671
rect 20992 7625 21038 7671
rect 3281 7401 3327 7447
rect 3384 7401 3430 7447
rect 3487 7401 3533 7447
rect 3590 7401 3636 7447
rect 3693 7401 3739 7447
rect 3796 7401 3842 7447
rect 3899 7401 3945 7447
rect 4002 7401 4048 7447
rect 4105 7401 4151 7447
rect 4209 7401 4255 7447
rect 9337 7401 9383 7447
rect 9459 7401 9505 7447
rect 9582 7401 9628 7447
rect 9705 7401 9751 7447
rect 3281 7177 3327 7223
rect 3384 7177 3430 7223
rect 3487 7177 3533 7223
rect 3590 7177 3636 7223
rect 3693 7177 3739 7223
rect 3796 7177 3842 7223
rect 3899 7177 3945 7223
rect 4002 7177 4048 7223
rect 4105 7177 4151 7223
rect 4209 7177 4255 7223
rect 9337 7177 9383 7223
rect 9459 7177 9505 7223
rect 9582 7177 9628 7223
rect 9705 7177 9751 7223
rect 20064 7401 20110 7447
rect 20168 7401 20214 7447
rect 20271 7401 20317 7447
rect 20374 7401 20420 7447
rect 20477 7401 20523 7447
rect 20580 7401 20626 7447
rect 20683 7401 20729 7447
rect 20786 7401 20832 7447
rect 20889 7401 20935 7447
rect 20992 7401 21038 7447
rect 3281 6953 3327 6999
rect 3384 6953 3430 6999
rect 3487 6953 3533 6999
rect 3590 6953 3636 6999
rect 3693 6953 3739 6999
rect 3796 6953 3842 6999
rect 3899 6953 3945 6999
rect 4002 6953 4048 6999
rect 4105 6953 4151 6999
rect 4209 6953 4255 6999
rect 9337 6953 9383 6999
rect 9459 6953 9505 6999
rect 9582 6953 9628 6999
rect 9705 6953 9751 6999
rect 20064 7177 20110 7223
rect 20168 7177 20214 7223
rect 20271 7177 20317 7223
rect 20374 7177 20420 7223
rect 20477 7177 20523 7223
rect 20580 7177 20626 7223
rect 20683 7177 20729 7223
rect 20786 7177 20832 7223
rect 20889 7177 20935 7223
rect 20992 7177 21038 7223
rect 20064 6953 20110 6999
rect 20168 6953 20214 6999
rect 20271 6953 20317 6999
rect 20374 6953 20420 6999
rect 20477 6953 20523 6999
rect 20580 6953 20626 6999
rect 20683 6953 20729 6999
rect 20786 6953 20832 6999
rect 20889 6953 20935 6999
rect 20992 6953 21038 6999
rect 7506 6866 7552 6912
rect 7623 6866 7669 6912
rect 7740 6866 7786 6912
rect 7858 6866 7904 6912
rect 7976 6866 8022 6912
rect 8094 6866 8140 6912
rect 3281 6729 3327 6775
rect 3384 6729 3430 6775
rect 3487 6729 3533 6775
rect 3590 6729 3636 6775
rect 3693 6729 3739 6775
rect 3796 6729 3842 6775
rect 3899 6729 3945 6775
rect 4002 6729 4048 6775
rect 4105 6729 4151 6775
rect 4209 6729 4255 6775
rect 7506 6642 7552 6688
rect 7623 6642 7669 6688
rect 7740 6642 7786 6688
rect 7858 6642 7904 6688
rect 7976 6642 8022 6688
rect 8094 6642 8140 6688
rect 9238 6642 9284 6688
rect 20064 6729 20110 6775
rect 20168 6729 20214 6775
rect 20271 6729 20317 6775
rect 20374 6729 20420 6775
rect 20477 6729 20523 6775
rect 20580 6729 20626 6775
rect 20683 6729 20729 6775
rect 20786 6729 20832 6775
rect 20889 6729 20935 6775
rect 20992 6729 21038 6775
rect 7506 6418 7552 6464
rect 7623 6418 7669 6464
rect 7740 6418 7786 6464
rect 7858 6418 7904 6464
rect 7976 6418 8022 6464
rect 8094 6418 8140 6464
rect 9238 6418 9284 6464
rect 7506 6136 7552 6182
rect 7623 6136 7669 6182
rect 7740 6136 7786 6182
rect 7858 6136 7904 6182
rect 7976 6136 8022 6182
rect 8094 6136 8140 6182
rect 9238 6136 9284 6182
rect 3281 5825 3327 5871
rect 3384 5825 3430 5871
rect 3487 5825 3533 5871
rect 3590 5825 3636 5871
rect 3693 5825 3739 5871
rect 3796 5825 3842 5871
rect 3899 5825 3945 5871
rect 4002 5825 4048 5871
rect 4105 5825 4151 5871
rect 4209 5825 4255 5871
rect 7506 5912 7552 5958
rect 7623 5912 7669 5958
rect 7740 5912 7786 5958
rect 7858 5912 7904 5958
rect 7976 5912 8022 5958
rect 8094 5912 8140 5958
rect 9238 5912 9284 5958
rect 7506 5688 7552 5734
rect 7623 5688 7669 5734
rect 7740 5688 7786 5734
rect 7858 5688 7904 5734
rect 7976 5688 8022 5734
rect 8094 5688 8140 5734
rect 20064 5825 20110 5871
rect 20168 5825 20214 5871
rect 20271 5825 20317 5871
rect 20374 5825 20420 5871
rect 20477 5825 20523 5871
rect 20580 5825 20626 5871
rect 20683 5825 20729 5871
rect 20786 5825 20832 5871
rect 20889 5825 20935 5871
rect 20992 5825 21038 5871
rect 3281 5601 3327 5647
rect 3384 5601 3430 5647
rect 3487 5601 3533 5647
rect 3590 5601 3636 5647
rect 3693 5601 3739 5647
rect 3796 5601 3842 5647
rect 3899 5601 3945 5647
rect 4002 5601 4048 5647
rect 4105 5601 4151 5647
rect 4209 5601 4255 5647
rect 9337 5601 9383 5647
rect 9459 5601 9505 5647
rect 9582 5601 9628 5647
rect 9705 5601 9751 5647
rect 3281 5377 3327 5423
rect 3384 5377 3430 5423
rect 3487 5377 3533 5423
rect 3590 5377 3636 5423
rect 3693 5377 3739 5423
rect 3796 5377 3842 5423
rect 3899 5377 3945 5423
rect 4002 5377 4048 5423
rect 4105 5377 4151 5423
rect 4209 5377 4255 5423
rect 9337 5377 9383 5423
rect 9459 5377 9505 5423
rect 9582 5377 9628 5423
rect 9705 5377 9751 5423
rect 20064 5601 20110 5647
rect 20168 5601 20214 5647
rect 20271 5601 20317 5647
rect 20374 5601 20420 5647
rect 20477 5601 20523 5647
rect 20580 5601 20626 5647
rect 20683 5601 20729 5647
rect 20786 5601 20832 5647
rect 20889 5601 20935 5647
rect 20992 5601 21038 5647
rect 3281 5153 3327 5199
rect 3384 5153 3430 5199
rect 3487 5153 3533 5199
rect 3590 5153 3636 5199
rect 3693 5153 3739 5199
rect 3796 5153 3842 5199
rect 3899 5153 3945 5199
rect 4002 5153 4048 5199
rect 4105 5153 4151 5199
rect 4209 5153 4255 5199
rect 9337 5153 9383 5199
rect 9459 5153 9505 5199
rect 9582 5153 9628 5199
rect 9705 5153 9751 5199
rect 20064 5377 20110 5423
rect 20168 5377 20214 5423
rect 20271 5377 20317 5423
rect 20374 5377 20420 5423
rect 20477 5377 20523 5423
rect 20580 5377 20626 5423
rect 20683 5377 20729 5423
rect 20786 5377 20832 5423
rect 20889 5377 20935 5423
rect 20992 5377 21038 5423
rect 20064 5153 20110 5199
rect 20168 5153 20214 5199
rect 20271 5153 20317 5199
rect 20374 5153 20420 5199
rect 20477 5153 20523 5199
rect 20580 5153 20626 5199
rect 20683 5153 20729 5199
rect 20786 5153 20832 5199
rect 20889 5153 20935 5199
rect 20992 5153 21038 5199
rect 7506 5066 7552 5112
rect 7623 5066 7669 5112
rect 7740 5066 7786 5112
rect 7858 5066 7904 5112
rect 7976 5066 8022 5112
rect 8094 5066 8140 5112
rect 3281 4929 3327 4975
rect 3384 4929 3430 4975
rect 3487 4929 3533 4975
rect 3590 4929 3636 4975
rect 3693 4929 3739 4975
rect 3796 4929 3842 4975
rect 3899 4929 3945 4975
rect 4002 4929 4048 4975
rect 4105 4929 4151 4975
rect 4209 4929 4255 4975
rect 7506 4842 7552 4888
rect 7623 4842 7669 4888
rect 7740 4842 7786 4888
rect 7858 4842 7904 4888
rect 7976 4842 8022 4888
rect 8094 4842 8140 4888
rect 9238 4842 9284 4888
rect 20064 4929 20110 4975
rect 20168 4929 20214 4975
rect 20271 4929 20317 4975
rect 20374 4929 20420 4975
rect 20477 4929 20523 4975
rect 20580 4929 20626 4975
rect 20683 4929 20729 4975
rect 20786 4929 20832 4975
rect 20889 4929 20935 4975
rect 20992 4929 21038 4975
rect 7506 4618 7552 4664
rect 7623 4618 7669 4664
rect 7740 4618 7786 4664
rect 7858 4618 7904 4664
rect 7976 4618 8022 4664
rect 8094 4618 8140 4664
rect 9238 4618 9284 4664
rect 7506 4336 7552 4382
rect 7623 4336 7669 4382
rect 7740 4336 7786 4382
rect 7858 4336 7904 4382
rect 7976 4336 8022 4382
rect 8094 4336 8140 4382
rect 9238 4336 9284 4382
rect 3281 4025 3327 4071
rect 3384 4025 3430 4071
rect 3487 4025 3533 4071
rect 3590 4025 3636 4071
rect 3693 4025 3739 4071
rect 3796 4025 3842 4071
rect 3899 4025 3945 4071
rect 4002 4025 4048 4071
rect 4105 4025 4151 4071
rect 4209 4025 4255 4071
rect 7506 4112 7552 4158
rect 7623 4112 7669 4158
rect 7740 4112 7786 4158
rect 7858 4112 7904 4158
rect 7976 4112 8022 4158
rect 8094 4112 8140 4158
rect 9238 4112 9284 4158
rect 7506 3888 7552 3934
rect 7623 3888 7669 3934
rect 7740 3888 7786 3934
rect 7858 3888 7904 3934
rect 7976 3888 8022 3934
rect 8094 3888 8140 3934
rect 20064 4025 20110 4071
rect 20168 4025 20214 4071
rect 20271 4025 20317 4071
rect 20374 4025 20420 4071
rect 20477 4025 20523 4071
rect 20580 4025 20626 4071
rect 20683 4025 20729 4071
rect 20786 4025 20832 4071
rect 20889 4025 20935 4071
rect 20992 4025 21038 4071
rect 3281 3801 3327 3847
rect 3384 3801 3430 3847
rect 3487 3801 3533 3847
rect 3590 3801 3636 3847
rect 3693 3801 3739 3847
rect 3796 3801 3842 3847
rect 3899 3801 3945 3847
rect 4002 3801 4048 3847
rect 4105 3801 4151 3847
rect 4209 3801 4255 3847
rect 9337 3801 9383 3847
rect 9459 3801 9505 3847
rect 9582 3801 9628 3847
rect 9705 3801 9751 3847
rect 3281 3577 3327 3623
rect 3384 3577 3430 3623
rect 3487 3577 3533 3623
rect 3590 3577 3636 3623
rect 3693 3577 3739 3623
rect 3796 3577 3842 3623
rect 3899 3577 3945 3623
rect 4002 3577 4048 3623
rect 4105 3577 4151 3623
rect 4209 3577 4255 3623
rect 9337 3577 9383 3623
rect 9459 3577 9505 3623
rect 9582 3577 9628 3623
rect 9705 3577 9751 3623
rect 20064 3801 20110 3847
rect 20168 3801 20214 3847
rect 20271 3801 20317 3847
rect 20374 3801 20420 3847
rect 20477 3801 20523 3847
rect 20580 3801 20626 3847
rect 20683 3801 20729 3847
rect 20786 3801 20832 3847
rect 20889 3801 20935 3847
rect 20992 3801 21038 3847
rect 3281 3353 3327 3399
rect 3384 3353 3430 3399
rect 3487 3353 3533 3399
rect 3590 3353 3636 3399
rect 3693 3353 3739 3399
rect 3796 3353 3842 3399
rect 3899 3353 3945 3399
rect 4002 3353 4048 3399
rect 4105 3353 4151 3399
rect 4209 3353 4255 3399
rect 9337 3353 9383 3399
rect 9459 3353 9505 3399
rect 9582 3353 9628 3399
rect 9705 3353 9751 3399
rect 20064 3577 20110 3623
rect 20168 3577 20214 3623
rect 20271 3577 20317 3623
rect 20374 3577 20420 3623
rect 20477 3577 20523 3623
rect 20580 3577 20626 3623
rect 20683 3577 20729 3623
rect 20786 3577 20832 3623
rect 20889 3577 20935 3623
rect 20992 3577 21038 3623
rect 20064 3353 20110 3399
rect 20168 3353 20214 3399
rect 20271 3353 20317 3399
rect 20374 3353 20420 3399
rect 20477 3353 20523 3399
rect 20580 3353 20626 3399
rect 20683 3353 20729 3399
rect 20786 3353 20832 3399
rect 20889 3353 20935 3399
rect 20992 3353 21038 3399
rect 7506 3266 7552 3312
rect 7623 3266 7669 3312
rect 7740 3266 7786 3312
rect 7858 3266 7904 3312
rect 7976 3266 8022 3312
rect 8094 3266 8140 3312
rect 3281 3129 3327 3175
rect 3384 3129 3430 3175
rect 3487 3129 3533 3175
rect 3590 3129 3636 3175
rect 3693 3129 3739 3175
rect 3796 3129 3842 3175
rect 3899 3129 3945 3175
rect 4002 3129 4048 3175
rect 4105 3129 4151 3175
rect 4209 3129 4255 3175
rect 7506 3042 7552 3088
rect 7623 3042 7669 3088
rect 7740 3042 7786 3088
rect 7858 3042 7904 3088
rect 7976 3042 8022 3088
rect 8094 3042 8140 3088
rect 9238 3042 9284 3088
rect 20064 3129 20110 3175
rect 20168 3129 20214 3175
rect 20271 3129 20317 3175
rect 20374 3129 20420 3175
rect 20477 3129 20523 3175
rect 20580 3129 20626 3175
rect 20683 3129 20729 3175
rect 20786 3129 20832 3175
rect 20889 3129 20935 3175
rect 20992 3129 21038 3175
rect 7506 2818 7552 2864
rect 7623 2818 7669 2864
rect 7740 2818 7786 2864
rect 7858 2818 7904 2864
rect 7976 2818 8022 2864
rect 8094 2818 8140 2864
rect 9238 2818 9284 2864
rect 7506 2536 7552 2582
rect 7623 2536 7669 2582
rect 7740 2536 7786 2582
rect 7858 2536 7904 2582
rect 7976 2536 8022 2582
rect 8094 2536 8140 2582
rect 9238 2536 9284 2582
rect 3281 2225 3327 2271
rect 3384 2225 3430 2271
rect 3487 2225 3533 2271
rect 3590 2225 3636 2271
rect 3693 2225 3739 2271
rect 3796 2225 3842 2271
rect 3899 2225 3945 2271
rect 4002 2225 4048 2271
rect 4105 2225 4151 2271
rect 4209 2225 4255 2271
rect 7506 2312 7552 2358
rect 7623 2312 7669 2358
rect 7740 2312 7786 2358
rect 7858 2312 7904 2358
rect 7976 2312 8022 2358
rect 8094 2312 8140 2358
rect 9238 2312 9284 2358
rect 7506 2088 7552 2134
rect 7623 2088 7669 2134
rect 7740 2088 7786 2134
rect 7858 2088 7904 2134
rect 7976 2088 8022 2134
rect 8094 2088 8140 2134
rect 20064 2225 20110 2271
rect 20168 2225 20214 2271
rect 20271 2225 20317 2271
rect 20374 2225 20420 2271
rect 20477 2225 20523 2271
rect 20580 2225 20626 2271
rect 20683 2225 20729 2271
rect 20786 2225 20832 2271
rect 20889 2225 20935 2271
rect 20992 2225 21038 2271
rect 3281 2001 3327 2047
rect 3384 2001 3430 2047
rect 3487 2001 3533 2047
rect 3590 2001 3636 2047
rect 3693 2001 3739 2047
rect 3796 2001 3842 2047
rect 3899 2001 3945 2047
rect 4002 2001 4048 2047
rect 4105 2001 4151 2047
rect 4209 2001 4255 2047
rect 9337 2001 9383 2047
rect 9459 2001 9505 2047
rect 9582 2001 9628 2047
rect 9705 2001 9751 2047
rect 3281 1777 3327 1823
rect 3384 1777 3430 1823
rect 3487 1777 3533 1823
rect 3590 1777 3636 1823
rect 3693 1777 3739 1823
rect 3796 1777 3842 1823
rect 3899 1777 3945 1823
rect 4002 1777 4048 1823
rect 4105 1777 4151 1823
rect 4209 1777 4255 1823
rect 9337 1777 9383 1823
rect 9459 1777 9505 1823
rect 9582 1777 9628 1823
rect 9705 1777 9751 1823
rect 20064 2001 20110 2047
rect 20168 2001 20214 2047
rect 20271 2001 20317 2047
rect 20374 2001 20420 2047
rect 20477 2001 20523 2047
rect 20580 2001 20626 2047
rect 20683 2001 20729 2047
rect 20786 2001 20832 2047
rect 20889 2001 20935 2047
rect 20992 2001 21038 2047
rect 3281 1553 3327 1599
rect 3384 1553 3430 1599
rect 3487 1553 3533 1599
rect 3590 1553 3636 1599
rect 3693 1553 3739 1599
rect 3796 1553 3842 1599
rect 3899 1553 3945 1599
rect 4002 1553 4048 1599
rect 4105 1553 4151 1599
rect 4209 1553 4255 1599
rect 9337 1553 9383 1599
rect 9459 1553 9505 1599
rect 9582 1553 9628 1599
rect 9705 1553 9751 1599
rect 20064 1777 20110 1823
rect 20168 1777 20214 1823
rect 20271 1777 20317 1823
rect 20374 1777 20420 1823
rect 20477 1777 20523 1823
rect 20580 1777 20626 1823
rect 20683 1777 20729 1823
rect 20786 1777 20832 1823
rect 20889 1777 20935 1823
rect 20992 1777 21038 1823
rect 20064 1553 20110 1599
rect 20168 1553 20214 1599
rect 20271 1553 20317 1599
rect 20374 1553 20420 1599
rect 20477 1553 20523 1599
rect 20580 1553 20626 1599
rect 20683 1553 20729 1599
rect 20786 1553 20832 1599
rect 20889 1553 20935 1599
rect 20992 1553 21038 1599
rect 7506 1466 7552 1512
rect 7623 1466 7669 1512
rect 7740 1466 7786 1512
rect 7858 1466 7904 1512
rect 7976 1466 8022 1512
rect 8094 1466 8140 1512
rect 3281 1329 3327 1375
rect 3384 1329 3430 1375
rect 3487 1329 3533 1375
rect 3590 1329 3636 1375
rect 3693 1329 3739 1375
rect 3796 1329 3842 1375
rect 3899 1329 3945 1375
rect 4002 1329 4048 1375
rect 4105 1329 4151 1375
rect 4209 1329 4255 1375
rect 7506 1242 7552 1288
rect 7623 1242 7669 1288
rect 7740 1242 7786 1288
rect 7858 1242 7904 1288
rect 7976 1242 8022 1288
rect 8094 1242 8140 1288
rect 9238 1242 9284 1288
rect 20064 1329 20110 1375
rect 20168 1329 20214 1375
rect 20271 1329 20317 1375
rect 20374 1329 20420 1375
rect 20477 1329 20523 1375
rect 20580 1329 20626 1375
rect 20683 1329 20729 1375
rect 20786 1329 20832 1375
rect 20889 1329 20935 1375
rect 20992 1329 21038 1375
rect 7506 1018 7552 1064
rect 7623 1018 7669 1064
rect 7740 1018 7786 1064
rect 7858 1018 7904 1064
rect 7976 1018 8022 1064
rect 8094 1018 8140 1064
rect 9238 1018 9284 1064
rect 7506 736 7552 782
rect 7623 736 7669 782
rect 7740 736 7786 782
rect 7858 736 7904 782
rect 7976 736 8022 782
rect 8094 736 8140 782
rect 9238 736 9284 782
rect 3281 425 3327 471
rect 3384 425 3430 471
rect 3487 425 3533 471
rect 3590 425 3636 471
rect 3693 425 3739 471
rect 3796 425 3842 471
rect 3899 425 3945 471
rect 4002 425 4048 471
rect 4105 425 4151 471
rect 4209 425 4255 471
rect 7506 512 7552 558
rect 7623 512 7669 558
rect 7740 512 7786 558
rect 7858 512 7904 558
rect 7976 512 8022 558
rect 8094 512 8140 558
rect 9238 512 9284 558
rect 7506 288 7552 334
rect 7623 288 7669 334
rect 7740 288 7786 334
rect 7858 288 7904 334
rect 7976 288 8022 334
rect 8094 288 8140 334
rect 20064 425 20110 471
rect 20168 425 20214 471
rect 20271 425 20317 471
rect 20374 425 20420 471
rect 20477 425 20523 471
rect 20580 425 20626 471
rect 20683 425 20729 471
rect 20786 425 20832 471
rect 20889 425 20935 471
rect 20992 425 21038 471
rect 3281 201 3327 247
rect 3384 201 3430 247
rect 3487 201 3533 247
rect 3590 201 3636 247
rect 3693 201 3739 247
rect 3796 201 3842 247
rect 3899 201 3945 247
rect 4002 201 4048 247
rect 4105 201 4151 247
rect 4209 201 4255 247
rect 9337 201 9383 247
rect 9459 201 9505 247
rect 9582 201 9628 247
rect 9705 201 9751 247
rect 3281 -23 3327 23
rect 3384 -23 3430 23
rect 3487 -23 3533 23
rect 3590 -23 3636 23
rect 3693 -23 3739 23
rect 3796 -23 3842 23
rect 3899 -23 3945 23
rect 4002 -23 4048 23
rect 4105 -23 4151 23
rect 4209 -23 4255 23
rect 9337 -23 9383 23
rect 9459 -23 9505 23
rect 9582 -23 9628 23
rect 9705 -23 9751 23
rect 20064 201 20110 247
rect 20168 201 20214 247
rect 20271 201 20317 247
rect 20374 201 20420 247
rect 20477 201 20523 247
rect 20580 201 20626 247
rect 20683 201 20729 247
rect 20786 201 20832 247
rect 20889 201 20935 247
rect 20992 201 21038 247
rect 20064 -23 20110 23
rect 20168 -23 20214 23
rect 20271 -23 20317 23
rect 20374 -23 20420 23
rect 20477 -23 20523 23
rect 20580 -23 20626 23
rect 20683 -23 20729 23
rect 20786 -23 20832 23
rect 20889 -23 20935 23
rect 20992 -23 21038 23
<< mvpdiffc >>
rect 946 14377 2920 14423
rect 946 14153 2920 14199
rect 946 13929 2920 13975
rect 14409 14377 14455 14423
rect 14522 14377 14568 14423
rect 14635 14377 14681 14423
rect 14748 14377 14794 14423
rect 14861 14377 14907 14423
rect 21399 14377 23373 14423
rect 4870 14066 5120 14112
rect 5177 14066 5223 14112
rect 5280 14066 5326 14112
rect 5383 14066 5429 14112
rect 5486 14066 5532 14112
rect 5589 14066 5635 14112
rect 5692 14066 5738 14112
rect 5795 14066 5841 14112
rect 5898 14066 5944 14112
rect 6451 14066 6497 14112
rect 6568 14066 6614 14112
rect 6685 14066 6731 14112
rect 6803 14066 6849 14112
rect 6921 14066 6967 14112
rect 7039 14066 7085 14112
rect 14409 14153 14455 14199
rect 14522 14153 14568 14199
rect 14635 14153 14681 14199
rect 14748 14153 14794 14199
rect 14861 14153 14907 14199
rect 946 13705 2920 13751
rect 4870 13842 5120 13888
rect 5177 13842 5223 13888
rect 5280 13842 5326 13888
rect 5383 13842 5429 13888
rect 5486 13842 5532 13888
rect 5589 13842 5635 13888
rect 5692 13842 5738 13888
rect 5795 13842 5841 13888
rect 5898 13842 5944 13888
rect 18375 14066 18421 14112
rect 18478 14066 18524 14112
rect 18581 14066 18627 14112
rect 18684 14066 18730 14112
rect 18787 14066 18833 14112
rect 18890 14066 18936 14112
rect 18993 14066 19039 14112
rect 19096 14066 19142 14112
rect 19199 14066 19449 14112
rect 6451 13842 6497 13888
rect 6568 13842 6614 13888
rect 6685 13842 6731 13888
rect 6803 13842 6849 13888
rect 6921 13842 6967 13888
rect 7039 13842 7085 13888
rect 8618 13842 8664 13888
rect 8741 13842 8787 13888
rect 8864 13842 8910 13888
rect 14409 13929 14455 13975
rect 14522 13929 14568 13975
rect 14635 13929 14681 13975
rect 14748 13929 14794 13975
rect 14861 13929 14907 13975
rect 18375 13842 18421 13888
rect 18478 13842 18524 13888
rect 18581 13842 18627 13888
rect 18684 13842 18730 13888
rect 18787 13842 18833 13888
rect 18890 13842 18936 13888
rect 18993 13842 19039 13888
rect 19096 13842 19142 13888
rect 19199 13842 19449 13888
rect 4870 13618 5120 13664
rect 5177 13618 5223 13664
rect 5280 13618 5326 13664
rect 5383 13618 5429 13664
rect 5486 13618 5532 13664
rect 5589 13618 5635 13664
rect 5692 13618 5738 13664
rect 5795 13618 5841 13664
rect 5898 13618 5944 13664
rect 6451 13618 6497 13664
rect 6568 13618 6614 13664
rect 6685 13618 6731 13664
rect 6803 13618 6849 13664
rect 6921 13618 6967 13664
rect 7039 13618 7085 13664
rect 8618 13618 8664 13664
rect 8741 13618 8787 13664
rect 8864 13618 8910 13664
rect 14409 13705 14455 13751
rect 14522 13705 14568 13751
rect 14635 13705 14681 13751
rect 14748 13705 14794 13751
rect 14861 13705 14907 13751
rect 21399 14153 23373 14199
rect 21399 13929 23373 13975
rect 18375 13618 18421 13664
rect 18478 13618 18524 13664
rect 18581 13618 18627 13664
rect 18684 13618 18730 13664
rect 18787 13618 18833 13664
rect 18890 13618 18936 13664
rect 18993 13618 19039 13664
rect 19096 13618 19142 13664
rect 19199 13618 19449 13664
rect 21399 13705 23373 13751
rect 946 13249 2920 13295
rect 4870 13336 5120 13382
rect 5177 13336 5223 13382
rect 5280 13336 5326 13382
rect 5383 13336 5429 13382
rect 5486 13336 5532 13382
rect 5589 13336 5635 13382
rect 5692 13336 5738 13382
rect 5795 13336 5841 13382
rect 5898 13336 5944 13382
rect 6451 13336 6497 13382
rect 6568 13336 6614 13382
rect 6685 13336 6731 13382
rect 6803 13336 6849 13382
rect 6921 13336 6967 13382
rect 7039 13336 7085 13382
rect 8618 13336 8664 13382
rect 8741 13336 8787 13382
rect 8864 13336 8910 13382
rect 946 13025 2920 13071
rect 946 12801 2920 12847
rect 4870 13112 5120 13158
rect 5177 13112 5223 13158
rect 5280 13112 5326 13158
rect 5383 13112 5429 13158
rect 5486 13112 5532 13158
rect 5589 13112 5635 13158
rect 5692 13112 5738 13158
rect 5795 13112 5841 13158
rect 5898 13112 5944 13158
rect 6451 13112 6497 13158
rect 6568 13112 6614 13158
rect 6685 13112 6731 13158
rect 6803 13112 6849 13158
rect 6921 13112 6967 13158
rect 7039 13112 7085 13158
rect 18375 13336 18421 13382
rect 18478 13336 18524 13382
rect 18581 13336 18627 13382
rect 18684 13336 18730 13382
rect 18787 13336 18833 13382
rect 18890 13336 18936 13382
rect 18993 13336 19039 13382
rect 19096 13336 19142 13382
rect 19199 13336 19449 13382
rect 14409 13249 14455 13295
rect 14522 13249 14568 13295
rect 14635 13249 14681 13295
rect 14748 13249 14794 13295
rect 14861 13249 14907 13295
rect 8618 13112 8664 13158
rect 8741 13112 8787 13158
rect 8864 13112 8910 13158
rect 14409 13025 14455 13071
rect 14522 13025 14568 13071
rect 14635 13025 14681 13071
rect 14748 13025 14794 13071
rect 14861 13025 14907 13071
rect 18375 13112 18421 13158
rect 18478 13112 18524 13158
rect 18581 13112 18627 13158
rect 18684 13112 18730 13158
rect 18787 13112 18833 13158
rect 18890 13112 18936 13158
rect 18993 13112 19039 13158
rect 19096 13112 19142 13158
rect 19199 13112 19449 13158
rect 21399 13249 23373 13295
rect 4870 12888 5120 12934
rect 5177 12888 5223 12934
rect 5280 12888 5326 12934
rect 5383 12888 5429 12934
rect 5486 12888 5532 12934
rect 5589 12888 5635 12934
rect 5692 12888 5738 12934
rect 5795 12888 5841 12934
rect 5898 12888 5944 12934
rect 6451 12888 6497 12934
rect 6568 12888 6614 12934
rect 6685 12888 6731 12934
rect 6803 12888 6849 12934
rect 6921 12888 6967 12934
rect 7039 12888 7085 12934
rect 18375 12888 18421 12934
rect 18478 12888 18524 12934
rect 18581 12888 18627 12934
rect 18684 12888 18730 12934
rect 18787 12888 18833 12934
rect 18890 12888 18936 12934
rect 18993 12888 19039 12934
rect 19096 12888 19142 12934
rect 19199 12888 19449 12934
rect 14409 12801 14455 12847
rect 14522 12801 14568 12847
rect 14635 12801 14681 12847
rect 14748 12801 14794 12847
rect 14861 12801 14907 12847
rect 946 12577 2920 12623
rect 946 12353 2920 12399
rect 946 12129 2920 12175
rect 21399 13025 23373 13071
rect 21399 12801 23373 12847
rect 14409 12577 14455 12623
rect 14522 12577 14568 12623
rect 14635 12577 14681 12623
rect 14748 12577 14794 12623
rect 14861 12577 14907 12623
rect 21399 12577 23373 12623
rect 4870 12266 5120 12312
rect 5177 12266 5223 12312
rect 5280 12266 5326 12312
rect 5383 12266 5429 12312
rect 5486 12266 5532 12312
rect 5589 12266 5635 12312
rect 5692 12266 5738 12312
rect 5795 12266 5841 12312
rect 5898 12266 5944 12312
rect 6451 12266 6497 12312
rect 6568 12266 6614 12312
rect 6685 12266 6731 12312
rect 6803 12266 6849 12312
rect 6921 12266 6967 12312
rect 7039 12266 7085 12312
rect 14409 12353 14455 12399
rect 14522 12353 14568 12399
rect 14635 12353 14681 12399
rect 14748 12353 14794 12399
rect 14861 12353 14907 12399
rect 946 11905 2920 11951
rect 4870 12042 5120 12088
rect 5177 12042 5223 12088
rect 5280 12042 5326 12088
rect 5383 12042 5429 12088
rect 5486 12042 5532 12088
rect 5589 12042 5635 12088
rect 5692 12042 5738 12088
rect 5795 12042 5841 12088
rect 5898 12042 5944 12088
rect 18375 12266 18421 12312
rect 18478 12266 18524 12312
rect 18581 12266 18627 12312
rect 18684 12266 18730 12312
rect 18787 12266 18833 12312
rect 18890 12266 18936 12312
rect 18993 12266 19039 12312
rect 19096 12266 19142 12312
rect 19199 12266 19449 12312
rect 6451 12042 6497 12088
rect 6568 12042 6614 12088
rect 6685 12042 6731 12088
rect 6803 12042 6849 12088
rect 6921 12042 6967 12088
rect 7039 12042 7085 12088
rect 8618 12042 8664 12088
rect 8741 12042 8787 12088
rect 8864 12042 8910 12088
rect 14409 12129 14455 12175
rect 14522 12129 14568 12175
rect 14635 12129 14681 12175
rect 14748 12129 14794 12175
rect 14861 12129 14907 12175
rect 18375 12042 18421 12088
rect 18478 12042 18524 12088
rect 18581 12042 18627 12088
rect 18684 12042 18730 12088
rect 18787 12042 18833 12088
rect 18890 12042 18936 12088
rect 18993 12042 19039 12088
rect 19096 12042 19142 12088
rect 19199 12042 19449 12088
rect 4870 11818 5120 11864
rect 5177 11818 5223 11864
rect 5280 11818 5326 11864
rect 5383 11818 5429 11864
rect 5486 11818 5532 11864
rect 5589 11818 5635 11864
rect 5692 11818 5738 11864
rect 5795 11818 5841 11864
rect 5898 11818 5944 11864
rect 6451 11818 6497 11864
rect 6568 11818 6614 11864
rect 6685 11818 6731 11864
rect 6803 11818 6849 11864
rect 6921 11818 6967 11864
rect 7039 11818 7085 11864
rect 8618 11818 8664 11864
rect 8741 11818 8787 11864
rect 8864 11818 8910 11864
rect 14409 11905 14455 11951
rect 14522 11905 14568 11951
rect 14635 11905 14681 11951
rect 14748 11905 14794 11951
rect 14861 11905 14907 11951
rect 21399 12353 23373 12399
rect 21399 12129 23373 12175
rect 18375 11818 18421 11864
rect 18478 11818 18524 11864
rect 18581 11818 18627 11864
rect 18684 11818 18730 11864
rect 18787 11818 18833 11864
rect 18890 11818 18936 11864
rect 18993 11818 19039 11864
rect 19096 11818 19142 11864
rect 19199 11818 19449 11864
rect 21399 11905 23373 11951
rect 946 11449 2920 11495
rect 4870 11536 5120 11582
rect 5177 11536 5223 11582
rect 5280 11536 5326 11582
rect 5383 11536 5429 11582
rect 5486 11536 5532 11582
rect 5589 11536 5635 11582
rect 5692 11536 5738 11582
rect 5795 11536 5841 11582
rect 5898 11536 5944 11582
rect 6451 11536 6497 11582
rect 6568 11536 6614 11582
rect 6685 11536 6731 11582
rect 6803 11536 6849 11582
rect 6921 11536 6967 11582
rect 7039 11536 7085 11582
rect 8618 11536 8664 11582
rect 8741 11536 8787 11582
rect 8864 11536 8910 11582
rect 946 11225 2920 11271
rect 946 11001 2920 11047
rect 4870 11312 5120 11358
rect 5177 11312 5223 11358
rect 5280 11312 5326 11358
rect 5383 11312 5429 11358
rect 5486 11312 5532 11358
rect 5589 11312 5635 11358
rect 5692 11312 5738 11358
rect 5795 11312 5841 11358
rect 5898 11312 5944 11358
rect 6451 11312 6497 11358
rect 6568 11312 6614 11358
rect 6685 11312 6731 11358
rect 6803 11312 6849 11358
rect 6921 11312 6967 11358
rect 7039 11312 7085 11358
rect 18375 11536 18421 11582
rect 18478 11536 18524 11582
rect 18581 11536 18627 11582
rect 18684 11536 18730 11582
rect 18787 11536 18833 11582
rect 18890 11536 18936 11582
rect 18993 11536 19039 11582
rect 19096 11536 19142 11582
rect 19199 11536 19449 11582
rect 14409 11449 14455 11495
rect 14522 11449 14568 11495
rect 14635 11449 14681 11495
rect 14748 11449 14794 11495
rect 14861 11449 14907 11495
rect 8618 11312 8664 11358
rect 8741 11312 8787 11358
rect 8864 11312 8910 11358
rect 14409 11225 14455 11271
rect 14522 11225 14568 11271
rect 14635 11225 14681 11271
rect 14748 11225 14794 11271
rect 14861 11225 14907 11271
rect 18375 11312 18421 11358
rect 18478 11312 18524 11358
rect 18581 11312 18627 11358
rect 18684 11312 18730 11358
rect 18787 11312 18833 11358
rect 18890 11312 18936 11358
rect 18993 11312 19039 11358
rect 19096 11312 19142 11358
rect 19199 11312 19449 11358
rect 21399 11449 23373 11495
rect 4870 11088 5120 11134
rect 5177 11088 5223 11134
rect 5280 11088 5326 11134
rect 5383 11088 5429 11134
rect 5486 11088 5532 11134
rect 5589 11088 5635 11134
rect 5692 11088 5738 11134
rect 5795 11088 5841 11134
rect 5898 11088 5944 11134
rect 6451 11088 6497 11134
rect 6568 11088 6614 11134
rect 6685 11088 6731 11134
rect 6803 11088 6849 11134
rect 6921 11088 6967 11134
rect 7039 11088 7085 11134
rect 18375 11088 18421 11134
rect 18478 11088 18524 11134
rect 18581 11088 18627 11134
rect 18684 11088 18730 11134
rect 18787 11088 18833 11134
rect 18890 11088 18936 11134
rect 18993 11088 19039 11134
rect 19096 11088 19142 11134
rect 19199 11088 19449 11134
rect 14409 11001 14455 11047
rect 14522 11001 14568 11047
rect 14635 11001 14681 11047
rect 14748 11001 14794 11047
rect 14861 11001 14907 11047
rect 946 10777 2920 10823
rect 946 10553 2920 10599
rect 946 10329 2920 10375
rect 21399 11225 23373 11271
rect 21399 11001 23373 11047
rect 14409 10777 14455 10823
rect 14522 10777 14568 10823
rect 14635 10777 14681 10823
rect 14748 10777 14794 10823
rect 14861 10777 14907 10823
rect 21399 10777 23373 10823
rect 4870 10466 5120 10512
rect 5177 10466 5223 10512
rect 5280 10466 5326 10512
rect 5383 10466 5429 10512
rect 5486 10466 5532 10512
rect 5589 10466 5635 10512
rect 5692 10466 5738 10512
rect 5795 10466 5841 10512
rect 5898 10466 5944 10512
rect 6451 10466 6497 10512
rect 6568 10466 6614 10512
rect 6685 10466 6731 10512
rect 6803 10466 6849 10512
rect 6921 10466 6967 10512
rect 7039 10466 7085 10512
rect 14409 10553 14455 10599
rect 14522 10553 14568 10599
rect 14635 10553 14681 10599
rect 14748 10553 14794 10599
rect 14861 10553 14907 10599
rect 946 10105 2920 10151
rect 4870 10242 5120 10288
rect 5177 10242 5223 10288
rect 5280 10242 5326 10288
rect 5383 10242 5429 10288
rect 5486 10242 5532 10288
rect 5589 10242 5635 10288
rect 5692 10242 5738 10288
rect 5795 10242 5841 10288
rect 5898 10242 5944 10288
rect 18375 10466 18421 10512
rect 18478 10466 18524 10512
rect 18581 10466 18627 10512
rect 18684 10466 18730 10512
rect 18787 10466 18833 10512
rect 18890 10466 18936 10512
rect 18993 10466 19039 10512
rect 19096 10466 19142 10512
rect 19199 10466 19449 10512
rect 6451 10242 6497 10288
rect 6568 10242 6614 10288
rect 6685 10242 6731 10288
rect 6803 10242 6849 10288
rect 6921 10242 6967 10288
rect 7039 10242 7085 10288
rect 8618 10242 8664 10288
rect 8741 10242 8787 10288
rect 8864 10242 8910 10288
rect 14409 10329 14455 10375
rect 14522 10329 14568 10375
rect 14635 10329 14681 10375
rect 14748 10329 14794 10375
rect 14861 10329 14907 10375
rect 18375 10242 18421 10288
rect 18478 10242 18524 10288
rect 18581 10242 18627 10288
rect 18684 10242 18730 10288
rect 18787 10242 18833 10288
rect 18890 10242 18936 10288
rect 18993 10242 19039 10288
rect 19096 10242 19142 10288
rect 19199 10242 19449 10288
rect 4870 10018 5120 10064
rect 5177 10018 5223 10064
rect 5280 10018 5326 10064
rect 5383 10018 5429 10064
rect 5486 10018 5532 10064
rect 5589 10018 5635 10064
rect 5692 10018 5738 10064
rect 5795 10018 5841 10064
rect 5898 10018 5944 10064
rect 6451 10018 6497 10064
rect 6568 10018 6614 10064
rect 6685 10018 6731 10064
rect 6803 10018 6849 10064
rect 6921 10018 6967 10064
rect 7039 10018 7085 10064
rect 8618 10018 8664 10064
rect 8741 10018 8787 10064
rect 8864 10018 8910 10064
rect 14409 10105 14455 10151
rect 14522 10105 14568 10151
rect 14635 10105 14681 10151
rect 14748 10105 14794 10151
rect 14861 10105 14907 10151
rect 21399 10553 23373 10599
rect 21399 10329 23373 10375
rect 18375 10018 18421 10064
rect 18478 10018 18524 10064
rect 18581 10018 18627 10064
rect 18684 10018 18730 10064
rect 18787 10018 18833 10064
rect 18890 10018 18936 10064
rect 18993 10018 19039 10064
rect 19096 10018 19142 10064
rect 19199 10018 19449 10064
rect 21399 10105 23373 10151
rect 946 9649 2920 9695
rect 4870 9736 5120 9782
rect 5177 9736 5223 9782
rect 5280 9736 5326 9782
rect 5383 9736 5429 9782
rect 5486 9736 5532 9782
rect 5589 9736 5635 9782
rect 5692 9736 5738 9782
rect 5795 9736 5841 9782
rect 5898 9736 5944 9782
rect 6451 9736 6497 9782
rect 6568 9736 6614 9782
rect 6685 9736 6731 9782
rect 6803 9736 6849 9782
rect 6921 9736 6967 9782
rect 7039 9736 7085 9782
rect 8618 9736 8664 9782
rect 8741 9736 8787 9782
rect 8864 9736 8910 9782
rect 946 9425 2920 9471
rect 946 9201 2920 9247
rect 4870 9512 5120 9558
rect 5177 9512 5223 9558
rect 5280 9512 5326 9558
rect 5383 9512 5429 9558
rect 5486 9512 5532 9558
rect 5589 9512 5635 9558
rect 5692 9512 5738 9558
rect 5795 9512 5841 9558
rect 5898 9512 5944 9558
rect 6451 9512 6497 9558
rect 6568 9512 6614 9558
rect 6685 9512 6731 9558
rect 6803 9512 6849 9558
rect 6921 9512 6967 9558
rect 7039 9512 7085 9558
rect 18375 9736 18421 9782
rect 18478 9736 18524 9782
rect 18581 9736 18627 9782
rect 18684 9736 18730 9782
rect 18787 9736 18833 9782
rect 18890 9736 18936 9782
rect 18993 9736 19039 9782
rect 19096 9736 19142 9782
rect 19199 9736 19449 9782
rect 14409 9649 14455 9695
rect 14522 9649 14568 9695
rect 14635 9649 14681 9695
rect 14748 9649 14794 9695
rect 14861 9649 14907 9695
rect 8618 9512 8664 9558
rect 8741 9512 8787 9558
rect 8864 9512 8910 9558
rect 14409 9425 14455 9471
rect 14522 9425 14568 9471
rect 14635 9425 14681 9471
rect 14748 9425 14794 9471
rect 14861 9425 14907 9471
rect 18375 9512 18421 9558
rect 18478 9512 18524 9558
rect 18581 9512 18627 9558
rect 18684 9512 18730 9558
rect 18787 9512 18833 9558
rect 18890 9512 18936 9558
rect 18993 9512 19039 9558
rect 19096 9512 19142 9558
rect 19199 9512 19449 9558
rect 21399 9649 23373 9695
rect 4870 9288 5120 9334
rect 5177 9288 5223 9334
rect 5280 9288 5326 9334
rect 5383 9288 5429 9334
rect 5486 9288 5532 9334
rect 5589 9288 5635 9334
rect 5692 9288 5738 9334
rect 5795 9288 5841 9334
rect 5898 9288 5944 9334
rect 6451 9288 6497 9334
rect 6568 9288 6614 9334
rect 6685 9288 6731 9334
rect 6803 9288 6849 9334
rect 6921 9288 6967 9334
rect 7039 9288 7085 9334
rect 18375 9288 18421 9334
rect 18478 9288 18524 9334
rect 18581 9288 18627 9334
rect 18684 9288 18730 9334
rect 18787 9288 18833 9334
rect 18890 9288 18936 9334
rect 18993 9288 19039 9334
rect 19096 9288 19142 9334
rect 19199 9288 19449 9334
rect 14409 9201 14455 9247
rect 14522 9201 14568 9247
rect 14635 9201 14681 9247
rect 14748 9201 14794 9247
rect 14861 9201 14907 9247
rect 946 8977 2920 9023
rect 946 8753 2920 8799
rect 946 8529 2920 8575
rect 21399 9425 23373 9471
rect 21399 9201 23373 9247
rect 14409 8977 14455 9023
rect 14522 8977 14568 9023
rect 14635 8977 14681 9023
rect 14748 8977 14794 9023
rect 14861 8977 14907 9023
rect 21399 8977 23373 9023
rect 4870 8666 5120 8712
rect 5177 8666 5223 8712
rect 5280 8666 5326 8712
rect 5383 8666 5429 8712
rect 5486 8666 5532 8712
rect 5589 8666 5635 8712
rect 5692 8666 5738 8712
rect 5795 8666 5841 8712
rect 5898 8666 5944 8712
rect 6451 8666 6497 8712
rect 6568 8666 6614 8712
rect 6685 8666 6731 8712
rect 6803 8666 6849 8712
rect 6921 8666 6967 8712
rect 7039 8666 7085 8712
rect 14409 8753 14455 8799
rect 14522 8753 14568 8799
rect 14635 8753 14681 8799
rect 14748 8753 14794 8799
rect 14861 8753 14907 8799
rect 946 8305 2920 8351
rect 4870 8442 5120 8488
rect 5177 8442 5223 8488
rect 5280 8442 5326 8488
rect 5383 8442 5429 8488
rect 5486 8442 5532 8488
rect 5589 8442 5635 8488
rect 5692 8442 5738 8488
rect 5795 8442 5841 8488
rect 5898 8442 5944 8488
rect 18375 8666 18421 8712
rect 18478 8666 18524 8712
rect 18581 8666 18627 8712
rect 18684 8666 18730 8712
rect 18787 8666 18833 8712
rect 18890 8666 18936 8712
rect 18993 8666 19039 8712
rect 19096 8666 19142 8712
rect 19199 8666 19449 8712
rect 6451 8442 6497 8488
rect 6568 8442 6614 8488
rect 6685 8442 6731 8488
rect 6803 8442 6849 8488
rect 6921 8442 6967 8488
rect 7039 8442 7085 8488
rect 8618 8442 8664 8488
rect 8741 8442 8787 8488
rect 8864 8442 8910 8488
rect 14409 8529 14455 8575
rect 14522 8529 14568 8575
rect 14635 8529 14681 8575
rect 14748 8529 14794 8575
rect 14861 8529 14907 8575
rect 18375 8442 18421 8488
rect 18478 8442 18524 8488
rect 18581 8442 18627 8488
rect 18684 8442 18730 8488
rect 18787 8442 18833 8488
rect 18890 8442 18936 8488
rect 18993 8442 19039 8488
rect 19096 8442 19142 8488
rect 19199 8442 19449 8488
rect 4870 8218 5120 8264
rect 5177 8218 5223 8264
rect 5280 8218 5326 8264
rect 5383 8218 5429 8264
rect 5486 8218 5532 8264
rect 5589 8218 5635 8264
rect 5692 8218 5738 8264
rect 5795 8218 5841 8264
rect 5898 8218 5944 8264
rect 6451 8218 6497 8264
rect 6568 8218 6614 8264
rect 6685 8218 6731 8264
rect 6803 8218 6849 8264
rect 6921 8218 6967 8264
rect 7039 8218 7085 8264
rect 8618 8218 8664 8264
rect 8741 8218 8787 8264
rect 8864 8218 8910 8264
rect 14409 8305 14455 8351
rect 14522 8305 14568 8351
rect 14635 8305 14681 8351
rect 14748 8305 14794 8351
rect 14861 8305 14907 8351
rect 21399 8753 23373 8799
rect 21399 8529 23373 8575
rect 18375 8218 18421 8264
rect 18478 8218 18524 8264
rect 18581 8218 18627 8264
rect 18684 8218 18730 8264
rect 18787 8218 18833 8264
rect 18890 8218 18936 8264
rect 18993 8218 19039 8264
rect 19096 8218 19142 8264
rect 19199 8218 19449 8264
rect 21399 8305 23373 8351
rect 946 7849 2920 7895
rect 4870 7936 5120 7982
rect 5177 7936 5223 7982
rect 5280 7936 5326 7982
rect 5383 7936 5429 7982
rect 5486 7936 5532 7982
rect 5589 7936 5635 7982
rect 5692 7936 5738 7982
rect 5795 7936 5841 7982
rect 5898 7936 5944 7982
rect 6451 7936 6497 7982
rect 6568 7936 6614 7982
rect 6685 7936 6731 7982
rect 6803 7936 6849 7982
rect 6921 7936 6967 7982
rect 7039 7936 7085 7982
rect 8618 7936 8664 7982
rect 8741 7936 8787 7982
rect 8864 7936 8910 7982
rect 946 7625 2920 7671
rect 946 7401 2920 7447
rect 4870 7712 5120 7758
rect 5177 7712 5223 7758
rect 5280 7712 5326 7758
rect 5383 7712 5429 7758
rect 5486 7712 5532 7758
rect 5589 7712 5635 7758
rect 5692 7712 5738 7758
rect 5795 7712 5841 7758
rect 5898 7712 5944 7758
rect 6451 7712 6497 7758
rect 6568 7712 6614 7758
rect 6685 7712 6731 7758
rect 6803 7712 6849 7758
rect 6921 7712 6967 7758
rect 7039 7712 7085 7758
rect 18375 7936 18421 7982
rect 18478 7936 18524 7982
rect 18581 7936 18627 7982
rect 18684 7936 18730 7982
rect 18787 7936 18833 7982
rect 18890 7936 18936 7982
rect 18993 7936 19039 7982
rect 19096 7936 19142 7982
rect 19199 7936 19449 7982
rect 14409 7849 14455 7895
rect 14522 7849 14568 7895
rect 14635 7849 14681 7895
rect 14748 7849 14794 7895
rect 14861 7849 14907 7895
rect 8618 7712 8664 7758
rect 8741 7712 8787 7758
rect 8864 7712 8910 7758
rect 14409 7625 14455 7671
rect 14522 7625 14568 7671
rect 14635 7625 14681 7671
rect 14748 7625 14794 7671
rect 14861 7625 14907 7671
rect 18375 7712 18421 7758
rect 18478 7712 18524 7758
rect 18581 7712 18627 7758
rect 18684 7712 18730 7758
rect 18787 7712 18833 7758
rect 18890 7712 18936 7758
rect 18993 7712 19039 7758
rect 19096 7712 19142 7758
rect 19199 7712 19449 7758
rect 21399 7849 23373 7895
rect 4870 7488 5120 7534
rect 5177 7488 5223 7534
rect 5280 7488 5326 7534
rect 5383 7488 5429 7534
rect 5486 7488 5532 7534
rect 5589 7488 5635 7534
rect 5692 7488 5738 7534
rect 5795 7488 5841 7534
rect 5898 7488 5944 7534
rect 6451 7488 6497 7534
rect 6568 7488 6614 7534
rect 6685 7488 6731 7534
rect 6803 7488 6849 7534
rect 6921 7488 6967 7534
rect 7039 7488 7085 7534
rect 18375 7488 18421 7534
rect 18478 7488 18524 7534
rect 18581 7488 18627 7534
rect 18684 7488 18730 7534
rect 18787 7488 18833 7534
rect 18890 7488 18936 7534
rect 18993 7488 19039 7534
rect 19096 7488 19142 7534
rect 19199 7488 19449 7534
rect 14409 7401 14455 7447
rect 14522 7401 14568 7447
rect 14635 7401 14681 7447
rect 14748 7401 14794 7447
rect 14861 7401 14907 7447
rect 946 7177 2920 7223
rect 946 6953 2920 6999
rect 946 6729 2920 6775
rect 21399 7625 23373 7671
rect 21399 7401 23373 7447
rect 14409 7177 14455 7223
rect 14522 7177 14568 7223
rect 14635 7177 14681 7223
rect 14748 7177 14794 7223
rect 14861 7177 14907 7223
rect 21399 7177 23373 7223
rect 4870 6866 5120 6912
rect 5177 6866 5223 6912
rect 5280 6866 5326 6912
rect 5383 6866 5429 6912
rect 5486 6866 5532 6912
rect 5589 6866 5635 6912
rect 5692 6866 5738 6912
rect 5795 6866 5841 6912
rect 5898 6866 5944 6912
rect 6451 6866 6497 6912
rect 6568 6866 6614 6912
rect 6685 6866 6731 6912
rect 6803 6866 6849 6912
rect 6921 6866 6967 6912
rect 7039 6866 7085 6912
rect 14409 6953 14455 6999
rect 14522 6953 14568 6999
rect 14635 6953 14681 6999
rect 14748 6953 14794 6999
rect 14861 6953 14907 6999
rect 946 6505 2920 6551
rect 4870 6642 5120 6688
rect 5177 6642 5223 6688
rect 5280 6642 5326 6688
rect 5383 6642 5429 6688
rect 5486 6642 5532 6688
rect 5589 6642 5635 6688
rect 5692 6642 5738 6688
rect 5795 6642 5841 6688
rect 5898 6642 5944 6688
rect 18375 6866 18421 6912
rect 18478 6866 18524 6912
rect 18581 6866 18627 6912
rect 18684 6866 18730 6912
rect 18787 6866 18833 6912
rect 18890 6866 18936 6912
rect 18993 6866 19039 6912
rect 19096 6866 19142 6912
rect 19199 6866 19449 6912
rect 6451 6642 6497 6688
rect 6568 6642 6614 6688
rect 6685 6642 6731 6688
rect 6803 6642 6849 6688
rect 6921 6642 6967 6688
rect 7039 6642 7085 6688
rect 8618 6642 8664 6688
rect 8741 6642 8787 6688
rect 8864 6642 8910 6688
rect 14409 6729 14455 6775
rect 14522 6729 14568 6775
rect 14635 6729 14681 6775
rect 14748 6729 14794 6775
rect 14861 6729 14907 6775
rect 18375 6642 18421 6688
rect 18478 6642 18524 6688
rect 18581 6642 18627 6688
rect 18684 6642 18730 6688
rect 18787 6642 18833 6688
rect 18890 6642 18936 6688
rect 18993 6642 19039 6688
rect 19096 6642 19142 6688
rect 19199 6642 19449 6688
rect 4870 6418 5120 6464
rect 5177 6418 5223 6464
rect 5280 6418 5326 6464
rect 5383 6418 5429 6464
rect 5486 6418 5532 6464
rect 5589 6418 5635 6464
rect 5692 6418 5738 6464
rect 5795 6418 5841 6464
rect 5898 6418 5944 6464
rect 6451 6418 6497 6464
rect 6568 6418 6614 6464
rect 6685 6418 6731 6464
rect 6803 6418 6849 6464
rect 6921 6418 6967 6464
rect 7039 6418 7085 6464
rect 8618 6418 8664 6464
rect 8741 6418 8787 6464
rect 8864 6418 8910 6464
rect 14409 6505 14455 6551
rect 14522 6505 14568 6551
rect 14635 6505 14681 6551
rect 14748 6505 14794 6551
rect 14861 6505 14907 6551
rect 21399 6953 23373 6999
rect 21399 6729 23373 6775
rect 18375 6418 18421 6464
rect 18478 6418 18524 6464
rect 18581 6418 18627 6464
rect 18684 6418 18730 6464
rect 18787 6418 18833 6464
rect 18890 6418 18936 6464
rect 18993 6418 19039 6464
rect 19096 6418 19142 6464
rect 19199 6418 19449 6464
rect 21399 6505 23373 6551
rect 946 6049 2920 6095
rect 4870 6136 5120 6182
rect 5177 6136 5223 6182
rect 5280 6136 5326 6182
rect 5383 6136 5429 6182
rect 5486 6136 5532 6182
rect 5589 6136 5635 6182
rect 5692 6136 5738 6182
rect 5795 6136 5841 6182
rect 5898 6136 5944 6182
rect 6451 6136 6497 6182
rect 6568 6136 6614 6182
rect 6685 6136 6731 6182
rect 6803 6136 6849 6182
rect 6921 6136 6967 6182
rect 7039 6136 7085 6182
rect 8618 6136 8664 6182
rect 8741 6136 8787 6182
rect 8864 6136 8910 6182
rect 946 5825 2920 5871
rect 946 5601 2920 5647
rect 4870 5912 5120 5958
rect 5177 5912 5223 5958
rect 5280 5912 5326 5958
rect 5383 5912 5429 5958
rect 5486 5912 5532 5958
rect 5589 5912 5635 5958
rect 5692 5912 5738 5958
rect 5795 5912 5841 5958
rect 5898 5912 5944 5958
rect 6451 5912 6497 5958
rect 6568 5912 6614 5958
rect 6685 5912 6731 5958
rect 6803 5912 6849 5958
rect 6921 5912 6967 5958
rect 7039 5912 7085 5958
rect 18375 6136 18421 6182
rect 18478 6136 18524 6182
rect 18581 6136 18627 6182
rect 18684 6136 18730 6182
rect 18787 6136 18833 6182
rect 18890 6136 18936 6182
rect 18993 6136 19039 6182
rect 19096 6136 19142 6182
rect 19199 6136 19449 6182
rect 14409 6049 14455 6095
rect 14522 6049 14568 6095
rect 14635 6049 14681 6095
rect 14748 6049 14794 6095
rect 14861 6049 14907 6095
rect 8618 5912 8664 5958
rect 8741 5912 8787 5958
rect 8864 5912 8910 5958
rect 14409 5825 14455 5871
rect 14522 5825 14568 5871
rect 14635 5825 14681 5871
rect 14748 5825 14794 5871
rect 14861 5825 14907 5871
rect 18375 5912 18421 5958
rect 18478 5912 18524 5958
rect 18581 5912 18627 5958
rect 18684 5912 18730 5958
rect 18787 5912 18833 5958
rect 18890 5912 18936 5958
rect 18993 5912 19039 5958
rect 19096 5912 19142 5958
rect 19199 5912 19449 5958
rect 21399 6049 23373 6095
rect 4870 5688 5120 5734
rect 5177 5688 5223 5734
rect 5280 5688 5326 5734
rect 5383 5688 5429 5734
rect 5486 5688 5532 5734
rect 5589 5688 5635 5734
rect 5692 5688 5738 5734
rect 5795 5688 5841 5734
rect 5898 5688 5944 5734
rect 6451 5688 6497 5734
rect 6568 5688 6614 5734
rect 6685 5688 6731 5734
rect 6803 5688 6849 5734
rect 6921 5688 6967 5734
rect 7039 5688 7085 5734
rect 18375 5688 18421 5734
rect 18478 5688 18524 5734
rect 18581 5688 18627 5734
rect 18684 5688 18730 5734
rect 18787 5688 18833 5734
rect 18890 5688 18936 5734
rect 18993 5688 19039 5734
rect 19096 5688 19142 5734
rect 19199 5688 19449 5734
rect 14409 5601 14455 5647
rect 14522 5601 14568 5647
rect 14635 5601 14681 5647
rect 14748 5601 14794 5647
rect 14861 5601 14907 5647
rect 946 5377 2920 5423
rect 946 5153 2920 5199
rect 946 4929 2920 4975
rect 21399 5825 23373 5871
rect 21399 5601 23373 5647
rect 14409 5377 14455 5423
rect 14522 5377 14568 5423
rect 14635 5377 14681 5423
rect 14748 5377 14794 5423
rect 14861 5377 14907 5423
rect 21399 5377 23373 5423
rect 4870 5066 5120 5112
rect 5177 5066 5223 5112
rect 5280 5066 5326 5112
rect 5383 5066 5429 5112
rect 5486 5066 5532 5112
rect 5589 5066 5635 5112
rect 5692 5066 5738 5112
rect 5795 5066 5841 5112
rect 5898 5066 5944 5112
rect 6451 5066 6497 5112
rect 6568 5066 6614 5112
rect 6685 5066 6731 5112
rect 6803 5066 6849 5112
rect 6921 5066 6967 5112
rect 7039 5066 7085 5112
rect 14409 5153 14455 5199
rect 14522 5153 14568 5199
rect 14635 5153 14681 5199
rect 14748 5153 14794 5199
rect 14861 5153 14907 5199
rect 946 4705 2920 4751
rect 4870 4842 5120 4888
rect 5177 4842 5223 4888
rect 5280 4842 5326 4888
rect 5383 4842 5429 4888
rect 5486 4842 5532 4888
rect 5589 4842 5635 4888
rect 5692 4842 5738 4888
rect 5795 4842 5841 4888
rect 5898 4842 5944 4888
rect 18375 5066 18421 5112
rect 18478 5066 18524 5112
rect 18581 5066 18627 5112
rect 18684 5066 18730 5112
rect 18787 5066 18833 5112
rect 18890 5066 18936 5112
rect 18993 5066 19039 5112
rect 19096 5066 19142 5112
rect 19199 5066 19449 5112
rect 6451 4842 6497 4888
rect 6568 4842 6614 4888
rect 6685 4842 6731 4888
rect 6803 4842 6849 4888
rect 6921 4842 6967 4888
rect 7039 4842 7085 4888
rect 8618 4842 8664 4888
rect 8741 4842 8787 4888
rect 8864 4842 8910 4888
rect 14409 4929 14455 4975
rect 14522 4929 14568 4975
rect 14635 4929 14681 4975
rect 14748 4929 14794 4975
rect 14861 4929 14907 4975
rect 18375 4842 18421 4888
rect 18478 4842 18524 4888
rect 18581 4842 18627 4888
rect 18684 4842 18730 4888
rect 18787 4842 18833 4888
rect 18890 4842 18936 4888
rect 18993 4842 19039 4888
rect 19096 4842 19142 4888
rect 19199 4842 19449 4888
rect 4870 4618 5120 4664
rect 5177 4618 5223 4664
rect 5280 4618 5326 4664
rect 5383 4618 5429 4664
rect 5486 4618 5532 4664
rect 5589 4618 5635 4664
rect 5692 4618 5738 4664
rect 5795 4618 5841 4664
rect 5898 4618 5944 4664
rect 6451 4618 6497 4664
rect 6568 4618 6614 4664
rect 6685 4618 6731 4664
rect 6803 4618 6849 4664
rect 6921 4618 6967 4664
rect 7039 4618 7085 4664
rect 8618 4618 8664 4664
rect 8741 4618 8787 4664
rect 8864 4618 8910 4664
rect 14409 4705 14455 4751
rect 14522 4705 14568 4751
rect 14635 4705 14681 4751
rect 14748 4705 14794 4751
rect 14861 4705 14907 4751
rect 21399 5153 23373 5199
rect 21399 4929 23373 4975
rect 18375 4618 18421 4664
rect 18478 4618 18524 4664
rect 18581 4618 18627 4664
rect 18684 4618 18730 4664
rect 18787 4618 18833 4664
rect 18890 4618 18936 4664
rect 18993 4618 19039 4664
rect 19096 4618 19142 4664
rect 19199 4618 19449 4664
rect 21399 4705 23373 4751
rect 946 4249 2920 4295
rect 4870 4336 5120 4382
rect 5177 4336 5223 4382
rect 5280 4336 5326 4382
rect 5383 4336 5429 4382
rect 5486 4336 5532 4382
rect 5589 4336 5635 4382
rect 5692 4336 5738 4382
rect 5795 4336 5841 4382
rect 5898 4336 5944 4382
rect 6451 4336 6497 4382
rect 6568 4336 6614 4382
rect 6685 4336 6731 4382
rect 6803 4336 6849 4382
rect 6921 4336 6967 4382
rect 7039 4336 7085 4382
rect 8618 4336 8664 4382
rect 8741 4336 8787 4382
rect 8864 4336 8910 4382
rect 946 4025 2920 4071
rect 946 3801 2920 3847
rect 4870 4112 5120 4158
rect 5177 4112 5223 4158
rect 5280 4112 5326 4158
rect 5383 4112 5429 4158
rect 5486 4112 5532 4158
rect 5589 4112 5635 4158
rect 5692 4112 5738 4158
rect 5795 4112 5841 4158
rect 5898 4112 5944 4158
rect 6451 4112 6497 4158
rect 6568 4112 6614 4158
rect 6685 4112 6731 4158
rect 6803 4112 6849 4158
rect 6921 4112 6967 4158
rect 7039 4112 7085 4158
rect 18375 4336 18421 4382
rect 18478 4336 18524 4382
rect 18581 4336 18627 4382
rect 18684 4336 18730 4382
rect 18787 4336 18833 4382
rect 18890 4336 18936 4382
rect 18993 4336 19039 4382
rect 19096 4336 19142 4382
rect 19199 4336 19449 4382
rect 14409 4249 14455 4295
rect 14522 4249 14568 4295
rect 14635 4249 14681 4295
rect 14748 4249 14794 4295
rect 14861 4249 14907 4295
rect 8618 4112 8664 4158
rect 8741 4112 8787 4158
rect 8864 4112 8910 4158
rect 14409 4025 14455 4071
rect 14522 4025 14568 4071
rect 14635 4025 14681 4071
rect 14748 4025 14794 4071
rect 14861 4025 14907 4071
rect 18375 4112 18421 4158
rect 18478 4112 18524 4158
rect 18581 4112 18627 4158
rect 18684 4112 18730 4158
rect 18787 4112 18833 4158
rect 18890 4112 18936 4158
rect 18993 4112 19039 4158
rect 19096 4112 19142 4158
rect 19199 4112 19449 4158
rect 21399 4249 23373 4295
rect 4870 3888 5120 3934
rect 5177 3888 5223 3934
rect 5280 3888 5326 3934
rect 5383 3888 5429 3934
rect 5486 3888 5532 3934
rect 5589 3888 5635 3934
rect 5692 3888 5738 3934
rect 5795 3888 5841 3934
rect 5898 3888 5944 3934
rect 6451 3888 6497 3934
rect 6568 3888 6614 3934
rect 6685 3888 6731 3934
rect 6803 3888 6849 3934
rect 6921 3888 6967 3934
rect 7039 3888 7085 3934
rect 18375 3888 18421 3934
rect 18478 3888 18524 3934
rect 18581 3888 18627 3934
rect 18684 3888 18730 3934
rect 18787 3888 18833 3934
rect 18890 3888 18936 3934
rect 18993 3888 19039 3934
rect 19096 3888 19142 3934
rect 19199 3888 19449 3934
rect 14409 3801 14455 3847
rect 14522 3801 14568 3847
rect 14635 3801 14681 3847
rect 14748 3801 14794 3847
rect 14861 3801 14907 3847
rect 946 3577 2920 3623
rect 946 3353 2920 3399
rect 946 3129 2920 3175
rect 21399 4025 23373 4071
rect 21399 3801 23373 3847
rect 14409 3577 14455 3623
rect 14522 3577 14568 3623
rect 14635 3577 14681 3623
rect 14748 3577 14794 3623
rect 14861 3577 14907 3623
rect 21399 3577 23373 3623
rect 4870 3266 5120 3312
rect 5177 3266 5223 3312
rect 5280 3266 5326 3312
rect 5383 3266 5429 3312
rect 5486 3266 5532 3312
rect 5589 3266 5635 3312
rect 5692 3266 5738 3312
rect 5795 3266 5841 3312
rect 5898 3266 5944 3312
rect 6451 3266 6497 3312
rect 6568 3266 6614 3312
rect 6685 3266 6731 3312
rect 6803 3266 6849 3312
rect 6921 3266 6967 3312
rect 7039 3266 7085 3312
rect 14409 3353 14455 3399
rect 14522 3353 14568 3399
rect 14635 3353 14681 3399
rect 14748 3353 14794 3399
rect 14861 3353 14907 3399
rect 946 2905 2920 2951
rect 4870 3042 5120 3088
rect 5177 3042 5223 3088
rect 5280 3042 5326 3088
rect 5383 3042 5429 3088
rect 5486 3042 5532 3088
rect 5589 3042 5635 3088
rect 5692 3042 5738 3088
rect 5795 3042 5841 3088
rect 5898 3042 5944 3088
rect 18375 3266 18421 3312
rect 18478 3266 18524 3312
rect 18581 3266 18627 3312
rect 18684 3266 18730 3312
rect 18787 3266 18833 3312
rect 18890 3266 18936 3312
rect 18993 3266 19039 3312
rect 19096 3266 19142 3312
rect 19199 3266 19449 3312
rect 6451 3042 6497 3088
rect 6568 3042 6614 3088
rect 6685 3042 6731 3088
rect 6803 3042 6849 3088
rect 6921 3042 6967 3088
rect 7039 3042 7085 3088
rect 8618 3042 8664 3088
rect 8741 3042 8787 3088
rect 8864 3042 8910 3088
rect 14409 3129 14455 3175
rect 14522 3129 14568 3175
rect 14635 3129 14681 3175
rect 14748 3129 14794 3175
rect 14861 3129 14907 3175
rect 18375 3042 18421 3088
rect 18478 3042 18524 3088
rect 18581 3042 18627 3088
rect 18684 3042 18730 3088
rect 18787 3042 18833 3088
rect 18890 3042 18936 3088
rect 18993 3042 19039 3088
rect 19096 3042 19142 3088
rect 19199 3042 19449 3088
rect 4870 2818 5120 2864
rect 5177 2818 5223 2864
rect 5280 2818 5326 2864
rect 5383 2818 5429 2864
rect 5486 2818 5532 2864
rect 5589 2818 5635 2864
rect 5692 2818 5738 2864
rect 5795 2818 5841 2864
rect 5898 2818 5944 2864
rect 6451 2818 6497 2864
rect 6568 2818 6614 2864
rect 6685 2818 6731 2864
rect 6803 2818 6849 2864
rect 6921 2818 6967 2864
rect 7039 2818 7085 2864
rect 8618 2818 8664 2864
rect 8741 2818 8787 2864
rect 8864 2818 8910 2864
rect 14409 2905 14455 2951
rect 14522 2905 14568 2951
rect 14635 2905 14681 2951
rect 14748 2905 14794 2951
rect 14861 2905 14907 2951
rect 21399 3353 23373 3399
rect 21399 3129 23373 3175
rect 18375 2818 18421 2864
rect 18478 2818 18524 2864
rect 18581 2818 18627 2864
rect 18684 2818 18730 2864
rect 18787 2818 18833 2864
rect 18890 2818 18936 2864
rect 18993 2818 19039 2864
rect 19096 2818 19142 2864
rect 19199 2818 19449 2864
rect 21399 2905 23373 2951
rect 946 2449 2920 2495
rect 4870 2536 5120 2582
rect 5177 2536 5223 2582
rect 5280 2536 5326 2582
rect 5383 2536 5429 2582
rect 5486 2536 5532 2582
rect 5589 2536 5635 2582
rect 5692 2536 5738 2582
rect 5795 2536 5841 2582
rect 5898 2536 5944 2582
rect 6451 2536 6497 2582
rect 6568 2536 6614 2582
rect 6685 2536 6731 2582
rect 6803 2536 6849 2582
rect 6921 2536 6967 2582
rect 7039 2536 7085 2582
rect 8618 2536 8664 2582
rect 8741 2536 8787 2582
rect 8864 2536 8910 2582
rect 946 2225 2920 2271
rect 946 2001 2920 2047
rect 4870 2312 5120 2358
rect 5177 2312 5223 2358
rect 5280 2312 5326 2358
rect 5383 2312 5429 2358
rect 5486 2312 5532 2358
rect 5589 2312 5635 2358
rect 5692 2312 5738 2358
rect 5795 2312 5841 2358
rect 5898 2312 5944 2358
rect 6451 2312 6497 2358
rect 6568 2312 6614 2358
rect 6685 2312 6731 2358
rect 6803 2312 6849 2358
rect 6921 2312 6967 2358
rect 7039 2312 7085 2358
rect 18375 2536 18421 2582
rect 18478 2536 18524 2582
rect 18581 2536 18627 2582
rect 18684 2536 18730 2582
rect 18787 2536 18833 2582
rect 18890 2536 18936 2582
rect 18993 2536 19039 2582
rect 19096 2536 19142 2582
rect 19199 2536 19449 2582
rect 14409 2449 14455 2495
rect 14522 2449 14568 2495
rect 14635 2449 14681 2495
rect 14748 2449 14794 2495
rect 14861 2449 14907 2495
rect 8618 2312 8664 2358
rect 8741 2312 8787 2358
rect 8864 2312 8910 2358
rect 14409 2225 14455 2271
rect 14522 2225 14568 2271
rect 14635 2225 14681 2271
rect 14748 2225 14794 2271
rect 14861 2225 14907 2271
rect 18375 2312 18421 2358
rect 18478 2312 18524 2358
rect 18581 2312 18627 2358
rect 18684 2312 18730 2358
rect 18787 2312 18833 2358
rect 18890 2312 18936 2358
rect 18993 2312 19039 2358
rect 19096 2312 19142 2358
rect 19199 2312 19449 2358
rect 21399 2449 23373 2495
rect 4870 2088 5120 2134
rect 5177 2088 5223 2134
rect 5280 2088 5326 2134
rect 5383 2088 5429 2134
rect 5486 2088 5532 2134
rect 5589 2088 5635 2134
rect 5692 2088 5738 2134
rect 5795 2088 5841 2134
rect 5898 2088 5944 2134
rect 6451 2088 6497 2134
rect 6568 2088 6614 2134
rect 6685 2088 6731 2134
rect 6803 2088 6849 2134
rect 6921 2088 6967 2134
rect 7039 2088 7085 2134
rect 18375 2088 18421 2134
rect 18478 2088 18524 2134
rect 18581 2088 18627 2134
rect 18684 2088 18730 2134
rect 18787 2088 18833 2134
rect 18890 2088 18936 2134
rect 18993 2088 19039 2134
rect 19096 2088 19142 2134
rect 19199 2088 19449 2134
rect 14409 2001 14455 2047
rect 14522 2001 14568 2047
rect 14635 2001 14681 2047
rect 14748 2001 14794 2047
rect 14861 2001 14907 2047
rect 946 1777 2920 1823
rect 946 1553 2920 1599
rect 946 1329 2920 1375
rect 21399 2225 23373 2271
rect 21399 2001 23373 2047
rect 14409 1777 14455 1823
rect 14522 1777 14568 1823
rect 14635 1777 14681 1823
rect 14748 1777 14794 1823
rect 14861 1777 14907 1823
rect 21399 1777 23373 1823
rect 4870 1466 5120 1512
rect 5177 1466 5223 1512
rect 5280 1466 5326 1512
rect 5383 1466 5429 1512
rect 5486 1466 5532 1512
rect 5589 1466 5635 1512
rect 5692 1466 5738 1512
rect 5795 1466 5841 1512
rect 5898 1466 5944 1512
rect 6451 1466 6497 1512
rect 6568 1466 6614 1512
rect 6685 1466 6731 1512
rect 6803 1466 6849 1512
rect 6921 1466 6967 1512
rect 7039 1466 7085 1512
rect 14409 1553 14455 1599
rect 14522 1553 14568 1599
rect 14635 1553 14681 1599
rect 14748 1553 14794 1599
rect 14861 1553 14907 1599
rect 946 1105 2920 1151
rect 4870 1242 5120 1288
rect 5177 1242 5223 1288
rect 5280 1242 5326 1288
rect 5383 1242 5429 1288
rect 5486 1242 5532 1288
rect 5589 1242 5635 1288
rect 5692 1242 5738 1288
rect 5795 1242 5841 1288
rect 5898 1242 5944 1288
rect 18375 1466 18421 1512
rect 18478 1466 18524 1512
rect 18581 1466 18627 1512
rect 18684 1466 18730 1512
rect 18787 1466 18833 1512
rect 18890 1466 18936 1512
rect 18993 1466 19039 1512
rect 19096 1466 19142 1512
rect 19199 1466 19449 1512
rect 6451 1242 6497 1288
rect 6568 1242 6614 1288
rect 6685 1242 6731 1288
rect 6803 1242 6849 1288
rect 6921 1242 6967 1288
rect 7039 1242 7085 1288
rect 8618 1242 8664 1288
rect 8741 1242 8787 1288
rect 8864 1242 8910 1288
rect 14409 1329 14455 1375
rect 14522 1329 14568 1375
rect 14635 1329 14681 1375
rect 14748 1329 14794 1375
rect 14861 1329 14907 1375
rect 18375 1242 18421 1288
rect 18478 1242 18524 1288
rect 18581 1242 18627 1288
rect 18684 1242 18730 1288
rect 18787 1242 18833 1288
rect 18890 1242 18936 1288
rect 18993 1242 19039 1288
rect 19096 1242 19142 1288
rect 19199 1242 19449 1288
rect 4870 1018 5120 1064
rect 5177 1018 5223 1064
rect 5280 1018 5326 1064
rect 5383 1018 5429 1064
rect 5486 1018 5532 1064
rect 5589 1018 5635 1064
rect 5692 1018 5738 1064
rect 5795 1018 5841 1064
rect 5898 1018 5944 1064
rect 6451 1018 6497 1064
rect 6568 1018 6614 1064
rect 6685 1018 6731 1064
rect 6803 1018 6849 1064
rect 6921 1018 6967 1064
rect 7039 1018 7085 1064
rect 8618 1018 8664 1064
rect 8741 1018 8787 1064
rect 8864 1018 8910 1064
rect 14409 1105 14455 1151
rect 14522 1105 14568 1151
rect 14635 1105 14681 1151
rect 14748 1105 14794 1151
rect 14861 1105 14907 1151
rect 21399 1553 23373 1599
rect 21399 1329 23373 1375
rect 18375 1018 18421 1064
rect 18478 1018 18524 1064
rect 18581 1018 18627 1064
rect 18684 1018 18730 1064
rect 18787 1018 18833 1064
rect 18890 1018 18936 1064
rect 18993 1018 19039 1064
rect 19096 1018 19142 1064
rect 19199 1018 19449 1064
rect 21399 1105 23373 1151
rect 946 649 2920 695
rect 4870 736 5120 782
rect 5177 736 5223 782
rect 5280 736 5326 782
rect 5383 736 5429 782
rect 5486 736 5532 782
rect 5589 736 5635 782
rect 5692 736 5738 782
rect 5795 736 5841 782
rect 5898 736 5944 782
rect 6451 736 6497 782
rect 6568 736 6614 782
rect 6685 736 6731 782
rect 6803 736 6849 782
rect 6921 736 6967 782
rect 7039 736 7085 782
rect 8618 736 8664 782
rect 8741 736 8787 782
rect 8864 736 8910 782
rect 946 425 2920 471
rect 946 201 2920 247
rect 4870 512 5120 558
rect 5177 512 5223 558
rect 5280 512 5326 558
rect 5383 512 5429 558
rect 5486 512 5532 558
rect 5589 512 5635 558
rect 5692 512 5738 558
rect 5795 512 5841 558
rect 5898 512 5944 558
rect 6451 512 6497 558
rect 6568 512 6614 558
rect 6685 512 6731 558
rect 6803 512 6849 558
rect 6921 512 6967 558
rect 7039 512 7085 558
rect 18375 736 18421 782
rect 18478 736 18524 782
rect 18581 736 18627 782
rect 18684 736 18730 782
rect 18787 736 18833 782
rect 18890 736 18936 782
rect 18993 736 19039 782
rect 19096 736 19142 782
rect 19199 736 19449 782
rect 14409 649 14455 695
rect 14522 649 14568 695
rect 14635 649 14681 695
rect 14748 649 14794 695
rect 14861 649 14907 695
rect 8618 512 8664 558
rect 8741 512 8787 558
rect 8864 512 8910 558
rect 14409 425 14455 471
rect 14522 425 14568 471
rect 14635 425 14681 471
rect 14748 425 14794 471
rect 14861 425 14907 471
rect 18375 512 18421 558
rect 18478 512 18524 558
rect 18581 512 18627 558
rect 18684 512 18730 558
rect 18787 512 18833 558
rect 18890 512 18936 558
rect 18993 512 19039 558
rect 19096 512 19142 558
rect 19199 512 19449 558
rect 21399 649 23373 695
rect 4870 288 5120 334
rect 5177 288 5223 334
rect 5280 288 5326 334
rect 5383 288 5429 334
rect 5486 288 5532 334
rect 5589 288 5635 334
rect 5692 288 5738 334
rect 5795 288 5841 334
rect 5898 288 5944 334
rect 6451 288 6497 334
rect 6568 288 6614 334
rect 6685 288 6731 334
rect 6803 288 6849 334
rect 6921 288 6967 334
rect 7039 288 7085 334
rect 18375 288 18421 334
rect 18478 288 18524 334
rect 18581 288 18627 334
rect 18684 288 18730 334
rect 18787 288 18833 334
rect 18890 288 18936 334
rect 18993 288 19039 334
rect 19096 288 19142 334
rect 19199 288 19449 334
rect 14409 201 14455 247
rect 14522 201 14568 247
rect 14635 201 14681 247
rect 14748 201 14794 247
rect 14861 201 14907 247
rect 946 -23 2920 23
rect 21399 425 23373 471
rect 21399 201 23373 247
rect 14409 -23 14455 23
rect 14522 -23 14568 23
rect 14635 -23 14681 23
rect 14748 -23 14794 23
rect 14861 -23 14907 23
rect 21399 -23 23373 23
<< psubdiff >>
rect 7535 14423 8089 14442
rect 7535 14377 7554 14423
rect 8070 14377 8089 14423
rect 7535 14358 8089 14377
rect 10376 14423 12592 14483
rect 10376 14377 10433 14423
rect 10479 14377 10591 14423
rect 10637 14377 10749 14423
rect 10795 14377 10907 14423
rect 10953 14377 11066 14423
rect 11112 14377 11224 14423
rect 11270 14377 11382 14423
rect 11428 14377 11540 14423
rect 11586 14377 11698 14423
rect 11744 14377 11856 14423
rect 11902 14377 12015 14423
rect 12061 14377 12173 14423
rect 12219 14377 12331 14423
rect 12377 14377 12489 14423
rect 12535 14377 12592 14423
rect 10376 14317 12592 14377
rect 4458 13523 4614 13580
rect 4458 13477 4513 13523
rect 4559 13477 4614 13523
rect 4458 13420 4614 13477
rect 19700 13523 19860 13583
rect 19700 13477 19757 13523
rect 19803 13477 19860 13523
rect 19700 13417 19860 13477
rect 7535 12623 8089 12642
rect 7535 12577 7554 12623
rect 8070 12577 8089 12623
rect 7535 12558 8089 12577
rect 10376 12623 12592 12683
rect 10376 12577 10433 12623
rect 10479 12577 10591 12623
rect 10637 12577 10749 12623
rect 10795 12577 10907 12623
rect 10953 12577 11066 12623
rect 11112 12577 11224 12623
rect 11270 12577 11382 12623
rect 11428 12577 11540 12623
rect 11586 12577 11698 12623
rect 11744 12577 11856 12623
rect 11902 12577 12015 12623
rect 12061 12577 12173 12623
rect 12219 12577 12331 12623
rect 12377 12577 12489 12623
rect 12535 12577 12592 12623
rect 10376 12517 12592 12577
rect 4458 11723 4614 11780
rect 4458 11677 4513 11723
rect 4559 11677 4614 11723
rect 4458 11620 4614 11677
rect 19700 11723 19860 11783
rect 19700 11677 19757 11723
rect 19803 11677 19860 11723
rect 19700 11617 19860 11677
rect 7535 10823 8089 10842
rect 7535 10777 7554 10823
rect 8070 10777 8089 10823
rect 7535 10758 8089 10777
rect 10376 10823 12592 10883
rect 10376 10777 10433 10823
rect 10479 10777 10591 10823
rect 10637 10777 10749 10823
rect 10795 10777 10907 10823
rect 10953 10777 11066 10823
rect 11112 10777 11224 10823
rect 11270 10777 11382 10823
rect 11428 10777 11540 10823
rect 11586 10777 11698 10823
rect 11744 10777 11856 10823
rect 11902 10777 12015 10823
rect 12061 10777 12173 10823
rect 12219 10777 12331 10823
rect 12377 10777 12489 10823
rect 12535 10777 12592 10823
rect 10376 10717 12592 10777
rect 4458 9923 4614 9980
rect 4458 9877 4513 9923
rect 4559 9877 4614 9923
rect 4458 9820 4614 9877
rect 19700 9923 19860 9983
rect 19700 9877 19757 9923
rect 19803 9877 19860 9923
rect 19700 9817 19860 9877
rect 7535 9023 8089 9042
rect 7535 8977 7554 9023
rect 8070 8977 8089 9023
rect 7535 8958 8089 8977
rect 10376 9023 12592 9083
rect 10376 8977 10433 9023
rect 10479 8977 10591 9023
rect 10637 8977 10749 9023
rect 10795 8977 10907 9023
rect 10953 8977 11066 9023
rect 11112 8977 11224 9023
rect 11270 8977 11382 9023
rect 11428 8977 11540 9023
rect 11586 8977 11698 9023
rect 11744 8977 11856 9023
rect 11902 8977 12015 9023
rect 12061 8977 12173 9023
rect 12219 8977 12331 9023
rect 12377 8977 12489 9023
rect 12535 8977 12592 9023
rect 10376 8917 12592 8977
rect 4458 8123 4614 8180
rect 4458 8077 4513 8123
rect 4559 8077 4614 8123
rect 4458 8020 4614 8077
rect 19700 8123 19860 8183
rect 19700 8077 19757 8123
rect 19803 8077 19860 8123
rect 19700 8017 19860 8077
rect 7535 7223 8089 7242
rect 7535 7177 7554 7223
rect 8070 7177 8089 7223
rect 7535 7158 8089 7177
rect 10376 7223 12592 7283
rect 10376 7177 10433 7223
rect 10479 7177 10591 7223
rect 10637 7177 10749 7223
rect 10795 7177 10907 7223
rect 10953 7177 11066 7223
rect 11112 7177 11224 7223
rect 11270 7177 11382 7223
rect 11428 7177 11540 7223
rect 11586 7177 11698 7223
rect 11744 7177 11856 7223
rect 11902 7177 12015 7223
rect 12061 7177 12173 7223
rect 12219 7177 12331 7223
rect 12377 7177 12489 7223
rect 12535 7177 12592 7223
rect 10376 7117 12592 7177
rect 4458 6323 4614 6380
rect 4458 6277 4513 6323
rect 4559 6277 4614 6323
rect 4458 6220 4614 6277
rect 19700 6323 19860 6383
rect 19700 6277 19757 6323
rect 19803 6277 19860 6323
rect 19700 6217 19860 6277
rect 7535 5423 8089 5442
rect 7535 5377 7554 5423
rect 8070 5377 8089 5423
rect 7535 5358 8089 5377
rect 10376 5423 12592 5483
rect 10376 5377 10433 5423
rect 10479 5377 10591 5423
rect 10637 5377 10749 5423
rect 10795 5377 10907 5423
rect 10953 5377 11066 5423
rect 11112 5377 11224 5423
rect 11270 5377 11382 5423
rect 11428 5377 11540 5423
rect 11586 5377 11698 5423
rect 11744 5377 11856 5423
rect 11902 5377 12015 5423
rect 12061 5377 12173 5423
rect 12219 5377 12331 5423
rect 12377 5377 12489 5423
rect 12535 5377 12592 5423
rect 10376 5317 12592 5377
rect 4458 4523 4614 4580
rect 4458 4477 4513 4523
rect 4559 4477 4614 4523
rect 4458 4420 4614 4477
rect 19700 4523 19860 4583
rect 19700 4477 19757 4523
rect 19803 4477 19860 4523
rect 19700 4417 19860 4477
rect 7535 3623 8089 3642
rect 7535 3577 7554 3623
rect 8070 3577 8089 3623
rect 7535 3558 8089 3577
rect 10376 3623 12592 3683
rect 10376 3577 10433 3623
rect 10479 3577 10591 3623
rect 10637 3577 10749 3623
rect 10795 3577 10907 3623
rect 10953 3577 11066 3623
rect 11112 3577 11224 3623
rect 11270 3577 11382 3623
rect 11428 3577 11540 3623
rect 11586 3577 11698 3623
rect 11744 3577 11856 3623
rect 11902 3577 12015 3623
rect 12061 3577 12173 3623
rect 12219 3577 12331 3623
rect 12377 3577 12489 3623
rect 12535 3577 12592 3623
rect 10376 3517 12592 3577
rect 4458 2723 4614 2780
rect 4458 2677 4513 2723
rect 4559 2677 4614 2723
rect 4458 2620 4614 2677
rect 19700 2723 19860 2783
rect 19700 2677 19757 2723
rect 19803 2677 19860 2723
rect 19700 2617 19860 2677
rect 7535 1823 8089 1842
rect 7535 1777 7554 1823
rect 8070 1777 8089 1823
rect 7535 1758 8089 1777
rect 10376 1823 12592 1883
rect 10376 1777 10433 1823
rect 10479 1777 10591 1823
rect 10637 1777 10749 1823
rect 10795 1777 10907 1823
rect 10953 1777 11066 1823
rect 11112 1777 11224 1823
rect 11270 1777 11382 1823
rect 11428 1777 11540 1823
rect 11586 1777 11698 1823
rect 11744 1777 11856 1823
rect 11902 1777 12015 1823
rect 12061 1777 12173 1823
rect 12219 1777 12331 1823
rect 12377 1777 12489 1823
rect 12535 1777 12592 1823
rect 10376 1717 12592 1777
rect 4458 923 4614 980
rect 4458 877 4513 923
rect 4559 877 4614 923
rect 4458 820 4614 877
rect 19700 923 19860 983
rect 19700 877 19757 923
rect 19803 877 19860 923
rect 19700 817 19860 877
rect 7535 23 8089 42
rect 7535 -23 7554 23
rect 8070 -23 8089 23
rect 7535 -42 8089 -23
rect 10376 23 12592 83
rect 10376 -23 10433 23
rect 10479 -23 10591 23
rect 10637 -23 10749 23
rect 10795 -23 10907 23
rect 10953 -23 11066 23
rect 11112 -23 11224 23
rect 11270 -23 11382 23
rect 11428 -23 11540 23
rect 11586 -23 11698 23
rect 11744 -23 11856 23
rect 11902 -23 12015 23
rect 12061 -23 12173 23
rect 12219 -23 12331 23
rect 12377 -23 12489 23
rect 12535 -23 12592 23
rect 10376 -83 12592 -23
<< nsubdiff >>
rect 397 14299 553 14462
rect 5945 14423 6458 14469
rect 5945 14377 6086 14423
rect 6320 14377 6458 14423
rect 397 14253 452 14299
rect 498 14253 553 14299
rect 397 14135 553 14253
rect 397 14089 452 14135
rect 498 14089 553 14135
rect 397 13972 553 14089
rect 397 13926 452 13972
rect 498 13926 553 13972
rect 397 13809 553 13926
rect 397 13763 452 13809
rect 498 13763 553 13809
rect 5945 14331 6458 14377
rect 8604 14423 8918 14480
rect 8604 14377 8659 14423
rect 8705 14377 8817 14423
rect 8863 14377 8918 14423
rect 8604 14320 8918 14377
rect 15161 14469 18163 14480
rect 15161 14423 18363 14469
rect 15161 14377 15216 14423
rect 15262 14377 15374 14423
rect 15420 14377 15532 14423
rect 15578 14377 15690 14423
rect 15736 14377 15848 14423
rect 15894 14377 16006 14423
rect 16052 14377 16165 14423
rect 16211 14377 16323 14423
rect 16369 14377 16481 14423
rect 16527 14377 16639 14423
rect 16685 14377 16797 14423
rect 16843 14377 16955 14423
rect 17001 14377 17113 14423
rect 17159 14377 17272 14423
rect 17318 14377 17430 14423
rect 17476 14377 17588 14423
rect 17634 14377 17746 14423
rect 17792 14377 17904 14423
rect 17950 14377 18062 14423
rect 18108 14377 18363 14423
rect 15161 14331 18363 14377
rect 15161 14259 18163 14331
rect 15161 14213 15216 14259
rect 15262 14213 15374 14259
rect 15420 14213 15532 14259
rect 15578 14213 15690 14259
rect 15736 14213 15848 14259
rect 15894 14213 16006 14259
rect 16052 14213 16165 14259
rect 16211 14213 16323 14259
rect 16369 14213 16481 14259
rect 16527 14213 16639 14259
rect 16685 14213 16797 14259
rect 16843 14213 16955 14259
rect 17001 14213 17113 14259
rect 17159 14213 17272 14259
rect 17318 14213 17430 14259
rect 17476 14213 17588 14259
rect 17634 14213 17746 14259
rect 17792 14213 17904 14259
rect 17950 14213 18062 14259
rect 18108 14213 18163 14259
rect 23765 14299 23921 14462
rect 23765 14253 23820 14299
rect 23866 14253 23921 14299
rect 15161 14156 18163 14213
rect 397 13646 553 13763
rect 397 13600 452 13646
rect 498 13600 553 13646
rect 23765 14135 23921 14253
rect 23765 14089 23820 14135
rect 23866 14089 23921 14135
rect 23765 13646 23921 14089
rect 397 13400 553 13600
rect 23765 13600 23820 13646
rect 23866 13600 23921 13646
rect 397 13354 452 13400
rect 498 13354 553 13400
rect 23765 13400 23921 13600
rect 397 13237 553 13354
rect 397 13191 452 13237
rect 498 13191 553 13237
rect 397 13074 553 13191
rect 397 13028 452 13074
rect 498 13028 553 13074
rect 397 12911 553 13028
rect 397 12865 452 12911
rect 498 12865 553 12911
rect 397 12747 553 12865
rect 397 12701 452 12747
rect 498 12701 553 12747
rect 397 12499 553 12701
rect 23765 13354 23820 13400
rect 23866 13354 23921 13400
rect 5945 12623 6458 12669
rect 5945 12577 6086 12623
rect 6320 12577 6458 12623
rect 397 12453 452 12499
rect 498 12453 553 12499
rect 397 12335 553 12453
rect 397 12289 452 12335
rect 498 12289 553 12335
rect 397 12172 553 12289
rect 397 12126 452 12172
rect 498 12126 553 12172
rect 397 12009 553 12126
rect 397 11963 452 12009
rect 498 11963 553 12009
rect 5945 12531 6458 12577
rect 8604 12623 8918 12680
rect 8604 12577 8659 12623
rect 8705 12577 8817 12623
rect 8863 12577 8918 12623
rect 8604 12520 8918 12577
rect 15161 12787 18163 12844
rect 15161 12741 15216 12787
rect 15262 12741 15374 12787
rect 15420 12741 15532 12787
rect 15578 12741 15690 12787
rect 15736 12741 15848 12787
rect 15894 12741 16006 12787
rect 16052 12741 16165 12787
rect 16211 12741 16323 12787
rect 16369 12741 16481 12787
rect 16527 12741 16639 12787
rect 16685 12741 16797 12787
rect 16843 12741 16955 12787
rect 17001 12741 17113 12787
rect 17159 12741 17272 12787
rect 17318 12741 17430 12787
rect 17476 12741 17588 12787
rect 17634 12741 17746 12787
rect 17792 12741 17904 12787
rect 17950 12741 18062 12787
rect 18108 12741 18163 12787
rect 23765 12911 23921 13354
rect 23765 12865 23820 12911
rect 23866 12865 23921 12911
rect 15161 12669 18163 12741
rect 15161 12623 18363 12669
rect 23765 12747 23921 12865
rect 23765 12701 23820 12747
rect 23866 12701 23921 12747
rect 15161 12577 15216 12623
rect 15262 12577 15374 12623
rect 15420 12577 15532 12623
rect 15578 12577 15690 12623
rect 15736 12577 15848 12623
rect 15894 12577 16006 12623
rect 16052 12577 16165 12623
rect 16211 12577 16323 12623
rect 16369 12577 16481 12623
rect 16527 12577 16639 12623
rect 16685 12577 16797 12623
rect 16843 12577 16955 12623
rect 17001 12577 17113 12623
rect 17159 12577 17272 12623
rect 17318 12577 17430 12623
rect 17476 12577 17588 12623
rect 17634 12577 17746 12623
rect 17792 12577 17904 12623
rect 17950 12577 18062 12623
rect 18108 12577 18363 12623
rect 15161 12531 18363 12577
rect 15161 12459 18163 12531
rect 15161 12413 15216 12459
rect 15262 12413 15374 12459
rect 15420 12413 15532 12459
rect 15578 12413 15690 12459
rect 15736 12413 15848 12459
rect 15894 12413 16006 12459
rect 16052 12413 16165 12459
rect 16211 12413 16323 12459
rect 16369 12413 16481 12459
rect 16527 12413 16639 12459
rect 16685 12413 16797 12459
rect 16843 12413 16955 12459
rect 17001 12413 17113 12459
rect 17159 12413 17272 12459
rect 17318 12413 17430 12459
rect 17476 12413 17588 12459
rect 17634 12413 17746 12459
rect 17792 12413 17904 12459
rect 17950 12413 18062 12459
rect 18108 12413 18163 12459
rect 23765 12499 23921 12701
rect 23765 12453 23820 12499
rect 23866 12453 23921 12499
rect 15161 12356 18163 12413
rect 397 11846 553 11963
rect 397 11800 452 11846
rect 498 11800 553 11846
rect 23765 12335 23921 12453
rect 23765 12289 23820 12335
rect 23866 12289 23921 12335
rect 23765 11846 23921 12289
rect 397 11600 553 11800
rect 23765 11800 23820 11846
rect 23866 11800 23921 11846
rect 397 11554 452 11600
rect 498 11554 553 11600
rect 23765 11600 23921 11800
rect 397 11437 553 11554
rect 397 11391 452 11437
rect 498 11391 553 11437
rect 397 11274 553 11391
rect 397 11228 452 11274
rect 498 11228 553 11274
rect 397 11111 553 11228
rect 397 11065 452 11111
rect 498 11065 553 11111
rect 397 10947 553 11065
rect 397 10901 452 10947
rect 498 10901 553 10947
rect 397 10699 553 10901
rect 23765 11554 23820 11600
rect 23866 11554 23921 11600
rect 5945 10823 6458 10869
rect 5945 10777 6086 10823
rect 6320 10777 6458 10823
rect 397 10653 452 10699
rect 498 10653 553 10699
rect 397 10535 553 10653
rect 397 10489 452 10535
rect 498 10489 553 10535
rect 397 10372 553 10489
rect 397 10326 452 10372
rect 498 10326 553 10372
rect 397 10209 553 10326
rect 397 10163 452 10209
rect 498 10163 553 10209
rect 5945 10731 6458 10777
rect 8604 10823 8918 10880
rect 8604 10777 8659 10823
rect 8705 10777 8817 10823
rect 8863 10777 8918 10823
rect 8604 10720 8918 10777
rect 15161 10987 18163 11044
rect 15161 10941 15216 10987
rect 15262 10941 15374 10987
rect 15420 10941 15532 10987
rect 15578 10941 15690 10987
rect 15736 10941 15848 10987
rect 15894 10941 16006 10987
rect 16052 10941 16165 10987
rect 16211 10941 16323 10987
rect 16369 10941 16481 10987
rect 16527 10941 16639 10987
rect 16685 10941 16797 10987
rect 16843 10941 16955 10987
rect 17001 10941 17113 10987
rect 17159 10941 17272 10987
rect 17318 10941 17430 10987
rect 17476 10941 17588 10987
rect 17634 10941 17746 10987
rect 17792 10941 17904 10987
rect 17950 10941 18062 10987
rect 18108 10941 18163 10987
rect 23765 11111 23921 11554
rect 23765 11065 23820 11111
rect 23866 11065 23921 11111
rect 15161 10869 18163 10941
rect 15161 10823 18363 10869
rect 23765 10947 23921 11065
rect 23765 10901 23820 10947
rect 23866 10901 23921 10947
rect 15161 10777 15216 10823
rect 15262 10777 15374 10823
rect 15420 10777 15532 10823
rect 15578 10777 15690 10823
rect 15736 10777 15848 10823
rect 15894 10777 16006 10823
rect 16052 10777 16165 10823
rect 16211 10777 16323 10823
rect 16369 10777 16481 10823
rect 16527 10777 16639 10823
rect 16685 10777 16797 10823
rect 16843 10777 16955 10823
rect 17001 10777 17113 10823
rect 17159 10777 17272 10823
rect 17318 10777 17430 10823
rect 17476 10777 17588 10823
rect 17634 10777 17746 10823
rect 17792 10777 17904 10823
rect 17950 10777 18062 10823
rect 18108 10777 18363 10823
rect 15161 10731 18363 10777
rect 15161 10659 18163 10731
rect 15161 10613 15216 10659
rect 15262 10613 15374 10659
rect 15420 10613 15532 10659
rect 15578 10613 15690 10659
rect 15736 10613 15848 10659
rect 15894 10613 16006 10659
rect 16052 10613 16165 10659
rect 16211 10613 16323 10659
rect 16369 10613 16481 10659
rect 16527 10613 16639 10659
rect 16685 10613 16797 10659
rect 16843 10613 16955 10659
rect 17001 10613 17113 10659
rect 17159 10613 17272 10659
rect 17318 10613 17430 10659
rect 17476 10613 17588 10659
rect 17634 10613 17746 10659
rect 17792 10613 17904 10659
rect 17950 10613 18062 10659
rect 18108 10613 18163 10659
rect 23765 10699 23921 10901
rect 23765 10653 23820 10699
rect 23866 10653 23921 10699
rect 15161 10556 18163 10613
rect 397 10046 553 10163
rect 397 10000 452 10046
rect 498 10000 553 10046
rect 23765 10535 23921 10653
rect 23765 10489 23820 10535
rect 23866 10489 23921 10535
rect 23765 10046 23921 10489
rect 397 9800 553 10000
rect 23765 10000 23820 10046
rect 23866 10000 23921 10046
rect 397 9754 452 9800
rect 498 9754 553 9800
rect 23765 9800 23921 10000
rect 397 9637 553 9754
rect 397 9591 452 9637
rect 498 9591 553 9637
rect 397 9474 553 9591
rect 397 9428 452 9474
rect 498 9428 553 9474
rect 397 9311 553 9428
rect 397 9265 452 9311
rect 498 9265 553 9311
rect 397 9147 553 9265
rect 397 9101 452 9147
rect 498 9101 553 9147
rect 397 8899 553 9101
rect 23765 9754 23820 9800
rect 23866 9754 23921 9800
rect 5945 9023 6458 9069
rect 5945 8977 6086 9023
rect 6320 8977 6458 9023
rect 397 8853 452 8899
rect 498 8853 553 8899
rect 397 8735 553 8853
rect 397 8689 452 8735
rect 498 8689 553 8735
rect 397 8572 553 8689
rect 397 8526 452 8572
rect 498 8526 553 8572
rect 397 8409 553 8526
rect 397 8363 452 8409
rect 498 8363 553 8409
rect 5945 8931 6458 8977
rect 8604 9023 8918 9080
rect 8604 8977 8659 9023
rect 8705 8977 8817 9023
rect 8863 8977 8918 9023
rect 8604 8920 8918 8977
rect 15161 9187 18163 9244
rect 15161 9141 15216 9187
rect 15262 9141 15374 9187
rect 15420 9141 15532 9187
rect 15578 9141 15690 9187
rect 15736 9141 15848 9187
rect 15894 9141 16006 9187
rect 16052 9141 16165 9187
rect 16211 9141 16323 9187
rect 16369 9141 16481 9187
rect 16527 9141 16639 9187
rect 16685 9141 16797 9187
rect 16843 9141 16955 9187
rect 17001 9141 17113 9187
rect 17159 9141 17272 9187
rect 17318 9141 17430 9187
rect 17476 9141 17588 9187
rect 17634 9141 17746 9187
rect 17792 9141 17904 9187
rect 17950 9141 18062 9187
rect 18108 9141 18163 9187
rect 23765 9311 23921 9754
rect 23765 9265 23820 9311
rect 23866 9265 23921 9311
rect 15161 9069 18163 9141
rect 15161 9023 18363 9069
rect 23765 9147 23921 9265
rect 23765 9101 23820 9147
rect 23866 9101 23921 9147
rect 15161 8977 15216 9023
rect 15262 8977 15374 9023
rect 15420 8977 15532 9023
rect 15578 8977 15690 9023
rect 15736 8977 15848 9023
rect 15894 8977 16006 9023
rect 16052 8977 16165 9023
rect 16211 8977 16323 9023
rect 16369 8977 16481 9023
rect 16527 8977 16639 9023
rect 16685 8977 16797 9023
rect 16843 8977 16955 9023
rect 17001 8977 17113 9023
rect 17159 8977 17272 9023
rect 17318 8977 17430 9023
rect 17476 8977 17588 9023
rect 17634 8977 17746 9023
rect 17792 8977 17904 9023
rect 17950 8977 18062 9023
rect 18108 8977 18363 9023
rect 15161 8931 18363 8977
rect 15161 8859 18163 8931
rect 15161 8813 15216 8859
rect 15262 8813 15374 8859
rect 15420 8813 15532 8859
rect 15578 8813 15690 8859
rect 15736 8813 15848 8859
rect 15894 8813 16006 8859
rect 16052 8813 16165 8859
rect 16211 8813 16323 8859
rect 16369 8813 16481 8859
rect 16527 8813 16639 8859
rect 16685 8813 16797 8859
rect 16843 8813 16955 8859
rect 17001 8813 17113 8859
rect 17159 8813 17272 8859
rect 17318 8813 17430 8859
rect 17476 8813 17588 8859
rect 17634 8813 17746 8859
rect 17792 8813 17904 8859
rect 17950 8813 18062 8859
rect 18108 8813 18163 8859
rect 23765 8899 23921 9101
rect 23765 8853 23820 8899
rect 23866 8853 23921 8899
rect 15161 8756 18163 8813
rect 397 8246 553 8363
rect 397 8200 452 8246
rect 498 8200 553 8246
rect 23765 8735 23921 8853
rect 23765 8689 23820 8735
rect 23866 8689 23921 8735
rect 23765 8246 23921 8689
rect 397 8000 553 8200
rect 23765 8200 23820 8246
rect 23866 8200 23921 8246
rect 397 7954 452 8000
rect 498 7954 553 8000
rect 23765 8000 23921 8200
rect 397 7837 553 7954
rect 397 7791 452 7837
rect 498 7791 553 7837
rect 397 7674 553 7791
rect 397 7628 452 7674
rect 498 7628 553 7674
rect 397 7511 553 7628
rect 397 7465 452 7511
rect 498 7465 553 7511
rect 397 7347 553 7465
rect 397 7301 452 7347
rect 498 7301 553 7347
rect 397 7099 553 7301
rect 23765 7954 23820 8000
rect 23866 7954 23921 8000
rect 5945 7223 6458 7269
rect 5945 7177 6086 7223
rect 6320 7177 6458 7223
rect 397 7053 452 7099
rect 498 7053 553 7099
rect 397 6935 553 7053
rect 397 6889 452 6935
rect 498 6889 553 6935
rect 397 6772 553 6889
rect 397 6726 452 6772
rect 498 6726 553 6772
rect 397 6609 553 6726
rect 397 6563 452 6609
rect 498 6563 553 6609
rect 5945 7131 6458 7177
rect 8604 7223 8918 7280
rect 8604 7177 8659 7223
rect 8705 7177 8817 7223
rect 8863 7177 8918 7223
rect 8604 7120 8918 7177
rect 15161 7387 18163 7444
rect 15161 7341 15216 7387
rect 15262 7341 15374 7387
rect 15420 7341 15532 7387
rect 15578 7341 15690 7387
rect 15736 7341 15848 7387
rect 15894 7341 16006 7387
rect 16052 7341 16165 7387
rect 16211 7341 16323 7387
rect 16369 7341 16481 7387
rect 16527 7341 16639 7387
rect 16685 7341 16797 7387
rect 16843 7341 16955 7387
rect 17001 7341 17113 7387
rect 17159 7341 17272 7387
rect 17318 7341 17430 7387
rect 17476 7341 17588 7387
rect 17634 7341 17746 7387
rect 17792 7341 17904 7387
rect 17950 7341 18062 7387
rect 18108 7341 18163 7387
rect 23765 7511 23921 7954
rect 23765 7465 23820 7511
rect 23866 7465 23921 7511
rect 15161 7269 18163 7341
rect 15161 7223 18363 7269
rect 23765 7347 23921 7465
rect 23765 7301 23820 7347
rect 23866 7301 23921 7347
rect 15161 7177 15216 7223
rect 15262 7177 15374 7223
rect 15420 7177 15532 7223
rect 15578 7177 15690 7223
rect 15736 7177 15848 7223
rect 15894 7177 16006 7223
rect 16052 7177 16165 7223
rect 16211 7177 16323 7223
rect 16369 7177 16481 7223
rect 16527 7177 16639 7223
rect 16685 7177 16797 7223
rect 16843 7177 16955 7223
rect 17001 7177 17113 7223
rect 17159 7177 17272 7223
rect 17318 7177 17430 7223
rect 17476 7177 17588 7223
rect 17634 7177 17746 7223
rect 17792 7177 17904 7223
rect 17950 7177 18062 7223
rect 18108 7177 18363 7223
rect 15161 7131 18363 7177
rect 15161 7059 18163 7131
rect 15161 7013 15216 7059
rect 15262 7013 15374 7059
rect 15420 7013 15532 7059
rect 15578 7013 15690 7059
rect 15736 7013 15848 7059
rect 15894 7013 16006 7059
rect 16052 7013 16165 7059
rect 16211 7013 16323 7059
rect 16369 7013 16481 7059
rect 16527 7013 16639 7059
rect 16685 7013 16797 7059
rect 16843 7013 16955 7059
rect 17001 7013 17113 7059
rect 17159 7013 17272 7059
rect 17318 7013 17430 7059
rect 17476 7013 17588 7059
rect 17634 7013 17746 7059
rect 17792 7013 17904 7059
rect 17950 7013 18062 7059
rect 18108 7013 18163 7059
rect 23765 7099 23921 7301
rect 23765 7053 23820 7099
rect 23866 7053 23921 7099
rect 15161 6956 18163 7013
rect 397 6446 553 6563
rect 397 6400 452 6446
rect 498 6400 553 6446
rect 23765 6935 23921 7053
rect 23765 6889 23820 6935
rect 23866 6889 23921 6935
rect 23765 6446 23921 6889
rect 397 6200 553 6400
rect 23765 6400 23820 6446
rect 23866 6400 23921 6446
rect 397 6154 452 6200
rect 498 6154 553 6200
rect 23765 6200 23921 6400
rect 397 6037 553 6154
rect 397 5991 452 6037
rect 498 5991 553 6037
rect 397 5874 553 5991
rect 397 5828 452 5874
rect 498 5828 553 5874
rect 397 5711 553 5828
rect 397 5665 452 5711
rect 498 5665 553 5711
rect 397 5547 553 5665
rect 397 5501 452 5547
rect 498 5501 553 5547
rect 397 5299 553 5501
rect 23765 6154 23820 6200
rect 23866 6154 23921 6200
rect 5945 5423 6458 5469
rect 5945 5377 6086 5423
rect 6320 5377 6458 5423
rect 397 5253 452 5299
rect 498 5253 553 5299
rect 397 5135 553 5253
rect 397 5089 452 5135
rect 498 5089 553 5135
rect 397 4972 553 5089
rect 397 4926 452 4972
rect 498 4926 553 4972
rect 397 4809 553 4926
rect 397 4763 452 4809
rect 498 4763 553 4809
rect 5945 5331 6458 5377
rect 8604 5423 8918 5480
rect 8604 5377 8659 5423
rect 8705 5377 8817 5423
rect 8863 5377 8918 5423
rect 8604 5320 8918 5377
rect 15161 5587 18163 5644
rect 15161 5541 15216 5587
rect 15262 5541 15374 5587
rect 15420 5541 15532 5587
rect 15578 5541 15690 5587
rect 15736 5541 15848 5587
rect 15894 5541 16006 5587
rect 16052 5541 16165 5587
rect 16211 5541 16323 5587
rect 16369 5541 16481 5587
rect 16527 5541 16639 5587
rect 16685 5541 16797 5587
rect 16843 5541 16955 5587
rect 17001 5541 17113 5587
rect 17159 5541 17272 5587
rect 17318 5541 17430 5587
rect 17476 5541 17588 5587
rect 17634 5541 17746 5587
rect 17792 5541 17904 5587
rect 17950 5541 18062 5587
rect 18108 5541 18163 5587
rect 23765 5711 23921 6154
rect 23765 5665 23820 5711
rect 23866 5665 23921 5711
rect 15161 5469 18163 5541
rect 15161 5423 18363 5469
rect 23765 5547 23921 5665
rect 23765 5501 23820 5547
rect 23866 5501 23921 5547
rect 15161 5377 15216 5423
rect 15262 5377 15374 5423
rect 15420 5377 15532 5423
rect 15578 5377 15690 5423
rect 15736 5377 15848 5423
rect 15894 5377 16006 5423
rect 16052 5377 16165 5423
rect 16211 5377 16323 5423
rect 16369 5377 16481 5423
rect 16527 5377 16639 5423
rect 16685 5377 16797 5423
rect 16843 5377 16955 5423
rect 17001 5377 17113 5423
rect 17159 5377 17272 5423
rect 17318 5377 17430 5423
rect 17476 5377 17588 5423
rect 17634 5377 17746 5423
rect 17792 5377 17904 5423
rect 17950 5377 18062 5423
rect 18108 5377 18363 5423
rect 15161 5331 18363 5377
rect 15161 5259 18163 5331
rect 15161 5213 15216 5259
rect 15262 5213 15374 5259
rect 15420 5213 15532 5259
rect 15578 5213 15690 5259
rect 15736 5213 15848 5259
rect 15894 5213 16006 5259
rect 16052 5213 16165 5259
rect 16211 5213 16323 5259
rect 16369 5213 16481 5259
rect 16527 5213 16639 5259
rect 16685 5213 16797 5259
rect 16843 5213 16955 5259
rect 17001 5213 17113 5259
rect 17159 5213 17272 5259
rect 17318 5213 17430 5259
rect 17476 5213 17588 5259
rect 17634 5213 17746 5259
rect 17792 5213 17904 5259
rect 17950 5213 18062 5259
rect 18108 5213 18163 5259
rect 23765 5299 23921 5501
rect 23765 5253 23820 5299
rect 23866 5253 23921 5299
rect 15161 5156 18163 5213
rect 397 4646 553 4763
rect 397 4600 452 4646
rect 498 4600 553 4646
rect 23765 5135 23921 5253
rect 23765 5089 23820 5135
rect 23866 5089 23921 5135
rect 23765 4646 23921 5089
rect 397 4400 553 4600
rect 23765 4600 23820 4646
rect 23866 4600 23921 4646
rect 397 4354 452 4400
rect 498 4354 553 4400
rect 23765 4400 23921 4600
rect 397 4237 553 4354
rect 397 4191 452 4237
rect 498 4191 553 4237
rect 397 4074 553 4191
rect 397 4028 452 4074
rect 498 4028 553 4074
rect 397 3911 553 4028
rect 397 3865 452 3911
rect 498 3865 553 3911
rect 397 3747 553 3865
rect 397 3701 452 3747
rect 498 3701 553 3747
rect 397 3499 553 3701
rect 23765 4354 23820 4400
rect 23866 4354 23921 4400
rect 5945 3623 6458 3669
rect 5945 3577 6086 3623
rect 6320 3577 6458 3623
rect 397 3453 452 3499
rect 498 3453 553 3499
rect 397 3335 553 3453
rect 397 3289 452 3335
rect 498 3289 553 3335
rect 397 3172 553 3289
rect 397 3126 452 3172
rect 498 3126 553 3172
rect 397 3009 553 3126
rect 397 2963 452 3009
rect 498 2963 553 3009
rect 5945 3531 6458 3577
rect 8604 3623 8918 3680
rect 8604 3577 8659 3623
rect 8705 3577 8817 3623
rect 8863 3577 8918 3623
rect 8604 3520 8918 3577
rect 15161 3787 18163 3844
rect 15161 3741 15216 3787
rect 15262 3741 15374 3787
rect 15420 3741 15532 3787
rect 15578 3741 15690 3787
rect 15736 3741 15848 3787
rect 15894 3741 16006 3787
rect 16052 3741 16165 3787
rect 16211 3741 16323 3787
rect 16369 3741 16481 3787
rect 16527 3741 16639 3787
rect 16685 3741 16797 3787
rect 16843 3741 16955 3787
rect 17001 3741 17113 3787
rect 17159 3741 17272 3787
rect 17318 3741 17430 3787
rect 17476 3741 17588 3787
rect 17634 3741 17746 3787
rect 17792 3741 17904 3787
rect 17950 3741 18062 3787
rect 18108 3741 18163 3787
rect 23765 3911 23921 4354
rect 23765 3865 23820 3911
rect 23866 3865 23921 3911
rect 15161 3669 18163 3741
rect 15161 3623 18363 3669
rect 23765 3747 23921 3865
rect 23765 3701 23820 3747
rect 23866 3701 23921 3747
rect 15161 3577 15216 3623
rect 15262 3577 15374 3623
rect 15420 3577 15532 3623
rect 15578 3577 15690 3623
rect 15736 3577 15848 3623
rect 15894 3577 16006 3623
rect 16052 3577 16165 3623
rect 16211 3577 16323 3623
rect 16369 3577 16481 3623
rect 16527 3577 16639 3623
rect 16685 3577 16797 3623
rect 16843 3577 16955 3623
rect 17001 3577 17113 3623
rect 17159 3577 17272 3623
rect 17318 3577 17430 3623
rect 17476 3577 17588 3623
rect 17634 3577 17746 3623
rect 17792 3577 17904 3623
rect 17950 3577 18062 3623
rect 18108 3577 18363 3623
rect 15161 3531 18363 3577
rect 15161 3459 18163 3531
rect 15161 3413 15216 3459
rect 15262 3413 15374 3459
rect 15420 3413 15532 3459
rect 15578 3413 15690 3459
rect 15736 3413 15848 3459
rect 15894 3413 16006 3459
rect 16052 3413 16165 3459
rect 16211 3413 16323 3459
rect 16369 3413 16481 3459
rect 16527 3413 16639 3459
rect 16685 3413 16797 3459
rect 16843 3413 16955 3459
rect 17001 3413 17113 3459
rect 17159 3413 17272 3459
rect 17318 3413 17430 3459
rect 17476 3413 17588 3459
rect 17634 3413 17746 3459
rect 17792 3413 17904 3459
rect 17950 3413 18062 3459
rect 18108 3413 18163 3459
rect 23765 3499 23921 3701
rect 23765 3453 23820 3499
rect 23866 3453 23921 3499
rect 15161 3356 18163 3413
rect 397 2846 553 2963
rect 397 2800 452 2846
rect 498 2800 553 2846
rect 23765 3335 23921 3453
rect 23765 3289 23820 3335
rect 23866 3289 23921 3335
rect 23765 2846 23921 3289
rect 397 2600 553 2800
rect 23765 2800 23820 2846
rect 23866 2800 23921 2846
rect 397 2554 452 2600
rect 498 2554 553 2600
rect 23765 2600 23921 2800
rect 397 2437 553 2554
rect 397 2391 452 2437
rect 498 2391 553 2437
rect 397 2274 553 2391
rect 397 2228 452 2274
rect 498 2228 553 2274
rect 397 2111 553 2228
rect 397 2065 452 2111
rect 498 2065 553 2111
rect 397 1947 553 2065
rect 397 1901 452 1947
rect 498 1901 553 1947
rect 397 1699 553 1901
rect 23765 2554 23820 2600
rect 23866 2554 23921 2600
rect 5945 1823 6458 1869
rect 5945 1777 6086 1823
rect 6320 1777 6458 1823
rect 397 1653 452 1699
rect 498 1653 553 1699
rect 397 1535 553 1653
rect 397 1489 452 1535
rect 498 1489 553 1535
rect 397 1372 553 1489
rect 397 1326 452 1372
rect 498 1326 553 1372
rect 397 1209 553 1326
rect 397 1163 452 1209
rect 498 1163 553 1209
rect 5945 1731 6458 1777
rect 8604 1823 8918 1880
rect 8604 1777 8659 1823
rect 8705 1777 8817 1823
rect 8863 1777 8918 1823
rect 8604 1720 8918 1777
rect 15161 1987 18163 2044
rect 15161 1941 15216 1987
rect 15262 1941 15374 1987
rect 15420 1941 15532 1987
rect 15578 1941 15690 1987
rect 15736 1941 15848 1987
rect 15894 1941 16006 1987
rect 16052 1941 16165 1987
rect 16211 1941 16323 1987
rect 16369 1941 16481 1987
rect 16527 1941 16639 1987
rect 16685 1941 16797 1987
rect 16843 1941 16955 1987
rect 17001 1941 17113 1987
rect 17159 1941 17272 1987
rect 17318 1941 17430 1987
rect 17476 1941 17588 1987
rect 17634 1941 17746 1987
rect 17792 1941 17904 1987
rect 17950 1941 18062 1987
rect 18108 1941 18163 1987
rect 23765 2111 23921 2554
rect 23765 2065 23820 2111
rect 23866 2065 23921 2111
rect 15161 1869 18163 1941
rect 15161 1823 18363 1869
rect 23765 1947 23921 2065
rect 23765 1901 23820 1947
rect 23866 1901 23921 1947
rect 15161 1777 15216 1823
rect 15262 1777 15374 1823
rect 15420 1777 15532 1823
rect 15578 1777 15690 1823
rect 15736 1777 15848 1823
rect 15894 1777 16006 1823
rect 16052 1777 16165 1823
rect 16211 1777 16323 1823
rect 16369 1777 16481 1823
rect 16527 1777 16639 1823
rect 16685 1777 16797 1823
rect 16843 1777 16955 1823
rect 17001 1777 17113 1823
rect 17159 1777 17272 1823
rect 17318 1777 17430 1823
rect 17476 1777 17588 1823
rect 17634 1777 17746 1823
rect 17792 1777 17904 1823
rect 17950 1777 18062 1823
rect 18108 1777 18363 1823
rect 15161 1731 18363 1777
rect 15161 1659 18163 1731
rect 15161 1613 15216 1659
rect 15262 1613 15374 1659
rect 15420 1613 15532 1659
rect 15578 1613 15690 1659
rect 15736 1613 15848 1659
rect 15894 1613 16006 1659
rect 16052 1613 16165 1659
rect 16211 1613 16323 1659
rect 16369 1613 16481 1659
rect 16527 1613 16639 1659
rect 16685 1613 16797 1659
rect 16843 1613 16955 1659
rect 17001 1613 17113 1659
rect 17159 1613 17272 1659
rect 17318 1613 17430 1659
rect 17476 1613 17588 1659
rect 17634 1613 17746 1659
rect 17792 1613 17904 1659
rect 17950 1613 18062 1659
rect 18108 1613 18163 1659
rect 23765 1699 23921 1901
rect 23765 1653 23820 1699
rect 23866 1653 23921 1699
rect 15161 1556 18163 1613
rect 397 1046 553 1163
rect 397 1000 452 1046
rect 498 1000 553 1046
rect 23765 1535 23921 1653
rect 23765 1489 23820 1535
rect 23866 1489 23921 1535
rect 23765 1046 23921 1489
rect 397 800 553 1000
rect 23765 1000 23820 1046
rect 23866 1000 23921 1046
rect 397 754 452 800
rect 498 754 553 800
rect 23765 800 23921 1000
rect 397 637 553 754
rect 397 591 452 637
rect 498 591 553 637
rect 397 474 553 591
rect 397 428 452 474
rect 498 428 553 474
rect 397 311 553 428
rect 397 265 452 311
rect 498 265 553 311
rect 397 147 553 265
rect 397 101 452 147
rect 498 101 553 147
rect 397 -62 553 101
rect 23765 754 23820 800
rect 23866 754 23921 800
rect 5945 23 6458 69
rect 5945 -23 6086 23
rect 6320 -23 6458 23
rect 5945 -69 6458 -23
rect 8604 23 8918 80
rect 8604 -23 8659 23
rect 8705 -23 8817 23
rect 8863 -23 8918 23
rect 8604 -80 8918 -23
rect 15161 187 18163 244
rect 15161 141 15216 187
rect 15262 141 15374 187
rect 15420 141 15532 187
rect 15578 141 15690 187
rect 15736 141 15848 187
rect 15894 141 16006 187
rect 16052 141 16165 187
rect 16211 141 16323 187
rect 16369 141 16481 187
rect 16527 141 16639 187
rect 16685 141 16797 187
rect 16843 141 16955 187
rect 17001 141 17113 187
rect 17159 141 17272 187
rect 17318 141 17430 187
rect 17476 141 17588 187
rect 17634 141 17746 187
rect 17792 141 17904 187
rect 17950 141 18062 187
rect 18108 141 18163 187
rect 23765 311 23921 754
rect 23765 265 23820 311
rect 23866 265 23921 311
rect 15161 69 18163 141
rect 15161 23 18363 69
rect 23765 147 23921 265
rect 23765 101 23820 147
rect 23866 101 23921 147
rect 15161 -23 15216 23
rect 15262 -23 15374 23
rect 15420 -23 15532 23
rect 15578 -23 15690 23
rect 15736 -23 15848 23
rect 15894 -23 16006 23
rect 16052 -23 16165 23
rect 16211 -23 16323 23
rect 16369 -23 16481 23
rect 16527 -23 16639 23
rect 16685 -23 16797 23
rect 16843 -23 16955 23
rect 17001 -23 17113 23
rect 17159 -23 17272 23
rect 17318 -23 17430 23
rect 17476 -23 17588 23
rect 17634 -23 17746 23
rect 17792 -23 17904 23
rect 17950 -23 18062 23
rect 18108 -23 18363 23
rect 15161 -69 18363 -23
rect 23765 -62 23921 101
rect 15161 -80 18163 -69
<< psubdiffcont >>
rect 7554 14377 8070 14423
rect 10433 14377 10479 14423
rect 10591 14377 10637 14423
rect 10749 14377 10795 14423
rect 10907 14377 10953 14423
rect 11066 14377 11112 14423
rect 11224 14377 11270 14423
rect 11382 14377 11428 14423
rect 11540 14377 11586 14423
rect 11698 14377 11744 14423
rect 11856 14377 11902 14423
rect 12015 14377 12061 14423
rect 12173 14377 12219 14423
rect 12331 14377 12377 14423
rect 12489 14377 12535 14423
rect 4513 13477 4559 13523
rect 19757 13477 19803 13523
rect 7554 12577 8070 12623
rect 10433 12577 10479 12623
rect 10591 12577 10637 12623
rect 10749 12577 10795 12623
rect 10907 12577 10953 12623
rect 11066 12577 11112 12623
rect 11224 12577 11270 12623
rect 11382 12577 11428 12623
rect 11540 12577 11586 12623
rect 11698 12577 11744 12623
rect 11856 12577 11902 12623
rect 12015 12577 12061 12623
rect 12173 12577 12219 12623
rect 12331 12577 12377 12623
rect 12489 12577 12535 12623
rect 4513 11677 4559 11723
rect 19757 11677 19803 11723
rect 7554 10777 8070 10823
rect 10433 10777 10479 10823
rect 10591 10777 10637 10823
rect 10749 10777 10795 10823
rect 10907 10777 10953 10823
rect 11066 10777 11112 10823
rect 11224 10777 11270 10823
rect 11382 10777 11428 10823
rect 11540 10777 11586 10823
rect 11698 10777 11744 10823
rect 11856 10777 11902 10823
rect 12015 10777 12061 10823
rect 12173 10777 12219 10823
rect 12331 10777 12377 10823
rect 12489 10777 12535 10823
rect 4513 9877 4559 9923
rect 19757 9877 19803 9923
rect 7554 8977 8070 9023
rect 10433 8977 10479 9023
rect 10591 8977 10637 9023
rect 10749 8977 10795 9023
rect 10907 8977 10953 9023
rect 11066 8977 11112 9023
rect 11224 8977 11270 9023
rect 11382 8977 11428 9023
rect 11540 8977 11586 9023
rect 11698 8977 11744 9023
rect 11856 8977 11902 9023
rect 12015 8977 12061 9023
rect 12173 8977 12219 9023
rect 12331 8977 12377 9023
rect 12489 8977 12535 9023
rect 4513 8077 4559 8123
rect 19757 8077 19803 8123
rect 7554 7177 8070 7223
rect 10433 7177 10479 7223
rect 10591 7177 10637 7223
rect 10749 7177 10795 7223
rect 10907 7177 10953 7223
rect 11066 7177 11112 7223
rect 11224 7177 11270 7223
rect 11382 7177 11428 7223
rect 11540 7177 11586 7223
rect 11698 7177 11744 7223
rect 11856 7177 11902 7223
rect 12015 7177 12061 7223
rect 12173 7177 12219 7223
rect 12331 7177 12377 7223
rect 12489 7177 12535 7223
rect 4513 6277 4559 6323
rect 19757 6277 19803 6323
rect 7554 5377 8070 5423
rect 10433 5377 10479 5423
rect 10591 5377 10637 5423
rect 10749 5377 10795 5423
rect 10907 5377 10953 5423
rect 11066 5377 11112 5423
rect 11224 5377 11270 5423
rect 11382 5377 11428 5423
rect 11540 5377 11586 5423
rect 11698 5377 11744 5423
rect 11856 5377 11902 5423
rect 12015 5377 12061 5423
rect 12173 5377 12219 5423
rect 12331 5377 12377 5423
rect 12489 5377 12535 5423
rect 4513 4477 4559 4523
rect 19757 4477 19803 4523
rect 7554 3577 8070 3623
rect 10433 3577 10479 3623
rect 10591 3577 10637 3623
rect 10749 3577 10795 3623
rect 10907 3577 10953 3623
rect 11066 3577 11112 3623
rect 11224 3577 11270 3623
rect 11382 3577 11428 3623
rect 11540 3577 11586 3623
rect 11698 3577 11744 3623
rect 11856 3577 11902 3623
rect 12015 3577 12061 3623
rect 12173 3577 12219 3623
rect 12331 3577 12377 3623
rect 12489 3577 12535 3623
rect 4513 2677 4559 2723
rect 19757 2677 19803 2723
rect 7554 1777 8070 1823
rect 10433 1777 10479 1823
rect 10591 1777 10637 1823
rect 10749 1777 10795 1823
rect 10907 1777 10953 1823
rect 11066 1777 11112 1823
rect 11224 1777 11270 1823
rect 11382 1777 11428 1823
rect 11540 1777 11586 1823
rect 11698 1777 11744 1823
rect 11856 1777 11902 1823
rect 12015 1777 12061 1823
rect 12173 1777 12219 1823
rect 12331 1777 12377 1823
rect 12489 1777 12535 1823
rect 4513 877 4559 923
rect 19757 877 19803 923
rect 7554 -23 8070 23
rect 10433 -23 10479 23
rect 10591 -23 10637 23
rect 10749 -23 10795 23
rect 10907 -23 10953 23
rect 11066 -23 11112 23
rect 11224 -23 11270 23
rect 11382 -23 11428 23
rect 11540 -23 11586 23
rect 11698 -23 11744 23
rect 11856 -23 11902 23
rect 12015 -23 12061 23
rect 12173 -23 12219 23
rect 12331 -23 12377 23
rect 12489 -23 12535 23
<< nsubdiffcont >>
rect 6086 14377 6320 14423
rect 452 14253 498 14299
rect 452 14089 498 14135
rect 452 13926 498 13972
rect 452 13763 498 13809
rect 8659 14377 8705 14423
rect 8817 14377 8863 14423
rect 15216 14377 15262 14423
rect 15374 14377 15420 14423
rect 15532 14377 15578 14423
rect 15690 14377 15736 14423
rect 15848 14377 15894 14423
rect 16006 14377 16052 14423
rect 16165 14377 16211 14423
rect 16323 14377 16369 14423
rect 16481 14377 16527 14423
rect 16639 14377 16685 14423
rect 16797 14377 16843 14423
rect 16955 14377 17001 14423
rect 17113 14377 17159 14423
rect 17272 14377 17318 14423
rect 17430 14377 17476 14423
rect 17588 14377 17634 14423
rect 17746 14377 17792 14423
rect 17904 14377 17950 14423
rect 18062 14377 18108 14423
rect 15216 14213 15262 14259
rect 15374 14213 15420 14259
rect 15532 14213 15578 14259
rect 15690 14213 15736 14259
rect 15848 14213 15894 14259
rect 16006 14213 16052 14259
rect 16165 14213 16211 14259
rect 16323 14213 16369 14259
rect 16481 14213 16527 14259
rect 16639 14213 16685 14259
rect 16797 14213 16843 14259
rect 16955 14213 17001 14259
rect 17113 14213 17159 14259
rect 17272 14213 17318 14259
rect 17430 14213 17476 14259
rect 17588 14213 17634 14259
rect 17746 14213 17792 14259
rect 17904 14213 17950 14259
rect 18062 14213 18108 14259
rect 23820 14253 23866 14299
rect 452 13600 498 13646
rect 23820 14089 23866 14135
rect 23820 13600 23866 13646
rect 452 13354 498 13400
rect 452 13191 498 13237
rect 452 13028 498 13074
rect 452 12865 498 12911
rect 452 12701 498 12747
rect 23820 13354 23866 13400
rect 6086 12577 6320 12623
rect 452 12453 498 12499
rect 452 12289 498 12335
rect 452 12126 498 12172
rect 452 11963 498 12009
rect 8659 12577 8705 12623
rect 8817 12577 8863 12623
rect 15216 12741 15262 12787
rect 15374 12741 15420 12787
rect 15532 12741 15578 12787
rect 15690 12741 15736 12787
rect 15848 12741 15894 12787
rect 16006 12741 16052 12787
rect 16165 12741 16211 12787
rect 16323 12741 16369 12787
rect 16481 12741 16527 12787
rect 16639 12741 16685 12787
rect 16797 12741 16843 12787
rect 16955 12741 17001 12787
rect 17113 12741 17159 12787
rect 17272 12741 17318 12787
rect 17430 12741 17476 12787
rect 17588 12741 17634 12787
rect 17746 12741 17792 12787
rect 17904 12741 17950 12787
rect 18062 12741 18108 12787
rect 23820 12865 23866 12911
rect 23820 12701 23866 12747
rect 15216 12577 15262 12623
rect 15374 12577 15420 12623
rect 15532 12577 15578 12623
rect 15690 12577 15736 12623
rect 15848 12577 15894 12623
rect 16006 12577 16052 12623
rect 16165 12577 16211 12623
rect 16323 12577 16369 12623
rect 16481 12577 16527 12623
rect 16639 12577 16685 12623
rect 16797 12577 16843 12623
rect 16955 12577 17001 12623
rect 17113 12577 17159 12623
rect 17272 12577 17318 12623
rect 17430 12577 17476 12623
rect 17588 12577 17634 12623
rect 17746 12577 17792 12623
rect 17904 12577 17950 12623
rect 18062 12577 18108 12623
rect 15216 12413 15262 12459
rect 15374 12413 15420 12459
rect 15532 12413 15578 12459
rect 15690 12413 15736 12459
rect 15848 12413 15894 12459
rect 16006 12413 16052 12459
rect 16165 12413 16211 12459
rect 16323 12413 16369 12459
rect 16481 12413 16527 12459
rect 16639 12413 16685 12459
rect 16797 12413 16843 12459
rect 16955 12413 17001 12459
rect 17113 12413 17159 12459
rect 17272 12413 17318 12459
rect 17430 12413 17476 12459
rect 17588 12413 17634 12459
rect 17746 12413 17792 12459
rect 17904 12413 17950 12459
rect 18062 12413 18108 12459
rect 23820 12453 23866 12499
rect 452 11800 498 11846
rect 23820 12289 23866 12335
rect 23820 11800 23866 11846
rect 452 11554 498 11600
rect 452 11391 498 11437
rect 452 11228 498 11274
rect 452 11065 498 11111
rect 452 10901 498 10947
rect 23820 11554 23866 11600
rect 6086 10777 6320 10823
rect 452 10653 498 10699
rect 452 10489 498 10535
rect 452 10326 498 10372
rect 452 10163 498 10209
rect 8659 10777 8705 10823
rect 8817 10777 8863 10823
rect 15216 10941 15262 10987
rect 15374 10941 15420 10987
rect 15532 10941 15578 10987
rect 15690 10941 15736 10987
rect 15848 10941 15894 10987
rect 16006 10941 16052 10987
rect 16165 10941 16211 10987
rect 16323 10941 16369 10987
rect 16481 10941 16527 10987
rect 16639 10941 16685 10987
rect 16797 10941 16843 10987
rect 16955 10941 17001 10987
rect 17113 10941 17159 10987
rect 17272 10941 17318 10987
rect 17430 10941 17476 10987
rect 17588 10941 17634 10987
rect 17746 10941 17792 10987
rect 17904 10941 17950 10987
rect 18062 10941 18108 10987
rect 23820 11065 23866 11111
rect 23820 10901 23866 10947
rect 15216 10777 15262 10823
rect 15374 10777 15420 10823
rect 15532 10777 15578 10823
rect 15690 10777 15736 10823
rect 15848 10777 15894 10823
rect 16006 10777 16052 10823
rect 16165 10777 16211 10823
rect 16323 10777 16369 10823
rect 16481 10777 16527 10823
rect 16639 10777 16685 10823
rect 16797 10777 16843 10823
rect 16955 10777 17001 10823
rect 17113 10777 17159 10823
rect 17272 10777 17318 10823
rect 17430 10777 17476 10823
rect 17588 10777 17634 10823
rect 17746 10777 17792 10823
rect 17904 10777 17950 10823
rect 18062 10777 18108 10823
rect 15216 10613 15262 10659
rect 15374 10613 15420 10659
rect 15532 10613 15578 10659
rect 15690 10613 15736 10659
rect 15848 10613 15894 10659
rect 16006 10613 16052 10659
rect 16165 10613 16211 10659
rect 16323 10613 16369 10659
rect 16481 10613 16527 10659
rect 16639 10613 16685 10659
rect 16797 10613 16843 10659
rect 16955 10613 17001 10659
rect 17113 10613 17159 10659
rect 17272 10613 17318 10659
rect 17430 10613 17476 10659
rect 17588 10613 17634 10659
rect 17746 10613 17792 10659
rect 17904 10613 17950 10659
rect 18062 10613 18108 10659
rect 23820 10653 23866 10699
rect 452 10000 498 10046
rect 23820 10489 23866 10535
rect 23820 10000 23866 10046
rect 452 9754 498 9800
rect 452 9591 498 9637
rect 452 9428 498 9474
rect 452 9265 498 9311
rect 452 9101 498 9147
rect 23820 9754 23866 9800
rect 6086 8977 6320 9023
rect 452 8853 498 8899
rect 452 8689 498 8735
rect 452 8526 498 8572
rect 452 8363 498 8409
rect 8659 8977 8705 9023
rect 8817 8977 8863 9023
rect 15216 9141 15262 9187
rect 15374 9141 15420 9187
rect 15532 9141 15578 9187
rect 15690 9141 15736 9187
rect 15848 9141 15894 9187
rect 16006 9141 16052 9187
rect 16165 9141 16211 9187
rect 16323 9141 16369 9187
rect 16481 9141 16527 9187
rect 16639 9141 16685 9187
rect 16797 9141 16843 9187
rect 16955 9141 17001 9187
rect 17113 9141 17159 9187
rect 17272 9141 17318 9187
rect 17430 9141 17476 9187
rect 17588 9141 17634 9187
rect 17746 9141 17792 9187
rect 17904 9141 17950 9187
rect 18062 9141 18108 9187
rect 23820 9265 23866 9311
rect 23820 9101 23866 9147
rect 15216 8977 15262 9023
rect 15374 8977 15420 9023
rect 15532 8977 15578 9023
rect 15690 8977 15736 9023
rect 15848 8977 15894 9023
rect 16006 8977 16052 9023
rect 16165 8977 16211 9023
rect 16323 8977 16369 9023
rect 16481 8977 16527 9023
rect 16639 8977 16685 9023
rect 16797 8977 16843 9023
rect 16955 8977 17001 9023
rect 17113 8977 17159 9023
rect 17272 8977 17318 9023
rect 17430 8977 17476 9023
rect 17588 8977 17634 9023
rect 17746 8977 17792 9023
rect 17904 8977 17950 9023
rect 18062 8977 18108 9023
rect 15216 8813 15262 8859
rect 15374 8813 15420 8859
rect 15532 8813 15578 8859
rect 15690 8813 15736 8859
rect 15848 8813 15894 8859
rect 16006 8813 16052 8859
rect 16165 8813 16211 8859
rect 16323 8813 16369 8859
rect 16481 8813 16527 8859
rect 16639 8813 16685 8859
rect 16797 8813 16843 8859
rect 16955 8813 17001 8859
rect 17113 8813 17159 8859
rect 17272 8813 17318 8859
rect 17430 8813 17476 8859
rect 17588 8813 17634 8859
rect 17746 8813 17792 8859
rect 17904 8813 17950 8859
rect 18062 8813 18108 8859
rect 23820 8853 23866 8899
rect 452 8200 498 8246
rect 23820 8689 23866 8735
rect 23820 8200 23866 8246
rect 452 7954 498 8000
rect 452 7791 498 7837
rect 452 7628 498 7674
rect 452 7465 498 7511
rect 452 7301 498 7347
rect 23820 7954 23866 8000
rect 6086 7177 6320 7223
rect 452 7053 498 7099
rect 452 6889 498 6935
rect 452 6726 498 6772
rect 452 6563 498 6609
rect 8659 7177 8705 7223
rect 8817 7177 8863 7223
rect 15216 7341 15262 7387
rect 15374 7341 15420 7387
rect 15532 7341 15578 7387
rect 15690 7341 15736 7387
rect 15848 7341 15894 7387
rect 16006 7341 16052 7387
rect 16165 7341 16211 7387
rect 16323 7341 16369 7387
rect 16481 7341 16527 7387
rect 16639 7341 16685 7387
rect 16797 7341 16843 7387
rect 16955 7341 17001 7387
rect 17113 7341 17159 7387
rect 17272 7341 17318 7387
rect 17430 7341 17476 7387
rect 17588 7341 17634 7387
rect 17746 7341 17792 7387
rect 17904 7341 17950 7387
rect 18062 7341 18108 7387
rect 23820 7465 23866 7511
rect 23820 7301 23866 7347
rect 15216 7177 15262 7223
rect 15374 7177 15420 7223
rect 15532 7177 15578 7223
rect 15690 7177 15736 7223
rect 15848 7177 15894 7223
rect 16006 7177 16052 7223
rect 16165 7177 16211 7223
rect 16323 7177 16369 7223
rect 16481 7177 16527 7223
rect 16639 7177 16685 7223
rect 16797 7177 16843 7223
rect 16955 7177 17001 7223
rect 17113 7177 17159 7223
rect 17272 7177 17318 7223
rect 17430 7177 17476 7223
rect 17588 7177 17634 7223
rect 17746 7177 17792 7223
rect 17904 7177 17950 7223
rect 18062 7177 18108 7223
rect 15216 7013 15262 7059
rect 15374 7013 15420 7059
rect 15532 7013 15578 7059
rect 15690 7013 15736 7059
rect 15848 7013 15894 7059
rect 16006 7013 16052 7059
rect 16165 7013 16211 7059
rect 16323 7013 16369 7059
rect 16481 7013 16527 7059
rect 16639 7013 16685 7059
rect 16797 7013 16843 7059
rect 16955 7013 17001 7059
rect 17113 7013 17159 7059
rect 17272 7013 17318 7059
rect 17430 7013 17476 7059
rect 17588 7013 17634 7059
rect 17746 7013 17792 7059
rect 17904 7013 17950 7059
rect 18062 7013 18108 7059
rect 23820 7053 23866 7099
rect 452 6400 498 6446
rect 23820 6889 23866 6935
rect 23820 6400 23866 6446
rect 452 6154 498 6200
rect 452 5991 498 6037
rect 452 5828 498 5874
rect 452 5665 498 5711
rect 452 5501 498 5547
rect 23820 6154 23866 6200
rect 6086 5377 6320 5423
rect 452 5253 498 5299
rect 452 5089 498 5135
rect 452 4926 498 4972
rect 452 4763 498 4809
rect 8659 5377 8705 5423
rect 8817 5377 8863 5423
rect 15216 5541 15262 5587
rect 15374 5541 15420 5587
rect 15532 5541 15578 5587
rect 15690 5541 15736 5587
rect 15848 5541 15894 5587
rect 16006 5541 16052 5587
rect 16165 5541 16211 5587
rect 16323 5541 16369 5587
rect 16481 5541 16527 5587
rect 16639 5541 16685 5587
rect 16797 5541 16843 5587
rect 16955 5541 17001 5587
rect 17113 5541 17159 5587
rect 17272 5541 17318 5587
rect 17430 5541 17476 5587
rect 17588 5541 17634 5587
rect 17746 5541 17792 5587
rect 17904 5541 17950 5587
rect 18062 5541 18108 5587
rect 23820 5665 23866 5711
rect 23820 5501 23866 5547
rect 15216 5377 15262 5423
rect 15374 5377 15420 5423
rect 15532 5377 15578 5423
rect 15690 5377 15736 5423
rect 15848 5377 15894 5423
rect 16006 5377 16052 5423
rect 16165 5377 16211 5423
rect 16323 5377 16369 5423
rect 16481 5377 16527 5423
rect 16639 5377 16685 5423
rect 16797 5377 16843 5423
rect 16955 5377 17001 5423
rect 17113 5377 17159 5423
rect 17272 5377 17318 5423
rect 17430 5377 17476 5423
rect 17588 5377 17634 5423
rect 17746 5377 17792 5423
rect 17904 5377 17950 5423
rect 18062 5377 18108 5423
rect 15216 5213 15262 5259
rect 15374 5213 15420 5259
rect 15532 5213 15578 5259
rect 15690 5213 15736 5259
rect 15848 5213 15894 5259
rect 16006 5213 16052 5259
rect 16165 5213 16211 5259
rect 16323 5213 16369 5259
rect 16481 5213 16527 5259
rect 16639 5213 16685 5259
rect 16797 5213 16843 5259
rect 16955 5213 17001 5259
rect 17113 5213 17159 5259
rect 17272 5213 17318 5259
rect 17430 5213 17476 5259
rect 17588 5213 17634 5259
rect 17746 5213 17792 5259
rect 17904 5213 17950 5259
rect 18062 5213 18108 5259
rect 23820 5253 23866 5299
rect 452 4600 498 4646
rect 23820 5089 23866 5135
rect 23820 4600 23866 4646
rect 452 4354 498 4400
rect 452 4191 498 4237
rect 452 4028 498 4074
rect 452 3865 498 3911
rect 452 3701 498 3747
rect 23820 4354 23866 4400
rect 6086 3577 6320 3623
rect 452 3453 498 3499
rect 452 3289 498 3335
rect 452 3126 498 3172
rect 452 2963 498 3009
rect 8659 3577 8705 3623
rect 8817 3577 8863 3623
rect 15216 3741 15262 3787
rect 15374 3741 15420 3787
rect 15532 3741 15578 3787
rect 15690 3741 15736 3787
rect 15848 3741 15894 3787
rect 16006 3741 16052 3787
rect 16165 3741 16211 3787
rect 16323 3741 16369 3787
rect 16481 3741 16527 3787
rect 16639 3741 16685 3787
rect 16797 3741 16843 3787
rect 16955 3741 17001 3787
rect 17113 3741 17159 3787
rect 17272 3741 17318 3787
rect 17430 3741 17476 3787
rect 17588 3741 17634 3787
rect 17746 3741 17792 3787
rect 17904 3741 17950 3787
rect 18062 3741 18108 3787
rect 23820 3865 23866 3911
rect 23820 3701 23866 3747
rect 15216 3577 15262 3623
rect 15374 3577 15420 3623
rect 15532 3577 15578 3623
rect 15690 3577 15736 3623
rect 15848 3577 15894 3623
rect 16006 3577 16052 3623
rect 16165 3577 16211 3623
rect 16323 3577 16369 3623
rect 16481 3577 16527 3623
rect 16639 3577 16685 3623
rect 16797 3577 16843 3623
rect 16955 3577 17001 3623
rect 17113 3577 17159 3623
rect 17272 3577 17318 3623
rect 17430 3577 17476 3623
rect 17588 3577 17634 3623
rect 17746 3577 17792 3623
rect 17904 3577 17950 3623
rect 18062 3577 18108 3623
rect 15216 3413 15262 3459
rect 15374 3413 15420 3459
rect 15532 3413 15578 3459
rect 15690 3413 15736 3459
rect 15848 3413 15894 3459
rect 16006 3413 16052 3459
rect 16165 3413 16211 3459
rect 16323 3413 16369 3459
rect 16481 3413 16527 3459
rect 16639 3413 16685 3459
rect 16797 3413 16843 3459
rect 16955 3413 17001 3459
rect 17113 3413 17159 3459
rect 17272 3413 17318 3459
rect 17430 3413 17476 3459
rect 17588 3413 17634 3459
rect 17746 3413 17792 3459
rect 17904 3413 17950 3459
rect 18062 3413 18108 3459
rect 23820 3453 23866 3499
rect 452 2800 498 2846
rect 23820 3289 23866 3335
rect 23820 2800 23866 2846
rect 452 2554 498 2600
rect 452 2391 498 2437
rect 452 2228 498 2274
rect 452 2065 498 2111
rect 452 1901 498 1947
rect 23820 2554 23866 2600
rect 6086 1777 6320 1823
rect 452 1653 498 1699
rect 452 1489 498 1535
rect 452 1326 498 1372
rect 452 1163 498 1209
rect 8659 1777 8705 1823
rect 8817 1777 8863 1823
rect 15216 1941 15262 1987
rect 15374 1941 15420 1987
rect 15532 1941 15578 1987
rect 15690 1941 15736 1987
rect 15848 1941 15894 1987
rect 16006 1941 16052 1987
rect 16165 1941 16211 1987
rect 16323 1941 16369 1987
rect 16481 1941 16527 1987
rect 16639 1941 16685 1987
rect 16797 1941 16843 1987
rect 16955 1941 17001 1987
rect 17113 1941 17159 1987
rect 17272 1941 17318 1987
rect 17430 1941 17476 1987
rect 17588 1941 17634 1987
rect 17746 1941 17792 1987
rect 17904 1941 17950 1987
rect 18062 1941 18108 1987
rect 23820 2065 23866 2111
rect 23820 1901 23866 1947
rect 15216 1777 15262 1823
rect 15374 1777 15420 1823
rect 15532 1777 15578 1823
rect 15690 1777 15736 1823
rect 15848 1777 15894 1823
rect 16006 1777 16052 1823
rect 16165 1777 16211 1823
rect 16323 1777 16369 1823
rect 16481 1777 16527 1823
rect 16639 1777 16685 1823
rect 16797 1777 16843 1823
rect 16955 1777 17001 1823
rect 17113 1777 17159 1823
rect 17272 1777 17318 1823
rect 17430 1777 17476 1823
rect 17588 1777 17634 1823
rect 17746 1777 17792 1823
rect 17904 1777 17950 1823
rect 18062 1777 18108 1823
rect 15216 1613 15262 1659
rect 15374 1613 15420 1659
rect 15532 1613 15578 1659
rect 15690 1613 15736 1659
rect 15848 1613 15894 1659
rect 16006 1613 16052 1659
rect 16165 1613 16211 1659
rect 16323 1613 16369 1659
rect 16481 1613 16527 1659
rect 16639 1613 16685 1659
rect 16797 1613 16843 1659
rect 16955 1613 17001 1659
rect 17113 1613 17159 1659
rect 17272 1613 17318 1659
rect 17430 1613 17476 1659
rect 17588 1613 17634 1659
rect 17746 1613 17792 1659
rect 17904 1613 17950 1659
rect 18062 1613 18108 1659
rect 23820 1653 23866 1699
rect 452 1000 498 1046
rect 23820 1489 23866 1535
rect 23820 1000 23866 1046
rect 452 754 498 800
rect 452 591 498 637
rect 452 428 498 474
rect 452 265 498 311
rect 452 101 498 147
rect 23820 754 23866 800
rect 6086 -23 6320 23
rect 8659 -23 8705 23
rect 8817 -23 8863 23
rect 15216 141 15262 187
rect 15374 141 15420 187
rect 15532 141 15578 187
rect 15690 141 15736 187
rect 15848 141 15894 187
rect 16006 141 16052 187
rect 16165 141 16211 187
rect 16323 141 16369 187
rect 16481 141 16527 187
rect 16639 141 16685 187
rect 16797 141 16843 187
rect 16955 141 17001 187
rect 17113 141 17159 187
rect 17272 141 17318 187
rect 17430 141 17476 187
rect 17588 141 17634 187
rect 17746 141 17792 187
rect 17904 141 17950 187
rect 18062 141 18108 187
rect 23820 265 23866 311
rect 23820 101 23866 147
rect 15216 -23 15262 23
rect 15374 -23 15420 23
rect 15532 -23 15578 23
rect 15690 -23 15736 23
rect 15848 -23 15894 23
rect 16006 -23 16052 23
rect 16165 -23 16211 23
rect 16323 -23 16369 23
rect 16481 -23 16527 23
rect 16639 -23 16685 23
rect 16797 -23 16843 23
rect 16955 -23 17001 23
rect 17113 -23 17159 23
rect 17272 -23 17318 23
rect 17430 -23 17476 23
rect 17588 -23 17634 23
rect 17746 -23 17792 23
rect 17904 -23 17950 23
rect 18062 -23 18108 23
<< polysilicon >>
rect 889 14228 933 14348
rect 2933 14257 3268 14348
rect 2933 14228 3092 14257
rect 3073 14124 3092 14228
rect 889 14004 933 14124
rect 2933 14004 3092 14124
rect 3055 13900 3092 14004
rect 889 13780 933 13900
rect 2933 13835 3092 13900
rect 3138 14228 3268 14257
rect 4268 14228 4312 14348
rect 9254 14228 9324 14348
rect 9764 14228 9943 14348
rect 14048 14337 14396 14348
rect 3138 14124 3157 14228
rect 9859 14210 9943 14228
rect 12951 14282 13292 14337
rect 12951 14236 12970 14282
rect 13110 14236 13292 14282
rect 12951 14217 13292 14236
rect 13922 14228 14396 14337
rect 14920 14228 14990 14348
rect 13922 14217 14149 14228
rect 9859 14164 9878 14210
rect 9924 14164 9943 14210
rect 9859 14145 9943 14164
rect 3138 14004 3268 14124
rect 4268 14004 4312 14124
rect 20007 14228 20051 14348
rect 21051 14228 21386 14348
rect 23386 14228 23430 14348
rect 3138 13835 3157 14004
rect 4730 13917 4857 14037
rect 5957 13938 6137 14037
rect 5957 13917 6072 13938
rect 4730 13868 4789 13917
rect 2933 13780 3157 13835
rect 3217 13748 3268 13868
rect 4268 13813 4789 13868
rect 6028 13813 6072 13917
rect 4268 13748 4857 13813
rect 4730 13693 4857 13748
rect 5957 13798 6072 13813
rect 6118 13798 6137 13938
rect 5957 13693 6137 13798
rect 6275 13938 6438 14037
rect 6275 13798 6294 13938
rect 6340 13917 6438 13938
rect 7098 13917 7169 14037
rect 7423 13917 7493 14037
rect 8153 13940 8331 14037
rect 13222 14004 13292 14124
rect 13922 14087 14396 14124
rect 13922 14041 13955 14087
rect 14095 14041 14396 14087
rect 13922 14004 14396 14041
rect 14920 14004 14964 14124
rect 21153 14227 21262 14228
rect 21153 14124 21197 14227
rect 8153 13917 8266 13940
rect 6340 13813 6370 13917
rect 8224 13813 8266 13917
rect 6340 13798 6438 13813
rect 6275 13693 6438 13798
rect 7098 13693 7169 13813
rect 7423 13693 7493 13813
rect 8153 13800 8266 13813
rect 8312 13800 8331 13940
rect 18200 13965 18362 14037
rect 8153 13693 8331 13800
rect 8536 13693 8605 13813
rect 8923 13693 9195 13813
rect 9327 13779 9506 13813
rect 13222 13780 13292 13900
rect 13922 13780 14396 13900
rect 14920 13856 15220 13900
rect 14920 13810 15061 13856
rect 15201 13810 15220 13856
rect 14920 13780 15220 13810
rect 18200 13825 18219 13965
rect 18265 13917 18362 13965
rect 19462 13917 19588 14037
rect 20007 14004 20051 14124
rect 21051 14004 21197 14124
rect 18265 13825 18302 13917
rect 18200 13813 18302 13825
rect 19529 13868 19588 13917
rect 19529 13813 20051 13868
rect 9327 13733 9441 13779
rect 9487 13733 9506 13779
rect 9327 13693 9506 13733
rect 18200 13693 18362 13813
rect 19462 13748 20051 13813
rect 21051 13748 21095 13868
rect 21178 13805 21197 14004
rect 21243 14124 21262 14227
rect 21243 14004 21386 14124
rect 23386 14004 23430 14124
rect 21243 13900 21264 14004
rect 21243 13805 21386 13900
rect 21178 13780 21386 13805
rect 23386 13780 23430 13900
rect 19462 13693 19588 13748
rect 4730 13252 4857 13307
rect 889 13100 933 13220
rect 2933 13165 3157 13220
rect 2933 13100 3092 13165
rect 3055 12996 3092 13100
rect 889 12876 933 12996
rect 2933 12876 3092 12996
rect 3073 12772 3092 12876
rect 889 12652 933 12772
rect 2933 12743 3092 12772
rect 3138 12996 3157 13165
rect 3217 13132 3268 13252
rect 4268 13187 4857 13252
rect 5957 13202 6137 13307
rect 5957 13187 6072 13202
rect 4268 13132 4789 13187
rect 4730 13083 4789 13132
rect 6028 13083 6072 13187
rect 3138 12876 3268 12996
rect 4268 12876 4312 12996
rect 4730 12963 4857 13083
rect 5957 13062 6072 13083
rect 6118 13062 6137 13202
rect 5957 12963 6137 13062
rect 6275 13202 6438 13307
rect 6275 13062 6294 13202
rect 6340 13187 6438 13202
rect 7098 13187 7169 13307
rect 7423 13187 7493 13307
rect 8153 13200 8331 13307
rect 8153 13187 8266 13200
rect 6340 13083 6370 13187
rect 8224 13083 8266 13187
rect 6340 13062 6438 13083
rect 6275 12963 6438 13062
rect 7098 12963 7169 13083
rect 7423 12963 7493 13083
rect 8153 13060 8266 13083
rect 8312 13060 8331 13200
rect 8536 13187 8605 13307
rect 8923 13187 9195 13307
rect 9327 13267 9506 13307
rect 9327 13221 9441 13267
rect 9487 13221 9506 13267
rect 9327 13187 9506 13221
rect 13222 13100 13292 13220
rect 13922 13100 14396 13220
rect 14920 13190 15220 13220
rect 14920 13144 15061 13190
rect 15201 13144 15220 13190
rect 14920 13100 15220 13144
rect 18200 13187 18362 13307
rect 19462 13252 19588 13307
rect 19462 13187 20051 13252
rect 18200 13175 18302 13187
rect 8153 12963 8331 13060
rect 18200 13035 18219 13175
rect 18265 13083 18302 13175
rect 19529 13132 20051 13187
rect 21051 13132 21095 13252
rect 21178 13195 21386 13220
rect 19529 13083 19588 13132
rect 18265 13035 18362 13083
rect 3138 12772 3157 12876
rect 13222 12876 13292 12996
rect 13922 12959 14396 12996
rect 13922 12913 13955 12959
rect 14095 12913 14396 12959
rect 13922 12876 14396 12913
rect 14920 12876 14964 12996
rect 18200 12963 18362 13035
rect 19462 12963 19588 13083
rect 21178 12996 21197 13195
rect 9859 12836 9943 12855
rect 9859 12790 9878 12836
rect 9924 12790 9943 12836
rect 9859 12772 9943 12790
rect 20007 12876 20051 12996
rect 21051 12876 21197 12996
rect 3138 12743 3268 12772
rect 2933 12652 3268 12743
rect 4268 12652 4312 12772
rect 889 12428 933 12548
rect 2933 12457 3268 12548
rect 2933 12428 3092 12457
rect 3073 12324 3092 12428
rect 889 12204 933 12324
rect 2933 12204 3092 12324
rect 3055 12100 3092 12204
rect 889 11980 933 12100
rect 2933 12035 3092 12100
rect 3138 12428 3268 12457
rect 4268 12428 4312 12548
rect 9254 12652 9324 12772
rect 9764 12652 9943 12772
rect 12951 12764 13292 12783
rect 12951 12718 12970 12764
rect 13110 12718 13292 12764
rect 12951 12663 13292 12718
rect 13922 12772 14149 12783
rect 13922 12663 14396 12772
rect 9254 12428 9324 12548
rect 9764 12428 9943 12548
rect 14048 12652 14396 12663
rect 14920 12652 14990 12772
rect 21153 12773 21197 12876
rect 21243 13100 21386 13195
rect 23386 13100 23430 13220
rect 21243 12996 21264 13100
rect 21243 12876 21386 12996
rect 23386 12876 23430 12996
rect 21243 12773 21262 12876
rect 21153 12772 21262 12773
rect 20007 12652 20051 12772
rect 21051 12652 21386 12772
rect 23386 12652 23430 12772
rect 14048 12537 14396 12548
rect 3138 12324 3157 12428
rect 9859 12410 9943 12428
rect 12951 12482 13292 12537
rect 12951 12436 12970 12482
rect 13110 12436 13292 12482
rect 12951 12417 13292 12436
rect 13922 12428 14396 12537
rect 14920 12428 14990 12548
rect 13922 12417 14149 12428
rect 9859 12364 9878 12410
rect 9924 12364 9943 12410
rect 9859 12345 9943 12364
rect 3138 12204 3268 12324
rect 4268 12204 4312 12324
rect 20007 12428 20051 12548
rect 21051 12428 21386 12548
rect 23386 12428 23430 12548
rect 3138 12035 3157 12204
rect 4730 12117 4857 12237
rect 5957 12138 6137 12237
rect 5957 12117 6072 12138
rect 4730 12068 4789 12117
rect 2933 11980 3157 12035
rect 3217 11948 3268 12068
rect 4268 12013 4789 12068
rect 6028 12013 6072 12117
rect 4268 11948 4857 12013
rect 4730 11893 4857 11948
rect 5957 11998 6072 12013
rect 6118 11998 6137 12138
rect 5957 11893 6137 11998
rect 6275 12138 6438 12237
rect 6275 11998 6294 12138
rect 6340 12117 6438 12138
rect 7098 12117 7169 12237
rect 7423 12117 7493 12237
rect 8153 12140 8331 12237
rect 13222 12204 13292 12324
rect 13922 12287 14396 12324
rect 13922 12241 13955 12287
rect 14095 12241 14396 12287
rect 13922 12204 14396 12241
rect 14920 12204 14964 12324
rect 21153 12427 21262 12428
rect 21153 12324 21197 12427
rect 8153 12117 8266 12140
rect 6340 12013 6370 12117
rect 8224 12013 8266 12117
rect 6340 11998 6438 12013
rect 6275 11893 6438 11998
rect 7098 11893 7169 12013
rect 7423 11893 7493 12013
rect 8153 12000 8266 12013
rect 8312 12000 8331 12140
rect 18200 12165 18362 12237
rect 8153 11893 8331 12000
rect 8536 11893 8605 12013
rect 8923 11893 9195 12013
rect 9327 11979 9506 12013
rect 13222 11980 13292 12100
rect 13922 11980 14396 12100
rect 14920 12056 15220 12100
rect 14920 12010 15061 12056
rect 15201 12010 15220 12056
rect 14920 11980 15220 12010
rect 18200 12025 18219 12165
rect 18265 12117 18362 12165
rect 19462 12117 19588 12237
rect 20007 12204 20051 12324
rect 21051 12204 21197 12324
rect 18265 12025 18302 12117
rect 18200 12013 18302 12025
rect 19529 12068 19588 12117
rect 19529 12013 20051 12068
rect 9327 11933 9441 11979
rect 9487 11933 9506 11979
rect 9327 11893 9506 11933
rect 18200 11893 18362 12013
rect 19462 11948 20051 12013
rect 21051 11948 21095 12068
rect 21178 12005 21197 12204
rect 21243 12324 21262 12427
rect 21243 12204 21386 12324
rect 23386 12204 23430 12324
rect 21243 12100 21264 12204
rect 21243 12005 21386 12100
rect 21178 11980 21386 12005
rect 23386 11980 23430 12100
rect 19462 11893 19588 11948
rect 4730 11452 4857 11507
rect 889 11300 933 11420
rect 2933 11365 3157 11420
rect 2933 11300 3092 11365
rect 3055 11196 3092 11300
rect 889 11076 933 11196
rect 2933 11076 3092 11196
rect 3073 10972 3092 11076
rect 889 10852 933 10972
rect 2933 10943 3092 10972
rect 3138 11196 3157 11365
rect 3217 11332 3268 11452
rect 4268 11387 4857 11452
rect 5957 11402 6137 11507
rect 5957 11387 6072 11402
rect 4268 11332 4789 11387
rect 4730 11283 4789 11332
rect 6028 11283 6072 11387
rect 3138 11076 3268 11196
rect 4268 11076 4312 11196
rect 4730 11163 4857 11283
rect 5957 11262 6072 11283
rect 6118 11262 6137 11402
rect 5957 11163 6137 11262
rect 6275 11402 6438 11507
rect 6275 11262 6294 11402
rect 6340 11387 6438 11402
rect 7098 11387 7169 11507
rect 7423 11387 7493 11507
rect 8153 11400 8331 11507
rect 8153 11387 8266 11400
rect 6340 11283 6370 11387
rect 8224 11283 8266 11387
rect 6340 11262 6438 11283
rect 6275 11163 6438 11262
rect 7098 11163 7169 11283
rect 7423 11163 7493 11283
rect 8153 11260 8266 11283
rect 8312 11260 8331 11400
rect 8536 11387 8605 11507
rect 8923 11387 9195 11507
rect 9327 11467 9506 11507
rect 9327 11421 9441 11467
rect 9487 11421 9506 11467
rect 9327 11387 9506 11421
rect 13222 11300 13292 11420
rect 13922 11300 14396 11420
rect 14920 11390 15220 11420
rect 14920 11344 15061 11390
rect 15201 11344 15220 11390
rect 14920 11300 15220 11344
rect 18200 11387 18362 11507
rect 19462 11452 19588 11507
rect 19462 11387 20051 11452
rect 18200 11375 18302 11387
rect 8153 11163 8331 11260
rect 18200 11235 18219 11375
rect 18265 11283 18302 11375
rect 19529 11332 20051 11387
rect 21051 11332 21095 11452
rect 21178 11395 21386 11420
rect 19529 11283 19588 11332
rect 18265 11235 18362 11283
rect 3138 10972 3157 11076
rect 13222 11076 13292 11196
rect 13922 11159 14396 11196
rect 13922 11113 13955 11159
rect 14095 11113 14396 11159
rect 13922 11076 14396 11113
rect 14920 11076 14964 11196
rect 18200 11163 18362 11235
rect 19462 11163 19588 11283
rect 21178 11196 21197 11395
rect 9859 11036 9943 11055
rect 9859 10990 9878 11036
rect 9924 10990 9943 11036
rect 9859 10972 9943 10990
rect 20007 11076 20051 11196
rect 21051 11076 21197 11196
rect 3138 10943 3268 10972
rect 2933 10852 3268 10943
rect 4268 10852 4312 10972
rect 889 10628 933 10748
rect 2933 10657 3268 10748
rect 2933 10628 3092 10657
rect 3073 10524 3092 10628
rect 889 10404 933 10524
rect 2933 10404 3092 10524
rect 3055 10300 3092 10404
rect 889 10180 933 10300
rect 2933 10235 3092 10300
rect 3138 10628 3268 10657
rect 4268 10628 4312 10748
rect 9254 10852 9324 10972
rect 9764 10852 9943 10972
rect 12951 10964 13292 10983
rect 12951 10918 12970 10964
rect 13110 10918 13292 10964
rect 12951 10863 13292 10918
rect 13922 10972 14149 10983
rect 13922 10863 14396 10972
rect 9254 10628 9324 10748
rect 9764 10628 9943 10748
rect 14048 10852 14396 10863
rect 14920 10852 14990 10972
rect 21153 10973 21197 11076
rect 21243 11300 21386 11395
rect 23386 11300 23430 11420
rect 21243 11196 21264 11300
rect 21243 11076 21386 11196
rect 23386 11076 23430 11196
rect 21243 10973 21262 11076
rect 21153 10972 21262 10973
rect 20007 10852 20051 10972
rect 21051 10852 21386 10972
rect 23386 10852 23430 10972
rect 14048 10737 14396 10748
rect 3138 10524 3157 10628
rect 9859 10610 9943 10628
rect 12951 10682 13292 10737
rect 12951 10636 12970 10682
rect 13110 10636 13292 10682
rect 12951 10617 13292 10636
rect 13922 10628 14396 10737
rect 14920 10628 14990 10748
rect 13922 10617 14149 10628
rect 9859 10564 9878 10610
rect 9924 10564 9943 10610
rect 9859 10545 9943 10564
rect 3138 10404 3268 10524
rect 4268 10404 4312 10524
rect 20007 10628 20051 10748
rect 21051 10628 21386 10748
rect 23386 10628 23430 10748
rect 3138 10235 3157 10404
rect 4730 10317 4857 10437
rect 5957 10338 6137 10437
rect 5957 10317 6072 10338
rect 4730 10268 4789 10317
rect 2933 10180 3157 10235
rect 3217 10148 3268 10268
rect 4268 10213 4789 10268
rect 6028 10213 6072 10317
rect 4268 10148 4857 10213
rect 4730 10093 4857 10148
rect 5957 10198 6072 10213
rect 6118 10198 6137 10338
rect 5957 10093 6137 10198
rect 6275 10338 6438 10437
rect 6275 10198 6294 10338
rect 6340 10317 6438 10338
rect 7098 10317 7169 10437
rect 7423 10317 7493 10437
rect 8153 10340 8331 10437
rect 13222 10404 13292 10524
rect 13922 10487 14396 10524
rect 13922 10441 13955 10487
rect 14095 10441 14396 10487
rect 13922 10404 14396 10441
rect 14920 10404 14964 10524
rect 21153 10627 21262 10628
rect 21153 10524 21197 10627
rect 8153 10317 8266 10340
rect 6340 10213 6370 10317
rect 8224 10213 8266 10317
rect 6340 10198 6438 10213
rect 6275 10093 6438 10198
rect 7098 10093 7169 10213
rect 7423 10093 7493 10213
rect 8153 10200 8266 10213
rect 8312 10200 8331 10340
rect 18200 10365 18362 10437
rect 8153 10093 8331 10200
rect 8536 10093 8605 10213
rect 8923 10093 9195 10213
rect 9327 10179 9506 10213
rect 13222 10180 13292 10300
rect 13922 10180 14396 10300
rect 14920 10256 15220 10300
rect 14920 10210 15061 10256
rect 15201 10210 15220 10256
rect 14920 10180 15220 10210
rect 18200 10225 18219 10365
rect 18265 10317 18362 10365
rect 19462 10317 19588 10437
rect 20007 10404 20051 10524
rect 21051 10404 21197 10524
rect 18265 10225 18302 10317
rect 18200 10213 18302 10225
rect 19529 10268 19588 10317
rect 19529 10213 20051 10268
rect 9327 10133 9441 10179
rect 9487 10133 9506 10179
rect 9327 10093 9506 10133
rect 18200 10093 18362 10213
rect 19462 10148 20051 10213
rect 21051 10148 21095 10268
rect 21178 10205 21197 10404
rect 21243 10524 21262 10627
rect 21243 10404 21386 10524
rect 23386 10404 23430 10524
rect 21243 10300 21264 10404
rect 21243 10205 21386 10300
rect 21178 10180 21386 10205
rect 23386 10180 23430 10300
rect 19462 10093 19588 10148
rect 4730 9652 4857 9707
rect 889 9500 933 9620
rect 2933 9565 3157 9620
rect 2933 9500 3092 9565
rect 3055 9396 3092 9500
rect 889 9276 933 9396
rect 2933 9276 3092 9396
rect 3073 9172 3092 9276
rect 889 9052 933 9172
rect 2933 9143 3092 9172
rect 3138 9396 3157 9565
rect 3217 9532 3268 9652
rect 4268 9587 4857 9652
rect 5957 9602 6137 9707
rect 5957 9587 6072 9602
rect 4268 9532 4789 9587
rect 4730 9483 4789 9532
rect 6028 9483 6072 9587
rect 3138 9276 3268 9396
rect 4268 9276 4312 9396
rect 4730 9363 4857 9483
rect 5957 9462 6072 9483
rect 6118 9462 6137 9602
rect 5957 9363 6137 9462
rect 6275 9602 6438 9707
rect 6275 9462 6294 9602
rect 6340 9587 6438 9602
rect 7098 9587 7169 9707
rect 7423 9587 7493 9707
rect 8153 9600 8331 9707
rect 8153 9587 8266 9600
rect 6340 9483 6370 9587
rect 8224 9483 8266 9587
rect 6340 9462 6438 9483
rect 6275 9363 6438 9462
rect 7098 9363 7169 9483
rect 7423 9363 7493 9483
rect 8153 9460 8266 9483
rect 8312 9460 8331 9600
rect 8536 9587 8605 9707
rect 8923 9587 9195 9707
rect 9327 9667 9506 9707
rect 9327 9621 9441 9667
rect 9487 9621 9506 9667
rect 9327 9587 9506 9621
rect 13222 9500 13292 9620
rect 13922 9500 14396 9620
rect 14920 9590 15220 9620
rect 14920 9544 15061 9590
rect 15201 9544 15220 9590
rect 14920 9500 15220 9544
rect 18200 9587 18362 9707
rect 19462 9652 19588 9707
rect 19462 9587 20051 9652
rect 18200 9575 18302 9587
rect 8153 9363 8331 9460
rect 18200 9435 18219 9575
rect 18265 9483 18302 9575
rect 19529 9532 20051 9587
rect 21051 9532 21095 9652
rect 21178 9595 21386 9620
rect 19529 9483 19588 9532
rect 18265 9435 18362 9483
rect 3138 9172 3157 9276
rect 13222 9276 13292 9396
rect 13922 9359 14396 9396
rect 13922 9313 13955 9359
rect 14095 9313 14396 9359
rect 13922 9276 14396 9313
rect 14920 9276 14964 9396
rect 18200 9363 18362 9435
rect 19462 9363 19588 9483
rect 21178 9396 21197 9595
rect 9859 9236 9943 9255
rect 9859 9190 9878 9236
rect 9924 9190 9943 9236
rect 9859 9172 9943 9190
rect 20007 9276 20051 9396
rect 21051 9276 21197 9396
rect 3138 9143 3268 9172
rect 2933 9052 3268 9143
rect 4268 9052 4312 9172
rect 889 8828 933 8948
rect 2933 8857 3268 8948
rect 2933 8828 3092 8857
rect 3073 8724 3092 8828
rect 889 8604 933 8724
rect 2933 8604 3092 8724
rect 3055 8500 3092 8604
rect 889 8380 933 8500
rect 2933 8435 3092 8500
rect 3138 8828 3268 8857
rect 4268 8828 4312 8948
rect 9254 9052 9324 9172
rect 9764 9052 9943 9172
rect 12951 9164 13292 9183
rect 12951 9118 12970 9164
rect 13110 9118 13292 9164
rect 12951 9063 13292 9118
rect 13922 9172 14149 9183
rect 13922 9063 14396 9172
rect 9254 8828 9324 8948
rect 9764 8828 9943 8948
rect 14048 9052 14396 9063
rect 14920 9052 14990 9172
rect 21153 9173 21197 9276
rect 21243 9500 21386 9595
rect 23386 9500 23430 9620
rect 21243 9396 21264 9500
rect 21243 9276 21386 9396
rect 23386 9276 23430 9396
rect 21243 9173 21262 9276
rect 21153 9172 21262 9173
rect 20007 9052 20051 9172
rect 21051 9052 21386 9172
rect 23386 9052 23430 9172
rect 14048 8937 14396 8948
rect 3138 8724 3157 8828
rect 9859 8810 9943 8828
rect 12951 8882 13292 8937
rect 12951 8836 12970 8882
rect 13110 8836 13292 8882
rect 12951 8817 13292 8836
rect 13922 8828 14396 8937
rect 14920 8828 14990 8948
rect 13922 8817 14149 8828
rect 9859 8764 9878 8810
rect 9924 8764 9943 8810
rect 9859 8745 9943 8764
rect 3138 8604 3268 8724
rect 4268 8604 4312 8724
rect 20007 8828 20051 8948
rect 21051 8828 21386 8948
rect 23386 8828 23430 8948
rect 3138 8435 3157 8604
rect 4730 8517 4857 8637
rect 5957 8538 6137 8637
rect 5957 8517 6072 8538
rect 4730 8468 4789 8517
rect 2933 8380 3157 8435
rect 3217 8348 3268 8468
rect 4268 8413 4789 8468
rect 6028 8413 6072 8517
rect 4268 8348 4857 8413
rect 4730 8293 4857 8348
rect 5957 8398 6072 8413
rect 6118 8398 6137 8538
rect 5957 8293 6137 8398
rect 6275 8538 6438 8637
rect 6275 8398 6294 8538
rect 6340 8517 6438 8538
rect 7098 8517 7169 8637
rect 7423 8517 7493 8637
rect 8153 8540 8331 8637
rect 13222 8604 13292 8724
rect 13922 8687 14396 8724
rect 13922 8641 13955 8687
rect 14095 8641 14396 8687
rect 13922 8604 14396 8641
rect 14920 8604 14964 8724
rect 21153 8827 21262 8828
rect 21153 8724 21197 8827
rect 8153 8517 8266 8540
rect 6340 8413 6370 8517
rect 8224 8413 8266 8517
rect 6340 8398 6438 8413
rect 6275 8293 6438 8398
rect 7098 8293 7169 8413
rect 7423 8293 7493 8413
rect 8153 8400 8266 8413
rect 8312 8400 8331 8540
rect 18200 8565 18362 8637
rect 8153 8293 8331 8400
rect 8536 8293 8605 8413
rect 8923 8293 9195 8413
rect 9327 8379 9506 8413
rect 13222 8380 13292 8500
rect 13922 8380 14396 8500
rect 14920 8456 15220 8500
rect 14920 8410 15061 8456
rect 15201 8410 15220 8456
rect 14920 8380 15220 8410
rect 18200 8425 18219 8565
rect 18265 8517 18362 8565
rect 19462 8517 19588 8637
rect 20007 8604 20051 8724
rect 21051 8604 21197 8724
rect 18265 8425 18302 8517
rect 18200 8413 18302 8425
rect 19529 8468 19588 8517
rect 19529 8413 20051 8468
rect 9327 8333 9441 8379
rect 9487 8333 9506 8379
rect 9327 8293 9506 8333
rect 18200 8293 18362 8413
rect 19462 8348 20051 8413
rect 21051 8348 21095 8468
rect 21178 8405 21197 8604
rect 21243 8724 21262 8827
rect 21243 8604 21386 8724
rect 23386 8604 23430 8724
rect 21243 8500 21264 8604
rect 21243 8405 21386 8500
rect 21178 8380 21386 8405
rect 23386 8380 23430 8500
rect 19462 8293 19588 8348
rect 4730 7852 4857 7907
rect 889 7700 933 7820
rect 2933 7765 3157 7820
rect 2933 7700 3092 7765
rect 3055 7596 3092 7700
rect 889 7476 933 7596
rect 2933 7476 3092 7596
rect 3073 7372 3092 7476
rect 889 7252 933 7372
rect 2933 7343 3092 7372
rect 3138 7596 3157 7765
rect 3217 7732 3268 7852
rect 4268 7787 4857 7852
rect 5957 7802 6137 7907
rect 5957 7787 6072 7802
rect 4268 7732 4789 7787
rect 4730 7683 4789 7732
rect 6028 7683 6072 7787
rect 3138 7476 3268 7596
rect 4268 7476 4312 7596
rect 4730 7563 4857 7683
rect 5957 7662 6072 7683
rect 6118 7662 6137 7802
rect 5957 7563 6137 7662
rect 6275 7802 6438 7907
rect 6275 7662 6294 7802
rect 6340 7787 6438 7802
rect 7098 7787 7169 7907
rect 7423 7787 7493 7907
rect 8153 7800 8331 7907
rect 8153 7787 8266 7800
rect 6340 7683 6370 7787
rect 8224 7683 8266 7787
rect 6340 7662 6438 7683
rect 6275 7563 6438 7662
rect 7098 7563 7169 7683
rect 7423 7563 7493 7683
rect 8153 7660 8266 7683
rect 8312 7660 8331 7800
rect 8536 7787 8605 7907
rect 8923 7787 9195 7907
rect 9327 7867 9506 7907
rect 9327 7821 9441 7867
rect 9487 7821 9506 7867
rect 9327 7787 9506 7821
rect 13222 7700 13292 7820
rect 13922 7700 14396 7820
rect 14920 7790 15220 7820
rect 14920 7744 15061 7790
rect 15201 7744 15220 7790
rect 14920 7700 15220 7744
rect 18200 7787 18362 7907
rect 19462 7852 19588 7907
rect 19462 7787 20051 7852
rect 18200 7775 18302 7787
rect 8153 7563 8331 7660
rect 18200 7635 18219 7775
rect 18265 7683 18302 7775
rect 19529 7732 20051 7787
rect 21051 7732 21095 7852
rect 21178 7795 21386 7820
rect 19529 7683 19588 7732
rect 18265 7635 18362 7683
rect 3138 7372 3157 7476
rect 13222 7476 13292 7596
rect 13922 7559 14396 7596
rect 13922 7513 13955 7559
rect 14095 7513 14396 7559
rect 13922 7476 14396 7513
rect 14920 7476 14964 7596
rect 18200 7563 18362 7635
rect 19462 7563 19588 7683
rect 21178 7596 21197 7795
rect 9859 7436 9943 7455
rect 9859 7390 9878 7436
rect 9924 7390 9943 7436
rect 9859 7372 9943 7390
rect 20007 7476 20051 7596
rect 21051 7476 21197 7596
rect 3138 7343 3268 7372
rect 2933 7252 3268 7343
rect 4268 7252 4312 7372
rect 889 7028 933 7148
rect 2933 7057 3268 7148
rect 2933 7028 3092 7057
rect 3073 6924 3092 7028
rect 889 6804 933 6924
rect 2933 6804 3092 6924
rect 3055 6700 3092 6804
rect 889 6580 933 6700
rect 2933 6635 3092 6700
rect 3138 7028 3268 7057
rect 4268 7028 4312 7148
rect 9254 7252 9324 7372
rect 9764 7252 9943 7372
rect 12951 7364 13292 7383
rect 12951 7318 12970 7364
rect 13110 7318 13292 7364
rect 12951 7263 13292 7318
rect 13922 7372 14149 7383
rect 13922 7263 14396 7372
rect 9254 7028 9324 7148
rect 9764 7028 9943 7148
rect 14048 7252 14396 7263
rect 14920 7252 14990 7372
rect 21153 7373 21197 7476
rect 21243 7700 21386 7795
rect 23386 7700 23430 7820
rect 21243 7596 21264 7700
rect 21243 7476 21386 7596
rect 23386 7476 23430 7596
rect 21243 7373 21262 7476
rect 21153 7372 21262 7373
rect 20007 7252 20051 7372
rect 21051 7252 21386 7372
rect 23386 7252 23430 7372
rect 14048 7137 14396 7148
rect 3138 6924 3157 7028
rect 9859 7010 9943 7028
rect 12951 7082 13292 7137
rect 12951 7036 12970 7082
rect 13110 7036 13292 7082
rect 12951 7017 13292 7036
rect 13922 7028 14396 7137
rect 14920 7028 14990 7148
rect 13922 7017 14149 7028
rect 9859 6964 9878 7010
rect 9924 6964 9943 7010
rect 9859 6945 9943 6964
rect 3138 6804 3268 6924
rect 4268 6804 4312 6924
rect 20007 7028 20051 7148
rect 21051 7028 21386 7148
rect 23386 7028 23430 7148
rect 3138 6635 3157 6804
rect 4730 6717 4857 6837
rect 5957 6738 6137 6837
rect 5957 6717 6072 6738
rect 4730 6668 4789 6717
rect 2933 6580 3157 6635
rect 3217 6548 3268 6668
rect 4268 6613 4789 6668
rect 6028 6613 6072 6717
rect 4268 6548 4857 6613
rect 4730 6493 4857 6548
rect 5957 6598 6072 6613
rect 6118 6598 6137 6738
rect 5957 6493 6137 6598
rect 6275 6738 6438 6837
rect 6275 6598 6294 6738
rect 6340 6717 6438 6738
rect 7098 6717 7169 6837
rect 7423 6717 7493 6837
rect 8153 6740 8331 6837
rect 13222 6804 13292 6924
rect 13922 6887 14396 6924
rect 13922 6841 13955 6887
rect 14095 6841 14396 6887
rect 13922 6804 14396 6841
rect 14920 6804 14964 6924
rect 21153 7027 21262 7028
rect 21153 6924 21197 7027
rect 8153 6717 8266 6740
rect 6340 6613 6370 6717
rect 8224 6613 8266 6717
rect 6340 6598 6438 6613
rect 6275 6493 6438 6598
rect 7098 6493 7169 6613
rect 7423 6493 7493 6613
rect 8153 6600 8266 6613
rect 8312 6600 8331 6740
rect 18200 6765 18362 6837
rect 8153 6493 8331 6600
rect 8536 6493 8605 6613
rect 8923 6493 9195 6613
rect 9327 6579 9506 6613
rect 13222 6580 13292 6700
rect 13922 6580 14396 6700
rect 14920 6656 15220 6700
rect 14920 6610 15061 6656
rect 15201 6610 15220 6656
rect 14920 6580 15220 6610
rect 18200 6625 18219 6765
rect 18265 6717 18362 6765
rect 19462 6717 19588 6837
rect 20007 6804 20051 6924
rect 21051 6804 21197 6924
rect 18265 6625 18302 6717
rect 18200 6613 18302 6625
rect 19529 6668 19588 6717
rect 19529 6613 20051 6668
rect 9327 6533 9441 6579
rect 9487 6533 9506 6579
rect 9327 6493 9506 6533
rect 18200 6493 18362 6613
rect 19462 6548 20051 6613
rect 21051 6548 21095 6668
rect 21178 6605 21197 6804
rect 21243 6924 21262 7027
rect 21243 6804 21386 6924
rect 23386 6804 23430 6924
rect 21243 6700 21264 6804
rect 21243 6605 21386 6700
rect 21178 6580 21386 6605
rect 23386 6580 23430 6700
rect 19462 6493 19588 6548
rect 4730 6052 4857 6107
rect 889 5900 933 6020
rect 2933 5965 3157 6020
rect 2933 5900 3092 5965
rect 3055 5796 3092 5900
rect 889 5676 933 5796
rect 2933 5676 3092 5796
rect 3073 5572 3092 5676
rect 889 5452 933 5572
rect 2933 5543 3092 5572
rect 3138 5796 3157 5965
rect 3217 5932 3268 6052
rect 4268 5987 4857 6052
rect 5957 6002 6137 6107
rect 5957 5987 6072 6002
rect 4268 5932 4789 5987
rect 4730 5883 4789 5932
rect 6028 5883 6072 5987
rect 3138 5676 3268 5796
rect 4268 5676 4312 5796
rect 4730 5763 4857 5883
rect 5957 5862 6072 5883
rect 6118 5862 6137 6002
rect 5957 5763 6137 5862
rect 6275 6002 6438 6107
rect 6275 5862 6294 6002
rect 6340 5987 6438 6002
rect 7098 5987 7169 6107
rect 7423 5987 7493 6107
rect 8153 6000 8331 6107
rect 8153 5987 8266 6000
rect 6340 5883 6370 5987
rect 8224 5883 8266 5987
rect 6340 5862 6438 5883
rect 6275 5763 6438 5862
rect 7098 5763 7169 5883
rect 7423 5763 7493 5883
rect 8153 5860 8266 5883
rect 8312 5860 8331 6000
rect 8536 5987 8605 6107
rect 8923 5987 9195 6107
rect 9327 6067 9506 6107
rect 9327 6021 9441 6067
rect 9487 6021 9506 6067
rect 9327 5987 9506 6021
rect 13222 5900 13292 6020
rect 13922 5900 14396 6020
rect 14920 5990 15220 6020
rect 14920 5944 15061 5990
rect 15201 5944 15220 5990
rect 14920 5900 15220 5944
rect 18200 5987 18362 6107
rect 19462 6052 19588 6107
rect 19462 5987 20051 6052
rect 18200 5975 18302 5987
rect 8153 5763 8331 5860
rect 18200 5835 18219 5975
rect 18265 5883 18302 5975
rect 19529 5932 20051 5987
rect 21051 5932 21095 6052
rect 21178 5995 21386 6020
rect 19529 5883 19588 5932
rect 18265 5835 18362 5883
rect 3138 5572 3157 5676
rect 13222 5676 13292 5796
rect 13922 5759 14396 5796
rect 13922 5713 13955 5759
rect 14095 5713 14396 5759
rect 13922 5676 14396 5713
rect 14920 5676 14964 5796
rect 18200 5763 18362 5835
rect 19462 5763 19588 5883
rect 21178 5796 21197 5995
rect 9859 5636 9943 5655
rect 9859 5590 9878 5636
rect 9924 5590 9943 5636
rect 9859 5572 9943 5590
rect 20007 5676 20051 5796
rect 21051 5676 21197 5796
rect 3138 5543 3268 5572
rect 2933 5452 3268 5543
rect 4268 5452 4312 5572
rect 889 5228 933 5348
rect 2933 5257 3268 5348
rect 2933 5228 3092 5257
rect 3073 5124 3092 5228
rect 889 5004 933 5124
rect 2933 5004 3092 5124
rect 3055 4900 3092 5004
rect 889 4780 933 4900
rect 2933 4835 3092 4900
rect 3138 5228 3268 5257
rect 4268 5228 4312 5348
rect 9254 5452 9324 5572
rect 9764 5452 9943 5572
rect 12951 5564 13292 5583
rect 12951 5518 12970 5564
rect 13110 5518 13292 5564
rect 12951 5463 13292 5518
rect 13922 5572 14149 5583
rect 13922 5463 14396 5572
rect 9254 5228 9324 5348
rect 9764 5228 9943 5348
rect 14048 5452 14396 5463
rect 14920 5452 14990 5572
rect 21153 5573 21197 5676
rect 21243 5900 21386 5995
rect 23386 5900 23430 6020
rect 21243 5796 21264 5900
rect 21243 5676 21386 5796
rect 23386 5676 23430 5796
rect 21243 5573 21262 5676
rect 21153 5572 21262 5573
rect 20007 5452 20051 5572
rect 21051 5452 21386 5572
rect 23386 5452 23430 5572
rect 14048 5337 14396 5348
rect 3138 5124 3157 5228
rect 9859 5210 9943 5228
rect 12951 5282 13292 5337
rect 12951 5236 12970 5282
rect 13110 5236 13292 5282
rect 12951 5217 13292 5236
rect 13922 5228 14396 5337
rect 14920 5228 14990 5348
rect 13922 5217 14149 5228
rect 9859 5164 9878 5210
rect 9924 5164 9943 5210
rect 9859 5145 9943 5164
rect 3138 5004 3268 5124
rect 4268 5004 4312 5124
rect 20007 5228 20051 5348
rect 21051 5228 21386 5348
rect 23386 5228 23430 5348
rect 3138 4835 3157 5004
rect 4730 4917 4857 5037
rect 5957 4938 6137 5037
rect 5957 4917 6072 4938
rect 4730 4868 4789 4917
rect 2933 4780 3157 4835
rect 3217 4748 3268 4868
rect 4268 4813 4789 4868
rect 6028 4813 6072 4917
rect 4268 4748 4857 4813
rect 4730 4693 4857 4748
rect 5957 4798 6072 4813
rect 6118 4798 6137 4938
rect 5957 4693 6137 4798
rect 6275 4938 6438 5037
rect 6275 4798 6294 4938
rect 6340 4917 6438 4938
rect 7098 4917 7169 5037
rect 7423 4917 7493 5037
rect 8153 4940 8331 5037
rect 13222 5004 13292 5124
rect 13922 5087 14396 5124
rect 13922 5041 13955 5087
rect 14095 5041 14396 5087
rect 13922 5004 14396 5041
rect 14920 5004 14964 5124
rect 21153 5227 21262 5228
rect 21153 5124 21197 5227
rect 8153 4917 8266 4940
rect 6340 4813 6370 4917
rect 8224 4813 8266 4917
rect 6340 4798 6438 4813
rect 6275 4693 6438 4798
rect 7098 4693 7169 4813
rect 7423 4693 7493 4813
rect 8153 4800 8266 4813
rect 8312 4800 8331 4940
rect 18200 4965 18362 5037
rect 8153 4693 8331 4800
rect 8536 4693 8605 4813
rect 8923 4693 9195 4813
rect 9327 4779 9506 4813
rect 13222 4780 13292 4900
rect 13922 4780 14396 4900
rect 14920 4856 15220 4900
rect 14920 4810 15061 4856
rect 15201 4810 15220 4856
rect 14920 4780 15220 4810
rect 18200 4825 18219 4965
rect 18265 4917 18362 4965
rect 19462 4917 19588 5037
rect 20007 5004 20051 5124
rect 21051 5004 21197 5124
rect 18265 4825 18302 4917
rect 18200 4813 18302 4825
rect 19529 4868 19588 4917
rect 19529 4813 20051 4868
rect 9327 4733 9441 4779
rect 9487 4733 9506 4779
rect 9327 4693 9506 4733
rect 18200 4693 18362 4813
rect 19462 4748 20051 4813
rect 21051 4748 21095 4868
rect 21178 4805 21197 5004
rect 21243 5124 21262 5227
rect 21243 5004 21386 5124
rect 23386 5004 23430 5124
rect 21243 4900 21264 5004
rect 21243 4805 21386 4900
rect 21178 4780 21386 4805
rect 23386 4780 23430 4900
rect 19462 4693 19588 4748
rect 4730 4252 4857 4307
rect 889 4100 933 4220
rect 2933 4165 3157 4220
rect 2933 4100 3092 4165
rect 3055 3996 3092 4100
rect 889 3876 933 3996
rect 2933 3876 3092 3996
rect 3073 3772 3092 3876
rect 889 3652 933 3772
rect 2933 3743 3092 3772
rect 3138 3996 3157 4165
rect 3217 4132 3268 4252
rect 4268 4187 4857 4252
rect 5957 4202 6137 4307
rect 5957 4187 6072 4202
rect 4268 4132 4789 4187
rect 4730 4083 4789 4132
rect 6028 4083 6072 4187
rect 3138 3876 3268 3996
rect 4268 3876 4312 3996
rect 4730 3963 4857 4083
rect 5957 4062 6072 4083
rect 6118 4062 6137 4202
rect 5957 3963 6137 4062
rect 6275 4202 6438 4307
rect 6275 4062 6294 4202
rect 6340 4187 6438 4202
rect 7098 4187 7169 4307
rect 7423 4187 7493 4307
rect 8153 4200 8331 4307
rect 8153 4187 8266 4200
rect 6340 4083 6370 4187
rect 8224 4083 8266 4187
rect 6340 4062 6438 4083
rect 6275 3963 6438 4062
rect 7098 3963 7169 4083
rect 7423 3963 7493 4083
rect 8153 4060 8266 4083
rect 8312 4060 8331 4200
rect 8536 4187 8605 4307
rect 8923 4187 9195 4307
rect 9327 4267 9506 4307
rect 9327 4221 9441 4267
rect 9487 4221 9506 4267
rect 9327 4187 9506 4221
rect 13222 4100 13292 4220
rect 13922 4100 14396 4220
rect 14920 4190 15220 4220
rect 14920 4144 15061 4190
rect 15201 4144 15220 4190
rect 14920 4100 15220 4144
rect 18200 4187 18362 4307
rect 19462 4252 19588 4307
rect 19462 4187 20051 4252
rect 18200 4175 18302 4187
rect 8153 3963 8331 4060
rect 18200 4035 18219 4175
rect 18265 4083 18302 4175
rect 19529 4132 20051 4187
rect 21051 4132 21095 4252
rect 21178 4195 21386 4220
rect 19529 4083 19588 4132
rect 18265 4035 18362 4083
rect 3138 3772 3157 3876
rect 13222 3876 13292 3996
rect 13922 3959 14396 3996
rect 13922 3913 13955 3959
rect 14095 3913 14396 3959
rect 13922 3876 14396 3913
rect 14920 3876 14964 3996
rect 18200 3963 18362 4035
rect 19462 3963 19588 4083
rect 21178 3996 21197 4195
rect 9859 3836 9943 3855
rect 9859 3790 9878 3836
rect 9924 3790 9943 3836
rect 9859 3772 9943 3790
rect 20007 3876 20051 3996
rect 21051 3876 21197 3996
rect 3138 3743 3268 3772
rect 2933 3652 3268 3743
rect 4268 3652 4312 3772
rect 889 3428 933 3548
rect 2933 3457 3268 3548
rect 2933 3428 3092 3457
rect 3073 3324 3092 3428
rect 889 3204 933 3324
rect 2933 3204 3092 3324
rect 3055 3100 3092 3204
rect 889 2980 933 3100
rect 2933 3035 3092 3100
rect 3138 3428 3268 3457
rect 4268 3428 4312 3548
rect 9254 3652 9324 3772
rect 9764 3652 9943 3772
rect 12951 3764 13292 3783
rect 12951 3718 12970 3764
rect 13110 3718 13292 3764
rect 12951 3663 13292 3718
rect 13922 3772 14149 3783
rect 13922 3663 14396 3772
rect 9254 3428 9324 3548
rect 9764 3428 9943 3548
rect 14048 3652 14396 3663
rect 14920 3652 14990 3772
rect 21153 3773 21197 3876
rect 21243 4100 21386 4195
rect 23386 4100 23430 4220
rect 21243 3996 21264 4100
rect 21243 3876 21386 3996
rect 23386 3876 23430 3996
rect 21243 3773 21262 3876
rect 21153 3772 21262 3773
rect 20007 3652 20051 3772
rect 21051 3652 21386 3772
rect 23386 3652 23430 3772
rect 14048 3537 14396 3548
rect 3138 3324 3157 3428
rect 9859 3410 9943 3428
rect 12951 3482 13292 3537
rect 12951 3436 12970 3482
rect 13110 3436 13292 3482
rect 12951 3417 13292 3436
rect 13922 3428 14396 3537
rect 14920 3428 14990 3548
rect 13922 3417 14149 3428
rect 9859 3364 9878 3410
rect 9924 3364 9943 3410
rect 9859 3345 9943 3364
rect 3138 3204 3268 3324
rect 4268 3204 4312 3324
rect 20007 3428 20051 3548
rect 21051 3428 21386 3548
rect 23386 3428 23430 3548
rect 3138 3035 3157 3204
rect 4730 3117 4857 3237
rect 5957 3138 6137 3237
rect 5957 3117 6072 3138
rect 4730 3068 4789 3117
rect 2933 2980 3157 3035
rect 3217 2948 3268 3068
rect 4268 3013 4789 3068
rect 6028 3013 6072 3117
rect 4268 2948 4857 3013
rect 4730 2893 4857 2948
rect 5957 2998 6072 3013
rect 6118 2998 6137 3138
rect 5957 2893 6137 2998
rect 6275 3138 6438 3237
rect 6275 2998 6294 3138
rect 6340 3117 6438 3138
rect 7098 3117 7169 3237
rect 7423 3117 7493 3237
rect 8153 3140 8331 3237
rect 13222 3204 13292 3324
rect 13922 3287 14396 3324
rect 13922 3241 13955 3287
rect 14095 3241 14396 3287
rect 13922 3204 14396 3241
rect 14920 3204 14964 3324
rect 21153 3427 21262 3428
rect 21153 3324 21197 3427
rect 8153 3117 8266 3140
rect 6340 3013 6370 3117
rect 8224 3013 8266 3117
rect 6340 2998 6438 3013
rect 6275 2893 6438 2998
rect 7098 2893 7169 3013
rect 7423 2893 7493 3013
rect 8153 3000 8266 3013
rect 8312 3000 8331 3140
rect 18200 3165 18362 3237
rect 8153 2893 8331 3000
rect 8536 2893 8605 3013
rect 8923 2893 9195 3013
rect 9327 2979 9506 3013
rect 13222 2980 13292 3100
rect 13922 2980 14396 3100
rect 14920 3056 15220 3100
rect 14920 3010 15061 3056
rect 15201 3010 15220 3056
rect 14920 2980 15220 3010
rect 18200 3025 18219 3165
rect 18265 3117 18362 3165
rect 19462 3117 19588 3237
rect 20007 3204 20051 3324
rect 21051 3204 21197 3324
rect 18265 3025 18302 3117
rect 18200 3013 18302 3025
rect 19529 3068 19588 3117
rect 19529 3013 20051 3068
rect 9327 2933 9441 2979
rect 9487 2933 9506 2979
rect 9327 2893 9506 2933
rect 18200 2893 18362 3013
rect 19462 2948 20051 3013
rect 21051 2948 21095 3068
rect 21178 3005 21197 3204
rect 21243 3324 21262 3427
rect 21243 3204 21386 3324
rect 23386 3204 23430 3324
rect 21243 3100 21264 3204
rect 21243 3005 21386 3100
rect 21178 2980 21386 3005
rect 23386 2980 23430 3100
rect 19462 2893 19588 2948
rect 4730 2452 4857 2507
rect 889 2300 933 2420
rect 2933 2365 3157 2420
rect 2933 2300 3092 2365
rect 3055 2196 3092 2300
rect 889 2076 933 2196
rect 2933 2076 3092 2196
rect 3073 1972 3092 2076
rect 889 1852 933 1972
rect 2933 1943 3092 1972
rect 3138 2196 3157 2365
rect 3217 2332 3268 2452
rect 4268 2387 4857 2452
rect 5957 2402 6137 2507
rect 5957 2387 6072 2402
rect 4268 2332 4789 2387
rect 4730 2283 4789 2332
rect 6028 2283 6072 2387
rect 3138 2076 3268 2196
rect 4268 2076 4312 2196
rect 4730 2163 4857 2283
rect 5957 2262 6072 2283
rect 6118 2262 6137 2402
rect 5957 2163 6137 2262
rect 6275 2402 6438 2507
rect 6275 2262 6294 2402
rect 6340 2387 6438 2402
rect 7098 2387 7169 2507
rect 7423 2387 7493 2507
rect 8153 2400 8331 2507
rect 8153 2387 8266 2400
rect 6340 2283 6370 2387
rect 8224 2283 8266 2387
rect 6340 2262 6438 2283
rect 6275 2163 6438 2262
rect 7098 2163 7169 2283
rect 7423 2163 7493 2283
rect 8153 2260 8266 2283
rect 8312 2260 8331 2400
rect 8536 2387 8605 2507
rect 8923 2387 9195 2507
rect 9327 2467 9506 2507
rect 9327 2421 9441 2467
rect 9487 2421 9506 2467
rect 9327 2387 9506 2421
rect 13222 2300 13292 2420
rect 13922 2300 14396 2420
rect 14920 2390 15220 2420
rect 14920 2344 15061 2390
rect 15201 2344 15220 2390
rect 14920 2300 15220 2344
rect 18200 2387 18362 2507
rect 19462 2452 19588 2507
rect 19462 2387 20051 2452
rect 18200 2375 18302 2387
rect 8153 2163 8331 2260
rect 18200 2235 18219 2375
rect 18265 2283 18302 2375
rect 19529 2332 20051 2387
rect 21051 2332 21095 2452
rect 21178 2395 21386 2420
rect 19529 2283 19588 2332
rect 18265 2235 18362 2283
rect 3138 1972 3157 2076
rect 13222 2076 13292 2196
rect 13922 2159 14396 2196
rect 13922 2113 13955 2159
rect 14095 2113 14396 2159
rect 13922 2076 14396 2113
rect 14920 2076 14964 2196
rect 18200 2163 18362 2235
rect 19462 2163 19588 2283
rect 21178 2196 21197 2395
rect 9859 2036 9943 2055
rect 9859 1990 9878 2036
rect 9924 1990 9943 2036
rect 9859 1972 9943 1990
rect 20007 2076 20051 2196
rect 21051 2076 21197 2196
rect 3138 1943 3268 1972
rect 2933 1852 3268 1943
rect 4268 1852 4312 1972
rect 889 1628 933 1748
rect 2933 1657 3268 1748
rect 2933 1628 3092 1657
rect 3073 1524 3092 1628
rect 889 1404 933 1524
rect 2933 1404 3092 1524
rect 3055 1300 3092 1404
rect 889 1180 933 1300
rect 2933 1235 3092 1300
rect 3138 1628 3268 1657
rect 4268 1628 4312 1748
rect 9254 1852 9324 1972
rect 9764 1852 9943 1972
rect 12951 1964 13292 1983
rect 12951 1918 12970 1964
rect 13110 1918 13292 1964
rect 12951 1863 13292 1918
rect 13922 1972 14149 1983
rect 13922 1863 14396 1972
rect 9254 1628 9324 1748
rect 9764 1628 9943 1748
rect 14048 1852 14396 1863
rect 14920 1852 14990 1972
rect 21153 1973 21197 2076
rect 21243 2300 21386 2395
rect 23386 2300 23430 2420
rect 21243 2196 21264 2300
rect 21243 2076 21386 2196
rect 23386 2076 23430 2196
rect 21243 1973 21262 2076
rect 21153 1972 21262 1973
rect 20007 1852 20051 1972
rect 21051 1852 21386 1972
rect 23386 1852 23430 1972
rect 14048 1737 14396 1748
rect 3138 1524 3157 1628
rect 9859 1610 9943 1628
rect 12951 1682 13292 1737
rect 12951 1636 12970 1682
rect 13110 1636 13292 1682
rect 12951 1617 13292 1636
rect 13922 1628 14396 1737
rect 14920 1628 14990 1748
rect 13922 1617 14149 1628
rect 9859 1564 9878 1610
rect 9924 1564 9943 1610
rect 9859 1545 9943 1564
rect 3138 1404 3268 1524
rect 4268 1404 4312 1524
rect 20007 1628 20051 1748
rect 21051 1628 21386 1748
rect 23386 1628 23430 1748
rect 3138 1235 3157 1404
rect 4730 1317 4857 1437
rect 5957 1338 6137 1437
rect 5957 1317 6072 1338
rect 4730 1268 4789 1317
rect 2933 1180 3157 1235
rect 3217 1148 3268 1268
rect 4268 1213 4789 1268
rect 6028 1213 6072 1317
rect 4268 1148 4857 1213
rect 4730 1093 4857 1148
rect 5957 1198 6072 1213
rect 6118 1198 6137 1338
rect 5957 1093 6137 1198
rect 6275 1338 6438 1437
rect 6275 1198 6294 1338
rect 6340 1317 6438 1338
rect 7098 1317 7169 1437
rect 7423 1317 7493 1437
rect 8153 1340 8331 1437
rect 13222 1404 13292 1524
rect 13922 1487 14396 1524
rect 13922 1441 13955 1487
rect 14095 1441 14396 1487
rect 13922 1404 14396 1441
rect 14920 1404 14964 1524
rect 21153 1627 21262 1628
rect 21153 1524 21197 1627
rect 8153 1317 8266 1340
rect 6340 1213 6370 1317
rect 8224 1213 8266 1317
rect 6340 1198 6438 1213
rect 6275 1093 6438 1198
rect 7098 1093 7169 1213
rect 7423 1093 7493 1213
rect 8153 1200 8266 1213
rect 8312 1200 8331 1340
rect 18200 1365 18362 1437
rect 8153 1093 8331 1200
rect 8536 1093 8605 1213
rect 8923 1093 9195 1213
rect 9327 1179 9506 1213
rect 13222 1180 13292 1300
rect 13922 1180 14396 1300
rect 14920 1256 15220 1300
rect 14920 1210 15061 1256
rect 15201 1210 15220 1256
rect 14920 1180 15220 1210
rect 18200 1225 18219 1365
rect 18265 1317 18362 1365
rect 19462 1317 19588 1437
rect 20007 1404 20051 1524
rect 21051 1404 21197 1524
rect 18265 1225 18302 1317
rect 18200 1213 18302 1225
rect 19529 1268 19588 1317
rect 19529 1213 20051 1268
rect 9327 1133 9441 1179
rect 9487 1133 9506 1179
rect 9327 1093 9506 1133
rect 18200 1093 18362 1213
rect 19462 1148 20051 1213
rect 21051 1148 21095 1268
rect 21178 1205 21197 1404
rect 21243 1524 21262 1627
rect 21243 1404 21386 1524
rect 23386 1404 23430 1524
rect 21243 1300 21264 1404
rect 21243 1205 21386 1300
rect 21178 1180 21386 1205
rect 23386 1180 23430 1300
rect 19462 1093 19588 1148
rect 4730 652 4857 707
rect 889 500 933 620
rect 2933 565 3157 620
rect 2933 500 3092 565
rect 3055 396 3092 500
rect 889 276 933 396
rect 2933 276 3092 396
rect 3073 172 3092 276
rect 889 52 933 172
rect 2933 143 3092 172
rect 3138 396 3157 565
rect 3217 532 3268 652
rect 4268 587 4857 652
rect 5957 602 6137 707
rect 5957 587 6072 602
rect 4268 532 4789 587
rect 4730 483 4789 532
rect 6028 483 6072 587
rect 3138 276 3268 396
rect 4268 276 4312 396
rect 4730 363 4857 483
rect 5957 462 6072 483
rect 6118 462 6137 602
rect 5957 363 6137 462
rect 6275 602 6438 707
rect 6275 462 6294 602
rect 6340 587 6438 602
rect 7098 587 7169 707
rect 7423 587 7493 707
rect 8153 600 8331 707
rect 8153 587 8266 600
rect 6340 483 6370 587
rect 8224 483 8266 587
rect 6340 462 6438 483
rect 6275 363 6438 462
rect 7098 363 7169 483
rect 7423 363 7493 483
rect 8153 460 8266 483
rect 8312 460 8331 600
rect 8536 587 8605 707
rect 8923 587 9195 707
rect 9327 667 9506 707
rect 9327 621 9441 667
rect 9487 621 9506 667
rect 9327 587 9506 621
rect 13222 500 13292 620
rect 13922 500 14396 620
rect 14920 590 15220 620
rect 14920 544 15061 590
rect 15201 544 15220 590
rect 14920 500 15220 544
rect 18200 587 18362 707
rect 19462 652 19588 707
rect 19462 587 20051 652
rect 18200 575 18302 587
rect 8153 363 8331 460
rect 18200 435 18219 575
rect 18265 483 18302 575
rect 19529 532 20051 587
rect 21051 532 21095 652
rect 21178 595 21386 620
rect 19529 483 19588 532
rect 18265 435 18362 483
rect 3138 172 3157 276
rect 13222 276 13292 396
rect 13922 359 14396 396
rect 13922 313 13955 359
rect 14095 313 14396 359
rect 13922 276 14396 313
rect 14920 276 14964 396
rect 18200 363 18362 435
rect 19462 363 19588 483
rect 21178 396 21197 595
rect 9859 236 9943 255
rect 9859 190 9878 236
rect 9924 190 9943 236
rect 9859 172 9943 190
rect 20007 276 20051 396
rect 21051 276 21197 396
rect 3138 143 3268 172
rect 2933 52 3268 143
rect 4268 52 4312 172
rect 9254 52 9324 172
rect 9764 52 9943 172
rect 12951 164 13292 183
rect 12951 118 12970 164
rect 13110 118 13292 164
rect 12951 63 13292 118
rect 13922 172 14149 183
rect 13922 63 14396 172
rect 14048 52 14396 63
rect 14920 52 14990 172
rect 21153 173 21197 276
rect 21243 500 21386 595
rect 23386 500 23430 620
rect 21243 396 21264 500
rect 21243 276 21386 396
rect 23386 276 23430 396
rect 21243 173 21262 276
rect 21153 172 21262 173
rect 20007 52 20051 172
rect 21051 52 21386 172
rect 23386 52 23430 172
<< polycontact >>
rect 3092 13835 3138 14257
rect 12970 14236 13110 14282
rect 9878 14164 9924 14210
rect 6072 13798 6118 13938
rect 6294 13798 6340 13938
rect 13955 14041 14095 14087
rect 8266 13800 8312 13940
rect 15061 13810 15201 13856
rect 18219 13825 18265 13965
rect 9441 13733 9487 13779
rect 21197 13805 21243 14227
rect 3092 12743 3138 13165
rect 6072 13062 6118 13202
rect 6294 13062 6340 13202
rect 8266 13060 8312 13200
rect 9441 13221 9487 13267
rect 15061 13144 15201 13190
rect 18219 13035 18265 13175
rect 13955 12913 14095 12959
rect 9878 12790 9924 12836
rect 3092 12035 3138 12457
rect 12970 12718 13110 12764
rect 21197 12773 21243 13195
rect 12970 12436 13110 12482
rect 9878 12364 9924 12410
rect 6072 11998 6118 12138
rect 6294 11998 6340 12138
rect 13955 12241 14095 12287
rect 8266 12000 8312 12140
rect 15061 12010 15201 12056
rect 18219 12025 18265 12165
rect 9441 11933 9487 11979
rect 21197 12005 21243 12427
rect 3092 10943 3138 11365
rect 6072 11262 6118 11402
rect 6294 11262 6340 11402
rect 8266 11260 8312 11400
rect 9441 11421 9487 11467
rect 15061 11344 15201 11390
rect 18219 11235 18265 11375
rect 13955 11113 14095 11159
rect 9878 10990 9924 11036
rect 3092 10235 3138 10657
rect 12970 10918 13110 10964
rect 21197 10973 21243 11395
rect 12970 10636 13110 10682
rect 9878 10564 9924 10610
rect 6072 10198 6118 10338
rect 6294 10198 6340 10338
rect 13955 10441 14095 10487
rect 8266 10200 8312 10340
rect 15061 10210 15201 10256
rect 18219 10225 18265 10365
rect 9441 10133 9487 10179
rect 21197 10205 21243 10627
rect 3092 9143 3138 9565
rect 6072 9462 6118 9602
rect 6294 9462 6340 9602
rect 8266 9460 8312 9600
rect 9441 9621 9487 9667
rect 15061 9544 15201 9590
rect 18219 9435 18265 9575
rect 13955 9313 14095 9359
rect 9878 9190 9924 9236
rect 3092 8435 3138 8857
rect 12970 9118 13110 9164
rect 21197 9173 21243 9595
rect 12970 8836 13110 8882
rect 9878 8764 9924 8810
rect 6072 8398 6118 8538
rect 6294 8398 6340 8538
rect 13955 8641 14095 8687
rect 8266 8400 8312 8540
rect 15061 8410 15201 8456
rect 18219 8425 18265 8565
rect 9441 8333 9487 8379
rect 21197 8405 21243 8827
rect 3092 7343 3138 7765
rect 6072 7662 6118 7802
rect 6294 7662 6340 7802
rect 8266 7660 8312 7800
rect 9441 7821 9487 7867
rect 15061 7744 15201 7790
rect 18219 7635 18265 7775
rect 13955 7513 14095 7559
rect 9878 7390 9924 7436
rect 3092 6635 3138 7057
rect 12970 7318 13110 7364
rect 21197 7373 21243 7795
rect 12970 7036 13110 7082
rect 9878 6964 9924 7010
rect 6072 6598 6118 6738
rect 6294 6598 6340 6738
rect 13955 6841 14095 6887
rect 8266 6600 8312 6740
rect 15061 6610 15201 6656
rect 18219 6625 18265 6765
rect 9441 6533 9487 6579
rect 21197 6605 21243 7027
rect 3092 5543 3138 5965
rect 6072 5862 6118 6002
rect 6294 5862 6340 6002
rect 8266 5860 8312 6000
rect 9441 6021 9487 6067
rect 15061 5944 15201 5990
rect 18219 5835 18265 5975
rect 13955 5713 14095 5759
rect 9878 5590 9924 5636
rect 3092 4835 3138 5257
rect 12970 5518 13110 5564
rect 21197 5573 21243 5995
rect 12970 5236 13110 5282
rect 9878 5164 9924 5210
rect 6072 4798 6118 4938
rect 6294 4798 6340 4938
rect 13955 5041 14095 5087
rect 8266 4800 8312 4940
rect 15061 4810 15201 4856
rect 18219 4825 18265 4965
rect 9441 4733 9487 4779
rect 21197 4805 21243 5227
rect 3092 3743 3138 4165
rect 6072 4062 6118 4202
rect 6294 4062 6340 4202
rect 8266 4060 8312 4200
rect 9441 4221 9487 4267
rect 15061 4144 15201 4190
rect 18219 4035 18265 4175
rect 13955 3913 14095 3959
rect 9878 3790 9924 3836
rect 3092 3035 3138 3457
rect 12970 3718 13110 3764
rect 21197 3773 21243 4195
rect 12970 3436 13110 3482
rect 9878 3364 9924 3410
rect 6072 2998 6118 3138
rect 6294 2998 6340 3138
rect 13955 3241 14095 3287
rect 8266 3000 8312 3140
rect 15061 3010 15201 3056
rect 18219 3025 18265 3165
rect 9441 2933 9487 2979
rect 21197 3005 21243 3427
rect 3092 1943 3138 2365
rect 6072 2262 6118 2402
rect 6294 2262 6340 2402
rect 8266 2260 8312 2400
rect 9441 2421 9487 2467
rect 15061 2344 15201 2390
rect 18219 2235 18265 2375
rect 13955 2113 14095 2159
rect 9878 1990 9924 2036
rect 3092 1235 3138 1657
rect 12970 1918 13110 1964
rect 21197 1973 21243 2395
rect 12970 1636 13110 1682
rect 9878 1564 9924 1610
rect 6072 1198 6118 1338
rect 6294 1198 6340 1338
rect 13955 1441 14095 1487
rect 8266 1200 8312 1340
rect 15061 1210 15201 1256
rect 18219 1225 18265 1365
rect 9441 1133 9487 1179
rect 21197 1205 21243 1627
rect 3092 143 3138 565
rect 6072 462 6118 602
rect 6294 462 6340 602
rect 8266 460 8312 600
rect 9441 621 9487 667
rect 15061 544 15201 590
rect 18219 435 18265 575
rect 13955 313 14095 359
rect 9878 190 9924 236
rect 12970 118 13110 164
rect 21197 173 21243 595
<< metal1 >>
rect 345 14426 2439 14467
rect 3844 14460 4605 14466
rect 345 14374 451 14426
rect 503 14374 662 14426
rect 714 14374 873 14426
rect 925 14423 1083 14426
rect 1135 14423 1294 14426
rect 1346 14423 1506 14426
rect 1558 14423 1717 14426
rect 1769 14423 1927 14426
rect 1979 14423 2138 14426
rect 2190 14423 2349 14426
rect 2401 14423 2439 14426
rect 3843 14426 4605 14460
rect 3843 14423 3881 14426
rect 3933 14423 4092 14426
rect 4144 14423 4304 14426
rect 925 14377 946 14423
rect 2920 14377 2933 14423
rect 3268 14377 3281 14423
rect 3327 14377 3384 14423
rect 3430 14377 3487 14423
rect 3533 14377 3590 14423
rect 3636 14377 3693 14423
rect 3739 14377 3796 14423
rect 3842 14377 3881 14423
rect 3945 14377 4002 14423
rect 4048 14377 4092 14423
rect 4151 14377 4209 14423
rect 4255 14377 4304 14423
rect 925 14374 1083 14377
rect 1135 14374 1294 14377
rect 1346 14374 1506 14377
rect 1558 14374 1717 14377
rect 1769 14374 1927 14377
rect 1979 14374 2138 14377
rect 2190 14374 2349 14377
rect 2401 14374 2439 14377
rect 345 14333 2439 14374
rect 3843 14374 3881 14377
rect 3933 14374 4092 14377
rect 4144 14374 4304 14377
rect 4356 14374 4515 14426
rect 4567 14374 4605 14426
rect 3843 14340 4605 14374
rect 3844 14333 4605 14340
rect 4779 14460 5961 14467
rect 7543 14466 7921 14467
rect 4779 14426 6555 14460
rect 4779 14374 4817 14426
rect 4869 14374 5027 14426
rect 5079 14374 5238 14426
rect 5290 14374 5450 14426
rect 5502 14374 5661 14426
rect 5713 14374 5871 14426
rect 5923 14423 6555 14426
rect 5923 14377 6086 14423
rect 6320 14377 6555 14423
rect 5923 14374 6555 14377
rect 4779 14340 6555 14374
rect 7543 14426 8439 14466
rect 7543 14423 7927 14426
rect 7979 14423 8138 14426
rect 7543 14377 7554 14423
rect 8070 14377 8138 14423
rect 7543 14374 7927 14377
rect 7979 14374 8138 14377
rect 8190 14374 8349 14426
rect 8401 14374 8439 14426
rect 4779 14333 5961 14340
rect 7543 14333 8439 14374
rect 8611 14460 8919 14467
rect 9812 14460 10120 14467
rect 10385 14460 12583 14474
rect 13350 14460 14111 14466
rect 8611 14426 8920 14460
rect 8611 14374 8649 14426
rect 8701 14423 8829 14426
rect 8705 14377 8817 14423
rect 8701 14374 8829 14377
rect 8881 14374 8920 14426
rect 345 14299 637 14333
rect 345 14253 452 14299
rect 498 14253 637 14299
rect 345 14135 637 14253
rect 3081 14257 3149 14268
rect 2616 14202 2924 14243
rect 2616 14199 2654 14202
rect 2706 14199 2834 14202
rect 2886 14199 2924 14202
rect 933 14153 946 14199
rect 2920 14153 2933 14199
rect 345 14089 452 14135
rect 498 14089 637 14135
rect 2616 14150 2654 14153
rect 2706 14150 2834 14153
rect 2886 14150 2924 14153
rect 2616 14110 2924 14150
rect 345 13997 637 14089
rect 345 13975 1090 13997
rect 345 13972 946 13975
rect 345 13926 452 13972
rect 498 13929 946 13972
rect 2920 13929 2933 13975
rect 498 13926 1090 13929
rect 345 13878 1090 13926
rect 345 13809 637 13878
rect 345 13763 452 13809
rect 498 13763 637 13809
rect 3081 13835 3092 14257
rect 3138 13835 3149 14257
rect 3378 14210 3686 14251
rect 3378 14199 3416 14210
rect 3468 14199 3596 14210
rect 3648 14199 3686 14210
rect 3268 14153 3281 14199
rect 3327 14153 3384 14199
rect 3468 14158 3487 14199
rect 3430 14153 3487 14158
rect 3533 14153 3590 14199
rect 3648 14158 3693 14199
rect 3636 14153 3693 14158
rect 3739 14153 3796 14199
rect 3842 14153 3899 14199
rect 3945 14153 4002 14199
rect 4048 14153 4105 14199
rect 4151 14153 4209 14199
rect 4255 14153 4268 14199
rect 3378 14118 3686 14153
rect 4891 14124 5863 14164
rect 7450 14161 7758 14177
rect 4891 14112 4929 14124
rect 4981 14112 5140 14124
rect 5192 14112 5351 14124
rect 5403 14112 5562 14124
rect 5614 14112 5773 14124
rect 5825 14112 5863 14124
rect 6035 14112 6550 14161
rect 7036 14136 7758 14161
rect 7036 14112 7488 14136
rect 7540 14112 7668 14136
rect 7720 14112 7758 14136
rect 4857 14066 4870 14112
rect 5120 14072 5140 14112
rect 5120 14066 5177 14072
rect 5223 14066 5280 14112
rect 5326 14072 5351 14112
rect 5326 14066 5383 14072
rect 5429 14066 5486 14112
rect 5532 14072 5562 14112
rect 5532 14066 5589 14072
rect 5635 14066 5692 14112
rect 5738 14072 5773 14112
rect 5738 14066 5795 14072
rect 5841 14066 5898 14112
rect 5944 14066 5957 14112
rect 6035 14066 6451 14112
rect 6497 14066 6568 14112
rect 6614 14066 6685 14112
rect 6731 14066 6803 14112
rect 6849 14066 6921 14112
rect 6967 14066 7039 14112
rect 7085 14084 7488 14112
rect 7085 14066 7506 14084
rect 7552 14066 7623 14112
rect 7720 14084 7740 14112
rect 7669 14066 7740 14084
rect 7786 14066 7858 14112
rect 7904 14066 7976 14112
rect 8022 14066 8094 14112
rect 8140 14066 8153 14112
rect 4891 14032 5863 14066
rect 6035 14041 6550 14066
rect 7036 14044 7758 14066
rect 7036 14041 7528 14044
rect 3825 13975 4315 14004
rect 3268 13929 3281 13975
rect 3327 13929 3384 13975
rect 3430 13929 3487 13975
rect 3533 13929 3590 13975
rect 3636 13929 3693 13975
rect 3739 13929 3796 13975
rect 3842 13964 3899 13975
rect 3842 13929 3864 13964
rect 3945 13929 4002 13975
rect 4048 13964 4105 13975
rect 4096 13929 4105 13964
rect 4151 13929 4209 13975
rect 4255 13964 4315 13975
rect 3825 13912 3864 13929
rect 3916 13912 4044 13929
rect 4096 13912 4224 13929
rect 4276 13912 4315 13964
rect 6035 13938 6151 14041
rect 3825 13871 4315 13912
rect 4561 13888 5957 13932
rect 345 13646 637 13763
rect 2616 13754 2924 13795
rect 2616 13751 2654 13754
rect 2706 13751 2834 13754
rect 2886 13751 2924 13754
rect 3081 13753 3149 13835
rect 4561 13842 4870 13888
rect 5120 13842 5177 13888
rect 5223 13842 5280 13888
rect 5326 13842 5383 13888
rect 5429 13842 5486 13888
rect 5532 13842 5589 13888
rect 5635 13842 5692 13888
rect 5738 13842 5795 13888
rect 5841 13842 5898 13888
rect 5944 13842 5957 13888
rect 4561 13810 5957 13842
rect 4561 13753 4679 13810
rect 933 13705 946 13751
rect 2920 13705 2933 13751
rect 3081 13716 4679 13753
rect 2616 13702 2654 13705
rect 2706 13702 2834 13705
rect 2886 13702 2924 13705
rect 2616 13662 2924 13702
rect 3081 13670 3413 13716
rect 3459 13670 3599 13716
rect 3645 13670 3786 13716
rect 3832 13670 3973 13716
rect 4019 13670 4159 13716
rect 4205 13670 4679 13716
rect 6035 13798 6072 13938
rect 6118 13798 6151 13938
rect 3081 13662 4679 13670
rect 4891 13664 5863 13704
rect 6035 13698 6151 13798
rect 6237 13938 6370 13961
rect 6237 13889 6294 13938
rect 6237 13837 6275 13889
rect 6237 13798 6294 13837
rect 6340 13798 6370 13938
rect 8255 13940 8323 13951
rect 6521 13930 7282 13936
rect 6520 13929 7282 13930
rect 6520 13896 7528 13929
rect 6520 13888 6558 13896
rect 6610 13888 6769 13896
rect 6821 13888 6981 13896
rect 6438 13842 6451 13888
rect 6497 13844 6558 13888
rect 6497 13842 6568 13844
rect 6614 13842 6685 13888
rect 6731 13844 6769 13888
rect 6731 13842 6803 13844
rect 6849 13842 6921 13888
rect 6967 13844 6981 13888
rect 7033 13888 7192 13896
rect 7033 13844 7039 13888
rect 6967 13842 7039 13844
rect 7085 13844 7192 13888
rect 7244 13888 7528 13896
rect 7244 13844 7506 13888
rect 7085 13842 7506 13844
rect 7552 13842 7623 13888
rect 7669 13842 7740 13888
rect 7786 13842 7858 13888
rect 7904 13842 7976 13888
rect 8022 13842 8094 13888
rect 8140 13842 8153 13888
rect 6520 13810 7528 13842
rect 6521 13803 7282 13810
rect 6237 13778 6370 13798
rect 8255 13800 8266 13940
rect 8312 13800 8323 13940
rect 8611 13888 8920 14374
rect 9089 14437 12583 14460
rect 13301 14437 14111 14460
rect 9089 14426 14111 14437
rect 9089 14423 9850 14426
rect 9089 14377 9337 14423
rect 9383 14377 9459 14423
rect 9505 14377 9582 14423
rect 9628 14377 9705 14423
rect 9751 14377 9850 14423
rect 9089 14374 9850 14377
rect 9902 14374 10030 14426
rect 10082 14423 13387 14426
rect 10082 14377 10433 14423
rect 10479 14377 10591 14423
rect 10637 14377 10749 14423
rect 10795 14377 10907 14423
rect 10953 14377 11066 14423
rect 11112 14377 11224 14423
rect 11270 14377 11382 14423
rect 11428 14377 11540 14423
rect 11586 14377 11698 14423
rect 11744 14377 11856 14423
rect 11902 14377 12015 14423
rect 12061 14377 12173 14423
rect 12219 14377 12331 14423
rect 12377 14377 12489 14423
rect 12535 14377 13336 14423
rect 13382 14377 13387 14423
rect 10082 14374 13387 14377
rect 13439 14423 13598 14426
rect 13439 14377 13503 14423
rect 13549 14377 13598 14423
rect 13439 14374 13598 14377
rect 13650 14423 13810 14426
rect 13862 14423 14021 14426
rect 13650 14377 13668 14423
rect 13714 14377 13810 14423
rect 13879 14377 14021 14423
rect 13650 14374 13810 14377
rect 13862 14374 14021 14377
rect 14073 14374 14111 14426
rect 9089 14363 14111 14374
rect 9089 14340 12583 14363
rect 13301 14340 14111 14363
rect 9089 13888 9205 14340
rect 9812 14334 10120 14340
rect 10385 14326 12583 14340
rect 13350 14333 14111 14340
rect 14393 14460 14943 14466
rect 18397 14460 19579 14467
rect 19905 14460 20456 14467
rect 14393 14426 19579 14460
rect 14393 14423 14431 14426
rect 14483 14423 14642 14426
rect 14694 14423 14853 14426
rect 14905 14423 18435 14426
rect 14393 14377 14409 14423
rect 14483 14377 14522 14423
rect 14568 14377 14635 14423
rect 14694 14377 14748 14423
rect 14794 14377 14853 14423
rect 14907 14377 15216 14423
rect 15262 14377 15374 14423
rect 15420 14377 15532 14423
rect 15578 14377 15690 14423
rect 15736 14377 15848 14423
rect 15894 14377 16006 14423
rect 16052 14377 16165 14423
rect 16211 14377 16323 14423
rect 16369 14377 16481 14423
rect 16527 14377 16639 14423
rect 16685 14377 16797 14423
rect 16843 14377 16955 14423
rect 17001 14377 17113 14423
rect 17159 14377 17272 14423
rect 17318 14377 17430 14423
rect 17476 14377 17588 14423
rect 17634 14377 17746 14423
rect 17792 14377 17904 14423
rect 17950 14377 18062 14423
rect 18108 14377 18435 14423
rect 14393 14374 14431 14377
rect 14483 14374 14642 14377
rect 14694 14374 14853 14377
rect 14905 14374 18435 14377
rect 18487 14374 18645 14426
rect 18697 14374 18856 14426
rect 18908 14374 19068 14426
rect 19120 14374 19279 14426
rect 19331 14374 19489 14426
rect 19541 14374 19579 14426
rect 14393 14340 19579 14374
rect 19904 14426 20456 14460
rect 19904 14374 19943 14426
rect 19995 14423 20154 14426
rect 20206 14423 20365 14426
rect 20417 14423 20456 14426
rect 21875 14426 23974 14467
rect 21875 14423 21913 14426
rect 21965 14423 22124 14426
rect 22176 14423 22335 14426
rect 22387 14423 22545 14426
rect 22597 14423 22756 14426
rect 22808 14423 22968 14426
rect 23020 14423 23179 14426
rect 23231 14423 23389 14426
rect 19995 14377 20064 14423
rect 20110 14377 20154 14423
rect 20214 14377 20271 14423
rect 20317 14377 20365 14423
rect 20420 14377 20477 14423
rect 20523 14377 20580 14423
rect 20626 14377 20683 14423
rect 20729 14377 20786 14423
rect 20832 14377 20889 14423
rect 20935 14377 20992 14423
rect 21038 14377 21051 14423
rect 21386 14377 21399 14423
rect 23373 14377 23389 14423
rect 19995 14374 20154 14377
rect 20206 14374 20365 14377
rect 20417 14374 20456 14377
rect 19904 14340 20456 14374
rect 14393 14333 14943 14340
rect 12959 14282 13121 14293
rect 9334 14199 9463 14228
rect 9843 14210 9959 14247
rect 12959 14236 12970 14282
rect 13110 14236 13121 14282
rect 12959 14229 13121 14236
rect 9324 14153 9337 14199
rect 9383 14188 9459 14199
rect 9424 14153 9459 14188
rect 9505 14153 9582 14199
rect 9628 14153 9705 14199
rect 9751 14153 9764 14199
rect 9843 14164 9878 14210
rect 9924 14164 9959 14210
rect 9334 14136 9372 14153
rect 9424 14136 9463 14153
rect 9334 14109 9463 14136
rect 9334 14096 9462 14109
rect 9520 13973 9682 14013
rect 9520 13921 9591 13973
rect 9643 13921 9682 13973
rect 8605 13842 8618 13888
rect 8664 13842 8741 13888
rect 8787 13842 8864 13888
rect 8910 13842 8923 13888
rect 9089 13842 9238 13888
rect 9284 13842 9327 13888
rect 8611 13810 8920 13842
rect 9089 13810 9205 13842
rect 7450 13698 7758 13703
rect 6035 13664 6550 13698
rect 7036 13664 7758 13698
rect 8255 13678 8323 13800
rect 9520 13790 9682 13921
rect 9406 13787 9682 13790
rect 9406 13779 9591 13787
rect 9406 13733 9441 13779
rect 9487 13735 9591 13779
rect 9643 13766 9682 13787
rect 9843 13766 9959 14164
rect 10315 14188 13121 14229
rect 15181 14259 18143 14340
rect 18397 14333 19579 14340
rect 19905 14333 20456 14340
rect 21875 14374 21913 14377
rect 21965 14374 22124 14377
rect 22176 14374 22335 14377
rect 22387 14374 22545 14377
rect 22597 14374 22756 14377
rect 22808 14374 22968 14377
rect 23020 14374 23179 14377
rect 23231 14374 23389 14377
rect 23441 14374 23600 14426
rect 23652 14374 23811 14426
rect 23863 14374 23974 14426
rect 21875 14333 23974 14374
rect 15181 14213 15216 14259
rect 15262 14213 15374 14259
rect 15420 14213 15532 14259
rect 15578 14213 15690 14259
rect 15736 14213 15848 14259
rect 15894 14213 16006 14259
rect 16052 14213 16165 14259
rect 16211 14213 16323 14259
rect 16369 14213 16481 14259
rect 16527 14213 16639 14259
rect 16685 14213 16797 14259
rect 16843 14213 16955 14259
rect 17001 14213 17113 14259
rect 17159 14213 17272 14259
rect 17318 14213 17430 14259
rect 17476 14213 17588 14259
rect 17634 14213 17746 14259
rect 17792 14213 17904 14259
rect 17950 14213 18062 14259
rect 18108 14213 18143 14259
rect 23682 14299 23974 14333
rect 23682 14253 23820 14299
rect 23866 14253 23974 14299
rect 10315 14136 11532 14188
rect 11584 14136 13121 14188
rect 10315 14095 13121 14136
rect 14202 14153 14409 14199
rect 14455 14153 14522 14199
rect 14568 14153 14635 14199
rect 14681 14153 14748 14199
rect 14794 14153 14861 14199
rect 14907 14153 14920 14199
rect 15181 14177 18143 14213
rect 20632 14202 20940 14243
rect 20632 14199 20670 14202
rect 20722 14199 20850 14202
rect 20902 14199 20940 14202
rect 21186 14227 21254 14238
rect 13938 14087 14106 14098
rect 13938 14041 13955 14087
rect 14095 14041 14106 14087
rect 13938 13997 14106 14041
rect 11826 13957 14106 13997
rect 11826 13905 12665 13957
rect 12717 13905 14106 13957
rect 11826 13864 14106 13905
rect 14202 13766 14318 14153
rect 18502 14127 19474 14167
rect 20051 14153 20064 14199
rect 20110 14153 20168 14199
rect 20214 14153 20271 14199
rect 20317 14153 20374 14199
rect 20420 14153 20477 14199
rect 20523 14153 20580 14199
rect 20626 14153 20670 14199
rect 20729 14153 20786 14199
rect 20832 14153 20850 14199
rect 20935 14153 20992 14199
rect 21038 14153 21051 14199
rect 18502 14112 18540 14127
rect 18592 14112 18751 14127
rect 18803 14112 18962 14127
rect 19014 14112 19173 14127
rect 19225 14112 19384 14127
rect 19436 14112 19474 14127
rect 18362 14066 18375 14112
rect 18421 14066 18478 14112
rect 18524 14075 18540 14112
rect 18524 14066 18581 14075
rect 18627 14066 18684 14112
rect 18730 14075 18751 14112
rect 18730 14066 18787 14075
rect 18833 14066 18890 14112
rect 18936 14075 18962 14112
rect 18936 14066 18993 14075
rect 19039 14066 19096 14112
rect 19142 14075 19173 14112
rect 19142 14066 19199 14075
rect 19449 14066 19474 14112
rect 20632 14150 20670 14153
rect 20722 14150 20850 14153
rect 20902 14150 20940 14153
rect 20632 14110 20940 14150
rect 18154 14020 18284 14061
rect 18502 14035 19474 14066
rect 14498 13975 14838 14004
rect 14396 13929 14409 13975
rect 14455 13929 14522 13975
rect 14568 13964 14635 13975
rect 14588 13929 14635 13964
rect 14681 13929 14748 13975
rect 14794 13964 14861 13975
rect 14800 13929 14861 13964
rect 14907 13929 14920 13975
rect 18154 13968 18193 14020
rect 18245 13968 18284 14020
rect 18154 13965 18284 13968
rect 14498 13912 14536 13929
rect 14588 13912 14748 13929
rect 14800 13912 14838 13929
rect 14498 13871 14838 13912
rect 14997 13856 17976 13889
rect 14997 13810 15061 13856
rect 15201 13848 17976 13856
rect 14997 13796 15194 13810
rect 15246 13796 17976 13848
rect 9643 13751 14515 13766
rect 14997 13755 17976 13796
rect 18154 13825 18219 13965
rect 18265 13825 18284 13965
rect 19859 13975 20409 14004
rect 19859 13964 20064 13975
rect 20110 13964 20168 13975
rect 19417 13888 19757 13929
rect 18362 13842 18375 13888
rect 18421 13842 18478 13888
rect 18524 13842 18581 13888
rect 18627 13842 18684 13888
rect 18730 13842 18787 13888
rect 18833 13842 18890 13888
rect 18936 13842 18993 13888
rect 19039 13842 19096 13888
rect 19142 13842 19199 13888
rect 19449 13842 19757 13888
rect 19859 13912 19897 13964
rect 19949 13929 20064 13964
rect 20160 13929 20168 13964
rect 20214 13929 20271 13975
rect 20317 13964 20374 13975
rect 20317 13929 20319 13964
rect 19949 13912 20108 13929
rect 20160 13912 20319 13929
rect 20371 13929 20374 13964
rect 20420 13929 20477 13975
rect 20523 13929 20580 13975
rect 20626 13929 20683 13975
rect 20729 13929 20786 13975
rect 20832 13929 20889 13975
rect 20935 13929 20992 13975
rect 21038 13929 21051 13975
rect 20371 13912 20409 13929
rect 19859 13871 20409 13912
rect 18154 13802 18284 13825
rect 19417 13810 19757 13842
rect 9643 13735 14409 13751
rect 9487 13733 14409 13735
rect 9406 13730 14409 13733
rect 9406 13684 13336 13730
rect 13382 13684 13503 13730
rect 13549 13684 13668 13730
rect 13714 13684 13833 13730
rect 13879 13705 14409 13730
rect 14455 13705 14522 13751
rect 14568 13705 14635 13751
rect 14681 13705 14748 13751
rect 14794 13705 14861 13751
rect 14907 13705 14920 13751
rect 18154 13750 18193 13802
rect 18245 13750 18284 13802
rect 18154 13710 18284 13750
rect 19641 13753 19757 13810
rect 21186 13805 21197 14227
rect 21243 13805 21254 14227
rect 21394 14199 21702 14236
rect 21386 14153 21399 14199
rect 23373 14153 23386 14199
rect 21394 14143 21432 14153
rect 21484 14143 21612 14153
rect 21664 14143 21702 14153
rect 21394 14103 21702 14143
rect 23682 14135 23974 14253
rect 23682 14089 23820 14135
rect 23866 14089 23974 14135
rect 23682 13997 23974 14089
rect 23182 13975 23974 13997
rect 21386 13929 21399 13975
rect 23373 13929 23974 13975
rect 23182 13878 23974 13929
rect 21186 13753 21254 13805
rect 19641 13716 21254 13753
rect 21394 13751 21702 13773
rect 13879 13684 14515 13705
rect 8255 13664 9320 13678
rect 345 13600 452 13646
rect 498 13600 637 13646
rect 3081 13633 4240 13662
rect 4857 13618 4870 13664
rect 5120 13618 5140 13664
rect 5223 13618 5280 13664
rect 5326 13618 5351 13664
rect 5429 13618 5486 13664
rect 5532 13618 5562 13664
rect 5635 13618 5692 13664
rect 5738 13618 5773 13664
rect 5841 13618 5898 13664
rect 5944 13618 5957 13664
rect 6035 13618 6451 13664
rect 6497 13618 6568 13664
rect 6614 13618 6685 13664
rect 6731 13618 6803 13664
rect 6849 13618 6921 13664
rect 6967 13618 7039 13664
rect 7085 13662 7506 13664
rect 7085 13618 7488 13662
rect 7552 13618 7623 13664
rect 7669 13662 7740 13664
rect 7720 13618 7740 13662
rect 7786 13618 7858 13664
rect 7904 13618 7976 13664
rect 8022 13618 8094 13664
rect 8140 13618 8153 13664
rect 8255 13618 8618 13664
rect 8664 13618 8741 13664
rect 8787 13618 8864 13664
rect 8910 13618 9238 13664
rect 9284 13618 9327 13664
rect 9406 13646 14515 13684
rect 18502 13664 19474 13704
rect 18362 13618 18375 13664
rect 18421 13618 18478 13664
rect 18524 13618 18540 13664
rect 18627 13618 18684 13664
rect 18730 13618 18751 13664
rect 18833 13618 18890 13664
rect 18936 13618 18962 13664
rect 19039 13618 19096 13664
rect 19142 13618 19173 13664
rect 19449 13618 19474 13664
rect 19641 13670 20113 13716
rect 20159 13670 20300 13716
rect 20346 13670 20487 13716
rect 20533 13670 20673 13716
rect 20719 13670 20860 13716
rect 20906 13670 21254 13716
rect 21386 13705 21399 13751
rect 23373 13705 23386 13751
rect 19641 13660 21254 13670
rect 20078 13633 21254 13660
rect 21394 13680 21432 13705
rect 21484 13680 21612 13705
rect 21664 13680 21702 13705
rect 21394 13640 21702 13680
rect 23682 13646 23974 13878
rect 345 13567 637 13600
rect 4891 13612 4929 13618
rect 4981 13612 5140 13618
rect 5192 13612 5351 13618
rect 5403 13612 5562 13618
rect 5614 13612 5773 13618
rect 5825 13612 5863 13618
rect 4467 13567 4622 13574
rect 4891 13572 5863 13612
rect 6035 13578 6550 13618
rect 7036 13610 7488 13618
rect 7540 13610 7668 13618
rect 7720 13610 7758 13618
rect 7036 13578 7758 13610
rect 7450 13570 7758 13578
rect 345 13526 2439 13567
rect 345 13474 451 13526
rect 503 13474 662 13526
rect 714 13474 873 13526
rect 925 13474 1083 13526
rect 1135 13474 1294 13526
rect 1346 13474 1506 13526
rect 1558 13474 1717 13526
rect 1769 13474 1927 13526
rect 1979 13474 2138 13526
rect 2190 13474 2349 13526
rect 2401 13474 2439 13526
rect 345 13433 2439 13474
rect 4314 13526 4622 13567
rect 8255 13558 9320 13618
rect 18502 13612 18540 13618
rect 18592 13612 18751 13618
rect 18803 13612 18962 13618
rect 19014 13612 19173 13618
rect 19225 13612 19384 13618
rect 19436 13612 19474 13618
rect 18502 13572 19474 13612
rect 23682 13600 23820 13646
rect 23866 13600 23974 13646
rect 19696 13567 19852 13574
rect 23682 13567 23974 13600
rect 4314 13474 4352 13526
rect 4404 13523 4532 13526
rect 4404 13477 4513 13523
rect 4404 13474 4532 13477
rect 4584 13474 4622 13526
rect 4314 13433 4622 13474
rect 19696 13526 20005 13567
rect 19696 13474 19735 13526
rect 19787 13523 19915 13526
rect 19803 13477 19915 13523
rect 19787 13474 19915 13477
rect 19967 13474 20005 13526
rect 345 13400 637 13433
rect 4467 13426 4622 13433
rect 345 13354 452 13400
rect 498 13354 637 13400
rect 4891 13388 5863 13428
rect 7450 13422 7758 13430
rect 4891 13382 4929 13388
rect 4981 13382 5140 13388
rect 5192 13382 5351 13388
rect 5403 13382 5562 13388
rect 5614 13382 5773 13388
rect 5825 13382 5863 13388
rect 6035 13382 6550 13422
rect 7036 13390 7758 13422
rect 7036 13382 7488 13390
rect 7540 13382 7668 13390
rect 7720 13382 7758 13390
rect 8255 13382 9320 13442
rect 19696 13433 20005 13474
rect 21875 13526 23974 13567
rect 21875 13474 21913 13526
rect 21965 13474 22124 13526
rect 22176 13474 22335 13526
rect 22387 13474 22545 13526
rect 22597 13474 22756 13526
rect 22808 13474 22968 13526
rect 23020 13474 23179 13526
rect 23231 13474 23389 13526
rect 23441 13474 23600 13526
rect 23652 13474 23811 13526
rect 23863 13474 23974 13526
rect 21875 13433 23974 13474
rect 18502 13388 19474 13428
rect 19696 13426 19852 13433
rect 18502 13382 18540 13388
rect 18592 13382 18751 13388
rect 18803 13382 18962 13388
rect 19014 13382 19173 13388
rect 19225 13382 19384 13388
rect 19436 13382 19474 13388
rect 345 13237 637 13354
rect 3081 13338 4240 13367
rect 2616 13298 2924 13338
rect 2616 13295 2654 13298
rect 2706 13295 2834 13298
rect 2886 13295 2924 13298
rect 3081 13330 4679 13338
rect 4857 13336 4870 13382
rect 5120 13336 5140 13382
rect 5223 13336 5280 13382
rect 5326 13336 5351 13382
rect 5429 13336 5486 13382
rect 5532 13336 5562 13382
rect 5635 13336 5692 13382
rect 5738 13336 5773 13382
rect 5841 13336 5898 13382
rect 5944 13336 5957 13382
rect 6035 13336 6451 13382
rect 6497 13336 6568 13382
rect 6614 13336 6685 13382
rect 6731 13336 6803 13382
rect 6849 13336 6921 13382
rect 6967 13336 7039 13382
rect 7085 13338 7488 13382
rect 7085 13336 7506 13338
rect 7552 13336 7623 13382
rect 7720 13338 7740 13382
rect 7669 13336 7740 13338
rect 7786 13336 7858 13382
rect 7904 13336 7976 13382
rect 8022 13336 8094 13382
rect 8140 13336 8153 13382
rect 8255 13336 8618 13382
rect 8664 13336 8741 13382
rect 8787 13336 8864 13382
rect 8910 13336 9238 13382
rect 9284 13336 9327 13382
rect 933 13249 946 13295
rect 2920 13249 2933 13295
rect 3081 13284 3413 13330
rect 3459 13284 3599 13330
rect 3645 13284 3786 13330
rect 3832 13284 3973 13330
rect 4019 13284 4159 13330
rect 4205 13284 4679 13330
rect 4891 13296 5863 13336
rect 6035 13302 6550 13336
rect 7036 13302 7758 13336
rect 345 13191 452 13237
rect 498 13191 637 13237
rect 2616 13246 2654 13249
rect 2706 13246 2834 13249
rect 2886 13246 2924 13249
rect 2616 13205 2924 13246
rect 3081 13247 4679 13284
rect 345 13122 637 13191
rect 3081 13165 3149 13247
rect 345 13074 1090 13122
rect 345 13028 452 13074
rect 498 13071 1090 13074
rect 498 13028 946 13071
rect 345 13025 946 13028
rect 2920 13025 2933 13071
rect 345 13003 1090 13025
rect 345 12911 637 13003
rect 345 12865 452 12911
rect 498 12865 637 12911
rect 345 12747 637 12865
rect 2616 12850 2924 12890
rect 2616 12847 2654 12850
rect 2706 12847 2834 12850
rect 2886 12847 2924 12850
rect 933 12801 946 12847
rect 2920 12801 2933 12847
rect 2616 12798 2654 12801
rect 2706 12798 2834 12801
rect 2886 12798 2924 12801
rect 2616 12757 2924 12798
rect 345 12701 452 12747
rect 498 12701 637 12747
rect 3081 12743 3092 13165
rect 3138 12743 3149 13165
rect 4561 13190 4679 13247
rect 6035 13202 6151 13302
rect 7450 13297 7758 13302
rect 8255 13322 9320 13336
rect 4561 13158 5957 13190
rect 3825 13088 4315 13129
rect 3825 13071 3864 13088
rect 3916 13071 4044 13088
rect 4096 13071 4224 13088
rect 3268 13025 3281 13071
rect 3327 13025 3384 13071
rect 3430 13025 3487 13071
rect 3533 13025 3590 13071
rect 3636 13025 3693 13071
rect 3739 13025 3796 13071
rect 3842 13036 3864 13071
rect 3842 13025 3899 13036
rect 3945 13025 4002 13071
rect 4096 13036 4105 13071
rect 4048 13025 4105 13036
rect 4151 13025 4209 13071
rect 4276 13036 4315 13088
rect 4561 13112 4870 13158
rect 5120 13112 5177 13158
rect 5223 13112 5280 13158
rect 5326 13112 5383 13158
rect 5429 13112 5486 13158
rect 5532 13112 5589 13158
rect 5635 13112 5692 13158
rect 5738 13112 5795 13158
rect 5841 13112 5898 13158
rect 5944 13112 5957 13158
rect 4561 13068 5957 13112
rect 4255 13025 4315 13036
rect 3825 12996 4315 13025
rect 6035 13062 6072 13202
rect 6118 13062 6151 13202
rect 4891 12934 5863 12968
rect 6035 12959 6151 13062
rect 6237 13202 6370 13222
rect 6237 13163 6294 13202
rect 6237 13111 6275 13163
rect 6237 13062 6294 13111
rect 6340 13062 6370 13202
rect 8255 13200 8323 13322
rect 9406 13316 14515 13354
rect 18362 13336 18375 13382
rect 18421 13336 18478 13382
rect 18524 13336 18540 13382
rect 18627 13336 18684 13382
rect 18730 13336 18751 13382
rect 18833 13336 18890 13382
rect 18936 13336 18962 13382
rect 19039 13336 19096 13382
rect 19142 13336 19173 13382
rect 19449 13336 19474 13382
rect 23682 13400 23974 13433
rect 20078 13340 21254 13367
rect 9406 13270 13336 13316
rect 13382 13270 13503 13316
rect 13549 13270 13668 13316
rect 13714 13270 13833 13316
rect 13879 13295 14515 13316
rect 18502 13296 19474 13336
rect 19641 13330 21254 13340
rect 13879 13270 14409 13295
rect 9406 13267 14409 13270
rect 9406 13221 9441 13267
rect 9487 13265 14409 13267
rect 9487 13221 9591 13265
rect 9406 13213 9591 13221
rect 9643 13249 14409 13265
rect 14455 13249 14522 13295
rect 14568 13249 14635 13295
rect 14681 13249 14748 13295
rect 14794 13249 14861 13295
rect 14907 13249 14920 13295
rect 18154 13250 18284 13290
rect 9643 13234 14515 13249
rect 9643 13213 9682 13234
rect 9406 13210 9682 13213
rect 6521 13190 7282 13197
rect 6520 13158 7528 13190
rect 6438 13112 6451 13158
rect 6497 13156 6568 13158
rect 6497 13112 6558 13156
rect 6614 13112 6685 13158
rect 6731 13156 6803 13158
rect 6731 13112 6769 13156
rect 6849 13112 6921 13158
rect 6967 13156 7039 13158
rect 6967 13112 6981 13156
rect 6520 13104 6558 13112
rect 6610 13104 6769 13112
rect 6821 13104 6981 13112
rect 7033 13112 7039 13156
rect 7085 13156 7506 13158
rect 7085 13112 7192 13156
rect 7033 13104 7192 13112
rect 7244 13112 7506 13156
rect 7552 13112 7623 13158
rect 7669 13112 7740 13158
rect 7786 13112 7858 13158
rect 7904 13112 7976 13158
rect 8022 13112 8094 13158
rect 8140 13112 8153 13158
rect 7244 13104 7528 13112
rect 6520 13071 7528 13104
rect 6520 13070 7282 13071
rect 6521 13064 7282 13070
rect 6237 13039 6370 13062
rect 8255 13060 8266 13200
rect 8312 13060 8323 13200
rect 8611 13158 8920 13190
rect 9089 13158 9205 13190
rect 8605 13112 8618 13158
rect 8664 13112 8741 13158
rect 8787 13112 8864 13158
rect 8910 13112 8923 13158
rect 9089 13112 9238 13158
rect 9284 13112 9327 13158
rect 8255 13049 8323 13060
rect 6035 12934 6550 12959
rect 7036 12956 7528 12959
rect 7036 12934 7758 12956
rect 4857 12888 4870 12934
rect 5120 12928 5177 12934
rect 5120 12888 5140 12928
rect 5223 12888 5280 12934
rect 5326 12928 5383 12934
rect 5326 12888 5351 12928
rect 5429 12888 5486 12934
rect 5532 12928 5589 12934
rect 5532 12888 5562 12928
rect 5635 12888 5692 12934
rect 5738 12928 5795 12934
rect 5738 12888 5773 12928
rect 5841 12888 5898 12934
rect 5944 12888 5957 12934
rect 6035 12888 6451 12934
rect 6497 12888 6568 12934
rect 6614 12888 6685 12934
rect 6731 12888 6803 12934
rect 6849 12888 6921 12934
rect 6967 12888 7039 12934
rect 7085 12916 7506 12934
rect 7085 12888 7488 12916
rect 7552 12888 7623 12934
rect 7669 12916 7740 12934
rect 7720 12888 7740 12916
rect 7786 12888 7858 12934
rect 7904 12888 7976 12934
rect 8022 12888 8094 12934
rect 8140 12888 8153 12934
rect 3378 12847 3686 12882
rect 4891 12876 4929 12888
rect 4981 12876 5140 12888
rect 5192 12876 5351 12888
rect 5403 12876 5562 12888
rect 5614 12876 5773 12888
rect 5825 12876 5863 12888
rect 3268 12801 3281 12847
rect 3327 12801 3384 12847
rect 3430 12842 3487 12847
rect 3468 12801 3487 12842
rect 3533 12801 3590 12847
rect 3636 12842 3693 12847
rect 3648 12801 3693 12842
rect 3739 12801 3796 12847
rect 3842 12801 3899 12847
rect 3945 12801 4002 12847
rect 4048 12801 4105 12847
rect 4151 12801 4209 12847
rect 4255 12801 4268 12847
rect 4891 12836 5863 12876
rect 6035 12839 6550 12888
rect 7036 12864 7488 12888
rect 7540 12864 7668 12888
rect 7720 12864 7758 12888
rect 7036 12839 7758 12864
rect 7450 12823 7758 12839
rect 3378 12790 3416 12801
rect 3468 12790 3596 12801
rect 3648 12790 3686 12801
rect 3378 12749 3686 12790
rect 3081 12732 3149 12743
rect 345 12667 637 12701
rect 345 12626 2439 12667
rect 3844 12660 4605 12667
rect 345 12574 451 12626
rect 503 12574 662 12626
rect 714 12574 873 12626
rect 925 12623 1083 12626
rect 1135 12623 1294 12626
rect 1346 12623 1506 12626
rect 1558 12623 1717 12626
rect 1769 12623 1927 12626
rect 1979 12623 2138 12626
rect 2190 12623 2349 12626
rect 2401 12623 2439 12626
rect 3843 12626 4605 12660
rect 3843 12623 3881 12626
rect 3933 12623 4092 12626
rect 4144 12623 4304 12626
rect 925 12577 946 12623
rect 2920 12577 2933 12623
rect 3268 12577 3281 12623
rect 3327 12577 3384 12623
rect 3430 12577 3487 12623
rect 3533 12577 3590 12623
rect 3636 12577 3693 12623
rect 3739 12577 3796 12623
rect 3842 12577 3881 12623
rect 3945 12577 4002 12623
rect 4048 12577 4092 12623
rect 4151 12577 4209 12623
rect 4255 12577 4304 12623
rect 925 12574 1083 12577
rect 1135 12574 1294 12577
rect 1346 12574 1506 12577
rect 1558 12574 1717 12577
rect 1769 12574 1927 12577
rect 1979 12574 2138 12577
rect 2190 12574 2349 12577
rect 2401 12574 2439 12577
rect 345 12533 2439 12574
rect 3843 12574 3881 12577
rect 3933 12574 4092 12577
rect 4144 12574 4304 12577
rect 4356 12574 4515 12626
rect 4567 12574 4605 12626
rect 3843 12540 4605 12574
rect 3844 12533 4605 12540
rect 4779 12660 5961 12667
rect 4779 12626 6555 12660
rect 4779 12574 4817 12626
rect 4869 12574 5027 12626
rect 5079 12574 5238 12626
rect 5290 12574 5450 12626
rect 5502 12574 5661 12626
rect 5713 12574 5871 12626
rect 5923 12623 6555 12626
rect 5923 12577 6086 12623
rect 6320 12577 6555 12623
rect 5923 12574 6555 12577
rect 4779 12540 6555 12574
rect 7543 12626 8439 12667
rect 7543 12623 7927 12626
rect 7979 12623 8138 12626
rect 7543 12577 7554 12623
rect 8070 12577 8138 12623
rect 7543 12574 7927 12577
rect 7979 12574 8138 12577
rect 8190 12574 8349 12626
rect 8401 12574 8439 12626
rect 4779 12533 5961 12540
rect 7543 12533 8439 12574
rect 8611 12626 8920 13112
rect 8611 12574 8649 12626
rect 8701 12623 8829 12626
rect 8705 12577 8817 12623
rect 8701 12574 8829 12577
rect 8881 12574 8920 12626
rect 345 12499 637 12533
rect 345 12453 452 12499
rect 498 12453 637 12499
rect 345 12335 637 12453
rect 3081 12457 3149 12468
rect 2616 12402 2924 12443
rect 2616 12399 2654 12402
rect 2706 12399 2834 12402
rect 2886 12399 2924 12402
rect 933 12353 946 12399
rect 2920 12353 2933 12399
rect 345 12289 452 12335
rect 498 12289 637 12335
rect 2616 12350 2654 12353
rect 2706 12350 2834 12353
rect 2886 12350 2924 12353
rect 2616 12310 2924 12350
rect 345 12197 637 12289
rect 345 12175 1090 12197
rect 345 12172 946 12175
rect 345 12126 452 12172
rect 498 12129 946 12172
rect 2920 12129 2933 12175
rect 498 12126 1090 12129
rect 345 12078 1090 12126
rect 345 12009 637 12078
rect 345 11963 452 12009
rect 498 11963 637 12009
rect 3081 12035 3092 12457
rect 3138 12035 3149 12457
rect 3378 12410 3686 12451
rect 3378 12399 3416 12410
rect 3468 12399 3596 12410
rect 3648 12399 3686 12410
rect 3268 12353 3281 12399
rect 3327 12353 3384 12399
rect 3468 12358 3487 12399
rect 3430 12353 3487 12358
rect 3533 12353 3590 12399
rect 3648 12358 3693 12399
rect 3636 12353 3693 12358
rect 3739 12353 3796 12399
rect 3842 12353 3899 12399
rect 3945 12353 4002 12399
rect 4048 12353 4105 12399
rect 4151 12353 4209 12399
rect 4255 12353 4268 12399
rect 3378 12318 3686 12353
rect 4891 12324 5863 12364
rect 7450 12361 7758 12377
rect 4891 12312 4929 12324
rect 4981 12312 5140 12324
rect 5192 12312 5351 12324
rect 5403 12312 5562 12324
rect 5614 12312 5773 12324
rect 5825 12312 5863 12324
rect 6035 12312 6550 12361
rect 7036 12336 7758 12361
rect 7036 12312 7488 12336
rect 7540 12312 7668 12336
rect 7720 12312 7758 12336
rect 4857 12266 4870 12312
rect 5120 12272 5140 12312
rect 5120 12266 5177 12272
rect 5223 12266 5280 12312
rect 5326 12272 5351 12312
rect 5326 12266 5383 12272
rect 5429 12266 5486 12312
rect 5532 12272 5562 12312
rect 5532 12266 5589 12272
rect 5635 12266 5692 12312
rect 5738 12272 5773 12312
rect 5738 12266 5795 12272
rect 5841 12266 5898 12312
rect 5944 12266 5957 12312
rect 6035 12266 6451 12312
rect 6497 12266 6568 12312
rect 6614 12266 6685 12312
rect 6731 12266 6803 12312
rect 6849 12266 6921 12312
rect 6967 12266 7039 12312
rect 7085 12284 7488 12312
rect 7085 12266 7506 12284
rect 7552 12266 7623 12312
rect 7720 12284 7740 12312
rect 7669 12266 7740 12284
rect 7786 12266 7858 12312
rect 7904 12266 7976 12312
rect 8022 12266 8094 12312
rect 8140 12266 8153 12312
rect 4891 12232 5863 12266
rect 6035 12241 6550 12266
rect 7036 12244 7758 12266
rect 7036 12241 7528 12244
rect 3825 12175 4315 12204
rect 3268 12129 3281 12175
rect 3327 12129 3384 12175
rect 3430 12129 3487 12175
rect 3533 12129 3590 12175
rect 3636 12129 3693 12175
rect 3739 12129 3796 12175
rect 3842 12164 3899 12175
rect 3842 12129 3864 12164
rect 3945 12129 4002 12175
rect 4048 12164 4105 12175
rect 4096 12129 4105 12164
rect 4151 12129 4209 12175
rect 4255 12164 4315 12175
rect 3825 12112 3864 12129
rect 3916 12112 4044 12129
rect 4096 12112 4224 12129
rect 4276 12112 4315 12164
rect 6035 12138 6151 12241
rect 3825 12071 4315 12112
rect 4561 12088 5957 12132
rect 345 11846 637 11963
rect 2616 11954 2924 11995
rect 2616 11951 2654 11954
rect 2706 11951 2834 11954
rect 2886 11951 2924 11954
rect 3081 11953 3149 12035
rect 4561 12042 4870 12088
rect 5120 12042 5177 12088
rect 5223 12042 5280 12088
rect 5326 12042 5383 12088
rect 5429 12042 5486 12088
rect 5532 12042 5589 12088
rect 5635 12042 5692 12088
rect 5738 12042 5795 12088
rect 5841 12042 5898 12088
rect 5944 12042 5957 12088
rect 4561 12010 5957 12042
rect 4561 11953 4679 12010
rect 933 11905 946 11951
rect 2920 11905 2933 11951
rect 3081 11916 4679 11953
rect 2616 11902 2654 11905
rect 2706 11902 2834 11905
rect 2886 11902 2924 11905
rect 2616 11862 2924 11902
rect 3081 11870 3413 11916
rect 3459 11870 3599 11916
rect 3645 11870 3786 11916
rect 3832 11870 3973 11916
rect 4019 11870 4159 11916
rect 4205 11870 4679 11916
rect 6035 11998 6072 12138
rect 6118 11998 6151 12138
rect 3081 11862 4679 11870
rect 4891 11864 5863 11904
rect 6035 11898 6151 11998
rect 6237 12138 6370 12161
rect 6237 12089 6294 12138
rect 6237 12037 6275 12089
rect 6237 11998 6294 12037
rect 6340 11998 6370 12138
rect 8255 12140 8323 12151
rect 6521 12130 7282 12136
rect 6520 12129 7282 12130
rect 6520 12096 7528 12129
rect 6520 12088 6558 12096
rect 6610 12088 6769 12096
rect 6821 12088 6981 12096
rect 6438 12042 6451 12088
rect 6497 12044 6558 12088
rect 6497 12042 6568 12044
rect 6614 12042 6685 12088
rect 6731 12044 6769 12088
rect 6731 12042 6803 12044
rect 6849 12042 6921 12088
rect 6967 12044 6981 12088
rect 7033 12088 7192 12096
rect 7033 12044 7039 12088
rect 6967 12042 7039 12044
rect 7085 12044 7192 12088
rect 7244 12088 7528 12096
rect 7244 12044 7506 12088
rect 7085 12042 7506 12044
rect 7552 12042 7623 12088
rect 7669 12042 7740 12088
rect 7786 12042 7858 12088
rect 7904 12042 7976 12088
rect 8022 12042 8094 12088
rect 8140 12042 8153 12088
rect 6520 12010 7528 12042
rect 6521 12003 7282 12010
rect 6237 11978 6370 11998
rect 8255 12000 8266 12140
rect 8312 12000 8323 12140
rect 8611 12088 8920 12574
rect 9089 12660 9205 13112
rect 9520 13079 9682 13210
rect 9520 13027 9591 13079
rect 9643 13027 9682 13079
rect 9520 12987 9682 13027
rect 9334 12891 9462 12904
rect 9334 12864 9463 12891
rect 9334 12847 9372 12864
rect 9424 12847 9463 12864
rect 9324 12801 9337 12847
rect 9424 12812 9459 12847
rect 9383 12801 9459 12812
rect 9505 12801 9582 12847
rect 9628 12801 9705 12847
rect 9751 12801 9764 12847
rect 9843 12836 9959 13234
rect 11826 13095 14106 13136
rect 11826 13043 12665 13095
rect 12717 13043 14106 13095
rect 11826 13003 14106 13043
rect 13938 12959 14106 13003
rect 13938 12913 13955 12959
rect 14095 12913 14106 12959
rect 9334 12772 9463 12801
rect 9843 12790 9878 12836
rect 9924 12790 9959 12836
rect 9843 12753 9959 12790
rect 10315 12864 13121 12905
rect 13938 12902 14106 12913
rect 10315 12812 11532 12864
rect 11584 12812 13121 12864
rect 10315 12771 13121 12812
rect 14202 12847 14318 13234
rect 14997 13204 17976 13245
rect 14997 13190 15572 13204
rect 14997 13144 15061 13190
rect 15201 13152 15572 13190
rect 15624 13152 17976 13204
rect 15201 13144 17976 13152
rect 14498 13088 14838 13129
rect 14997 13111 17976 13144
rect 18154 13198 18193 13250
rect 18245 13198 18284 13250
rect 18154 13175 18284 13198
rect 19641 13284 20113 13330
rect 20159 13284 20300 13330
rect 20346 13284 20487 13330
rect 20533 13284 20673 13330
rect 20719 13284 20860 13330
rect 20906 13284 21254 13330
rect 21394 13320 21702 13360
rect 21394 13295 21432 13320
rect 21484 13295 21612 13320
rect 21664 13295 21702 13320
rect 23682 13354 23820 13400
rect 23866 13354 23974 13400
rect 19641 13247 21254 13284
rect 21386 13249 21399 13295
rect 23373 13249 23386 13295
rect 19641 13190 19757 13247
rect 14498 13071 14536 13088
rect 14588 13071 14748 13088
rect 14800 13071 14838 13088
rect 14396 13025 14409 13071
rect 14455 13025 14522 13071
rect 14588 13036 14635 13071
rect 14568 13025 14635 13036
rect 14681 13025 14748 13071
rect 14800 13036 14861 13071
rect 14794 13025 14861 13036
rect 14907 13025 14920 13071
rect 18154 13035 18219 13175
rect 18265 13035 18284 13175
rect 19417 13158 19757 13190
rect 18362 13112 18375 13158
rect 18421 13112 18478 13158
rect 18524 13112 18581 13158
rect 18627 13112 18684 13158
rect 18730 13112 18787 13158
rect 18833 13112 18890 13158
rect 18936 13112 18993 13158
rect 19039 13112 19096 13158
rect 19142 13112 19199 13158
rect 19449 13112 19757 13158
rect 21186 13195 21254 13247
rect 21394 13227 21702 13249
rect 19417 13071 19757 13112
rect 19859 13088 20409 13129
rect 18154 13032 18284 13035
rect 14498 12996 14838 13025
rect 18154 12980 18193 13032
rect 18245 12980 18284 13032
rect 19859 13036 19897 13088
rect 19949 13071 20108 13088
rect 20160 13071 20319 13088
rect 19949 13036 20064 13071
rect 20160 13036 20168 13071
rect 19859 13025 20064 13036
rect 20110 13025 20168 13036
rect 20214 13025 20271 13071
rect 20317 13036 20319 13071
rect 20371 13071 20409 13088
rect 20371 13036 20374 13071
rect 20317 13025 20374 13036
rect 20420 13025 20477 13071
rect 20523 13025 20580 13071
rect 20626 13025 20683 13071
rect 20729 13025 20786 13071
rect 20832 13025 20889 13071
rect 20935 13025 20992 13071
rect 21038 13025 21051 13071
rect 19859 12996 20409 13025
rect 18154 12939 18284 12980
rect 18502 12934 19474 12965
rect 18362 12888 18375 12934
rect 18421 12888 18478 12934
rect 18524 12925 18581 12934
rect 18524 12888 18540 12925
rect 18627 12888 18684 12934
rect 18730 12925 18787 12934
rect 18730 12888 18751 12925
rect 18833 12888 18890 12934
rect 18936 12925 18993 12934
rect 18936 12888 18962 12925
rect 19039 12888 19096 12934
rect 19142 12925 19199 12934
rect 19142 12888 19173 12925
rect 19449 12888 19474 12934
rect 18502 12873 18540 12888
rect 18592 12873 18751 12888
rect 18803 12873 18962 12888
rect 19014 12873 19173 12888
rect 19225 12873 19384 12888
rect 19436 12873 19474 12888
rect 14202 12801 14409 12847
rect 14455 12801 14522 12847
rect 14568 12801 14635 12847
rect 14681 12801 14748 12847
rect 14794 12801 14861 12847
rect 14907 12801 14920 12847
rect 18502 12833 19474 12873
rect 20632 12850 20940 12890
rect 20632 12847 20670 12850
rect 20722 12847 20850 12850
rect 20902 12847 20940 12850
rect 12959 12764 13121 12771
rect 12959 12718 12970 12764
rect 13110 12718 13121 12764
rect 12959 12707 13121 12718
rect 15181 12787 18143 12823
rect 20051 12801 20064 12847
rect 20110 12801 20168 12847
rect 20214 12801 20271 12847
rect 20317 12801 20374 12847
rect 20420 12801 20477 12847
rect 20523 12801 20580 12847
rect 20626 12801 20670 12847
rect 20729 12801 20786 12847
rect 20832 12801 20850 12847
rect 20935 12801 20992 12847
rect 21038 12801 21051 12847
rect 15181 12741 15216 12787
rect 15262 12741 15374 12787
rect 15420 12741 15532 12787
rect 15578 12741 15690 12787
rect 15736 12741 15848 12787
rect 15894 12741 16006 12787
rect 16052 12741 16165 12787
rect 16211 12741 16323 12787
rect 16369 12741 16481 12787
rect 16527 12741 16639 12787
rect 16685 12741 16797 12787
rect 16843 12741 16955 12787
rect 17001 12741 17113 12787
rect 17159 12741 17272 12787
rect 17318 12741 17430 12787
rect 17476 12741 17588 12787
rect 17634 12741 17746 12787
rect 17792 12741 17904 12787
rect 17950 12741 18062 12787
rect 18108 12741 18143 12787
rect 20632 12798 20670 12801
rect 20722 12798 20850 12801
rect 20902 12798 20940 12801
rect 20632 12757 20940 12798
rect 21186 12773 21197 13195
rect 21243 12773 21254 13195
rect 23682 13122 23974 13354
rect 23182 13071 23974 13122
rect 21386 13025 21399 13071
rect 23373 13025 23974 13071
rect 23182 13003 23974 13025
rect 23682 12911 23974 13003
rect 21394 12857 21702 12897
rect 21394 12847 21432 12857
rect 21484 12847 21612 12857
rect 21664 12847 21702 12857
rect 23682 12865 23820 12911
rect 23866 12865 23974 12911
rect 21386 12801 21399 12847
rect 23373 12801 23386 12847
rect 21186 12762 21254 12773
rect 21394 12764 21702 12801
rect 9812 12660 10120 12667
rect 10385 12660 12583 12674
rect 13350 12660 14111 12667
rect 9089 12637 12583 12660
rect 13301 12637 14111 12660
rect 9089 12626 14111 12637
rect 9089 12623 9850 12626
rect 9089 12577 9337 12623
rect 9383 12577 9459 12623
rect 9505 12577 9582 12623
rect 9628 12577 9705 12623
rect 9751 12577 9850 12623
rect 9089 12574 9850 12577
rect 9902 12574 10030 12626
rect 10082 12623 13387 12626
rect 10082 12577 10433 12623
rect 10479 12577 10591 12623
rect 10637 12577 10749 12623
rect 10795 12577 10907 12623
rect 10953 12577 11066 12623
rect 11112 12577 11224 12623
rect 11270 12577 11382 12623
rect 11428 12577 11540 12623
rect 11586 12577 11698 12623
rect 11744 12577 11856 12623
rect 11902 12577 12015 12623
rect 12061 12577 12173 12623
rect 12219 12577 12331 12623
rect 12377 12577 12489 12623
rect 12535 12577 13336 12623
rect 13382 12577 13387 12623
rect 10082 12574 13387 12577
rect 13439 12623 13598 12626
rect 13439 12577 13503 12623
rect 13549 12577 13598 12623
rect 13439 12574 13598 12577
rect 13650 12623 13810 12626
rect 13862 12623 14021 12626
rect 13650 12577 13668 12623
rect 13714 12577 13810 12623
rect 13879 12577 14021 12623
rect 13650 12574 13810 12577
rect 13862 12574 14021 12577
rect 14073 12574 14111 12626
rect 9089 12563 14111 12574
rect 9089 12540 12583 12563
rect 13301 12540 14111 12563
rect 9089 12088 9205 12540
rect 9812 12533 10120 12540
rect 10385 12526 12583 12540
rect 13350 12533 14111 12540
rect 14393 12660 14943 12667
rect 15181 12660 18143 12741
rect 23682 12747 23974 12865
rect 23682 12701 23820 12747
rect 23866 12701 23974 12747
rect 23682 12667 23974 12701
rect 18397 12660 19579 12667
rect 19905 12660 20456 12667
rect 14393 12626 19579 12660
rect 14393 12623 14431 12626
rect 14483 12623 14642 12626
rect 14694 12623 14853 12626
rect 14905 12623 18435 12626
rect 14393 12577 14409 12623
rect 14483 12577 14522 12623
rect 14568 12577 14635 12623
rect 14694 12577 14748 12623
rect 14794 12577 14853 12623
rect 14907 12577 15216 12623
rect 15262 12577 15374 12623
rect 15420 12577 15532 12623
rect 15578 12577 15690 12623
rect 15736 12577 15848 12623
rect 15894 12577 16006 12623
rect 16052 12577 16165 12623
rect 16211 12577 16323 12623
rect 16369 12577 16481 12623
rect 16527 12577 16639 12623
rect 16685 12577 16797 12623
rect 16843 12577 16955 12623
rect 17001 12577 17113 12623
rect 17159 12577 17272 12623
rect 17318 12577 17430 12623
rect 17476 12577 17588 12623
rect 17634 12577 17746 12623
rect 17792 12577 17904 12623
rect 17950 12577 18062 12623
rect 18108 12577 18435 12623
rect 14393 12574 14431 12577
rect 14483 12574 14642 12577
rect 14694 12574 14853 12577
rect 14905 12574 18435 12577
rect 18487 12574 18645 12626
rect 18697 12574 18856 12626
rect 18908 12574 19068 12626
rect 19120 12574 19279 12626
rect 19331 12574 19489 12626
rect 19541 12574 19579 12626
rect 14393 12540 19579 12574
rect 19904 12626 20456 12660
rect 19904 12574 19943 12626
rect 19995 12623 20154 12626
rect 20206 12623 20365 12626
rect 20417 12623 20456 12626
rect 21875 12626 23974 12667
rect 21875 12623 21913 12626
rect 21965 12623 22124 12626
rect 22176 12623 22335 12626
rect 22387 12623 22545 12626
rect 22597 12623 22756 12626
rect 22808 12623 22968 12626
rect 23020 12623 23179 12626
rect 23231 12623 23389 12626
rect 19995 12577 20064 12623
rect 20110 12577 20154 12623
rect 20214 12577 20271 12623
rect 20317 12577 20365 12623
rect 20420 12577 20477 12623
rect 20523 12577 20580 12623
rect 20626 12577 20683 12623
rect 20729 12577 20786 12623
rect 20832 12577 20889 12623
rect 20935 12577 20992 12623
rect 21038 12577 21051 12623
rect 21386 12577 21399 12623
rect 23373 12577 23389 12623
rect 19995 12574 20154 12577
rect 20206 12574 20365 12577
rect 20417 12574 20456 12577
rect 19904 12540 20456 12574
rect 14393 12533 14943 12540
rect 12959 12482 13121 12493
rect 9334 12399 9463 12428
rect 9843 12410 9959 12447
rect 12959 12436 12970 12482
rect 13110 12436 13121 12482
rect 12959 12429 13121 12436
rect 9324 12353 9337 12399
rect 9383 12388 9459 12399
rect 9424 12353 9459 12388
rect 9505 12353 9582 12399
rect 9628 12353 9705 12399
rect 9751 12353 9764 12399
rect 9843 12364 9878 12410
rect 9924 12364 9959 12410
rect 9334 12336 9372 12353
rect 9424 12336 9463 12353
rect 9334 12309 9463 12336
rect 9334 12296 9462 12309
rect 9520 12173 9682 12213
rect 9520 12121 9591 12173
rect 9643 12121 9682 12173
rect 8605 12042 8618 12088
rect 8664 12042 8741 12088
rect 8787 12042 8864 12088
rect 8910 12042 8923 12088
rect 9089 12042 9238 12088
rect 9284 12042 9327 12088
rect 8611 12010 8920 12042
rect 9089 12010 9205 12042
rect 7450 11898 7758 11903
rect 6035 11864 6550 11898
rect 7036 11864 7758 11898
rect 8255 11878 8323 12000
rect 9520 11990 9682 12121
rect 9406 11987 9682 11990
rect 9406 11979 9591 11987
rect 9406 11933 9441 11979
rect 9487 11935 9591 11979
rect 9643 11966 9682 11987
rect 9843 11966 9959 12364
rect 10315 12388 13121 12429
rect 15181 12459 18143 12540
rect 18397 12533 19579 12540
rect 19905 12533 20456 12540
rect 21875 12574 21913 12577
rect 21965 12574 22124 12577
rect 22176 12574 22335 12577
rect 22387 12574 22545 12577
rect 22597 12574 22756 12577
rect 22808 12574 22968 12577
rect 23020 12574 23179 12577
rect 23231 12574 23389 12577
rect 23441 12574 23600 12626
rect 23652 12574 23811 12626
rect 23863 12574 23974 12626
rect 21875 12533 23974 12574
rect 15181 12413 15216 12459
rect 15262 12413 15374 12459
rect 15420 12413 15532 12459
rect 15578 12413 15690 12459
rect 15736 12413 15848 12459
rect 15894 12413 16006 12459
rect 16052 12413 16165 12459
rect 16211 12413 16323 12459
rect 16369 12413 16481 12459
rect 16527 12413 16639 12459
rect 16685 12413 16797 12459
rect 16843 12413 16955 12459
rect 17001 12413 17113 12459
rect 17159 12413 17272 12459
rect 17318 12413 17430 12459
rect 17476 12413 17588 12459
rect 17634 12413 17746 12459
rect 17792 12413 17904 12459
rect 17950 12413 18062 12459
rect 18108 12413 18143 12459
rect 23682 12499 23974 12533
rect 23682 12453 23820 12499
rect 23866 12453 23974 12499
rect 10315 12336 11532 12388
rect 11584 12336 13121 12388
rect 10315 12295 13121 12336
rect 14202 12353 14409 12399
rect 14455 12353 14522 12399
rect 14568 12353 14635 12399
rect 14681 12353 14748 12399
rect 14794 12353 14861 12399
rect 14907 12353 14920 12399
rect 15181 12377 18143 12413
rect 20632 12402 20940 12443
rect 20632 12399 20670 12402
rect 20722 12399 20850 12402
rect 20902 12399 20940 12402
rect 21186 12427 21254 12438
rect 13938 12287 14106 12298
rect 13938 12241 13955 12287
rect 14095 12241 14106 12287
rect 13938 12197 14106 12241
rect 11826 12157 14106 12197
rect 11826 12105 12665 12157
rect 12717 12105 14106 12157
rect 11826 12064 14106 12105
rect 14202 11966 14318 12353
rect 18502 12327 19474 12367
rect 20051 12353 20064 12399
rect 20110 12353 20168 12399
rect 20214 12353 20271 12399
rect 20317 12353 20374 12399
rect 20420 12353 20477 12399
rect 20523 12353 20580 12399
rect 20626 12353 20670 12399
rect 20729 12353 20786 12399
rect 20832 12353 20850 12399
rect 20935 12353 20992 12399
rect 21038 12353 21051 12399
rect 18502 12312 18540 12327
rect 18592 12312 18751 12327
rect 18803 12312 18962 12327
rect 19014 12312 19173 12327
rect 19225 12312 19384 12327
rect 19436 12312 19474 12327
rect 18362 12266 18375 12312
rect 18421 12266 18478 12312
rect 18524 12275 18540 12312
rect 18524 12266 18581 12275
rect 18627 12266 18684 12312
rect 18730 12275 18751 12312
rect 18730 12266 18787 12275
rect 18833 12266 18890 12312
rect 18936 12275 18962 12312
rect 18936 12266 18993 12275
rect 19039 12266 19096 12312
rect 19142 12275 19173 12312
rect 19142 12266 19199 12275
rect 19449 12266 19474 12312
rect 20632 12350 20670 12353
rect 20722 12350 20850 12353
rect 20902 12350 20940 12353
rect 20632 12310 20940 12350
rect 18154 12220 18284 12261
rect 18502 12235 19474 12266
rect 14498 12175 14838 12204
rect 14396 12129 14409 12175
rect 14455 12129 14522 12175
rect 14568 12164 14635 12175
rect 14588 12129 14635 12164
rect 14681 12129 14748 12175
rect 14794 12164 14861 12175
rect 14800 12129 14861 12164
rect 14907 12129 14920 12175
rect 18154 12168 18193 12220
rect 18245 12168 18284 12220
rect 18154 12165 18284 12168
rect 14498 12112 14536 12129
rect 14588 12112 14748 12129
rect 14800 12112 14838 12129
rect 14498 12071 14838 12112
rect 14997 12056 17976 12089
rect 14997 12010 15061 12056
rect 15201 12048 17976 12056
rect 15201 12010 15950 12048
rect 14997 11996 15950 12010
rect 16002 11996 17976 12048
rect 9643 11951 14515 11966
rect 14997 11955 17976 11996
rect 18154 12025 18219 12165
rect 18265 12025 18284 12165
rect 19859 12175 20409 12204
rect 19859 12164 20064 12175
rect 20110 12164 20168 12175
rect 19417 12088 19757 12129
rect 18362 12042 18375 12088
rect 18421 12042 18478 12088
rect 18524 12042 18581 12088
rect 18627 12042 18684 12088
rect 18730 12042 18787 12088
rect 18833 12042 18890 12088
rect 18936 12042 18993 12088
rect 19039 12042 19096 12088
rect 19142 12042 19199 12088
rect 19449 12042 19757 12088
rect 19859 12112 19897 12164
rect 19949 12129 20064 12164
rect 20160 12129 20168 12164
rect 20214 12129 20271 12175
rect 20317 12164 20374 12175
rect 20317 12129 20319 12164
rect 19949 12112 20108 12129
rect 20160 12112 20319 12129
rect 20371 12129 20374 12164
rect 20420 12129 20477 12175
rect 20523 12129 20580 12175
rect 20626 12129 20683 12175
rect 20729 12129 20786 12175
rect 20832 12129 20889 12175
rect 20935 12129 20992 12175
rect 21038 12129 21051 12175
rect 20371 12112 20409 12129
rect 19859 12071 20409 12112
rect 18154 12002 18284 12025
rect 19417 12010 19757 12042
rect 9643 11935 14409 11951
rect 9487 11933 14409 11935
rect 9406 11930 14409 11933
rect 9406 11884 13336 11930
rect 13382 11884 13503 11930
rect 13549 11884 13668 11930
rect 13714 11884 13833 11930
rect 13879 11905 14409 11930
rect 14455 11905 14522 11951
rect 14568 11905 14635 11951
rect 14681 11905 14748 11951
rect 14794 11905 14861 11951
rect 14907 11905 14920 11951
rect 18154 11950 18193 12002
rect 18245 11950 18284 12002
rect 18154 11910 18284 11950
rect 19641 11953 19757 12010
rect 21186 12005 21197 12427
rect 21243 12005 21254 12427
rect 21394 12399 21702 12436
rect 21386 12353 21399 12399
rect 23373 12353 23386 12399
rect 21394 12343 21432 12353
rect 21484 12343 21612 12353
rect 21664 12343 21702 12353
rect 21394 12303 21702 12343
rect 23682 12335 23974 12453
rect 23682 12289 23820 12335
rect 23866 12289 23974 12335
rect 23682 12197 23974 12289
rect 23182 12175 23974 12197
rect 21386 12129 21399 12175
rect 23373 12129 23974 12175
rect 23182 12078 23974 12129
rect 21186 11953 21254 12005
rect 19641 11916 21254 11953
rect 21394 11951 21702 11973
rect 13879 11884 14515 11905
rect 8255 11864 9320 11878
rect 345 11800 452 11846
rect 498 11800 637 11846
rect 3081 11833 4240 11862
rect 4857 11818 4870 11864
rect 5120 11818 5140 11864
rect 5223 11818 5280 11864
rect 5326 11818 5351 11864
rect 5429 11818 5486 11864
rect 5532 11818 5562 11864
rect 5635 11818 5692 11864
rect 5738 11818 5773 11864
rect 5841 11818 5898 11864
rect 5944 11818 5957 11864
rect 6035 11818 6451 11864
rect 6497 11818 6568 11864
rect 6614 11818 6685 11864
rect 6731 11818 6803 11864
rect 6849 11818 6921 11864
rect 6967 11818 7039 11864
rect 7085 11862 7506 11864
rect 7085 11818 7488 11862
rect 7552 11818 7623 11864
rect 7669 11862 7740 11864
rect 7720 11818 7740 11862
rect 7786 11818 7858 11864
rect 7904 11818 7976 11864
rect 8022 11818 8094 11864
rect 8140 11818 8153 11864
rect 8255 11818 8618 11864
rect 8664 11818 8741 11864
rect 8787 11818 8864 11864
rect 8910 11818 9238 11864
rect 9284 11818 9327 11864
rect 9406 11846 14515 11884
rect 18502 11864 19474 11904
rect 18362 11818 18375 11864
rect 18421 11818 18478 11864
rect 18524 11818 18540 11864
rect 18627 11818 18684 11864
rect 18730 11818 18751 11864
rect 18833 11818 18890 11864
rect 18936 11818 18962 11864
rect 19039 11818 19096 11864
rect 19142 11818 19173 11864
rect 19449 11818 19474 11864
rect 19641 11870 20113 11916
rect 20159 11870 20300 11916
rect 20346 11870 20487 11916
rect 20533 11870 20673 11916
rect 20719 11870 20860 11916
rect 20906 11870 21254 11916
rect 21386 11905 21399 11951
rect 23373 11905 23386 11951
rect 19641 11860 21254 11870
rect 20078 11833 21254 11860
rect 21394 11880 21432 11905
rect 21484 11880 21612 11905
rect 21664 11880 21702 11905
rect 21394 11840 21702 11880
rect 23682 11846 23974 12078
rect 345 11767 637 11800
rect 4891 11812 4929 11818
rect 4981 11812 5140 11818
rect 5192 11812 5351 11818
rect 5403 11812 5562 11818
rect 5614 11812 5773 11818
rect 5825 11812 5863 11818
rect 4467 11767 4622 11774
rect 4891 11772 5863 11812
rect 6035 11778 6550 11818
rect 7036 11810 7488 11818
rect 7540 11810 7668 11818
rect 7720 11810 7758 11818
rect 7036 11778 7758 11810
rect 7450 11770 7758 11778
rect 345 11726 2439 11767
rect 345 11674 451 11726
rect 503 11674 662 11726
rect 714 11674 873 11726
rect 925 11674 1083 11726
rect 1135 11674 1294 11726
rect 1346 11674 1506 11726
rect 1558 11674 1717 11726
rect 1769 11674 1927 11726
rect 1979 11674 2138 11726
rect 2190 11674 2349 11726
rect 2401 11674 2439 11726
rect 345 11633 2439 11674
rect 4314 11726 4622 11767
rect 8255 11758 9320 11818
rect 18502 11812 18540 11818
rect 18592 11812 18751 11818
rect 18803 11812 18962 11818
rect 19014 11812 19173 11818
rect 19225 11812 19384 11818
rect 19436 11812 19474 11818
rect 18502 11772 19474 11812
rect 23682 11800 23820 11846
rect 23866 11800 23974 11846
rect 19696 11767 19852 11774
rect 23682 11767 23974 11800
rect 4314 11674 4352 11726
rect 4404 11723 4532 11726
rect 4404 11677 4513 11723
rect 4404 11674 4532 11677
rect 4584 11674 4622 11726
rect 4314 11633 4622 11674
rect 19696 11726 20005 11767
rect 19696 11674 19735 11726
rect 19787 11723 19915 11726
rect 19803 11677 19915 11723
rect 19787 11674 19915 11677
rect 19967 11674 20005 11726
rect 345 11600 637 11633
rect 4467 11626 4622 11633
rect 345 11554 452 11600
rect 498 11554 637 11600
rect 4891 11588 5863 11628
rect 7450 11622 7758 11630
rect 4891 11582 4929 11588
rect 4981 11582 5140 11588
rect 5192 11582 5351 11588
rect 5403 11582 5562 11588
rect 5614 11582 5773 11588
rect 5825 11582 5863 11588
rect 6035 11582 6550 11622
rect 7036 11590 7758 11622
rect 7036 11582 7488 11590
rect 7540 11582 7668 11590
rect 7720 11582 7758 11590
rect 8255 11582 9320 11642
rect 19696 11633 20005 11674
rect 21875 11726 23974 11767
rect 21875 11674 21913 11726
rect 21965 11674 22124 11726
rect 22176 11674 22335 11726
rect 22387 11674 22545 11726
rect 22597 11674 22756 11726
rect 22808 11674 22968 11726
rect 23020 11674 23179 11726
rect 23231 11674 23389 11726
rect 23441 11674 23600 11726
rect 23652 11674 23811 11726
rect 23863 11674 23974 11726
rect 21875 11633 23974 11674
rect 18502 11588 19474 11628
rect 19696 11626 19852 11633
rect 18502 11582 18540 11588
rect 18592 11582 18751 11588
rect 18803 11582 18962 11588
rect 19014 11582 19173 11588
rect 19225 11582 19384 11588
rect 19436 11582 19474 11588
rect 345 11437 637 11554
rect 3081 11538 4240 11567
rect 2616 11498 2924 11538
rect 2616 11495 2654 11498
rect 2706 11495 2834 11498
rect 2886 11495 2924 11498
rect 3081 11530 4679 11538
rect 4857 11536 4870 11582
rect 5120 11536 5140 11582
rect 5223 11536 5280 11582
rect 5326 11536 5351 11582
rect 5429 11536 5486 11582
rect 5532 11536 5562 11582
rect 5635 11536 5692 11582
rect 5738 11536 5773 11582
rect 5841 11536 5898 11582
rect 5944 11536 5957 11582
rect 6035 11536 6451 11582
rect 6497 11536 6568 11582
rect 6614 11536 6685 11582
rect 6731 11536 6803 11582
rect 6849 11536 6921 11582
rect 6967 11536 7039 11582
rect 7085 11538 7488 11582
rect 7085 11536 7506 11538
rect 7552 11536 7623 11582
rect 7720 11538 7740 11582
rect 7669 11536 7740 11538
rect 7786 11536 7858 11582
rect 7904 11536 7976 11582
rect 8022 11536 8094 11582
rect 8140 11536 8153 11582
rect 8255 11536 8618 11582
rect 8664 11536 8741 11582
rect 8787 11536 8864 11582
rect 8910 11536 9238 11582
rect 9284 11536 9327 11582
rect 933 11449 946 11495
rect 2920 11449 2933 11495
rect 3081 11484 3413 11530
rect 3459 11484 3599 11530
rect 3645 11484 3786 11530
rect 3832 11484 3973 11530
rect 4019 11484 4159 11530
rect 4205 11484 4679 11530
rect 4891 11496 5863 11536
rect 6035 11502 6550 11536
rect 7036 11502 7758 11536
rect 345 11391 452 11437
rect 498 11391 637 11437
rect 2616 11446 2654 11449
rect 2706 11446 2834 11449
rect 2886 11446 2924 11449
rect 2616 11405 2924 11446
rect 3081 11447 4679 11484
rect 345 11322 637 11391
rect 3081 11365 3149 11447
rect 345 11274 1090 11322
rect 345 11228 452 11274
rect 498 11271 1090 11274
rect 498 11228 946 11271
rect 345 11225 946 11228
rect 2920 11225 2933 11271
rect 345 11203 1090 11225
rect 345 11111 637 11203
rect 345 11065 452 11111
rect 498 11065 637 11111
rect 345 10947 637 11065
rect 2616 11050 2924 11090
rect 2616 11047 2654 11050
rect 2706 11047 2834 11050
rect 2886 11047 2924 11050
rect 933 11001 946 11047
rect 2920 11001 2933 11047
rect 2616 10998 2654 11001
rect 2706 10998 2834 11001
rect 2886 10998 2924 11001
rect 2616 10957 2924 10998
rect 345 10901 452 10947
rect 498 10901 637 10947
rect 3081 10943 3092 11365
rect 3138 10943 3149 11365
rect 4561 11390 4679 11447
rect 6035 11402 6151 11502
rect 7450 11497 7758 11502
rect 8255 11522 9320 11536
rect 4561 11358 5957 11390
rect 3825 11288 4315 11329
rect 3825 11271 3864 11288
rect 3916 11271 4044 11288
rect 4096 11271 4224 11288
rect 3268 11225 3281 11271
rect 3327 11225 3384 11271
rect 3430 11225 3487 11271
rect 3533 11225 3590 11271
rect 3636 11225 3693 11271
rect 3739 11225 3796 11271
rect 3842 11236 3864 11271
rect 3842 11225 3899 11236
rect 3945 11225 4002 11271
rect 4096 11236 4105 11271
rect 4048 11225 4105 11236
rect 4151 11225 4209 11271
rect 4276 11236 4315 11288
rect 4561 11312 4870 11358
rect 5120 11312 5177 11358
rect 5223 11312 5280 11358
rect 5326 11312 5383 11358
rect 5429 11312 5486 11358
rect 5532 11312 5589 11358
rect 5635 11312 5692 11358
rect 5738 11312 5795 11358
rect 5841 11312 5898 11358
rect 5944 11312 5957 11358
rect 4561 11268 5957 11312
rect 4255 11225 4315 11236
rect 3825 11196 4315 11225
rect 6035 11262 6072 11402
rect 6118 11262 6151 11402
rect 4891 11134 5863 11168
rect 6035 11159 6151 11262
rect 6237 11402 6370 11422
rect 6237 11363 6294 11402
rect 6237 11311 6275 11363
rect 6237 11262 6294 11311
rect 6340 11262 6370 11402
rect 8255 11400 8323 11522
rect 9406 11516 14515 11554
rect 18362 11536 18375 11582
rect 18421 11536 18478 11582
rect 18524 11536 18540 11582
rect 18627 11536 18684 11582
rect 18730 11536 18751 11582
rect 18833 11536 18890 11582
rect 18936 11536 18962 11582
rect 19039 11536 19096 11582
rect 19142 11536 19173 11582
rect 19449 11536 19474 11582
rect 23682 11600 23974 11633
rect 20078 11540 21254 11567
rect 9406 11470 13336 11516
rect 13382 11470 13503 11516
rect 13549 11470 13668 11516
rect 13714 11470 13833 11516
rect 13879 11495 14515 11516
rect 18502 11496 19474 11536
rect 19641 11530 21254 11540
rect 13879 11470 14409 11495
rect 9406 11467 14409 11470
rect 9406 11421 9441 11467
rect 9487 11465 14409 11467
rect 9487 11421 9591 11465
rect 9406 11413 9591 11421
rect 9643 11449 14409 11465
rect 14455 11449 14522 11495
rect 14568 11449 14635 11495
rect 14681 11449 14748 11495
rect 14794 11449 14861 11495
rect 14907 11449 14920 11495
rect 18154 11450 18284 11490
rect 9643 11434 14515 11449
rect 9643 11413 9682 11434
rect 9406 11410 9682 11413
rect 6521 11390 7282 11397
rect 6520 11358 7528 11390
rect 6438 11312 6451 11358
rect 6497 11356 6568 11358
rect 6497 11312 6558 11356
rect 6614 11312 6685 11358
rect 6731 11356 6803 11358
rect 6731 11312 6769 11356
rect 6849 11312 6921 11358
rect 6967 11356 7039 11358
rect 6967 11312 6981 11356
rect 6520 11304 6558 11312
rect 6610 11304 6769 11312
rect 6821 11304 6981 11312
rect 7033 11312 7039 11356
rect 7085 11356 7506 11358
rect 7085 11312 7192 11356
rect 7033 11304 7192 11312
rect 7244 11312 7506 11356
rect 7552 11312 7623 11358
rect 7669 11312 7740 11358
rect 7786 11312 7858 11358
rect 7904 11312 7976 11358
rect 8022 11312 8094 11358
rect 8140 11312 8153 11358
rect 7244 11304 7528 11312
rect 6520 11271 7528 11304
rect 6520 11270 7282 11271
rect 6521 11264 7282 11270
rect 6237 11239 6370 11262
rect 8255 11260 8266 11400
rect 8312 11260 8323 11400
rect 8611 11358 8920 11390
rect 9089 11358 9205 11390
rect 8605 11312 8618 11358
rect 8664 11312 8741 11358
rect 8787 11312 8864 11358
rect 8910 11312 8923 11358
rect 9089 11312 9238 11358
rect 9284 11312 9327 11358
rect 8255 11249 8323 11260
rect 6035 11134 6550 11159
rect 7036 11156 7528 11159
rect 7036 11134 7758 11156
rect 4857 11088 4870 11134
rect 5120 11128 5177 11134
rect 5120 11088 5140 11128
rect 5223 11088 5280 11134
rect 5326 11128 5383 11134
rect 5326 11088 5351 11128
rect 5429 11088 5486 11134
rect 5532 11128 5589 11134
rect 5532 11088 5562 11128
rect 5635 11088 5692 11134
rect 5738 11128 5795 11134
rect 5738 11088 5773 11128
rect 5841 11088 5898 11134
rect 5944 11088 5957 11134
rect 6035 11088 6451 11134
rect 6497 11088 6568 11134
rect 6614 11088 6685 11134
rect 6731 11088 6803 11134
rect 6849 11088 6921 11134
rect 6967 11088 7039 11134
rect 7085 11116 7506 11134
rect 7085 11088 7488 11116
rect 7552 11088 7623 11134
rect 7669 11116 7740 11134
rect 7720 11088 7740 11116
rect 7786 11088 7858 11134
rect 7904 11088 7976 11134
rect 8022 11088 8094 11134
rect 8140 11088 8153 11134
rect 3378 11047 3686 11082
rect 4891 11076 4929 11088
rect 4981 11076 5140 11088
rect 5192 11076 5351 11088
rect 5403 11076 5562 11088
rect 5614 11076 5773 11088
rect 5825 11076 5863 11088
rect 3268 11001 3281 11047
rect 3327 11001 3384 11047
rect 3430 11042 3487 11047
rect 3468 11001 3487 11042
rect 3533 11001 3590 11047
rect 3636 11042 3693 11047
rect 3648 11001 3693 11042
rect 3739 11001 3796 11047
rect 3842 11001 3899 11047
rect 3945 11001 4002 11047
rect 4048 11001 4105 11047
rect 4151 11001 4209 11047
rect 4255 11001 4268 11047
rect 4891 11036 5863 11076
rect 6035 11039 6550 11088
rect 7036 11064 7488 11088
rect 7540 11064 7668 11088
rect 7720 11064 7758 11088
rect 7036 11039 7758 11064
rect 7450 11023 7758 11039
rect 3378 10990 3416 11001
rect 3468 10990 3596 11001
rect 3648 10990 3686 11001
rect 3378 10949 3686 10990
rect 3081 10932 3149 10943
rect 345 10867 637 10901
rect 345 10826 2439 10867
rect 3844 10860 4605 10867
rect 345 10774 451 10826
rect 503 10774 662 10826
rect 714 10774 873 10826
rect 925 10823 1083 10826
rect 1135 10823 1294 10826
rect 1346 10823 1506 10826
rect 1558 10823 1717 10826
rect 1769 10823 1927 10826
rect 1979 10823 2138 10826
rect 2190 10823 2349 10826
rect 2401 10823 2439 10826
rect 3843 10826 4605 10860
rect 3843 10823 3881 10826
rect 3933 10823 4092 10826
rect 4144 10823 4304 10826
rect 925 10777 946 10823
rect 2920 10777 2933 10823
rect 3268 10777 3281 10823
rect 3327 10777 3384 10823
rect 3430 10777 3487 10823
rect 3533 10777 3590 10823
rect 3636 10777 3693 10823
rect 3739 10777 3796 10823
rect 3842 10777 3881 10823
rect 3945 10777 4002 10823
rect 4048 10777 4092 10823
rect 4151 10777 4209 10823
rect 4255 10777 4304 10823
rect 925 10774 1083 10777
rect 1135 10774 1294 10777
rect 1346 10774 1506 10777
rect 1558 10774 1717 10777
rect 1769 10774 1927 10777
rect 1979 10774 2138 10777
rect 2190 10774 2349 10777
rect 2401 10774 2439 10777
rect 345 10733 2439 10774
rect 3843 10774 3881 10777
rect 3933 10774 4092 10777
rect 4144 10774 4304 10777
rect 4356 10774 4515 10826
rect 4567 10774 4605 10826
rect 3843 10740 4605 10774
rect 3844 10733 4605 10740
rect 4779 10860 5961 10867
rect 4779 10826 6555 10860
rect 4779 10774 4817 10826
rect 4869 10774 5027 10826
rect 5079 10774 5238 10826
rect 5290 10774 5450 10826
rect 5502 10774 5661 10826
rect 5713 10774 5871 10826
rect 5923 10823 6555 10826
rect 5923 10777 6086 10823
rect 6320 10777 6555 10823
rect 5923 10774 6555 10777
rect 4779 10740 6555 10774
rect 7543 10826 8439 10867
rect 7543 10823 7927 10826
rect 7979 10823 8138 10826
rect 7543 10777 7554 10823
rect 8070 10777 8138 10823
rect 7543 10774 7927 10777
rect 7979 10774 8138 10777
rect 8190 10774 8349 10826
rect 8401 10774 8439 10826
rect 4779 10733 5961 10740
rect 7543 10733 8439 10774
rect 8611 10826 8920 11312
rect 8611 10774 8649 10826
rect 8701 10823 8829 10826
rect 8705 10777 8817 10823
rect 8701 10774 8829 10777
rect 8881 10774 8920 10826
rect 345 10699 637 10733
rect 345 10653 452 10699
rect 498 10653 637 10699
rect 345 10535 637 10653
rect 3081 10657 3149 10668
rect 2616 10602 2924 10643
rect 2616 10599 2654 10602
rect 2706 10599 2834 10602
rect 2886 10599 2924 10602
rect 933 10553 946 10599
rect 2920 10553 2933 10599
rect 345 10489 452 10535
rect 498 10489 637 10535
rect 2616 10550 2654 10553
rect 2706 10550 2834 10553
rect 2886 10550 2924 10553
rect 2616 10510 2924 10550
rect 345 10397 637 10489
rect 345 10375 1090 10397
rect 345 10372 946 10375
rect 345 10326 452 10372
rect 498 10329 946 10372
rect 2920 10329 2933 10375
rect 498 10326 1090 10329
rect 345 10278 1090 10326
rect 345 10209 637 10278
rect 345 10163 452 10209
rect 498 10163 637 10209
rect 3081 10235 3092 10657
rect 3138 10235 3149 10657
rect 3378 10610 3686 10651
rect 3378 10599 3416 10610
rect 3468 10599 3596 10610
rect 3648 10599 3686 10610
rect 3268 10553 3281 10599
rect 3327 10553 3384 10599
rect 3468 10558 3487 10599
rect 3430 10553 3487 10558
rect 3533 10553 3590 10599
rect 3648 10558 3693 10599
rect 3636 10553 3693 10558
rect 3739 10553 3796 10599
rect 3842 10553 3899 10599
rect 3945 10553 4002 10599
rect 4048 10553 4105 10599
rect 4151 10553 4209 10599
rect 4255 10553 4268 10599
rect 3378 10518 3686 10553
rect 4891 10524 5863 10564
rect 7450 10561 7758 10577
rect 4891 10512 4929 10524
rect 4981 10512 5140 10524
rect 5192 10512 5351 10524
rect 5403 10512 5562 10524
rect 5614 10512 5773 10524
rect 5825 10512 5863 10524
rect 6035 10512 6550 10561
rect 7036 10536 7758 10561
rect 7036 10512 7488 10536
rect 7540 10512 7668 10536
rect 7720 10512 7758 10536
rect 4857 10466 4870 10512
rect 5120 10472 5140 10512
rect 5120 10466 5177 10472
rect 5223 10466 5280 10512
rect 5326 10472 5351 10512
rect 5326 10466 5383 10472
rect 5429 10466 5486 10512
rect 5532 10472 5562 10512
rect 5532 10466 5589 10472
rect 5635 10466 5692 10512
rect 5738 10472 5773 10512
rect 5738 10466 5795 10472
rect 5841 10466 5898 10512
rect 5944 10466 5957 10512
rect 6035 10466 6451 10512
rect 6497 10466 6568 10512
rect 6614 10466 6685 10512
rect 6731 10466 6803 10512
rect 6849 10466 6921 10512
rect 6967 10466 7039 10512
rect 7085 10484 7488 10512
rect 7085 10466 7506 10484
rect 7552 10466 7623 10512
rect 7720 10484 7740 10512
rect 7669 10466 7740 10484
rect 7786 10466 7858 10512
rect 7904 10466 7976 10512
rect 8022 10466 8094 10512
rect 8140 10466 8153 10512
rect 4891 10432 5863 10466
rect 6035 10441 6550 10466
rect 7036 10444 7758 10466
rect 7036 10441 7528 10444
rect 3825 10375 4315 10404
rect 3268 10329 3281 10375
rect 3327 10329 3384 10375
rect 3430 10329 3487 10375
rect 3533 10329 3590 10375
rect 3636 10329 3693 10375
rect 3739 10329 3796 10375
rect 3842 10364 3899 10375
rect 3842 10329 3864 10364
rect 3945 10329 4002 10375
rect 4048 10364 4105 10375
rect 4096 10329 4105 10364
rect 4151 10329 4209 10375
rect 4255 10364 4315 10375
rect 3825 10312 3864 10329
rect 3916 10312 4044 10329
rect 4096 10312 4224 10329
rect 4276 10312 4315 10364
rect 6035 10338 6151 10441
rect 3825 10271 4315 10312
rect 4561 10288 5957 10332
rect 345 10046 637 10163
rect 2616 10154 2924 10195
rect 2616 10151 2654 10154
rect 2706 10151 2834 10154
rect 2886 10151 2924 10154
rect 3081 10153 3149 10235
rect 4561 10242 4870 10288
rect 5120 10242 5177 10288
rect 5223 10242 5280 10288
rect 5326 10242 5383 10288
rect 5429 10242 5486 10288
rect 5532 10242 5589 10288
rect 5635 10242 5692 10288
rect 5738 10242 5795 10288
rect 5841 10242 5898 10288
rect 5944 10242 5957 10288
rect 4561 10210 5957 10242
rect 4561 10153 4679 10210
rect 933 10105 946 10151
rect 2920 10105 2933 10151
rect 3081 10116 4679 10153
rect 2616 10102 2654 10105
rect 2706 10102 2834 10105
rect 2886 10102 2924 10105
rect 2616 10062 2924 10102
rect 3081 10070 3413 10116
rect 3459 10070 3599 10116
rect 3645 10070 3786 10116
rect 3832 10070 3973 10116
rect 4019 10070 4159 10116
rect 4205 10070 4679 10116
rect 6035 10198 6072 10338
rect 6118 10198 6151 10338
rect 3081 10062 4679 10070
rect 4891 10064 5863 10104
rect 6035 10098 6151 10198
rect 6237 10338 6370 10361
rect 6237 10289 6294 10338
rect 6237 10237 6275 10289
rect 6237 10198 6294 10237
rect 6340 10198 6370 10338
rect 8255 10340 8323 10351
rect 6521 10330 7282 10336
rect 6520 10329 7282 10330
rect 6520 10296 7528 10329
rect 6520 10288 6558 10296
rect 6610 10288 6769 10296
rect 6821 10288 6981 10296
rect 6438 10242 6451 10288
rect 6497 10244 6558 10288
rect 6497 10242 6568 10244
rect 6614 10242 6685 10288
rect 6731 10244 6769 10288
rect 6731 10242 6803 10244
rect 6849 10242 6921 10288
rect 6967 10244 6981 10288
rect 7033 10288 7192 10296
rect 7033 10244 7039 10288
rect 6967 10242 7039 10244
rect 7085 10244 7192 10288
rect 7244 10288 7528 10296
rect 7244 10244 7506 10288
rect 7085 10242 7506 10244
rect 7552 10242 7623 10288
rect 7669 10242 7740 10288
rect 7786 10242 7858 10288
rect 7904 10242 7976 10288
rect 8022 10242 8094 10288
rect 8140 10242 8153 10288
rect 6520 10210 7528 10242
rect 6521 10203 7282 10210
rect 6237 10178 6370 10198
rect 8255 10200 8266 10340
rect 8312 10200 8323 10340
rect 8611 10288 8920 10774
rect 9089 10860 9205 11312
rect 9520 11279 9682 11410
rect 9520 11227 9591 11279
rect 9643 11227 9682 11279
rect 9520 11187 9682 11227
rect 9334 11091 9462 11104
rect 9334 11064 9463 11091
rect 9334 11047 9372 11064
rect 9424 11047 9463 11064
rect 9324 11001 9337 11047
rect 9424 11012 9459 11047
rect 9383 11001 9459 11012
rect 9505 11001 9582 11047
rect 9628 11001 9705 11047
rect 9751 11001 9764 11047
rect 9843 11036 9959 11434
rect 11826 11295 14106 11336
rect 11826 11243 12665 11295
rect 12717 11243 14106 11295
rect 11826 11203 14106 11243
rect 13938 11159 14106 11203
rect 13938 11113 13955 11159
rect 14095 11113 14106 11159
rect 9334 10972 9463 11001
rect 9843 10990 9878 11036
rect 9924 10990 9959 11036
rect 9843 10953 9959 10990
rect 10315 11064 13121 11105
rect 13938 11102 14106 11113
rect 10315 11012 11532 11064
rect 11584 11012 13121 11064
rect 10315 10971 13121 11012
rect 14202 11047 14318 11434
rect 14997 11404 17976 11445
rect 14997 11390 16328 11404
rect 14997 11344 15061 11390
rect 15201 11352 16328 11390
rect 16380 11352 17976 11404
rect 15201 11344 17976 11352
rect 14498 11288 14838 11329
rect 14997 11311 17976 11344
rect 18154 11398 18193 11450
rect 18245 11398 18284 11450
rect 18154 11375 18284 11398
rect 19641 11484 20113 11530
rect 20159 11484 20300 11530
rect 20346 11484 20487 11530
rect 20533 11484 20673 11530
rect 20719 11484 20860 11530
rect 20906 11484 21254 11530
rect 21394 11520 21702 11560
rect 21394 11495 21432 11520
rect 21484 11495 21612 11520
rect 21664 11495 21702 11520
rect 23682 11554 23820 11600
rect 23866 11554 23974 11600
rect 19641 11447 21254 11484
rect 21386 11449 21399 11495
rect 23373 11449 23386 11495
rect 19641 11390 19757 11447
rect 14498 11271 14536 11288
rect 14588 11271 14748 11288
rect 14800 11271 14838 11288
rect 14396 11225 14409 11271
rect 14455 11225 14522 11271
rect 14588 11236 14635 11271
rect 14568 11225 14635 11236
rect 14681 11225 14748 11271
rect 14800 11236 14861 11271
rect 14794 11225 14861 11236
rect 14907 11225 14920 11271
rect 18154 11235 18219 11375
rect 18265 11235 18284 11375
rect 19417 11358 19757 11390
rect 18362 11312 18375 11358
rect 18421 11312 18478 11358
rect 18524 11312 18581 11358
rect 18627 11312 18684 11358
rect 18730 11312 18787 11358
rect 18833 11312 18890 11358
rect 18936 11312 18993 11358
rect 19039 11312 19096 11358
rect 19142 11312 19199 11358
rect 19449 11312 19757 11358
rect 21186 11395 21254 11447
rect 21394 11427 21702 11449
rect 19417 11271 19757 11312
rect 19859 11288 20409 11329
rect 18154 11232 18284 11235
rect 14498 11196 14838 11225
rect 18154 11180 18193 11232
rect 18245 11180 18284 11232
rect 19859 11236 19897 11288
rect 19949 11271 20108 11288
rect 20160 11271 20319 11288
rect 19949 11236 20064 11271
rect 20160 11236 20168 11271
rect 19859 11225 20064 11236
rect 20110 11225 20168 11236
rect 20214 11225 20271 11271
rect 20317 11236 20319 11271
rect 20371 11271 20409 11288
rect 20371 11236 20374 11271
rect 20317 11225 20374 11236
rect 20420 11225 20477 11271
rect 20523 11225 20580 11271
rect 20626 11225 20683 11271
rect 20729 11225 20786 11271
rect 20832 11225 20889 11271
rect 20935 11225 20992 11271
rect 21038 11225 21051 11271
rect 19859 11196 20409 11225
rect 18154 11139 18284 11180
rect 18502 11134 19474 11165
rect 18362 11088 18375 11134
rect 18421 11088 18478 11134
rect 18524 11125 18581 11134
rect 18524 11088 18540 11125
rect 18627 11088 18684 11134
rect 18730 11125 18787 11134
rect 18730 11088 18751 11125
rect 18833 11088 18890 11134
rect 18936 11125 18993 11134
rect 18936 11088 18962 11125
rect 19039 11088 19096 11134
rect 19142 11125 19199 11134
rect 19142 11088 19173 11125
rect 19449 11088 19474 11134
rect 18502 11073 18540 11088
rect 18592 11073 18751 11088
rect 18803 11073 18962 11088
rect 19014 11073 19173 11088
rect 19225 11073 19384 11088
rect 19436 11073 19474 11088
rect 14202 11001 14409 11047
rect 14455 11001 14522 11047
rect 14568 11001 14635 11047
rect 14681 11001 14748 11047
rect 14794 11001 14861 11047
rect 14907 11001 14920 11047
rect 18502 11033 19474 11073
rect 20632 11050 20940 11090
rect 20632 11047 20670 11050
rect 20722 11047 20850 11050
rect 20902 11047 20940 11050
rect 12959 10964 13121 10971
rect 12959 10918 12970 10964
rect 13110 10918 13121 10964
rect 12959 10907 13121 10918
rect 15181 10987 18143 11023
rect 20051 11001 20064 11047
rect 20110 11001 20168 11047
rect 20214 11001 20271 11047
rect 20317 11001 20374 11047
rect 20420 11001 20477 11047
rect 20523 11001 20580 11047
rect 20626 11001 20670 11047
rect 20729 11001 20786 11047
rect 20832 11001 20850 11047
rect 20935 11001 20992 11047
rect 21038 11001 21051 11047
rect 15181 10941 15216 10987
rect 15262 10941 15374 10987
rect 15420 10941 15532 10987
rect 15578 10941 15690 10987
rect 15736 10941 15848 10987
rect 15894 10941 16006 10987
rect 16052 10941 16165 10987
rect 16211 10941 16323 10987
rect 16369 10941 16481 10987
rect 16527 10941 16639 10987
rect 16685 10941 16797 10987
rect 16843 10941 16955 10987
rect 17001 10941 17113 10987
rect 17159 10941 17272 10987
rect 17318 10941 17430 10987
rect 17476 10941 17588 10987
rect 17634 10941 17746 10987
rect 17792 10941 17904 10987
rect 17950 10941 18062 10987
rect 18108 10941 18143 10987
rect 20632 10998 20670 11001
rect 20722 10998 20850 11001
rect 20902 10998 20940 11001
rect 20632 10957 20940 10998
rect 21186 10973 21197 11395
rect 21243 10973 21254 11395
rect 23682 11322 23974 11554
rect 23182 11271 23974 11322
rect 21386 11225 21399 11271
rect 23373 11225 23974 11271
rect 23182 11203 23974 11225
rect 23682 11111 23974 11203
rect 21394 11057 21702 11097
rect 21394 11047 21432 11057
rect 21484 11047 21612 11057
rect 21664 11047 21702 11057
rect 23682 11065 23820 11111
rect 23866 11065 23974 11111
rect 21386 11001 21399 11047
rect 23373 11001 23386 11047
rect 21186 10962 21254 10973
rect 21394 10964 21702 11001
rect 9812 10860 10120 10867
rect 10385 10860 12583 10874
rect 13350 10860 14111 10867
rect 9089 10837 12583 10860
rect 13301 10837 14111 10860
rect 9089 10826 14111 10837
rect 9089 10823 9850 10826
rect 9089 10777 9337 10823
rect 9383 10777 9459 10823
rect 9505 10777 9582 10823
rect 9628 10777 9705 10823
rect 9751 10777 9850 10823
rect 9089 10774 9850 10777
rect 9902 10774 10030 10826
rect 10082 10823 13387 10826
rect 10082 10777 10433 10823
rect 10479 10777 10591 10823
rect 10637 10777 10749 10823
rect 10795 10777 10907 10823
rect 10953 10777 11066 10823
rect 11112 10777 11224 10823
rect 11270 10777 11382 10823
rect 11428 10777 11540 10823
rect 11586 10777 11698 10823
rect 11744 10777 11856 10823
rect 11902 10777 12015 10823
rect 12061 10777 12173 10823
rect 12219 10777 12331 10823
rect 12377 10777 12489 10823
rect 12535 10777 13336 10823
rect 13382 10777 13387 10823
rect 10082 10774 13387 10777
rect 13439 10823 13598 10826
rect 13439 10777 13503 10823
rect 13549 10777 13598 10823
rect 13439 10774 13598 10777
rect 13650 10823 13810 10826
rect 13862 10823 14021 10826
rect 13650 10777 13668 10823
rect 13714 10777 13810 10823
rect 13879 10777 14021 10823
rect 13650 10774 13810 10777
rect 13862 10774 14021 10777
rect 14073 10774 14111 10826
rect 9089 10763 14111 10774
rect 9089 10740 12583 10763
rect 13301 10740 14111 10763
rect 9089 10288 9205 10740
rect 9812 10733 10120 10740
rect 10385 10726 12583 10740
rect 13350 10733 14111 10740
rect 14393 10860 14943 10867
rect 15181 10860 18143 10941
rect 23682 10947 23974 11065
rect 23682 10901 23820 10947
rect 23866 10901 23974 10947
rect 23682 10867 23974 10901
rect 18397 10860 19579 10867
rect 19905 10860 20456 10867
rect 14393 10826 19579 10860
rect 14393 10823 14431 10826
rect 14483 10823 14642 10826
rect 14694 10823 14853 10826
rect 14905 10823 18435 10826
rect 14393 10777 14409 10823
rect 14483 10777 14522 10823
rect 14568 10777 14635 10823
rect 14694 10777 14748 10823
rect 14794 10777 14853 10823
rect 14907 10777 15216 10823
rect 15262 10777 15374 10823
rect 15420 10777 15532 10823
rect 15578 10777 15690 10823
rect 15736 10777 15848 10823
rect 15894 10777 16006 10823
rect 16052 10777 16165 10823
rect 16211 10777 16323 10823
rect 16369 10777 16481 10823
rect 16527 10777 16639 10823
rect 16685 10777 16797 10823
rect 16843 10777 16955 10823
rect 17001 10777 17113 10823
rect 17159 10777 17272 10823
rect 17318 10777 17430 10823
rect 17476 10777 17588 10823
rect 17634 10777 17746 10823
rect 17792 10777 17904 10823
rect 17950 10777 18062 10823
rect 18108 10777 18435 10823
rect 14393 10774 14431 10777
rect 14483 10774 14642 10777
rect 14694 10774 14853 10777
rect 14905 10774 18435 10777
rect 18487 10774 18645 10826
rect 18697 10774 18856 10826
rect 18908 10774 19068 10826
rect 19120 10774 19279 10826
rect 19331 10774 19489 10826
rect 19541 10774 19579 10826
rect 14393 10740 19579 10774
rect 19904 10826 20456 10860
rect 19904 10774 19943 10826
rect 19995 10823 20154 10826
rect 20206 10823 20365 10826
rect 20417 10823 20456 10826
rect 21875 10826 23974 10867
rect 21875 10823 21913 10826
rect 21965 10823 22124 10826
rect 22176 10823 22335 10826
rect 22387 10823 22545 10826
rect 22597 10823 22756 10826
rect 22808 10823 22968 10826
rect 23020 10823 23179 10826
rect 23231 10823 23389 10826
rect 19995 10777 20064 10823
rect 20110 10777 20154 10823
rect 20214 10777 20271 10823
rect 20317 10777 20365 10823
rect 20420 10777 20477 10823
rect 20523 10777 20580 10823
rect 20626 10777 20683 10823
rect 20729 10777 20786 10823
rect 20832 10777 20889 10823
rect 20935 10777 20992 10823
rect 21038 10777 21051 10823
rect 21386 10777 21399 10823
rect 23373 10777 23389 10823
rect 19995 10774 20154 10777
rect 20206 10774 20365 10777
rect 20417 10774 20456 10777
rect 19904 10740 20456 10774
rect 14393 10733 14943 10740
rect 12959 10682 13121 10693
rect 9334 10599 9463 10628
rect 9843 10610 9959 10647
rect 12959 10636 12970 10682
rect 13110 10636 13121 10682
rect 12959 10629 13121 10636
rect 9324 10553 9337 10599
rect 9383 10588 9459 10599
rect 9424 10553 9459 10588
rect 9505 10553 9582 10599
rect 9628 10553 9705 10599
rect 9751 10553 9764 10599
rect 9843 10564 9878 10610
rect 9924 10564 9959 10610
rect 9334 10536 9372 10553
rect 9424 10536 9463 10553
rect 9334 10509 9463 10536
rect 9334 10496 9462 10509
rect 9520 10373 9682 10413
rect 9520 10321 9591 10373
rect 9643 10321 9682 10373
rect 8605 10242 8618 10288
rect 8664 10242 8741 10288
rect 8787 10242 8864 10288
rect 8910 10242 8923 10288
rect 9089 10242 9238 10288
rect 9284 10242 9327 10288
rect 8611 10210 8920 10242
rect 9089 10210 9205 10242
rect 7450 10098 7758 10103
rect 6035 10064 6550 10098
rect 7036 10064 7758 10098
rect 8255 10078 8323 10200
rect 9520 10190 9682 10321
rect 9406 10187 9682 10190
rect 9406 10179 9591 10187
rect 9406 10133 9441 10179
rect 9487 10135 9591 10179
rect 9643 10166 9682 10187
rect 9843 10166 9959 10564
rect 10315 10588 13121 10629
rect 15181 10659 18143 10740
rect 18397 10733 19579 10740
rect 19905 10733 20456 10740
rect 21875 10774 21913 10777
rect 21965 10774 22124 10777
rect 22176 10774 22335 10777
rect 22387 10774 22545 10777
rect 22597 10774 22756 10777
rect 22808 10774 22968 10777
rect 23020 10774 23179 10777
rect 23231 10774 23389 10777
rect 23441 10774 23600 10826
rect 23652 10774 23811 10826
rect 23863 10774 23974 10826
rect 21875 10733 23974 10774
rect 15181 10613 15216 10659
rect 15262 10613 15374 10659
rect 15420 10613 15532 10659
rect 15578 10613 15690 10659
rect 15736 10613 15848 10659
rect 15894 10613 16006 10659
rect 16052 10613 16165 10659
rect 16211 10613 16323 10659
rect 16369 10613 16481 10659
rect 16527 10613 16639 10659
rect 16685 10613 16797 10659
rect 16843 10613 16955 10659
rect 17001 10613 17113 10659
rect 17159 10613 17272 10659
rect 17318 10613 17430 10659
rect 17476 10613 17588 10659
rect 17634 10613 17746 10659
rect 17792 10613 17904 10659
rect 17950 10613 18062 10659
rect 18108 10613 18143 10659
rect 23682 10699 23974 10733
rect 23682 10653 23820 10699
rect 23866 10653 23974 10699
rect 10315 10536 11532 10588
rect 11584 10536 13121 10588
rect 10315 10495 13121 10536
rect 14202 10553 14409 10599
rect 14455 10553 14522 10599
rect 14568 10553 14635 10599
rect 14681 10553 14748 10599
rect 14794 10553 14861 10599
rect 14907 10553 14920 10599
rect 15181 10577 18143 10613
rect 20632 10602 20940 10643
rect 20632 10599 20670 10602
rect 20722 10599 20850 10602
rect 20902 10599 20940 10602
rect 21186 10627 21254 10638
rect 13938 10487 14106 10498
rect 13938 10441 13955 10487
rect 14095 10441 14106 10487
rect 13938 10397 14106 10441
rect 11826 10357 14106 10397
rect 11826 10305 12665 10357
rect 12717 10305 14106 10357
rect 11826 10264 14106 10305
rect 14202 10166 14318 10553
rect 18502 10527 19474 10567
rect 20051 10553 20064 10599
rect 20110 10553 20168 10599
rect 20214 10553 20271 10599
rect 20317 10553 20374 10599
rect 20420 10553 20477 10599
rect 20523 10553 20580 10599
rect 20626 10553 20670 10599
rect 20729 10553 20786 10599
rect 20832 10553 20850 10599
rect 20935 10553 20992 10599
rect 21038 10553 21051 10599
rect 18502 10512 18540 10527
rect 18592 10512 18751 10527
rect 18803 10512 18962 10527
rect 19014 10512 19173 10527
rect 19225 10512 19384 10527
rect 19436 10512 19474 10527
rect 18362 10466 18375 10512
rect 18421 10466 18478 10512
rect 18524 10475 18540 10512
rect 18524 10466 18581 10475
rect 18627 10466 18684 10512
rect 18730 10475 18751 10512
rect 18730 10466 18787 10475
rect 18833 10466 18890 10512
rect 18936 10475 18962 10512
rect 18936 10466 18993 10475
rect 19039 10466 19096 10512
rect 19142 10475 19173 10512
rect 19142 10466 19199 10475
rect 19449 10466 19474 10512
rect 20632 10550 20670 10553
rect 20722 10550 20850 10553
rect 20902 10550 20940 10553
rect 20632 10510 20940 10550
rect 18154 10420 18284 10461
rect 18502 10435 19474 10466
rect 14498 10375 14838 10404
rect 14396 10329 14409 10375
rect 14455 10329 14522 10375
rect 14568 10364 14635 10375
rect 14588 10329 14635 10364
rect 14681 10329 14748 10375
rect 14794 10364 14861 10375
rect 14800 10329 14861 10364
rect 14907 10329 14920 10375
rect 18154 10368 18193 10420
rect 18245 10368 18284 10420
rect 18154 10365 18284 10368
rect 14498 10312 14536 10329
rect 14588 10312 14748 10329
rect 14800 10312 14838 10329
rect 14498 10271 14838 10312
rect 14997 10256 17976 10289
rect 14997 10210 15061 10256
rect 15201 10248 17976 10256
rect 15201 10210 16705 10248
rect 14997 10196 16705 10210
rect 16757 10196 17976 10248
rect 9643 10151 14515 10166
rect 14997 10155 17976 10196
rect 18154 10225 18219 10365
rect 18265 10225 18284 10365
rect 19859 10375 20409 10404
rect 19859 10364 20064 10375
rect 20110 10364 20168 10375
rect 19417 10288 19757 10329
rect 18362 10242 18375 10288
rect 18421 10242 18478 10288
rect 18524 10242 18581 10288
rect 18627 10242 18684 10288
rect 18730 10242 18787 10288
rect 18833 10242 18890 10288
rect 18936 10242 18993 10288
rect 19039 10242 19096 10288
rect 19142 10242 19199 10288
rect 19449 10242 19757 10288
rect 19859 10312 19897 10364
rect 19949 10329 20064 10364
rect 20160 10329 20168 10364
rect 20214 10329 20271 10375
rect 20317 10364 20374 10375
rect 20317 10329 20319 10364
rect 19949 10312 20108 10329
rect 20160 10312 20319 10329
rect 20371 10329 20374 10364
rect 20420 10329 20477 10375
rect 20523 10329 20580 10375
rect 20626 10329 20683 10375
rect 20729 10329 20786 10375
rect 20832 10329 20889 10375
rect 20935 10329 20992 10375
rect 21038 10329 21051 10375
rect 20371 10312 20409 10329
rect 19859 10271 20409 10312
rect 18154 10202 18284 10225
rect 19417 10210 19757 10242
rect 9643 10135 14409 10151
rect 9487 10133 14409 10135
rect 9406 10130 14409 10133
rect 9406 10084 13336 10130
rect 13382 10084 13503 10130
rect 13549 10084 13668 10130
rect 13714 10084 13833 10130
rect 13879 10105 14409 10130
rect 14455 10105 14522 10151
rect 14568 10105 14635 10151
rect 14681 10105 14748 10151
rect 14794 10105 14861 10151
rect 14907 10105 14920 10151
rect 18154 10150 18193 10202
rect 18245 10150 18284 10202
rect 18154 10110 18284 10150
rect 19641 10153 19757 10210
rect 21186 10205 21197 10627
rect 21243 10205 21254 10627
rect 21394 10599 21702 10636
rect 21386 10553 21399 10599
rect 23373 10553 23386 10599
rect 21394 10543 21432 10553
rect 21484 10543 21612 10553
rect 21664 10543 21702 10553
rect 21394 10503 21702 10543
rect 23682 10535 23974 10653
rect 23682 10489 23820 10535
rect 23866 10489 23974 10535
rect 23682 10397 23974 10489
rect 23182 10375 23974 10397
rect 21386 10329 21399 10375
rect 23373 10329 23974 10375
rect 23182 10278 23974 10329
rect 21186 10153 21254 10205
rect 19641 10116 21254 10153
rect 21394 10151 21702 10173
rect 13879 10084 14515 10105
rect 8255 10064 9320 10078
rect 345 10000 452 10046
rect 498 10000 637 10046
rect 3081 10033 4240 10062
rect 4857 10018 4870 10064
rect 5120 10018 5140 10064
rect 5223 10018 5280 10064
rect 5326 10018 5351 10064
rect 5429 10018 5486 10064
rect 5532 10018 5562 10064
rect 5635 10018 5692 10064
rect 5738 10018 5773 10064
rect 5841 10018 5898 10064
rect 5944 10018 5957 10064
rect 6035 10018 6451 10064
rect 6497 10018 6568 10064
rect 6614 10018 6685 10064
rect 6731 10018 6803 10064
rect 6849 10018 6921 10064
rect 6967 10018 7039 10064
rect 7085 10062 7506 10064
rect 7085 10018 7488 10062
rect 7552 10018 7623 10064
rect 7669 10062 7740 10064
rect 7720 10018 7740 10062
rect 7786 10018 7858 10064
rect 7904 10018 7976 10064
rect 8022 10018 8094 10064
rect 8140 10018 8153 10064
rect 8255 10018 8618 10064
rect 8664 10018 8741 10064
rect 8787 10018 8864 10064
rect 8910 10018 9238 10064
rect 9284 10018 9327 10064
rect 9406 10046 14515 10084
rect 18502 10064 19474 10104
rect 18362 10018 18375 10064
rect 18421 10018 18478 10064
rect 18524 10018 18540 10064
rect 18627 10018 18684 10064
rect 18730 10018 18751 10064
rect 18833 10018 18890 10064
rect 18936 10018 18962 10064
rect 19039 10018 19096 10064
rect 19142 10018 19173 10064
rect 19449 10018 19474 10064
rect 19641 10070 20113 10116
rect 20159 10070 20300 10116
rect 20346 10070 20487 10116
rect 20533 10070 20673 10116
rect 20719 10070 20860 10116
rect 20906 10070 21254 10116
rect 21386 10105 21399 10151
rect 23373 10105 23386 10151
rect 19641 10060 21254 10070
rect 20078 10033 21254 10060
rect 21394 10080 21432 10105
rect 21484 10080 21612 10105
rect 21664 10080 21702 10105
rect 21394 10040 21702 10080
rect 23682 10046 23974 10278
rect 345 9967 637 10000
rect 4891 10012 4929 10018
rect 4981 10012 5140 10018
rect 5192 10012 5351 10018
rect 5403 10012 5562 10018
rect 5614 10012 5773 10018
rect 5825 10012 5863 10018
rect 4467 9967 4622 9974
rect 4891 9972 5863 10012
rect 6035 9978 6550 10018
rect 7036 10010 7488 10018
rect 7540 10010 7668 10018
rect 7720 10010 7758 10018
rect 7036 9978 7758 10010
rect 7450 9970 7758 9978
rect 345 9926 2439 9967
rect 345 9874 451 9926
rect 503 9874 662 9926
rect 714 9874 873 9926
rect 925 9874 1083 9926
rect 1135 9874 1294 9926
rect 1346 9874 1506 9926
rect 1558 9874 1717 9926
rect 1769 9874 1927 9926
rect 1979 9874 2138 9926
rect 2190 9874 2349 9926
rect 2401 9874 2439 9926
rect 345 9833 2439 9874
rect 4314 9926 4622 9967
rect 8255 9958 9320 10018
rect 18502 10012 18540 10018
rect 18592 10012 18751 10018
rect 18803 10012 18962 10018
rect 19014 10012 19173 10018
rect 19225 10012 19384 10018
rect 19436 10012 19474 10018
rect 18502 9972 19474 10012
rect 23682 10000 23820 10046
rect 23866 10000 23974 10046
rect 19696 9967 19852 9974
rect 23682 9967 23974 10000
rect 4314 9874 4352 9926
rect 4404 9923 4532 9926
rect 4404 9877 4513 9923
rect 4404 9874 4532 9877
rect 4584 9874 4622 9926
rect 4314 9833 4622 9874
rect 19696 9926 20005 9967
rect 19696 9874 19735 9926
rect 19787 9923 19915 9926
rect 19803 9877 19915 9923
rect 19787 9874 19915 9877
rect 19967 9874 20005 9926
rect 345 9800 637 9833
rect 4467 9826 4622 9833
rect 345 9754 452 9800
rect 498 9754 637 9800
rect 4891 9788 5863 9828
rect 7450 9822 7758 9830
rect 4891 9782 4929 9788
rect 4981 9782 5140 9788
rect 5192 9782 5351 9788
rect 5403 9782 5562 9788
rect 5614 9782 5773 9788
rect 5825 9782 5863 9788
rect 6035 9782 6550 9822
rect 7036 9790 7758 9822
rect 7036 9782 7488 9790
rect 7540 9782 7668 9790
rect 7720 9782 7758 9790
rect 8255 9782 9320 9842
rect 19696 9833 20005 9874
rect 21875 9926 23974 9967
rect 21875 9874 21913 9926
rect 21965 9874 22124 9926
rect 22176 9874 22335 9926
rect 22387 9874 22545 9926
rect 22597 9874 22756 9926
rect 22808 9874 22968 9926
rect 23020 9874 23179 9926
rect 23231 9874 23389 9926
rect 23441 9874 23600 9926
rect 23652 9874 23811 9926
rect 23863 9874 23974 9926
rect 21875 9833 23974 9874
rect 18502 9788 19474 9828
rect 19696 9826 19852 9833
rect 18502 9782 18540 9788
rect 18592 9782 18751 9788
rect 18803 9782 18962 9788
rect 19014 9782 19173 9788
rect 19225 9782 19384 9788
rect 19436 9782 19474 9788
rect 345 9637 637 9754
rect 3081 9738 4240 9767
rect 2616 9698 2924 9738
rect 2616 9695 2654 9698
rect 2706 9695 2834 9698
rect 2886 9695 2924 9698
rect 3081 9730 4679 9738
rect 4857 9736 4870 9782
rect 5120 9736 5140 9782
rect 5223 9736 5280 9782
rect 5326 9736 5351 9782
rect 5429 9736 5486 9782
rect 5532 9736 5562 9782
rect 5635 9736 5692 9782
rect 5738 9736 5773 9782
rect 5841 9736 5898 9782
rect 5944 9736 5957 9782
rect 6035 9736 6451 9782
rect 6497 9736 6568 9782
rect 6614 9736 6685 9782
rect 6731 9736 6803 9782
rect 6849 9736 6921 9782
rect 6967 9736 7039 9782
rect 7085 9738 7488 9782
rect 7085 9736 7506 9738
rect 7552 9736 7623 9782
rect 7720 9738 7740 9782
rect 7669 9736 7740 9738
rect 7786 9736 7858 9782
rect 7904 9736 7976 9782
rect 8022 9736 8094 9782
rect 8140 9736 8153 9782
rect 8255 9736 8618 9782
rect 8664 9736 8741 9782
rect 8787 9736 8864 9782
rect 8910 9736 9238 9782
rect 9284 9736 9327 9782
rect 933 9649 946 9695
rect 2920 9649 2933 9695
rect 3081 9684 3413 9730
rect 3459 9684 3599 9730
rect 3645 9684 3786 9730
rect 3832 9684 3973 9730
rect 4019 9684 4159 9730
rect 4205 9684 4679 9730
rect 4891 9696 5863 9736
rect 6035 9702 6550 9736
rect 7036 9702 7758 9736
rect 345 9591 452 9637
rect 498 9591 637 9637
rect 2616 9646 2654 9649
rect 2706 9646 2834 9649
rect 2886 9646 2924 9649
rect 2616 9605 2924 9646
rect 3081 9647 4679 9684
rect 345 9522 637 9591
rect 3081 9565 3149 9647
rect 345 9474 1090 9522
rect 345 9428 452 9474
rect 498 9471 1090 9474
rect 498 9428 946 9471
rect 345 9425 946 9428
rect 2920 9425 2933 9471
rect 345 9403 1090 9425
rect 345 9311 637 9403
rect 345 9265 452 9311
rect 498 9265 637 9311
rect 345 9147 637 9265
rect 2616 9250 2924 9290
rect 2616 9247 2654 9250
rect 2706 9247 2834 9250
rect 2886 9247 2924 9250
rect 933 9201 946 9247
rect 2920 9201 2933 9247
rect 2616 9198 2654 9201
rect 2706 9198 2834 9201
rect 2886 9198 2924 9201
rect 2616 9157 2924 9198
rect 345 9101 452 9147
rect 498 9101 637 9147
rect 3081 9143 3092 9565
rect 3138 9143 3149 9565
rect 4561 9590 4679 9647
rect 6035 9602 6151 9702
rect 7450 9697 7758 9702
rect 8255 9722 9320 9736
rect 4561 9558 5957 9590
rect 3825 9488 4315 9529
rect 3825 9471 3864 9488
rect 3916 9471 4044 9488
rect 4096 9471 4224 9488
rect 3268 9425 3281 9471
rect 3327 9425 3384 9471
rect 3430 9425 3487 9471
rect 3533 9425 3590 9471
rect 3636 9425 3693 9471
rect 3739 9425 3796 9471
rect 3842 9436 3864 9471
rect 3842 9425 3899 9436
rect 3945 9425 4002 9471
rect 4096 9436 4105 9471
rect 4048 9425 4105 9436
rect 4151 9425 4209 9471
rect 4276 9436 4315 9488
rect 4561 9512 4870 9558
rect 5120 9512 5177 9558
rect 5223 9512 5280 9558
rect 5326 9512 5383 9558
rect 5429 9512 5486 9558
rect 5532 9512 5589 9558
rect 5635 9512 5692 9558
rect 5738 9512 5795 9558
rect 5841 9512 5898 9558
rect 5944 9512 5957 9558
rect 4561 9468 5957 9512
rect 4255 9425 4315 9436
rect 3825 9396 4315 9425
rect 6035 9462 6072 9602
rect 6118 9462 6151 9602
rect 4891 9334 5863 9368
rect 6035 9359 6151 9462
rect 6237 9602 6370 9622
rect 6237 9563 6294 9602
rect 6237 9511 6275 9563
rect 6237 9462 6294 9511
rect 6340 9462 6370 9602
rect 8255 9600 8323 9722
rect 9406 9716 14515 9754
rect 18362 9736 18375 9782
rect 18421 9736 18478 9782
rect 18524 9736 18540 9782
rect 18627 9736 18684 9782
rect 18730 9736 18751 9782
rect 18833 9736 18890 9782
rect 18936 9736 18962 9782
rect 19039 9736 19096 9782
rect 19142 9736 19173 9782
rect 19449 9736 19474 9782
rect 23682 9800 23974 9833
rect 20078 9740 21254 9767
rect 9406 9670 13336 9716
rect 13382 9670 13503 9716
rect 13549 9670 13668 9716
rect 13714 9670 13833 9716
rect 13879 9695 14515 9716
rect 18502 9696 19474 9736
rect 19641 9730 21254 9740
rect 13879 9670 14409 9695
rect 9406 9667 14409 9670
rect 9406 9621 9441 9667
rect 9487 9665 14409 9667
rect 9487 9621 9591 9665
rect 9406 9613 9591 9621
rect 9643 9649 14409 9665
rect 14455 9649 14522 9695
rect 14568 9649 14635 9695
rect 14681 9649 14748 9695
rect 14794 9649 14861 9695
rect 14907 9649 14920 9695
rect 18154 9650 18284 9690
rect 9643 9634 14515 9649
rect 9643 9613 9682 9634
rect 9406 9610 9682 9613
rect 6521 9590 7282 9597
rect 6520 9558 7528 9590
rect 6438 9512 6451 9558
rect 6497 9556 6568 9558
rect 6497 9512 6558 9556
rect 6614 9512 6685 9558
rect 6731 9556 6803 9558
rect 6731 9512 6769 9556
rect 6849 9512 6921 9558
rect 6967 9556 7039 9558
rect 6967 9512 6981 9556
rect 6520 9504 6558 9512
rect 6610 9504 6769 9512
rect 6821 9504 6981 9512
rect 7033 9512 7039 9556
rect 7085 9556 7506 9558
rect 7085 9512 7192 9556
rect 7033 9504 7192 9512
rect 7244 9512 7506 9556
rect 7552 9512 7623 9558
rect 7669 9512 7740 9558
rect 7786 9512 7858 9558
rect 7904 9512 7976 9558
rect 8022 9512 8094 9558
rect 8140 9512 8153 9558
rect 7244 9504 7528 9512
rect 6520 9471 7528 9504
rect 6520 9470 7282 9471
rect 6521 9464 7282 9470
rect 6237 9439 6370 9462
rect 8255 9460 8266 9600
rect 8312 9460 8323 9600
rect 8611 9558 8920 9590
rect 9089 9558 9205 9590
rect 8605 9512 8618 9558
rect 8664 9512 8741 9558
rect 8787 9512 8864 9558
rect 8910 9512 8923 9558
rect 9089 9512 9238 9558
rect 9284 9512 9327 9558
rect 8255 9449 8323 9460
rect 6035 9334 6550 9359
rect 7036 9356 7528 9359
rect 7036 9334 7758 9356
rect 4857 9288 4870 9334
rect 5120 9328 5177 9334
rect 5120 9288 5140 9328
rect 5223 9288 5280 9334
rect 5326 9328 5383 9334
rect 5326 9288 5351 9328
rect 5429 9288 5486 9334
rect 5532 9328 5589 9334
rect 5532 9288 5562 9328
rect 5635 9288 5692 9334
rect 5738 9328 5795 9334
rect 5738 9288 5773 9328
rect 5841 9288 5898 9334
rect 5944 9288 5957 9334
rect 6035 9288 6451 9334
rect 6497 9288 6568 9334
rect 6614 9288 6685 9334
rect 6731 9288 6803 9334
rect 6849 9288 6921 9334
rect 6967 9288 7039 9334
rect 7085 9316 7506 9334
rect 7085 9288 7488 9316
rect 7552 9288 7623 9334
rect 7669 9316 7740 9334
rect 7720 9288 7740 9316
rect 7786 9288 7858 9334
rect 7904 9288 7976 9334
rect 8022 9288 8094 9334
rect 8140 9288 8153 9334
rect 3378 9247 3686 9282
rect 4891 9276 4929 9288
rect 4981 9276 5140 9288
rect 5192 9276 5351 9288
rect 5403 9276 5562 9288
rect 5614 9276 5773 9288
rect 5825 9276 5863 9288
rect 3268 9201 3281 9247
rect 3327 9201 3384 9247
rect 3430 9242 3487 9247
rect 3468 9201 3487 9242
rect 3533 9201 3590 9247
rect 3636 9242 3693 9247
rect 3648 9201 3693 9242
rect 3739 9201 3796 9247
rect 3842 9201 3899 9247
rect 3945 9201 4002 9247
rect 4048 9201 4105 9247
rect 4151 9201 4209 9247
rect 4255 9201 4268 9247
rect 4891 9236 5863 9276
rect 6035 9239 6550 9288
rect 7036 9264 7488 9288
rect 7540 9264 7668 9288
rect 7720 9264 7758 9288
rect 7036 9239 7758 9264
rect 7450 9223 7758 9239
rect 3378 9190 3416 9201
rect 3468 9190 3596 9201
rect 3648 9190 3686 9201
rect 3378 9149 3686 9190
rect 3081 9132 3149 9143
rect 345 9067 637 9101
rect 345 9026 2439 9067
rect 3844 9060 4605 9067
rect 345 8974 451 9026
rect 503 8974 662 9026
rect 714 8974 873 9026
rect 925 9023 1083 9026
rect 1135 9023 1294 9026
rect 1346 9023 1506 9026
rect 1558 9023 1717 9026
rect 1769 9023 1927 9026
rect 1979 9023 2138 9026
rect 2190 9023 2349 9026
rect 2401 9023 2439 9026
rect 3843 9026 4605 9060
rect 3843 9023 3881 9026
rect 3933 9023 4092 9026
rect 4144 9023 4304 9026
rect 925 8977 946 9023
rect 2920 8977 2933 9023
rect 3268 8977 3281 9023
rect 3327 8977 3384 9023
rect 3430 8977 3487 9023
rect 3533 8977 3590 9023
rect 3636 8977 3693 9023
rect 3739 8977 3796 9023
rect 3842 8977 3881 9023
rect 3945 8977 4002 9023
rect 4048 8977 4092 9023
rect 4151 8977 4209 9023
rect 4255 8977 4304 9023
rect 925 8974 1083 8977
rect 1135 8974 1294 8977
rect 1346 8974 1506 8977
rect 1558 8974 1717 8977
rect 1769 8974 1927 8977
rect 1979 8974 2138 8977
rect 2190 8974 2349 8977
rect 2401 8974 2439 8977
rect 345 8933 2439 8974
rect 3843 8974 3881 8977
rect 3933 8974 4092 8977
rect 4144 8974 4304 8977
rect 4356 8974 4515 9026
rect 4567 8974 4605 9026
rect 3843 8940 4605 8974
rect 3844 8933 4605 8940
rect 4779 9060 5961 9067
rect 4779 9026 6555 9060
rect 4779 8974 4817 9026
rect 4869 8974 5027 9026
rect 5079 8974 5238 9026
rect 5290 8974 5450 9026
rect 5502 8974 5661 9026
rect 5713 8974 5871 9026
rect 5923 9023 6555 9026
rect 5923 8977 6086 9023
rect 6320 8977 6555 9023
rect 5923 8974 6555 8977
rect 4779 8940 6555 8974
rect 7543 9026 8439 9067
rect 7543 9023 7927 9026
rect 7979 9023 8138 9026
rect 7543 8977 7554 9023
rect 8070 8977 8138 9023
rect 7543 8974 7927 8977
rect 7979 8974 8138 8977
rect 8190 8974 8349 9026
rect 8401 8974 8439 9026
rect 4779 8933 5961 8940
rect 7543 8933 8439 8974
rect 8611 9026 8920 9512
rect 8611 8974 8649 9026
rect 8701 9023 8829 9026
rect 8705 8977 8817 9023
rect 8701 8974 8829 8977
rect 8881 8974 8920 9026
rect 345 8899 637 8933
rect 345 8853 452 8899
rect 498 8853 637 8899
rect 345 8735 637 8853
rect 3081 8857 3149 8868
rect 2616 8802 2924 8843
rect 2616 8799 2654 8802
rect 2706 8799 2834 8802
rect 2886 8799 2924 8802
rect 933 8753 946 8799
rect 2920 8753 2933 8799
rect 345 8689 452 8735
rect 498 8689 637 8735
rect 2616 8750 2654 8753
rect 2706 8750 2834 8753
rect 2886 8750 2924 8753
rect 2616 8710 2924 8750
rect 345 8597 637 8689
rect 345 8575 1090 8597
rect 345 8572 946 8575
rect 345 8526 452 8572
rect 498 8529 946 8572
rect 2920 8529 2933 8575
rect 498 8526 1090 8529
rect 345 8478 1090 8526
rect 345 8409 637 8478
rect 345 8363 452 8409
rect 498 8363 637 8409
rect 3081 8435 3092 8857
rect 3138 8435 3149 8857
rect 3378 8810 3686 8851
rect 3378 8799 3416 8810
rect 3468 8799 3596 8810
rect 3648 8799 3686 8810
rect 3268 8753 3281 8799
rect 3327 8753 3384 8799
rect 3468 8758 3487 8799
rect 3430 8753 3487 8758
rect 3533 8753 3590 8799
rect 3648 8758 3693 8799
rect 3636 8753 3693 8758
rect 3739 8753 3796 8799
rect 3842 8753 3899 8799
rect 3945 8753 4002 8799
rect 4048 8753 4105 8799
rect 4151 8753 4209 8799
rect 4255 8753 4268 8799
rect 3378 8718 3686 8753
rect 4891 8724 5863 8764
rect 7450 8761 7758 8777
rect 4891 8712 4929 8724
rect 4981 8712 5140 8724
rect 5192 8712 5351 8724
rect 5403 8712 5562 8724
rect 5614 8712 5773 8724
rect 5825 8712 5863 8724
rect 6035 8712 6550 8761
rect 7036 8736 7758 8761
rect 7036 8712 7488 8736
rect 7540 8712 7668 8736
rect 7720 8712 7758 8736
rect 4857 8666 4870 8712
rect 5120 8672 5140 8712
rect 5120 8666 5177 8672
rect 5223 8666 5280 8712
rect 5326 8672 5351 8712
rect 5326 8666 5383 8672
rect 5429 8666 5486 8712
rect 5532 8672 5562 8712
rect 5532 8666 5589 8672
rect 5635 8666 5692 8712
rect 5738 8672 5773 8712
rect 5738 8666 5795 8672
rect 5841 8666 5898 8712
rect 5944 8666 5957 8712
rect 6035 8666 6451 8712
rect 6497 8666 6568 8712
rect 6614 8666 6685 8712
rect 6731 8666 6803 8712
rect 6849 8666 6921 8712
rect 6967 8666 7039 8712
rect 7085 8684 7488 8712
rect 7085 8666 7506 8684
rect 7552 8666 7623 8712
rect 7720 8684 7740 8712
rect 7669 8666 7740 8684
rect 7786 8666 7858 8712
rect 7904 8666 7976 8712
rect 8022 8666 8094 8712
rect 8140 8666 8153 8712
rect 4891 8632 5863 8666
rect 6035 8641 6550 8666
rect 7036 8644 7758 8666
rect 7036 8641 7528 8644
rect 3825 8575 4315 8604
rect 3268 8529 3281 8575
rect 3327 8529 3384 8575
rect 3430 8529 3487 8575
rect 3533 8529 3590 8575
rect 3636 8529 3693 8575
rect 3739 8529 3796 8575
rect 3842 8564 3899 8575
rect 3842 8529 3864 8564
rect 3945 8529 4002 8575
rect 4048 8564 4105 8575
rect 4096 8529 4105 8564
rect 4151 8529 4209 8575
rect 4255 8564 4315 8575
rect 3825 8512 3864 8529
rect 3916 8512 4044 8529
rect 4096 8512 4224 8529
rect 4276 8512 4315 8564
rect 6035 8538 6151 8641
rect 3825 8471 4315 8512
rect 4561 8488 5957 8532
rect 345 8246 637 8363
rect 2616 8354 2924 8395
rect 2616 8351 2654 8354
rect 2706 8351 2834 8354
rect 2886 8351 2924 8354
rect 3081 8353 3149 8435
rect 4561 8442 4870 8488
rect 5120 8442 5177 8488
rect 5223 8442 5280 8488
rect 5326 8442 5383 8488
rect 5429 8442 5486 8488
rect 5532 8442 5589 8488
rect 5635 8442 5692 8488
rect 5738 8442 5795 8488
rect 5841 8442 5898 8488
rect 5944 8442 5957 8488
rect 4561 8410 5957 8442
rect 4561 8353 4679 8410
rect 933 8305 946 8351
rect 2920 8305 2933 8351
rect 3081 8316 4679 8353
rect 2616 8302 2654 8305
rect 2706 8302 2834 8305
rect 2886 8302 2924 8305
rect 2616 8262 2924 8302
rect 3081 8270 3413 8316
rect 3459 8270 3599 8316
rect 3645 8270 3786 8316
rect 3832 8270 3973 8316
rect 4019 8270 4159 8316
rect 4205 8270 4679 8316
rect 6035 8398 6072 8538
rect 6118 8398 6151 8538
rect 3081 8262 4679 8270
rect 4891 8264 5863 8304
rect 6035 8298 6151 8398
rect 6237 8538 6370 8561
rect 6237 8489 6294 8538
rect 6237 8437 6275 8489
rect 6237 8398 6294 8437
rect 6340 8398 6370 8538
rect 8255 8540 8323 8551
rect 6521 8530 7282 8536
rect 6520 8529 7282 8530
rect 6520 8496 7528 8529
rect 6520 8488 6558 8496
rect 6610 8488 6769 8496
rect 6821 8488 6981 8496
rect 6438 8442 6451 8488
rect 6497 8444 6558 8488
rect 6497 8442 6568 8444
rect 6614 8442 6685 8488
rect 6731 8444 6769 8488
rect 6731 8442 6803 8444
rect 6849 8442 6921 8488
rect 6967 8444 6981 8488
rect 7033 8488 7192 8496
rect 7033 8444 7039 8488
rect 6967 8442 7039 8444
rect 7085 8444 7192 8488
rect 7244 8488 7528 8496
rect 7244 8444 7506 8488
rect 7085 8442 7506 8444
rect 7552 8442 7623 8488
rect 7669 8442 7740 8488
rect 7786 8442 7858 8488
rect 7904 8442 7976 8488
rect 8022 8442 8094 8488
rect 8140 8442 8153 8488
rect 6520 8410 7528 8442
rect 6521 8403 7282 8410
rect 6237 8378 6370 8398
rect 8255 8400 8266 8540
rect 8312 8400 8323 8540
rect 8611 8488 8920 8974
rect 9089 9060 9205 9512
rect 9520 9479 9682 9610
rect 9520 9427 9591 9479
rect 9643 9427 9682 9479
rect 9520 9387 9682 9427
rect 9334 9291 9462 9304
rect 9334 9264 9463 9291
rect 9334 9247 9372 9264
rect 9424 9247 9463 9264
rect 9324 9201 9337 9247
rect 9424 9212 9459 9247
rect 9383 9201 9459 9212
rect 9505 9201 9582 9247
rect 9628 9201 9705 9247
rect 9751 9201 9764 9247
rect 9843 9236 9959 9634
rect 11826 9495 14106 9536
rect 11826 9443 12665 9495
rect 12717 9443 14106 9495
rect 11826 9403 14106 9443
rect 13938 9359 14106 9403
rect 13938 9313 13955 9359
rect 14095 9313 14106 9359
rect 9334 9172 9463 9201
rect 9843 9190 9878 9236
rect 9924 9190 9959 9236
rect 9843 9153 9959 9190
rect 10315 9264 13121 9305
rect 13938 9302 14106 9313
rect 10315 9212 11532 9264
rect 11584 9212 13121 9264
rect 10315 9171 13121 9212
rect 14202 9247 14318 9634
rect 14997 9604 17976 9645
rect 14997 9590 17083 9604
rect 14997 9544 15061 9590
rect 15201 9552 17083 9590
rect 17135 9552 17976 9604
rect 15201 9544 17976 9552
rect 14498 9488 14838 9529
rect 14997 9511 17976 9544
rect 18154 9598 18193 9650
rect 18245 9598 18284 9650
rect 18154 9575 18284 9598
rect 19641 9684 20113 9730
rect 20159 9684 20300 9730
rect 20346 9684 20487 9730
rect 20533 9684 20673 9730
rect 20719 9684 20860 9730
rect 20906 9684 21254 9730
rect 21394 9720 21702 9760
rect 21394 9695 21432 9720
rect 21484 9695 21612 9720
rect 21664 9695 21702 9720
rect 23682 9754 23820 9800
rect 23866 9754 23974 9800
rect 19641 9647 21254 9684
rect 21386 9649 21399 9695
rect 23373 9649 23386 9695
rect 19641 9590 19757 9647
rect 14498 9471 14536 9488
rect 14588 9471 14748 9488
rect 14800 9471 14838 9488
rect 14396 9425 14409 9471
rect 14455 9425 14522 9471
rect 14588 9436 14635 9471
rect 14568 9425 14635 9436
rect 14681 9425 14748 9471
rect 14800 9436 14861 9471
rect 14794 9425 14861 9436
rect 14907 9425 14920 9471
rect 18154 9435 18219 9575
rect 18265 9435 18284 9575
rect 19417 9558 19757 9590
rect 18362 9512 18375 9558
rect 18421 9512 18478 9558
rect 18524 9512 18581 9558
rect 18627 9512 18684 9558
rect 18730 9512 18787 9558
rect 18833 9512 18890 9558
rect 18936 9512 18993 9558
rect 19039 9512 19096 9558
rect 19142 9512 19199 9558
rect 19449 9512 19757 9558
rect 21186 9595 21254 9647
rect 21394 9627 21702 9649
rect 19417 9471 19757 9512
rect 19859 9488 20409 9529
rect 18154 9432 18284 9435
rect 14498 9396 14838 9425
rect 18154 9380 18193 9432
rect 18245 9380 18284 9432
rect 19859 9436 19897 9488
rect 19949 9471 20108 9488
rect 20160 9471 20319 9488
rect 19949 9436 20064 9471
rect 20160 9436 20168 9471
rect 19859 9425 20064 9436
rect 20110 9425 20168 9436
rect 20214 9425 20271 9471
rect 20317 9436 20319 9471
rect 20371 9471 20409 9488
rect 20371 9436 20374 9471
rect 20317 9425 20374 9436
rect 20420 9425 20477 9471
rect 20523 9425 20580 9471
rect 20626 9425 20683 9471
rect 20729 9425 20786 9471
rect 20832 9425 20889 9471
rect 20935 9425 20992 9471
rect 21038 9425 21051 9471
rect 19859 9396 20409 9425
rect 18154 9339 18284 9380
rect 18502 9334 19474 9365
rect 18362 9288 18375 9334
rect 18421 9288 18478 9334
rect 18524 9325 18581 9334
rect 18524 9288 18540 9325
rect 18627 9288 18684 9334
rect 18730 9325 18787 9334
rect 18730 9288 18751 9325
rect 18833 9288 18890 9334
rect 18936 9325 18993 9334
rect 18936 9288 18962 9325
rect 19039 9288 19096 9334
rect 19142 9325 19199 9334
rect 19142 9288 19173 9325
rect 19449 9288 19474 9334
rect 18502 9273 18540 9288
rect 18592 9273 18751 9288
rect 18803 9273 18962 9288
rect 19014 9273 19173 9288
rect 19225 9273 19384 9288
rect 19436 9273 19474 9288
rect 14202 9201 14409 9247
rect 14455 9201 14522 9247
rect 14568 9201 14635 9247
rect 14681 9201 14748 9247
rect 14794 9201 14861 9247
rect 14907 9201 14920 9247
rect 18502 9233 19474 9273
rect 20632 9250 20940 9290
rect 20632 9247 20670 9250
rect 20722 9247 20850 9250
rect 20902 9247 20940 9250
rect 12959 9164 13121 9171
rect 12959 9118 12970 9164
rect 13110 9118 13121 9164
rect 12959 9107 13121 9118
rect 15181 9187 18143 9223
rect 20051 9201 20064 9247
rect 20110 9201 20168 9247
rect 20214 9201 20271 9247
rect 20317 9201 20374 9247
rect 20420 9201 20477 9247
rect 20523 9201 20580 9247
rect 20626 9201 20670 9247
rect 20729 9201 20786 9247
rect 20832 9201 20850 9247
rect 20935 9201 20992 9247
rect 21038 9201 21051 9247
rect 15181 9141 15216 9187
rect 15262 9141 15374 9187
rect 15420 9141 15532 9187
rect 15578 9141 15690 9187
rect 15736 9141 15848 9187
rect 15894 9141 16006 9187
rect 16052 9141 16165 9187
rect 16211 9141 16323 9187
rect 16369 9141 16481 9187
rect 16527 9141 16639 9187
rect 16685 9141 16797 9187
rect 16843 9141 16955 9187
rect 17001 9141 17113 9187
rect 17159 9141 17272 9187
rect 17318 9141 17430 9187
rect 17476 9141 17588 9187
rect 17634 9141 17746 9187
rect 17792 9141 17904 9187
rect 17950 9141 18062 9187
rect 18108 9141 18143 9187
rect 20632 9198 20670 9201
rect 20722 9198 20850 9201
rect 20902 9198 20940 9201
rect 20632 9157 20940 9198
rect 21186 9173 21197 9595
rect 21243 9173 21254 9595
rect 23682 9522 23974 9754
rect 23182 9471 23974 9522
rect 21386 9425 21399 9471
rect 23373 9425 23974 9471
rect 23182 9403 23974 9425
rect 23682 9311 23974 9403
rect 21394 9257 21702 9297
rect 21394 9247 21432 9257
rect 21484 9247 21612 9257
rect 21664 9247 21702 9257
rect 23682 9265 23820 9311
rect 23866 9265 23974 9311
rect 21386 9201 21399 9247
rect 23373 9201 23386 9247
rect 21186 9162 21254 9173
rect 21394 9164 21702 9201
rect 9812 9060 10120 9067
rect 10385 9060 12583 9074
rect 13350 9060 14111 9067
rect 9089 9037 12583 9060
rect 13301 9037 14111 9060
rect 9089 9026 14111 9037
rect 9089 9023 9850 9026
rect 9089 8977 9337 9023
rect 9383 8977 9459 9023
rect 9505 8977 9582 9023
rect 9628 8977 9705 9023
rect 9751 8977 9850 9023
rect 9089 8974 9850 8977
rect 9902 8974 10030 9026
rect 10082 9023 13387 9026
rect 10082 8977 10433 9023
rect 10479 8977 10591 9023
rect 10637 8977 10749 9023
rect 10795 8977 10907 9023
rect 10953 8977 11066 9023
rect 11112 8977 11224 9023
rect 11270 8977 11382 9023
rect 11428 8977 11540 9023
rect 11586 8977 11698 9023
rect 11744 8977 11856 9023
rect 11902 8977 12015 9023
rect 12061 8977 12173 9023
rect 12219 8977 12331 9023
rect 12377 8977 12489 9023
rect 12535 8977 13336 9023
rect 13382 8977 13387 9023
rect 10082 8974 13387 8977
rect 13439 9023 13598 9026
rect 13439 8977 13503 9023
rect 13549 8977 13598 9023
rect 13439 8974 13598 8977
rect 13650 9023 13810 9026
rect 13862 9023 14021 9026
rect 13650 8977 13668 9023
rect 13714 8977 13810 9023
rect 13879 8977 14021 9023
rect 13650 8974 13810 8977
rect 13862 8974 14021 8977
rect 14073 8974 14111 9026
rect 9089 8963 14111 8974
rect 9089 8940 12583 8963
rect 13301 8940 14111 8963
rect 9089 8488 9205 8940
rect 9812 8933 10120 8940
rect 10385 8926 12583 8940
rect 13350 8933 14111 8940
rect 14393 9060 14943 9067
rect 15181 9060 18143 9141
rect 23682 9147 23974 9265
rect 23682 9101 23820 9147
rect 23866 9101 23974 9147
rect 23682 9067 23974 9101
rect 18397 9060 19579 9067
rect 19905 9060 20456 9067
rect 14393 9026 19579 9060
rect 14393 9023 14431 9026
rect 14483 9023 14642 9026
rect 14694 9023 14853 9026
rect 14905 9023 18435 9026
rect 14393 8977 14409 9023
rect 14483 8977 14522 9023
rect 14568 8977 14635 9023
rect 14694 8977 14748 9023
rect 14794 8977 14853 9023
rect 14907 8977 15216 9023
rect 15262 8977 15374 9023
rect 15420 8977 15532 9023
rect 15578 8977 15690 9023
rect 15736 8977 15848 9023
rect 15894 8977 16006 9023
rect 16052 8977 16165 9023
rect 16211 8977 16323 9023
rect 16369 8977 16481 9023
rect 16527 8977 16639 9023
rect 16685 8977 16797 9023
rect 16843 8977 16955 9023
rect 17001 8977 17113 9023
rect 17159 8977 17272 9023
rect 17318 8977 17430 9023
rect 17476 8977 17588 9023
rect 17634 8977 17746 9023
rect 17792 8977 17904 9023
rect 17950 8977 18062 9023
rect 18108 8977 18435 9023
rect 14393 8974 14431 8977
rect 14483 8974 14642 8977
rect 14694 8974 14853 8977
rect 14905 8974 18435 8977
rect 18487 8974 18645 9026
rect 18697 8974 18856 9026
rect 18908 8974 19068 9026
rect 19120 8974 19279 9026
rect 19331 8974 19489 9026
rect 19541 8974 19579 9026
rect 14393 8940 19579 8974
rect 19904 9026 20456 9060
rect 19904 8974 19943 9026
rect 19995 9023 20154 9026
rect 20206 9023 20365 9026
rect 20417 9023 20456 9026
rect 21875 9026 23974 9067
rect 21875 9023 21913 9026
rect 21965 9023 22124 9026
rect 22176 9023 22335 9026
rect 22387 9023 22545 9026
rect 22597 9023 22756 9026
rect 22808 9023 22968 9026
rect 23020 9023 23179 9026
rect 23231 9023 23389 9026
rect 19995 8977 20064 9023
rect 20110 8977 20154 9023
rect 20214 8977 20271 9023
rect 20317 8977 20365 9023
rect 20420 8977 20477 9023
rect 20523 8977 20580 9023
rect 20626 8977 20683 9023
rect 20729 8977 20786 9023
rect 20832 8977 20889 9023
rect 20935 8977 20992 9023
rect 21038 8977 21051 9023
rect 21386 8977 21399 9023
rect 23373 8977 23389 9023
rect 19995 8974 20154 8977
rect 20206 8974 20365 8977
rect 20417 8974 20456 8977
rect 19904 8940 20456 8974
rect 14393 8933 14943 8940
rect 12959 8882 13121 8893
rect 9334 8799 9463 8828
rect 9843 8810 9959 8847
rect 12959 8836 12970 8882
rect 13110 8836 13121 8882
rect 12959 8829 13121 8836
rect 9324 8753 9337 8799
rect 9383 8788 9459 8799
rect 9424 8753 9459 8788
rect 9505 8753 9582 8799
rect 9628 8753 9705 8799
rect 9751 8753 9764 8799
rect 9843 8764 9878 8810
rect 9924 8764 9959 8810
rect 9334 8736 9372 8753
rect 9424 8736 9463 8753
rect 9334 8709 9463 8736
rect 9334 8696 9462 8709
rect 9520 8573 9682 8613
rect 9520 8521 9591 8573
rect 9643 8521 9682 8573
rect 8605 8442 8618 8488
rect 8664 8442 8741 8488
rect 8787 8442 8864 8488
rect 8910 8442 8923 8488
rect 9089 8442 9238 8488
rect 9284 8442 9327 8488
rect 8611 8410 8920 8442
rect 9089 8410 9205 8442
rect 7450 8298 7758 8303
rect 6035 8264 6550 8298
rect 7036 8264 7758 8298
rect 8255 8278 8323 8400
rect 9520 8390 9682 8521
rect 9406 8387 9682 8390
rect 9406 8379 9591 8387
rect 9406 8333 9441 8379
rect 9487 8335 9591 8379
rect 9643 8366 9682 8387
rect 9843 8366 9959 8764
rect 10315 8788 13121 8829
rect 15181 8859 18143 8940
rect 18397 8933 19579 8940
rect 19905 8933 20456 8940
rect 21875 8974 21913 8977
rect 21965 8974 22124 8977
rect 22176 8974 22335 8977
rect 22387 8974 22545 8977
rect 22597 8974 22756 8977
rect 22808 8974 22968 8977
rect 23020 8974 23179 8977
rect 23231 8974 23389 8977
rect 23441 8974 23600 9026
rect 23652 8974 23811 9026
rect 23863 8974 23974 9026
rect 21875 8933 23974 8974
rect 15181 8813 15216 8859
rect 15262 8813 15374 8859
rect 15420 8813 15532 8859
rect 15578 8813 15690 8859
rect 15736 8813 15848 8859
rect 15894 8813 16006 8859
rect 16052 8813 16165 8859
rect 16211 8813 16323 8859
rect 16369 8813 16481 8859
rect 16527 8813 16639 8859
rect 16685 8813 16797 8859
rect 16843 8813 16955 8859
rect 17001 8813 17113 8859
rect 17159 8813 17272 8859
rect 17318 8813 17430 8859
rect 17476 8813 17588 8859
rect 17634 8813 17746 8859
rect 17792 8813 17904 8859
rect 17950 8813 18062 8859
rect 18108 8813 18143 8859
rect 23682 8899 23974 8933
rect 23682 8853 23820 8899
rect 23866 8853 23974 8899
rect 10315 8736 11532 8788
rect 11584 8736 13121 8788
rect 10315 8695 13121 8736
rect 14202 8753 14409 8799
rect 14455 8753 14522 8799
rect 14568 8753 14635 8799
rect 14681 8753 14748 8799
rect 14794 8753 14861 8799
rect 14907 8753 14920 8799
rect 15181 8777 18143 8813
rect 20632 8802 20940 8843
rect 20632 8799 20670 8802
rect 20722 8799 20850 8802
rect 20902 8799 20940 8802
rect 21186 8827 21254 8838
rect 13938 8687 14106 8698
rect 13938 8641 13955 8687
rect 14095 8641 14106 8687
rect 13938 8597 14106 8641
rect 11826 8557 14106 8597
rect 11826 8505 12665 8557
rect 12717 8505 14106 8557
rect 11826 8464 14106 8505
rect 14202 8366 14318 8753
rect 18502 8727 19474 8767
rect 20051 8753 20064 8799
rect 20110 8753 20168 8799
rect 20214 8753 20271 8799
rect 20317 8753 20374 8799
rect 20420 8753 20477 8799
rect 20523 8753 20580 8799
rect 20626 8753 20670 8799
rect 20729 8753 20786 8799
rect 20832 8753 20850 8799
rect 20935 8753 20992 8799
rect 21038 8753 21051 8799
rect 18502 8712 18540 8727
rect 18592 8712 18751 8727
rect 18803 8712 18962 8727
rect 19014 8712 19173 8727
rect 19225 8712 19384 8727
rect 19436 8712 19474 8727
rect 18362 8666 18375 8712
rect 18421 8666 18478 8712
rect 18524 8675 18540 8712
rect 18524 8666 18581 8675
rect 18627 8666 18684 8712
rect 18730 8675 18751 8712
rect 18730 8666 18787 8675
rect 18833 8666 18890 8712
rect 18936 8675 18962 8712
rect 18936 8666 18993 8675
rect 19039 8666 19096 8712
rect 19142 8675 19173 8712
rect 19142 8666 19199 8675
rect 19449 8666 19474 8712
rect 20632 8750 20670 8753
rect 20722 8750 20850 8753
rect 20902 8750 20940 8753
rect 20632 8710 20940 8750
rect 18154 8620 18284 8661
rect 18502 8635 19474 8666
rect 14498 8575 14838 8604
rect 14396 8529 14409 8575
rect 14455 8529 14522 8575
rect 14568 8564 14635 8575
rect 14588 8529 14635 8564
rect 14681 8529 14748 8575
rect 14794 8564 14861 8575
rect 14800 8529 14861 8564
rect 14907 8529 14920 8575
rect 18154 8568 18193 8620
rect 18245 8568 18284 8620
rect 18154 8565 18284 8568
rect 14498 8512 14536 8529
rect 14588 8512 14748 8529
rect 14800 8512 14838 8529
rect 14498 8471 14838 8512
rect 14997 8456 17976 8489
rect 14997 8410 15061 8456
rect 15201 8448 17976 8456
rect 15201 8410 17461 8448
rect 14997 8396 17461 8410
rect 17513 8396 17976 8448
rect 9643 8351 14515 8366
rect 14997 8355 17976 8396
rect 18154 8425 18219 8565
rect 18265 8425 18284 8565
rect 19859 8575 20409 8604
rect 19859 8564 20064 8575
rect 20110 8564 20168 8575
rect 19417 8488 19757 8529
rect 18362 8442 18375 8488
rect 18421 8442 18478 8488
rect 18524 8442 18581 8488
rect 18627 8442 18684 8488
rect 18730 8442 18787 8488
rect 18833 8442 18890 8488
rect 18936 8442 18993 8488
rect 19039 8442 19096 8488
rect 19142 8442 19199 8488
rect 19449 8442 19757 8488
rect 19859 8512 19897 8564
rect 19949 8529 20064 8564
rect 20160 8529 20168 8564
rect 20214 8529 20271 8575
rect 20317 8564 20374 8575
rect 20317 8529 20319 8564
rect 19949 8512 20108 8529
rect 20160 8512 20319 8529
rect 20371 8529 20374 8564
rect 20420 8529 20477 8575
rect 20523 8529 20580 8575
rect 20626 8529 20683 8575
rect 20729 8529 20786 8575
rect 20832 8529 20889 8575
rect 20935 8529 20992 8575
rect 21038 8529 21051 8575
rect 20371 8512 20409 8529
rect 19859 8471 20409 8512
rect 18154 8402 18284 8425
rect 19417 8410 19757 8442
rect 9643 8335 14409 8351
rect 9487 8333 14409 8335
rect 9406 8330 14409 8333
rect 9406 8284 13336 8330
rect 13382 8284 13503 8330
rect 13549 8284 13668 8330
rect 13714 8284 13833 8330
rect 13879 8305 14409 8330
rect 14455 8305 14522 8351
rect 14568 8305 14635 8351
rect 14681 8305 14748 8351
rect 14794 8305 14861 8351
rect 14907 8305 14920 8351
rect 18154 8350 18193 8402
rect 18245 8350 18284 8402
rect 18154 8310 18284 8350
rect 19641 8353 19757 8410
rect 21186 8405 21197 8827
rect 21243 8405 21254 8827
rect 21394 8799 21702 8836
rect 21386 8753 21399 8799
rect 23373 8753 23386 8799
rect 21394 8743 21432 8753
rect 21484 8743 21612 8753
rect 21664 8743 21702 8753
rect 21394 8703 21702 8743
rect 23682 8735 23974 8853
rect 23682 8689 23820 8735
rect 23866 8689 23974 8735
rect 23682 8597 23974 8689
rect 23182 8575 23974 8597
rect 21386 8529 21399 8575
rect 23373 8529 23974 8575
rect 23182 8478 23974 8529
rect 21186 8353 21254 8405
rect 19641 8316 21254 8353
rect 21394 8351 21702 8373
rect 13879 8284 14515 8305
rect 8255 8264 9320 8278
rect 345 8200 452 8246
rect 498 8200 637 8246
rect 3081 8233 4240 8262
rect 4857 8218 4870 8264
rect 5120 8218 5140 8264
rect 5223 8218 5280 8264
rect 5326 8218 5351 8264
rect 5429 8218 5486 8264
rect 5532 8218 5562 8264
rect 5635 8218 5692 8264
rect 5738 8218 5773 8264
rect 5841 8218 5898 8264
rect 5944 8218 5957 8264
rect 6035 8218 6451 8264
rect 6497 8218 6568 8264
rect 6614 8218 6685 8264
rect 6731 8218 6803 8264
rect 6849 8218 6921 8264
rect 6967 8218 7039 8264
rect 7085 8262 7506 8264
rect 7085 8218 7488 8262
rect 7552 8218 7623 8264
rect 7669 8262 7740 8264
rect 7720 8218 7740 8262
rect 7786 8218 7858 8264
rect 7904 8218 7976 8264
rect 8022 8218 8094 8264
rect 8140 8218 8153 8264
rect 8255 8218 8618 8264
rect 8664 8218 8741 8264
rect 8787 8218 8864 8264
rect 8910 8218 9238 8264
rect 9284 8218 9327 8264
rect 9406 8246 14515 8284
rect 18502 8264 19474 8304
rect 18362 8218 18375 8264
rect 18421 8218 18478 8264
rect 18524 8218 18540 8264
rect 18627 8218 18684 8264
rect 18730 8218 18751 8264
rect 18833 8218 18890 8264
rect 18936 8218 18962 8264
rect 19039 8218 19096 8264
rect 19142 8218 19173 8264
rect 19449 8218 19474 8264
rect 19641 8270 20113 8316
rect 20159 8270 20300 8316
rect 20346 8270 20487 8316
rect 20533 8270 20673 8316
rect 20719 8270 20860 8316
rect 20906 8270 21254 8316
rect 21386 8305 21399 8351
rect 23373 8305 23386 8351
rect 19641 8260 21254 8270
rect 20078 8233 21254 8260
rect 21394 8280 21432 8305
rect 21484 8280 21612 8305
rect 21664 8280 21702 8305
rect 21394 8240 21702 8280
rect 23682 8246 23974 8478
rect 345 8167 637 8200
rect 4891 8212 4929 8218
rect 4981 8212 5140 8218
rect 5192 8212 5351 8218
rect 5403 8212 5562 8218
rect 5614 8212 5773 8218
rect 5825 8212 5863 8218
rect 4467 8167 4622 8174
rect 4891 8172 5863 8212
rect 6035 8178 6550 8218
rect 7036 8210 7488 8218
rect 7540 8210 7668 8218
rect 7720 8210 7758 8218
rect 7036 8178 7758 8210
rect 7450 8170 7758 8178
rect 345 8126 2439 8167
rect 345 8074 451 8126
rect 503 8074 662 8126
rect 714 8074 873 8126
rect 925 8074 1083 8126
rect 1135 8074 1294 8126
rect 1346 8074 1506 8126
rect 1558 8074 1717 8126
rect 1769 8074 1927 8126
rect 1979 8074 2138 8126
rect 2190 8074 2349 8126
rect 2401 8074 2439 8126
rect 345 8033 2439 8074
rect 4314 8126 4622 8167
rect 8255 8158 9320 8218
rect 18502 8212 18540 8218
rect 18592 8212 18751 8218
rect 18803 8212 18962 8218
rect 19014 8212 19173 8218
rect 19225 8212 19384 8218
rect 19436 8212 19474 8218
rect 18502 8172 19474 8212
rect 23682 8200 23820 8246
rect 23866 8200 23974 8246
rect 19696 8167 19852 8174
rect 23682 8167 23974 8200
rect 4314 8074 4352 8126
rect 4404 8123 4532 8126
rect 4404 8077 4513 8123
rect 4404 8074 4532 8077
rect 4584 8074 4622 8126
rect 4314 8033 4622 8074
rect 19696 8126 20005 8167
rect 19696 8074 19735 8126
rect 19787 8123 19915 8126
rect 19803 8077 19915 8123
rect 19787 8074 19915 8077
rect 19967 8074 20005 8126
rect 345 8000 637 8033
rect 4467 8026 4622 8033
rect 345 7954 452 8000
rect 498 7954 637 8000
rect 4891 7988 5863 8028
rect 7450 8022 7758 8030
rect 4891 7982 4929 7988
rect 4981 7982 5140 7988
rect 5192 7982 5351 7988
rect 5403 7982 5562 7988
rect 5614 7982 5773 7988
rect 5825 7982 5863 7988
rect 6035 7982 6550 8022
rect 7036 7990 7758 8022
rect 7036 7982 7488 7990
rect 7540 7982 7668 7990
rect 7720 7982 7758 7990
rect 8255 7982 9320 8042
rect 19696 8033 20005 8074
rect 21875 8126 23974 8167
rect 21875 8074 21913 8126
rect 21965 8074 22124 8126
rect 22176 8074 22335 8126
rect 22387 8074 22545 8126
rect 22597 8074 22756 8126
rect 22808 8074 22968 8126
rect 23020 8074 23179 8126
rect 23231 8074 23389 8126
rect 23441 8074 23600 8126
rect 23652 8074 23811 8126
rect 23863 8074 23974 8126
rect 21875 8033 23974 8074
rect 18502 7988 19474 8028
rect 19696 8026 19852 8033
rect 18502 7982 18540 7988
rect 18592 7982 18751 7988
rect 18803 7982 18962 7988
rect 19014 7982 19173 7988
rect 19225 7982 19384 7988
rect 19436 7982 19474 7988
rect 345 7837 637 7954
rect 3081 7938 4240 7967
rect 2616 7898 2924 7938
rect 2616 7895 2654 7898
rect 2706 7895 2834 7898
rect 2886 7895 2924 7898
rect 3081 7930 4679 7938
rect 4857 7936 4870 7982
rect 5120 7936 5140 7982
rect 5223 7936 5280 7982
rect 5326 7936 5351 7982
rect 5429 7936 5486 7982
rect 5532 7936 5562 7982
rect 5635 7936 5692 7982
rect 5738 7936 5773 7982
rect 5841 7936 5898 7982
rect 5944 7936 5957 7982
rect 6035 7936 6451 7982
rect 6497 7936 6568 7982
rect 6614 7936 6685 7982
rect 6731 7936 6803 7982
rect 6849 7936 6921 7982
rect 6967 7936 7039 7982
rect 7085 7938 7488 7982
rect 7085 7936 7506 7938
rect 7552 7936 7623 7982
rect 7720 7938 7740 7982
rect 7669 7936 7740 7938
rect 7786 7936 7858 7982
rect 7904 7936 7976 7982
rect 8022 7936 8094 7982
rect 8140 7936 8153 7982
rect 8255 7936 8618 7982
rect 8664 7936 8741 7982
rect 8787 7936 8864 7982
rect 8910 7936 9238 7982
rect 9284 7936 9327 7982
rect 933 7849 946 7895
rect 2920 7849 2933 7895
rect 3081 7884 3413 7930
rect 3459 7884 3599 7930
rect 3645 7884 3786 7930
rect 3832 7884 3973 7930
rect 4019 7884 4159 7930
rect 4205 7884 4679 7930
rect 4891 7896 5863 7936
rect 6035 7902 6550 7936
rect 7036 7902 7758 7936
rect 345 7791 452 7837
rect 498 7791 637 7837
rect 2616 7846 2654 7849
rect 2706 7846 2834 7849
rect 2886 7846 2924 7849
rect 2616 7805 2924 7846
rect 3081 7847 4679 7884
rect 345 7722 637 7791
rect 3081 7765 3149 7847
rect 345 7674 1090 7722
rect 345 7628 452 7674
rect 498 7671 1090 7674
rect 498 7628 946 7671
rect 345 7625 946 7628
rect 2920 7625 2933 7671
rect 345 7603 1090 7625
rect 345 7511 637 7603
rect 345 7465 452 7511
rect 498 7465 637 7511
rect 345 7347 637 7465
rect 2616 7450 2924 7490
rect 2616 7447 2654 7450
rect 2706 7447 2834 7450
rect 2886 7447 2924 7450
rect 933 7401 946 7447
rect 2920 7401 2933 7447
rect 2616 7398 2654 7401
rect 2706 7398 2834 7401
rect 2886 7398 2924 7401
rect 2616 7357 2924 7398
rect 345 7301 452 7347
rect 498 7301 637 7347
rect 3081 7343 3092 7765
rect 3138 7343 3149 7765
rect 4561 7790 4679 7847
rect 6035 7802 6151 7902
rect 7450 7897 7758 7902
rect 8255 7922 9320 7936
rect 4561 7758 5957 7790
rect 3825 7688 4315 7729
rect 3825 7671 3864 7688
rect 3916 7671 4044 7688
rect 4096 7671 4224 7688
rect 3268 7625 3281 7671
rect 3327 7625 3384 7671
rect 3430 7625 3487 7671
rect 3533 7625 3590 7671
rect 3636 7625 3693 7671
rect 3739 7625 3796 7671
rect 3842 7636 3864 7671
rect 3842 7625 3899 7636
rect 3945 7625 4002 7671
rect 4096 7636 4105 7671
rect 4048 7625 4105 7636
rect 4151 7625 4209 7671
rect 4276 7636 4315 7688
rect 4561 7712 4870 7758
rect 5120 7712 5177 7758
rect 5223 7712 5280 7758
rect 5326 7712 5383 7758
rect 5429 7712 5486 7758
rect 5532 7712 5589 7758
rect 5635 7712 5692 7758
rect 5738 7712 5795 7758
rect 5841 7712 5898 7758
rect 5944 7712 5957 7758
rect 4561 7668 5957 7712
rect 4255 7625 4315 7636
rect 3825 7596 4315 7625
rect 6035 7662 6072 7802
rect 6118 7662 6151 7802
rect 4891 7534 5863 7568
rect 6035 7559 6151 7662
rect 6237 7802 6370 7822
rect 6237 7763 6294 7802
rect 6237 7711 6275 7763
rect 6237 7662 6294 7711
rect 6340 7662 6370 7802
rect 8255 7800 8323 7922
rect 9406 7916 14515 7954
rect 18362 7936 18375 7982
rect 18421 7936 18478 7982
rect 18524 7936 18540 7982
rect 18627 7936 18684 7982
rect 18730 7936 18751 7982
rect 18833 7936 18890 7982
rect 18936 7936 18962 7982
rect 19039 7936 19096 7982
rect 19142 7936 19173 7982
rect 19449 7936 19474 7982
rect 23682 8000 23974 8033
rect 20078 7940 21254 7967
rect 9406 7870 13336 7916
rect 13382 7870 13503 7916
rect 13549 7870 13668 7916
rect 13714 7870 13833 7916
rect 13879 7895 14515 7916
rect 18502 7896 19474 7936
rect 19641 7930 21254 7940
rect 13879 7870 14409 7895
rect 9406 7867 14409 7870
rect 9406 7821 9441 7867
rect 9487 7865 14409 7867
rect 9487 7821 9591 7865
rect 9406 7813 9591 7821
rect 9643 7849 14409 7865
rect 14455 7849 14522 7895
rect 14568 7849 14635 7895
rect 14681 7849 14748 7895
rect 14794 7849 14861 7895
rect 14907 7849 14920 7895
rect 18154 7850 18284 7890
rect 9643 7834 14515 7849
rect 9643 7813 9682 7834
rect 9406 7810 9682 7813
rect 6521 7790 7282 7797
rect 6520 7758 7528 7790
rect 6438 7712 6451 7758
rect 6497 7756 6568 7758
rect 6497 7712 6558 7756
rect 6614 7712 6685 7758
rect 6731 7756 6803 7758
rect 6731 7712 6769 7756
rect 6849 7712 6921 7758
rect 6967 7756 7039 7758
rect 6967 7712 6981 7756
rect 6520 7704 6558 7712
rect 6610 7704 6769 7712
rect 6821 7704 6981 7712
rect 7033 7712 7039 7756
rect 7085 7756 7506 7758
rect 7085 7712 7192 7756
rect 7033 7704 7192 7712
rect 7244 7712 7506 7756
rect 7552 7712 7623 7758
rect 7669 7712 7740 7758
rect 7786 7712 7858 7758
rect 7904 7712 7976 7758
rect 8022 7712 8094 7758
rect 8140 7712 8153 7758
rect 7244 7704 7528 7712
rect 6520 7671 7528 7704
rect 6520 7670 7282 7671
rect 6521 7664 7282 7670
rect 6237 7639 6370 7662
rect 8255 7660 8266 7800
rect 8312 7660 8323 7800
rect 8611 7758 8920 7790
rect 9089 7758 9205 7790
rect 8605 7712 8618 7758
rect 8664 7712 8741 7758
rect 8787 7712 8864 7758
rect 8910 7712 8923 7758
rect 9089 7712 9238 7758
rect 9284 7712 9327 7758
rect 8255 7649 8323 7660
rect 6035 7534 6550 7559
rect 7036 7556 7528 7559
rect 7036 7534 7758 7556
rect 4857 7488 4870 7534
rect 5120 7528 5177 7534
rect 5120 7488 5140 7528
rect 5223 7488 5280 7534
rect 5326 7528 5383 7534
rect 5326 7488 5351 7528
rect 5429 7488 5486 7534
rect 5532 7528 5589 7534
rect 5532 7488 5562 7528
rect 5635 7488 5692 7534
rect 5738 7528 5795 7534
rect 5738 7488 5773 7528
rect 5841 7488 5898 7534
rect 5944 7488 5957 7534
rect 6035 7488 6451 7534
rect 6497 7488 6568 7534
rect 6614 7488 6685 7534
rect 6731 7488 6803 7534
rect 6849 7488 6921 7534
rect 6967 7488 7039 7534
rect 7085 7516 7506 7534
rect 7085 7488 7488 7516
rect 7552 7488 7623 7534
rect 7669 7516 7740 7534
rect 7720 7488 7740 7516
rect 7786 7488 7858 7534
rect 7904 7488 7976 7534
rect 8022 7488 8094 7534
rect 8140 7488 8153 7534
rect 3378 7447 3686 7482
rect 4891 7476 4929 7488
rect 4981 7476 5140 7488
rect 5192 7476 5351 7488
rect 5403 7476 5562 7488
rect 5614 7476 5773 7488
rect 5825 7476 5863 7488
rect 3268 7401 3281 7447
rect 3327 7401 3384 7447
rect 3430 7442 3487 7447
rect 3468 7401 3487 7442
rect 3533 7401 3590 7447
rect 3636 7442 3693 7447
rect 3648 7401 3693 7442
rect 3739 7401 3796 7447
rect 3842 7401 3899 7447
rect 3945 7401 4002 7447
rect 4048 7401 4105 7447
rect 4151 7401 4209 7447
rect 4255 7401 4268 7447
rect 4891 7436 5863 7476
rect 6035 7439 6550 7488
rect 7036 7464 7488 7488
rect 7540 7464 7668 7488
rect 7720 7464 7758 7488
rect 7036 7439 7758 7464
rect 7450 7423 7758 7439
rect 3378 7390 3416 7401
rect 3468 7390 3596 7401
rect 3648 7390 3686 7401
rect 3378 7349 3686 7390
rect 3081 7332 3149 7343
rect 345 7267 637 7301
rect 345 7226 2439 7267
rect 3844 7260 4605 7267
rect 345 7174 451 7226
rect 503 7174 662 7226
rect 714 7174 873 7226
rect 925 7223 1083 7226
rect 1135 7223 1294 7226
rect 1346 7223 1506 7226
rect 1558 7223 1717 7226
rect 1769 7223 1927 7226
rect 1979 7223 2138 7226
rect 2190 7223 2349 7226
rect 2401 7223 2439 7226
rect 3843 7226 4605 7260
rect 3843 7223 3881 7226
rect 3933 7223 4092 7226
rect 4144 7223 4304 7226
rect 925 7177 946 7223
rect 2920 7177 2933 7223
rect 3268 7177 3281 7223
rect 3327 7177 3384 7223
rect 3430 7177 3487 7223
rect 3533 7177 3590 7223
rect 3636 7177 3693 7223
rect 3739 7177 3796 7223
rect 3842 7177 3881 7223
rect 3945 7177 4002 7223
rect 4048 7177 4092 7223
rect 4151 7177 4209 7223
rect 4255 7177 4304 7223
rect 925 7174 1083 7177
rect 1135 7174 1294 7177
rect 1346 7174 1506 7177
rect 1558 7174 1717 7177
rect 1769 7174 1927 7177
rect 1979 7174 2138 7177
rect 2190 7174 2349 7177
rect 2401 7174 2439 7177
rect 345 7133 2439 7174
rect 3843 7174 3881 7177
rect 3933 7174 4092 7177
rect 4144 7174 4304 7177
rect 4356 7174 4515 7226
rect 4567 7174 4605 7226
rect 3843 7140 4605 7174
rect 3844 7133 4605 7140
rect 4779 7260 5961 7267
rect 4779 7226 6555 7260
rect 4779 7174 4817 7226
rect 4869 7174 5027 7226
rect 5079 7174 5238 7226
rect 5290 7174 5450 7226
rect 5502 7174 5661 7226
rect 5713 7174 5871 7226
rect 5923 7223 6555 7226
rect 5923 7177 6086 7223
rect 6320 7177 6555 7223
rect 5923 7174 6555 7177
rect 4779 7140 6555 7174
rect 7543 7226 8439 7267
rect 7543 7223 7927 7226
rect 7979 7223 8138 7226
rect 7543 7177 7554 7223
rect 8070 7177 8138 7223
rect 7543 7174 7927 7177
rect 7979 7174 8138 7177
rect 8190 7174 8349 7226
rect 8401 7174 8439 7226
rect 4779 7133 5961 7140
rect 7543 7133 8439 7174
rect 8611 7226 8920 7712
rect 8611 7174 8649 7226
rect 8701 7223 8829 7226
rect 8705 7177 8817 7223
rect 8701 7174 8829 7177
rect 8881 7174 8920 7226
rect 345 7099 637 7133
rect 345 7053 452 7099
rect 498 7053 637 7099
rect 345 6935 637 7053
rect 3081 7057 3149 7068
rect 2616 7002 2924 7043
rect 2616 6999 2654 7002
rect 2706 6999 2834 7002
rect 2886 6999 2924 7002
rect 933 6953 946 6999
rect 2920 6953 2933 6999
rect 345 6889 452 6935
rect 498 6889 637 6935
rect 2616 6950 2654 6953
rect 2706 6950 2834 6953
rect 2886 6950 2924 6953
rect 2616 6910 2924 6950
rect 345 6797 637 6889
rect 345 6775 1090 6797
rect 345 6772 946 6775
rect 345 6726 452 6772
rect 498 6729 946 6772
rect 2920 6729 2933 6775
rect 498 6726 1090 6729
rect 345 6678 1090 6726
rect 345 6609 637 6678
rect 345 6563 452 6609
rect 498 6563 637 6609
rect 3081 6635 3092 7057
rect 3138 6635 3149 7057
rect 3378 7010 3686 7051
rect 3378 6999 3416 7010
rect 3468 6999 3596 7010
rect 3648 6999 3686 7010
rect 3268 6953 3281 6999
rect 3327 6953 3384 6999
rect 3468 6958 3487 6999
rect 3430 6953 3487 6958
rect 3533 6953 3590 6999
rect 3648 6958 3693 6999
rect 3636 6953 3693 6958
rect 3739 6953 3796 6999
rect 3842 6953 3899 6999
rect 3945 6953 4002 6999
rect 4048 6953 4105 6999
rect 4151 6953 4209 6999
rect 4255 6953 4268 6999
rect 3378 6918 3686 6953
rect 4891 6924 5863 6964
rect 7450 6961 7758 6977
rect 4891 6912 4929 6924
rect 4981 6912 5140 6924
rect 5192 6912 5351 6924
rect 5403 6912 5562 6924
rect 5614 6912 5773 6924
rect 5825 6912 5863 6924
rect 6035 6912 6550 6961
rect 7036 6936 7758 6961
rect 7036 6912 7488 6936
rect 7540 6912 7668 6936
rect 7720 6912 7758 6936
rect 4857 6866 4870 6912
rect 5120 6872 5140 6912
rect 5120 6866 5177 6872
rect 5223 6866 5280 6912
rect 5326 6872 5351 6912
rect 5326 6866 5383 6872
rect 5429 6866 5486 6912
rect 5532 6872 5562 6912
rect 5532 6866 5589 6872
rect 5635 6866 5692 6912
rect 5738 6872 5773 6912
rect 5738 6866 5795 6872
rect 5841 6866 5898 6912
rect 5944 6866 5957 6912
rect 6035 6866 6451 6912
rect 6497 6866 6568 6912
rect 6614 6866 6685 6912
rect 6731 6866 6803 6912
rect 6849 6866 6921 6912
rect 6967 6866 7039 6912
rect 7085 6884 7488 6912
rect 7085 6866 7506 6884
rect 7552 6866 7623 6912
rect 7720 6884 7740 6912
rect 7669 6866 7740 6884
rect 7786 6866 7858 6912
rect 7904 6866 7976 6912
rect 8022 6866 8094 6912
rect 8140 6866 8153 6912
rect 4891 6832 5863 6866
rect 6035 6841 6550 6866
rect 7036 6844 7758 6866
rect 7036 6841 7528 6844
rect 3825 6775 4315 6804
rect 3268 6729 3281 6775
rect 3327 6729 3384 6775
rect 3430 6729 3487 6775
rect 3533 6729 3590 6775
rect 3636 6729 3693 6775
rect 3739 6729 3796 6775
rect 3842 6764 3899 6775
rect 3842 6729 3864 6764
rect 3945 6729 4002 6775
rect 4048 6764 4105 6775
rect 4096 6729 4105 6764
rect 4151 6729 4209 6775
rect 4255 6764 4315 6775
rect 3825 6712 3864 6729
rect 3916 6712 4044 6729
rect 4096 6712 4224 6729
rect 4276 6712 4315 6764
rect 6035 6738 6151 6841
rect 3825 6671 4315 6712
rect 4561 6688 5957 6732
rect 345 6446 637 6563
rect 2616 6554 2924 6595
rect 2616 6551 2654 6554
rect 2706 6551 2834 6554
rect 2886 6551 2924 6554
rect 3081 6553 3149 6635
rect 4561 6642 4870 6688
rect 5120 6642 5177 6688
rect 5223 6642 5280 6688
rect 5326 6642 5383 6688
rect 5429 6642 5486 6688
rect 5532 6642 5589 6688
rect 5635 6642 5692 6688
rect 5738 6642 5795 6688
rect 5841 6642 5898 6688
rect 5944 6642 5957 6688
rect 4561 6610 5957 6642
rect 4561 6553 4679 6610
rect 933 6505 946 6551
rect 2920 6505 2933 6551
rect 3081 6516 4679 6553
rect 2616 6502 2654 6505
rect 2706 6502 2834 6505
rect 2886 6502 2924 6505
rect 2616 6462 2924 6502
rect 3081 6470 3413 6516
rect 3459 6470 3599 6516
rect 3645 6470 3786 6516
rect 3832 6470 3973 6516
rect 4019 6470 4159 6516
rect 4205 6470 4679 6516
rect 6035 6598 6072 6738
rect 6118 6598 6151 6738
rect 3081 6462 4679 6470
rect 4891 6464 5863 6504
rect 6035 6498 6151 6598
rect 6237 6738 6370 6761
rect 6237 6689 6294 6738
rect 6237 6637 6275 6689
rect 6237 6598 6294 6637
rect 6340 6598 6370 6738
rect 8255 6740 8323 6751
rect 6521 6730 7282 6736
rect 6520 6729 7282 6730
rect 6520 6696 7528 6729
rect 6520 6688 6558 6696
rect 6610 6688 6769 6696
rect 6821 6688 6981 6696
rect 6438 6642 6451 6688
rect 6497 6644 6558 6688
rect 6497 6642 6568 6644
rect 6614 6642 6685 6688
rect 6731 6644 6769 6688
rect 6731 6642 6803 6644
rect 6849 6642 6921 6688
rect 6967 6644 6981 6688
rect 7033 6688 7192 6696
rect 7033 6644 7039 6688
rect 6967 6642 7039 6644
rect 7085 6644 7192 6688
rect 7244 6688 7528 6696
rect 7244 6644 7506 6688
rect 7085 6642 7506 6644
rect 7552 6642 7623 6688
rect 7669 6642 7740 6688
rect 7786 6642 7858 6688
rect 7904 6642 7976 6688
rect 8022 6642 8094 6688
rect 8140 6642 8153 6688
rect 6520 6610 7528 6642
rect 6521 6603 7282 6610
rect 6237 6578 6370 6598
rect 8255 6600 8266 6740
rect 8312 6600 8323 6740
rect 8611 6688 8920 7174
rect 9089 7260 9205 7712
rect 9520 7679 9682 7810
rect 9520 7627 9591 7679
rect 9643 7627 9682 7679
rect 9520 7587 9682 7627
rect 9334 7491 9462 7504
rect 9334 7464 9463 7491
rect 9334 7447 9372 7464
rect 9424 7447 9463 7464
rect 9324 7401 9337 7447
rect 9424 7412 9459 7447
rect 9383 7401 9459 7412
rect 9505 7401 9582 7447
rect 9628 7401 9705 7447
rect 9751 7401 9764 7447
rect 9843 7436 9959 7834
rect 11826 7695 14106 7736
rect 11826 7643 12665 7695
rect 12717 7643 14106 7695
rect 11826 7603 14106 7643
rect 13938 7559 14106 7603
rect 13938 7513 13955 7559
rect 14095 7513 14106 7559
rect 9334 7372 9463 7401
rect 9843 7390 9878 7436
rect 9924 7390 9959 7436
rect 9843 7353 9959 7390
rect 10315 7464 13121 7505
rect 13938 7502 14106 7513
rect 10315 7412 11532 7464
rect 11584 7412 13121 7464
rect 10315 7371 13121 7412
rect 14202 7447 14318 7834
rect 14997 7804 17976 7845
rect 14997 7790 17838 7804
rect 14997 7744 15061 7790
rect 15201 7752 17838 7790
rect 17890 7752 17976 7804
rect 15201 7744 17976 7752
rect 14498 7688 14838 7729
rect 14997 7711 17976 7744
rect 18154 7798 18193 7850
rect 18245 7798 18284 7850
rect 18154 7775 18284 7798
rect 19641 7884 20113 7930
rect 20159 7884 20300 7930
rect 20346 7884 20487 7930
rect 20533 7884 20673 7930
rect 20719 7884 20860 7930
rect 20906 7884 21254 7930
rect 21394 7920 21702 7960
rect 21394 7895 21432 7920
rect 21484 7895 21612 7920
rect 21664 7895 21702 7920
rect 23682 7954 23820 8000
rect 23866 7954 23974 8000
rect 19641 7847 21254 7884
rect 21386 7849 21399 7895
rect 23373 7849 23386 7895
rect 19641 7790 19757 7847
rect 14498 7671 14536 7688
rect 14588 7671 14748 7688
rect 14800 7671 14838 7688
rect 14396 7625 14409 7671
rect 14455 7625 14522 7671
rect 14588 7636 14635 7671
rect 14568 7625 14635 7636
rect 14681 7625 14748 7671
rect 14800 7636 14861 7671
rect 14794 7625 14861 7636
rect 14907 7625 14920 7671
rect 18154 7635 18219 7775
rect 18265 7635 18284 7775
rect 19417 7758 19757 7790
rect 18362 7712 18375 7758
rect 18421 7712 18478 7758
rect 18524 7712 18581 7758
rect 18627 7712 18684 7758
rect 18730 7712 18787 7758
rect 18833 7712 18890 7758
rect 18936 7712 18993 7758
rect 19039 7712 19096 7758
rect 19142 7712 19199 7758
rect 19449 7712 19757 7758
rect 21186 7795 21254 7847
rect 21394 7827 21702 7849
rect 19417 7671 19757 7712
rect 19859 7688 20409 7729
rect 18154 7632 18284 7635
rect 14498 7596 14838 7625
rect 18154 7580 18193 7632
rect 18245 7580 18284 7632
rect 19859 7636 19897 7688
rect 19949 7671 20108 7688
rect 20160 7671 20319 7688
rect 19949 7636 20064 7671
rect 20160 7636 20168 7671
rect 19859 7625 20064 7636
rect 20110 7625 20168 7636
rect 20214 7625 20271 7671
rect 20317 7636 20319 7671
rect 20371 7671 20409 7688
rect 20371 7636 20374 7671
rect 20317 7625 20374 7636
rect 20420 7625 20477 7671
rect 20523 7625 20580 7671
rect 20626 7625 20683 7671
rect 20729 7625 20786 7671
rect 20832 7625 20889 7671
rect 20935 7625 20992 7671
rect 21038 7625 21051 7671
rect 19859 7596 20409 7625
rect 18154 7539 18284 7580
rect 18502 7534 19474 7565
rect 18362 7488 18375 7534
rect 18421 7488 18478 7534
rect 18524 7525 18581 7534
rect 18524 7488 18540 7525
rect 18627 7488 18684 7534
rect 18730 7525 18787 7534
rect 18730 7488 18751 7525
rect 18833 7488 18890 7534
rect 18936 7525 18993 7534
rect 18936 7488 18962 7525
rect 19039 7488 19096 7534
rect 19142 7525 19199 7534
rect 19142 7488 19173 7525
rect 19449 7488 19474 7534
rect 18502 7473 18540 7488
rect 18592 7473 18751 7488
rect 18803 7473 18962 7488
rect 19014 7473 19173 7488
rect 19225 7473 19384 7488
rect 19436 7473 19474 7488
rect 14202 7401 14409 7447
rect 14455 7401 14522 7447
rect 14568 7401 14635 7447
rect 14681 7401 14748 7447
rect 14794 7401 14861 7447
rect 14907 7401 14920 7447
rect 18502 7433 19474 7473
rect 20632 7450 20940 7490
rect 20632 7447 20670 7450
rect 20722 7447 20850 7450
rect 20902 7447 20940 7450
rect 12959 7364 13121 7371
rect 12959 7318 12970 7364
rect 13110 7318 13121 7364
rect 12959 7307 13121 7318
rect 15181 7387 18143 7423
rect 20051 7401 20064 7447
rect 20110 7401 20168 7447
rect 20214 7401 20271 7447
rect 20317 7401 20374 7447
rect 20420 7401 20477 7447
rect 20523 7401 20580 7447
rect 20626 7401 20670 7447
rect 20729 7401 20786 7447
rect 20832 7401 20850 7447
rect 20935 7401 20992 7447
rect 21038 7401 21051 7447
rect 15181 7341 15216 7387
rect 15262 7341 15374 7387
rect 15420 7341 15532 7387
rect 15578 7341 15690 7387
rect 15736 7341 15848 7387
rect 15894 7341 16006 7387
rect 16052 7341 16165 7387
rect 16211 7341 16323 7387
rect 16369 7341 16481 7387
rect 16527 7341 16639 7387
rect 16685 7341 16797 7387
rect 16843 7341 16955 7387
rect 17001 7341 17113 7387
rect 17159 7341 17272 7387
rect 17318 7341 17430 7387
rect 17476 7341 17588 7387
rect 17634 7341 17746 7387
rect 17792 7341 17904 7387
rect 17950 7341 18062 7387
rect 18108 7341 18143 7387
rect 20632 7398 20670 7401
rect 20722 7398 20850 7401
rect 20902 7398 20940 7401
rect 20632 7357 20940 7398
rect 21186 7373 21197 7795
rect 21243 7373 21254 7795
rect 23682 7722 23974 7954
rect 23182 7671 23974 7722
rect 21386 7625 21399 7671
rect 23373 7625 23974 7671
rect 23182 7603 23974 7625
rect 23682 7511 23974 7603
rect 21394 7457 21702 7497
rect 21394 7447 21432 7457
rect 21484 7447 21612 7457
rect 21664 7447 21702 7457
rect 23682 7465 23820 7511
rect 23866 7465 23974 7511
rect 21386 7401 21399 7447
rect 23373 7401 23386 7447
rect 21186 7362 21254 7373
rect 21394 7364 21702 7401
rect 9812 7260 10120 7267
rect 10385 7260 12583 7274
rect 13350 7260 14111 7267
rect 9089 7237 12583 7260
rect 13301 7237 14111 7260
rect 9089 7226 14111 7237
rect 9089 7223 9850 7226
rect 9089 7177 9337 7223
rect 9383 7177 9459 7223
rect 9505 7177 9582 7223
rect 9628 7177 9705 7223
rect 9751 7177 9850 7223
rect 9089 7174 9850 7177
rect 9902 7174 10030 7226
rect 10082 7223 13387 7226
rect 10082 7177 10433 7223
rect 10479 7177 10591 7223
rect 10637 7177 10749 7223
rect 10795 7177 10907 7223
rect 10953 7177 11066 7223
rect 11112 7177 11224 7223
rect 11270 7177 11382 7223
rect 11428 7177 11540 7223
rect 11586 7177 11698 7223
rect 11744 7177 11856 7223
rect 11902 7177 12015 7223
rect 12061 7177 12173 7223
rect 12219 7177 12331 7223
rect 12377 7177 12489 7223
rect 12535 7177 13336 7223
rect 13382 7177 13387 7223
rect 10082 7174 13387 7177
rect 13439 7223 13598 7226
rect 13439 7177 13503 7223
rect 13549 7177 13598 7223
rect 13439 7174 13598 7177
rect 13650 7223 13810 7226
rect 13862 7223 14021 7226
rect 13650 7177 13668 7223
rect 13714 7177 13810 7223
rect 13879 7177 14021 7223
rect 13650 7174 13810 7177
rect 13862 7174 14021 7177
rect 14073 7174 14111 7226
rect 9089 7163 14111 7174
rect 9089 7140 12583 7163
rect 13301 7140 14111 7163
rect 9089 6688 9205 7140
rect 9812 7133 10120 7140
rect 10385 7126 12583 7140
rect 13350 7133 14111 7140
rect 14393 7260 14943 7267
rect 15181 7260 18143 7341
rect 23682 7347 23974 7465
rect 23682 7301 23820 7347
rect 23866 7301 23974 7347
rect 23682 7267 23974 7301
rect 18397 7260 19579 7267
rect 19905 7260 20456 7267
rect 14393 7226 19579 7260
rect 14393 7223 14431 7226
rect 14483 7223 14642 7226
rect 14694 7223 14853 7226
rect 14905 7223 18435 7226
rect 14393 7177 14409 7223
rect 14483 7177 14522 7223
rect 14568 7177 14635 7223
rect 14694 7177 14748 7223
rect 14794 7177 14853 7223
rect 14907 7177 15216 7223
rect 15262 7177 15374 7223
rect 15420 7177 15532 7223
rect 15578 7177 15690 7223
rect 15736 7177 15848 7223
rect 15894 7177 16006 7223
rect 16052 7177 16165 7223
rect 16211 7177 16323 7223
rect 16369 7177 16481 7223
rect 16527 7177 16639 7223
rect 16685 7177 16797 7223
rect 16843 7177 16955 7223
rect 17001 7177 17113 7223
rect 17159 7177 17272 7223
rect 17318 7177 17430 7223
rect 17476 7177 17588 7223
rect 17634 7177 17746 7223
rect 17792 7177 17904 7223
rect 17950 7177 18062 7223
rect 18108 7177 18435 7223
rect 14393 7174 14431 7177
rect 14483 7174 14642 7177
rect 14694 7174 14853 7177
rect 14905 7174 18435 7177
rect 18487 7174 18645 7226
rect 18697 7174 18856 7226
rect 18908 7174 19068 7226
rect 19120 7174 19279 7226
rect 19331 7174 19489 7226
rect 19541 7174 19579 7226
rect 14393 7140 19579 7174
rect 19904 7226 20456 7260
rect 19904 7174 19943 7226
rect 19995 7223 20154 7226
rect 20206 7223 20365 7226
rect 20417 7223 20456 7226
rect 21875 7226 23974 7267
rect 21875 7223 21913 7226
rect 21965 7223 22124 7226
rect 22176 7223 22335 7226
rect 22387 7223 22545 7226
rect 22597 7223 22756 7226
rect 22808 7223 22968 7226
rect 23020 7223 23179 7226
rect 23231 7223 23389 7226
rect 19995 7177 20064 7223
rect 20110 7177 20154 7223
rect 20214 7177 20271 7223
rect 20317 7177 20365 7223
rect 20420 7177 20477 7223
rect 20523 7177 20580 7223
rect 20626 7177 20683 7223
rect 20729 7177 20786 7223
rect 20832 7177 20889 7223
rect 20935 7177 20992 7223
rect 21038 7177 21051 7223
rect 21386 7177 21399 7223
rect 23373 7177 23389 7223
rect 19995 7174 20154 7177
rect 20206 7174 20365 7177
rect 20417 7174 20456 7177
rect 19904 7140 20456 7174
rect 14393 7133 14943 7140
rect 12959 7082 13121 7093
rect 9334 6999 9463 7028
rect 9843 7010 9959 7047
rect 12959 7036 12970 7082
rect 13110 7036 13121 7082
rect 12959 7029 13121 7036
rect 9324 6953 9337 6999
rect 9383 6988 9459 6999
rect 9424 6953 9459 6988
rect 9505 6953 9582 6999
rect 9628 6953 9705 6999
rect 9751 6953 9764 6999
rect 9843 6964 9878 7010
rect 9924 6964 9959 7010
rect 9334 6936 9372 6953
rect 9424 6936 9463 6953
rect 9334 6909 9463 6936
rect 9334 6896 9462 6909
rect 9520 6773 9682 6813
rect 9520 6721 9591 6773
rect 9643 6721 9682 6773
rect 8605 6642 8618 6688
rect 8664 6642 8741 6688
rect 8787 6642 8864 6688
rect 8910 6642 8923 6688
rect 9089 6642 9238 6688
rect 9284 6642 9327 6688
rect 8611 6610 8920 6642
rect 9089 6610 9205 6642
rect 7450 6498 7758 6503
rect 6035 6464 6550 6498
rect 7036 6464 7758 6498
rect 8255 6478 8323 6600
rect 9520 6590 9682 6721
rect 9406 6587 9682 6590
rect 9406 6579 9591 6587
rect 9406 6533 9441 6579
rect 9487 6535 9591 6579
rect 9643 6566 9682 6587
rect 9843 6566 9959 6964
rect 10315 6988 13121 7029
rect 15181 7059 18143 7140
rect 18397 7133 19579 7140
rect 19905 7133 20456 7140
rect 21875 7174 21913 7177
rect 21965 7174 22124 7177
rect 22176 7174 22335 7177
rect 22387 7174 22545 7177
rect 22597 7174 22756 7177
rect 22808 7174 22968 7177
rect 23020 7174 23179 7177
rect 23231 7174 23389 7177
rect 23441 7174 23600 7226
rect 23652 7174 23811 7226
rect 23863 7174 23974 7226
rect 21875 7133 23974 7174
rect 15181 7013 15216 7059
rect 15262 7013 15374 7059
rect 15420 7013 15532 7059
rect 15578 7013 15690 7059
rect 15736 7013 15848 7059
rect 15894 7013 16006 7059
rect 16052 7013 16165 7059
rect 16211 7013 16323 7059
rect 16369 7013 16481 7059
rect 16527 7013 16639 7059
rect 16685 7013 16797 7059
rect 16843 7013 16955 7059
rect 17001 7013 17113 7059
rect 17159 7013 17272 7059
rect 17318 7013 17430 7059
rect 17476 7013 17588 7059
rect 17634 7013 17746 7059
rect 17792 7013 17904 7059
rect 17950 7013 18062 7059
rect 18108 7013 18143 7059
rect 23682 7099 23974 7133
rect 23682 7053 23820 7099
rect 23866 7053 23974 7099
rect 10315 6936 11532 6988
rect 11584 6936 13121 6988
rect 10315 6895 13121 6936
rect 14202 6953 14409 6999
rect 14455 6953 14522 6999
rect 14568 6953 14635 6999
rect 14681 6953 14748 6999
rect 14794 6953 14861 6999
rect 14907 6953 14920 6999
rect 15181 6977 18143 7013
rect 20632 7002 20940 7043
rect 20632 6999 20670 7002
rect 20722 6999 20850 7002
rect 20902 6999 20940 7002
rect 21186 7027 21254 7038
rect 13938 6887 14106 6898
rect 13938 6841 13955 6887
rect 14095 6841 14106 6887
rect 13938 6797 14106 6841
rect 11826 6757 14106 6797
rect 11826 6705 13042 6757
rect 13094 6705 14106 6757
rect 11826 6664 14106 6705
rect 14202 6566 14318 6953
rect 18502 6927 19474 6967
rect 20051 6953 20064 6999
rect 20110 6953 20168 6999
rect 20214 6953 20271 6999
rect 20317 6953 20374 6999
rect 20420 6953 20477 6999
rect 20523 6953 20580 6999
rect 20626 6953 20670 6999
rect 20729 6953 20786 6999
rect 20832 6953 20850 6999
rect 20935 6953 20992 6999
rect 21038 6953 21051 6999
rect 18502 6912 18540 6927
rect 18592 6912 18751 6927
rect 18803 6912 18962 6927
rect 19014 6912 19173 6927
rect 19225 6912 19384 6927
rect 19436 6912 19474 6927
rect 18362 6866 18375 6912
rect 18421 6866 18478 6912
rect 18524 6875 18540 6912
rect 18524 6866 18581 6875
rect 18627 6866 18684 6912
rect 18730 6875 18751 6912
rect 18730 6866 18787 6875
rect 18833 6866 18890 6912
rect 18936 6875 18962 6912
rect 18936 6866 18993 6875
rect 19039 6866 19096 6912
rect 19142 6875 19173 6912
rect 19142 6866 19199 6875
rect 19449 6866 19474 6912
rect 20632 6950 20670 6953
rect 20722 6950 20850 6953
rect 20902 6950 20940 6953
rect 20632 6910 20940 6950
rect 18154 6820 18284 6861
rect 18502 6835 19474 6866
rect 14498 6775 14838 6804
rect 14396 6729 14409 6775
rect 14455 6729 14522 6775
rect 14568 6764 14635 6775
rect 14588 6729 14635 6764
rect 14681 6729 14748 6775
rect 14794 6764 14861 6775
rect 14800 6729 14861 6764
rect 14907 6729 14920 6775
rect 18154 6768 18193 6820
rect 18245 6768 18284 6820
rect 18154 6765 18284 6768
rect 14498 6712 14536 6729
rect 14588 6712 14748 6729
rect 14800 6712 14838 6729
rect 14498 6671 14838 6712
rect 14997 6656 17976 6689
rect 14997 6610 15061 6656
rect 15201 6648 17976 6656
rect 14997 6596 15194 6610
rect 15246 6596 17976 6648
rect 9643 6551 14515 6566
rect 14997 6555 17976 6596
rect 18154 6625 18219 6765
rect 18265 6625 18284 6765
rect 19859 6775 20409 6804
rect 19859 6764 20064 6775
rect 20110 6764 20168 6775
rect 19417 6688 19757 6729
rect 18362 6642 18375 6688
rect 18421 6642 18478 6688
rect 18524 6642 18581 6688
rect 18627 6642 18684 6688
rect 18730 6642 18787 6688
rect 18833 6642 18890 6688
rect 18936 6642 18993 6688
rect 19039 6642 19096 6688
rect 19142 6642 19199 6688
rect 19449 6642 19757 6688
rect 19859 6712 19897 6764
rect 19949 6729 20064 6764
rect 20160 6729 20168 6764
rect 20214 6729 20271 6775
rect 20317 6764 20374 6775
rect 20317 6729 20319 6764
rect 19949 6712 20108 6729
rect 20160 6712 20319 6729
rect 20371 6729 20374 6764
rect 20420 6729 20477 6775
rect 20523 6729 20580 6775
rect 20626 6729 20683 6775
rect 20729 6729 20786 6775
rect 20832 6729 20889 6775
rect 20935 6729 20992 6775
rect 21038 6729 21051 6775
rect 20371 6712 20409 6729
rect 19859 6671 20409 6712
rect 18154 6602 18284 6625
rect 19417 6610 19757 6642
rect 9643 6535 14409 6551
rect 9487 6533 14409 6535
rect 9406 6530 14409 6533
rect 9406 6484 13336 6530
rect 13382 6484 13503 6530
rect 13549 6484 13668 6530
rect 13714 6484 13833 6530
rect 13879 6505 14409 6530
rect 14455 6505 14522 6551
rect 14568 6505 14635 6551
rect 14681 6505 14748 6551
rect 14794 6505 14861 6551
rect 14907 6505 14920 6551
rect 18154 6550 18193 6602
rect 18245 6550 18284 6602
rect 18154 6510 18284 6550
rect 19641 6553 19757 6610
rect 21186 6605 21197 7027
rect 21243 6605 21254 7027
rect 21394 6999 21702 7036
rect 21386 6953 21399 6999
rect 23373 6953 23386 6999
rect 21394 6943 21432 6953
rect 21484 6943 21612 6953
rect 21664 6943 21702 6953
rect 21394 6903 21702 6943
rect 23682 6935 23974 7053
rect 23682 6889 23820 6935
rect 23866 6889 23974 6935
rect 23682 6797 23974 6889
rect 23182 6775 23974 6797
rect 21386 6729 21399 6775
rect 23373 6729 23974 6775
rect 23182 6678 23974 6729
rect 21186 6553 21254 6605
rect 19641 6516 21254 6553
rect 21394 6551 21702 6573
rect 13879 6484 14515 6505
rect 8255 6464 9320 6478
rect 345 6400 452 6446
rect 498 6400 637 6446
rect 3081 6433 4240 6462
rect 4857 6418 4870 6464
rect 5120 6418 5140 6464
rect 5223 6418 5280 6464
rect 5326 6418 5351 6464
rect 5429 6418 5486 6464
rect 5532 6418 5562 6464
rect 5635 6418 5692 6464
rect 5738 6418 5773 6464
rect 5841 6418 5898 6464
rect 5944 6418 5957 6464
rect 6035 6418 6451 6464
rect 6497 6418 6568 6464
rect 6614 6418 6685 6464
rect 6731 6418 6803 6464
rect 6849 6418 6921 6464
rect 6967 6418 7039 6464
rect 7085 6462 7506 6464
rect 7085 6418 7488 6462
rect 7552 6418 7623 6464
rect 7669 6462 7740 6464
rect 7720 6418 7740 6462
rect 7786 6418 7858 6464
rect 7904 6418 7976 6464
rect 8022 6418 8094 6464
rect 8140 6418 8153 6464
rect 8255 6418 8618 6464
rect 8664 6418 8741 6464
rect 8787 6418 8864 6464
rect 8910 6418 9238 6464
rect 9284 6418 9327 6464
rect 9406 6446 14515 6484
rect 18502 6464 19474 6504
rect 18362 6418 18375 6464
rect 18421 6418 18478 6464
rect 18524 6418 18540 6464
rect 18627 6418 18684 6464
rect 18730 6418 18751 6464
rect 18833 6418 18890 6464
rect 18936 6418 18962 6464
rect 19039 6418 19096 6464
rect 19142 6418 19173 6464
rect 19449 6418 19474 6464
rect 19641 6470 20113 6516
rect 20159 6470 20300 6516
rect 20346 6470 20487 6516
rect 20533 6470 20673 6516
rect 20719 6470 20860 6516
rect 20906 6470 21254 6516
rect 21386 6505 21399 6551
rect 23373 6505 23386 6551
rect 19641 6460 21254 6470
rect 20078 6433 21254 6460
rect 21394 6480 21432 6505
rect 21484 6480 21612 6505
rect 21664 6480 21702 6505
rect 21394 6440 21702 6480
rect 23682 6446 23974 6678
rect 345 6367 637 6400
rect 4891 6412 4929 6418
rect 4981 6412 5140 6418
rect 5192 6412 5351 6418
rect 5403 6412 5562 6418
rect 5614 6412 5773 6418
rect 5825 6412 5863 6418
rect 4467 6367 4622 6374
rect 4891 6372 5863 6412
rect 6035 6378 6550 6418
rect 7036 6410 7488 6418
rect 7540 6410 7668 6418
rect 7720 6410 7758 6418
rect 7036 6378 7758 6410
rect 7450 6370 7758 6378
rect 345 6326 2439 6367
rect 345 6274 451 6326
rect 503 6274 662 6326
rect 714 6274 873 6326
rect 925 6274 1083 6326
rect 1135 6274 1294 6326
rect 1346 6274 1506 6326
rect 1558 6274 1717 6326
rect 1769 6274 1927 6326
rect 1979 6274 2138 6326
rect 2190 6274 2349 6326
rect 2401 6274 2439 6326
rect 345 6233 2439 6274
rect 4314 6326 4622 6367
rect 8255 6358 9320 6418
rect 18502 6412 18540 6418
rect 18592 6412 18751 6418
rect 18803 6412 18962 6418
rect 19014 6412 19173 6418
rect 19225 6412 19384 6418
rect 19436 6412 19474 6418
rect 18502 6372 19474 6412
rect 23682 6400 23820 6446
rect 23866 6400 23974 6446
rect 19696 6367 19852 6374
rect 23682 6367 23974 6400
rect 4314 6274 4352 6326
rect 4404 6323 4532 6326
rect 4404 6277 4513 6323
rect 4404 6274 4532 6277
rect 4584 6274 4622 6326
rect 4314 6233 4622 6274
rect 19696 6326 20005 6367
rect 19696 6274 19735 6326
rect 19787 6323 19915 6326
rect 19803 6277 19915 6323
rect 19787 6274 19915 6277
rect 19967 6274 20005 6326
rect 345 6200 637 6233
rect 4467 6226 4622 6233
rect 345 6154 452 6200
rect 498 6154 637 6200
rect 4891 6188 5863 6228
rect 7450 6222 7758 6230
rect 4891 6182 4929 6188
rect 4981 6182 5140 6188
rect 5192 6182 5351 6188
rect 5403 6182 5562 6188
rect 5614 6182 5773 6188
rect 5825 6182 5863 6188
rect 6035 6182 6550 6222
rect 7036 6190 7758 6222
rect 7036 6182 7488 6190
rect 7540 6182 7668 6190
rect 7720 6182 7758 6190
rect 8255 6182 9320 6242
rect 19696 6233 20005 6274
rect 21875 6326 23974 6367
rect 21875 6274 21913 6326
rect 21965 6274 22124 6326
rect 22176 6274 22335 6326
rect 22387 6274 22545 6326
rect 22597 6274 22756 6326
rect 22808 6274 22968 6326
rect 23020 6274 23179 6326
rect 23231 6274 23389 6326
rect 23441 6274 23600 6326
rect 23652 6274 23811 6326
rect 23863 6274 23974 6326
rect 21875 6233 23974 6274
rect 18502 6188 19474 6228
rect 19696 6226 19852 6233
rect 18502 6182 18540 6188
rect 18592 6182 18751 6188
rect 18803 6182 18962 6188
rect 19014 6182 19173 6188
rect 19225 6182 19384 6188
rect 19436 6182 19474 6188
rect 345 6037 637 6154
rect 3081 6138 4240 6167
rect 2616 6098 2924 6138
rect 2616 6095 2654 6098
rect 2706 6095 2834 6098
rect 2886 6095 2924 6098
rect 3081 6130 4679 6138
rect 4857 6136 4870 6182
rect 5120 6136 5140 6182
rect 5223 6136 5280 6182
rect 5326 6136 5351 6182
rect 5429 6136 5486 6182
rect 5532 6136 5562 6182
rect 5635 6136 5692 6182
rect 5738 6136 5773 6182
rect 5841 6136 5898 6182
rect 5944 6136 5957 6182
rect 6035 6136 6451 6182
rect 6497 6136 6568 6182
rect 6614 6136 6685 6182
rect 6731 6136 6803 6182
rect 6849 6136 6921 6182
rect 6967 6136 7039 6182
rect 7085 6138 7488 6182
rect 7085 6136 7506 6138
rect 7552 6136 7623 6182
rect 7720 6138 7740 6182
rect 7669 6136 7740 6138
rect 7786 6136 7858 6182
rect 7904 6136 7976 6182
rect 8022 6136 8094 6182
rect 8140 6136 8153 6182
rect 8255 6136 8618 6182
rect 8664 6136 8741 6182
rect 8787 6136 8864 6182
rect 8910 6136 9238 6182
rect 9284 6136 9327 6182
rect 933 6049 946 6095
rect 2920 6049 2933 6095
rect 3081 6084 3413 6130
rect 3459 6084 3599 6130
rect 3645 6084 3786 6130
rect 3832 6084 3973 6130
rect 4019 6084 4159 6130
rect 4205 6084 4679 6130
rect 4891 6096 5863 6136
rect 6035 6102 6550 6136
rect 7036 6102 7758 6136
rect 345 5991 452 6037
rect 498 5991 637 6037
rect 2616 6046 2654 6049
rect 2706 6046 2834 6049
rect 2886 6046 2924 6049
rect 2616 6005 2924 6046
rect 3081 6047 4679 6084
rect 345 5922 637 5991
rect 3081 5965 3149 6047
rect 345 5874 1090 5922
rect 345 5828 452 5874
rect 498 5871 1090 5874
rect 498 5828 946 5871
rect 345 5825 946 5828
rect 2920 5825 2933 5871
rect 345 5803 1090 5825
rect 345 5711 637 5803
rect 345 5665 452 5711
rect 498 5665 637 5711
rect 345 5547 637 5665
rect 2616 5650 2924 5690
rect 2616 5647 2654 5650
rect 2706 5647 2834 5650
rect 2886 5647 2924 5650
rect 933 5601 946 5647
rect 2920 5601 2933 5647
rect 2616 5598 2654 5601
rect 2706 5598 2834 5601
rect 2886 5598 2924 5601
rect 2616 5557 2924 5598
rect 345 5501 452 5547
rect 498 5501 637 5547
rect 3081 5543 3092 5965
rect 3138 5543 3149 5965
rect 4561 5990 4679 6047
rect 6035 6002 6151 6102
rect 7450 6097 7758 6102
rect 8255 6122 9320 6136
rect 4561 5958 5957 5990
rect 3825 5888 4315 5929
rect 3825 5871 3864 5888
rect 3916 5871 4044 5888
rect 4096 5871 4224 5888
rect 3268 5825 3281 5871
rect 3327 5825 3384 5871
rect 3430 5825 3487 5871
rect 3533 5825 3590 5871
rect 3636 5825 3693 5871
rect 3739 5825 3796 5871
rect 3842 5836 3864 5871
rect 3842 5825 3899 5836
rect 3945 5825 4002 5871
rect 4096 5836 4105 5871
rect 4048 5825 4105 5836
rect 4151 5825 4209 5871
rect 4276 5836 4315 5888
rect 4561 5912 4870 5958
rect 5120 5912 5177 5958
rect 5223 5912 5280 5958
rect 5326 5912 5383 5958
rect 5429 5912 5486 5958
rect 5532 5912 5589 5958
rect 5635 5912 5692 5958
rect 5738 5912 5795 5958
rect 5841 5912 5898 5958
rect 5944 5912 5957 5958
rect 4561 5868 5957 5912
rect 4255 5825 4315 5836
rect 3825 5796 4315 5825
rect 6035 5862 6072 6002
rect 6118 5862 6151 6002
rect 4891 5734 5863 5768
rect 6035 5759 6151 5862
rect 6237 6002 6370 6022
rect 6237 5963 6294 6002
rect 6237 5911 6275 5963
rect 6237 5862 6294 5911
rect 6340 5862 6370 6002
rect 8255 6000 8323 6122
rect 9406 6116 14515 6154
rect 18362 6136 18375 6182
rect 18421 6136 18478 6182
rect 18524 6136 18540 6182
rect 18627 6136 18684 6182
rect 18730 6136 18751 6182
rect 18833 6136 18890 6182
rect 18936 6136 18962 6182
rect 19039 6136 19096 6182
rect 19142 6136 19173 6182
rect 19449 6136 19474 6182
rect 23682 6200 23974 6233
rect 20078 6140 21254 6167
rect 9406 6070 13336 6116
rect 13382 6070 13503 6116
rect 13549 6070 13668 6116
rect 13714 6070 13833 6116
rect 13879 6095 14515 6116
rect 18502 6096 19474 6136
rect 19641 6130 21254 6140
rect 13879 6070 14409 6095
rect 9406 6067 14409 6070
rect 9406 6021 9441 6067
rect 9487 6065 14409 6067
rect 9487 6021 9591 6065
rect 9406 6013 9591 6021
rect 9643 6049 14409 6065
rect 14455 6049 14522 6095
rect 14568 6049 14635 6095
rect 14681 6049 14748 6095
rect 14794 6049 14861 6095
rect 14907 6049 14920 6095
rect 18154 6050 18284 6090
rect 9643 6034 14515 6049
rect 9643 6013 9682 6034
rect 9406 6010 9682 6013
rect 6521 5990 7282 5997
rect 6520 5958 7528 5990
rect 6438 5912 6451 5958
rect 6497 5956 6568 5958
rect 6497 5912 6558 5956
rect 6614 5912 6685 5958
rect 6731 5956 6803 5958
rect 6731 5912 6769 5956
rect 6849 5912 6921 5958
rect 6967 5956 7039 5958
rect 6967 5912 6981 5956
rect 6520 5904 6558 5912
rect 6610 5904 6769 5912
rect 6821 5904 6981 5912
rect 7033 5912 7039 5956
rect 7085 5956 7506 5958
rect 7085 5912 7192 5956
rect 7033 5904 7192 5912
rect 7244 5912 7506 5956
rect 7552 5912 7623 5958
rect 7669 5912 7740 5958
rect 7786 5912 7858 5958
rect 7904 5912 7976 5958
rect 8022 5912 8094 5958
rect 8140 5912 8153 5958
rect 7244 5904 7528 5912
rect 6520 5871 7528 5904
rect 6520 5870 7282 5871
rect 6521 5864 7282 5870
rect 6237 5839 6370 5862
rect 8255 5860 8266 6000
rect 8312 5860 8323 6000
rect 8611 5958 8920 5990
rect 9089 5958 9205 5990
rect 8605 5912 8618 5958
rect 8664 5912 8741 5958
rect 8787 5912 8864 5958
rect 8910 5912 8923 5958
rect 9089 5912 9238 5958
rect 9284 5912 9327 5958
rect 8255 5849 8323 5860
rect 6035 5734 6550 5759
rect 7036 5756 7528 5759
rect 7036 5734 7758 5756
rect 4857 5688 4870 5734
rect 5120 5728 5177 5734
rect 5120 5688 5140 5728
rect 5223 5688 5280 5734
rect 5326 5728 5383 5734
rect 5326 5688 5351 5728
rect 5429 5688 5486 5734
rect 5532 5728 5589 5734
rect 5532 5688 5562 5728
rect 5635 5688 5692 5734
rect 5738 5728 5795 5734
rect 5738 5688 5773 5728
rect 5841 5688 5898 5734
rect 5944 5688 5957 5734
rect 6035 5688 6451 5734
rect 6497 5688 6568 5734
rect 6614 5688 6685 5734
rect 6731 5688 6803 5734
rect 6849 5688 6921 5734
rect 6967 5688 7039 5734
rect 7085 5716 7506 5734
rect 7085 5688 7488 5716
rect 7552 5688 7623 5734
rect 7669 5716 7740 5734
rect 7720 5688 7740 5716
rect 7786 5688 7858 5734
rect 7904 5688 7976 5734
rect 8022 5688 8094 5734
rect 8140 5688 8153 5734
rect 3378 5647 3686 5682
rect 4891 5676 4929 5688
rect 4981 5676 5140 5688
rect 5192 5676 5351 5688
rect 5403 5676 5562 5688
rect 5614 5676 5773 5688
rect 5825 5676 5863 5688
rect 3268 5601 3281 5647
rect 3327 5601 3384 5647
rect 3430 5642 3487 5647
rect 3468 5601 3487 5642
rect 3533 5601 3590 5647
rect 3636 5642 3693 5647
rect 3648 5601 3693 5642
rect 3739 5601 3796 5647
rect 3842 5601 3899 5647
rect 3945 5601 4002 5647
rect 4048 5601 4105 5647
rect 4151 5601 4209 5647
rect 4255 5601 4268 5647
rect 4891 5636 5863 5676
rect 6035 5639 6550 5688
rect 7036 5664 7488 5688
rect 7540 5664 7668 5688
rect 7720 5664 7758 5688
rect 7036 5639 7758 5664
rect 7450 5623 7758 5639
rect 3378 5590 3416 5601
rect 3468 5590 3596 5601
rect 3648 5590 3686 5601
rect 3378 5549 3686 5590
rect 3081 5532 3149 5543
rect 345 5467 637 5501
rect 345 5426 2439 5467
rect 3844 5460 4605 5467
rect 345 5374 451 5426
rect 503 5374 662 5426
rect 714 5374 873 5426
rect 925 5423 1083 5426
rect 1135 5423 1294 5426
rect 1346 5423 1506 5426
rect 1558 5423 1717 5426
rect 1769 5423 1927 5426
rect 1979 5423 2138 5426
rect 2190 5423 2349 5426
rect 2401 5423 2439 5426
rect 3843 5426 4605 5460
rect 3843 5423 3881 5426
rect 3933 5423 4092 5426
rect 4144 5423 4304 5426
rect 925 5377 946 5423
rect 2920 5377 2933 5423
rect 3268 5377 3281 5423
rect 3327 5377 3384 5423
rect 3430 5377 3487 5423
rect 3533 5377 3590 5423
rect 3636 5377 3693 5423
rect 3739 5377 3796 5423
rect 3842 5377 3881 5423
rect 3945 5377 4002 5423
rect 4048 5377 4092 5423
rect 4151 5377 4209 5423
rect 4255 5377 4304 5423
rect 925 5374 1083 5377
rect 1135 5374 1294 5377
rect 1346 5374 1506 5377
rect 1558 5374 1717 5377
rect 1769 5374 1927 5377
rect 1979 5374 2138 5377
rect 2190 5374 2349 5377
rect 2401 5374 2439 5377
rect 345 5333 2439 5374
rect 3843 5374 3881 5377
rect 3933 5374 4092 5377
rect 4144 5374 4304 5377
rect 4356 5374 4515 5426
rect 4567 5374 4605 5426
rect 3843 5340 4605 5374
rect 3844 5333 4605 5340
rect 4779 5460 5961 5467
rect 4779 5426 6555 5460
rect 4779 5374 4817 5426
rect 4869 5374 5027 5426
rect 5079 5374 5238 5426
rect 5290 5374 5450 5426
rect 5502 5374 5661 5426
rect 5713 5374 5871 5426
rect 5923 5423 6555 5426
rect 5923 5377 6086 5423
rect 6320 5377 6555 5423
rect 5923 5374 6555 5377
rect 4779 5340 6555 5374
rect 7543 5426 8439 5467
rect 7543 5423 7927 5426
rect 7979 5423 8138 5426
rect 7543 5377 7554 5423
rect 8070 5377 8138 5423
rect 7543 5374 7927 5377
rect 7979 5374 8138 5377
rect 8190 5374 8349 5426
rect 8401 5374 8439 5426
rect 4779 5333 5961 5340
rect 7543 5333 8439 5374
rect 8611 5426 8920 5912
rect 8611 5374 8649 5426
rect 8701 5423 8829 5426
rect 8705 5377 8817 5423
rect 8701 5374 8829 5377
rect 8881 5374 8920 5426
rect 345 5299 637 5333
rect 345 5253 452 5299
rect 498 5253 637 5299
rect 345 5135 637 5253
rect 3081 5257 3149 5268
rect 2616 5202 2924 5243
rect 2616 5199 2654 5202
rect 2706 5199 2834 5202
rect 2886 5199 2924 5202
rect 933 5153 946 5199
rect 2920 5153 2933 5199
rect 345 5089 452 5135
rect 498 5089 637 5135
rect 2616 5150 2654 5153
rect 2706 5150 2834 5153
rect 2886 5150 2924 5153
rect 2616 5110 2924 5150
rect 345 4997 637 5089
rect 345 4975 1090 4997
rect 345 4972 946 4975
rect 345 4926 452 4972
rect 498 4929 946 4972
rect 2920 4929 2933 4975
rect 498 4926 1090 4929
rect 345 4878 1090 4926
rect 345 4809 637 4878
rect 345 4763 452 4809
rect 498 4763 637 4809
rect 3081 4835 3092 5257
rect 3138 4835 3149 5257
rect 3378 5210 3686 5251
rect 3378 5199 3416 5210
rect 3468 5199 3596 5210
rect 3648 5199 3686 5210
rect 3268 5153 3281 5199
rect 3327 5153 3384 5199
rect 3468 5158 3487 5199
rect 3430 5153 3487 5158
rect 3533 5153 3590 5199
rect 3648 5158 3693 5199
rect 3636 5153 3693 5158
rect 3739 5153 3796 5199
rect 3842 5153 3899 5199
rect 3945 5153 4002 5199
rect 4048 5153 4105 5199
rect 4151 5153 4209 5199
rect 4255 5153 4268 5199
rect 3378 5118 3686 5153
rect 4891 5124 5863 5164
rect 7450 5161 7758 5177
rect 4891 5112 4929 5124
rect 4981 5112 5140 5124
rect 5192 5112 5351 5124
rect 5403 5112 5562 5124
rect 5614 5112 5773 5124
rect 5825 5112 5863 5124
rect 6035 5112 6550 5161
rect 7036 5136 7758 5161
rect 7036 5112 7488 5136
rect 7540 5112 7668 5136
rect 7720 5112 7758 5136
rect 4857 5066 4870 5112
rect 5120 5072 5140 5112
rect 5120 5066 5177 5072
rect 5223 5066 5280 5112
rect 5326 5072 5351 5112
rect 5326 5066 5383 5072
rect 5429 5066 5486 5112
rect 5532 5072 5562 5112
rect 5532 5066 5589 5072
rect 5635 5066 5692 5112
rect 5738 5072 5773 5112
rect 5738 5066 5795 5072
rect 5841 5066 5898 5112
rect 5944 5066 5957 5112
rect 6035 5066 6451 5112
rect 6497 5066 6568 5112
rect 6614 5066 6685 5112
rect 6731 5066 6803 5112
rect 6849 5066 6921 5112
rect 6967 5066 7039 5112
rect 7085 5084 7488 5112
rect 7085 5066 7506 5084
rect 7552 5066 7623 5112
rect 7720 5084 7740 5112
rect 7669 5066 7740 5084
rect 7786 5066 7858 5112
rect 7904 5066 7976 5112
rect 8022 5066 8094 5112
rect 8140 5066 8153 5112
rect 4891 5032 5863 5066
rect 6035 5041 6550 5066
rect 7036 5044 7758 5066
rect 7036 5041 7528 5044
rect 3825 4975 4315 5004
rect 3268 4929 3281 4975
rect 3327 4929 3384 4975
rect 3430 4929 3487 4975
rect 3533 4929 3590 4975
rect 3636 4929 3693 4975
rect 3739 4929 3796 4975
rect 3842 4964 3899 4975
rect 3842 4929 3864 4964
rect 3945 4929 4002 4975
rect 4048 4964 4105 4975
rect 4096 4929 4105 4964
rect 4151 4929 4209 4975
rect 4255 4964 4315 4975
rect 3825 4912 3864 4929
rect 3916 4912 4044 4929
rect 4096 4912 4224 4929
rect 4276 4912 4315 4964
rect 6035 4938 6151 5041
rect 3825 4871 4315 4912
rect 4561 4888 5957 4932
rect 345 4646 637 4763
rect 2616 4754 2924 4795
rect 2616 4751 2654 4754
rect 2706 4751 2834 4754
rect 2886 4751 2924 4754
rect 3081 4753 3149 4835
rect 4561 4842 4870 4888
rect 5120 4842 5177 4888
rect 5223 4842 5280 4888
rect 5326 4842 5383 4888
rect 5429 4842 5486 4888
rect 5532 4842 5589 4888
rect 5635 4842 5692 4888
rect 5738 4842 5795 4888
rect 5841 4842 5898 4888
rect 5944 4842 5957 4888
rect 4561 4810 5957 4842
rect 4561 4753 4679 4810
rect 933 4705 946 4751
rect 2920 4705 2933 4751
rect 3081 4716 4679 4753
rect 2616 4702 2654 4705
rect 2706 4702 2834 4705
rect 2886 4702 2924 4705
rect 2616 4662 2924 4702
rect 3081 4670 3413 4716
rect 3459 4670 3599 4716
rect 3645 4670 3786 4716
rect 3832 4670 3973 4716
rect 4019 4670 4159 4716
rect 4205 4670 4679 4716
rect 6035 4798 6072 4938
rect 6118 4798 6151 4938
rect 3081 4662 4679 4670
rect 4891 4664 5863 4704
rect 6035 4698 6151 4798
rect 6237 4938 6370 4961
rect 6237 4889 6294 4938
rect 6237 4837 6275 4889
rect 6237 4798 6294 4837
rect 6340 4798 6370 4938
rect 8255 4940 8323 4951
rect 6521 4930 7282 4936
rect 6520 4929 7282 4930
rect 6520 4896 7528 4929
rect 6520 4888 6558 4896
rect 6610 4888 6769 4896
rect 6821 4888 6981 4896
rect 6438 4842 6451 4888
rect 6497 4844 6558 4888
rect 6497 4842 6568 4844
rect 6614 4842 6685 4888
rect 6731 4844 6769 4888
rect 6731 4842 6803 4844
rect 6849 4842 6921 4888
rect 6967 4844 6981 4888
rect 7033 4888 7192 4896
rect 7033 4844 7039 4888
rect 6967 4842 7039 4844
rect 7085 4844 7192 4888
rect 7244 4888 7528 4896
rect 7244 4844 7506 4888
rect 7085 4842 7506 4844
rect 7552 4842 7623 4888
rect 7669 4842 7740 4888
rect 7786 4842 7858 4888
rect 7904 4842 7976 4888
rect 8022 4842 8094 4888
rect 8140 4842 8153 4888
rect 6520 4810 7528 4842
rect 6521 4803 7282 4810
rect 6237 4778 6370 4798
rect 8255 4800 8266 4940
rect 8312 4800 8323 4940
rect 8611 4888 8920 5374
rect 9089 5460 9205 5912
rect 9520 5879 9682 6010
rect 9520 5827 9591 5879
rect 9643 5827 9682 5879
rect 9520 5787 9682 5827
rect 9334 5691 9462 5704
rect 9334 5664 9463 5691
rect 9334 5647 9372 5664
rect 9424 5647 9463 5664
rect 9324 5601 9337 5647
rect 9424 5612 9459 5647
rect 9383 5601 9459 5612
rect 9505 5601 9582 5647
rect 9628 5601 9705 5647
rect 9751 5601 9764 5647
rect 9843 5636 9959 6034
rect 11826 5895 14106 5936
rect 11826 5843 13042 5895
rect 13094 5843 14106 5895
rect 11826 5803 14106 5843
rect 13938 5759 14106 5803
rect 13938 5713 13955 5759
rect 14095 5713 14106 5759
rect 9334 5572 9463 5601
rect 9843 5590 9878 5636
rect 9924 5590 9959 5636
rect 9843 5553 9959 5590
rect 10315 5664 13121 5705
rect 13938 5702 14106 5713
rect 10315 5612 11532 5664
rect 11584 5612 13121 5664
rect 10315 5571 13121 5612
rect 14202 5647 14318 6034
rect 14997 6004 17976 6045
rect 14997 5990 15572 6004
rect 14997 5944 15061 5990
rect 15201 5952 15572 5990
rect 15624 5952 17976 6004
rect 15201 5944 17976 5952
rect 14498 5888 14838 5929
rect 14997 5911 17976 5944
rect 18154 5998 18193 6050
rect 18245 5998 18284 6050
rect 18154 5975 18284 5998
rect 19641 6084 20113 6130
rect 20159 6084 20300 6130
rect 20346 6084 20487 6130
rect 20533 6084 20673 6130
rect 20719 6084 20860 6130
rect 20906 6084 21254 6130
rect 21394 6120 21702 6160
rect 21394 6095 21432 6120
rect 21484 6095 21612 6120
rect 21664 6095 21702 6120
rect 23682 6154 23820 6200
rect 23866 6154 23974 6200
rect 19641 6047 21254 6084
rect 21386 6049 21399 6095
rect 23373 6049 23386 6095
rect 19641 5990 19757 6047
rect 14498 5871 14536 5888
rect 14588 5871 14748 5888
rect 14800 5871 14838 5888
rect 14396 5825 14409 5871
rect 14455 5825 14522 5871
rect 14588 5836 14635 5871
rect 14568 5825 14635 5836
rect 14681 5825 14748 5871
rect 14800 5836 14861 5871
rect 14794 5825 14861 5836
rect 14907 5825 14920 5871
rect 18154 5835 18219 5975
rect 18265 5835 18284 5975
rect 19417 5958 19757 5990
rect 18362 5912 18375 5958
rect 18421 5912 18478 5958
rect 18524 5912 18581 5958
rect 18627 5912 18684 5958
rect 18730 5912 18787 5958
rect 18833 5912 18890 5958
rect 18936 5912 18993 5958
rect 19039 5912 19096 5958
rect 19142 5912 19199 5958
rect 19449 5912 19757 5958
rect 21186 5995 21254 6047
rect 21394 6027 21702 6049
rect 19417 5871 19757 5912
rect 19859 5888 20409 5929
rect 18154 5832 18284 5835
rect 14498 5796 14838 5825
rect 18154 5780 18193 5832
rect 18245 5780 18284 5832
rect 19859 5836 19897 5888
rect 19949 5871 20108 5888
rect 20160 5871 20319 5888
rect 19949 5836 20064 5871
rect 20160 5836 20168 5871
rect 19859 5825 20064 5836
rect 20110 5825 20168 5836
rect 20214 5825 20271 5871
rect 20317 5836 20319 5871
rect 20371 5871 20409 5888
rect 20371 5836 20374 5871
rect 20317 5825 20374 5836
rect 20420 5825 20477 5871
rect 20523 5825 20580 5871
rect 20626 5825 20683 5871
rect 20729 5825 20786 5871
rect 20832 5825 20889 5871
rect 20935 5825 20992 5871
rect 21038 5825 21051 5871
rect 19859 5796 20409 5825
rect 18154 5739 18284 5780
rect 18502 5734 19474 5765
rect 18362 5688 18375 5734
rect 18421 5688 18478 5734
rect 18524 5725 18581 5734
rect 18524 5688 18540 5725
rect 18627 5688 18684 5734
rect 18730 5725 18787 5734
rect 18730 5688 18751 5725
rect 18833 5688 18890 5734
rect 18936 5725 18993 5734
rect 18936 5688 18962 5725
rect 19039 5688 19096 5734
rect 19142 5725 19199 5734
rect 19142 5688 19173 5725
rect 19449 5688 19474 5734
rect 18502 5673 18540 5688
rect 18592 5673 18751 5688
rect 18803 5673 18962 5688
rect 19014 5673 19173 5688
rect 19225 5673 19384 5688
rect 19436 5673 19474 5688
rect 14202 5601 14409 5647
rect 14455 5601 14522 5647
rect 14568 5601 14635 5647
rect 14681 5601 14748 5647
rect 14794 5601 14861 5647
rect 14907 5601 14920 5647
rect 18502 5633 19474 5673
rect 20632 5650 20940 5690
rect 20632 5647 20670 5650
rect 20722 5647 20850 5650
rect 20902 5647 20940 5650
rect 12959 5564 13121 5571
rect 12959 5518 12970 5564
rect 13110 5518 13121 5564
rect 12959 5507 13121 5518
rect 15181 5587 18143 5623
rect 20051 5601 20064 5647
rect 20110 5601 20168 5647
rect 20214 5601 20271 5647
rect 20317 5601 20374 5647
rect 20420 5601 20477 5647
rect 20523 5601 20580 5647
rect 20626 5601 20670 5647
rect 20729 5601 20786 5647
rect 20832 5601 20850 5647
rect 20935 5601 20992 5647
rect 21038 5601 21051 5647
rect 15181 5541 15216 5587
rect 15262 5541 15374 5587
rect 15420 5541 15532 5587
rect 15578 5541 15690 5587
rect 15736 5541 15848 5587
rect 15894 5541 16006 5587
rect 16052 5541 16165 5587
rect 16211 5541 16323 5587
rect 16369 5541 16481 5587
rect 16527 5541 16639 5587
rect 16685 5541 16797 5587
rect 16843 5541 16955 5587
rect 17001 5541 17113 5587
rect 17159 5541 17272 5587
rect 17318 5541 17430 5587
rect 17476 5541 17588 5587
rect 17634 5541 17746 5587
rect 17792 5541 17904 5587
rect 17950 5541 18062 5587
rect 18108 5541 18143 5587
rect 20632 5598 20670 5601
rect 20722 5598 20850 5601
rect 20902 5598 20940 5601
rect 20632 5557 20940 5598
rect 21186 5573 21197 5995
rect 21243 5573 21254 5995
rect 23682 5922 23974 6154
rect 23182 5871 23974 5922
rect 21386 5825 21399 5871
rect 23373 5825 23974 5871
rect 23182 5803 23974 5825
rect 23682 5711 23974 5803
rect 21394 5657 21702 5697
rect 21394 5647 21432 5657
rect 21484 5647 21612 5657
rect 21664 5647 21702 5657
rect 23682 5665 23820 5711
rect 23866 5665 23974 5711
rect 21386 5601 21399 5647
rect 23373 5601 23386 5647
rect 21186 5562 21254 5573
rect 21394 5564 21702 5601
rect 9812 5460 10120 5467
rect 10385 5460 12583 5474
rect 13350 5460 14111 5467
rect 9089 5437 12583 5460
rect 13301 5437 14111 5460
rect 9089 5426 14111 5437
rect 9089 5423 9850 5426
rect 9089 5377 9337 5423
rect 9383 5377 9459 5423
rect 9505 5377 9582 5423
rect 9628 5377 9705 5423
rect 9751 5377 9850 5423
rect 9089 5374 9850 5377
rect 9902 5374 10030 5426
rect 10082 5423 13387 5426
rect 10082 5377 10433 5423
rect 10479 5377 10591 5423
rect 10637 5377 10749 5423
rect 10795 5377 10907 5423
rect 10953 5377 11066 5423
rect 11112 5377 11224 5423
rect 11270 5377 11382 5423
rect 11428 5377 11540 5423
rect 11586 5377 11698 5423
rect 11744 5377 11856 5423
rect 11902 5377 12015 5423
rect 12061 5377 12173 5423
rect 12219 5377 12331 5423
rect 12377 5377 12489 5423
rect 12535 5377 13336 5423
rect 13382 5377 13387 5423
rect 10082 5374 13387 5377
rect 13439 5423 13598 5426
rect 13439 5377 13503 5423
rect 13549 5377 13598 5423
rect 13439 5374 13598 5377
rect 13650 5423 13810 5426
rect 13862 5423 14021 5426
rect 13650 5377 13668 5423
rect 13714 5377 13810 5423
rect 13879 5377 14021 5423
rect 13650 5374 13810 5377
rect 13862 5374 14021 5377
rect 14073 5374 14111 5426
rect 9089 5363 14111 5374
rect 9089 5340 12583 5363
rect 13301 5340 14111 5363
rect 9089 4888 9205 5340
rect 9812 5333 10120 5340
rect 10385 5326 12583 5340
rect 13350 5333 14111 5340
rect 14393 5460 14943 5467
rect 15181 5460 18143 5541
rect 23682 5547 23974 5665
rect 23682 5501 23820 5547
rect 23866 5501 23974 5547
rect 23682 5467 23974 5501
rect 18397 5460 19579 5467
rect 19905 5460 20456 5467
rect 14393 5426 19579 5460
rect 14393 5423 14431 5426
rect 14483 5423 14642 5426
rect 14694 5423 14853 5426
rect 14905 5423 18435 5426
rect 14393 5377 14409 5423
rect 14483 5377 14522 5423
rect 14568 5377 14635 5423
rect 14694 5377 14748 5423
rect 14794 5377 14853 5423
rect 14907 5377 15216 5423
rect 15262 5377 15374 5423
rect 15420 5377 15532 5423
rect 15578 5377 15690 5423
rect 15736 5377 15848 5423
rect 15894 5377 16006 5423
rect 16052 5377 16165 5423
rect 16211 5377 16323 5423
rect 16369 5377 16481 5423
rect 16527 5377 16639 5423
rect 16685 5377 16797 5423
rect 16843 5377 16955 5423
rect 17001 5377 17113 5423
rect 17159 5377 17272 5423
rect 17318 5377 17430 5423
rect 17476 5377 17588 5423
rect 17634 5377 17746 5423
rect 17792 5377 17904 5423
rect 17950 5377 18062 5423
rect 18108 5377 18435 5423
rect 14393 5374 14431 5377
rect 14483 5374 14642 5377
rect 14694 5374 14853 5377
rect 14905 5374 18435 5377
rect 18487 5374 18645 5426
rect 18697 5374 18856 5426
rect 18908 5374 19068 5426
rect 19120 5374 19279 5426
rect 19331 5374 19489 5426
rect 19541 5374 19579 5426
rect 14393 5340 19579 5374
rect 19904 5426 20456 5460
rect 19904 5374 19943 5426
rect 19995 5423 20154 5426
rect 20206 5423 20365 5426
rect 20417 5423 20456 5426
rect 21875 5426 23974 5467
rect 21875 5423 21913 5426
rect 21965 5423 22124 5426
rect 22176 5423 22335 5426
rect 22387 5423 22545 5426
rect 22597 5423 22756 5426
rect 22808 5423 22968 5426
rect 23020 5423 23179 5426
rect 23231 5423 23389 5426
rect 19995 5377 20064 5423
rect 20110 5377 20154 5423
rect 20214 5377 20271 5423
rect 20317 5377 20365 5423
rect 20420 5377 20477 5423
rect 20523 5377 20580 5423
rect 20626 5377 20683 5423
rect 20729 5377 20786 5423
rect 20832 5377 20889 5423
rect 20935 5377 20992 5423
rect 21038 5377 21051 5423
rect 21386 5377 21399 5423
rect 23373 5377 23389 5423
rect 19995 5374 20154 5377
rect 20206 5374 20365 5377
rect 20417 5374 20456 5377
rect 19904 5340 20456 5374
rect 14393 5333 14943 5340
rect 12959 5282 13121 5293
rect 9334 5199 9463 5228
rect 9843 5210 9959 5247
rect 12959 5236 12970 5282
rect 13110 5236 13121 5282
rect 12959 5229 13121 5236
rect 9324 5153 9337 5199
rect 9383 5188 9459 5199
rect 9424 5153 9459 5188
rect 9505 5153 9582 5199
rect 9628 5153 9705 5199
rect 9751 5153 9764 5199
rect 9843 5164 9878 5210
rect 9924 5164 9959 5210
rect 9334 5136 9372 5153
rect 9424 5136 9463 5153
rect 9334 5109 9463 5136
rect 9334 5096 9462 5109
rect 9520 4973 9682 5013
rect 9520 4921 9591 4973
rect 9643 4921 9682 4973
rect 8605 4842 8618 4888
rect 8664 4842 8741 4888
rect 8787 4842 8864 4888
rect 8910 4842 8923 4888
rect 9089 4842 9238 4888
rect 9284 4842 9327 4888
rect 8611 4810 8920 4842
rect 9089 4810 9205 4842
rect 7450 4698 7758 4703
rect 6035 4664 6550 4698
rect 7036 4664 7758 4698
rect 8255 4678 8323 4800
rect 9520 4790 9682 4921
rect 9406 4787 9682 4790
rect 9406 4779 9591 4787
rect 9406 4733 9441 4779
rect 9487 4735 9591 4779
rect 9643 4766 9682 4787
rect 9843 4766 9959 5164
rect 10315 5188 13121 5229
rect 15181 5259 18143 5340
rect 18397 5333 19579 5340
rect 19905 5333 20456 5340
rect 21875 5374 21913 5377
rect 21965 5374 22124 5377
rect 22176 5374 22335 5377
rect 22387 5374 22545 5377
rect 22597 5374 22756 5377
rect 22808 5374 22968 5377
rect 23020 5374 23179 5377
rect 23231 5374 23389 5377
rect 23441 5374 23600 5426
rect 23652 5374 23811 5426
rect 23863 5374 23974 5426
rect 21875 5333 23974 5374
rect 15181 5213 15216 5259
rect 15262 5213 15374 5259
rect 15420 5213 15532 5259
rect 15578 5213 15690 5259
rect 15736 5213 15848 5259
rect 15894 5213 16006 5259
rect 16052 5213 16165 5259
rect 16211 5213 16323 5259
rect 16369 5213 16481 5259
rect 16527 5213 16639 5259
rect 16685 5213 16797 5259
rect 16843 5213 16955 5259
rect 17001 5213 17113 5259
rect 17159 5213 17272 5259
rect 17318 5213 17430 5259
rect 17476 5213 17588 5259
rect 17634 5213 17746 5259
rect 17792 5213 17904 5259
rect 17950 5213 18062 5259
rect 18108 5213 18143 5259
rect 23682 5299 23974 5333
rect 23682 5253 23820 5299
rect 23866 5253 23974 5299
rect 10315 5136 11532 5188
rect 11584 5136 13121 5188
rect 10315 5095 13121 5136
rect 14202 5153 14409 5199
rect 14455 5153 14522 5199
rect 14568 5153 14635 5199
rect 14681 5153 14748 5199
rect 14794 5153 14861 5199
rect 14907 5153 14920 5199
rect 15181 5177 18143 5213
rect 20632 5202 20940 5243
rect 20632 5199 20670 5202
rect 20722 5199 20850 5202
rect 20902 5199 20940 5202
rect 21186 5227 21254 5238
rect 13938 5087 14106 5098
rect 13938 5041 13955 5087
rect 14095 5041 14106 5087
rect 13938 4997 14106 5041
rect 11826 4957 14106 4997
rect 11826 4905 13042 4957
rect 13094 4905 14106 4957
rect 11826 4864 14106 4905
rect 14202 4766 14318 5153
rect 18502 5127 19474 5167
rect 20051 5153 20064 5199
rect 20110 5153 20168 5199
rect 20214 5153 20271 5199
rect 20317 5153 20374 5199
rect 20420 5153 20477 5199
rect 20523 5153 20580 5199
rect 20626 5153 20670 5199
rect 20729 5153 20786 5199
rect 20832 5153 20850 5199
rect 20935 5153 20992 5199
rect 21038 5153 21051 5199
rect 18502 5112 18540 5127
rect 18592 5112 18751 5127
rect 18803 5112 18962 5127
rect 19014 5112 19173 5127
rect 19225 5112 19384 5127
rect 19436 5112 19474 5127
rect 18362 5066 18375 5112
rect 18421 5066 18478 5112
rect 18524 5075 18540 5112
rect 18524 5066 18581 5075
rect 18627 5066 18684 5112
rect 18730 5075 18751 5112
rect 18730 5066 18787 5075
rect 18833 5066 18890 5112
rect 18936 5075 18962 5112
rect 18936 5066 18993 5075
rect 19039 5066 19096 5112
rect 19142 5075 19173 5112
rect 19142 5066 19199 5075
rect 19449 5066 19474 5112
rect 20632 5150 20670 5153
rect 20722 5150 20850 5153
rect 20902 5150 20940 5153
rect 20632 5110 20940 5150
rect 18154 5020 18284 5061
rect 18502 5035 19474 5066
rect 14498 4975 14838 5004
rect 14396 4929 14409 4975
rect 14455 4929 14522 4975
rect 14568 4964 14635 4975
rect 14588 4929 14635 4964
rect 14681 4929 14748 4975
rect 14794 4964 14861 4975
rect 14800 4929 14861 4964
rect 14907 4929 14920 4975
rect 18154 4968 18193 5020
rect 18245 4968 18284 5020
rect 18154 4965 18284 4968
rect 14498 4912 14536 4929
rect 14588 4912 14748 4929
rect 14800 4912 14838 4929
rect 14498 4871 14838 4912
rect 14997 4856 17976 4889
rect 14997 4810 15061 4856
rect 15201 4848 17976 4856
rect 15201 4810 15950 4848
rect 14997 4796 15950 4810
rect 16002 4796 17976 4848
rect 9643 4751 14515 4766
rect 14997 4755 17976 4796
rect 18154 4825 18219 4965
rect 18265 4825 18284 4965
rect 19859 4975 20409 5004
rect 19859 4964 20064 4975
rect 20110 4964 20168 4975
rect 19417 4888 19757 4929
rect 18362 4842 18375 4888
rect 18421 4842 18478 4888
rect 18524 4842 18581 4888
rect 18627 4842 18684 4888
rect 18730 4842 18787 4888
rect 18833 4842 18890 4888
rect 18936 4842 18993 4888
rect 19039 4842 19096 4888
rect 19142 4842 19199 4888
rect 19449 4842 19757 4888
rect 19859 4912 19897 4964
rect 19949 4929 20064 4964
rect 20160 4929 20168 4964
rect 20214 4929 20271 4975
rect 20317 4964 20374 4975
rect 20317 4929 20319 4964
rect 19949 4912 20108 4929
rect 20160 4912 20319 4929
rect 20371 4929 20374 4964
rect 20420 4929 20477 4975
rect 20523 4929 20580 4975
rect 20626 4929 20683 4975
rect 20729 4929 20786 4975
rect 20832 4929 20889 4975
rect 20935 4929 20992 4975
rect 21038 4929 21051 4975
rect 20371 4912 20409 4929
rect 19859 4871 20409 4912
rect 18154 4802 18284 4825
rect 19417 4810 19757 4842
rect 9643 4735 14409 4751
rect 9487 4733 14409 4735
rect 9406 4730 14409 4733
rect 9406 4684 13336 4730
rect 13382 4684 13503 4730
rect 13549 4684 13668 4730
rect 13714 4684 13833 4730
rect 13879 4705 14409 4730
rect 14455 4705 14522 4751
rect 14568 4705 14635 4751
rect 14681 4705 14748 4751
rect 14794 4705 14861 4751
rect 14907 4705 14920 4751
rect 18154 4750 18193 4802
rect 18245 4750 18284 4802
rect 18154 4710 18284 4750
rect 19641 4753 19757 4810
rect 21186 4805 21197 5227
rect 21243 4805 21254 5227
rect 21394 5199 21702 5236
rect 21386 5153 21399 5199
rect 23373 5153 23386 5199
rect 21394 5143 21432 5153
rect 21484 5143 21612 5153
rect 21664 5143 21702 5153
rect 21394 5103 21702 5143
rect 23682 5135 23974 5253
rect 23682 5089 23820 5135
rect 23866 5089 23974 5135
rect 23682 4997 23974 5089
rect 23182 4975 23974 4997
rect 21386 4929 21399 4975
rect 23373 4929 23974 4975
rect 23182 4878 23974 4929
rect 21186 4753 21254 4805
rect 19641 4716 21254 4753
rect 21394 4751 21702 4773
rect 13879 4684 14515 4705
rect 8255 4664 9320 4678
rect 345 4600 452 4646
rect 498 4600 637 4646
rect 3081 4633 4240 4662
rect 4857 4618 4870 4664
rect 5120 4618 5140 4664
rect 5223 4618 5280 4664
rect 5326 4618 5351 4664
rect 5429 4618 5486 4664
rect 5532 4618 5562 4664
rect 5635 4618 5692 4664
rect 5738 4618 5773 4664
rect 5841 4618 5898 4664
rect 5944 4618 5957 4664
rect 6035 4618 6451 4664
rect 6497 4618 6568 4664
rect 6614 4618 6685 4664
rect 6731 4618 6803 4664
rect 6849 4618 6921 4664
rect 6967 4618 7039 4664
rect 7085 4662 7506 4664
rect 7085 4618 7488 4662
rect 7552 4618 7623 4664
rect 7669 4662 7740 4664
rect 7720 4618 7740 4662
rect 7786 4618 7858 4664
rect 7904 4618 7976 4664
rect 8022 4618 8094 4664
rect 8140 4618 8153 4664
rect 8255 4618 8618 4664
rect 8664 4618 8741 4664
rect 8787 4618 8864 4664
rect 8910 4618 9238 4664
rect 9284 4618 9327 4664
rect 9406 4646 14515 4684
rect 18502 4664 19474 4704
rect 18362 4618 18375 4664
rect 18421 4618 18478 4664
rect 18524 4618 18540 4664
rect 18627 4618 18684 4664
rect 18730 4618 18751 4664
rect 18833 4618 18890 4664
rect 18936 4618 18962 4664
rect 19039 4618 19096 4664
rect 19142 4618 19173 4664
rect 19449 4618 19474 4664
rect 19641 4670 20113 4716
rect 20159 4670 20300 4716
rect 20346 4670 20487 4716
rect 20533 4670 20673 4716
rect 20719 4670 20860 4716
rect 20906 4670 21254 4716
rect 21386 4705 21399 4751
rect 23373 4705 23386 4751
rect 19641 4660 21254 4670
rect 20078 4633 21254 4660
rect 21394 4680 21432 4705
rect 21484 4680 21612 4705
rect 21664 4680 21702 4705
rect 21394 4640 21702 4680
rect 23682 4646 23974 4878
rect 345 4567 637 4600
rect 4891 4612 4929 4618
rect 4981 4612 5140 4618
rect 5192 4612 5351 4618
rect 5403 4612 5562 4618
rect 5614 4612 5773 4618
rect 5825 4612 5863 4618
rect 4467 4567 4622 4574
rect 4891 4572 5863 4612
rect 6035 4578 6550 4618
rect 7036 4610 7488 4618
rect 7540 4610 7668 4618
rect 7720 4610 7758 4618
rect 7036 4578 7758 4610
rect 7450 4570 7758 4578
rect 345 4526 2439 4567
rect 345 4474 451 4526
rect 503 4474 662 4526
rect 714 4474 873 4526
rect 925 4474 1083 4526
rect 1135 4474 1294 4526
rect 1346 4474 1506 4526
rect 1558 4474 1717 4526
rect 1769 4474 1927 4526
rect 1979 4474 2138 4526
rect 2190 4474 2349 4526
rect 2401 4474 2439 4526
rect 345 4433 2439 4474
rect 4314 4526 4622 4567
rect 8255 4558 9320 4618
rect 18502 4612 18540 4618
rect 18592 4612 18751 4618
rect 18803 4612 18962 4618
rect 19014 4612 19173 4618
rect 19225 4612 19384 4618
rect 19436 4612 19474 4618
rect 18502 4572 19474 4612
rect 23682 4600 23820 4646
rect 23866 4600 23974 4646
rect 19696 4567 19852 4574
rect 23682 4567 23974 4600
rect 4314 4474 4352 4526
rect 4404 4523 4532 4526
rect 4404 4477 4513 4523
rect 4404 4474 4532 4477
rect 4584 4474 4622 4526
rect 4314 4433 4622 4474
rect 19696 4526 20005 4567
rect 19696 4474 19735 4526
rect 19787 4523 19915 4526
rect 19803 4477 19915 4523
rect 19787 4474 19915 4477
rect 19967 4474 20005 4526
rect 345 4400 637 4433
rect 4467 4426 4622 4433
rect 345 4354 452 4400
rect 498 4354 637 4400
rect 4891 4388 5863 4428
rect 7450 4422 7758 4430
rect 4891 4382 4929 4388
rect 4981 4382 5140 4388
rect 5192 4382 5351 4388
rect 5403 4382 5562 4388
rect 5614 4382 5773 4388
rect 5825 4382 5863 4388
rect 6035 4382 6550 4422
rect 7036 4390 7758 4422
rect 7036 4382 7488 4390
rect 7540 4382 7668 4390
rect 7720 4382 7758 4390
rect 8255 4382 9320 4442
rect 19696 4433 20005 4474
rect 21875 4526 23974 4567
rect 21875 4474 21913 4526
rect 21965 4474 22124 4526
rect 22176 4474 22335 4526
rect 22387 4474 22545 4526
rect 22597 4474 22756 4526
rect 22808 4474 22968 4526
rect 23020 4474 23179 4526
rect 23231 4474 23389 4526
rect 23441 4474 23600 4526
rect 23652 4474 23811 4526
rect 23863 4474 23974 4526
rect 21875 4433 23974 4474
rect 18502 4388 19474 4428
rect 19696 4426 19852 4433
rect 18502 4382 18540 4388
rect 18592 4382 18751 4388
rect 18803 4382 18962 4388
rect 19014 4382 19173 4388
rect 19225 4382 19384 4388
rect 19436 4382 19474 4388
rect 345 4237 637 4354
rect 3081 4338 4240 4367
rect 2616 4298 2924 4338
rect 2616 4295 2654 4298
rect 2706 4295 2834 4298
rect 2886 4295 2924 4298
rect 3081 4330 4679 4338
rect 4857 4336 4870 4382
rect 5120 4336 5140 4382
rect 5223 4336 5280 4382
rect 5326 4336 5351 4382
rect 5429 4336 5486 4382
rect 5532 4336 5562 4382
rect 5635 4336 5692 4382
rect 5738 4336 5773 4382
rect 5841 4336 5898 4382
rect 5944 4336 5957 4382
rect 6035 4336 6451 4382
rect 6497 4336 6568 4382
rect 6614 4336 6685 4382
rect 6731 4336 6803 4382
rect 6849 4336 6921 4382
rect 6967 4336 7039 4382
rect 7085 4338 7488 4382
rect 7085 4336 7506 4338
rect 7552 4336 7623 4382
rect 7720 4338 7740 4382
rect 7669 4336 7740 4338
rect 7786 4336 7858 4382
rect 7904 4336 7976 4382
rect 8022 4336 8094 4382
rect 8140 4336 8153 4382
rect 8255 4336 8618 4382
rect 8664 4336 8741 4382
rect 8787 4336 8864 4382
rect 8910 4336 9238 4382
rect 9284 4336 9327 4382
rect 933 4249 946 4295
rect 2920 4249 2933 4295
rect 3081 4284 3413 4330
rect 3459 4284 3599 4330
rect 3645 4284 3786 4330
rect 3832 4284 3973 4330
rect 4019 4284 4159 4330
rect 4205 4284 4679 4330
rect 4891 4296 5863 4336
rect 6035 4302 6550 4336
rect 7036 4302 7758 4336
rect 345 4191 452 4237
rect 498 4191 637 4237
rect 2616 4246 2654 4249
rect 2706 4246 2834 4249
rect 2886 4246 2924 4249
rect 2616 4205 2924 4246
rect 3081 4247 4679 4284
rect 345 4122 637 4191
rect 3081 4165 3149 4247
rect 345 4074 1090 4122
rect 345 4028 452 4074
rect 498 4071 1090 4074
rect 498 4028 946 4071
rect 345 4025 946 4028
rect 2920 4025 2933 4071
rect 345 4003 1090 4025
rect 345 3911 637 4003
rect 345 3865 452 3911
rect 498 3865 637 3911
rect 345 3747 637 3865
rect 2616 3850 2924 3890
rect 2616 3847 2654 3850
rect 2706 3847 2834 3850
rect 2886 3847 2924 3850
rect 933 3801 946 3847
rect 2920 3801 2933 3847
rect 2616 3798 2654 3801
rect 2706 3798 2834 3801
rect 2886 3798 2924 3801
rect 2616 3757 2924 3798
rect 345 3701 452 3747
rect 498 3701 637 3747
rect 3081 3743 3092 4165
rect 3138 3743 3149 4165
rect 4561 4190 4679 4247
rect 6035 4202 6151 4302
rect 7450 4297 7758 4302
rect 8255 4322 9320 4336
rect 4561 4158 5957 4190
rect 3825 4088 4315 4129
rect 3825 4071 3864 4088
rect 3916 4071 4044 4088
rect 4096 4071 4224 4088
rect 3268 4025 3281 4071
rect 3327 4025 3384 4071
rect 3430 4025 3487 4071
rect 3533 4025 3590 4071
rect 3636 4025 3693 4071
rect 3739 4025 3796 4071
rect 3842 4036 3864 4071
rect 3842 4025 3899 4036
rect 3945 4025 4002 4071
rect 4096 4036 4105 4071
rect 4048 4025 4105 4036
rect 4151 4025 4209 4071
rect 4276 4036 4315 4088
rect 4561 4112 4870 4158
rect 5120 4112 5177 4158
rect 5223 4112 5280 4158
rect 5326 4112 5383 4158
rect 5429 4112 5486 4158
rect 5532 4112 5589 4158
rect 5635 4112 5692 4158
rect 5738 4112 5795 4158
rect 5841 4112 5898 4158
rect 5944 4112 5957 4158
rect 4561 4068 5957 4112
rect 4255 4025 4315 4036
rect 3825 3996 4315 4025
rect 6035 4062 6072 4202
rect 6118 4062 6151 4202
rect 4891 3934 5863 3968
rect 6035 3959 6151 4062
rect 6237 4202 6370 4222
rect 6237 4163 6294 4202
rect 6237 4111 6275 4163
rect 6237 4062 6294 4111
rect 6340 4062 6370 4202
rect 8255 4200 8323 4322
rect 9406 4316 14515 4354
rect 18362 4336 18375 4382
rect 18421 4336 18478 4382
rect 18524 4336 18540 4382
rect 18627 4336 18684 4382
rect 18730 4336 18751 4382
rect 18833 4336 18890 4382
rect 18936 4336 18962 4382
rect 19039 4336 19096 4382
rect 19142 4336 19173 4382
rect 19449 4336 19474 4382
rect 23682 4400 23974 4433
rect 20078 4340 21254 4367
rect 9406 4270 13336 4316
rect 13382 4270 13503 4316
rect 13549 4270 13668 4316
rect 13714 4270 13833 4316
rect 13879 4295 14515 4316
rect 18502 4296 19474 4336
rect 19641 4330 21254 4340
rect 13879 4270 14409 4295
rect 9406 4267 14409 4270
rect 9406 4221 9441 4267
rect 9487 4265 14409 4267
rect 9487 4221 9591 4265
rect 9406 4213 9591 4221
rect 9643 4249 14409 4265
rect 14455 4249 14522 4295
rect 14568 4249 14635 4295
rect 14681 4249 14748 4295
rect 14794 4249 14861 4295
rect 14907 4249 14920 4295
rect 18154 4250 18284 4290
rect 9643 4234 14515 4249
rect 9643 4213 9682 4234
rect 9406 4210 9682 4213
rect 6521 4190 7282 4197
rect 6520 4158 7528 4190
rect 6438 4112 6451 4158
rect 6497 4156 6568 4158
rect 6497 4112 6558 4156
rect 6614 4112 6685 4158
rect 6731 4156 6803 4158
rect 6731 4112 6769 4156
rect 6849 4112 6921 4158
rect 6967 4156 7039 4158
rect 6967 4112 6981 4156
rect 6520 4104 6558 4112
rect 6610 4104 6769 4112
rect 6821 4104 6981 4112
rect 7033 4112 7039 4156
rect 7085 4156 7506 4158
rect 7085 4112 7192 4156
rect 7033 4104 7192 4112
rect 7244 4112 7506 4156
rect 7552 4112 7623 4158
rect 7669 4112 7740 4158
rect 7786 4112 7858 4158
rect 7904 4112 7976 4158
rect 8022 4112 8094 4158
rect 8140 4112 8153 4158
rect 7244 4104 7528 4112
rect 6520 4071 7528 4104
rect 6520 4070 7282 4071
rect 6521 4064 7282 4070
rect 6237 4039 6370 4062
rect 8255 4060 8266 4200
rect 8312 4060 8323 4200
rect 8611 4158 8920 4190
rect 9089 4158 9205 4190
rect 8605 4112 8618 4158
rect 8664 4112 8741 4158
rect 8787 4112 8864 4158
rect 8910 4112 8923 4158
rect 9089 4112 9238 4158
rect 9284 4112 9327 4158
rect 8255 4049 8323 4060
rect 6035 3934 6550 3959
rect 7036 3956 7528 3959
rect 7036 3934 7758 3956
rect 4857 3888 4870 3934
rect 5120 3928 5177 3934
rect 5120 3888 5140 3928
rect 5223 3888 5280 3934
rect 5326 3928 5383 3934
rect 5326 3888 5351 3928
rect 5429 3888 5486 3934
rect 5532 3928 5589 3934
rect 5532 3888 5562 3928
rect 5635 3888 5692 3934
rect 5738 3928 5795 3934
rect 5738 3888 5773 3928
rect 5841 3888 5898 3934
rect 5944 3888 5957 3934
rect 6035 3888 6451 3934
rect 6497 3888 6568 3934
rect 6614 3888 6685 3934
rect 6731 3888 6803 3934
rect 6849 3888 6921 3934
rect 6967 3888 7039 3934
rect 7085 3916 7506 3934
rect 7085 3888 7488 3916
rect 7552 3888 7623 3934
rect 7669 3916 7740 3934
rect 7720 3888 7740 3916
rect 7786 3888 7858 3934
rect 7904 3888 7976 3934
rect 8022 3888 8094 3934
rect 8140 3888 8153 3934
rect 3378 3847 3686 3882
rect 4891 3876 4929 3888
rect 4981 3876 5140 3888
rect 5192 3876 5351 3888
rect 5403 3876 5562 3888
rect 5614 3876 5773 3888
rect 5825 3876 5863 3888
rect 3268 3801 3281 3847
rect 3327 3801 3384 3847
rect 3430 3842 3487 3847
rect 3468 3801 3487 3842
rect 3533 3801 3590 3847
rect 3636 3842 3693 3847
rect 3648 3801 3693 3842
rect 3739 3801 3796 3847
rect 3842 3801 3899 3847
rect 3945 3801 4002 3847
rect 4048 3801 4105 3847
rect 4151 3801 4209 3847
rect 4255 3801 4268 3847
rect 4891 3836 5863 3876
rect 6035 3839 6550 3888
rect 7036 3864 7488 3888
rect 7540 3864 7668 3888
rect 7720 3864 7758 3888
rect 7036 3839 7758 3864
rect 7450 3823 7758 3839
rect 3378 3790 3416 3801
rect 3468 3790 3596 3801
rect 3648 3790 3686 3801
rect 3378 3749 3686 3790
rect 3081 3732 3149 3743
rect 345 3667 637 3701
rect 345 3626 2439 3667
rect 3844 3660 4605 3667
rect 345 3574 451 3626
rect 503 3574 662 3626
rect 714 3574 873 3626
rect 925 3623 1083 3626
rect 1135 3623 1294 3626
rect 1346 3623 1506 3626
rect 1558 3623 1717 3626
rect 1769 3623 1927 3626
rect 1979 3623 2138 3626
rect 2190 3623 2349 3626
rect 2401 3623 2439 3626
rect 3843 3626 4605 3660
rect 3843 3623 3881 3626
rect 3933 3623 4092 3626
rect 4144 3623 4304 3626
rect 925 3577 946 3623
rect 2920 3577 2933 3623
rect 3268 3577 3281 3623
rect 3327 3577 3384 3623
rect 3430 3577 3487 3623
rect 3533 3577 3590 3623
rect 3636 3577 3693 3623
rect 3739 3577 3796 3623
rect 3842 3577 3881 3623
rect 3945 3577 4002 3623
rect 4048 3577 4092 3623
rect 4151 3577 4209 3623
rect 4255 3577 4304 3623
rect 925 3574 1083 3577
rect 1135 3574 1294 3577
rect 1346 3574 1506 3577
rect 1558 3574 1717 3577
rect 1769 3574 1927 3577
rect 1979 3574 2138 3577
rect 2190 3574 2349 3577
rect 2401 3574 2439 3577
rect 345 3533 2439 3574
rect 3843 3574 3881 3577
rect 3933 3574 4092 3577
rect 4144 3574 4304 3577
rect 4356 3574 4515 3626
rect 4567 3574 4605 3626
rect 3843 3540 4605 3574
rect 3844 3533 4605 3540
rect 4779 3660 5961 3667
rect 4779 3626 6555 3660
rect 4779 3574 4817 3626
rect 4869 3574 5027 3626
rect 5079 3574 5238 3626
rect 5290 3574 5450 3626
rect 5502 3574 5661 3626
rect 5713 3574 5871 3626
rect 5923 3623 6555 3626
rect 5923 3577 6086 3623
rect 6320 3577 6555 3623
rect 5923 3574 6555 3577
rect 4779 3540 6555 3574
rect 7543 3626 8439 3667
rect 7543 3623 7927 3626
rect 7979 3623 8138 3626
rect 7543 3577 7554 3623
rect 8070 3577 8138 3623
rect 7543 3574 7927 3577
rect 7979 3574 8138 3577
rect 8190 3574 8349 3626
rect 8401 3574 8439 3626
rect 4779 3533 5961 3540
rect 7543 3533 8439 3574
rect 8611 3626 8920 4112
rect 8611 3574 8649 3626
rect 8701 3623 8829 3626
rect 8705 3577 8817 3623
rect 8701 3574 8829 3577
rect 8881 3574 8920 3626
rect 345 3499 637 3533
rect 345 3453 452 3499
rect 498 3453 637 3499
rect 345 3335 637 3453
rect 3081 3457 3149 3468
rect 2616 3402 2924 3443
rect 2616 3399 2654 3402
rect 2706 3399 2834 3402
rect 2886 3399 2924 3402
rect 933 3353 946 3399
rect 2920 3353 2933 3399
rect 345 3289 452 3335
rect 498 3289 637 3335
rect 2616 3350 2654 3353
rect 2706 3350 2834 3353
rect 2886 3350 2924 3353
rect 2616 3310 2924 3350
rect 345 3197 637 3289
rect 345 3175 1090 3197
rect 345 3172 946 3175
rect 345 3126 452 3172
rect 498 3129 946 3172
rect 2920 3129 2933 3175
rect 498 3126 1090 3129
rect 345 3078 1090 3126
rect 345 3009 637 3078
rect 345 2963 452 3009
rect 498 2963 637 3009
rect 3081 3035 3092 3457
rect 3138 3035 3149 3457
rect 3378 3410 3686 3451
rect 3378 3399 3416 3410
rect 3468 3399 3596 3410
rect 3648 3399 3686 3410
rect 3268 3353 3281 3399
rect 3327 3353 3384 3399
rect 3468 3358 3487 3399
rect 3430 3353 3487 3358
rect 3533 3353 3590 3399
rect 3648 3358 3693 3399
rect 3636 3353 3693 3358
rect 3739 3353 3796 3399
rect 3842 3353 3899 3399
rect 3945 3353 4002 3399
rect 4048 3353 4105 3399
rect 4151 3353 4209 3399
rect 4255 3353 4268 3399
rect 3378 3318 3686 3353
rect 4891 3324 5863 3364
rect 7450 3361 7758 3377
rect 4891 3312 4929 3324
rect 4981 3312 5140 3324
rect 5192 3312 5351 3324
rect 5403 3312 5562 3324
rect 5614 3312 5773 3324
rect 5825 3312 5863 3324
rect 6035 3312 6550 3361
rect 7036 3336 7758 3361
rect 7036 3312 7488 3336
rect 7540 3312 7668 3336
rect 7720 3312 7758 3336
rect 4857 3266 4870 3312
rect 5120 3272 5140 3312
rect 5120 3266 5177 3272
rect 5223 3266 5280 3312
rect 5326 3272 5351 3312
rect 5326 3266 5383 3272
rect 5429 3266 5486 3312
rect 5532 3272 5562 3312
rect 5532 3266 5589 3272
rect 5635 3266 5692 3312
rect 5738 3272 5773 3312
rect 5738 3266 5795 3272
rect 5841 3266 5898 3312
rect 5944 3266 5957 3312
rect 6035 3266 6451 3312
rect 6497 3266 6568 3312
rect 6614 3266 6685 3312
rect 6731 3266 6803 3312
rect 6849 3266 6921 3312
rect 6967 3266 7039 3312
rect 7085 3284 7488 3312
rect 7085 3266 7506 3284
rect 7552 3266 7623 3312
rect 7720 3284 7740 3312
rect 7669 3266 7740 3284
rect 7786 3266 7858 3312
rect 7904 3266 7976 3312
rect 8022 3266 8094 3312
rect 8140 3266 8153 3312
rect 4891 3232 5863 3266
rect 6035 3241 6550 3266
rect 7036 3244 7758 3266
rect 7036 3241 7528 3244
rect 3825 3175 4315 3204
rect 3268 3129 3281 3175
rect 3327 3129 3384 3175
rect 3430 3129 3487 3175
rect 3533 3129 3590 3175
rect 3636 3129 3693 3175
rect 3739 3129 3796 3175
rect 3842 3164 3899 3175
rect 3842 3129 3864 3164
rect 3945 3129 4002 3175
rect 4048 3164 4105 3175
rect 4096 3129 4105 3164
rect 4151 3129 4209 3175
rect 4255 3164 4315 3175
rect 3825 3112 3864 3129
rect 3916 3112 4044 3129
rect 4096 3112 4224 3129
rect 4276 3112 4315 3164
rect 6035 3138 6151 3241
rect 3825 3071 4315 3112
rect 4561 3088 5957 3132
rect 345 2846 637 2963
rect 2616 2954 2924 2995
rect 2616 2951 2654 2954
rect 2706 2951 2834 2954
rect 2886 2951 2924 2954
rect 3081 2953 3149 3035
rect 4561 3042 4870 3088
rect 5120 3042 5177 3088
rect 5223 3042 5280 3088
rect 5326 3042 5383 3088
rect 5429 3042 5486 3088
rect 5532 3042 5589 3088
rect 5635 3042 5692 3088
rect 5738 3042 5795 3088
rect 5841 3042 5898 3088
rect 5944 3042 5957 3088
rect 4561 3010 5957 3042
rect 4561 2953 4679 3010
rect 933 2905 946 2951
rect 2920 2905 2933 2951
rect 3081 2916 4679 2953
rect 2616 2902 2654 2905
rect 2706 2902 2834 2905
rect 2886 2902 2924 2905
rect 2616 2862 2924 2902
rect 3081 2870 3413 2916
rect 3459 2870 3599 2916
rect 3645 2870 3786 2916
rect 3832 2870 3973 2916
rect 4019 2870 4159 2916
rect 4205 2870 4679 2916
rect 6035 2998 6072 3138
rect 6118 2998 6151 3138
rect 3081 2862 4679 2870
rect 4891 2864 5863 2904
rect 6035 2898 6151 2998
rect 6237 3138 6370 3161
rect 6237 3089 6294 3138
rect 6237 3037 6275 3089
rect 6237 2998 6294 3037
rect 6340 2998 6370 3138
rect 8255 3140 8323 3151
rect 6521 3130 7282 3136
rect 6520 3129 7282 3130
rect 6520 3096 7528 3129
rect 6520 3088 6558 3096
rect 6610 3088 6769 3096
rect 6821 3088 6981 3096
rect 6438 3042 6451 3088
rect 6497 3044 6558 3088
rect 6497 3042 6568 3044
rect 6614 3042 6685 3088
rect 6731 3044 6769 3088
rect 6731 3042 6803 3044
rect 6849 3042 6921 3088
rect 6967 3044 6981 3088
rect 7033 3088 7192 3096
rect 7033 3044 7039 3088
rect 6967 3042 7039 3044
rect 7085 3044 7192 3088
rect 7244 3088 7528 3096
rect 7244 3044 7506 3088
rect 7085 3042 7506 3044
rect 7552 3042 7623 3088
rect 7669 3042 7740 3088
rect 7786 3042 7858 3088
rect 7904 3042 7976 3088
rect 8022 3042 8094 3088
rect 8140 3042 8153 3088
rect 6520 3010 7528 3042
rect 6521 3003 7282 3010
rect 6237 2978 6370 2998
rect 8255 3000 8266 3140
rect 8312 3000 8323 3140
rect 8611 3088 8920 3574
rect 9089 3660 9205 4112
rect 9520 4079 9682 4210
rect 9520 4027 9591 4079
rect 9643 4027 9682 4079
rect 9520 3987 9682 4027
rect 9334 3891 9462 3904
rect 9334 3864 9463 3891
rect 9334 3847 9372 3864
rect 9424 3847 9463 3864
rect 9324 3801 9337 3847
rect 9424 3812 9459 3847
rect 9383 3801 9459 3812
rect 9505 3801 9582 3847
rect 9628 3801 9705 3847
rect 9751 3801 9764 3847
rect 9843 3836 9959 4234
rect 11826 4095 14106 4136
rect 11826 4043 13042 4095
rect 13094 4043 14106 4095
rect 11826 4003 14106 4043
rect 13938 3959 14106 4003
rect 13938 3913 13955 3959
rect 14095 3913 14106 3959
rect 9334 3772 9463 3801
rect 9843 3790 9878 3836
rect 9924 3790 9959 3836
rect 9843 3753 9959 3790
rect 10315 3864 13121 3905
rect 13938 3902 14106 3913
rect 10315 3812 11532 3864
rect 11584 3812 13121 3864
rect 10315 3771 13121 3812
rect 14202 3847 14318 4234
rect 14997 4204 17976 4245
rect 14997 4190 16328 4204
rect 14997 4144 15061 4190
rect 15201 4152 16328 4190
rect 16380 4152 17976 4204
rect 15201 4144 17976 4152
rect 14498 4088 14838 4129
rect 14997 4111 17976 4144
rect 18154 4198 18193 4250
rect 18245 4198 18284 4250
rect 18154 4175 18284 4198
rect 19641 4284 20113 4330
rect 20159 4284 20300 4330
rect 20346 4284 20487 4330
rect 20533 4284 20673 4330
rect 20719 4284 20860 4330
rect 20906 4284 21254 4330
rect 21394 4320 21702 4360
rect 21394 4295 21432 4320
rect 21484 4295 21612 4320
rect 21664 4295 21702 4320
rect 23682 4354 23820 4400
rect 23866 4354 23974 4400
rect 19641 4247 21254 4284
rect 21386 4249 21399 4295
rect 23373 4249 23386 4295
rect 19641 4190 19757 4247
rect 14498 4071 14536 4088
rect 14588 4071 14748 4088
rect 14800 4071 14838 4088
rect 14396 4025 14409 4071
rect 14455 4025 14522 4071
rect 14588 4036 14635 4071
rect 14568 4025 14635 4036
rect 14681 4025 14748 4071
rect 14800 4036 14861 4071
rect 14794 4025 14861 4036
rect 14907 4025 14920 4071
rect 18154 4035 18219 4175
rect 18265 4035 18284 4175
rect 19417 4158 19757 4190
rect 18362 4112 18375 4158
rect 18421 4112 18478 4158
rect 18524 4112 18581 4158
rect 18627 4112 18684 4158
rect 18730 4112 18787 4158
rect 18833 4112 18890 4158
rect 18936 4112 18993 4158
rect 19039 4112 19096 4158
rect 19142 4112 19199 4158
rect 19449 4112 19757 4158
rect 21186 4195 21254 4247
rect 21394 4227 21702 4249
rect 19417 4071 19757 4112
rect 19859 4088 20409 4129
rect 18154 4032 18284 4035
rect 14498 3996 14838 4025
rect 18154 3980 18193 4032
rect 18245 3980 18284 4032
rect 19859 4036 19897 4088
rect 19949 4071 20108 4088
rect 20160 4071 20319 4088
rect 19949 4036 20064 4071
rect 20160 4036 20168 4071
rect 19859 4025 20064 4036
rect 20110 4025 20168 4036
rect 20214 4025 20271 4071
rect 20317 4036 20319 4071
rect 20371 4071 20409 4088
rect 20371 4036 20374 4071
rect 20317 4025 20374 4036
rect 20420 4025 20477 4071
rect 20523 4025 20580 4071
rect 20626 4025 20683 4071
rect 20729 4025 20786 4071
rect 20832 4025 20889 4071
rect 20935 4025 20992 4071
rect 21038 4025 21051 4071
rect 19859 3996 20409 4025
rect 18154 3939 18284 3980
rect 18502 3934 19474 3965
rect 18362 3888 18375 3934
rect 18421 3888 18478 3934
rect 18524 3925 18581 3934
rect 18524 3888 18540 3925
rect 18627 3888 18684 3934
rect 18730 3925 18787 3934
rect 18730 3888 18751 3925
rect 18833 3888 18890 3934
rect 18936 3925 18993 3934
rect 18936 3888 18962 3925
rect 19039 3888 19096 3934
rect 19142 3925 19199 3934
rect 19142 3888 19173 3925
rect 19449 3888 19474 3934
rect 18502 3873 18540 3888
rect 18592 3873 18751 3888
rect 18803 3873 18962 3888
rect 19014 3873 19173 3888
rect 19225 3873 19384 3888
rect 19436 3873 19474 3888
rect 14202 3801 14409 3847
rect 14455 3801 14522 3847
rect 14568 3801 14635 3847
rect 14681 3801 14748 3847
rect 14794 3801 14861 3847
rect 14907 3801 14920 3847
rect 18502 3833 19474 3873
rect 20632 3850 20940 3890
rect 20632 3847 20670 3850
rect 20722 3847 20850 3850
rect 20902 3847 20940 3850
rect 12959 3764 13121 3771
rect 12959 3718 12970 3764
rect 13110 3718 13121 3764
rect 12959 3707 13121 3718
rect 15181 3787 18143 3823
rect 20051 3801 20064 3847
rect 20110 3801 20168 3847
rect 20214 3801 20271 3847
rect 20317 3801 20374 3847
rect 20420 3801 20477 3847
rect 20523 3801 20580 3847
rect 20626 3801 20670 3847
rect 20729 3801 20786 3847
rect 20832 3801 20850 3847
rect 20935 3801 20992 3847
rect 21038 3801 21051 3847
rect 15181 3741 15216 3787
rect 15262 3741 15374 3787
rect 15420 3741 15532 3787
rect 15578 3741 15690 3787
rect 15736 3741 15848 3787
rect 15894 3741 16006 3787
rect 16052 3741 16165 3787
rect 16211 3741 16323 3787
rect 16369 3741 16481 3787
rect 16527 3741 16639 3787
rect 16685 3741 16797 3787
rect 16843 3741 16955 3787
rect 17001 3741 17113 3787
rect 17159 3741 17272 3787
rect 17318 3741 17430 3787
rect 17476 3741 17588 3787
rect 17634 3741 17746 3787
rect 17792 3741 17904 3787
rect 17950 3741 18062 3787
rect 18108 3741 18143 3787
rect 20632 3798 20670 3801
rect 20722 3798 20850 3801
rect 20902 3798 20940 3801
rect 20632 3757 20940 3798
rect 21186 3773 21197 4195
rect 21243 3773 21254 4195
rect 23682 4122 23974 4354
rect 23182 4071 23974 4122
rect 21386 4025 21399 4071
rect 23373 4025 23974 4071
rect 23182 4003 23974 4025
rect 23682 3911 23974 4003
rect 21394 3857 21702 3897
rect 21394 3847 21432 3857
rect 21484 3847 21612 3857
rect 21664 3847 21702 3857
rect 23682 3865 23820 3911
rect 23866 3865 23974 3911
rect 21386 3801 21399 3847
rect 23373 3801 23386 3847
rect 21186 3762 21254 3773
rect 21394 3764 21702 3801
rect 9812 3660 10120 3667
rect 10385 3660 12583 3674
rect 13350 3660 14111 3667
rect 9089 3637 12583 3660
rect 13301 3637 14111 3660
rect 9089 3626 14111 3637
rect 9089 3623 9850 3626
rect 9089 3577 9337 3623
rect 9383 3577 9459 3623
rect 9505 3577 9582 3623
rect 9628 3577 9705 3623
rect 9751 3577 9850 3623
rect 9089 3574 9850 3577
rect 9902 3574 10030 3626
rect 10082 3623 13387 3626
rect 10082 3577 10433 3623
rect 10479 3577 10591 3623
rect 10637 3577 10749 3623
rect 10795 3577 10907 3623
rect 10953 3577 11066 3623
rect 11112 3577 11224 3623
rect 11270 3577 11382 3623
rect 11428 3577 11540 3623
rect 11586 3577 11698 3623
rect 11744 3577 11856 3623
rect 11902 3577 12015 3623
rect 12061 3577 12173 3623
rect 12219 3577 12331 3623
rect 12377 3577 12489 3623
rect 12535 3577 13336 3623
rect 13382 3577 13387 3623
rect 10082 3574 13387 3577
rect 13439 3623 13598 3626
rect 13439 3577 13503 3623
rect 13549 3577 13598 3623
rect 13439 3574 13598 3577
rect 13650 3623 13810 3626
rect 13862 3623 14021 3626
rect 13650 3577 13668 3623
rect 13714 3577 13810 3623
rect 13879 3577 14021 3623
rect 13650 3574 13810 3577
rect 13862 3574 14021 3577
rect 14073 3574 14111 3626
rect 9089 3563 14111 3574
rect 9089 3540 12583 3563
rect 13301 3540 14111 3563
rect 9089 3088 9205 3540
rect 9812 3533 10120 3540
rect 10385 3526 12583 3540
rect 13350 3533 14111 3540
rect 14393 3660 14943 3667
rect 15181 3660 18143 3741
rect 23682 3747 23974 3865
rect 23682 3701 23820 3747
rect 23866 3701 23974 3747
rect 23682 3667 23974 3701
rect 18397 3660 19579 3667
rect 19905 3660 20456 3667
rect 14393 3626 19579 3660
rect 14393 3623 14431 3626
rect 14483 3623 14642 3626
rect 14694 3623 14853 3626
rect 14905 3623 18435 3626
rect 14393 3577 14409 3623
rect 14483 3577 14522 3623
rect 14568 3577 14635 3623
rect 14694 3577 14748 3623
rect 14794 3577 14853 3623
rect 14907 3577 15216 3623
rect 15262 3577 15374 3623
rect 15420 3577 15532 3623
rect 15578 3577 15690 3623
rect 15736 3577 15848 3623
rect 15894 3577 16006 3623
rect 16052 3577 16165 3623
rect 16211 3577 16323 3623
rect 16369 3577 16481 3623
rect 16527 3577 16639 3623
rect 16685 3577 16797 3623
rect 16843 3577 16955 3623
rect 17001 3577 17113 3623
rect 17159 3577 17272 3623
rect 17318 3577 17430 3623
rect 17476 3577 17588 3623
rect 17634 3577 17746 3623
rect 17792 3577 17904 3623
rect 17950 3577 18062 3623
rect 18108 3577 18435 3623
rect 14393 3574 14431 3577
rect 14483 3574 14642 3577
rect 14694 3574 14853 3577
rect 14905 3574 18435 3577
rect 18487 3574 18645 3626
rect 18697 3574 18856 3626
rect 18908 3574 19068 3626
rect 19120 3574 19279 3626
rect 19331 3574 19489 3626
rect 19541 3574 19579 3626
rect 14393 3540 19579 3574
rect 19904 3626 20456 3660
rect 19904 3574 19943 3626
rect 19995 3623 20154 3626
rect 20206 3623 20365 3626
rect 20417 3623 20456 3626
rect 21875 3626 23974 3667
rect 21875 3623 21913 3626
rect 21965 3623 22124 3626
rect 22176 3623 22335 3626
rect 22387 3623 22545 3626
rect 22597 3623 22756 3626
rect 22808 3623 22968 3626
rect 23020 3623 23179 3626
rect 23231 3623 23389 3626
rect 19995 3577 20064 3623
rect 20110 3577 20154 3623
rect 20214 3577 20271 3623
rect 20317 3577 20365 3623
rect 20420 3577 20477 3623
rect 20523 3577 20580 3623
rect 20626 3577 20683 3623
rect 20729 3577 20786 3623
rect 20832 3577 20889 3623
rect 20935 3577 20992 3623
rect 21038 3577 21051 3623
rect 21386 3577 21399 3623
rect 23373 3577 23389 3623
rect 19995 3574 20154 3577
rect 20206 3574 20365 3577
rect 20417 3574 20456 3577
rect 19904 3540 20456 3574
rect 14393 3533 14943 3540
rect 12959 3482 13121 3493
rect 9334 3399 9463 3428
rect 9843 3410 9959 3447
rect 12959 3436 12970 3482
rect 13110 3436 13121 3482
rect 12959 3429 13121 3436
rect 9324 3353 9337 3399
rect 9383 3388 9459 3399
rect 9424 3353 9459 3388
rect 9505 3353 9582 3399
rect 9628 3353 9705 3399
rect 9751 3353 9764 3399
rect 9843 3364 9878 3410
rect 9924 3364 9959 3410
rect 9334 3336 9372 3353
rect 9424 3336 9463 3353
rect 9334 3309 9463 3336
rect 9334 3296 9462 3309
rect 9520 3173 9682 3213
rect 9520 3121 9591 3173
rect 9643 3121 9682 3173
rect 8605 3042 8618 3088
rect 8664 3042 8741 3088
rect 8787 3042 8864 3088
rect 8910 3042 8923 3088
rect 9089 3042 9238 3088
rect 9284 3042 9327 3088
rect 8611 3010 8920 3042
rect 9089 3010 9205 3042
rect 7450 2898 7758 2903
rect 6035 2864 6550 2898
rect 7036 2864 7758 2898
rect 8255 2878 8323 3000
rect 9520 2990 9682 3121
rect 9406 2987 9682 2990
rect 9406 2979 9591 2987
rect 9406 2933 9441 2979
rect 9487 2935 9591 2979
rect 9643 2966 9682 2987
rect 9843 2966 9959 3364
rect 10315 3388 13121 3429
rect 15181 3459 18143 3540
rect 18397 3533 19579 3540
rect 19905 3533 20456 3540
rect 21875 3574 21913 3577
rect 21965 3574 22124 3577
rect 22176 3574 22335 3577
rect 22387 3574 22545 3577
rect 22597 3574 22756 3577
rect 22808 3574 22968 3577
rect 23020 3574 23179 3577
rect 23231 3574 23389 3577
rect 23441 3574 23600 3626
rect 23652 3574 23811 3626
rect 23863 3574 23974 3626
rect 21875 3533 23974 3574
rect 15181 3413 15216 3459
rect 15262 3413 15374 3459
rect 15420 3413 15532 3459
rect 15578 3413 15690 3459
rect 15736 3413 15848 3459
rect 15894 3413 16006 3459
rect 16052 3413 16165 3459
rect 16211 3413 16323 3459
rect 16369 3413 16481 3459
rect 16527 3413 16639 3459
rect 16685 3413 16797 3459
rect 16843 3413 16955 3459
rect 17001 3413 17113 3459
rect 17159 3413 17272 3459
rect 17318 3413 17430 3459
rect 17476 3413 17588 3459
rect 17634 3413 17746 3459
rect 17792 3413 17904 3459
rect 17950 3413 18062 3459
rect 18108 3413 18143 3459
rect 23682 3499 23974 3533
rect 23682 3453 23820 3499
rect 23866 3453 23974 3499
rect 10315 3336 11532 3388
rect 11584 3336 13121 3388
rect 10315 3295 13121 3336
rect 14202 3353 14409 3399
rect 14455 3353 14522 3399
rect 14568 3353 14635 3399
rect 14681 3353 14748 3399
rect 14794 3353 14861 3399
rect 14907 3353 14920 3399
rect 15181 3377 18143 3413
rect 20632 3402 20940 3443
rect 20632 3399 20670 3402
rect 20722 3399 20850 3402
rect 20902 3399 20940 3402
rect 21186 3427 21254 3438
rect 13938 3287 14106 3298
rect 13938 3241 13955 3287
rect 14095 3241 14106 3287
rect 13938 3197 14106 3241
rect 11826 3157 14106 3197
rect 11826 3105 13042 3157
rect 13094 3105 14106 3157
rect 11826 3064 14106 3105
rect 14202 2966 14318 3353
rect 18502 3327 19474 3367
rect 20051 3353 20064 3399
rect 20110 3353 20168 3399
rect 20214 3353 20271 3399
rect 20317 3353 20374 3399
rect 20420 3353 20477 3399
rect 20523 3353 20580 3399
rect 20626 3353 20670 3399
rect 20729 3353 20786 3399
rect 20832 3353 20850 3399
rect 20935 3353 20992 3399
rect 21038 3353 21051 3399
rect 18502 3312 18540 3327
rect 18592 3312 18751 3327
rect 18803 3312 18962 3327
rect 19014 3312 19173 3327
rect 19225 3312 19384 3327
rect 19436 3312 19474 3327
rect 18362 3266 18375 3312
rect 18421 3266 18478 3312
rect 18524 3275 18540 3312
rect 18524 3266 18581 3275
rect 18627 3266 18684 3312
rect 18730 3275 18751 3312
rect 18730 3266 18787 3275
rect 18833 3266 18890 3312
rect 18936 3275 18962 3312
rect 18936 3266 18993 3275
rect 19039 3266 19096 3312
rect 19142 3275 19173 3312
rect 19142 3266 19199 3275
rect 19449 3266 19474 3312
rect 20632 3350 20670 3353
rect 20722 3350 20850 3353
rect 20902 3350 20940 3353
rect 20632 3310 20940 3350
rect 18154 3220 18284 3261
rect 18502 3235 19474 3266
rect 14498 3175 14838 3204
rect 14396 3129 14409 3175
rect 14455 3129 14522 3175
rect 14568 3164 14635 3175
rect 14588 3129 14635 3164
rect 14681 3129 14748 3175
rect 14794 3164 14861 3175
rect 14800 3129 14861 3164
rect 14907 3129 14920 3175
rect 18154 3168 18193 3220
rect 18245 3168 18284 3220
rect 18154 3165 18284 3168
rect 14498 3112 14536 3129
rect 14588 3112 14748 3129
rect 14800 3112 14838 3129
rect 14498 3071 14838 3112
rect 14997 3056 17976 3089
rect 14997 3010 15061 3056
rect 15201 3048 17976 3056
rect 15201 3010 16705 3048
rect 14997 2996 16705 3010
rect 16757 2996 17976 3048
rect 9643 2951 14515 2966
rect 14997 2955 17976 2996
rect 18154 3025 18219 3165
rect 18265 3025 18284 3165
rect 19859 3175 20409 3204
rect 19859 3164 20064 3175
rect 20110 3164 20168 3175
rect 19417 3088 19757 3129
rect 18362 3042 18375 3088
rect 18421 3042 18478 3088
rect 18524 3042 18581 3088
rect 18627 3042 18684 3088
rect 18730 3042 18787 3088
rect 18833 3042 18890 3088
rect 18936 3042 18993 3088
rect 19039 3042 19096 3088
rect 19142 3042 19199 3088
rect 19449 3042 19757 3088
rect 19859 3112 19897 3164
rect 19949 3129 20064 3164
rect 20160 3129 20168 3164
rect 20214 3129 20271 3175
rect 20317 3164 20374 3175
rect 20317 3129 20319 3164
rect 19949 3112 20108 3129
rect 20160 3112 20319 3129
rect 20371 3129 20374 3164
rect 20420 3129 20477 3175
rect 20523 3129 20580 3175
rect 20626 3129 20683 3175
rect 20729 3129 20786 3175
rect 20832 3129 20889 3175
rect 20935 3129 20992 3175
rect 21038 3129 21051 3175
rect 20371 3112 20409 3129
rect 19859 3071 20409 3112
rect 18154 3002 18284 3025
rect 19417 3010 19757 3042
rect 9643 2935 14409 2951
rect 9487 2933 14409 2935
rect 9406 2930 14409 2933
rect 9406 2884 13336 2930
rect 13382 2884 13503 2930
rect 13549 2884 13668 2930
rect 13714 2884 13833 2930
rect 13879 2905 14409 2930
rect 14455 2905 14522 2951
rect 14568 2905 14635 2951
rect 14681 2905 14748 2951
rect 14794 2905 14861 2951
rect 14907 2905 14920 2951
rect 18154 2950 18193 3002
rect 18245 2950 18284 3002
rect 18154 2910 18284 2950
rect 19641 2953 19757 3010
rect 21186 3005 21197 3427
rect 21243 3005 21254 3427
rect 21394 3399 21702 3436
rect 21386 3353 21399 3399
rect 23373 3353 23386 3399
rect 21394 3343 21432 3353
rect 21484 3343 21612 3353
rect 21664 3343 21702 3353
rect 21394 3303 21702 3343
rect 23682 3335 23974 3453
rect 23682 3289 23820 3335
rect 23866 3289 23974 3335
rect 23682 3197 23974 3289
rect 23182 3175 23974 3197
rect 21386 3129 21399 3175
rect 23373 3129 23974 3175
rect 23182 3078 23974 3129
rect 21186 2953 21254 3005
rect 19641 2916 21254 2953
rect 21394 2951 21702 2973
rect 13879 2884 14515 2905
rect 8255 2864 9320 2878
rect 345 2800 452 2846
rect 498 2800 637 2846
rect 3081 2833 4240 2862
rect 4857 2818 4870 2864
rect 5120 2818 5140 2864
rect 5223 2818 5280 2864
rect 5326 2818 5351 2864
rect 5429 2818 5486 2864
rect 5532 2818 5562 2864
rect 5635 2818 5692 2864
rect 5738 2818 5773 2864
rect 5841 2818 5898 2864
rect 5944 2818 5957 2864
rect 6035 2818 6451 2864
rect 6497 2818 6568 2864
rect 6614 2818 6685 2864
rect 6731 2818 6803 2864
rect 6849 2818 6921 2864
rect 6967 2818 7039 2864
rect 7085 2862 7506 2864
rect 7085 2818 7488 2862
rect 7552 2818 7623 2864
rect 7669 2862 7740 2864
rect 7720 2818 7740 2862
rect 7786 2818 7858 2864
rect 7904 2818 7976 2864
rect 8022 2818 8094 2864
rect 8140 2818 8153 2864
rect 8255 2818 8618 2864
rect 8664 2818 8741 2864
rect 8787 2818 8864 2864
rect 8910 2818 9238 2864
rect 9284 2818 9327 2864
rect 9406 2846 14515 2884
rect 18502 2864 19474 2904
rect 18362 2818 18375 2864
rect 18421 2818 18478 2864
rect 18524 2818 18540 2864
rect 18627 2818 18684 2864
rect 18730 2818 18751 2864
rect 18833 2818 18890 2864
rect 18936 2818 18962 2864
rect 19039 2818 19096 2864
rect 19142 2818 19173 2864
rect 19449 2818 19474 2864
rect 19641 2870 20113 2916
rect 20159 2870 20300 2916
rect 20346 2870 20487 2916
rect 20533 2870 20673 2916
rect 20719 2870 20860 2916
rect 20906 2870 21254 2916
rect 21386 2905 21399 2951
rect 23373 2905 23386 2951
rect 19641 2860 21254 2870
rect 20078 2833 21254 2860
rect 21394 2880 21432 2905
rect 21484 2880 21612 2905
rect 21664 2880 21702 2905
rect 21394 2840 21702 2880
rect 23682 2846 23974 3078
rect 345 2767 637 2800
rect 4891 2812 4929 2818
rect 4981 2812 5140 2818
rect 5192 2812 5351 2818
rect 5403 2812 5562 2818
rect 5614 2812 5773 2818
rect 5825 2812 5863 2818
rect 4467 2767 4622 2774
rect 4891 2772 5863 2812
rect 6035 2778 6550 2818
rect 7036 2810 7488 2818
rect 7540 2810 7668 2818
rect 7720 2810 7758 2818
rect 7036 2778 7758 2810
rect 7450 2770 7758 2778
rect 345 2726 2439 2767
rect 345 2674 451 2726
rect 503 2674 662 2726
rect 714 2674 873 2726
rect 925 2674 1083 2726
rect 1135 2674 1294 2726
rect 1346 2674 1506 2726
rect 1558 2674 1717 2726
rect 1769 2674 1927 2726
rect 1979 2674 2138 2726
rect 2190 2674 2349 2726
rect 2401 2674 2439 2726
rect 345 2633 2439 2674
rect 4314 2726 4622 2767
rect 8255 2758 9320 2818
rect 18502 2812 18540 2818
rect 18592 2812 18751 2818
rect 18803 2812 18962 2818
rect 19014 2812 19173 2818
rect 19225 2812 19384 2818
rect 19436 2812 19474 2818
rect 18502 2772 19474 2812
rect 23682 2800 23820 2846
rect 23866 2800 23974 2846
rect 19696 2767 19852 2774
rect 23682 2767 23974 2800
rect 4314 2674 4352 2726
rect 4404 2723 4532 2726
rect 4404 2677 4513 2723
rect 4404 2674 4532 2677
rect 4584 2674 4622 2726
rect 4314 2633 4622 2674
rect 19696 2726 20005 2767
rect 19696 2674 19735 2726
rect 19787 2723 19915 2726
rect 19803 2677 19915 2723
rect 19787 2674 19915 2677
rect 19967 2674 20005 2726
rect 345 2600 637 2633
rect 4467 2626 4622 2633
rect 345 2554 452 2600
rect 498 2554 637 2600
rect 4891 2588 5863 2628
rect 7450 2622 7758 2630
rect 4891 2582 4929 2588
rect 4981 2582 5140 2588
rect 5192 2582 5351 2588
rect 5403 2582 5562 2588
rect 5614 2582 5773 2588
rect 5825 2582 5863 2588
rect 6035 2582 6550 2622
rect 7036 2590 7758 2622
rect 7036 2582 7488 2590
rect 7540 2582 7668 2590
rect 7720 2582 7758 2590
rect 8255 2582 9320 2642
rect 19696 2633 20005 2674
rect 21875 2726 23974 2767
rect 21875 2674 21913 2726
rect 21965 2674 22124 2726
rect 22176 2674 22335 2726
rect 22387 2674 22545 2726
rect 22597 2674 22756 2726
rect 22808 2674 22968 2726
rect 23020 2674 23179 2726
rect 23231 2674 23389 2726
rect 23441 2674 23600 2726
rect 23652 2674 23811 2726
rect 23863 2674 23974 2726
rect 21875 2633 23974 2674
rect 18502 2588 19474 2628
rect 19696 2626 19852 2633
rect 18502 2582 18540 2588
rect 18592 2582 18751 2588
rect 18803 2582 18962 2588
rect 19014 2582 19173 2588
rect 19225 2582 19384 2588
rect 19436 2582 19474 2588
rect 345 2437 637 2554
rect 3081 2538 4240 2567
rect 2616 2498 2924 2538
rect 2616 2495 2654 2498
rect 2706 2495 2834 2498
rect 2886 2495 2924 2498
rect 3081 2530 4679 2538
rect 4857 2536 4870 2582
rect 5120 2536 5140 2582
rect 5223 2536 5280 2582
rect 5326 2536 5351 2582
rect 5429 2536 5486 2582
rect 5532 2536 5562 2582
rect 5635 2536 5692 2582
rect 5738 2536 5773 2582
rect 5841 2536 5898 2582
rect 5944 2536 5957 2582
rect 6035 2536 6451 2582
rect 6497 2536 6568 2582
rect 6614 2536 6685 2582
rect 6731 2536 6803 2582
rect 6849 2536 6921 2582
rect 6967 2536 7039 2582
rect 7085 2538 7488 2582
rect 7085 2536 7506 2538
rect 7552 2536 7623 2582
rect 7720 2538 7740 2582
rect 7669 2536 7740 2538
rect 7786 2536 7858 2582
rect 7904 2536 7976 2582
rect 8022 2536 8094 2582
rect 8140 2536 8153 2582
rect 8255 2536 8618 2582
rect 8664 2536 8741 2582
rect 8787 2536 8864 2582
rect 8910 2536 9238 2582
rect 9284 2536 9327 2582
rect 933 2449 946 2495
rect 2920 2449 2933 2495
rect 3081 2484 3413 2530
rect 3459 2484 3599 2530
rect 3645 2484 3786 2530
rect 3832 2484 3973 2530
rect 4019 2484 4159 2530
rect 4205 2484 4679 2530
rect 4891 2496 5863 2536
rect 6035 2502 6550 2536
rect 7036 2502 7758 2536
rect 345 2391 452 2437
rect 498 2391 637 2437
rect 2616 2446 2654 2449
rect 2706 2446 2834 2449
rect 2886 2446 2924 2449
rect 2616 2405 2924 2446
rect 3081 2447 4679 2484
rect 345 2322 637 2391
rect 3081 2365 3149 2447
rect 345 2274 1090 2322
rect 345 2228 452 2274
rect 498 2271 1090 2274
rect 498 2228 946 2271
rect 345 2225 946 2228
rect 2920 2225 2933 2271
rect 345 2203 1090 2225
rect 345 2111 637 2203
rect 345 2065 452 2111
rect 498 2065 637 2111
rect 345 1947 637 2065
rect 2616 2050 2924 2090
rect 2616 2047 2654 2050
rect 2706 2047 2834 2050
rect 2886 2047 2924 2050
rect 933 2001 946 2047
rect 2920 2001 2933 2047
rect 2616 1998 2654 2001
rect 2706 1998 2834 2001
rect 2886 1998 2924 2001
rect 2616 1957 2924 1998
rect 345 1901 452 1947
rect 498 1901 637 1947
rect 3081 1943 3092 2365
rect 3138 1943 3149 2365
rect 4561 2390 4679 2447
rect 6035 2402 6151 2502
rect 7450 2497 7758 2502
rect 8255 2522 9320 2536
rect 4561 2358 5957 2390
rect 3825 2288 4315 2329
rect 3825 2271 3864 2288
rect 3916 2271 4044 2288
rect 4096 2271 4224 2288
rect 3268 2225 3281 2271
rect 3327 2225 3384 2271
rect 3430 2225 3487 2271
rect 3533 2225 3590 2271
rect 3636 2225 3693 2271
rect 3739 2225 3796 2271
rect 3842 2236 3864 2271
rect 3842 2225 3899 2236
rect 3945 2225 4002 2271
rect 4096 2236 4105 2271
rect 4048 2225 4105 2236
rect 4151 2225 4209 2271
rect 4276 2236 4315 2288
rect 4561 2312 4870 2358
rect 5120 2312 5177 2358
rect 5223 2312 5280 2358
rect 5326 2312 5383 2358
rect 5429 2312 5486 2358
rect 5532 2312 5589 2358
rect 5635 2312 5692 2358
rect 5738 2312 5795 2358
rect 5841 2312 5898 2358
rect 5944 2312 5957 2358
rect 4561 2268 5957 2312
rect 4255 2225 4315 2236
rect 3825 2196 4315 2225
rect 6035 2262 6072 2402
rect 6118 2262 6151 2402
rect 4891 2134 5863 2168
rect 6035 2159 6151 2262
rect 6237 2402 6370 2422
rect 6237 2363 6294 2402
rect 6237 2311 6275 2363
rect 6237 2262 6294 2311
rect 6340 2262 6370 2402
rect 8255 2400 8323 2522
rect 9406 2516 14515 2554
rect 18362 2536 18375 2582
rect 18421 2536 18478 2582
rect 18524 2536 18540 2582
rect 18627 2536 18684 2582
rect 18730 2536 18751 2582
rect 18833 2536 18890 2582
rect 18936 2536 18962 2582
rect 19039 2536 19096 2582
rect 19142 2536 19173 2582
rect 19449 2536 19474 2582
rect 23682 2600 23974 2633
rect 20078 2540 21254 2567
rect 9406 2470 13336 2516
rect 13382 2470 13503 2516
rect 13549 2470 13668 2516
rect 13714 2470 13833 2516
rect 13879 2495 14515 2516
rect 18502 2496 19474 2536
rect 19641 2530 21254 2540
rect 13879 2470 14409 2495
rect 9406 2467 14409 2470
rect 9406 2421 9441 2467
rect 9487 2465 14409 2467
rect 9487 2421 9591 2465
rect 9406 2413 9591 2421
rect 9643 2449 14409 2465
rect 14455 2449 14522 2495
rect 14568 2449 14635 2495
rect 14681 2449 14748 2495
rect 14794 2449 14861 2495
rect 14907 2449 14920 2495
rect 18154 2450 18284 2490
rect 9643 2434 14515 2449
rect 9643 2413 9682 2434
rect 9406 2410 9682 2413
rect 6521 2390 7282 2397
rect 6520 2358 7528 2390
rect 6438 2312 6451 2358
rect 6497 2356 6568 2358
rect 6497 2312 6558 2356
rect 6614 2312 6685 2358
rect 6731 2356 6803 2358
rect 6731 2312 6769 2356
rect 6849 2312 6921 2358
rect 6967 2356 7039 2358
rect 6967 2312 6981 2356
rect 6520 2304 6558 2312
rect 6610 2304 6769 2312
rect 6821 2304 6981 2312
rect 7033 2312 7039 2356
rect 7085 2356 7506 2358
rect 7085 2312 7192 2356
rect 7033 2304 7192 2312
rect 7244 2312 7506 2356
rect 7552 2312 7623 2358
rect 7669 2312 7740 2358
rect 7786 2312 7858 2358
rect 7904 2312 7976 2358
rect 8022 2312 8094 2358
rect 8140 2312 8153 2358
rect 7244 2304 7528 2312
rect 6520 2271 7528 2304
rect 6520 2270 7282 2271
rect 6521 2264 7282 2270
rect 6237 2239 6370 2262
rect 8255 2260 8266 2400
rect 8312 2260 8323 2400
rect 8611 2358 8920 2390
rect 9089 2358 9205 2390
rect 8605 2312 8618 2358
rect 8664 2312 8741 2358
rect 8787 2312 8864 2358
rect 8910 2312 8923 2358
rect 9089 2312 9238 2358
rect 9284 2312 9327 2358
rect 8255 2249 8323 2260
rect 6035 2134 6550 2159
rect 7036 2156 7528 2159
rect 7036 2134 7758 2156
rect 4857 2088 4870 2134
rect 5120 2128 5177 2134
rect 5120 2088 5140 2128
rect 5223 2088 5280 2134
rect 5326 2128 5383 2134
rect 5326 2088 5351 2128
rect 5429 2088 5486 2134
rect 5532 2128 5589 2134
rect 5532 2088 5562 2128
rect 5635 2088 5692 2134
rect 5738 2128 5795 2134
rect 5738 2088 5773 2128
rect 5841 2088 5898 2134
rect 5944 2088 5957 2134
rect 6035 2088 6451 2134
rect 6497 2088 6568 2134
rect 6614 2088 6685 2134
rect 6731 2088 6803 2134
rect 6849 2088 6921 2134
rect 6967 2088 7039 2134
rect 7085 2116 7506 2134
rect 7085 2088 7488 2116
rect 7552 2088 7623 2134
rect 7669 2116 7740 2134
rect 7720 2088 7740 2116
rect 7786 2088 7858 2134
rect 7904 2088 7976 2134
rect 8022 2088 8094 2134
rect 8140 2088 8153 2134
rect 3378 2047 3686 2082
rect 4891 2076 4929 2088
rect 4981 2076 5140 2088
rect 5192 2076 5351 2088
rect 5403 2076 5562 2088
rect 5614 2076 5773 2088
rect 5825 2076 5863 2088
rect 3268 2001 3281 2047
rect 3327 2001 3384 2047
rect 3430 2042 3487 2047
rect 3468 2001 3487 2042
rect 3533 2001 3590 2047
rect 3636 2042 3693 2047
rect 3648 2001 3693 2042
rect 3739 2001 3796 2047
rect 3842 2001 3899 2047
rect 3945 2001 4002 2047
rect 4048 2001 4105 2047
rect 4151 2001 4209 2047
rect 4255 2001 4268 2047
rect 4891 2036 5863 2076
rect 6035 2039 6550 2088
rect 7036 2064 7488 2088
rect 7540 2064 7668 2088
rect 7720 2064 7758 2088
rect 7036 2039 7758 2064
rect 7450 2023 7758 2039
rect 3378 1990 3416 2001
rect 3468 1990 3596 2001
rect 3648 1990 3686 2001
rect 3378 1949 3686 1990
rect 3081 1932 3149 1943
rect 345 1867 637 1901
rect 345 1826 2439 1867
rect 3844 1860 4605 1867
rect 345 1774 451 1826
rect 503 1774 662 1826
rect 714 1774 873 1826
rect 925 1823 1083 1826
rect 1135 1823 1294 1826
rect 1346 1823 1506 1826
rect 1558 1823 1717 1826
rect 1769 1823 1927 1826
rect 1979 1823 2138 1826
rect 2190 1823 2349 1826
rect 2401 1823 2439 1826
rect 3843 1826 4605 1860
rect 3843 1823 3881 1826
rect 3933 1823 4092 1826
rect 4144 1823 4304 1826
rect 925 1777 946 1823
rect 2920 1777 2933 1823
rect 3268 1777 3281 1823
rect 3327 1777 3384 1823
rect 3430 1777 3487 1823
rect 3533 1777 3590 1823
rect 3636 1777 3693 1823
rect 3739 1777 3796 1823
rect 3842 1777 3881 1823
rect 3945 1777 4002 1823
rect 4048 1777 4092 1823
rect 4151 1777 4209 1823
rect 4255 1777 4304 1823
rect 925 1774 1083 1777
rect 1135 1774 1294 1777
rect 1346 1774 1506 1777
rect 1558 1774 1717 1777
rect 1769 1774 1927 1777
rect 1979 1774 2138 1777
rect 2190 1774 2349 1777
rect 2401 1774 2439 1777
rect 345 1733 2439 1774
rect 3843 1774 3881 1777
rect 3933 1774 4092 1777
rect 4144 1774 4304 1777
rect 4356 1774 4515 1826
rect 4567 1774 4605 1826
rect 3843 1740 4605 1774
rect 3844 1733 4605 1740
rect 4779 1860 5961 1867
rect 4779 1826 6555 1860
rect 4779 1774 4817 1826
rect 4869 1774 5027 1826
rect 5079 1774 5238 1826
rect 5290 1774 5450 1826
rect 5502 1774 5661 1826
rect 5713 1774 5871 1826
rect 5923 1823 6555 1826
rect 5923 1777 6086 1823
rect 6320 1777 6555 1823
rect 5923 1774 6555 1777
rect 4779 1740 6555 1774
rect 7543 1826 8439 1867
rect 7543 1823 7927 1826
rect 7979 1823 8138 1826
rect 7543 1777 7554 1823
rect 8070 1777 8138 1823
rect 7543 1774 7927 1777
rect 7979 1774 8138 1777
rect 8190 1774 8349 1826
rect 8401 1774 8439 1826
rect 4779 1733 5961 1740
rect 7543 1733 8439 1774
rect 8611 1826 8920 2312
rect 8611 1774 8649 1826
rect 8701 1823 8829 1826
rect 8705 1777 8817 1823
rect 8701 1774 8829 1777
rect 8881 1774 8920 1826
rect 345 1699 637 1733
rect 345 1653 452 1699
rect 498 1653 637 1699
rect 345 1535 637 1653
rect 3081 1657 3149 1668
rect 2616 1602 2924 1643
rect 2616 1599 2654 1602
rect 2706 1599 2834 1602
rect 2886 1599 2924 1602
rect 933 1553 946 1599
rect 2920 1553 2933 1599
rect 345 1489 452 1535
rect 498 1489 637 1535
rect 2616 1550 2654 1553
rect 2706 1550 2834 1553
rect 2886 1550 2924 1553
rect 2616 1510 2924 1550
rect 345 1397 637 1489
rect 345 1375 1090 1397
rect 345 1372 946 1375
rect 345 1326 452 1372
rect 498 1329 946 1372
rect 2920 1329 2933 1375
rect 498 1326 1090 1329
rect 345 1278 1090 1326
rect 345 1209 637 1278
rect 345 1163 452 1209
rect 498 1163 637 1209
rect 3081 1235 3092 1657
rect 3138 1235 3149 1657
rect 3378 1610 3686 1651
rect 3378 1599 3416 1610
rect 3468 1599 3596 1610
rect 3648 1599 3686 1610
rect 3268 1553 3281 1599
rect 3327 1553 3384 1599
rect 3468 1558 3487 1599
rect 3430 1553 3487 1558
rect 3533 1553 3590 1599
rect 3648 1558 3693 1599
rect 3636 1553 3693 1558
rect 3739 1553 3796 1599
rect 3842 1553 3899 1599
rect 3945 1553 4002 1599
rect 4048 1553 4105 1599
rect 4151 1553 4209 1599
rect 4255 1553 4268 1599
rect 3378 1518 3686 1553
rect 4891 1524 5863 1564
rect 7450 1561 7758 1577
rect 4891 1512 4929 1524
rect 4981 1512 5140 1524
rect 5192 1512 5351 1524
rect 5403 1512 5562 1524
rect 5614 1512 5773 1524
rect 5825 1512 5863 1524
rect 6035 1512 6550 1561
rect 7036 1536 7758 1561
rect 7036 1512 7488 1536
rect 7540 1512 7668 1536
rect 7720 1512 7758 1536
rect 4857 1466 4870 1512
rect 5120 1472 5140 1512
rect 5120 1466 5177 1472
rect 5223 1466 5280 1512
rect 5326 1472 5351 1512
rect 5326 1466 5383 1472
rect 5429 1466 5486 1512
rect 5532 1472 5562 1512
rect 5532 1466 5589 1472
rect 5635 1466 5692 1512
rect 5738 1472 5773 1512
rect 5738 1466 5795 1472
rect 5841 1466 5898 1512
rect 5944 1466 5957 1512
rect 6035 1466 6451 1512
rect 6497 1466 6568 1512
rect 6614 1466 6685 1512
rect 6731 1466 6803 1512
rect 6849 1466 6921 1512
rect 6967 1466 7039 1512
rect 7085 1484 7488 1512
rect 7085 1466 7506 1484
rect 7552 1466 7623 1512
rect 7720 1484 7740 1512
rect 7669 1466 7740 1484
rect 7786 1466 7858 1512
rect 7904 1466 7976 1512
rect 8022 1466 8094 1512
rect 8140 1466 8153 1512
rect 4891 1432 5863 1466
rect 6035 1441 6550 1466
rect 7036 1444 7758 1466
rect 7036 1441 7528 1444
rect 3825 1375 4315 1404
rect 3268 1329 3281 1375
rect 3327 1329 3384 1375
rect 3430 1329 3487 1375
rect 3533 1329 3590 1375
rect 3636 1329 3693 1375
rect 3739 1329 3796 1375
rect 3842 1364 3899 1375
rect 3842 1329 3864 1364
rect 3945 1329 4002 1375
rect 4048 1364 4105 1375
rect 4096 1329 4105 1364
rect 4151 1329 4209 1375
rect 4255 1364 4315 1375
rect 3825 1312 3864 1329
rect 3916 1312 4044 1329
rect 4096 1312 4224 1329
rect 4276 1312 4315 1364
rect 6035 1338 6151 1441
rect 3825 1271 4315 1312
rect 4561 1288 5957 1332
rect 345 1046 637 1163
rect 2616 1154 2924 1195
rect 2616 1151 2654 1154
rect 2706 1151 2834 1154
rect 2886 1151 2924 1154
rect 3081 1153 3149 1235
rect 4561 1242 4870 1288
rect 5120 1242 5177 1288
rect 5223 1242 5280 1288
rect 5326 1242 5383 1288
rect 5429 1242 5486 1288
rect 5532 1242 5589 1288
rect 5635 1242 5692 1288
rect 5738 1242 5795 1288
rect 5841 1242 5898 1288
rect 5944 1242 5957 1288
rect 4561 1210 5957 1242
rect 4561 1153 4679 1210
rect 933 1105 946 1151
rect 2920 1105 2933 1151
rect 3081 1116 4679 1153
rect 2616 1102 2654 1105
rect 2706 1102 2834 1105
rect 2886 1102 2924 1105
rect 2616 1062 2924 1102
rect 3081 1070 3413 1116
rect 3459 1070 3599 1116
rect 3645 1070 3786 1116
rect 3832 1070 3973 1116
rect 4019 1070 4159 1116
rect 4205 1070 4679 1116
rect 6035 1198 6072 1338
rect 6118 1198 6151 1338
rect 3081 1062 4679 1070
rect 4891 1064 5863 1104
rect 6035 1098 6151 1198
rect 6237 1338 6370 1361
rect 6237 1289 6294 1338
rect 6237 1237 6275 1289
rect 6237 1198 6294 1237
rect 6340 1198 6370 1338
rect 8255 1340 8323 1351
rect 6521 1330 7282 1336
rect 6520 1329 7282 1330
rect 6520 1296 7528 1329
rect 6520 1288 6558 1296
rect 6610 1288 6769 1296
rect 6821 1288 6981 1296
rect 6438 1242 6451 1288
rect 6497 1244 6558 1288
rect 6497 1242 6568 1244
rect 6614 1242 6685 1288
rect 6731 1244 6769 1288
rect 6731 1242 6803 1244
rect 6849 1242 6921 1288
rect 6967 1244 6981 1288
rect 7033 1288 7192 1296
rect 7033 1244 7039 1288
rect 6967 1242 7039 1244
rect 7085 1244 7192 1288
rect 7244 1288 7528 1296
rect 7244 1244 7506 1288
rect 7085 1242 7506 1244
rect 7552 1242 7623 1288
rect 7669 1242 7740 1288
rect 7786 1242 7858 1288
rect 7904 1242 7976 1288
rect 8022 1242 8094 1288
rect 8140 1242 8153 1288
rect 6520 1210 7528 1242
rect 6521 1203 7282 1210
rect 6237 1178 6370 1198
rect 8255 1200 8266 1340
rect 8312 1200 8323 1340
rect 8611 1288 8920 1774
rect 9089 1860 9205 2312
rect 9520 2279 9682 2410
rect 9520 2227 9591 2279
rect 9643 2227 9682 2279
rect 9520 2187 9682 2227
rect 9334 2091 9462 2104
rect 9334 2064 9463 2091
rect 9334 2047 9372 2064
rect 9424 2047 9463 2064
rect 9324 2001 9337 2047
rect 9424 2012 9459 2047
rect 9383 2001 9459 2012
rect 9505 2001 9582 2047
rect 9628 2001 9705 2047
rect 9751 2001 9764 2047
rect 9843 2036 9959 2434
rect 11826 2295 14106 2336
rect 11826 2243 13042 2295
rect 13094 2243 14106 2295
rect 11826 2203 14106 2243
rect 13938 2159 14106 2203
rect 13938 2113 13955 2159
rect 14095 2113 14106 2159
rect 9334 1972 9463 2001
rect 9843 1990 9878 2036
rect 9924 1990 9959 2036
rect 9843 1953 9959 1990
rect 10315 2064 13121 2105
rect 13938 2102 14106 2113
rect 10315 2012 11532 2064
rect 11584 2012 13121 2064
rect 10315 1971 13121 2012
rect 14202 2047 14318 2434
rect 14997 2404 17976 2445
rect 14997 2390 17083 2404
rect 14997 2344 15061 2390
rect 15201 2352 17083 2390
rect 17135 2352 17976 2404
rect 15201 2344 17976 2352
rect 14498 2288 14838 2329
rect 14997 2311 17976 2344
rect 18154 2398 18193 2450
rect 18245 2398 18284 2450
rect 18154 2375 18284 2398
rect 19641 2484 20113 2530
rect 20159 2484 20300 2530
rect 20346 2484 20487 2530
rect 20533 2484 20673 2530
rect 20719 2484 20860 2530
rect 20906 2484 21254 2530
rect 21394 2520 21702 2560
rect 21394 2495 21432 2520
rect 21484 2495 21612 2520
rect 21664 2495 21702 2520
rect 23682 2554 23820 2600
rect 23866 2554 23974 2600
rect 19641 2447 21254 2484
rect 21386 2449 21399 2495
rect 23373 2449 23386 2495
rect 19641 2390 19757 2447
rect 14498 2271 14536 2288
rect 14588 2271 14748 2288
rect 14800 2271 14838 2288
rect 14396 2225 14409 2271
rect 14455 2225 14522 2271
rect 14588 2236 14635 2271
rect 14568 2225 14635 2236
rect 14681 2225 14748 2271
rect 14800 2236 14861 2271
rect 14794 2225 14861 2236
rect 14907 2225 14920 2271
rect 18154 2235 18219 2375
rect 18265 2235 18284 2375
rect 19417 2358 19757 2390
rect 18362 2312 18375 2358
rect 18421 2312 18478 2358
rect 18524 2312 18581 2358
rect 18627 2312 18684 2358
rect 18730 2312 18787 2358
rect 18833 2312 18890 2358
rect 18936 2312 18993 2358
rect 19039 2312 19096 2358
rect 19142 2312 19199 2358
rect 19449 2312 19757 2358
rect 21186 2395 21254 2447
rect 21394 2427 21702 2449
rect 19417 2271 19757 2312
rect 19859 2288 20409 2329
rect 18154 2232 18284 2235
rect 14498 2196 14838 2225
rect 18154 2180 18193 2232
rect 18245 2180 18284 2232
rect 19859 2236 19897 2288
rect 19949 2271 20108 2288
rect 20160 2271 20319 2288
rect 19949 2236 20064 2271
rect 20160 2236 20168 2271
rect 19859 2225 20064 2236
rect 20110 2225 20168 2236
rect 20214 2225 20271 2271
rect 20317 2236 20319 2271
rect 20371 2271 20409 2288
rect 20371 2236 20374 2271
rect 20317 2225 20374 2236
rect 20420 2225 20477 2271
rect 20523 2225 20580 2271
rect 20626 2225 20683 2271
rect 20729 2225 20786 2271
rect 20832 2225 20889 2271
rect 20935 2225 20992 2271
rect 21038 2225 21051 2271
rect 19859 2196 20409 2225
rect 18154 2139 18284 2180
rect 18502 2134 19474 2165
rect 18362 2088 18375 2134
rect 18421 2088 18478 2134
rect 18524 2125 18581 2134
rect 18524 2088 18540 2125
rect 18627 2088 18684 2134
rect 18730 2125 18787 2134
rect 18730 2088 18751 2125
rect 18833 2088 18890 2134
rect 18936 2125 18993 2134
rect 18936 2088 18962 2125
rect 19039 2088 19096 2134
rect 19142 2125 19199 2134
rect 19142 2088 19173 2125
rect 19449 2088 19474 2134
rect 18502 2073 18540 2088
rect 18592 2073 18751 2088
rect 18803 2073 18962 2088
rect 19014 2073 19173 2088
rect 19225 2073 19384 2088
rect 19436 2073 19474 2088
rect 14202 2001 14409 2047
rect 14455 2001 14522 2047
rect 14568 2001 14635 2047
rect 14681 2001 14748 2047
rect 14794 2001 14861 2047
rect 14907 2001 14920 2047
rect 18502 2033 19474 2073
rect 20632 2050 20940 2090
rect 20632 2047 20670 2050
rect 20722 2047 20850 2050
rect 20902 2047 20940 2050
rect 12959 1964 13121 1971
rect 12959 1918 12970 1964
rect 13110 1918 13121 1964
rect 12959 1907 13121 1918
rect 15181 1987 18143 2023
rect 20051 2001 20064 2047
rect 20110 2001 20168 2047
rect 20214 2001 20271 2047
rect 20317 2001 20374 2047
rect 20420 2001 20477 2047
rect 20523 2001 20580 2047
rect 20626 2001 20670 2047
rect 20729 2001 20786 2047
rect 20832 2001 20850 2047
rect 20935 2001 20992 2047
rect 21038 2001 21051 2047
rect 15181 1941 15216 1987
rect 15262 1941 15374 1987
rect 15420 1941 15532 1987
rect 15578 1941 15690 1987
rect 15736 1941 15848 1987
rect 15894 1941 16006 1987
rect 16052 1941 16165 1987
rect 16211 1941 16323 1987
rect 16369 1941 16481 1987
rect 16527 1941 16639 1987
rect 16685 1941 16797 1987
rect 16843 1941 16955 1987
rect 17001 1941 17113 1987
rect 17159 1941 17272 1987
rect 17318 1941 17430 1987
rect 17476 1941 17588 1987
rect 17634 1941 17746 1987
rect 17792 1941 17904 1987
rect 17950 1941 18062 1987
rect 18108 1941 18143 1987
rect 20632 1998 20670 2001
rect 20722 1998 20850 2001
rect 20902 1998 20940 2001
rect 20632 1957 20940 1998
rect 21186 1973 21197 2395
rect 21243 1973 21254 2395
rect 23682 2322 23974 2554
rect 23182 2271 23974 2322
rect 21386 2225 21399 2271
rect 23373 2225 23974 2271
rect 23182 2203 23974 2225
rect 23682 2111 23974 2203
rect 21394 2057 21702 2097
rect 21394 2047 21432 2057
rect 21484 2047 21612 2057
rect 21664 2047 21702 2057
rect 23682 2065 23820 2111
rect 23866 2065 23974 2111
rect 21386 2001 21399 2047
rect 23373 2001 23386 2047
rect 21186 1962 21254 1973
rect 21394 1964 21702 2001
rect 9812 1860 10120 1867
rect 10385 1860 12583 1874
rect 13350 1860 14111 1867
rect 9089 1837 12583 1860
rect 13301 1837 14111 1860
rect 9089 1826 14111 1837
rect 9089 1823 9850 1826
rect 9089 1777 9337 1823
rect 9383 1777 9459 1823
rect 9505 1777 9582 1823
rect 9628 1777 9705 1823
rect 9751 1777 9850 1823
rect 9089 1774 9850 1777
rect 9902 1774 10030 1826
rect 10082 1823 13387 1826
rect 10082 1777 10433 1823
rect 10479 1777 10591 1823
rect 10637 1777 10749 1823
rect 10795 1777 10907 1823
rect 10953 1777 11066 1823
rect 11112 1777 11224 1823
rect 11270 1777 11382 1823
rect 11428 1777 11540 1823
rect 11586 1777 11698 1823
rect 11744 1777 11856 1823
rect 11902 1777 12015 1823
rect 12061 1777 12173 1823
rect 12219 1777 12331 1823
rect 12377 1777 12489 1823
rect 12535 1777 13336 1823
rect 13382 1777 13387 1823
rect 10082 1774 13387 1777
rect 13439 1823 13598 1826
rect 13439 1777 13503 1823
rect 13549 1777 13598 1823
rect 13439 1774 13598 1777
rect 13650 1823 13810 1826
rect 13862 1823 14021 1826
rect 13650 1777 13668 1823
rect 13714 1777 13810 1823
rect 13879 1777 14021 1823
rect 13650 1774 13810 1777
rect 13862 1774 14021 1777
rect 14073 1774 14111 1826
rect 9089 1763 14111 1774
rect 9089 1740 12583 1763
rect 13301 1740 14111 1763
rect 9089 1288 9205 1740
rect 9812 1733 10120 1740
rect 10385 1726 12583 1740
rect 13350 1733 14111 1740
rect 14393 1860 14943 1867
rect 15181 1860 18143 1941
rect 23682 1947 23974 2065
rect 23682 1901 23820 1947
rect 23866 1901 23974 1947
rect 23682 1867 23974 1901
rect 18397 1860 19579 1867
rect 19905 1860 20456 1867
rect 14393 1826 19579 1860
rect 14393 1823 14431 1826
rect 14483 1823 14642 1826
rect 14694 1823 14853 1826
rect 14905 1823 18435 1826
rect 14393 1777 14409 1823
rect 14483 1777 14522 1823
rect 14568 1777 14635 1823
rect 14694 1777 14748 1823
rect 14794 1777 14853 1823
rect 14907 1777 15216 1823
rect 15262 1777 15374 1823
rect 15420 1777 15532 1823
rect 15578 1777 15690 1823
rect 15736 1777 15848 1823
rect 15894 1777 16006 1823
rect 16052 1777 16165 1823
rect 16211 1777 16323 1823
rect 16369 1777 16481 1823
rect 16527 1777 16639 1823
rect 16685 1777 16797 1823
rect 16843 1777 16955 1823
rect 17001 1777 17113 1823
rect 17159 1777 17272 1823
rect 17318 1777 17430 1823
rect 17476 1777 17588 1823
rect 17634 1777 17746 1823
rect 17792 1777 17904 1823
rect 17950 1777 18062 1823
rect 18108 1777 18435 1823
rect 14393 1774 14431 1777
rect 14483 1774 14642 1777
rect 14694 1774 14853 1777
rect 14905 1774 18435 1777
rect 18487 1774 18645 1826
rect 18697 1774 18856 1826
rect 18908 1774 19068 1826
rect 19120 1774 19279 1826
rect 19331 1774 19489 1826
rect 19541 1774 19579 1826
rect 14393 1740 19579 1774
rect 19904 1826 20456 1860
rect 19904 1774 19943 1826
rect 19995 1823 20154 1826
rect 20206 1823 20365 1826
rect 20417 1823 20456 1826
rect 21875 1826 23974 1867
rect 21875 1823 21913 1826
rect 21965 1823 22124 1826
rect 22176 1823 22335 1826
rect 22387 1823 22545 1826
rect 22597 1823 22756 1826
rect 22808 1823 22968 1826
rect 23020 1823 23179 1826
rect 23231 1823 23389 1826
rect 19995 1777 20064 1823
rect 20110 1777 20154 1823
rect 20214 1777 20271 1823
rect 20317 1777 20365 1823
rect 20420 1777 20477 1823
rect 20523 1777 20580 1823
rect 20626 1777 20683 1823
rect 20729 1777 20786 1823
rect 20832 1777 20889 1823
rect 20935 1777 20992 1823
rect 21038 1777 21051 1823
rect 21386 1777 21399 1823
rect 23373 1777 23389 1823
rect 19995 1774 20154 1777
rect 20206 1774 20365 1777
rect 20417 1774 20456 1777
rect 19904 1740 20456 1774
rect 14393 1733 14943 1740
rect 12959 1682 13121 1693
rect 9334 1599 9463 1628
rect 9843 1610 9959 1647
rect 12959 1636 12970 1682
rect 13110 1636 13121 1682
rect 12959 1629 13121 1636
rect 9324 1553 9337 1599
rect 9383 1588 9459 1599
rect 9424 1553 9459 1588
rect 9505 1553 9582 1599
rect 9628 1553 9705 1599
rect 9751 1553 9764 1599
rect 9843 1564 9878 1610
rect 9924 1564 9959 1610
rect 9334 1536 9372 1553
rect 9424 1536 9463 1553
rect 9334 1509 9463 1536
rect 9334 1496 9462 1509
rect 9520 1373 9682 1413
rect 9520 1321 9591 1373
rect 9643 1321 9682 1373
rect 8605 1242 8618 1288
rect 8664 1242 8741 1288
rect 8787 1242 8864 1288
rect 8910 1242 8923 1288
rect 9089 1242 9238 1288
rect 9284 1242 9327 1288
rect 8611 1210 8920 1242
rect 9089 1210 9205 1242
rect 7450 1098 7758 1103
rect 6035 1064 6550 1098
rect 7036 1064 7758 1098
rect 8255 1078 8323 1200
rect 9520 1190 9682 1321
rect 9406 1187 9682 1190
rect 9406 1179 9591 1187
rect 9406 1133 9441 1179
rect 9487 1135 9591 1179
rect 9643 1166 9682 1187
rect 9843 1166 9959 1564
rect 10315 1588 13121 1629
rect 15181 1659 18143 1740
rect 18397 1733 19579 1740
rect 19905 1733 20456 1740
rect 21875 1774 21913 1777
rect 21965 1774 22124 1777
rect 22176 1774 22335 1777
rect 22387 1774 22545 1777
rect 22597 1774 22756 1777
rect 22808 1774 22968 1777
rect 23020 1774 23179 1777
rect 23231 1774 23389 1777
rect 23441 1774 23600 1826
rect 23652 1774 23811 1826
rect 23863 1774 23974 1826
rect 21875 1733 23974 1774
rect 15181 1613 15216 1659
rect 15262 1613 15374 1659
rect 15420 1613 15532 1659
rect 15578 1613 15690 1659
rect 15736 1613 15848 1659
rect 15894 1613 16006 1659
rect 16052 1613 16165 1659
rect 16211 1613 16323 1659
rect 16369 1613 16481 1659
rect 16527 1613 16639 1659
rect 16685 1613 16797 1659
rect 16843 1613 16955 1659
rect 17001 1613 17113 1659
rect 17159 1613 17272 1659
rect 17318 1613 17430 1659
rect 17476 1613 17588 1659
rect 17634 1613 17746 1659
rect 17792 1613 17904 1659
rect 17950 1613 18062 1659
rect 18108 1613 18143 1659
rect 23682 1699 23974 1733
rect 23682 1653 23820 1699
rect 23866 1653 23974 1699
rect 10315 1536 11532 1588
rect 11584 1536 13121 1588
rect 10315 1495 13121 1536
rect 14202 1553 14409 1599
rect 14455 1553 14522 1599
rect 14568 1553 14635 1599
rect 14681 1553 14748 1599
rect 14794 1553 14861 1599
rect 14907 1553 14920 1599
rect 15181 1577 18143 1613
rect 20632 1602 20940 1643
rect 20632 1599 20670 1602
rect 20722 1599 20850 1602
rect 20902 1599 20940 1602
rect 21186 1627 21254 1638
rect 13938 1487 14106 1498
rect 13938 1441 13955 1487
rect 14095 1441 14106 1487
rect 13938 1397 14106 1441
rect 11826 1357 14106 1397
rect 11826 1305 13042 1357
rect 13094 1305 14106 1357
rect 11826 1264 14106 1305
rect 14202 1166 14318 1553
rect 18502 1527 19474 1567
rect 20051 1553 20064 1599
rect 20110 1553 20168 1599
rect 20214 1553 20271 1599
rect 20317 1553 20374 1599
rect 20420 1553 20477 1599
rect 20523 1553 20580 1599
rect 20626 1553 20670 1599
rect 20729 1553 20786 1599
rect 20832 1553 20850 1599
rect 20935 1553 20992 1599
rect 21038 1553 21051 1599
rect 18502 1512 18540 1527
rect 18592 1512 18751 1527
rect 18803 1512 18962 1527
rect 19014 1512 19173 1527
rect 19225 1512 19384 1527
rect 19436 1512 19474 1527
rect 18362 1466 18375 1512
rect 18421 1466 18478 1512
rect 18524 1475 18540 1512
rect 18524 1466 18581 1475
rect 18627 1466 18684 1512
rect 18730 1475 18751 1512
rect 18730 1466 18787 1475
rect 18833 1466 18890 1512
rect 18936 1475 18962 1512
rect 18936 1466 18993 1475
rect 19039 1466 19096 1512
rect 19142 1475 19173 1512
rect 19142 1466 19199 1475
rect 19449 1466 19474 1512
rect 20632 1550 20670 1553
rect 20722 1550 20850 1553
rect 20902 1550 20940 1553
rect 20632 1510 20940 1550
rect 18154 1420 18284 1461
rect 18502 1435 19474 1466
rect 14498 1375 14838 1404
rect 14396 1329 14409 1375
rect 14455 1329 14522 1375
rect 14568 1364 14635 1375
rect 14588 1329 14635 1364
rect 14681 1329 14748 1375
rect 14794 1364 14861 1375
rect 14800 1329 14861 1364
rect 14907 1329 14920 1375
rect 18154 1368 18193 1420
rect 18245 1368 18284 1420
rect 18154 1365 18284 1368
rect 14498 1312 14536 1329
rect 14588 1312 14748 1329
rect 14800 1312 14838 1329
rect 14498 1271 14838 1312
rect 14997 1256 17976 1289
rect 14997 1210 15061 1256
rect 15201 1248 17976 1256
rect 15201 1210 17461 1248
rect 14997 1196 17461 1210
rect 17513 1196 17976 1248
rect 9643 1151 14515 1166
rect 14997 1155 17976 1196
rect 18154 1225 18219 1365
rect 18265 1225 18284 1365
rect 19859 1375 20409 1404
rect 19859 1364 20064 1375
rect 20110 1364 20168 1375
rect 19417 1288 19757 1329
rect 18362 1242 18375 1288
rect 18421 1242 18478 1288
rect 18524 1242 18581 1288
rect 18627 1242 18684 1288
rect 18730 1242 18787 1288
rect 18833 1242 18890 1288
rect 18936 1242 18993 1288
rect 19039 1242 19096 1288
rect 19142 1242 19199 1288
rect 19449 1242 19757 1288
rect 19859 1312 19897 1364
rect 19949 1329 20064 1364
rect 20160 1329 20168 1364
rect 20214 1329 20271 1375
rect 20317 1364 20374 1375
rect 20317 1329 20319 1364
rect 19949 1312 20108 1329
rect 20160 1312 20319 1329
rect 20371 1329 20374 1364
rect 20420 1329 20477 1375
rect 20523 1329 20580 1375
rect 20626 1329 20683 1375
rect 20729 1329 20786 1375
rect 20832 1329 20889 1375
rect 20935 1329 20992 1375
rect 21038 1329 21051 1375
rect 20371 1312 20409 1329
rect 19859 1271 20409 1312
rect 18154 1202 18284 1225
rect 19417 1210 19757 1242
rect 9643 1135 14409 1151
rect 9487 1133 14409 1135
rect 9406 1130 14409 1133
rect 9406 1084 13336 1130
rect 13382 1084 13503 1130
rect 13549 1084 13668 1130
rect 13714 1084 13833 1130
rect 13879 1105 14409 1130
rect 14455 1105 14522 1151
rect 14568 1105 14635 1151
rect 14681 1105 14748 1151
rect 14794 1105 14861 1151
rect 14907 1105 14920 1151
rect 18154 1150 18193 1202
rect 18245 1150 18284 1202
rect 18154 1110 18284 1150
rect 19641 1153 19757 1210
rect 21186 1205 21197 1627
rect 21243 1205 21254 1627
rect 21394 1599 21702 1636
rect 21386 1553 21399 1599
rect 23373 1553 23386 1599
rect 21394 1543 21432 1553
rect 21484 1543 21612 1553
rect 21664 1543 21702 1553
rect 21394 1503 21702 1543
rect 23682 1535 23974 1653
rect 23682 1489 23820 1535
rect 23866 1489 23974 1535
rect 23682 1397 23974 1489
rect 23182 1375 23974 1397
rect 21386 1329 21399 1375
rect 23373 1329 23974 1375
rect 23182 1278 23974 1329
rect 21186 1153 21254 1205
rect 19641 1116 21254 1153
rect 21394 1151 21702 1173
rect 13879 1084 14515 1105
rect 8255 1064 9320 1078
rect 345 1000 452 1046
rect 498 1000 637 1046
rect 3081 1033 4240 1062
rect 4857 1018 4870 1064
rect 5120 1018 5140 1064
rect 5223 1018 5280 1064
rect 5326 1018 5351 1064
rect 5429 1018 5486 1064
rect 5532 1018 5562 1064
rect 5635 1018 5692 1064
rect 5738 1018 5773 1064
rect 5841 1018 5898 1064
rect 5944 1018 5957 1064
rect 6035 1018 6451 1064
rect 6497 1018 6568 1064
rect 6614 1018 6685 1064
rect 6731 1018 6803 1064
rect 6849 1018 6921 1064
rect 6967 1018 7039 1064
rect 7085 1062 7506 1064
rect 7085 1018 7488 1062
rect 7552 1018 7623 1064
rect 7669 1062 7740 1064
rect 7720 1018 7740 1062
rect 7786 1018 7858 1064
rect 7904 1018 7976 1064
rect 8022 1018 8094 1064
rect 8140 1018 8153 1064
rect 8255 1018 8618 1064
rect 8664 1018 8741 1064
rect 8787 1018 8864 1064
rect 8910 1018 9238 1064
rect 9284 1018 9327 1064
rect 9406 1046 14515 1084
rect 18502 1064 19474 1104
rect 18362 1018 18375 1064
rect 18421 1018 18478 1064
rect 18524 1018 18540 1064
rect 18627 1018 18684 1064
rect 18730 1018 18751 1064
rect 18833 1018 18890 1064
rect 18936 1018 18962 1064
rect 19039 1018 19096 1064
rect 19142 1018 19173 1064
rect 19449 1018 19474 1064
rect 19641 1070 20113 1116
rect 20159 1070 20300 1116
rect 20346 1070 20487 1116
rect 20533 1070 20673 1116
rect 20719 1070 20860 1116
rect 20906 1070 21254 1116
rect 21386 1105 21399 1151
rect 23373 1105 23386 1151
rect 19641 1060 21254 1070
rect 20078 1033 21254 1060
rect 21394 1080 21432 1105
rect 21484 1080 21612 1105
rect 21664 1080 21702 1105
rect 21394 1040 21702 1080
rect 23682 1046 23974 1278
rect 345 967 637 1000
rect 4891 1012 4929 1018
rect 4981 1012 5140 1018
rect 5192 1012 5351 1018
rect 5403 1012 5562 1018
rect 5614 1012 5773 1018
rect 5825 1012 5863 1018
rect 4467 967 4622 974
rect 4891 972 5863 1012
rect 6035 978 6550 1018
rect 7036 1010 7488 1018
rect 7540 1010 7668 1018
rect 7720 1010 7758 1018
rect 7036 978 7758 1010
rect 7450 970 7758 978
rect 345 926 2439 967
rect 345 874 451 926
rect 503 874 662 926
rect 714 874 873 926
rect 925 874 1083 926
rect 1135 874 1294 926
rect 1346 874 1506 926
rect 1558 874 1717 926
rect 1769 874 1927 926
rect 1979 874 2138 926
rect 2190 874 2349 926
rect 2401 874 2439 926
rect 345 833 2439 874
rect 4314 926 4622 967
rect 8255 958 9320 1018
rect 18502 1012 18540 1018
rect 18592 1012 18751 1018
rect 18803 1012 18962 1018
rect 19014 1012 19173 1018
rect 19225 1012 19384 1018
rect 19436 1012 19474 1018
rect 18502 972 19474 1012
rect 23682 1000 23820 1046
rect 23866 1000 23974 1046
rect 19696 967 19852 974
rect 23682 967 23974 1000
rect 4314 874 4352 926
rect 4404 923 4532 926
rect 4404 877 4513 923
rect 4404 874 4532 877
rect 4584 874 4622 926
rect 4314 833 4622 874
rect 19696 926 20005 967
rect 19696 874 19735 926
rect 19787 923 19915 926
rect 19803 877 19915 923
rect 19787 874 19915 877
rect 19967 874 20005 926
rect 345 800 637 833
rect 4467 826 4622 833
rect 345 754 452 800
rect 498 754 637 800
rect 4891 788 5863 828
rect 7450 822 7758 830
rect 4891 782 4929 788
rect 4981 782 5140 788
rect 5192 782 5351 788
rect 5403 782 5562 788
rect 5614 782 5773 788
rect 5825 782 5863 788
rect 6035 782 6550 822
rect 7036 790 7758 822
rect 7036 782 7488 790
rect 7540 782 7668 790
rect 7720 782 7758 790
rect 8255 782 9320 842
rect 19696 833 20005 874
rect 21875 926 23974 967
rect 21875 874 21913 926
rect 21965 874 22124 926
rect 22176 874 22335 926
rect 22387 874 22545 926
rect 22597 874 22756 926
rect 22808 874 22968 926
rect 23020 874 23179 926
rect 23231 874 23389 926
rect 23441 874 23600 926
rect 23652 874 23811 926
rect 23863 874 23974 926
rect 21875 833 23974 874
rect 18502 788 19474 828
rect 19696 826 19852 833
rect 18502 782 18540 788
rect 18592 782 18751 788
rect 18803 782 18962 788
rect 19014 782 19173 788
rect 19225 782 19384 788
rect 19436 782 19474 788
rect 345 637 637 754
rect 3081 738 4240 767
rect 2616 698 2924 738
rect 2616 695 2654 698
rect 2706 695 2834 698
rect 2886 695 2924 698
rect 3081 730 4679 738
rect 4857 736 4870 782
rect 5120 736 5140 782
rect 5223 736 5280 782
rect 5326 736 5351 782
rect 5429 736 5486 782
rect 5532 736 5562 782
rect 5635 736 5692 782
rect 5738 736 5773 782
rect 5841 736 5898 782
rect 5944 736 5957 782
rect 6035 736 6451 782
rect 6497 736 6568 782
rect 6614 736 6685 782
rect 6731 736 6803 782
rect 6849 736 6921 782
rect 6967 736 7039 782
rect 7085 738 7488 782
rect 7085 736 7506 738
rect 7552 736 7623 782
rect 7720 738 7740 782
rect 7669 736 7740 738
rect 7786 736 7858 782
rect 7904 736 7976 782
rect 8022 736 8094 782
rect 8140 736 8153 782
rect 8255 736 8618 782
rect 8664 736 8741 782
rect 8787 736 8864 782
rect 8910 736 9238 782
rect 9284 736 9327 782
rect 933 649 946 695
rect 2920 649 2933 695
rect 3081 684 3413 730
rect 3459 684 3599 730
rect 3645 684 3786 730
rect 3832 684 3973 730
rect 4019 684 4159 730
rect 4205 684 4679 730
rect 4891 696 5863 736
rect 6035 702 6550 736
rect 7036 702 7758 736
rect 345 591 452 637
rect 498 591 637 637
rect 2616 646 2654 649
rect 2706 646 2834 649
rect 2886 646 2924 649
rect 2616 605 2924 646
rect 3081 647 4679 684
rect 345 522 637 591
rect 3081 565 3149 647
rect 345 474 1090 522
rect 345 428 452 474
rect 498 471 1090 474
rect 498 428 946 471
rect 345 425 946 428
rect 2920 425 2933 471
rect 345 403 1090 425
rect 345 311 637 403
rect 345 265 452 311
rect 498 265 637 311
rect 345 147 637 265
rect 2616 250 2924 290
rect 2616 247 2654 250
rect 2706 247 2834 250
rect 2886 247 2924 250
rect 933 201 946 247
rect 2920 201 2933 247
rect 2616 198 2654 201
rect 2706 198 2834 201
rect 2886 198 2924 201
rect 2616 157 2924 198
rect 345 101 452 147
rect 498 101 637 147
rect 3081 143 3092 565
rect 3138 143 3149 565
rect 4561 590 4679 647
rect 6035 602 6151 702
rect 7450 697 7758 702
rect 8255 722 9320 736
rect 4561 558 5957 590
rect 3825 488 4315 529
rect 3825 471 3864 488
rect 3916 471 4044 488
rect 4096 471 4224 488
rect 3268 425 3281 471
rect 3327 425 3384 471
rect 3430 425 3487 471
rect 3533 425 3590 471
rect 3636 425 3693 471
rect 3739 425 3796 471
rect 3842 436 3864 471
rect 3842 425 3899 436
rect 3945 425 4002 471
rect 4096 436 4105 471
rect 4048 425 4105 436
rect 4151 425 4209 471
rect 4276 436 4315 488
rect 4561 512 4870 558
rect 5120 512 5177 558
rect 5223 512 5280 558
rect 5326 512 5383 558
rect 5429 512 5486 558
rect 5532 512 5589 558
rect 5635 512 5692 558
rect 5738 512 5795 558
rect 5841 512 5898 558
rect 5944 512 5957 558
rect 4561 468 5957 512
rect 4255 425 4315 436
rect 3825 396 4315 425
rect 6035 462 6072 602
rect 6118 462 6151 602
rect 4891 334 5863 368
rect 6035 359 6151 462
rect 6237 602 6370 622
rect 6237 563 6294 602
rect 6237 511 6275 563
rect 6237 462 6294 511
rect 6340 462 6370 602
rect 8255 600 8323 722
rect 9406 716 14515 754
rect 18362 736 18375 782
rect 18421 736 18478 782
rect 18524 736 18540 782
rect 18627 736 18684 782
rect 18730 736 18751 782
rect 18833 736 18890 782
rect 18936 736 18962 782
rect 19039 736 19096 782
rect 19142 736 19173 782
rect 19449 736 19474 782
rect 23682 800 23974 833
rect 20078 740 21254 767
rect 9406 670 13336 716
rect 13382 670 13503 716
rect 13549 670 13668 716
rect 13714 670 13833 716
rect 13879 695 14515 716
rect 18502 696 19474 736
rect 19641 730 21254 740
rect 13879 670 14409 695
rect 9406 667 14409 670
rect 9406 621 9441 667
rect 9487 665 14409 667
rect 9487 621 9591 665
rect 9406 613 9591 621
rect 9643 649 14409 665
rect 14455 649 14522 695
rect 14568 649 14635 695
rect 14681 649 14748 695
rect 14794 649 14861 695
rect 14907 649 14920 695
rect 18154 650 18284 690
rect 9643 634 14515 649
rect 9643 613 9682 634
rect 9406 610 9682 613
rect 6521 590 7282 597
rect 6520 558 7528 590
rect 6438 512 6451 558
rect 6497 556 6568 558
rect 6497 512 6558 556
rect 6614 512 6685 558
rect 6731 556 6803 558
rect 6731 512 6769 556
rect 6849 512 6921 558
rect 6967 556 7039 558
rect 6967 512 6981 556
rect 6520 504 6558 512
rect 6610 504 6769 512
rect 6821 504 6981 512
rect 7033 512 7039 556
rect 7085 556 7506 558
rect 7085 512 7192 556
rect 7033 504 7192 512
rect 7244 512 7506 556
rect 7552 512 7623 558
rect 7669 512 7740 558
rect 7786 512 7858 558
rect 7904 512 7976 558
rect 8022 512 8094 558
rect 8140 512 8153 558
rect 7244 504 7528 512
rect 6520 471 7528 504
rect 6520 470 7282 471
rect 6521 464 7282 470
rect 6237 439 6370 462
rect 8255 460 8266 600
rect 8312 460 8323 600
rect 8611 558 8920 590
rect 9089 558 9205 590
rect 8605 512 8618 558
rect 8664 512 8741 558
rect 8787 512 8864 558
rect 8910 512 8923 558
rect 9089 512 9238 558
rect 9284 512 9327 558
rect 8255 449 8323 460
rect 6035 334 6550 359
rect 7036 356 7528 359
rect 7036 334 7758 356
rect 4857 288 4870 334
rect 5120 328 5177 334
rect 5120 288 5140 328
rect 5223 288 5280 334
rect 5326 328 5383 334
rect 5326 288 5351 328
rect 5429 288 5486 334
rect 5532 328 5589 334
rect 5532 288 5562 328
rect 5635 288 5692 334
rect 5738 328 5795 334
rect 5738 288 5773 328
rect 5841 288 5898 334
rect 5944 288 5957 334
rect 6035 288 6451 334
rect 6497 288 6568 334
rect 6614 288 6685 334
rect 6731 288 6803 334
rect 6849 288 6921 334
rect 6967 288 7039 334
rect 7085 316 7506 334
rect 7085 288 7488 316
rect 7552 288 7623 334
rect 7669 316 7740 334
rect 7720 288 7740 316
rect 7786 288 7858 334
rect 7904 288 7976 334
rect 8022 288 8094 334
rect 8140 288 8153 334
rect 3378 247 3686 282
rect 4891 276 4929 288
rect 4981 276 5140 288
rect 5192 276 5351 288
rect 5403 276 5562 288
rect 5614 276 5773 288
rect 5825 276 5863 288
rect 3268 201 3281 247
rect 3327 201 3384 247
rect 3430 242 3487 247
rect 3468 201 3487 242
rect 3533 201 3590 247
rect 3636 242 3693 247
rect 3648 201 3693 242
rect 3739 201 3796 247
rect 3842 201 3899 247
rect 3945 201 4002 247
rect 4048 201 4105 247
rect 4151 201 4209 247
rect 4255 201 4268 247
rect 4891 236 5863 276
rect 6035 239 6550 288
rect 7036 264 7488 288
rect 7540 264 7668 288
rect 7720 264 7758 288
rect 7036 239 7758 264
rect 7450 223 7758 239
rect 3378 190 3416 201
rect 3468 190 3596 201
rect 3648 190 3686 201
rect 3378 149 3686 190
rect 3081 132 3149 143
rect 345 67 637 101
rect 345 26 2439 67
rect 3844 60 4605 67
rect 345 -26 451 26
rect 503 -26 662 26
rect 714 -26 873 26
rect 925 23 1083 26
rect 1135 23 1294 26
rect 1346 23 1506 26
rect 1558 23 1717 26
rect 1769 23 1927 26
rect 1979 23 2138 26
rect 2190 23 2349 26
rect 2401 23 2439 26
rect 3843 26 4605 60
rect 3843 23 3881 26
rect 3933 23 4092 26
rect 4144 23 4304 26
rect 925 -23 946 23
rect 2920 -23 2933 23
rect 3268 -23 3281 23
rect 3327 -23 3384 23
rect 3430 -23 3487 23
rect 3533 -23 3590 23
rect 3636 -23 3693 23
rect 3739 -23 3796 23
rect 3842 -23 3881 23
rect 3945 -23 4002 23
rect 4048 -23 4092 23
rect 4151 -23 4209 23
rect 4255 -23 4304 23
rect 925 -26 1083 -23
rect 1135 -26 1294 -23
rect 1346 -26 1506 -23
rect 1558 -26 1717 -23
rect 1769 -26 1927 -23
rect 1979 -26 2138 -23
rect 2190 -26 2349 -23
rect 2401 -26 2439 -23
rect 345 -67 2439 -26
rect 3843 -26 3881 -23
rect 3933 -26 4092 -23
rect 4144 -26 4304 -23
rect 4356 -26 4515 26
rect 4567 -26 4605 26
rect 3843 -60 4605 -26
rect 3844 -66 4605 -60
rect 4779 60 5961 67
rect 4779 26 6555 60
rect 4779 -26 4817 26
rect 4869 -26 5027 26
rect 5079 -26 5238 26
rect 5290 -26 5450 26
rect 5502 -26 5661 26
rect 5713 -26 5871 26
rect 5923 23 6555 26
rect 5923 -23 6086 23
rect 6320 -23 6555 23
rect 5923 -26 6555 -23
rect 4779 -60 6555 -26
rect 7543 26 8439 67
rect 7543 23 7927 26
rect 7979 23 8138 26
rect 7543 -23 7554 23
rect 8070 -23 8138 23
rect 7543 -26 7927 -23
rect 7979 -26 8138 -23
rect 8190 -26 8349 26
rect 8401 -26 8439 26
rect 4779 -67 5961 -60
rect 7543 -66 8439 -26
rect 8611 26 8920 512
rect 8611 -26 8649 26
rect 8701 23 8829 26
rect 8705 -23 8817 23
rect 8701 -26 8829 -23
rect 8881 -26 8920 26
rect 8611 -60 8920 -26
rect 9089 60 9205 512
rect 9520 479 9682 610
rect 9520 427 9591 479
rect 9643 427 9682 479
rect 9520 387 9682 427
rect 9334 291 9462 304
rect 9334 264 9463 291
rect 9334 247 9372 264
rect 9424 247 9463 264
rect 9324 201 9337 247
rect 9424 212 9459 247
rect 9383 201 9459 212
rect 9505 201 9582 247
rect 9628 201 9705 247
rect 9751 201 9764 247
rect 9843 236 9959 634
rect 11826 495 14106 536
rect 11826 443 13042 495
rect 13094 443 14106 495
rect 11826 403 14106 443
rect 13938 359 14106 403
rect 13938 313 13955 359
rect 14095 313 14106 359
rect 9334 172 9463 201
rect 9843 190 9878 236
rect 9924 190 9959 236
rect 9843 153 9959 190
rect 10315 264 13121 305
rect 13938 302 14106 313
rect 10315 212 11532 264
rect 11584 212 13121 264
rect 10315 171 13121 212
rect 14202 247 14318 634
rect 14997 604 17976 645
rect 14997 590 17838 604
rect 14997 544 15061 590
rect 15201 552 17838 590
rect 17890 552 17976 604
rect 15201 544 17976 552
rect 14498 488 14838 529
rect 14997 511 17976 544
rect 18154 598 18193 650
rect 18245 598 18284 650
rect 18154 575 18284 598
rect 19641 684 20113 730
rect 20159 684 20300 730
rect 20346 684 20487 730
rect 20533 684 20673 730
rect 20719 684 20860 730
rect 20906 684 21254 730
rect 21394 720 21702 760
rect 21394 695 21432 720
rect 21484 695 21612 720
rect 21664 695 21702 720
rect 23682 754 23820 800
rect 23866 754 23974 800
rect 19641 647 21254 684
rect 21386 649 21399 695
rect 23373 649 23386 695
rect 19641 590 19757 647
rect 14498 471 14536 488
rect 14588 471 14748 488
rect 14800 471 14838 488
rect 14396 425 14409 471
rect 14455 425 14522 471
rect 14588 436 14635 471
rect 14568 425 14635 436
rect 14681 425 14748 471
rect 14800 436 14861 471
rect 14794 425 14861 436
rect 14907 425 14920 471
rect 18154 435 18219 575
rect 18265 435 18284 575
rect 19417 558 19757 590
rect 18362 512 18375 558
rect 18421 512 18478 558
rect 18524 512 18581 558
rect 18627 512 18684 558
rect 18730 512 18787 558
rect 18833 512 18890 558
rect 18936 512 18993 558
rect 19039 512 19096 558
rect 19142 512 19199 558
rect 19449 512 19757 558
rect 21186 595 21254 647
rect 21394 627 21702 649
rect 19417 471 19757 512
rect 19859 488 20409 529
rect 18154 432 18284 435
rect 14498 396 14838 425
rect 18154 380 18193 432
rect 18245 380 18284 432
rect 19859 436 19897 488
rect 19949 471 20108 488
rect 20160 471 20319 488
rect 19949 436 20064 471
rect 20160 436 20168 471
rect 19859 425 20064 436
rect 20110 425 20168 436
rect 20214 425 20271 471
rect 20317 436 20319 471
rect 20371 471 20409 488
rect 20371 436 20374 471
rect 20317 425 20374 436
rect 20420 425 20477 471
rect 20523 425 20580 471
rect 20626 425 20683 471
rect 20729 425 20786 471
rect 20832 425 20889 471
rect 20935 425 20992 471
rect 21038 425 21051 471
rect 19859 396 20409 425
rect 18154 339 18284 380
rect 18502 334 19474 365
rect 18362 288 18375 334
rect 18421 288 18478 334
rect 18524 325 18581 334
rect 18524 288 18540 325
rect 18627 288 18684 334
rect 18730 325 18787 334
rect 18730 288 18751 325
rect 18833 288 18890 334
rect 18936 325 18993 334
rect 18936 288 18962 325
rect 19039 288 19096 334
rect 19142 325 19199 334
rect 19142 288 19173 325
rect 19449 288 19474 334
rect 18502 273 18540 288
rect 18592 273 18751 288
rect 18803 273 18962 288
rect 19014 273 19173 288
rect 19225 273 19384 288
rect 19436 273 19474 288
rect 14202 201 14409 247
rect 14455 201 14522 247
rect 14568 201 14635 247
rect 14681 201 14748 247
rect 14794 201 14861 247
rect 14907 201 14920 247
rect 18502 233 19474 273
rect 20632 250 20940 290
rect 20632 247 20670 250
rect 20722 247 20850 250
rect 20902 247 20940 250
rect 12959 164 13121 171
rect 12959 118 12970 164
rect 13110 118 13121 164
rect 12959 107 13121 118
rect 15181 187 18143 223
rect 20051 201 20064 247
rect 20110 201 20168 247
rect 20214 201 20271 247
rect 20317 201 20374 247
rect 20420 201 20477 247
rect 20523 201 20580 247
rect 20626 201 20670 247
rect 20729 201 20786 247
rect 20832 201 20850 247
rect 20935 201 20992 247
rect 21038 201 21051 247
rect 15181 141 15216 187
rect 15262 141 15374 187
rect 15420 141 15532 187
rect 15578 141 15690 187
rect 15736 141 15848 187
rect 15894 141 16006 187
rect 16052 141 16165 187
rect 16211 141 16323 187
rect 16369 141 16481 187
rect 16527 141 16639 187
rect 16685 141 16797 187
rect 16843 141 16955 187
rect 17001 141 17113 187
rect 17159 141 17272 187
rect 17318 141 17430 187
rect 17476 141 17588 187
rect 17634 141 17746 187
rect 17792 141 17904 187
rect 17950 141 18062 187
rect 18108 141 18143 187
rect 20632 198 20670 201
rect 20722 198 20850 201
rect 20902 198 20940 201
rect 20632 157 20940 198
rect 21186 173 21197 595
rect 21243 173 21254 595
rect 23682 522 23974 754
rect 23182 471 23974 522
rect 21386 425 21399 471
rect 23373 425 23974 471
rect 23182 403 23974 425
rect 23682 311 23974 403
rect 21394 257 21702 297
rect 21394 247 21432 257
rect 21484 247 21612 257
rect 21664 247 21702 257
rect 23682 265 23820 311
rect 23866 265 23974 311
rect 21386 201 21399 247
rect 23373 201 23386 247
rect 21186 162 21254 173
rect 21394 164 21702 201
rect 9812 60 10120 66
rect 10385 60 12583 74
rect 13350 60 14111 67
rect 9089 37 12583 60
rect 13301 37 14111 60
rect 9089 26 14111 37
rect 9089 23 9850 26
rect 9089 -23 9337 23
rect 9383 -23 9459 23
rect 9505 -23 9582 23
rect 9628 -23 9705 23
rect 9751 -23 9850 23
rect 9089 -26 9850 -23
rect 9902 -26 10030 26
rect 10082 23 13387 26
rect 10082 -23 10433 23
rect 10479 -23 10591 23
rect 10637 -23 10749 23
rect 10795 -23 10907 23
rect 10953 -23 11066 23
rect 11112 -23 11224 23
rect 11270 -23 11382 23
rect 11428 -23 11540 23
rect 11586 -23 11698 23
rect 11744 -23 11856 23
rect 11902 -23 12015 23
rect 12061 -23 12173 23
rect 12219 -23 12331 23
rect 12377 -23 12489 23
rect 12535 -23 13336 23
rect 13382 -23 13387 23
rect 10082 -26 13387 -23
rect 13439 23 13598 26
rect 13439 -23 13503 23
rect 13549 -23 13598 23
rect 13439 -26 13598 -23
rect 13650 23 13810 26
rect 13862 23 14021 26
rect 13650 -23 13668 23
rect 13714 -23 13810 23
rect 13879 -23 14021 23
rect 13650 -26 13810 -23
rect 13862 -26 14021 -23
rect 14073 -26 14111 26
rect 9089 -37 14111 -26
rect 9089 -60 12583 -37
rect 13301 -60 14111 -37
rect 7543 -67 7921 -66
rect 8611 -67 8919 -60
rect 9812 -67 10120 -60
rect 10385 -74 12583 -60
rect 13350 -66 14111 -60
rect 14393 60 14943 67
rect 15181 60 18143 141
rect 23682 147 23974 265
rect 23682 101 23820 147
rect 23866 101 23974 147
rect 23682 67 23974 101
rect 18397 60 19579 67
rect 19905 60 20456 67
rect 14393 26 19579 60
rect 14393 23 14431 26
rect 14483 23 14642 26
rect 14694 23 14853 26
rect 14905 23 18435 26
rect 14393 -23 14409 23
rect 14483 -23 14522 23
rect 14568 -23 14635 23
rect 14694 -23 14748 23
rect 14794 -23 14853 23
rect 14907 -23 15216 23
rect 15262 -23 15374 23
rect 15420 -23 15532 23
rect 15578 -23 15690 23
rect 15736 -23 15848 23
rect 15894 -23 16006 23
rect 16052 -23 16165 23
rect 16211 -23 16323 23
rect 16369 -23 16481 23
rect 16527 -23 16639 23
rect 16685 -23 16797 23
rect 16843 -23 16955 23
rect 17001 -23 17113 23
rect 17159 -23 17272 23
rect 17318 -23 17430 23
rect 17476 -23 17588 23
rect 17634 -23 17746 23
rect 17792 -23 17904 23
rect 17950 -23 18062 23
rect 18108 -23 18435 23
rect 14393 -26 14431 -23
rect 14483 -26 14642 -23
rect 14694 -26 14853 -23
rect 14905 -26 18435 -23
rect 18487 -26 18645 26
rect 18697 -26 18856 26
rect 18908 -26 19068 26
rect 19120 -26 19279 26
rect 19331 -26 19489 26
rect 19541 -26 19579 26
rect 14393 -60 19579 -26
rect 19904 26 20456 60
rect 19904 -26 19943 26
rect 19995 23 20154 26
rect 20206 23 20365 26
rect 20417 23 20456 26
rect 21875 26 23974 67
rect 21875 23 21913 26
rect 21965 23 22124 26
rect 22176 23 22335 26
rect 22387 23 22545 26
rect 22597 23 22756 26
rect 22808 23 22968 26
rect 23020 23 23179 26
rect 23231 23 23389 26
rect 19995 -23 20064 23
rect 20110 -23 20154 23
rect 20214 -23 20271 23
rect 20317 -23 20365 23
rect 20420 -23 20477 23
rect 20523 -23 20580 23
rect 20626 -23 20683 23
rect 20729 -23 20786 23
rect 20832 -23 20889 23
rect 20935 -23 20992 23
rect 21038 -23 21051 23
rect 21386 -23 21399 23
rect 23373 -23 23389 23
rect 19995 -26 20154 -23
rect 20206 -26 20365 -23
rect 20417 -26 20456 -23
rect 19904 -60 20456 -26
rect 14393 -66 14943 -60
rect 18397 -67 19579 -60
rect 19905 -67 20456 -60
rect 21875 -26 21913 -23
rect 21965 -26 22124 -23
rect 22176 -26 22335 -23
rect 22387 -26 22545 -23
rect 22597 -26 22756 -23
rect 22808 -26 22968 -23
rect 23020 -26 23179 -23
rect 23231 -26 23389 -23
rect 23441 -26 23600 26
rect 23652 -26 23811 26
rect 23863 -26 23974 26
rect 21875 -67 23974 -26
<< via1 >>
rect 451 14374 503 14426
rect 662 14374 714 14426
rect 873 14374 925 14426
rect 1083 14423 1135 14426
rect 1294 14423 1346 14426
rect 1506 14423 1558 14426
rect 1717 14423 1769 14426
rect 1927 14423 1979 14426
rect 2138 14423 2190 14426
rect 2349 14423 2401 14426
rect 3881 14423 3933 14426
rect 4092 14423 4144 14426
rect 1083 14377 1135 14423
rect 1294 14377 1346 14423
rect 1506 14377 1558 14423
rect 1717 14377 1769 14423
rect 1927 14377 1979 14423
rect 2138 14377 2190 14423
rect 2349 14377 2401 14423
rect 3881 14377 3899 14423
rect 3899 14377 3933 14423
rect 4092 14377 4105 14423
rect 4105 14377 4144 14423
rect 1083 14374 1135 14377
rect 1294 14374 1346 14377
rect 1506 14374 1558 14377
rect 1717 14374 1769 14377
rect 1927 14374 1979 14377
rect 2138 14374 2190 14377
rect 2349 14374 2401 14377
rect 3881 14374 3933 14377
rect 4092 14374 4144 14377
rect 4304 14374 4356 14426
rect 4515 14374 4567 14426
rect 4817 14374 4869 14426
rect 5027 14374 5079 14426
rect 5238 14374 5290 14426
rect 5450 14374 5502 14426
rect 5661 14374 5713 14426
rect 5871 14374 5923 14426
rect 7927 14423 7979 14426
rect 7927 14377 7979 14423
rect 7927 14374 7979 14377
rect 8138 14374 8190 14426
rect 8349 14374 8401 14426
rect 8649 14423 8701 14426
rect 8829 14423 8881 14426
rect 8649 14377 8659 14423
rect 8659 14377 8701 14423
rect 8829 14377 8863 14423
rect 8863 14377 8881 14423
rect 8649 14374 8701 14377
rect 8829 14374 8881 14377
rect 2654 14199 2706 14202
rect 2834 14199 2886 14202
rect 2654 14153 2706 14199
rect 2834 14153 2886 14199
rect 2654 14150 2706 14153
rect 2834 14150 2886 14153
rect 3416 14199 3468 14210
rect 3596 14199 3648 14210
rect 3416 14158 3430 14199
rect 3430 14158 3468 14199
rect 3596 14158 3636 14199
rect 3636 14158 3648 14199
rect 4929 14112 4981 14124
rect 5140 14112 5192 14124
rect 5351 14112 5403 14124
rect 5562 14112 5614 14124
rect 5773 14112 5825 14124
rect 7488 14112 7540 14136
rect 7668 14112 7720 14136
rect 4929 14072 4981 14112
rect 5140 14072 5177 14112
rect 5177 14072 5192 14112
rect 5351 14072 5383 14112
rect 5383 14072 5403 14112
rect 5562 14072 5589 14112
rect 5589 14072 5614 14112
rect 5773 14072 5795 14112
rect 5795 14072 5825 14112
rect 7488 14084 7506 14112
rect 7506 14084 7540 14112
rect 7668 14084 7669 14112
rect 7669 14084 7720 14112
rect 3864 13929 3899 13964
rect 3899 13929 3916 13964
rect 4044 13929 4048 13964
rect 4048 13929 4096 13964
rect 4224 13929 4255 13964
rect 4255 13929 4276 13964
rect 3864 13912 3916 13929
rect 4044 13912 4096 13929
rect 4224 13912 4276 13929
rect 2654 13751 2706 13754
rect 2834 13751 2886 13754
rect 2654 13705 2706 13751
rect 2834 13705 2886 13751
rect 2654 13702 2706 13705
rect 2834 13702 2886 13705
rect 6275 13837 6294 13889
rect 6294 13837 6327 13889
rect 6558 13888 6610 13896
rect 6769 13888 6821 13896
rect 6558 13844 6568 13888
rect 6568 13844 6610 13888
rect 6769 13844 6803 13888
rect 6803 13844 6821 13888
rect 6981 13844 7033 13896
rect 7192 13844 7244 13896
rect 9850 14374 9902 14426
rect 10030 14374 10082 14426
rect 13387 14374 13439 14426
rect 13598 14374 13650 14426
rect 13810 14423 13862 14426
rect 13810 14377 13833 14423
rect 13833 14377 13862 14423
rect 13810 14374 13862 14377
rect 14021 14374 14073 14426
rect 14431 14423 14483 14426
rect 14642 14423 14694 14426
rect 14853 14423 14905 14426
rect 14431 14377 14455 14423
rect 14455 14377 14483 14423
rect 14642 14377 14681 14423
rect 14681 14377 14694 14423
rect 14853 14377 14861 14423
rect 14861 14377 14905 14423
rect 14431 14374 14483 14377
rect 14642 14374 14694 14377
rect 14853 14374 14905 14377
rect 18435 14374 18487 14426
rect 18645 14374 18697 14426
rect 18856 14374 18908 14426
rect 19068 14374 19120 14426
rect 19279 14374 19331 14426
rect 19489 14374 19541 14426
rect 19943 14374 19995 14426
rect 20154 14423 20206 14426
rect 20365 14423 20417 14426
rect 21913 14423 21965 14426
rect 22124 14423 22176 14426
rect 22335 14423 22387 14426
rect 22545 14423 22597 14426
rect 22756 14423 22808 14426
rect 22968 14423 23020 14426
rect 23179 14423 23231 14426
rect 20154 14377 20168 14423
rect 20168 14377 20206 14423
rect 20365 14377 20374 14423
rect 20374 14377 20417 14423
rect 21913 14377 21965 14423
rect 22124 14377 22176 14423
rect 22335 14377 22387 14423
rect 22545 14377 22597 14423
rect 22756 14377 22808 14423
rect 22968 14377 23020 14423
rect 23179 14377 23231 14423
rect 20154 14374 20206 14377
rect 20365 14374 20417 14377
rect 9372 14153 9383 14188
rect 9383 14153 9424 14188
rect 9372 14136 9424 14153
rect 9591 13921 9643 13973
rect 9591 13735 9643 13787
rect 21913 14374 21965 14377
rect 22124 14374 22176 14377
rect 22335 14374 22387 14377
rect 22545 14374 22597 14377
rect 22756 14374 22808 14377
rect 22968 14374 23020 14377
rect 23179 14374 23231 14377
rect 23389 14374 23441 14426
rect 23600 14374 23652 14426
rect 23811 14374 23863 14426
rect 11532 14136 11584 14188
rect 20670 14199 20722 14202
rect 20850 14199 20902 14202
rect 12665 13905 12717 13957
rect 20670 14153 20683 14199
rect 20683 14153 20722 14199
rect 20850 14153 20889 14199
rect 20889 14153 20902 14199
rect 18540 14112 18592 14127
rect 18751 14112 18803 14127
rect 18962 14112 19014 14127
rect 19173 14112 19225 14127
rect 19384 14112 19436 14127
rect 18540 14075 18581 14112
rect 18581 14075 18592 14112
rect 18751 14075 18787 14112
rect 18787 14075 18803 14112
rect 18962 14075 18993 14112
rect 18993 14075 19014 14112
rect 19173 14075 19199 14112
rect 19199 14075 19225 14112
rect 19384 14075 19436 14112
rect 20670 14150 20722 14153
rect 20850 14150 20902 14153
rect 14536 13929 14568 13964
rect 14568 13929 14588 13964
rect 14748 13929 14794 13964
rect 14794 13929 14800 13964
rect 18193 13968 18245 14020
rect 14536 13912 14588 13929
rect 14748 13912 14800 13929
rect 15194 13810 15201 13848
rect 15201 13810 15246 13848
rect 15194 13796 15246 13810
rect 19897 13912 19949 13964
rect 20108 13929 20110 13964
rect 20110 13929 20160 13964
rect 20108 13912 20160 13929
rect 20319 13912 20371 13964
rect 18193 13750 18245 13802
rect 21432 14153 21484 14195
rect 21612 14153 21664 14195
rect 21432 14143 21484 14153
rect 21612 14143 21664 14153
rect 4929 13618 4981 13664
rect 5140 13618 5177 13664
rect 5177 13618 5192 13664
rect 5351 13618 5383 13664
rect 5383 13618 5403 13664
rect 5562 13618 5589 13664
rect 5589 13618 5614 13664
rect 5773 13618 5795 13664
rect 5795 13618 5825 13664
rect 7488 13618 7506 13662
rect 7506 13618 7540 13662
rect 7668 13618 7669 13662
rect 7669 13618 7720 13662
rect 18540 13618 18581 13664
rect 18581 13618 18592 13664
rect 18751 13618 18787 13664
rect 18787 13618 18803 13664
rect 18962 13618 18993 13664
rect 18993 13618 19014 13664
rect 19173 13618 19199 13664
rect 19199 13618 19225 13664
rect 19384 13618 19436 13664
rect 21432 13705 21484 13732
rect 21612 13705 21664 13732
rect 21432 13680 21484 13705
rect 21612 13680 21664 13705
rect 4929 13612 4981 13618
rect 5140 13612 5192 13618
rect 5351 13612 5403 13618
rect 5562 13612 5614 13618
rect 5773 13612 5825 13618
rect 7488 13610 7540 13618
rect 7668 13610 7720 13618
rect 451 13474 503 13526
rect 662 13474 714 13526
rect 873 13474 925 13526
rect 1083 13474 1135 13526
rect 1294 13474 1346 13526
rect 1506 13474 1558 13526
rect 1717 13474 1769 13526
rect 1927 13474 1979 13526
rect 2138 13474 2190 13526
rect 2349 13474 2401 13526
rect 18540 13612 18592 13618
rect 18751 13612 18803 13618
rect 18962 13612 19014 13618
rect 19173 13612 19225 13618
rect 19384 13612 19436 13618
rect 4352 13474 4404 13526
rect 4532 13523 4584 13526
rect 4532 13477 4559 13523
rect 4559 13477 4584 13523
rect 4532 13474 4584 13477
rect 19735 13523 19787 13526
rect 19735 13477 19757 13523
rect 19757 13477 19787 13523
rect 19735 13474 19787 13477
rect 19915 13474 19967 13526
rect 4929 13382 4981 13388
rect 5140 13382 5192 13388
rect 5351 13382 5403 13388
rect 5562 13382 5614 13388
rect 5773 13382 5825 13388
rect 7488 13382 7540 13390
rect 7668 13382 7720 13390
rect 21913 13474 21965 13526
rect 22124 13474 22176 13526
rect 22335 13474 22387 13526
rect 22545 13474 22597 13526
rect 22756 13474 22808 13526
rect 22968 13474 23020 13526
rect 23179 13474 23231 13526
rect 23389 13474 23441 13526
rect 23600 13474 23652 13526
rect 23811 13474 23863 13526
rect 18540 13382 18592 13388
rect 18751 13382 18803 13388
rect 18962 13382 19014 13388
rect 19173 13382 19225 13388
rect 19384 13382 19436 13388
rect 2654 13295 2706 13298
rect 2834 13295 2886 13298
rect 4929 13336 4981 13382
rect 5140 13336 5177 13382
rect 5177 13336 5192 13382
rect 5351 13336 5383 13382
rect 5383 13336 5403 13382
rect 5562 13336 5589 13382
rect 5589 13336 5614 13382
rect 5773 13336 5795 13382
rect 5795 13336 5825 13382
rect 7488 13338 7506 13382
rect 7506 13338 7540 13382
rect 7668 13338 7669 13382
rect 7669 13338 7720 13382
rect 2654 13249 2706 13295
rect 2834 13249 2886 13295
rect 2654 13246 2706 13249
rect 2834 13246 2886 13249
rect 2654 12847 2706 12850
rect 2834 12847 2886 12850
rect 2654 12801 2706 12847
rect 2834 12801 2886 12847
rect 2654 12798 2706 12801
rect 2834 12798 2886 12801
rect 3864 13071 3916 13088
rect 4044 13071 4096 13088
rect 4224 13071 4276 13088
rect 3864 13036 3899 13071
rect 3899 13036 3916 13071
rect 4044 13036 4048 13071
rect 4048 13036 4096 13071
rect 4224 13036 4255 13071
rect 4255 13036 4276 13071
rect 6275 13111 6294 13163
rect 6294 13111 6327 13163
rect 18540 13336 18581 13382
rect 18581 13336 18592 13382
rect 18751 13336 18787 13382
rect 18787 13336 18803 13382
rect 18962 13336 18993 13382
rect 18993 13336 19014 13382
rect 19173 13336 19199 13382
rect 19199 13336 19225 13382
rect 19384 13336 19436 13382
rect 9591 13213 9643 13265
rect 6558 13112 6568 13156
rect 6568 13112 6610 13156
rect 6769 13112 6803 13156
rect 6803 13112 6821 13156
rect 6558 13104 6610 13112
rect 6769 13104 6821 13112
rect 6981 13104 7033 13156
rect 7192 13104 7244 13156
rect 4929 12888 4981 12928
rect 5140 12888 5177 12928
rect 5177 12888 5192 12928
rect 5351 12888 5383 12928
rect 5383 12888 5403 12928
rect 5562 12888 5589 12928
rect 5589 12888 5614 12928
rect 5773 12888 5795 12928
rect 5795 12888 5825 12928
rect 7488 12888 7506 12916
rect 7506 12888 7540 12916
rect 7668 12888 7669 12916
rect 7669 12888 7720 12916
rect 4929 12876 4981 12888
rect 5140 12876 5192 12888
rect 5351 12876 5403 12888
rect 5562 12876 5614 12888
rect 5773 12876 5825 12888
rect 3416 12801 3430 12842
rect 3430 12801 3468 12842
rect 3596 12801 3636 12842
rect 3636 12801 3648 12842
rect 7488 12864 7540 12888
rect 7668 12864 7720 12888
rect 3416 12790 3468 12801
rect 3596 12790 3648 12801
rect 451 12574 503 12626
rect 662 12574 714 12626
rect 873 12574 925 12626
rect 1083 12623 1135 12626
rect 1294 12623 1346 12626
rect 1506 12623 1558 12626
rect 1717 12623 1769 12626
rect 1927 12623 1979 12626
rect 2138 12623 2190 12626
rect 2349 12623 2401 12626
rect 3881 12623 3933 12626
rect 4092 12623 4144 12626
rect 1083 12577 1135 12623
rect 1294 12577 1346 12623
rect 1506 12577 1558 12623
rect 1717 12577 1769 12623
rect 1927 12577 1979 12623
rect 2138 12577 2190 12623
rect 2349 12577 2401 12623
rect 3881 12577 3899 12623
rect 3899 12577 3933 12623
rect 4092 12577 4105 12623
rect 4105 12577 4144 12623
rect 1083 12574 1135 12577
rect 1294 12574 1346 12577
rect 1506 12574 1558 12577
rect 1717 12574 1769 12577
rect 1927 12574 1979 12577
rect 2138 12574 2190 12577
rect 2349 12574 2401 12577
rect 3881 12574 3933 12577
rect 4092 12574 4144 12577
rect 4304 12574 4356 12626
rect 4515 12574 4567 12626
rect 4817 12574 4869 12626
rect 5027 12574 5079 12626
rect 5238 12574 5290 12626
rect 5450 12574 5502 12626
rect 5661 12574 5713 12626
rect 5871 12574 5923 12626
rect 7927 12623 7979 12626
rect 7927 12577 7979 12623
rect 7927 12574 7979 12577
rect 8138 12574 8190 12626
rect 8349 12574 8401 12626
rect 8649 12623 8701 12626
rect 8829 12623 8881 12626
rect 8649 12577 8659 12623
rect 8659 12577 8701 12623
rect 8829 12577 8863 12623
rect 8863 12577 8881 12623
rect 8649 12574 8701 12577
rect 8829 12574 8881 12577
rect 2654 12399 2706 12402
rect 2834 12399 2886 12402
rect 2654 12353 2706 12399
rect 2834 12353 2886 12399
rect 2654 12350 2706 12353
rect 2834 12350 2886 12353
rect 3416 12399 3468 12410
rect 3596 12399 3648 12410
rect 3416 12358 3430 12399
rect 3430 12358 3468 12399
rect 3596 12358 3636 12399
rect 3636 12358 3648 12399
rect 4929 12312 4981 12324
rect 5140 12312 5192 12324
rect 5351 12312 5403 12324
rect 5562 12312 5614 12324
rect 5773 12312 5825 12324
rect 7488 12312 7540 12336
rect 7668 12312 7720 12336
rect 4929 12272 4981 12312
rect 5140 12272 5177 12312
rect 5177 12272 5192 12312
rect 5351 12272 5383 12312
rect 5383 12272 5403 12312
rect 5562 12272 5589 12312
rect 5589 12272 5614 12312
rect 5773 12272 5795 12312
rect 5795 12272 5825 12312
rect 7488 12284 7506 12312
rect 7506 12284 7540 12312
rect 7668 12284 7669 12312
rect 7669 12284 7720 12312
rect 3864 12129 3899 12164
rect 3899 12129 3916 12164
rect 4044 12129 4048 12164
rect 4048 12129 4096 12164
rect 4224 12129 4255 12164
rect 4255 12129 4276 12164
rect 3864 12112 3916 12129
rect 4044 12112 4096 12129
rect 4224 12112 4276 12129
rect 2654 11951 2706 11954
rect 2834 11951 2886 11954
rect 2654 11905 2706 11951
rect 2834 11905 2886 11951
rect 2654 11902 2706 11905
rect 2834 11902 2886 11905
rect 6275 12037 6294 12089
rect 6294 12037 6327 12089
rect 6558 12088 6610 12096
rect 6769 12088 6821 12096
rect 6558 12044 6568 12088
rect 6568 12044 6610 12088
rect 6769 12044 6803 12088
rect 6803 12044 6821 12088
rect 6981 12044 7033 12096
rect 7192 12044 7244 12096
rect 9591 13027 9643 13079
rect 9372 12847 9424 12864
rect 9372 12812 9383 12847
rect 9383 12812 9424 12847
rect 12665 13043 12717 13095
rect 11532 12812 11584 12864
rect 15572 13152 15624 13204
rect 18193 13198 18245 13250
rect 21432 13295 21484 13320
rect 21612 13295 21664 13320
rect 21432 13268 21484 13295
rect 21612 13268 21664 13295
rect 14536 13071 14588 13088
rect 14748 13071 14800 13088
rect 14536 13036 14568 13071
rect 14568 13036 14588 13071
rect 14748 13036 14794 13071
rect 14794 13036 14800 13071
rect 18193 12980 18245 13032
rect 19897 13036 19949 13088
rect 20108 13071 20160 13088
rect 20108 13036 20110 13071
rect 20110 13036 20160 13071
rect 20319 13036 20371 13088
rect 18540 12888 18581 12925
rect 18581 12888 18592 12925
rect 18751 12888 18787 12925
rect 18787 12888 18803 12925
rect 18962 12888 18993 12925
rect 18993 12888 19014 12925
rect 19173 12888 19199 12925
rect 19199 12888 19225 12925
rect 19384 12888 19436 12925
rect 18540 12873 18592 12888
rect 18751 12873 18803 12888
rect 18962 12873 19014 12888
rect 19173 12873 19225 12888
rect 19384 12873 19436 12888
rect 20670 12847 20722 12850
rect 20850 12847 20902 12850
rect 20670 12801 20683 12847
rect 20683 12801 20722 12847
rect 20850 12801 20889 12847
rect 20889 12801 20902 12847
rect 20670 12798 20722 12801
rect 20850 12798 20902 12801
rect 21432 12847 21484 12857
rect 21612 12847 21664 12857
rect 21432 12805 21484 12847
rect 21612 12805 21664 12847
rect 9850 12574 9902 12626
rect 10030 12574 10082 12626
rect 13387 12574 13439 12626
rect 13598 12574 13650 12626
rect 13810 12623 13862 12626
rect 13810 12577 13833 12623
rect 13833 12577 13862 12623
rect 13810 12574 13862 12577
rect 14021 12574 14073 12626
rect 14431 12623 14483 12626
rect 14642 12623 14694 12626
rect 14853 12623 14905 12626
rect 14431 12577 14455 12623
rect 14455 12577 14483 12623
rect 14642 12577 14681 12623
rect 14681 12577 14694 12623
rect 14853 12577 14861 12623
rect 14861 12577 14905 12623
rect 14431 12574 14483 12577
rect 14642 12574 14694 12577
rect 14853 12574 14905 12577
rect 18435 12574 18487 12626
rect 18645 12574 18697 12626
rect 18856 12574 18908 12626
rect 19068 12574 19120 12626
rect 19279 12574 19331 12626
rect 19489 12574 19541 12626
rect 19943 12574 19995 12626
rect 20154 12623 20206 12626
rect 20365 12623 20417 12626
rect 21913 12623 21965 12626
rect 22124 12623 22176 12626
rect 22335 12623 22387 12626
rect 22545 12623 22597 12626
rect 22756 12623 22808 12626
rect 22968 12623 23020 12626
rect 23179 12623 23231 12626
rect 20154 12577 20168 12623
rect 20168 12577 20206 12623
rect 20365 12577 20374 12623
rect 20374 12577 20417 12623
rect 21913 12577 21965 12623
rect 22124 12577 22176 12623
rect 22335 12577 22387 12623
rect 22545 12577 22597 12623
rect 22756 12577 22808 12623
rect 22968 12577 23020 12623
rect 23179 12577 23231 12623
rect 20154 12574 20206 12577
rect 20365 12574 20417 12577
rect 9372 12353 9383 12388
rect 9383 12353 9424 12388
rect 9372 12336 9424 12353
rect 9591 12121 9643 12173
rect 9591 11935 9643 11987
rect 21913 12574 21965 12577
rect 22124 12574 22176 12577
rect 22335 12574 22387 12577
rect 22545 12574 22597 12577
rect 22756 12574 22808 12577
rect 22968 12574 23020 12577
rect 23179 12574 23231 12577
rect 23389 12574 23441 12626
rect 23600 12574 23652 12626
rect 23811 12574 23863 12626
rect 11532 12336 11584 12388
rect 20670 12399 20722 12402
rect 20850 12399 20902 12402
rect 12665 12105 12717 12157
rect 20670 12353 20683 12399
rect 20683 12353 20722 12399
rect 20850 12353 20889 12399
rect 20889 12353 20902 12399
rect 18540 12312 18592 12327
rect 18751 12312 18803 12327
rect 18962 12312 19014 12327
rect 19173 12312 19225 12327
rect 19384 12312 19436 12327
rect 18540 12275 18581 12312
rect 18581 12275 18592 12312
rect 18751 12275 18787 12312
rect 18787 12275 18803 12312
rect 18962 12275 18993 12312
rect 18993 12275 19014 12312
rect 19173 12275 19199 12312
rect 19199 12275 19225 12312
rect 19384 12275 19436 12312
rect 20670 12350 20722 12353
rect 20850 12350 20902 12353
rect 14536 12129 14568 12164
rect 14568 12129 14588 12164
rect 14748 12129 14794 12164
rect 14794 12129 14800 12164
rect 18193 12168 18245 12220
rect 14536 12112 14588 12129
rect 14748 12112 14800 12129
rect 15950 11996 16002 12048
rect 19897 12112 19949 12164
rect 20108 12129 20110 12164
rect 20110 12129 20160 12164
rect 20108 12112 20160 12129
rect 20319 12112 20371 12164
rect 18193 11950 18245 12002
rect 21432 12353 21484 12395
rect 21612 12353 21664 12395
rect 21432 12343 21484 12353
rect 21612 12343 21664 12353
rect 4929 11818 4981 11864
rect 5140 11818 5177 11864
rect 5177 11818 5192 11864
rect 5351 11818 5383 11864
rect 5383 11818 5403 11864
rect 5562 11818 5589 11864
rect 5589 11818 5614 11864
rect 5773 11818 5795 11864
rect 5795 11818 5825 11864
rect 7488 11818 7506 11862
rect 7506 11818 7540 11862
rect 7668 11818 7669 11862
rect 7669 11818 7720 11862
rect 18540 11818 18581 11864
rect 18581 11818 18592 11864
rect 18751 11818 18787 11864
rect 18787 11818 18803 11864
rect 18962 11818 18993 11864
rect 18993 11818 19014 11864
rect 19173 11818 19199 11864
rect 19199 11818 19225 11864
rect 19384 11818 19436 11864
rect 21432 11905 21484 11932
rect 21612 11905 21664 11932
rect 21432 11880 21484 11905
rect 21612 11880 21664 11905
rect 4929 11812 4981 11818
rect 5140 11812 5192 11818
rect 5351 11812 5403 11818
rect 5562 11812 5614 11818
rect 5773 11812 5825 11818
rect 7488 11810 7540 11818
rect 7668 11810 7720 11818
rect 451 11674 503 11726
rect 662 11674 714 11726
rect 873 11674 925 11726
rect 1083 11674 1135 11726
rect 1294 11674 1346 11726
rect 1506 11674 1558 11726
rect 1717 11674 1769 11726
rect 1927 11674 1979 11726
rect 2138 11674 2190 11726
rect 2349 11674 2401 11726
rect 18540 11812 18592 11818
rect 18751 11812 18803 11818
rect 18962 11812 19014 11818
rect 19173 11812 19225 11818
rect 19384 11812 19436 11818
rect 4352 11674 4404 11726
rect 4532 11723 4584 11726
rect 4532 11677 4559 11723
rect 4559 11677 4584 11723
rect 4532 11674 4584 11677
rect 19735 11723 19787 11726
rect 19735 11677 19757 11723
rect 19757 11677 19787 11723
rect 19735 11674 19787 11677
rect 19915 11674 19967 11726
rect 4929 11582 4981 11588
rect 5140 11582 5192 11588
rect 5351 11582 5403 11588
rect 5562 11582 5614 11588
rect 5773 11582 5825 11588
rect 7488 11582 7540 11590
rect 7668 11582 7720 11590
rect 21913 11674 21965 11726
rect 22124 11674 22176 11726
rect 22335 11674 22387 11726
rect 22545 11674 22597 11726
rect 22756 11674 22808 11726
rect 22968 11674 23020 11726
rect 23179 11674 23231 11726
rect 23389 11674 23441 11726
rect 23600 11674 23652 11726
rect 23811 11674 23863 11726
rect 18540 11582 18592 11588
rect 18751 11582 18803 11588
rect 18962 11582 19014 11588
rect 19173 11582 19225 11588
rect 19384 11582 19436 11588
rect 2654 11495 2706 11498
rect 2834 11495 2886 11498
rect 4929 11536 4981 11582
rect 5140 11536 5177 11582
rect 5177 11536 5192 11582
rect 5351 11536 5383 11582
rect 5383 11536 5403 11582
rect 5562 11536 5589 11582
rect 5589 11536 5614 11582
rect 5773 11536 5795 11582
rect 5795 11536 5825 11582
rect 7488 11538 7506 11582
rect 7506 11538 7540 11582
rect 7668 11538 7669 11582
rect 7669 11538 7720 11582
rect 2654 11449 2706 11495
rect 2834 11449 2886 11495
rect 2654 11446 2706 11449
rect 2834 11446 2886 11449
rect 2654 11047 2706 11050
rect 2834 11047 2886 11050
rect 2654 11001 2706 11047
rect 2834 11001 2886 11047
rect 2654 10998 2706 11001
rect 2834 10998 2886 11001
rect 3864 11271 3916 11288
rect 4044 11271 4096 11288
rect 4224 11271 4276 11288
rect 3864 11236 3899 11271
rect 3899 11236 3916 11271
rect 4044 11236 4048 11271
rect 4048 11236 4096 11271
rect 4224 11236 4255 11271
rect 4255 11236 4276 11271
rect 6275 11311 6294 11363
rect 6294 11311 6327 11363
rect 18540 11536 18581 11582
rect 18581 11536 18592 11582
rect 18751 11536 18787 11582
rect 18787 11536 18803 11582
rect 18962 11536 18993 11582
rect 18993 11536 19014 11582
rect 19173 11536 19199 11582
rect 19199 11536 19225 11582
rect 19384 11536 19436 11582
rect 9591 11413 9643 11465
rect 6558 11312 6568 11356
rect 6568 11312 6610 11356
rect 6769 11312 6803 11356
rect 6803 11312 6821 11356
rect 6558 11304 6610 11312
rect 6769 11304 6821 11312
rect 6981 11304 7033 11356
rect 7192 11304 7244 11356
rect 4929 11088 4981 11128
rect 5140 11088 5177 11128
rect 5177 11088 5192 11128
rect 5351 11088 5383 11128
rect 5383 11088 5403 11128
rect 5562 11088 5589 11128
rect 5589 11088 5614 11128
rect 5773 11088 5795 11128
rect 5795 11088 5825 11128
rect 7488 11088 7506 11116
rect 7506 11088 7540 11116
rect 7668 11088 7669 11116
rect 7669 11088 7720 11116
rect 4929 11076 4981 11088
rect 5140 11076 5192 11088
rect 5351 11076 5403 11088
rect 5562 11076 5614 11088
rect 5773 11076 5825 11088
rect 3416 11001 3430 11042
rect 3430 11001 3468 11042
rect 3596 11001 3636 11042
rect 3636 11001 3648 11042
rect 7488 11064 7540 11088
rect 7668 11064 7720 11088
rect 3416 10990 3468 11001
rect 3596 10990 3648 11001
rect 451 10774 503 10826
rect 662 10774 714 10826
rect 873 10774 925 10826
rect 1083 10823 1135 10826
rect 1294 10823 1346 10826
rect 1506 10823 1558 10826
rect 1717 10823 1769 10826
rect 1927 10823 1979 10826
rect 2138 10823 2190 10826
rect 2349 10823 2401 10826
rect 3881 10823 3933 10826
rect 4092 10823 4144 10826
rect 1083 10777 1135 10823
rect 1294 10777 1346 10823
rect 1506 10777 1558 10823
rect 1717 10777 1769 10823
rect 1927 10777 1979 10823
rect 2138 10777 2190 10823
rect 2349 10777 2401 10823
rect 3881 10777 3899 10823
rect 3899 10777 3933 10823
rect 4092 10777 4105 10823
rect 4105 10777 4144 10823
rect 1083 10774 1135 10777
rect 1294 10774 1346 10777
rect 1506 10774 1558 10777
rect 1717 10774 1769 10777
rect 1927 10774 1979 10777
rect 2138 10774 2190 10777
rect 2349 10774 2401 10777
rect 3881 10774 3933 10777
rect 4092 10774 4144 10777
rect 4304 10774 4356 10826
rect 4515 10774 4567 10826
rect 4817 10774 4869 10826
rect 5027 10774 5079 10826
rect 5238 10774 5290 10826
rect 5450 10774 5502 10826
rect 5661 10774 5713 10826
rect 5871 10774 5923 10826
rect 7927 10823 7979 10826
rect 7927 10777 7979 10823
rect 7927 10774 7979 10777
rect 8138 10774 8190 10826
rect 8349 10774 8401 10826
rect 8649 10823 8701 10826
rect 8829 10823 8881 10826
rect 8649 10777 8659 10823
rect 8659 10777 8701 10823
rect 8829 10777 8863 10823
rect 8863 10777 8881 10823
rect 8649 10774 8701 10777
rect 8829 10774 8881 10777
rect 2654 10599 2706 10602
rect 2834 10599 2886 10602
rect 2654 10553 2706 10599
rect 2834 10553 2886 10599
rect 2654 10550 2706 10553
rect 2834 10550 2886 10553
rect 3416 10599 3468 10610
rect 3596 10599 3648 10610
rect 3416 10558 3430 10599
rect 3430 10558 3468 10599
rect 3596 10558 3636 10599
rect 3636 10558 3648 10599
rect 4929 10512 4981 10524
rect 5140 10512 5192 10524
rect 5351 10512 5403 10524
rect 5562 10512 5614 10524
rect 5773 10512 5825 10524
rect 7488 10512 7540 10536
rect 7668 10512 7720 10536
rect 4929 10472 4981 10512
rect 5140 10472 5177 10512
rect 5177 10472 5192 10512
rect 5351 10472 5383 10512
rect 5383 10472 5403 10512
rect 5562 10472 5589 10512
rect 5589 10472 5614 10512
rect 5773 10472 5795 10512
rect 5795 10472 5825 10512
rect 7488 10484 7506 10512
rect 7506 10484 7540 10512
rect 7668 10484 7669 10512
rect 7669 10484 7720 10512
rect 3864 10329 3899 10364
rect 3899 10329 3916 10364
rect 4044 10329 4048 10364
rect 4048 10329 4096 10364
rect 4224 10329 4255 10364
rect 4255 10329 4276 10364
rect 3864 10312 3916 10329
rect 4044 10312 4096 10329
rect 4224 10312 4276 10329
rect 2654 10151 2706 10154
rect 2834 10151 2886 10154
rect 2654 10105 2706 10151
rect 2834 10105 2886 10151
rect 2654 10102 2706 10105
rect 2834 10102 2886 10105
rect 6275 10237 6294 10289
rect 6294 10237 6327 10289
rect 6558 10288 6610 10296
rect 6769 10288 6821 10296
rect 6558 10244 6568 10288
rect 6568 10244 6610 10288
rect 6769 10244 6803 10288
rect 6803 10244 6821 10288
rect 6981 10244 7033 10296
rect 7192 10244 7244 10296
rect 9591 11227 9643 11279
rect 9372 11047 9424 11064
rect 9372 11012 9383 11047
rect 9383 11012 9424 11047
rect 12665 11243 12717 11295
rect 11532 11012 11584 11064
rect 16328 11352 16380 11404
rect 18193 11398 18245 11450
rect 21432 11495 21484 11520
rect 21612 11495 21664 11520
rect 21432 11468 21484 11495
rect 21612 11468 21664 11495
rect 14536 11271 14588 11288
rect 14748 11271 14800 11288
rect 14536 11236 14568 11271
rect 14568 11236 14588 11271
rect 14748 11236 14794 11271
rect 14794 11236 14800 11271
rect 18193 11180 18245 11232
rect 19897 11236 19949 11288
rect 20108 11271 20160 11288
rect 20108 11236 20110 11271
rect 20110 11236 20160 11271
rect 20319 11236 20371 11288
rect 18540 11088 18581 11125
rect 18581 11088 18592 11125
rect 18751 11088 18787 11125
rect 18787 11088 18803 11125
rect 18962 11088 18993 11125
rect 18993 11088 19014 11125
rect 19173 11088 19199 11125
rect 19199 11088 19225 11125
rect 19384 11088 19436 11125
rect 18540 11073 18592 11088
rect 18751 11073 18803 11088
rect 18962 11073 19014 11088
rect 19173 11073 19225 11088
rect 19384 11073 19436 11088
rect 20670 11047 20722 11050
rect 20850 11047 20902 11050
rect 20670 11001 20683 11047
rect 20683 11001 20722 11047
rect 20850 11001 20889 11047
rect 20889 11001 20902 11047
rect 20670 10998 20722 11001
rect 20850 10998 20902 11001
rect 21432 11047 21484 11057
rect 21612 11047 21664 11057
rect 21432 11005 21484 11047
rect 21612 11005 21664 11047
rect 9850 10774 9902 10826
rect 10030 10774 10082 10826
rect 13387 10774 13439 10826
rect 13598 10774 13650 10826
rect 13810 10823 13862 10826
rect 13810 10777 13833 10823
rect 13833 10777 13862 10823
rect 13810 10774 13862 10777
rect 14021 10774 14073 10826
rect 14431 10823 14483 10826
rect 14642 10823 14694 10826
rect 14853 10823 14905 10826
rect 14431 10777 14455 10823
rect 14455 10777 14483 10823
rect 14642 10777 14681 10823
rect 14681 10777 14694 10823
rect 14853 10777 14861 10823
rect 14861 10777 14905 10823
rect 14431 10774 14483 10777
rect 14642 10774 14694 10777
rect 14853 10774 14905 10777
rect 18435 10774 18487 10826
rect 18645 10774 18697 10826
rect 18856 10774 18908 10826
rect 19068 10774 19120 10826
rect 19279 10774 19331 10826
rect 19489 10774 19541 10826
rect 19943 10774 19995 10826
rect 20154 10823 20206 10826
rect 20365 10823 20417 10826
rect 21913 10823 21965 10826
rect 22124 10823 22176 10826
rect 22335 10823 22387 10826
rect 22545 10823 22597 10826
rect 22756 10823 22808 10826
rect 22968 10823 23020 10826
rect 23179 10823 23231 10826
rect 20154 10777 20168 10823
rect 20168 10777 20206 10823
rect 20365 10777 20374 10823
rect 20374 10777 20417 10823
rect 21913 10777 21965 10823
rect 22124 10777 22176 10823
rect 22335 10777 22387 10823
rect 22545 10777 22597 10823
rect 22756 10777 22808 10823
rect 22968 10777 23020 10823
rect 23179 10777 23231 10823
rect 20154 10774 20206 10777
rect 20365 10774 20417 10777
rect 9372 10553 9383 10588
rect 9383 10553 9424 10588
rect 9372 10536 9424 10553
rect 9591 10321 9643 10373
rect 9591 10135 9643 10187
rect 21913 10774 21965 10777
rect 22124 10774 22176 10777
rect 22335 10774 22387 10777
rect 22545 10774 22597 10777
rect 22756 10774 22808 10777
rect 22968 10774 23020 10777
rect 23179 10774 23231 10777
rect 23389 10774 23441 10826
rect 23600 10774 23652 10826
rect 23811 10774 23863 10826
rect 11532 10536 11584 10588
rect 20670 10599 20722 10602
rect 20850 10599 20902 10602
rect 12665 10305 12717 10357
rect 20670 10553 20683 10599
rect 20683 10553 20722 10599
rect 20850 10553 20889 10599
rect 20889 10553 20902 10599
rect 18540 10512 18592 10527
rect 18751 10512 18803 10527
rect 18962 10512 19014 10527
rect 19173 10512 19225 10527
rect 19384 10512 19436 10527
rect 18540 10475 18581 10512
rect 18581 10475 18592 10512
rect 18751 10475 18787 10512
rect 18787 10475 18803 10512
rect 18962 10475 18993 10512
rect 18993 10475 19014 10512
rect 19173 10475 19199 10512
rect 19199 10475 19225 10512
rect 19384 10475 19436 10512
rect 20670 10550 20722 10553
rect 20850 10550 20902 10553
rect 14536 10329 14568 10364
rect 14568 10329 14588 10364
rect 14748 10329 14794 10364
rect 14794 10329 14800 10364
rect 18193 10368 18245 10420
rect 14536 10312 14588 10329
rect 14748 10312 14800 10329
rect 16705 10196 16757 10248
rect 19897 10312 19949 10364
rect 20108 10329 20110 10364
rect 20110 10329 20160 10364
rect 20108 10312 20160 10329
rect 20319 10312 20371 10364
rect 18193 10150 18245 10202
rect 21432 10553 21484 10595
rect 21612 10553 21664 10595
rect 21432 10543 21484 10553
rect 21612 10543 21664 10553
rect 4929 10018 4981 10064
rect 5140 10018 5177 10064
rect 5177 10018 5192 10064
rect 5351 10018 5383 10064
rect 5383 10018 5403 10064
rect 5562 10018 5589 10064
rect 5589 10018 5614 10064
rect 5773 10018 5795 10064
rect 5795 10018 5825 10064
rect 7488 10018 7506 10062
rect 7506 10018 7540 10062
rect 7668 10018 7669 10062
rect 7669 10018 7720 10062
rect 18540 10018 18581 10064
rect 18581 10018 18592 10064
rect 18751 10018 18787 10064
rect 18787 10018 18803 10064
rect 18962 10018 18993 10064
rect 18993 10018 19014 10064
rect 19173 10018 19199 10064
rect 19199 10018 19225 10064
rect 19384 10018 19436 10064
rect 21432 10105 21484 10132
rect 21612 10105 21664 10132
rect 21432 10080 21484 10105
rect 21612 10080 21664 10105
rect 4929 10012 4981 10018
rect 5140 10012 5192 10018
rect 5351 10012 5403 10018
rect 5562 10012 5614 10018
rect 5773 10012 5825 10018
rect 7488 10010 7540 10018
rect 7668 10010 7720 10018
rect 451 9874 503 9926
rect 662 9874 714 9926
rect 873 9874 925 9926
rect 1083 9874 1135 9926
rect 1294 9874 1346 9926
rect 1506 9874 1558 9926
rect 1717 9874 1769 9926
rect 1927 9874 1979 9926
rect 2138 9874 2190 9926
rect 2349 9874 2401 9926
rect 18540 10012 18592 10018
rect 18751 10012 18803 10018
rect 18962 10012 19014 10018
rect 19173 10012 19225 10018
rect 19384 10012 19436 10018
rect 4352 9874 4404 9926
rect 4532 9923 4584 9926
rect 4532 9877 4559 9923
rect 4559 9877 4584 9923
rect 4532 9874 4584 9877
rect 19735 9923 19787 9926
rect 19735 9877 19757 9923
rect 19757 9877 19787 9923
rect 19735 9874 19787 9877
rect 19915 9874 19967 9926
rect 4929 9782 4981 9788
rect 5140 9782 5192 9788
rect 5351 9782 5403 9788
rect 5562 9782 5614 9788
rect 5773 9782 5825 9788
rect 7488 9782 7540 9790
rect 7668 9782 7720 9790
rect 21913 9874 21965 9926
rect 22124 9874 22176 9926
rect 22335 9874 22387 9926
rect 22545 9874 22597 9926
rect 22756 9874 22808 9926
rect 22968 9874 23020 9926
rect 23179 9874 23231 9926
rect 23389 9874 23441 9926
rect 23600 9874 23652 9926
rect 23811 9874 23863 9926
rect 18540 9782 18592 9788
rect 18751 9782 18803 9788
rect 18962 9782 19014 9788
rect 19173 9782 19225 9788
rect 19384 9782 19436 9788
rect 2654 9695 2706 9698
rect 2834 9695 2886 9698
rect 4929 9736 4981 9782
rect 5140 9736 5177 9782
rect 5177 9736 5192 9782
rect 5351 9736 5383 9782
rect 5383 9736 5403 9782
rect 5562 9736 5589 9782
rect 5589 9736 5614 9782
rect 5773 9736 5795 9782
rect 5795 9736 5825 9782
rect 7488 9738 7506 9782
rect 7506 9738 7540 9782
rect 7668 9738 7669 9782
rect 7669 9738 7720 9782
rect 2654 9649 2706 9695
rect 2834 9649 2886 9695
rect 2654 9646 2706 9649
rect 2834 9646 2886 9649
rect 2654 9247 2706 9250
rect 2834 9247 2886 9250
rect 2654 9201 2706 9247
rect 2834 9201 2886 9247
rect 2654 9198 2706 9201
rect 2834 9198 2886 9201
rect 3864 9471 3916 9488
rect 4044 9471 4096 9488
rect 4224 9471 4276 9488
rect 3864 9436 3899 9471
rect 3899 9436 3916 9471
rect 4044 9436 4048 9471
rect 4048 9436 4096 9471
rect 4224 9436 4255 9471
rect 4255 9436 4276 9471
rect 6275 9511 6294 9563
rect 6294 9511 6327 9563
rect 18540 9736 18581 9782
rect 18581 9736 18592 9782
rect 18751 9736 18787 9782
rect 18787 9736 18803 9782
rect 18962 9736 18993 9782
rect 18993 9736 19014 9782
rect 19173 9736 19199 9782
rect 19199 9736 19225 9782
rect 19384 9736 19436 9782
rect 9591 9613 9643 9665
rect 6558 9512 6568 9556
rect 6568 9512 6610 9556
rect 6769 9512 6803 9556
rect 6803 9512 6821 9556
rect 6558 9504 6610 9512
rect 6769 9504 6821 9512
rect 6981 9504 7033 9556
rect 7192 9504 7244 9556
rect 4929 9288 4981 9328
rect 5140 9288 5177 9328
rect 5177 9288 5192 9328
rect 5351 9288 5383 9328
rect 5383 9288 5403 9328
rect 5562 9288 5589 9328
rect 5589 9288 5614 9328
rect 5773 9288 5795 9328
rect 5795 9288 5825 9328
rect 7488 9288 7506 9316
rect 7506 9288 7540 9316
rect 7668 9288 7669 9316
rect 7669 9288 7720 9316
rect 4929 9276 4981 9288
rect 5140 9276 5192 9288
rect 5351 9276 5403 9288
rect 5562 9276 5614 9288
rect 5773 9276 5825 9288
rect 3416 9201 3430 9242
rect 3430 9201 3468 9242
rect 3596 9201 3636 9242
rect 3636 9201 3648 9242
rect 7488 9264 7540 9288
rect 7668 9264 7720 9288
rect 3416 9190 3468 9201
rect 3596 9190 3648 9201
rect 451 8974 503 9026
rect 662 8974 714 9026
rect 873 8974 925 9026
rect 1083 9023 1135 9026
rect 1294 9023 1346 9026
rect 1506 9023 1558 9026
rect 1717 9023 1769 9026
rect 1927 9023 1979 9026
rect 2138 9023 2190 9026
rect 2349 9023 2401 9026
rect 3881 9023 3933 9026
rect 4092 9023 4144 9026
rect 1083 8977 1135 9023
rect 1294 8977 1346 9023
rect 1506 8977 1558 9023
rect 1717 8977 1769 9023
rect 1927 8977 1979 9023
rect 2138 8977 2190 9023
rect 2349 8977 2401 9023
rect 3881 8977 3899 9023
rect 3899 8977 3933 9023
rect 4092 8977 4105 9023
rect 4105 8977 4144 9023
rect 1083 8974 1135 8977
rect 1294 8974 1346 8977
rect 1506 8974 1558 8977
rect 1717 8974 1769 8977
rect 1927 8974 1979 8977
rect 2138 8974 2190 8977
rect 2349 8974 2401 8977
rect 3881 8974 3933 8977
rect 4092 8974 4144 8977
rect 4304 8974 4356 9026
rect 4515 8974 4567 9026
rect 4817 8974 4869 9026
rect 5027 8974 5079 9026
rect 5238 8974 5290 9026
rect 5450 8974 5502 9026
rect 5661 8974 5713 9026
rect 5871 8974 5923 9026
rect 7927 9023 7979 9026
rect 7927 8977 7979 9023
rect 7927 8974 7979 8977
rect 8138 8974 8190 9026
rect 8349 8974 8401 9026
rect 8649 9023 8701 9026
rect 8829 9023 8881 9026
rect 8649 8977 8659 9023
rect 8659 8977 8701 9023
rect 8829 8977 8863 9023
rect 8863 8977 8881 9023
rect 8649 8974 8701 8977
rect 8829 8974 8881 8977
rect 2654 8799 2706 8802
rect 2834 8799 2886 8802
rect 2654 8753 2706 8799
rect 2834 8753 2886 8799
rect 2654 8750 2706 8753
rect 2834 8750 2886 8753
rect 3416 8799 3468 8810
rect 3596 8799 3648 8810
rect 3416 8758 3430 8799
rect 3430 8758 3468 8799
rect 3596 8758 3636 8799
rect 3636 8758 3648 8799
rect 4929 8712 4981 8724
rect 5140 8712 5192 8724
rect 5351 8712 5403 8724
rect 5562 8712 5614 8724
rect 5773 8712 5825 8724
rect 7488 8712 7540 8736
rect 7668 8712 7720 8736
rect 4929 8672 4981 8712
rect 5140 8672 5177 8712
rect 5177 8672 5192 8712
rect 5351 8672 5383 8712
rect 5383 8672 5403 8712
rect 5562 8672 5589 8712
rect 5589 8672 5614 8712
rect 5773 8672 5795 8712
rect 5795 8672 5825 8712
rect 7488 8684 7506 8712
rect 7506 8684 7540 8712
rect 7668 8684 7669 8712
rect 7669 8684 7720 8712
rect 3864 8529 3899 8564
rect 3899 8529 3916 8564
rect 4044 8529 4048 8564
rect 4048 8529 4096 8564
rect 4224 8529 4255 8564
rect 4255 8529 4276 8564
rect 3864 8512 3916 8529
rect 4044 8512 4096 8529
rect 4224 8512 4276 8529
rect 2654 8351 2706 8354
rect 2834 8351 2886 8354
rect 2654 8305 2706 8351
rect 2834 8305 2886 8351
rect 2654 8302 2706 8305
rect 2834 8302 2886 8305
rect 6275 8437 6294 8489
rect 6294 8437 6327 8489
rect 6558 8488 6610 8496
rect 6769 8488 6821 8496
rect 6558 8444 6568 8488
rect 6568 8444 6610 8488
rect 6769 8444 6803 8488
rect 6803 8444 6821 8488
rect 6981 8444 7033 8496
rect 7192 8444 7244 8496
rect 9591 9427 9643 9479
rect 9372 9247 9424 9264
rect 9372 9212 9383 9247
rect 9383 9212 9424 9247
rect 12665 9443 12717 9495
rect 11532 9212 11584 9264
rect 17083 9552 17135 9604
rect 18193 9598 18245 9650
rect 21432 9695 21484 9720
rect 21612 9695 21664 9720
rect 21432 9668 21484 9695
rect 21612 9668 21664 9695
rect 14536 9471 14588 9488
rect 14748 9471 14800 9488
rect 14536 9436 14568 9471
rect 14568 9436 14588 9471
rect 14748 9436 14794 9471
rect 14794 9436 14800 9471
rect 18193 9380 18245 9432
rect 19897 9436 19949 9488
rect 20108 9471 20160 9488
rect 20108 9436 20110 9471
rect 20110 9436 20160 9471
rect 20319 9436 20371 9488
rect 18540 9288 18581 9325
rect 18581 9288 18592 9325
rect 18751 9288 18787 9325
rect 18787 9288 18803 9325
rect 18962 9288 18993 9325
rect 18993 9288 19014 9325
rect 19173 9288 19199 9325
rect 19199 9288 19225 9325
rect 19384 9288 19436 9325
rect 18540 9273 18592 9288
rect 18751 9273 18803 9288
rect 18962 9273 19014 9288
rect 19173 9273 19225 9288
rect 19384 9273 19436 9288
rect 20670 9247 20722 9250
rect 20850 9247 20902 9250
rect 20670 9201 20683 9247
rect 20683 9201 20722 9247
rect 20850 9201 20889 9247
rect 20889 9201 20902 9247
rect 20670 9198 20722 9201
rect 20850 9198 20902 9201
rect 21432 9247 21484 9257
rect 21612 9247 21664 9257
rect 21432 9205 21484 9247
rect 21612 9205 21664 9247
rect 9850 8974 9902 9026
rect 10030 8974 10082 9026
rect 13387 8974 13439 9026
rect 13598 8974 13650 9026
rect 13810 9023 13862 9026
rect 13810 8977 13833 9023
rect 13833 8977 13862 9023
rect 13810 8974 13862 8977
rect 14021 8974 14073 9026
rect 14431 9023 14483 9026
rect 14642 9023 14694 9026
rect 14853 9023 14905 9026
rect 14431 8977 14455 9023
rect 14455 8977 14483 9023
rect 14642 8977 14681 9023
rect 14681 8977 14694 9023
rect 14853 8977 14861 9023
rect 14861 8977 14905 9023
rect 14431 8974 14483 8977
rect 14642 8974 14694 8977
rect 14853 8974 14905 8977
rect 18435 8974 18487 9026
rect 18645 8974 18697 9026
rect 18856 8974 18908 9026
rect 19068 8974 19120 9026
rect 19279 8974 19331 9026
rect 19489 8974 19541 9026
rect 19943 8974 19995 9026
rect 20154 9023 20206 9026
rect 20365 9023 20417 9026
rect 21913 9023 21965 9026
rect 22124 9023 22176 9026
rect 22335 9023 22387 9026
rect 22545 9023 22597 9026
rect 22756 9023 22808 9026
rect 22968 9023 23020 9026
rect 23179 9023 23231 9026
rect 20154 8977 20168 9023
rect 20168 8977 20206 9023
rect 20365 8977 20374 9023
rect 20374 8977 20417 9023
rect 21913 8977 21965 9023
rect 22124 8977 22176 9023
rect 22335 8977 22387 9023
rect 22545 8977 22597 9023
rect 22756 8977 22808 9023
rect 22968 8977 23020 9023
rect 23179 8977 23231 9023
rect 20154 8974 20206 8977
rect 20365 8974 20417 8977
rect 9372 8753 9383 8788
rect 9383 8753 9424 8788
rect 9372 8736 9424 8753
rect 9591 8521 9643 8573
rect 9591 8335 9643 8387
rect 21913 8974 21965 8977
rect 22124 8974 22176 8977
rect 22335 8974 22387 8977
rect 22545 8974 22597 8977
rect 22756 8974 22808 8977
rect 22968 8974 23020 8977
rect 23179 8974 23231 8977
rect 23389 8974 23441 9026
rect 23600 8974 23652 9026
rect 23811 8974 23863 9026
rect 11532 8736 11584 8788
rect 20670 8799 20722 8802
rect 20850 8799 20902 8802
rect 12665 8505 12717 8557
rect 20670 8753 20683 8799
rect 20683 8753 20722 8799
rect 20850 8753 20889 8799
rect 20889 8753 20902 8799
rect 18540 8712 18592 8727
rect 18751 8712 18803 8727
rect 18962 8712 19014 8727
rect 19173 8712 19225 8727
rect 19384 8712 19436 8727
rect 18540 8675 18581 8712
rect 18581 8675 18592 8712
rect 18751 8675 18787 8712
rect 18787 8675 18803 8712
rect 18962 8675 18993 8712
rect 18993 8675 19014 8712
rect 19173 8675 19199 8712
rect 19199 8675 19225 8712
rect 19384 8675 19436 8712
rect 20670 8750 20722 8753
rect 20850 8750 20902 8753
rect 14536 8529 14568 8564
rect 14568 8529 14588 8564
rect 14748 8529 14794 8564
rect 14794 8529 14800 8564
rect 18193 8568 18245 8620
rect 14536 8512 14588 8529
rect 14748 8512 14800 8529
rect 17461 8396 17513 8448
rect 19897 8512 19949 8564
rect 20108 8529 20110 8564
rect 20110 8529 20160 8564
rect 20108 8512 20160 8529
rect 20319 8512 20371 8564
rect 18193 8350 18245 8402
rect 21432 8753 21484 8795
rect 21612 8753 21664 8795
rect 21432 8743 21484 8753
rect 21612 8743 21664 8753
rect 4929 8218 4981 8264
rect 5140 8218 5177 8264
rect 5177 8218 5192 8264
rect 5351 8218 5383 8264
rect 5383 8218 5403 8264
rect 5562 8218 5589 8264
rect 5589 8218 5614 8264
rect 5773 8218 5795 8264
rect 5795 8218 5825 8264
rect 7488 8218 7506 8262
rect 7506 8218 7540 8262
rect 7668 8218 7669 8262
rect 7669 8218 7720 8262
rect 18540 8218 18581 8264
rect 18581 8218 18592 8264
rect 18751 8218 18787 8264
rect 18787 8218 18803 8264
rect 18962 8218 18993 8264
rect 18993 8218 19014 8264
rect 19173 8218 19199 8264
rect 19199 8218 19225 8264
rect 19384 8218 19436 8264
rect 21432 8305 21484 8332
rect 21612 8305 21664 8332
rect 21432 8280 21484 8305
rect 21612 8280 21664 8305
rect 4929 8212 4981 8218
rect 5140 8212 5192 8218
rect 5351 8212 5403 8218
rect 5562 8212 5614 8218
rect 5773 8212 5825 8218
rect 7488 8210 7540 8218
rect 7668 8210 7720 8218
rect 451 8074 503 8126
rect 662 8074 714 8126
rect 873 8074 925 8126
rect 1083 8074 1135 8126
rect 1294 8074 1346 8126
rect 1506 8074 1558 8126
rect 1717 8074 1769 8126
rect 1927 8074 1979 8126
rect 2138 8074 2190 8126
rect 2349 8074 2401 8126
rect 18540 8212 18592 8218
rect 18751 8212 18803 8218
rect 18962 8212 19014 8218
rect 19173 8212 19225 8218
rect 19384 8212 19436 8218
rect 4352 8074 4404 8126
rect 4532 8123 4584 8126
rect 4532 8077 4559 8123
rect 4559 8077 4584 8123
rect 4532 8074 4584 8077
rect 19735 8123 19787 8126
rect 19735 8077 19757 8123
rect 19757 8077 19787 8123
rect 19735 8074 19787 8077
rect 19915 8074 19967 8126
rect 4929 7982 4981 7988
rect 5140 7982 5192 7988
rect 5351 7982 5403 7988
rect 5562 7982 5614 7988
rect 5773 7982 5825 7988
rect 7488 7982 7540 7990
rect 7668 7982 7720 7990
rect 21913 8074 21965 8126
rect 22124 8074 22176 8126
rect 22335 8074 22387 8126
rect 22545 8074 22597 8126
rect 22756 8074 22808 8126
rect 22968 8074 23020 8126
rect 23179 8074 23231 8126
rect 23389 8074 23441 8126
rect 23600 8074 23652 8126
rect 23811 8074 23863 8126
rect 18540 7982 18592 7988
rect 18751 7982 18803 7988
rect 18962 7982 19014 7988
rect 19173 7982 19225 7988
rect 19384 7982 19436 7988
rect 2654 7895 2706 7898
rect 2834 7895 2886 7898
rect 4929 7936 4981 7982
rect 5140 7936 5177 7982
rect 5177 7936 5192 7982
rect 5351 7936 5383 7982
rect 5383 7936 5403 7982
rect 5562 7936 5589 7982
rect 5589 7936 5614 7982
rect 5773 7936 5795 7982
rect 5795 7936 5825 7982
rect 7488 7938 7506 7982
rect 7506 7938 7540 7982
rect 7668 7938 7669 7982
rect 7669 7938 7720 7982
rect 2654 7849 2706 7895
rect 2834 7849 2886 7895
rect 2654 7846 2706 7849
rect 2834 7846 2886 7849
rect 2654 7447 2706 7450
rect 2834 7447 2886 7450
rect 2654 7401 2706 7447
rect 2834 7401 2886 7447
rect 2654 7398 2706 7401
rect 2834 7398 2886 7401
rect 3864 7671 3916 7688
rect 4044 7671 4096 7688
rect 4224 7671 4276 7688
rect 3864 7636 3899 7671
rect 3899 7636 3916 7671
rect 4044 7636 4048 7671
rect 4048 7636 4096 7671
rect 4224 7636 4255 7671
rect 4255 7636 4276 7671
rect 6275 7711 6294 7763
rect 6294 7711 6327 7763
rect 18540 7936 18581 7982
rect 18581 7936 18592 7982
rect 18751 7936 18787 7982
rect 18787 7936 18803 7982
rect 18962 7936 18993 7982
rect 18993 7936 19014 7982
rect 19173 7936 19199 7982
rect 19199 7936 19225 7982
rect 19384 7936 19436 7982
rect 9591 7813 9643 7865
rect 6558 7712 6568 7756
rect 6568 7712 6610 7756
rect 6769 7712 6803 7756
rect 6803 7712 6821 7756
rect 6558 7704 6610 7712
rect 6769 7704 6821 7712
rect 6981 7704 7033 7756
rect 7192 7704 7244 7756
rect 4929 7488 4981 7528
rect 5140 7488 5177 7528
rect 5177 7488 5192 7528
rect 5351 7488 5383 7528
rect 5383 7488 5403 7528
rect 5562 7488 5589 7528
rect 5589 7488 5614 7528
rect 5773 7488 5795 7528
rect 5795 7488 5825 7528
rect 7488 7488 7506 7516
rect 7506 7488 7540 7516
rect 7668 7488 7669 7516
rect 7669 7488 7720 7516
rect 4929 7476 4981 7488
rect 5140 7476 5192 7488
rect 5351 7476 5403 7488
rect 5562 7476 5614 7488
rect 5773 7476 5825 7488
rect 3416 7401 3430 7442
rect 3430 7401 3468 7442
rect 3596 7401 3636 7442
rect 3636 7401 3648 7442
rect 7488 7464 7540 7488
rect 7668 7464 7720 7488
rect 3416 7390 3468 7401
rect 3596 7390 3648 7401
rect 451 7174 503 7226
rect 662 7174 714 7226
rect 873 7174 925 7226
rect 1083 7223 1135 7226
rect 1294 7223 1346 7226
rect 1506 7223 1558 7226
rect 1717 7223 1769 7226
rect 1927 7223 1979 7226
rect 2138 7223 2190 7226
rect 2349 7223 2401 7226
rect 3881 7223 3933 7226
rect 4092 7223 4144 7226
rect 1083 7177 1135 7223
rect 1294 7177 1346 7223
rect 1506 7177 1558 7223
rect 1717 7177 1769 7223
rect 1927 7177 1979 7223
rect 2138 7177 2190 7223
rect 2349 7177 2401 7223
rect 3881 7177 3899 7223
rect 3899 7177 3933 7223
rect 4092 7177 4105 7223
rect 4105 7177 4144 7223
rect 1083 7174 1135 7177
rect 1294 7174 1346 7177
rect 1506 7174 1558 7177
rect 1717 7174 1769 7177
rect 1927 7174 1979 7177
rect 2138 7174 2190 7177
rect 2349 7174 2401 7177
rect 3881 7174 3933 7177
rect 4092 7174 4144 7177
rect 4304 7174 4356 7226
rect 4515 7174 4567 7226
rect 4817 7174 4869 7226
rect 5027 7174 5079 7226
rect 5238 7174 5290 7226
rect 5450 7174 5502 7226
rect 5661 7174 5713 7226
rect 5871 7174 5923 7226
rect 7927 7223 7979 7226
rect 7927 7177 7979 7223
rect 7927 7174 7979 7177
rect 8138 7174 8190 7226
rect 8349 7174 8401 7226
rect 8649 7223 8701 7226
rect 8829 7223 8881 7226
rect 8649 7177 8659 7223
rect 8659 7177 8701 7223
rect 8829 7177 8863 7223
rect 8863 7177 8881 7223
rect 8649 7174 8701 7177
rect 8829 7174 8881 7177
rect 2654 6999 2706 7002
rect 2834 6999 2886 7002
rect 2654 6953 2706 6999
rect 2834 6953 2886 6999
rect 2654 6950 2706 6953
rect 2834 6950 2886 6953
rect 3416 6999 3468 7010
rect 3596 6999 3648 7010
rect 3416 6958 3430 6999
rect 3430 6958 3468 6999
rect 3596 6958 3636 6999
rect 3636 6958 3648 6999
rect 4929 6912 4981 6924
rect 5140 6912 5192 6924
rect 5351 6912 5403 6924
rect 5562 6912 5614 6924
rect 5773 6912 5825 6924
rect 7488 6912 7540 6936
rect 7668 6912 7720 6936
rect 4929 6872 4981 6912
rect 5140 6872 5177 6912
rect 5177 6872 5192 6912
rect 5351 6872 5383 6912
rect 5383 6872 5403 6912
rect 5562 6872 5589 6912
rect 5589 6872 5614 6912
rect 5773 6872 5795 6912
rect 5795 6872 5825 6912
rect 7488 6884 7506 6912
rect 7506 6884 7540 6912
rect 7668 6884 7669 6912
rect 7669 6884 7720 6912
rect 3864 6729 3899 6764
rect 3899 6729 3916 6764
rect 4044 6729 4048 6764
rect 4048 6729 4096 6764
rect 4224 6729 4255 6764
rect 4255 6729 4276 6764
rect 3864 6712 3916 6729
rect 4044 6712 4096 6729
rect 4224 6712 4276 6729
rect 2654 6551 2706 6554
rect 2834 6551 2886 6554
rect 2654 6505 2706 6551
rect 2834 6505 2886 6551
rect 2654 6502 2706 6505
rect 2834 6502 2886 6505
rect 6275 6637 6294 6689
rect 6294 6637 6327 6689
rect 6558 6688 6610 6696
rect 6769 6688 6821 6696
rect 6558 6644 6568 6688
rect 6568 6644 6610 6688
rect 6769 6644 6803 6688
rect 6803 6644 6821 6688
rect 6981 6644 7033 6696
rect 7192 6644 7244 6696
rect 9591 7627 9643 7679
rect 9372 7447 9424 7464
rect 9372 7412 9383 7447
rect 9383 7412 9424 7447
rect 12665 7643 12717 7695
rect 11532 7412 11584 7464
rect 17838 7752 17890 7804
rect 18193 7798 18245 7850
rect 21432 7895 21484 7920
rect 21612 7895 21664 7920
rect 21432 7868 21484 7895
rect 21612 7868 21664 7895
rect 14536 7671 14588 7688
rect 14748 7671 14800 7688
rect 14536 7636 14568 7671
rect 14568 7636 14588 7671
rect 14748 7636 14794 7671
rect 14794 7636 14800 7671
rect 18193 7580 18245 7632
rect 19897 7636 19949 7688
rect 20108 7671 20160 7688
rect 20108 7636 20110 7671
rect 20110 7636 20160 7671
rect 20319 7636 20371 7688
rect 18540 7488 18581 7525
rect 18581 7488 18592 7525
rect 18751 7488 18787 7525
rect 18787 7488 18803 7525
rect 18962 7488 18993 7525
rect 18993 7488 19014 7525
rect 19173 7488 19199 7525
rect 19199 7488 19225 7525
rect 19384 7488 19436 7525
rect 18540 7473 18592 7488
rect 18751 7473 18803 7488
rect 18962 7473 19014 7488
rect 19173 7473 19225 7488
rect 19384 7473 19436 7488
rect 20670 7447 20722 7450
rect 20850 7447 20902 7450
rect 20670 7401 20683 7447
rect 20683 7401 20722 7447
rect 20850 7401 20889 7447
rect 20889 7401 20902 7447
rect 20670 7398 20722 7401
rect 20850 7398 20902 7401
rect 21432 7447 21484 7457
rect 21612 7447 21664 7457
rect 21432 7405 21484 7447
rect 21612 7405 21664 7447
rect 9850 7174 9902 7226
rect 10030 7174 10082 7226
rect 13387 7174 13439 7226
rect 13598 7174 13650 7226
rect 13810 7223 13862 7226
rect 13810 7177 13833 7223
rect 13833 7177 13862 7223
rect 13810 7174 13862 7177
rect 14021 7174 14073 7226
rect 14431 7223 14483 7226
rect 14642 7223 14694 7226
rect 14853 7223 14905 7226
rect 14431 7177 14455 7223
rect 14455 7177 14483 7223
rect 14642 7177 14681 7223
rect 14681 7177 14694 7223
rect 14853 7177 14861 7223
rect 14861 7177 14905 7223
rect 14431 7174 14483 7177
rect 14642 7174 14694 7177
rect 14853 7174 14905 7177
rect 18435 7174 18487 7226
rect 18645 7174 18697 7226
rect 18856 7174 18908 7226
rect 19068 7174 19120 7226
rect 19279 7174 19331 7226
rect 19489 7174 19541 7226
rect 19943 7174 19995 7226
rect 20154 7223 20206 7226
rect 20365 7223 20417 7226
rect 21913 7223 21965 7226
rect 22124 7223 22176 7226
rect 22335 7223 22387 7226
rect 22545 7223 22597 7226
rect 22756 7223 22808 7226
rect 22968 7223 23020 7226
rect 23179 7223 23231 7226
rect 20154 7177 20168 7223
rect 20168 7177 20206 7223
rect 20365 7177 20374 7223
rect 20374 7177 20417 7223
rect 21913 7177 21965 7223
rect 22124 7177 22176 7223
rect 22335 7177 22387 7223
rect 22545 7177 22597 7223
rect 22756 7177 22808 7223
rect 22968 7177 23020 7223
rect 23179 7177 23231 7223
rect 20154 7174 20206 7177
rect 20365 7174 20417 7177
rect 9372 6953 9383 6988
rect 9383 6953 9424 6988
rect 9372 6936 9424 6953
rect 9591 6721 9643 6773
rect 9591 6535 9643 6587
rect 21913 7174 21965 7177
rect 22124 7174 22176 7177
rect 22335 7174 22387 7177
rect 22545 7174 22597 7177
rect 22756 7174 22808 7177
rect 22968 7174 23020 7177
rect 23179 7174 23231 7177
rect 23389 7174 23441 7226
rect 23600 7174 23652 7226
rect 23811 7174 23863 7226
rect 11532 6936 11584 6988
rect 20670 6999 20722 7002
rect 20850 6999 20902 7002
rect 13042 6705 13094 6757
rect 20670 6953 20683 6999
rect 20683 6953 20722 6999
rect 20850 6953 20889 6999
rect 20889 6953 20902 6999
rect 18540 6912 18592 6927
rect 18751 6912 18803 6927
rect 18962 6912 19014 6927
rect 19173 6912 19225 6927
rect 19384 6912 19436 6927
rect 18540 6875 18581 6912
rect 18581 6875 18592 6912
rect 18751 6875 18787 6912
rect 18787 6875 18803 6912
rect 18962 6875 18993 6912
rect 18993 6875 19014 6912
rect 19173 6875 19199 6912
rect 19199 6875 19225 6912
rect 19384 6875 19436 6912
rect 20670 6950 20722 6953
rect 20850 6950 20902 6953
rect 14536 6729 14568 6764
rect 14568 6729 14588 6764
rect 14748 6729 14794 6764
rect 14794 6729 14800 6764
rect 18193 6768 18245 6820
rect 14536 6712 14588 6729
rect 14748 6712 14800 6729
rect 15194 6610 15201 6648
rect 15201 6610 15246 6648
rect 15194 6596 15246 6610
rect 19897 6712 19949 6764
rect 20108 6729 20110 6764
rect 20110 6729 20160 6764
rect 20108 6712 20160 6729
rect 20319 6712 20371 6764
rect 18193 6550 18245 6602
rect 21432 6953 21484 6995
rect 21612 6953 21664 6995
rect 21432 6943 21484 6953
rect 21612 6943 21664 6953
rect 4929 6418 4981 6464
rect 5140 6418 5177 6464
rect 5177 6418 5192 6464
rect 5351 6418 5383 6464
rect 5383 6418 5403 6464
rect 5562 6418 5589 6464
rect 5589 6418 5614 6464
rect 5773 6418 5795 6464
rect 5795 6418 5825 6464
rect 7488 6418 7506 6462
rect 7506 6418 7540 6462
rect 7668 6418 7669 6462
rect 7669 6418 7720 6462
rect 18540 6418 18581 6464
rect 18581 6418 18592 6464
rect 18751 6418 18787 6464
rect 18787 6418 18803 6464
rect 18962 6418 18993 6464
rect 18993 6418 19014 6464
rect 19173 6418 19199 6464
rect 19199 6418 19225 6464
rect 19384 6418 19436 6464
rect 21432 6505 21484 6532
rect 21612 6505 21664 6532
rect 21432 6480 21484 6505
rect 21612 6480 21664 6505
rect 4929 6412 4981 6418
rect 5140 6412 5192 6418
rect 5351 6412 5403 6418
rect 5562 6412 5614 6418
rect 5773 6412 5825 6418
rect 7488 6410 7540 6418
rect 7668 6410 7720 6418
rect 451 6274 503 6326
rect 662 6274 714 6326
rect 873 6274 925 6326
rect 1083 6274 1135 6326
rect 1294 6274 1346 6326
rect 1506 6274 1558 6326
rect 1717 6274 1769 6326
rect 1927 6274 1979 6326
rect 2138 6274 2190 6326
rect 2349 6274 2401 6326
rect 18540 6412 18592 6418
rect 18751 6412 18803 6418
rect 18962 6412 19014 6418
rect 19173 6412 19225 6418
rect 19384 6412 19436 6418
rect 4352 6274 4404 6326
rect 4532 6323 4584 6326
rect 4532 6277 4559 6323
rect 4559 6277 4584 6323
rect 4532 6274 4584 6277
rect 19735 6323 19787 6326
rect 19735 6277 19757 6323
rect 19757 6277 19787 6323
rect 19735 6274 19787 6277
rect 19915 6274 19967 6326
rect 4929 6182 4981 6188
rect 5140 6182 5192 6188
rect 5351 6182 5403 6188
rect 5562 6182 5614 6188
rect 5773 6182 5825 6188
rect 7488 6182 7540 6190
rect 7668 6182 7720 6190
rect 21913 6274 21965 6326
rect 22124 6274 22176 6326
rect 22335 6274 22387 6326
rect 22545 6274 22597 6326
rect 22756 6274 22808 6326
rect 22968 6274 23020 6326
rect 23179 6274 23231 6326
rect 23389 6274 23441 6326
rect 23600 6274 23652 6326
rect 23811 6274 23863 6326
rect 18540 6182 18592 6188
rect 18751 6182 18803 6188
rect 18962 6182 19014 6188
rect 19173 6182 19225 6188
rect 19384 6182 19436 6188
rect 2654 6095 2706 6098
rect 2834 6095 2886 6098
rect 4929 6136 4981 6182
rect 5140 6136 5177 6182
rect 5177 6136 5192 6182
rect 5351 6136 5383 6182
rect 5383 6136 5403 6182
rect 5562 6136 5589 6182
rect 5589 6136 5614 6182
rect 5773 6136 5795 6182
rect 5795 6136 5825 6182
rect 7488 6138 7506 6182
rect 7506 6138 7540 6182
rect 7668 6138 7669 6182
rect 7669 6138 7720 6182
rect 2654 6049 2706 6095
rect 2834 6049 2886 6095
rect 2654 6046 2706 6049
rect 2834 6046 2886 6049
rect 2654 5647 2706 5650
rect 2834 5647 2886 5650
rect 2654 5601 2706 5647
rect 2834 5601 2886 5647
rect 2654 5598 2706 5601
rect 2834 5598 2886 5601
rect 3864 5871 3916 5888
rect 4044 5871 4096 5888
rect 4224 5871 4276 5888
rect 3864 5836 3899 5871
rect 3899 5836 3916 5871
rect 4044 5836 4048 5871
rect 4048 5836 4096 5871
rect 4224 5836 4255 5871
rect 4255 5836 4276 5871
rect 6275 5911 6294 5963
rect 6294 5911 6327 5963
rect 18540 6136 18581 6182
rect 18581 6136 18592 6182
rect 18751 6136 18787 6182
rect 18787 6136 18803 6182
rect 18962 6136 18993 6182
rect 18993 6136 19014 6182
rect 19173 6136 19199 6182
rect 19199 6136 19225 6182
rect 19384 6136 19436 6182
rect 9591 6013 9643 6065
rect 6558 5912 6568 5956
rect 6568 5912 6610 5956
rect 6769 5912 6803 5956
rect 6803 5912 6821 5956
rect 6558 5904 6610 5912
rect 6769 5904 6821 5912
rect 6981 5904 7033 5956
rect 7192 5904 7244 5956
rect 4929 5688 4981 5728
rect 5140 5688 5177 5728
rect 5177 5688 5192 5728
rect 5351 5688 5383 5728
rect 5383 5688 5403 5728
rect 5562 5688 5589 5728
rect 5589 5688 5614 5728
rect 5773 5688 5795 5728
rect 5795 5688 5825 5728
rect 7488 5688 7506 5716
rect 7506 5688 7540 5716
rect 7668 5688 7669 5716
rect 7669 5688 7720 5716
rect 4929 5676 4981 5688
rect 5140 5676 5192 5688
rect 5351 5676 5403 5688
rect 5562 5676 5614 5688
rect 5773 5676 5825 5688
rect 3416 5601 3430 5642
rect 3430 5601 3468 5642
rect 3596 5601 3636 5642
rect 3636 5601 3648 5642
rect 7488 5664 7540 5688
rect 7668 5664 7720 5688
rect 3416 5590 3468 5601
rect 3596 5590 3648 5601
rect 451 5374 503 5426
rect 662 5374 714 5426
rect 873 5374 925 5426
rect 1083 5423 1135 5426
rect 1294 5423 1346 5426
rect 1506 5423 1558 5426
rect 1717 5423 1769 5426
rect 1927 5423 1979 5426
rect 2138 5423 2190 5426
rect 2349 5423 2401 5426
rect 3881 5423 3933 5426
rect 4092 5423 4144 5426
rect 1083 5377 1135 5423
rect 1294 5377 1346 5423
rect 1506 5377 1558 5423
rect 1717 5377 1769 5423
rect 1927 5377 1979 5423
rect 2138 5377 2190 5423
rect 2349 5377 2401 5423
rect 3881 5377 3899 5423
rect 3899 5377 3933 5423
rect 4092 5377 4105 5423
rect 4105 5377 4144 5423
rect 1083 5374 1135 5377
rect 1294 5374 1346 5377
rect 1506 5374 1558 5377
rect 1717 5374 1769 5377
rect 1927 5374 1979 5377
rect 2138 5374 2190 5377
rect 2349 5374 2401 5377
rect 3881 5374 3933 5377
rect 4092 5374 4144 5377
rect 4304 5374 4356 5426
rect 4515 5374 4567 5426
rect 4817 5374 4869 5426
rect 5027 5374 5079 5426
rect 5238 5374 5290 5426
rect 5450 5374 5502 5426
rect 5661 5374 5713 5426
rect 5871 5374 5923 5426
rect 7927 5423 7979 5426
rect 7927 5377 7979 5423
rect 7927 5374 7979 5377
rect 8138 5374 8190 5426
rect 8349 5374 8401 5426
rect 8649 5423 8701 5426
rect 8829 5423 8881 5426
rect 8649 5377 8659 5423
rect 8659 5377 8701 5423
rect 8829 5377 8863 5423
rect 8863 5377 8881 5423
rect 8649 5374 8701 5377
rect 8829 5374 8881 5377
rect 2654 5199 2706 5202
rect 2834 5199 2886 5202
rect 2654 5153 2706 5199
rect 2834 5153 2886 5199
rect 2654 5150 2706 5153
rect 2834 5150 2886 5153
rect 3416 5199 3468 5210
rect 3596 5199 3648 5210
rect 3416 5158 3430 5199
rect 3430 5158 3468 5199
rect 3596 5158 3636 5199
rect 3636 5158 3648 5199
rect 4929 5112 4981 5124
rect 5140 5112 5192 5124
rect 5351 5112 5403 5124
rect 5562 5112 5614 5124
rect 5773 5112 5825 5124
rect 7488 5112 7540 5136
rect 7668 5112 7720 5136
rect 4929 5072 4981 5112
rect 5140 5072 5177 5112
rect 5177 5072 5192 5112
rect 5351 5072 5383 5112
rect 5383 5072 5403 5112
rect 5562 5072 5589 5112
rect 5589 5072 5614 5112
rect 5773 5072 5795 5112
rect 5795 5072 5825 5112
rect 7488 5084 7506 5112
rect 7506 5084 7540 5112
rect 7668 5084 7669 5112
rect 7669 5084 7720 5112
rect 3864 4929 3899 4964
rect 3899 4929 3916 4964
rect 4044 4929 4048 4964
rect 4048 4929 4096 4964
rect 4224 4929 4255 4964
rect 4255 4929 4276 4964
rect 3864 4912 3916 4929
rect 4044 4912 4096 4929
rect 4224 4912 4276 4929
rect 2654 4751 2706 4754
rect 2834 4751 2886 4754
rect 2654 4705 2706 4751
rect 2834 4705 2886 4751
rect 2654 4702 2706 4705
rect 2834 4702 2886 4705
rect 6275 4837 6294 4889
rect 6294 4837 6327 4889
rect 6558 4888 6610 4896
rect 6769 4888 6821 4896
rect 6558 4844 6568 4888
rect 6568 4844 6610 4888
rect 6769 4844 6803 4888
rect 6803 4844 6821 4888
rect 6981 4844 7033 4896
rect 7192 4844 7244 4896
rect 9591 5827 9643 5879
rect 9372 5647 9424 5664
rect 9372 5612 9383 5647
rect 9383 5612 9424 5647
rect 13042 5843 13094 5895
rect 11532 5612 11584 5664
rect 15572 5952 15624 6004
rect 18193 5998 18245 6050
rect 21432 6095 21484 6120
rect 21612 6095 21664 6120
rect 21432 6068 21484 6095
rect 21612 6068 21664 6095
rect 14536 5871 14588 5888
rect 14748 5871 14800 5888
rect 14536 5836 14568 5871
rect 14568 5836 14588 5871
rect 14748 5836 14794 5871
rect 14794 5836 14800 5871
rect 18193 5780 18245 5832
rect 19897 5836 19949 5888
rect 20108 5871 20160 5888
rect 20108 5836 20110 5871
rect 20110 5836 20160 5871
rect 20319 5836 20371 5888
rect 18540 5688 18581 5725
rect 18581 5688 18592 5725
rect 18751 5688 18787 5725
rect 18787 5688 18803 5725
rect 18962 5688 18993 5725
rect 18993 5688 19014 5725
rect 19173 5688 19199 5725
rect 19199 5688 19225 5725
rect 19384 5688 19436 5725
rect 18540 5673 18592 5688
rect 18751 5673 18803 5688
rect 18962 5673 19014 5688
rect 19173 5673 19225 5688
rect 19384 5673 19436 5688
rect 20670 5647 20722 5650
rect 20850 5647 20902 5650
rect 20670 5601 20683 5647
rect 20683 5601 20722 5647
rect 20850 5601 20889 5647
rect 20889 5601 20902 5647
rect 20670 5598 20722 5601
rect 20850 5598 20902 5601
rect 21432 5647 21484 5657
rect 21612 5647 21664 5657
rect 21432 5605 21484 5647
rect 21612 5605 21664 5647
rect 9850 5374 9902 5426
rect 10030 5374 10082 5426
rect 13387 5374 13439 5426
rect 13598 5374 13650 5426
rect 13810 5423 13862 5426
rect 13810 5377 13833 5423
rect 13833 5377 13862 5423
rect 13810 5374 13862 5377
rect 14021 5374 14073 5426
rect 14431 5423 14483 5426
rect 14642 5423 14694 5426
rect 14853 5423 14905 5426
rect 14431 5377 14455 5423
rect 14455 5377 14483 5423
rect 14642 5377 14681 5423
rect 14681 5377 14694 5423
rect 14853 5377 14861 5423
rect 14861 5377 14905 5423
rect 14431 5374 14483 5377
rect 14642 5374 14694 5377
rect 14853 5374 14905 5377
rect 18435 5374 18487 5426
rect 18645 5374 18697 5426
rect 18856 5374 18908 5426
rect 19068 5374 19120 5426
rect 19279 5374 19331 5426
rect 19489 5374 19541 5426
rect 19943 5374 19995 5426
rect 20154 5423 20206 5426
rect 20365 5423 20417 5426
rect 21913 5423 21965 5426
rect 22124 5423 22176 5426
rect 22335 5423 22387 5426
rect 22545 5423 22597 5426
rect 22756 5423 22808 5426
rect 22968 5423 23020 5426
rect 23179 5423 23231 5426
rect 20154 5377 20168 5423
rect 20168 5377 20206 5423
rect 20365 5377 20374 5423
rect 20374 5377 20417 5423
rect 21913 5377 21965 5423
rect 22124 5377 22176 5423
rect 22335 5377 22387 5423
rect 22545 5377 22597 5423
rect 22756 5377 22808 5423
rect 22968 5377 23020 5423
rect 23179 5377 23231 5423
rect 20154 5374 20206 5377
rect 20365 5374 20417 5377
rect 9372 5153 9383 5188
rect 9383 5153 9424 5188
rect 9372 5136 9424 5153
rect 9591 4921 9643 4973
rect 9591 4735 9643 4787
rect 21913 5374 21965 5377
rect 22124 5374 22176 5377
rect 22335 5374 22387 5377
rect 22545 5374 22597 5377
rect 22756 5374 22808 5377
rect 22968 5374 23020 5377
rect 23179 5374 23231 5377
rect 23389 5374 23441 5426
rect 23600 5374 23652 5426
rect 23811 5374 23863 5426
rect 11532 5136 11584 5188
rect 20670 5199 20722 5202
rect 20850 5199 20902 5202
rect 13042 4905 13094 4957
rect 20670 5153 20683 5199
rect 20683 5153 20722 5199
rect 20850 5153 20889 5199
rect 20889 5153 20902 5199
rect 18540 5112 18592 5127
rect 18751 5112 18803 5127
rect 18962 5112 19014 5127
rect 19173 5112 19225 5127
rect 19384 5112 19436 5127
rect 18540 5075 18581 5112
rect 18581 5075 18592 5112
rect 18751 5075 18787 5112
rect 18787 5075 18803 5112
rect 18962 5075 18993 5112
rect 18993 5075 19014 5112
rect 19173 5075 19199 5112
rect 19199 5075 19225 5112
rect 19384 5075 19436 5112
rect 20670 5150 20722 5153
rect 20850 5150 20902 5153
rect 14536 4929 14568 4964
rect 14568 4929 14588 4964
rect 14748 4929 14794 4964
rect 14794 4929 14800 4964
rect 18193 4968 18245 5020
rect 14536 4912 14588 4929
rect 14748 4912 14800 4929
rect 15950 4796 16002 4848
rect 19897 4912 19949 4964
rect 20108 4929 20110 4964
rect 20110 4929 20160 4964
rect 20108 4912 20160 4929
rect 20319 4912 20371 4964
rect 18193 4750 18245 4802
rect 21432 5153 21484 5195
rect 21612 5153 21664 5195
rect 21432 5143 21484 5153
rect 21612 5143 21664 5153
rect 4929 4618 4981 4664
rect 5140 4618 5177 4664
rect 5177 4618 5192 4664
rect 5351 4618 5383 4664
rect 5383 4618 5403 4664
rect 5562 4618 5589 4664
rect 5589 4618 5614 4664
rect 5773 4618 5795 4664
rect 5795 4618 5825 4664
rect 7488 4618 7506 4662
rect 7506 4618 7540 4662
rect 7668 4618 7669 4662
rect 7669 4618 7720 4662
rect 18540 4618 18581 4664
rect 18581 4618 18592 4664
rect 18751 4618 18787 4664
rect 18787 4618 18803 4664
rect 18962 4618 18993 4664
rect 18993 4618 19014 4664
rect 19173 4618 19199 4664
rect 19199 4618 19225 4664
rect 19384 4618 19436 4664
rect 21432 4705 21484 4732
rect 21612 4705 21664 4732
rect 21432 4680 21484 4705
rect 21612 4680 21664 4705
rect 4929 4612 4981 4618
rect 5140 4612 5192 4618
rect 5351 4612 5403 4618
rect 5562 4612 5614 4618
rect 5773 4612 5825 4618
rect 7488 4610 7540 4618
rect 7668 4610 7720 4618
rect 451 4474 503 4526
rect 662 4474 714 4526
rect 873 4474 925 4526
rect 1083 4474 1135 4526
rect 1294 4474 1346 4526
rect 1506 4474 1558 4526
rect 1717 4474 1769 4526
rect 1927 4474 1979 4526
rect 2138 4474 2190 4526
rect 2349 4474 2401 4526
rect 18540 4612 18592 4618
rect 18751 4612 18803 4618
rect 18962 4612 19014 4618
rect 19173 4612 19225 4618
rect 19384 4612 19436 4618
rect 4352 4474 4404 4526
rect 4532 4523 4584 4526
rect 4532 4477 4559 4523
rect 4559 4477 4584 4523
rect 4532 4474 4584 4477
rect 19735 4523 19787 4526
rect 19735 4477 19757 4523
rect 19757 4477 19787 4523
rect 19735 4474 19787 4477
rect 19915 4474 19967 4526
rect 4929 4382 4981 4388
rect 5140 4382 5192 4388
rect 5351 4382 5403 4388
rect 5562 4382 5614 4388
rect 5773 4382 5825 4388
rect 7488 4382 7540 4390
rect 7668 4382 7720 4390
rect 21913 4474 21965 4526
rect 22124 4474 22176 4526
rect 22335 4474 22387 4526
rect 22545 4474 22597 4526
rect 22756 4474 22808 4526
rect 22968 4474 23020 4526
rect 23179 4474 23231 4526
rect 23389 4474 23441 4526
rect 23600 4474 23652 4526
rect 23811 4474 23863 4526
rect 18540 4382 18592 4388
rect 18751 4382 18803 4388
rect 18962 4382 19014 4388
rect 19173 4382 19225 4388
rect 19384 4382 19436 4388
rect 2654 4295 2706 4298
rect 2834 4295 2886 4298
rect 4929 4336 4981 4382
rect 5140 4336 5177 4382
rect 5177 4336 5192 4382
rect 5351 4336 5383 4382
rect 5383 4336 5403 4382
rect 5562 4336 5589 4382
rect 5589 4336 5614 4382
rect 5773 4336 5795 4382
rect 5795 4336 5825 4382
rect 7488 4338 7506 4382
rect 7506 4338 7540 4382
rect 7668 4338 7669 4382
rect 7669 4338 7720 4382
rect 2654 4249 2706 4295
rect 2834 4249 2886 4295
rect 2654 4246 2706 4249
rect 2834 4246 2886 4249
rect 2654 3847 2706 3850
rect 2834 3847 2886 3850
rect 2654 3801 2706 3847
rect 2834 3801 2886 3847
rect 2654 3798 2706 3801
rect 2834 3798 2886 3801
rect 3864 4071 3916 4088
rect 4044 4071 4096 4088
rect 4224 4071 4276 4088
rect 3864 4036 3899 4071
rect 3899 4036 3916 4071
rect 4044 4036 4048 4071
rect 4048 4036 4096 4071
rect 4224 4036 4255 4071
rect 4255 4036 4276 4071
rect 6275 4111 6294 4163
rect 6294 4111 6327 4163
rect 18540 4336 18581 4382
rect 18581 4336 18592 4382
rect 18751 4336 18787 4382
rect 18787 4336 18803 4382
rect 18962 4336 18993 4382
rect 18993 4336 19014 4382
rect 19173 4336 19199 4382
rect 19199 4336 19225 4382
rect 19384 4336 19436 4382
rect 9591 4213 9643 4265
rect 6558 4112 6568 4156
rect 6568 4112 6610 4156
rect 6769 4112 6803 4156
rect 6803 4112 6821 4156
rect 6558 4104 6610 4112
rect 6769 4104 6821 4112
rect 6981 4104 7033 4156
rect 7192 4104 7244 4156
rect 4929 3888 4981 3928
rect 5140 3888 5177 3928
rect 5177 3888 5192 3928
rect 5351 3888 5383 3928
rect 5383 3888 5403 3928
rect 5562 3888 5589 3928
rect 5589 3888 5614 3928
rect 5773 3888 5795 3928
rect 5795 3888 5825 3928
rect 7488 3888 7506 3916
rect 7506 3888 7540 3916
rect 7668 3888 7669 3916
rect 7669 3888 7720 3916
rect 4929 3876 4981 3888
rect 5140 3876 5192 3888
rect 5351 3876 5403 3888
rect 5562 3876 5614 3888
rect 5773 3876 5825 3888
rect 3416 3801 3430 3842
rect 3430 3801 3468 3842
rect 3596 3801 3636 3842
rect 3636 3801 3648 3842
rect 7488 3864 7540 3888
rect 7668 3864 7720 3888
rect 3416 3790 3468 3801
rect 3596 3790 3648 3801
rect 451 3574 503 3626
rect 662 3574 714 3626
rect 873 3574 925 3626
rect 1083 3623 1135 3626
rect 1294 3623 1346 3626
rect 1506 3623 1558 3626
rect 1717 3623 1769 3626
rect 1927 3623 1979 3626
rect 2138 3623 2190 3626
rect 2349 3623 2401 3626
rect 3881 3623 3933 3626
rect 4092 3623 4144 3626
rect 1083 3577 1135 3623
rect 1294 3577 1346 3623
rect 1506 3577 1558 3623
rect 1717 3577 1769 3623
rect 1927 3577 1979 3623
rect 2138 3577 2190 3623
rect 2349 3577 2401 3623
rect 3881 3577 3899 3623
rect 3899 3577 3933 3623
rect 4092 3577 4105 3623
rect 4105 3577 4144 3623
rect 1083 3574 1135 3577
rect 1294 3574 1346 3577
rect 1506 3574 1558 3577
rect 1717 3574 1769 3577
rect 1927 3574 1979 3577
rect 2138 3574 2190 3577
rect 2349 3574 2401 3577
rect 3881 3574 3933 3577
rect 4092 3574 4144 3577
rect 4304 3574 4356 3626
rect 4515 3574 4567 3626
rect 4817 3574 4869 3626
rect 5027 3574 5079 3626
rect 5238 3574 5290 3626
rect 5450 3574 5502 3626
rect 5661 3574 5713 3626
rect 5871 3574 5923 3626
rect 7927 3623 7979 3626
rect 7927 3577 7979 3623
rect 7927 3574 7979 3577
rect 8138 3574 8190 3626
rect 8349 3574 8401 3626
rect 8649 3623 8701 3626
rect 8829 3623 8881 3626
rect 8649 3577 8659 3623
rect 8659 3577 8701 3623
rect 8829 3577 8863 3623
rect 8863 3577 8881 3623
rect 8649 3574 8701 3577
rect 8829 3574 8881 3577
rect 2654 3399 2706 3402
rect 2834 3399 2886 3402
rect 2654 3353 2706 3399
rect 2834 3353 2886 3399
rect 2654 3350 2706 3353
rect 2834 3350 2886 3353
rect 3416 3399 3468 3410
rect 3596 3399 3648 3410
rect 3416 3358 3430 3399
rect 3430 3358 3468 3399
rect 3596 3358 3636 3399
rect 3636 3358 3648 3399
rect 4929 3312 4981 3324
rect 5140 3312 5192 3324
rect 5351 3312 5403 3324
rect 5562 3312 5614 3324
rect 5773 3312 5825 3324
rect 7488 3312 7540 3336
rect 7668 3312 7720 3336
rect 4929 3272 4981 3312
rect 5140 3272 5177 3312
rect 5177 3272 5192 3312
rect 5351 3272 5383 3312
rect 5383 3272 5403 3312
rect 5562 3272 5589 3312
rect 5589 3272 5614 3312
rect 5773 3272 5795 3312
rect 5795 3272 5825 3312
rect 7488 3284 7506 3312
rect 7506 3284 7540 3312
rect 7668 3284 7669 3312
rect 7669 3284 7720 3312
rect 3864 3129 3899 3164
rect 3899 3129 3916 3164
rect 4044 3129 4048 3164
rect 4048 3129 4096 3164
rect 4224 3129 4255 3164
rect 4255 3129 4276 3164
rect 3864 3112 3916 3129
rect 4044 3112 4096 3129
rect 4224 3112 4276 3129
rect 2654 2951 2706 2954
rect 2834 2951 2886 2954
rect 2654 2905 2706 2951
rect 2834 2905 2886 2951
rect 2654 2902 2706 2905
rect 2834 2902 2886 2905
rect 6275 3037 6294 3089
rect 6294 3037 6327 3089
rect 6558 3088 6610 3096
rect 6769 3088 6821 3096
rect 6558 3044 6568 3088
rect 6568 3044 6610 3088
rect 6769 3044 6803 3088
rect 6803 3044 6821 3088
rect 6981 3044 7033 3096
rect 7192 3044 7244 3096
rect 9591 4027 9643 4079
rect 9372 3847 9424 3864
rect 9372 3812 9383 3847
rect 9383 3812 9424 3847
rect 13042 4043 13094 4095
rect 11532 3812 11584 3864
rect 16328 4152 16380 4204
rect 18193 4198 18245 4250
rect 21432 4295 21484 4320
rect 21612 4295 21664 4320
rect 21432 4268 21484 4295
rect 21612 4268 21664 4295
rect 14536 4071 14588 4088
rect 14748 4071 14800 4088
rect 14536 4036 14568 4071
rect 14568 4036 14588 4071
rect 14748 4036 14794 4071
rect 14794 4036 14800 4071
rect 18193 3980 18245 4032
rect 19897 4036 19949 4088
rect 20108 4071 20160 4088
rect 20108 4036 20110 4071
rect 20110 4036 20160 4071
rect 20319 4036 20371 4088
rect 18540 3888 18581 3925
rect 18581 3888 18592 3925
rect 18751 3888 18787 3925
rect 18787 3888 18803 3925
rect 18962 3888 18993 3925
rect 18993 3888 19014 3925
rect 19173 3888 19199 3925
rect 19199 3888 19225 3925
rect 19384 3888 19436 3925
rect 18540 3873 18592 3888
rect 18751 3873 18803 3888
rect 18962 3873 19014 3888
rect 19173 3873 19225 3888
rect 19384 3873 19436 3888
rect 20670 3847 20722 3850
rect 20850 3847 20902 3850
rect 20670 3801 20683 3847
rect 20683 3801 20722 3847
rect 20850 3801 20889 3847
rect 20889 3801 20902 3847
rect 20670 3798 20722 3801
rect 20850 3798 20902 3801
rect 21432 3847 21484 3857
rect 21612 3847 21664 3857
rect 21432 3805 21484 3847
rect 21612 3805 21664 3847
rect 9850 3574 9902 3626
rect 10030 3574 10082 3626
rect 13387 3574 13439 3626
rect 13598 3574 13650 3626
rect 13810 3623 13862 3626
rect 13810 3577 13833 3623
rect 13833 3577 13862 3623
rect 13810 3574 13862 3577
rect 14021 3574 14073 3626
rect 14431 3623 14483 3626
rect 14642 3623 14694 3626
rect 14853 3623 14905 3626
rect 14431 3577 14455 3623
rect 14455 3577 14483 3623
rect 14642 3577 14681 3623
rect 14681 3577 14694 3623
rect 14853 3577 14861 3623
rect 14861 3577 14905 3623
rect 14431 3574 14483 3577
rect 14642 3574 14694 3577
rect 14853 3574 14905 3577
rect 18435 3574 18487 3626
rect 18645 3574 18697 3626
rect 18856 3574 18908 3626
rect 19068 3574 19120 3626
rect 19279 3574 19331 3626
rect 19489 3574 19541 3626
rect 19943 3574 19995 3626
rect 20154 3623 20206 3626
rect 20365 3623 20417 3626
rect 21913 3623 21965 3626
rect 22124 3623 22176 3626
rect 22335 3623 22387 3626
rect 22545 3623 22597 3626
rect 22756 3623 22808 3626
rect 22968 3623 23020 3626
rect 23179 3623 23231 3626
rect 20154 3577 20168 3623
rect 20168 3577 20206 3623
rect 20365 3577 20374 3623
rect 20374 3577 20417 3623
rect 21913 3577 21965 3623
rect 22124 3577 22176 3623
rect 22335 3577 22387 3623
rect 22545 3577 22597 3623
rect 22756 3577 22808 3623
rect 22968 3577 23020 3623
rect 23179 3577 23231 3623
rect 20154 3574 20206 3577
rect 20365 3574 20417 3577
rect 9372 3353 9383 3388
rect 9383 3353 9424 3388
rect 9372 3336 9424 3353
rect 9591 3121 9643 3173
rect 9591 2935 9643 2987
rect 21913 3574 21965 3577
rect 22124 3574 22176 3577
rect 22335 3574 22387 3577
rect 22545 3574 22597 3577
rect 22756 3574 22808 3577
rect 22968 3574 23020 3577
rect 23179 3574 23231 3577
rect 23389 3574 23441 3626
rect 23600 3574 23652 3626
rect 23811 3574 23863 3626
rect 11532 3336 11584 3388
rect 20670 3399 20722 3402
rect 20850 3399 20902 3402
rect 13042 3105 13094 3157
rect 20670 3353 20683 3399
rect 20683 3353 20722 3399
rect 20850 3353 20889 3399
rect 20889 3353 20902 3399
rect 18540 3312 18592 3327
rect 18751 3312 18803 3327
rect 18962 3312 19014 3327
rect 19173 3312 19225 3327
rect 19384 3312 19436 3327
rect 18540 3275 18581 3312
rect 18581 3275 18592 3312
rect 18751 3275 18787 3312
rect 18787 3275 18803 3312
rect 18962 3275 18993 3312
rect 18993 3275 19014 3312
rect 19173 3275 19199 3312
rect 19199 3275 19225 3312
rect 19384 3275 19436 3312
rect 20670 3350 20722 3353
rect 20850 3350 20902 3353
rect 14536 3129 14568 3164
rect 14568 3129 14588 3164
rect 14748 3129 14794 3164
rect 14794 3129 14800 3164
rect 18193 3168 18245 3220
rect 14536 3112 14588 3129
rect 14748 3112 14800 3129
rect 16705 2996 16757 3048
rect 19897 3112 19949 3164
rect 20108 3129 20110 3164
rect 20110 3129 20160 3164
rect 20108 3112 20160 3129
rect 20319 3112 20371 3164
rect 18193 2950 18245 3002
rect 21432 3353 21484 3395
rect 21612 3353 21664 3395
rect 21432 3343 21484 3353
rect 21612 3343 21664 3353
rect 4929 2818 4981 2864
rect 5140 2818 5177 2864
rect 5177 2818 5192 2864
rect 5351 2818 5383 2864
rect 5383 2818 5403 2864
rect 5562 2818 5589 2864
rect 5589 2818 5614 2864
rect 5773 2818 5795 2864
rect 5795 2818 5825 2864
rect 7488 2818 7506 2862
rect 7506 2818 7540 2862
rect 7668 2818 7669 2862
rect 7669 2818 7720 2862
rect 18540 2818 18581 2864
rect 18581 2818 18592 2864
rect 18751 2818 18787 2864
rect 18787 2818 18803 2864
rect 18962 2818 18993 2864
rect 18993 2818 19014 2864
rect 19173 2818 19199 2864
rect 19199 2818 19225 2864
rect 19384 2818 19436 2864
rect 21432 2905 21484 2932
rect 21612 2905 21664 2932
rect 21432 2880 21484 2905
rect 21612 2880 21664 2905
rect 4929 2812 4981 2818
rect 5140 2812 5192 2818
rect 5351 2812 5403 2818
rect 5562 2812 5614 2818
rect 5773 2812 5825 2818
rect 7488 2810 7540 2818
rect 7668 2810 7720 2818
rect 451 2674 503 2726
rect 662 2674 714 2726
rect 873 2674 925 2726
rect 1083 2674 1135 2726
rect 1294 2674 1346 2726
rect 1506 2674 1558 2726
rect 1717 2674 1769 2726
rect 1927 2674 1979 2726
rect 2138 2674 2190 2726
rect 2349 2674 2401 2726
rect 18540 2812 18592 2818
rect 18751 2812 18803 2818
rect 18962 2812 19014 2818
rect 19173 2812 19225 2818
rect 19384 2812 19436 2818
rect 4352 2674 4404 2726
rect 4532 2723 4584 2726
rect 4532 2677 4559 2723
rect 4559 2677 4584 2723
rect 4532 2674 4584 2677
rect 19735 2723 19787 2726
rect 19735 2677 19757 2723
rect 19757 2677 19787 2723
rect 19735 2674 19787 2677
rect 19915 2674 19967 2726
rect 4929 2582 4981 2588
rect 5140 2582 5192 2588
rect 5351 2582 5403 2588
rect 5562 2582 5614 2588
rect 5773 2582 5825 2588
rect 7488 2582 7540 2590
rect 7668 2582 7720 2590
rect 21913 2674 21965 2726
rect 22124 2674 22176 2726
rect 22335 2674 22387 2726
rect 22545 2674 22597 2726
rect 22756 2674 22808 2726
rect 22968 2674 23020 2726
rect 23179 2674 23231 2726
rect 23389 2674 23441 2726
rect 23600 2674 23652 2726
rect 23811 2674 23863 2726
rect 18540 2582 18592 2588
rect 18751 2582 18803 2588
rect 18962 2582 19014 2588
rect 19173 2582 19225 2588
rect 19384 2582 19436 2588
rect 2654 2495 2706 2498
rect 2834 2495 2886 2498
rect 4929 2536 4981 2582
rect 5140 2536 5177 2582
rect 5177 2536 5192 2582
rect 5351 2536 5383 2582
rect 5383 2536 5403 2582
rect 5562 2536 5589 2582
rect 5589 2536 5614 2582
rect 5773 2536 5795 2582
rect 5795 2536 5825 2582
rect 7488 2538 7506 2582
rect 7506 2538 7540 2582
rect 7668 2538 7669 2582
rect 7669 2538 7720 2582
rect 2654 2449 2706 2495
rect 2834 2449 2886 2495
rect 2654 2446 2706 2449
rect 2834 2446 2886 2449
rect 2654 2047 2706 2050
rect 2834 2047 2886 2050
rect 2654 2001 2706 2047
rect 2834 2001 2886 2047
rect 2654 1998 2706 2001
rect 2834 1998 2886 2001
rect 3864 2271 3916 2288
rect 4044 2271 4096 2288
rect 4224 2271 4276 2288
rect 3864 2236 3899 2271
rect 3899 2236 3916 2271
rect 4044 2236 4048 2271
rect 4048 2236 4096 2271
rect 4224 2236 4255 2271
rect 4255 2236 4276 2271
rect 6275 2311 6294 2363
rect 6294 2311 6327 2363
rect 18540 2536 18581 2582
rect 18581 2536 18592 2582
rect 18751 2536 18787 2582
rect 18787 2536 18803 2582
rect 18962 2536 18993 2582
rect 18993 2536 19014 2582
rect 19173 2536 19199 2582
rect 19199 2536 19225 2582
rect 19384 2536 19436 2582
rect 9591 2413 9643 2465
rect 6558 2312 6568 2356
rect 6568 2312 6610 2356
rect 6769 2312 6803 2356
rect 6803 2312 6821 2356
rect 6558 2304 6610 2312
rect 6769 2304 6821 2312
rect 6981 2304 7033 2356
rect 7192 2304 7244 2356
rect 4929 2088 4981 2128
rect 5140 2088 5177 2128
rect 5177 2088 5192 2128
rect 5351 2088 5383 2128
rect 5383 2088 5403 2128
rect 5562 2088 5589 2128
rect 5589 2088 5614 2128
rect 5773 2088 5795 2128
rect 5795 2088 5825 2128
rect 7488 2088 7506 2116
rect 7506 2088 7540 2116
rect 7668 2088 7669 2116
rect 7669 2088 7720 2116
rect 4929 2076 4981 2088
rect 5140 2076 5192 2088
rect 5351 2076 5403 2088
rect 5562 2076 5614 2088
rect 5773 2076 5825 2088
rect 3416 2001 3430 2042
rect 3430 2001 3468 2042
rect 3596 2001 3636 2042
rect 3636 2001 3648 2042
rect 7488 2064 7540 2088
rect 7668 2064 7720 2088
rect 3416 1990 3468 2001
rect 3596 1990 3648 2001
rect 451 1774 503 1826
rect 662 1774 714 1826
rect 873 1774 925 1826
rect 1083 1823 1135 1826
rect 1294 1823 1346 1826
rect 1506 1823 1558 1826
rect 1717 1823 1769 1826
rect 1927 1823 1979 1826
rect 2138 1823 2190 1826
rect 2349 1823 2401 1826
rect 3881 1823 3933 1826
rect 4092 1823 4144 1826
rect 1083 1777 1135 1823
rect 1294 1777 1346 1823
rect 1506 1777 1558 1823
rect 1717 1777 1769 1823
rect 1927 1777 1979 1823
rect 2138 1777 2190 1823
rect 2349 1777 2401 1823
rect 3881 1777 3899 1823
rect 3899 1777 3933 1823
rect 4092 1777 4105 1823
rect 4105 1777 4144 1823
rect 1083 1774 1135 1777
rect 1294 1774 1346 1777
rect 1506 1774 1558 1777
rect 1717 1774 1769 1777
rect 1927 1774 1979 1777
rect 2138 1774 2190 1777
rect 2349 1774 2401 1777
rect 3881 1774 3933 1777
rect 4092 1774 4144 1777
rect 4304 1774 4356 1826
rect 4515 1774 4567 1826
rect 4817 1774 4869 1826
rect 5027 1774 5079 1826
rect 5238 1774 5290 1826
rect 5450 1774 5502 1826
rect 5661 1774 5713 1826
rect 5871 1774 5923 1826
rect 7927 1823 7979 1826
rect 7927 1777 7979 1823
rect 7927 1774 7979 1777
rect 8138 1774 8190 1826
rect 8349 1774 8401 1826
rect 8649 1823 8701 1826
rect 8829 1823 8881 1826
rect 8649 1777 8659 1823
rect 8659 1777 8701 1823
rect 8829 1777 8863 1823
rect 8863 1777 8881 1823
rect 8649 1774 8701 1777
rect 8829 1774 8881 1777
rect 2654 1599 2706 1602
rect 2834 1599 2886 1602
rect 2654 1553 2706 1599
rect 2834 1553 2886 1599
rect 2654 1550 2706 1553
rect 2834 1550 2886 1553
rect 3416 1599 3468 1610
rect 3596 1599 3648 1610
rect 3416 1558 3430 1599
rect 3430 1558 3468 1599
rect 3596 1558 3636 1599
rect 3636 1558 3648 1599
rect 4929 1512 4981 1524
rect 5140 1512 5192 1524
rect 5351 1512 5403 1524
rect 5562 1512 5614 1524
rect 5773 1512 5825 1524
rect 7488 1512 7540 1536
rect 7668 1512 7720 1536
rect 4929 1472 4981 1512
rect 5140 1472 5177 1512
rect 5177 1472 5192 1512
rect 5351 1472 5383 1512
rect 5383 1472 5403 1512
rect 5562 1472 5589 1512
rect 5589 1472 5614 1512
rect 5773 1472 5795 1512
rect 5795 1472 5825 1512
rect 7488 1484 7506 1512
rect 7506 1484 7540 1512
rect 7668 1484 7669 1512
rect 7669 1484 7720 1512
rect 3864 1329 3899 1364
rect 3899 1329 3916 1364
rect 4044 1329 4048 1364
rect 4048 1329 4096 1364
rect 4224 1329 4255 1364
rect 4255 1329 4276 1364
rect 3864 1312 3916 1329
rect 4044 1312 4096 1329
rect 4224 1312 4276 1329
rect 2654 1151 2706 1154
rect 2834 1151 2886 1154
rect 2654 1105 2706 1151
rect 2834 1105 2886 1151
rect 2654 1102 2706 1105
rect 2834 1102 2886 1105
rect 6275 1237 6294 1289
rect 6294 1237 6327 1289
rect 6558 1288 6610 1296
rect 6769 1288 6821 1296
rect 6558 1244 6568 1288
rect 6568 1244 6610 1288
rect 6769 1244 6803 1288
rect 6803 1244 6821 1288
rect 6981 1244 7033 1296
rect 7192 1244 7244 1296
rect 9591 2227 9643 2279
rect 9372 2047 9424 2064
rect 9372 2012 9383 2047
rect 9383 2012 9424 2047
rect 13042 2243 13094 2295
rect 11532 2012 11584 2064
rect 17083 2352 17135 2404
rect 18193 2398 18245 2450
rect 21432 2495 21484 2520
rect 21612 2495 21664 2520
rect 21432 2468 21484 2495
rect 21612 2468 21664 2495
rect 14536 2271 14588 2288
rect 14748 2271 14800 2288
rect 14536 2236 14568 2271
rect 14568 2236 14588 2271
rect 14748 2236 14794 2271
rect 14794 2236 14800 2271
rect 18193 2180 18245 2232
rect 19897 2236 19949 2288
rect 20108 2271 20160 2288
rect 20108 2236 20110 2271
rect 20110 2236 20160 2271
rect 20319 2236 20371 2288
rect 18540 2088 18581 2125
rect 18581 2088 18592 2125
rect 18751 2088 18787 2125
rect 18787 2088 18803 2125
rect 18962 2088 18993 2125
rect 18993 2088 19014 2125
rect 19173 2088 19199 2125
rect 19199 2088 19225 2125
rect 19384 2088 19436 2125
rect 18540 2073 18592 2088
rect 18751 2073 18803 2088
rect 18962 2073 19014 2088
rect 19173 2073 19225 2088
rect 19384 2073 19436 2088
rect 20670 2047 20722 2050
rect 20850 2047 20902 2050
rect 20670 2001 20683 2047
rect 20683 2001 20722 2047
rect 20850 2001 20889 2047
rect 20889 2001 20902 2047
rect 20670 1998 20722 2001
rect 20850 1998 20902 2001
rect 21432 2047 21484 2057
rect 21612 2047 21664 2057
rect 21432 2005 21484 2047
rect 21612 2005 21664 2047
rect 9850 1774 9902 1826
rect 10030 1774 10082 1826
rect 13387 1774 13439 1826
rect 13598 1774 13650 1826
rect 13810 1823 13862 1826
rect 13810 1777 13833 1823
rect 13833 1777 13862 1823
rect 13810 1774 13862 1777
rect 14021 1774 14073 1826
rect 14431 1823 14483 1826
rect 14642 1823 14694 1826
rect 14853 1823 14905 1826
rect 14431 1777 14455 1823
rect 14455 1777 14483 1823
rect 14642 1777 14681 1823
rect 14681 1777 14694 1823
rect 14853 1777 14861 1823
rect 14861 1777 14905 1823
rect 14431 1774 14483 1777
rect 14642 1774 14694 1777
rect 14853 1774 14905 1777
rect 18435 1774 18487 1826
rect 18645 1774 18697 1826
rect 18856 1774 18908 1826
rect 19068 1774 19120 1826
rect 19279 1774 19331 1826
rect 19489 1774 19541 1826
rect 19943 1774 19995 1826
rect 20154 1823 20206 1826
rect 20365 1823 20417 1826
rect 21913 1823 21965 1826
rect 22124 1823 22176 1826
rect 22335 1823 22387 1826
rect 22545 1823 22597 1826
rect 22756 1823 22808 1826
rect 22968 1823 23020 1826
rect 23179 1823 23231 1826
rect 20154 1777 20168 1823
rect 20168 1777 20206 1823
rect 20365 1777 20374 1823
rect 20374 1777 20417 1823
rect 21913 1777 21965 1823
rect 22124 1777 22176 1823
rect 22335 1777 22387 1823
rect 22545 1777 22597 1823
rect 22756 1777 22808 1823
rect 22968 1777 23020 1823
rect 23179 1777 23231 1823
rect 20154 1774 20206 1777
rect 20365 1774 20417 1777
rect 9372 1553 9383 1588
rect 9383 1553 9424 1588
rect 9372 1536 9424 1553
rect 9591 1321 9643 1373
rect 9591 1135 9643 1187
rect 21913 1774 21965 1777
rect 22124 1774 22176 1777
rect 22335 1774 22387 1777
rect 22545 1774 22597 1777
rect 22756 1774 22808 1777
rect 22968 1774 23020 1777
rect 23179 1774 23231 1777
rect 23389 1774 23441 1826
rect 23600 1774 23652 1826
rect 23811 1774 23863 1826
rect 11532 1536 11584 1588
rect 20670 1599 20722 1602
rect 20850 1599 20902 1602
rect 13042 1305 13094 1357
rect 20670 1553 20683 1599
rect 20683 1553 20722 1599
rect 20850 1553 20889 1599
rect 20889 1553 20902 1599
rect 18540 1512 18592 1527
rect 18751 1512 18803 1527
rect 18962 1512 19014 1527
rect 19173 1512 19225 1527
rect 19384 1512 19436 1527
rect 18540 1475 18581 1512
rect 18581 1475 18592 1512
rect 18751 1475 18787 1512
rect 18787 1475 18803 1512
rect 18962 1475 18993 1512
rect 18993 1475 19014 1512
rect 19173 1475 19199 1512
rect 19199 1475 19225 1512
rect 19384 1475 19436 1512
rect 20670 1550 20722 1553
rect 20850 1550 20902 1553
rect 14536 1329 14568 1364
rect 14568 1329 14588 1364
rect 14748 1329 14794 1364
rect 14794 1329 14800 1364
rect 18193 1368 18245 1420
rect 14536 1312 14588 1329
rect 14748 1312 14800 1329
rect 17461 1196 17513 1248
rect 19897 1312 19949 1364
rect 20108 1329 20110 1364
rect 20110 1329 20160 1364
rect 20108 1312 20160 1329
rect 20319 1312 20371 1364
rect 18193 1150 18245 1202
rect 21432 1553 21484 1595
rect 21612 1553 21664 1595
rect 21432 1543 21484 1553
rect 21612 1543 21664 1553
rect 4929 1018 4981 1064
rect 5140 1018 5177 1064
rect 5177 1018 5192 1064
rect 5351 1018 5383 1064
rect 5383 1018 5403 1064
rect 5562 1018 5589 1064
rect 5589 1018 5614 1064
rect 5773 1018 5795 1064
rect 5795 1018 5825 1064
rect 7488 1018 7506 1062
rect 7506 1018 7540 1062
rect 7668 1018 7669 1062
rect 7669 1018 7720 1062
rect 18540 1018 18581 1064
rect 18581 1018 18592 1064
rect 18751 1018 18787 1064
rect 18787 1018 18803 1064
rect 18962 1018 18993 1064
rect 18993 1018 19014 1064
rect 19173 1018 19199 1064
rect 19199 1018 19225 1064
rect 19384 1018 19436 1064
rect 21432 1105 21484 1132
rect 21612 1105 21664 1132
rect 21432 1080 21484 1105
rect 21612 1080 21664 1105
rect 4929 1012 4981 1018
rect 5140 1012 5192 1018
rect 5351 1012 5403 1018
rect 5562 1012 5614 1018
rect 5773 1012 5825 1018
rect 7488 1010 7540 1018
rect 7668 1010 7720 1018
rect 451 874 503 926
rect 662 874 714 926
rect 873 874 925 926
rect 1083 874 1135 926
rect 1294 874 1346 926
rect 1506 874 1558 926
rect 1717 874 1769 926
rect 1927 874 1979 926
rect 2138 874 2190 926
rect 2349 874 2401 926
rect 18540 1012 18592 1018
rect 18751 1012 18803 1018
rect 18962 1012 19014 1018
rect 19173 1012 19225 1018
rect 19384 1012 19436 1018
rect 4352 874 4404 926
rect 4532 923 4584 926
rect 4532 877 4559 923
rect 4559 877 4584 923
rect 4532 874 4584 877
rect 19735 923 19787 926
rect 19735 877 19757 923
rect 19757 877 19787 923
rect 19735 874 19787 877
rect 19915 874 19967 926
rect 4929 782 4981 788
rect 5140 782 5192 788
rect 5351 782 5403 788
rect 5562 782 5614 788
rect 5773 782 5825 788
rect 7488 782 7540 790
rect 7668 782 7720 790
rect 21913 874 21965 926
rect 22124 874 22176 926
rect 22335 874 22387 926
rect 22545 874 22597 926
rect 22756 874 22808 926
rect 22968 874 23020 926
rect 23179 874 23231 926
rect 23389 874 23441 926
rect 23600 874 23652 926
rect 23811 874 23863 926
rect 18540 782 18592 788
rect 18751 782 18803 788
rect 18962 782 19014 788
rect 19173 782 19225 788
rect 19384 782 19436 788
rect 2654 695 2706 698
rect 2834 695 2886 698
rect 4929 736 4981 782
rect 5140 736 5177 782
rect 5177 736 5192 782
rect 5351 736 5383 782
rect 5383 736 5403 782
rect 5562 736 5589 782
rect 5589 736 5614 782
rect 5773 736 5795 782
rect 5795 736 5825 782
rect 7488 738 7506 782
rect 7506 738 7540 782
rect 7668 738 7669 782
rect 7669 738 7720 782
rect 2654 649 2706 695
rect 2834 649 2886 695
rect 2654 646 2706 649
rect 2834 646 2886 649
rect 2654 247 2706 250
rect 2834 247 2886 250
rect 2654 201 2706 247
rect 2834 201 2886 247
rect 2654 198 2706 201
rect 2834 198 2886 201
rect 3864 471 3916 488
rect 4044 471 4096 488
rect 4224 471 4276 488
rect 3864 436 3899 471
rect 3899 436 3916 471
rect 4044 436 4048 471
rect 4048 436 4096 471
rect 4224 436 4255 471
rect 4255 436 4276 471
rect 6275 511 6294 563
rect 6294 511 6327 563
rect 18540 736 18581 782
rect 18581 736 18592 782
rect 18751 736 18787 782
rect 18787 736 18803 782
rect 18962 736 18993 782
rect 18993 736 19014 782
rect 19173 736 19199 782
rect 19199 736 19225 782
rect 19384 736 19436 782
rect 9591 613 9643 665
rect 6558 512 6568 556
rect 6568 512 6610 556
rect 6769 512 6803 556
rect 6803 512 6821 556
rect 6558 504 6610 512
rect 6769 504 6821 512
rect 6981 504 7033 556
rect 7192 504 7244 556
rect 4929 288 4981 328
rect 5140 288 5177 328
rect 5177 288 5192 328
rect 5351 288 5383 328
rect 5383 288 5403 328
rect 5562 288 5589 328
rect 5589 288 5614 328
rect 5773 288 5795 328
rect 5795 288 5825 328
rect 7488 288 7506 316
rect 7506 288 7540 316
rect 7668 288 7669 316
rect 7669 288 7720 316
rect 4929 276 4981 288
rect 5140 276 5192 288
rect 5351 276 5403 288
rect 5562 276 5614 288
rect 5773 276 5825 288
rect 3416 201 3430 242
rect 3430 201 3468 242
rect 3596 201 3636 242
rect 3636 201 3648 242
rect 7488 264 7540 288
rect 7668 264 7720 288
rect 3416 190 3468 201
rect 3596 190 3648 201
rect 451 -26 503 26
rect 662 -26 714 26
rect 873 -26 925 26
rect 1083 23 1135 26
rect 1294 23 1346 26
rect 1506 23 1558 26
rect 1717 23 1769 26
rect 1927 23 1979 26
rect 2138 23 2190 26
rect 2349 23 2401 26
rect 3881 23 3933 26
rect 4092 23 4144 26
rect 1083 -23 1135 23
rect 1294 -23 1346 23
rect 1506 -23 1558 23
rect 1717 -23 1769 23
rect 1927 -23 1979 23
rect 2138 -23 2190 23
rect 2349 -23 2401 23
rect 3881 -23 3899 23
rect 3899 -23 3933 23
rect 4092 -23 4105 23
rect 4105 -23 4144 23
rect 1083 -26 1135 -23
rect 1294 -26 1346 -23
rect 1506 -26 1558 -23
rect 1717 -26 1769 -23
rect 1927 -26 1979 -23
rect 2138 -26 2190 -23
rect 2349 -26 2401 -23
rect 3881 -26 3933 -23
rect 4092 -26 4144 -23
rect 4304 -26 4356 26
rect 4515 -26 4567 26
rect 4817 -26 4869 26
rect 5027 -26 5079 26
rect 5238 -26 5290 26
rect 5450 -26 5502 26
rect 5661 -26 5713 26
rect 5871 -26 5923 26
rect 7927 23 7979 26
rect 7927 -23 7979 23
rect 7927 -26 7979 -23
rect 8138 -26 8190 26
rect 8349 -26 8401 26
rect 8649 23 8701 26
rect 8829 23 8881 26
rect 8649 -23 8659 23
rect 8659 -23 8701 23
rect 8829 -23 8863 23
rect 8863 -23 8881 23
rect 8649 -26 8701 -23
rect 8829 -26 8881 -23
rect 9591 427 9643 479
rect 9372 247 9424 264
rect 9372 212 9383 247
rect 9383 212 9424 247
rect 13042 443 13094 495
rect 11532 212 11584 264
rect 17838 552 17890 604
rect 18193 598 18245 650
rect 21432 695 21484 720
rect 21612 695 21664 720
rect 21432 668 21484 695
rect 21612 668 21664 695
rect 14536 471 14588 488
rect 14748 471 14800 488
rect 14536 436 14568 471
rect 14568 436 14588 471
rect 14748 436 14794 471
rect 14794 436 14800 471
rect 18193 380 18245 432
rect 19897 436 19949 488
rect 20108 471 20160 488
rect 20108 436 20110 471
rect 20110 436 20160 471
rect 20319 436 20371 488
rect 18540 288 18581 325
rect 18581 288 18592 325
rect 18751 288 18787 325
rect 18787 288 18803 325
rect 18962 288 18993 325
rect 18993 288 19014 325
rect 19173 288 19199 325
rect 19199 288 19225 325
rect 19384 288 19436 325
rect 18540 273 18592 288
rect 18751 273 18803 288
rect 18962 273 19014 288
rect 19173 273 19225 288
rect 19384 273 19436 288
rect 20670 247 20722 250
rect 20850 247 20902 250
rect 20670 201 20683 247
rect 20683 201 20722 247
rect 20850 201 20889 247
rect 20889 201 20902 247
rect 20670 198 20722 201
rect 20850 198 20902 201
rect 21432 247 21484 257
rect 21612 247 21664 257
rect 21432 205 21484 247
rect 21612 205 21664 247
rect 9850 -26 9902 26
rect 10030 -26 10082 26
rect 13387 -26 13439 26
rect 13598 -26 13650 26
rect 13810 23 13862 26
rect 13810 -23 13833 23
rect 13833 -23 13862 23
rect 13810 -26 13862 -23
rect 14021 -26 14073 26
rect 14431 23 14483 26
rect 14642 23 14694 26
rect 14853 23 14905 26
rect 14431 -23 14455 23
rect 14455 -23 14483 23
rect 14642 -23 14681 23
rect 14681 -23 14694 23
rect 14853 -23 14861 23
rect 14861 -23 14905 23
rect 14431 -26 14483 -23
rect 14642 -26 14694 -23
rect 14853 -26 14905 -23
rect 18435 -26 18487 26
rect 18645 -26 18697 26
rect 18856 -26 18908 26
rect 19068 -26 19120 26
rect 19279 -26 19331 26
rect 19489 -26 19541 26
rect 19943 -26 19995 26
rect 20154 23 20206 26
rect 20365 23 20417 26
rect 21913 23 21965 26
rect 22124 23 22176 26
rect 22335 23 22387 26
rect 22545 23 22597 26
rect 22756 23 22808 26
rect 22968 23 23020 26
rect 23179 23 23231 26
rect 20154 -23 20168 23
rect 20168 -23 20206 23
rect 20365 -23 20374 23
rect 20374 -23 20417 23
rect 21913 -23 21965 23
rect 22124 -23 22176 23
rect 22335 -23 22387 23
rect 22545 -23 22597 23
rect 22756 -23 22808 23
rect 22968 -23 23020 23
rect 23179 -23 23231 23
rect 20154 -26 20206 -23
rect 20365 -26 20417 -23
rect 21913 -26 21965 -23
rect 22124 -26 22176 -23
rect 22335 -26 22387 -23
rect 22545 -26 22597 -23
rect 22756 -26 22808 -23
rect 22968 -26 23020 -23
rect 23179 -26 23231 -23
rect 23389 -26 23441 26
rect 23600 -26 23652 26
rect 23811 -26 23863 26
<< metal2 >>
rect 367 14428 2486 14551
rect 367 14372 449 14428
rect 505 14372 660 14428
rect 716 14372 871 14428
rect 927 14372 1081 14428
rect 1137 14372 1292 14428
rect 1348 14372 1504 14428
rect 1560 14372 1715 14428
rect 1771 14372 1925 14428
rect 1981 14372 2136 14428
rect 2192 14372 2347 14428
rect 2403 14372 2486 14428
rect 367 13526 2486 14372
rect 3825 14426 4622 14551
rect 3825 14374 3881 14426
rect 3933 14374 4092 14426
rect 4144 14374 4304 14426
rect 4356 14374 4515 14426
rect 4567 14374 4622 14426
rect 2616 14202 2924 14243
rect 2616 14150 2654 14202
rect 2706 14150 2834 14202
rect 2886 14150 2924 14202
rect 2616 13995 2924 14150
rect 2616 13939 2652 13995
rect 2708 13939 2832 13995
rect 2888 13939 2924 13995
rect 2616 13754 2924 13939
rect 3328 14210 3687 14251
rect 3328 14158 3416 14210
rect 3468 14158 3596 14210
rect 3648 14158 3687 14210
rect 3328 13988 3687 14158
rect 3328 13932 3414 13988
rect 3470 13932 3594 13988
rect 3650 13932 3687 13988
rect 3328 13859 3687 13932
rect 3825 13964 4622 14374
rect 3825 13912 3864 13964
rect 3916 13912 4044 13964
rect 4096 13912 4224 13964
rect 4276 13912 4622 13964
rect 2616 13702 2654 13754
rect 2706 13702 2834 13754
rect 2886 13702 2924 13754
rect 2616 13662 2924 13702
rect 367 13474 451 13526
rect 503 13474 662 13526
rect 714 13474 873 13526
rect 925 13474 1083 13526
rect 1135 13474 1294 13526
rect 1346 13474 1506 13526
rect 1558 13474 1717 13526
rect 1769 13474 1927 13526
rect 1979 13474 2138 13526
rect 2190 13474 2349 13526
rect 2401 13474 2486 13526
rect 367 12628 2486 13474
rect 3825 13528 4622 13912
rect 3825 13472 3879 13528
rect 3935 13472 4090 13528
rect 4146 13472 4302 13528
rect 4358 13526 4513 13528
rect 4569 13526 4622 13528
rect 4404 13474 4513 13526
rect 4584 13474 4622 13526
rect 4358 13472 4513 13474
rect 4569 13472 4622 13474
rect 2616 13298 2924 13338
rect 2616 13246 2654 13298
rect 2706 13246 2834 13298
rect 2886 13246 2924 13298
rect 2616 13061 2924 13246
rect 2616 13005 2652 13061
rect 2708 13005 2832 13061
rect 2888 13005 2924 13061
rect 2616 12850 2924 13005
rect 2616 12798 2654 12850
rect 2706 12798 2834 12850
rect 2886 12798 2924 12850
rect 2616 12757 2924 12798
rect 3328 13068 3687 13141
rect 3328 13012 3414 13068
rect 3470 13012 3594 13068
rect 3650 13012 3687 13068
rect 3328 12842 3687 13012
rect 3328 12790 3416 12842
rect 3468 12790 3596 12842
rect 3648 12790 3687 12842
rect 3328 12749 3687 12790
rect 3825 13088 4622 13472
rect 3825 13036 3864 13088
rect 3916 13036 4044 13088
rect 4096 13036 4224 13088
rect 4276 13036 4622 13088
rect 367 12572 449 12628
rect 505 12572 660 12628
rect 716 12572 871 12628
rect 927 12572 1081 12628
rect 1137 12572 1292 12628
rect 1348 12572 1504 12628
rect 1560 12572 1715 12628
rect 1771 12572 1925 12628
rect 1981 12572 2136 12628
rect 2192 12572 2347 12628
rect 2403 12572 2486 12628
rect 367 11726 2486 12572
rect 3825 12626 4622 13036
rect 3825 12574 3881 12626
rect 3933 12574 4092 12626
rect 4144 12574 4304 12626
rect 4356 12574 4515 12626
rect 4567 12574 4622 12626
rect 2616 12402 2924 12443
rect 2616 12350 2654 12402
rect 2706 12350 2834 12402
rect 2886 12350 2924 12402
rect 2616 12195 2924 12350
rect 2616 12139 2652 12195
rect 2708 12139 2832 12195
rect 2888 12139 2924 12195
rect 2616 11954 2924 12139
rect 3328 12410 3687 12451
rect 3328 12358 3416 12410
rect 3468 12358 3596 12410
rect 3648 12358 3687 12410
rect 3328 12188 3687 12358
rect 3328 12132 3414 12188
rect 3470 12132 3594 12188
rect 3650 12132 3687 12188
rect 3328 12059 3687 12132
rect 3825 12164 4622 12574
rect 3825 12112 3864 12164
rect 3916 12112 4044 12164
rect 4096 12112 4224 12164
rect 4276 12112 4622 12164
rect 2616 11902 2654 11954
rect 2706 11902 2834 11954
rect 2886 11902 2924 11954
rect 2616 11862 2924 11902
rect 367 11674 451 11726
rect 503 11674 662 11726
rect 714 11674 873 11726
rect 925 11674 1083 11726
rect 1135 11674 1294 11726
rect 1346 11674 1506 11726
rect 1558 11674 1717 11726
rect 1769 11674 1927 11726
rect 1979 11674 2138 11726
rect 2190 11674 2349 11726
rect 2401 11674 2486 11726
rect 367 10828 2486 11674
rect 3825 11728 4622 12112
rect 3825 11672 3879 11728
rect 3935 11672 4090 11728
rect 4146 11672 4302 11728
rect 4358 11726 4513 11728
rect 4569 11726 4622 11728
rect 4404 11674 4513 11726
rect 4584 11674 4622 11726
rect 4358 11672 4513 11674
rect 4569 11672 4622 11674
rect 2616 11498 2924 11538
rect 2616 11446 2654 11498
rect 2706 11446 2834 11498
rect 2886 11446 2924 11498
rect 2616 11261 2924 11446
rect 2616 11205 2652 11261
rect 2708 11205 2832 11261
rect 2888 11205 2924 11261
rect 2616 11050 2924 11205
rect 2616 10998 2654 11050
rect 2706 10998 2834 11050
rect 2886 10998 2924 11050
rect 2616 10957 2924 10998
rect 3328 11268 3687 11341
rect 3328 11212 3414 11268
rect 3470 11212 3594 11268
rect 3650 11212 3687 11268
rect 3328 11042 3687 11212
rect 3328 10990 3416 11042
rect 3468 10990 3596 11042
rect 3648 10990 3687 11042
rect 3328 10949 3687 10990
rect 3825 11288 4622 11672
rect 3825 11236 3864 11288
rect 3916 11236 4044 11288
rect 4096 11236 4224 11288
rect 4276 11236 4622 11288
rect 367 10772 449 10828
rect 505 10772 660 10828
rect 716 10772 871 10828
rect 927 10772 1081 10828
rect 1137 10772 1292 10828
rect 1348 10772 1504 10828
rect 1560 10772 1715 10828
rect 1771 10772 1925 10828
rect 1981 10772 2136 10828
rect 2192 10772 2347 10828
rect 2403 10772 2486 10828
rect 367 9926 2486 10772
rect 3825 10826 4622 11236
rect 3825 10774 3881 10826
rect 3933 10774 4092 10826
rect 4144 10774 4304 10826
rect 4356 10774 4515 10826
rect 4567 10774 4622 10826
rect 2616 10602 2924 10643
rect 2616 10550 2654 10602
rect 2706 10550 2834 10602
rect 2886 10550 2924 10602
rect 2616 10395 2924 10550
rect 2616 10339 2652 10395
rect 2708 10339 2832 10395
rect 2888 10339 2924 10395
rect 2616 10154 2924 10339
rect 3328 10610 3687 10651
rect 3328 10558 3416 10610
rect 3468 10558 3596 10610
rect 3648 10558 3687 10610
rect 3328 10388 3687 10558
rect 3328 10332 3414 10388
rect 3470 10332 3594 10388
rect 3650 10332 3687 10388
rect 3328 10259 3687 10332
rect 3825 10364 4622 10774
rect 3825 10312 3864 10364
rect 3916 10312 4044 10364
rect 4096 10312 4224 10364
rect 4276 10312 4622 10364
rect 2616 10102 2654 10154
rect 2706 10102 2834 10154
rect 2886 10102 2924 10154
rect 2616 10062 2924 10102
rect 367 9874 451 9926
rect 503 9874 662 9926
rect 714 9874 873 9926
rect 925 9874 1083 9926
rect 1135 9874 1294 9926
rect 1346 9874 1506 9926
rect 1558 9874 1717 9926
rect 1769 9874 1927 9926
rect 1979 9874 2138 9926
rect 2190 9874 2349 9926
rect 2401 9874 2486 9926
rect 367 9028 2486 9874
rect 3825 9928 4622 10312
rect 3825 9872 3879 9928
rect 3935 9872 4090 9928
rect 4146 9872 4302 9928
rect 4358 9926 4513 9928
rect 4569 9926 4622 9928
rect 4404 9874 4513 9926
rect 4584 9874 4622 9926
rect 4358 9872 4513 9874
rect 4569 9872 4622 9874
rect 2616 9698 2924 9738
rect 2616 9646 2654 9698
rect 2706 9646 2834 9698
rect 2886 9646 2924 9698
rect 2616 9461 2924 9646
rect 2616 9405 2652 9461
rect 2708 9405 2832 9461
rect 2888 9405 2924 9461
rect 2616 9250 2924 9405
rect 2616 9198 2654 9250
rect 2706 9198 2834 9250
rect 2886 9198 2924 9250
rect 2616 9157 2924 9198
rect 3328 9468 3687 9541
rect 3328 9412 3414 9468
rect 3470 9412 3594 9468
rect 3650 9412 3687 9468
rect 3328 9242 3687 9412
rect 3328 9190 3416 9242
rect 3468 9190 3596 9242
rect 3648 9190 3687 9242
rect 3328 9149 3687 9190
rect 3825 9488 4622 9872
rect 3825 9436 3864 9488
rect 3916 9436 4044 9488
rect 4096 9436 4224 9488
rect 4276 9436 4622 9488
rect 367 8972 449 9028
rect 505 8972 660 9028
rect 716 8972 871 9028
rect 927 8972 1081 9028
rect 1137 8972 1292 9028
rect 1348 8972 1504 9028
rect 1560 8972 1715 9028
rect 1771 8972 1925 9028
rect 1981 8972 2136 9028
rect 2192 8972 2347 9028
rect 2403 8972 2486 9028
rect 367 8126 2486 8972
rect 3825 9026 4622 9436
rect 3825 8974 3881 9026
rect 3933 8974 4092 9026
rect 4144 8974 4304 9026
rect 4356 8974 4515 9026
rect 4567 8974 4622 9026
rect 2616 8802 2924 8843
rect 2616 8750 2654 8802
rect 2706 8750 2834 8802
rect 2886 8750 2924 8802
rect 2616 8595 2924 8750
rect 2616 8539 2652 8595
rect 2708 8539 2832 8595
rect 2888 8539 2924 8595
rect 2616 8354 2924 8539
rect 3328 8810 3687 8851
rect 3328 8758 3416 8810
rect 3468 8758 3596 8810
rect 3648 8758 3687 8810
rect 3328 8588 3687 8758
rect 3328 8532 3414 8588
rect 3470 8532 3594 8588
rect 3650 8532 3687 8588
rect 3328 8459 3687 8532
rect 3825 8564 4622 8974
rect 3825 8512 3864 8564
rect 3916 8512 4044 8564
rect 4096 8512 4224 8564
rect 4276 8512 4622 8564
rect 2616 8302 2654 8354
rect 2706 8302 2834 8354
rect 2886 8302 2924 8354
rect 2616 8262 2924 8302
rect 367 8074 451 8126
rect 503 8074 662 8126
rect 714 8074 873 8126
rect 925 8074 1083 8126
rect 1135 8074 1294 8126
rect 1346 8074 1506 8126
rect 1558 8074 1717 8126
rect 1769 8074 1927 8126
rect 1979 8074 2138 8126
rect 2190 8074 2349 8126
rect 2401 8074 2486 8126
rect 367 7228 2486 8074
rect 3825 8128 4622 8512
rect 3825 8072 3879 8128
rect 3935 8072 4090 8128
rect 4146 8072 4302 8128
rect 4358 8126 4513 8128
rect 4569 8126 4622 8128
rect 4404 8074 4513 8126
rect 4584 8074 4622 8126
rect 4358 8072 4513 8074
rect 4569 8072 4622 8074
rect 2616 7898 2924 7938
rect 2616 7846 2654 7898
rect 2706 7846 2834 7898
rect 2886 7846 2924 7898
rect 2616 7661 2924 7846
rect 2616 7605 2652 7661
rect 2708 7605 2832 7661
rect 2888 7605 2924 7661
rect 2616 7450 2924 7605
rect 2616 7398 2654 7450
rect 2706 7398 2834 7450
rect 2886 7398 2924 7450
rect 2616 7357 2924 7398
rect 3328 7668 3687 7741
rect 3328 7612 3414 7668
rect 3470 7612 3594 7668
rect 3650 7612 3687 7668
rect 3328 7442 3687 7612
rect 3328 7390 3416 7442
rect 3468 7390 3596 7442
rect 3648 7390 3687 7442
rect 3328 7349 3687 7390
rect 3825 7688 4622 8072
rect 3825 7636 3864 7688
rect 3916 7636 4044 7688
rect 4096 7636 4224 7688
rect 4276 7636 4622 7688
rect 367 7172 449 7228
rect 505 7172 660 7228
rect 716 7172 871 7228
rect 927 7172 1081 7228
rect 1137 7172 1292 7228
rect 1348 7172 1504 7228
rect 1560 7172 1715 7228
rect 1771 7172 1925 7228
rect 1981 7172 2136 7228
rect 2192 7172 2347 7228
rect 2403 7172 2486 7228
rect 367 6326 2486 7172
rect 3825 7226 4622 7636
rect 3825 7174 3881 7226
rect 3933 7174 4092 7226
rect 4144 7174 4304 7226
rect 4356 7174 4515 7226
rect 4567 7174 4622 7226
rect 2616 7002 2924 7043
rect 2616 6950 2654 7002
rect 2706 6950 2834 7002
rect 2886 6950 2924 7002
rect 2616 6795 2924 6950
rect 2616 6739 2652 6795
rect 2708 6739 2832 6795
rect 2888 6739 2924 6795
rect 2616 6554 2924 6739
rect 3328 7010 3687 7051
rect 3328 6958 3416 7010
rect 3468 6958 3596 7010
rect 3648 6958 3687 7010
rect 3328 6788 3687 6958
rect 3328 6732 3414 6788
rect 3470 6732 3594 6788
rect 3650 6732 3687 6788
rect 3328 6659 3687 6732
rect 3825 6764 4622 7174
rect 3825 6712 3864 6764
rect 3916 6712 4044 6764
rect 4096 6712 4224 6764
rect 4276 6712 4622 6764
rect 2616 6502 2654 6554
rect 2706 6502 2834 6554
rect 2886 6502 2924 6554
rect 2616 6462 2924 6502
rect 367 6274 451 6326
rect 503 6274 662 6326
rect 714 6274 873 6326
rect 925 6274 1083 6326
rect 1135 6274 1294 6326
rect 1346 6274 1506 6326
rect 1558 6274 1717 6326
rect 1769 6274 1927 6326
rect 1979 6274 2138 6326
rect 2190 6274 2349 6326
rect 2401 6274 2486 6326
rect 367 5428 2486 6274
rect 3825 6328 4622 6712
rect 3825 6272 3879 6328
rect 3935 6272 4090 6328
rect 4146 6272 4302 6328
rect 4358 6326 4513 6328
rect 4569 6326 4622 6328
rect 4404 6274 4513 6326
rect 4584 6274 4622 6326
rect 4358 6272 4513 6274
rect 4569 6272 4622 6274
rect 2616 6098 2924 6138
rect 2616 6046 2654 6098
rect 2706 6046 2834 6098
rect 2886 6046 2924 6098
rect 2616 5861 2924 6046
rect 2616 5805 2652 5861
rect 2708 5805 2832 5861
rect 2888 5805 2924 5861
rect 2616 5650 2924 5805
rect 2616 5598 2654 5650
rect 2706 5598 2834 5650
rect 2886 5598 2924 5650
rect 2616 5557 2924 5598
rect 3328 5868 3687 5941
rect 3328 5812 3414 5868
rect 3470 5812 3594 5868
rect 3650 5812 3687 5868
rect 3328 5642 3687 5812
rect 3328 5590 3416 5642
rect 3468 5590 3596 5642
rect 3648 5590 3687 5642
rect 3328 5549 3687 5590
rect 3825 5888 4622 6272
rect 3825 5836 3864 5888
rect 3916 5836 4044 5888
rect 4096 5836 4224 5888
rect 4276 5836 4622 5888
rect 367 5372 449 5428
rect 505 5372 660 5428
rect 716 5372 871 5428
rect 927 5372 1081 5428
rect 1137 5372 1292 5428
rect 1348 5372 1504 5428
rect 1560 5372 1715 5428
rect 1771 5372 1925 5428
rect 1981 5372 2136 5428
rect 2192 5372 2347 5428
rect 2403 5372 2486 5428
rect 367 4526 2486 5372
rect 3825 5426 4622 5836
rect 3825 5374 3881 5426
rect 3933 5374 4092 5426
rect 4144 5374 4304 5426
rect 4356 5374 4515 5426
rect 4567 5374 4622 5426
rect 2616 5202 2924 5243
rect 2616 5150 2654 5202
rect 2706 5150 2834 5202
rect 2886 5150 2924 5202
rect 2616 4995 2924 5150
rect 2616 4939 2652 4995
rect 2708 4939 2832 4995
rect 2888 4939 2924 4995
rect 2616 4754 2924 4939
rect 3328 5210 3687 5251
rect 3328 5158 3416 5210
rect 3468 5158 3596 5210
rect 3648 5158 3687 5210
rect 3328 4988 3687 5158
rect 3328 4932 3414 4988
rect 3470 4932 3594 4988
rect 3650 4932 3687 4988
rect 3328 4859 3687 4932
rect 3825 4964 4622 5374
rect 3825 4912 3864 4964
rect 3916 4912 4044 4964
rect 4096 4912 4224 4964
rect 4276 4912 4622 4964
rect 2616 4702 2654 4754
rect 2706 4702 2834 4754
rect 2886 4702 2924 4754
rect 2616 4662 2924 4702
rect 367 4474 451 4526
rect 503 4474 662 4526
rect 714 4474 873 4526
rect 925 4474 1083 4526
rect 1135 4474 1294 4526
rect 1346 4474 1506 4526
rect 1558 4474 1717 4526
rect 1769 4474 1927 4526
rect 1979 4474 2138 4526
rect 2190 4474 2349 4526
rect 2401 4474 2486 4526
rect 367 3628 2486 4474
rect 3825 4528 4622 4912
rect 3825 4472 3879 4528
rect 3935 4472 4090 4528
rect 4146 4472 4302 4528
rect 4358 4526 4513 4528
rect 4569 4526 4622 4528
rect 4404 4474 4513 4526
rect 4584 4474 4622 4526
rect 4358 4472 4513 4474
rect 4569 4472 4622 4474
rect 2616 4298 2924 4338
rect 2616 4246 2654 4298
rect 2706 4246 2834 4298
rect 2886 4246 2924 4298
rect 2616 4061 2924 4246
rect 2616 4005 2652 4061
rect 2708 4005 2832 4061
rect 2888 4005 2924 4061
rect 2616 3850 2924 4005
rect 2616 3798 2654 3850
rect 2706 3798 2834 3850
rect 2886 3798 2924 3850
rect 2616 3757 2924 3798
rect 3328 4068 3687 4141
rect 3328 4012 3414 4068
rect 3470 4012 3594 4068
rect 3650 4012 3687 4068
rect 3328 3842 3687 4012
rect 3328 3790 3416 3842
rect 3468 3790 3596 3842
rect 3648 3790 3687 3842
rect 3328 3749 3687 3790
rect 3825 4088 4622 4472
rect 3825 4036 3864 4088
rect 3916 4036 4044 4088
rect 4096 4036 4224 4088
rect 4276 4036 4622 4088
rect 367 3572 449 3628
rect 505 3572 660 3628
rect 716 3572 871 3628
rect 927 3572 1081 3628
rect 1137 3572 1292 3628
rect 1348 3572 1504 3628
rect 1560 3572 1715 3628
rect 1771 3572 1925 3628
rect 1981 3572 2136 3628
rect 2192 3572 2347 3628
rect 2403 3572 2486 3628
rect 367 2726 2486 3572
rect 3825 3626 4622 4036
rect 3825 3574 3881 3626
rect 3933 3574 4092 3626
rect 4144 3574 4304 3626
rect 4356 3574 4515 3626
rect 4567 3574 4622 3626
rect 2616 3402 2924 3443
rect 2616 3350 2654 3402
rect 2706 3350 2834 3402
rect 2886 3350 2924 3402
rect 2616 3195 2924 3350
rect 2616 3139 2652 3195
rect 2708 3139 2832 3195
rect 2888 3139 2924 3195
rect 2616 2954 2924 3139
rect 3328 3410 3687 3451
rect 3328 3358 3416 3410
rect 3468 3358 3596 3410
rect 3648 3358 3687 3410
rect 3328 3188 3687 3358
rect 3328 3132 3414 3188
rect 3470 3132 3594 3188
rect 3650 3132 3687 3188
rect 3328 3059 3687 3132
rect 3825 3164 4622 3574
rect 3825 3112 3864 3164
rect 3916 3112 4044 3164
rect 4096 3112 4224 3164
rect 4276 3112 4622 3164
rect 2616 2902 2654 2954
rect 2706 2902 2834 2954
rect 2886 2902 2924 2954
rect 2616 2862 2924 2902
rect 367 2674 451 2726
rect 503 2674 662 2726
rect 714 2674 873 2726
rect 925 2674 1083 2726
rect 1135 2674 1294 2726
rect 1346 2674 1506 2726
rect 1558 2674 1717 2726
rect 1769 2674 1927 2726
rect 1979 2674 2138 2726
rect 2190 2674 2349 2726
rect 2401 2674 2486 2726
rect 367 1828 2486 2674
rect 3825 2728 4622 3112
rect 3825 2672 3879 2728
rect 3935 2672 4090 2728
rect 4146 2672 4302 2728
rect 4358 2726 4513 2728
rect 4569 2726 4622 2728
rect 4404 2674 4513 2726
rect 4584 2674 4622 2726
rect 4358 2672 4513 2674
rect 4569 2672 4622 2674
rect 2616 2498 2924 2538
rect 2616 2446 2654 2498
rect 2706 2446 2834 2498
rect 2886 2446 2924 2498
rect 2616 2261 2924 2446
rect 2616 2205 2652 2261
rect 2708 2205 2832 2261
rect 2888 2205 2924 2261
rect 2616 2050 2924 2205
rect 2616 1998 2654 2050
rect 2706 1998 2834 2050
rect 2886 1998 2924 2050
rect 2616 1957 2924 1998
rect 3328 2268 3687 2341
rect 3328 2212 3414 2268
rect 3470 2212 3594 2268
rect 3650 2212 3687 2268
rect 3328 2042 3687 2212
rect 3328 1990 3416 2042
rect 3468 1990 3596 2042
rect 3648 1990 3687 2042
rect 3328 1949 3687 1990
rect 3825 2288 4622 2672
rect 3825 2236 3864 2288
rect 3916 2236 4044 2288
rect 4096 2236 4224 2288
rect 4276 2236 4622 2288
rect 367 1772 449 1828
rect 505 1772 660 1828
rect 716 1772 871 1828
rect 927 1772 1081 1828
rect 1137 1772 1292 1828
rect 1348 1772 1504 1828
rect 1560 1772 1715 1828
rect 1771 1772 1925 1828
rect 1981 1772 2136 1828
rect 2192 1772 2347 1828
rect 2403 1772 2486 1828
rect 367 926 2486 1772
rect 3825 1826 4622 2236
rect 3825 1774 3881 1826
rect 3933 1774 4092 1826
rect 4144 1774 4304 1826
rect 4356 1774 4515 1826
rect 4567 1774 4622 1826
rect 2616 1602 2924 1643
rect 2616 1550 2654 1602
rect 2706 1550 2834 1602
rect 2886 1550 2924 1602
rect 2616 1395 2924 1550
rect 2616 1339 2652 1395
rect 2708 1339 2832 1395
rect 2888 1339 2924 1395
rect 2616 1154 2924 1339
rect 3328 1610 3687 1651
rect 3328 1558 3416 1610
rect 3468 1558 3596 1610
rect 3648 1558 3687 1610
rect 3328 1388 3687 1558
rect 3328 1332 3414 1388
rect 3470 1332 3594 1388
rect 3650 1332 3687 1388
rect 3328 1259 3687 1332
rect 3825 1364 4622 1774
rect 3825 1312 3864 1364
rect 3916 1312 4044 1364
rect 4096 1312 4224 1364
rect 4276 1312 4622 1364
rect 2616 1102 2654 1154
rect 2706 1102 2834 1154
rect 2886 1102 2924 1154
rect 2616 1062 2924 1102
rect 367 874 451 926
rect 503 874 662 926
rect 714 874 873 926
rect 925 874 1083 926
rect 1135 874 1294 926
rect 1346 874 1506 926
rect 1558 874 1717 926
rect 1769 874 1927 926
rect 1979 874 2138 926
rect 2190 874 2349 926
rect 2401 874 2486 926
rect 367 28 2486 874
rect 3825 928 4622 1312
rect 3825 872 3879 928
rect 3935 872 4090 928
rect 4146 872 4302 928
rect 4358 926 4513 928
rect 4569 926 4622 928
rect 4404 874 4513 926
rect 4584 874 4622 926
rect 4358 872 4513 874
rect 4569 872 4622 874
rect 2616 698 2924 738
rect 2616 646 2654 698
rect 2706 646 2834 698
rect 2886 646 2924 698
rect 2616 461 2924 646
rect 2616 405 2652 461
rect 2708 405 2832 461
rect 2888 405 2924 461
rect 2616 250 2924 405
rect 2616 198 2654 250
rect 2706 198 2834 250
rect 2886 198 2924 250
rect 2616 157 2924 198
rect 3328 468 3687 541
rect 3328 412 3414 468
rect 3470 412 3594 468
rect 3650 412 3687 468
rect 3328 242 3687 412
rect 3328 190 3416 242
rect 3468 190 3596 242
rect 3648 190 3687 242
rect 3328 149 3687 190
rect 3825 488 4622 872
rect 3825 436 3864 488
rect 3916 436 4044 488
rect 4096 436 4224 488
rect 4276 436 4622 488
rect 367 -28 449 28
rect 505 -28 660 28
rect 716 -28 871 28
rect 927 -28 1081 28
rect 1137 -28 1292 28
rect 1348 -28 1504 28
rect 1560 -28 1715 28
rect 1771 -28 1925 28
rect 1981 -28 2136 28
rect 2192 -28 2347 28
rect 2403 -28 2486 28
rect 367 -151 2486 -28
rect 3825 26 4622 436
rect 3825 -26 3881 26
rect 3933 -26 4092 26
rect 4144 -26 4304 26
rect 4356 -26 4515 26
rect 4567 -26 4622 26
rect 3825 -151 4622 -26
rect 4728 14428 6012 14551
rect 4728 14372 4815 14428
rect 4871 14372 5025 14428
rect 5081 14372 5236 14428
rect 5292 14372 5448 14428
rect 5504 14372 5659 14428
rect 5715 14372 5869 14428
rect 5925 14372 6012 14428
rect 4728 14124 6012 14372
rect 4728 14072 4929 14124
rect 4981 14072 5140 14124
rect 5192 14072 5351 14124
rect 5403 14072 5562 14124
rect 5614 14072 5773 14124
rect 5825 14072 6012 14124
rect 4728 13664 6012 14072
rect 6237 14036 6365 14075
rect 6237 13980 6273 14036
rect 6329 14013 6365 14036
rect 6329 13980 6366 14013
rect 6237 13889 6366 13980
rect 6237 13837 6275 13889
rect 6327 13837 6366 13889
rect 6237 13796 6366 13837
rect 6461 13896 7341 14551
rect 7866 14426 8461 14551
rect 7866 14374 7927 14426
rect 7979 14374 8138 14426
rect 8190 14374 8349 14426
rect 8401 14374 8461 14426
rect 6461 13844 6558 13896
rect 6610 13844 6769 13896
rect 6821 13844 6981 13896
rect 7033 13844 7192 13896
rect 7244 13844 7341 13896
rect 4728 13612 4929 13664
rect 4981 13612 5140 13664
rect 5192 13612 5351 13664
rect 5403 13612 5562 13664
rect 5614 13612 5773 13664
rect 5825 13612 6012 13664
rect 4728 13388 6012 13612
rect 4728 13336 4929 13388
rect 4981 13336 5140 13388
rect 5192 13336 5351 13388
rect 5403 13336 5562 13388
rect 5614 13336 5773 13388
rect 5825 13336 6012 13388
rect 4728 12928 6012 13336
rect 4728 12876 4929 12928
rect 4981 12876 5140 12928
rect 5192 12876 5351 12928
rect 5403 12876 5562 12928
rect 5614 12876 5773 12928
rect 5825 12876 6012 12928
rect 6237 13163 6366 13204
rect 6237 13111 6275 13163
rect 6327 13111 6366 13163
rect 6237 13020 6366 13111
rect 6237 12964 6273 13020
rect 6329 12987 6366 13020
rect 6461 13156 7341 13844
rect 7449 14136 7758 14177
rect 7449 14084 7488 14136
rect 7540 14084 7668 14136
rect 7720 14084 7758 14136
rect 7449 13805 7758 14084
rect 7449 13749 7486 13805
rect 7542 13749 7666 13805
rect 7722 13749 7758 13805
rect 7449 13662 7758 13749
rect 7449 13610 7488 13662
rect 7540 13610 7668 13662
rect 7720 13610 7758 13662
rect 7449 13569 7758 13610
rect 7866 13528 8461 14374
rect 7866 13472 7925 13528
rect 7981 13472 8136 13528
rect 8192 13472 8347 13528
rect 8403 13472 8461 13528
rect 6461 13104 6558 13156
rect 6610 13104 6769 13156
rect 6821 13104 6981 13156
rect 7033 13104 7192 13156
rect 7244 13104 7341 13156
rect 6329 12964 6365 12987
rect 6237 12925 6365 12964
rect 4728 12628 6012 12876
rect 4728 12572 4815 12628
rect 4871 12572 5025 12628
rect 5081 12572 5236 12628
rect 5292 12572 5448 12628
rect 5504 12572 5659 12628
rect 5715 12572 5869 12628
rect 5925 12572 6012 12628
rect 4728 12324 6012 12572
rect 4728 12272 4929 12324
rect 4981 12272 5140 12324
rect 5192 12272 5351 12324
rect 5403 12272 5562 12324
rect 5614 12272 5773 12324
rect 5825 12272 6012 12324
rect 4728 11864 6012 12272
rect 6237 12236 6365 12275
rect 6237 12180 6273 12236
rect 6329 12213 6365 12236
rect 6329 12180 6366 12213
rect 6237 12089 6366 12180
rect 6237 12037 6275 12089
rect 6327 12037 6366 12089
rect 6237 11996 6366 12037
rect 6461 12096 7341 13104
rect 7449 13390 7758 13431
rect 7449 13338 7488 13390
rect 7540 13338 7668 13390
rect 7720 13338 7758 13390
rect 7449 13251 7758 13338
rect 7449 13195 7486 13251
rect 7542 13195 7666 13251
rect 7722 13195 7758 13251
rect 7449 12916 7758 13195
rect 7449 12864 7488 12916
rect 7540 12864 7668 12916
rect 7720 12864 7758 12916
rect 7449 12823 7758 12864
rect 7866 12626 8461 13472
rect 7866 12574 7927 12626
rect 7979 12574 8138 12626
rect 8190 12574 8349 12626
rect 8401 12574 8461 12626
rect 6461 12044 6558 12096
rect 6610 12044 6769 12096
rect 6821 12044 6981 12096
rect 7033 12044 7192 12096
rect 7244 12044 7341 12096
rect 4728 11812 4929 11864
rect 4981 11812 5140 11864
rect 5192 11812 5351 11864
rect 5403 11812 5562 11864
rect 5614 11812 5773 11864
rect 5825 11812 6012 11864
rect 4728 11588 6012 11812
rect 4728 11536 4929 11588
rect 4981 11536 5140 11588
rect 5192 11536 5351 11588
rect 5403 11536 5562 11588
rect 5614 11536 5773 11588
rect 5825 11536 6012 11588
rect 4728 11128 6012 11536
rect 4728 11076 4929 11128
rect 4981 11076 5140 11128
rect 5192 11076 5351 11128
rect 5403 11076 5562 11128
rect 5614 11076 5773 11128
rect 5825 11076 6012 11128
rect 6237 11363 6366 11404
rect 6237 11311 6275 11363
rect 6327 11311 6366 11363
rect 6237 11220 6366 11311
rect 6237 11164 6273 11220
rect 6329 11187 6366 11220
rect 6461 11356 7341 12044
rect 7449 12336 7758 12377
rect 7449 12284 7488 12336
rect 7540 12284 7668 12336
rect 7720 12284 7758 12336
rect 7449 12005 7758 12284
rect 7449 11949 7486 12005
rect 7542 11949 7666 12005
rect 7722 11949 7758 12005
rect 7449 11862 7758 11949
rect 7449 11810 7488 11862
rect 7540 11810 7668 11862
rect 7720 11810 7758 11862
rect 7449 11769 7758 11810
rect 7866 11728 8461 12574
rect 7866 11672 7925 11728
rect 7981 11672 8136 11728
rect 8192 11672 8347 11728
rect 8403 11672 8461 11728
rect 6461 11304 6558 11356
rect 6610 11304 6769 11356
rect 6821 11304 6981 11356
rect 7033 11304 7192 11356
rect 7244 11304 7341 11356
rect 6329 11164 6365 11187
rect 6237 11125 6365 11164
rect 4728 10828 6012 11076
rect 4728 10772 4815 10828
rect 4871 10772 5025 10828
rect 5081 10772 5236 10828
rect 5292 10772 5448 10828
rect 5504 10772 5659 10828
rect 5715 10772 5869 10828
rect 5925 10772 6012 10828
rect 4728 10524 6012 10772
rect 4728 10472 4929 10524
rect 4981 10472 5140 10524
rect 5192 10472 5351 10524
rect 5403 10472 5562 10524
rect 5614 10472 5773 10524
rect 5825 10472 6012 10524
rect 4728 10064 6012 10472
rect 6237 10436 6365 10475
rect 6237 10380 6273 10436
rect 6329 10413 6365 10436
rect 6329 10380 6366 10413
rect 6237 10289 6366 10380
rect 6237 10237 6275 10289
rect 6327 10237 6366 10289
rect 6237 10196 6366 10237
rect 6461 10296 7341 11304
rect 7449 11590 7758 11631
rect 7449 11538 7488 11590
rect 7540 11538 7668 11590
rect 7720 11538 7758 11590
rect 7449 11451 7758 11538
rect 7449 11395 7486 11451
rect 7542 11395 7666 11451
rect 7722 11395 7758 11451
rect 7449 11116 7758 11395
rect 7449 11064 7488 11116
rect 7540 11064 7668 11116
rect 7720 11064 7758 11116
rect 7449 11023 7758 11064
rect 7866 10826 8461 11672
rect 7866 10774 7927 10826
rect 7979 10774 8138 10826
rect 8190 10774 8349 10826
rect 8401 10774 8461 10826
rect 6461 10244 6558 10296
rect 6610 10244 6769 10296
rect 6821 10244 6981 10296
rect 7033 10244 7192 10296
rect 7244 10244 7341 10296
rect 4728 10012 4929 10064
rect 4981 10012 5140 10064
rect 5192 10012 5351 10064
rect 5403 10012 5562 10064
rect 5614 10012 5773 10064
rect 5825 10012 6012 10064
rect 4728 9788 6012 10012
rect 4728 9736 4929 9788
rect 4981 9736 5140 9788
rect 5192 9736 5351 9788
rect 5403 9736 5562 9788
rect 5614 9736 5773 9788
rect 5825 9736 6012 9788
rect 4728 9328 6012 9736
rect 4728 9276 4929 9328
rect 4981 9276 5140 9328
rect 5192 9276 5351 9328
rect 5403 9276 5562 9328
rect 5614 9276 5773 9328
rect 5825 9276 6012 9328
rect 6237 9563 6366 9604
rect 6237 9511 6275 9563
rect 6327 9511 6366 9563
rect 6237 9420 6366 9511
rect 6237 9364 6273 9420
rect 6329 9387 6366 9420
rect 6461 9556 7341 10244
rect 7449 10536 7758 10577
rect 7449 10484 7488 10536
rect 7540 10484 7668 10536
rect 7720 10484 7758 10536
rect 7449 10205 7758 10484
rect 7449 10149 7486 10205
rect 7542 10149 7666 10205
rect 7722 10149 7758 10205
rect 7449 10062 7758 10149
rect 7449 10010 7488 10062
rect 7540 10010 7668 10062
rect 7720 10010 7758 10062
rect 7449 9969 7758 10010
rect 7866 9928 8461 10774
rect 7866 9872 7925 9928
rect 7981 9872 8136 9928
rect 8192 9872 8347 9928
rect 8403 9872 8461 9928
rect 6461 9504 6558 9556
rect 6610 9504 6769 9556
rect 6821 9504 6981 9556
rect 7033 9504 7192 9556
rect 7244 9504 7341 9556
rect 6329 9364 6365 9387
rect 6237 9325 6365 9364
rect 4728 9028 6012 9276
rect 4728 8972 4815 9028
rect 4871 8972 5025 9028
rect 5081 8972 5236 9028
rect 5292 8972 5448 9028
rect 5504 8972 5659 9028
rect 5715 8972 5869 9028
rect 5925 8972 6012 9028
rect 4728 8724 6012 8972
rect 4728 8672 4929 8724
rect 4981 8672 5140 8724
rect 5192 8672 5351 8724
rect 5403 8672 5562 8724
rect 5614 8672 5773 8724
rect 5825 8672 6012 8724
rect 4728 8264 6012 8672
rect 6237 8636 6365 8675
rect 6237 8580 6273 8636
rect 6329 8613 6365 8636
rect 6329 8580 6366 8613
rect 6237 8489 6366 8580
rect 6237 8437 6275 8489
rect 6327 8437 6366 8489
rect 6237 8396 6366 8437
rect 6461 8496 7341 9504
rect 7449 9790 7758 9831
rect 7449 9738 7488 9790
rect 7540 9738 7668 9790
rect 7720 9738 7758 9790
rect 7449 9651 7758 9738
rect 7449 9595 7486 9651
rect 7542 9595 7666 9651
rect 7722 9595 7758 9651
rect 7449 9316 7758 9595
rect 7449 9264 7488 9316
rect 7540 9264 7668 9316
rect 7720 9264 7758 9316
rect 7449 9223 7758 9264
rect 7866 9026 8461 9872
rect 7866 8974 7927 9026
rect 7979 8974 8138 9026
rect 8190 8974 8349 9026
rect 8401 8974 8461 9026
rect 6461 8444 6558 8496
rect 6610 8444 6769 8496
rect 6821 8444 6981 8496
rect 7033 8444 7192 8496
rect 7244 8444 7341 8496
rect 4728 8212 4929 8264
rect 4981 8212 5140 8264
rect 5192 8212 5351 8264
rect 5403 8212 5562 8264
rect 5614 8212 5773 8264
rect 5825 8212 6012 8264
rect 4728 7988 6012 8212
rect 4728 7936 4929 7988
rect 4981 7936 5140 7988
rect 5192 7936 5351 7988
rect 5403 7936 5562 7988
rect 5614 7936 5773 7988
rect 5825 7936 6012 7988
rect 4728 7528 6012 7936
rect 4728 7476 4929 7528
rect 4981 7476 5140 7528
rect 5192 7476 5351 7528
rect 5403 7476 5562 7528
rect 5614 7476 5773 7528
rect 5825 7476 6012 7528
rect 6237 7763 6366 7804
rect 6237 7711 6275 7763
rect 6327 7711 6366 7763
rect 6237 7620 6366 7711
rect 6237 7564 6273 7620
rect 6329 7587 6366 7620
rect 6461 7756 7341 8444
rect 7449 8736 7758 8777
rect 7449 8684 7488 8736
rect 7540 8684 7668 8736
rect 7720 8684 7758 8736
rect 7449 8405 7758 8684
rect 7449 8349 7486 8405
rect 7542 8349 7666 8405
rect 7722 8349 7758 8405
rect 7449 8262 7758 8349
rect 7449 8210 7488 8262
rect 7540 8210 7668 8262
rect 7720 8210 7758 8262
rect 7449 8169 7758 8210
rect 7866 8128 8461 8974
rect 7866 8072 7925 8128
rect 7981 8072 8136 8128
rect 8192 8072 8347 8128
rect 8403 8072 8461 8128
rect 6461 7704 6558 7756
rect 6610 7704 6769 7756
rect 6821 7704 6981 7756
rect 7033 7704 7192 7756
rect 7244 7704 7341 7756
rect 6329 7564 6365 7587
rect 6237 7525 6365 7564
rect 4728 7228 6012 7476
rect 4728 7172 4815 7228
rect 4871 7172 5025 7228
rect 5081 7172 5236 7228
rect 5292 7172 5448 7228
rect 5504 7172 5659 7228
rect 5715 7172 5869 7228
rect 5925 7172 6012 7228
rect 4728 6924 6012 7172
rect 4728 6872 4929 6924
rect 4981 6872 5140 6924
rect 5192 6872 5351 6924
rect 5403 6872 5562 6924
rect 5614 6872 5773 6924
rect 5825 6872 6012 6924
rect 4728 6464 6012 6872
rect 6237 6836 6365 6875
rect 6237 6780 6273 6836
rect 6329 6813 6365 6836
rect 6329 6780 6366 6813
rect 6237 6689 6366 6780
rect 6237 6637 6275 6689
rect 6327 6637 6366 6689
rect 6237 6596 6366 6637
rect 6461 6696 7341 7704
rect 7449 7990 7758 8031
rect 7449 7938 7488 7990
rect 7540 7938 7668 7990
rect 7720 7938 7758 7990
rect 7449 7851 7758 7938
rect 7449 7795 7486 7851
rect 7542 7795 7666 7851
rect 7722 7795 7758 7851
rect 7449 7516 7758 7795
rect 7449 7464 7488 7516
rect 7540 7464 7668 7516
rect 7720 7464 7758 7516
rect 7449 7423 7758 7464
rect 7866 7226 8461 8072
rect 7866 7174 7927 7226
rect 7979 7174 8138 7226
rect 8190 7174 8349 7226
rect 8401 7174 8461 7226
rect 6461 6644 6558 6696
rect 6610 6644 6769 6696
rect 6821 6644 6981 6696
rect 7033 6644 7192 6696
rect 7244 6644 7341 6696
rect 4728 6412 4929 6464
rect 4981 6412 5140 6464
rect 5192 6412 5351 6464
rect 5403 6412 5562 6464
rect 5614 6412 5773 6464
rect 5825 6412 6012 6464
rect 4728 6188 6012 6412
rect 4728 6136 4929 6188
rect 4981 6136 5140 6188
rect 5192 6136 5351 6188
rect 5403 6136 5562 6188
rect 5614 6136 5773 6188
rect 5825 6136 6012 6188
rect 4728 5728 6012 6136
rect 4728 5676 4929 5728
rect 4981 5676 5140 5728
rect 5192 5676 5351 5728
rect 5403 5676 5562 5728
rect 5614 5676 5773 5728
rect 5825 5676 6012 5728
rect 6237 5963 6366 6004
rect 6237 5911 6275 5963
rect 6327 5911 6366 5963
rect 6237 5820 6366 5911
rect 6237 5764 6273 5820
rect 6329 5787 6366 5820
rect 6461 5956 7341 6644
rect 7449 6936 7758 6977
rect 7449 6884 7488 6936
rect 7540 6884 7668 6936
rect 7720 6884 7758 6936
rect 7449 6605 7758 6884
rect 7449 6549 7486 6605
rect 7542 6549 7666 6605
rect 7722 6549 7758 6605
rect 7449 6462 7758 6549
rect 7449 6410 7488 6462
rect 7540 6410 7668 6462
rect 7720 6410 7758 6462
rect 7449 6369 7758 6410
rect 7866 6328 8461 7174
rect 7866 6272 7925 6328
rect 7981 6272 8136 6328
rect 8192 6272 8347 6328
rect 8403 6272 8461 6328
rect 6461 5904 6558 5956
rect 6610 5904 6769 5956
rect 6821 5904 6981 5956
rect 7033 5904 7192 5956
rect 7244 5904 7341 5956
rect 6329 5764 6365 5787
rect 6237 5725 6365 5764
rect 4728 5428 6012 5676
rect 4728 5372 4815 5428
rect 4871 5372 5025 5428
rect 5081 5372 5236 5428
rect 5292 5372 5448 5428
rect 5504 5372 5659 5428
rect 5715 5372 5869 5428
rect 5925 5372 6012 5428
rect 4728 5124 6012 5372
rect 4728 5072 4929 5124
rect 4981 5072 5140 5124
rect 5192 5072 5351 5124
rect 5403 5072 5562 5124
rect 5614 5072 5773 5124
rect 5825 5072 6012 5124
rect 4728 4664 6012 5072
rect 6237 5036 6365 5075
rect 6237 4980 6273 5036
rect 6329 5013 6365 5036
rect 6329 4980 6366 5013
rect 6237 4889 6366 4980
rect 6237 4837 6275 4889
rect 6327 4837 6366 4889
rect 6237 4796 6366 4837
rect 6461 4896 7341 5904
rect 7449 6190 7758 6231
rect 7449 6138 7488 6190
rect 7540 6138 7668 6190
rect 7720 6138 7758 6190
rect 7449 6051 7758 6138
rect 7449 5995 7486 6051
rect 7542 5995 7666 6051
rect 7722 5995 7758 6051
rect 7449 5716 7758 5995
rect 7449 5664 7488 5716
rect 7540 5664 7668 5716
rect 7720 5664 7758 5716
rect 7449 5623 7758 5664
rect 7866 5426 8461 6272
rect 7866 5374 7927 5426
rect 7979 5374 8138 5426
rect 8190 5374 8349 5426
rect 8401 5374 8461 5426
rect 6461 4844 6558 4896
rect 6610 4844 6769 4896
rect 6821 4844 6981 4896
rect 7033 4844 7192 4896
rect 7244 4844 7341 4896
rect 4728 4612 4929 4664
rect 4981 4612 5140 4664
rect 5192 4612 5351 4664
rect 5403 4612 5562 4664
rect 5614 4612 5773 4664
rect 5825 4612 6012 4664
rect 4728 4388 6012 4612
rect 4728 4336 4929 4388
rect 4981 4336 5140 4388
rect 5192 4336 5351 4388
rect 5403 4336 5562 4388
rect 5614 4336 5773 4388
rect 5825 4336 6012 4388
rect 4728 3928 6012 4336
rect 4728 3876 4929 3928
rect 4981 3876 5140 3928
rect 5192 3876 5351 3928
rect 5403 3876 5562 3928
rect 5614 3876 5773 3928
rect 5825 3876 6012 3928
rect 6237 4163 6366 4204
rect 6237 4111 6275 4163
rect 6327 4111 6366 4163
rect 6237 4020 6366 4111
rect 6237 3964 6273 4020
rect 6329 3987 6366 4020
rect 6461 4156 7341 4844
rect 7449 5136 7758 5177
rect 7449 5084 7488 5136
rect 7540 5084 7668 5136
rect 7720 5084 7758 5136
rect 7449 4805 7758 5084
rect 7449 4749 7486 4805
rect 7542 4749 7666 4805
rect 7722 4749 7758 4805
rect 7449 4662 7758 4749
rect 7449 4610 7488 4662
rect 7540 4610 7668 4662
rect 7720 4610 7758 4662
rect 7449 4569 7758 4610
rect 7866 4528 8461 5374
rect 7866 4472 7925 4528
rect 7981 4472 8136 4528
rect 8192 4472 8347 4528
rect 8403 4472 8461 4528
rect 6461 4104 6558 4156
rect 6610 4104 6769 4156
rect 6821 4104 6981 4156
rect 7033 4104 7192 4156
rect 7244 4104 7341 4156
rect 6329 3964 6365 3987
rect 6237 3925 6365 3964
rect 4728 3628 6012 3876
rect 4728 3572 4815 3628
rect 4871 3572 5025 3628
rect 5081 3572 5236 3628
rect 5292 3572 5448 3628
rect 5504 3572 5659 3628
rect 5715 3572 5869 3628
rect 5925 3572 6012 3628
rect 4728 3324 6012 3572
rect 4728 3272 4929 3324
rect 4981 3272 5140 3324
rect 5192 3272 5351 3324
rect 5403 3272 5562 3324
rect 5614 3272 5773 3324
rect 5825 3272 6012 3324
rect 4728 2864 6012 3272
rect 6237 3236 6365 3275
rect 6237 3180 6273 3236
rect 6329 3213 6365 3236
rect 6329 3180 6366 3213
rect 6237 3089 6366 3180
rect 6237 3037 6275 3089
rect 6327 3037 6366 3089
rect 6237 2996 6366 3037
rect 6461 3096 7341 4104
rect 7449 4390 7758 4431
rect 7449 4338 7488 4390
rect 7540 4338 7668 4390
rect 7720 4338 7758 4390
rect 7449 4251 7758 4338
rect 7449 4195 7486 4251
rect 7542 4195 7666 4251
rect 7722 4195 7758 4251
rect 7449 3916 7758 4195
rect 7449 3864 7488 3916
rect 7540 3864 7668 3916
rect 7720 3864 7758 3916
rect 7449 3823 7758 3864
rect 7866 3626 8461 4472
rect 7866 3574 7927 3626
rect 7979 3574 8138 3626
rect 8190 3574 8349 3626
rect 8401 3574 8461 3626
rect 6461 3044 6558 3096
rect 6610 3044 6769 3096
rect 6821 3044 6981 3096
rect 7033 3044 7192 3096
rect 7244 3044 7341 3096
rect 4728 2812 4929 2864
rect 4981 2812 5140 2864
rect 5192 2812 5351 2864
rect 5403 2812 5562 2864
rect 5614 2812 5773 2864
rect 5825 2812 6012 2864
rect 4728 2588 6012 2812
rect 4728 2536 4929 2588
rect 4981 2536 5140 2588
rect 5192 2536 5351 2588
rect 5403 2536 5562 2588
rect 5614 2536 5773 2588
rect 5825 2536 6012 2588
rect 4728 2128 6012 2536
rect 4728 2076 4929 2128
rect 4981 2076 5140 2128
rect 5192 2076 5351 2128
rect 5403 2076 5562 2128
rect 5614 2076 5773 2128
rect 5825 2076 6012 2128
rect 6237 2363 6366 2404
rect 6237 2311 6275 2363
rect 6327 2311 6366 2363
rect 6237 2220 6366 2311
rect 6237 2164 6273 2220
rect 6329 2187 6366 2220
rect 6461 2356 7341 3044
rect 7449 3336 7758 3377
rect 7449 3284 7488 3336
rect 7540 3284 7668 3336
rect 7720 3284 7758 3336
rect 7449 3005 7758 3284
rect 7449 2949 7486 3005
rect 7542 2949 7666 3005
rect 7722 2949 7758 3005
rect 7449 2862 7758 2949
rect 7449 2810 7488 2862
rect 7540 2810 7668 2862
rect 7720 2810 7758 2862
rect 7449 2769 7758 2810
rect 7866 2728 8461 3574
rect 7866 2672 7925 2728
rect 7981 2672 8136 2728
rect 8192 2672 8347 2728
rect 8403 2672 8461 2728
rect 6461 2304 6558 2356
rect 6610 2304 6769 2356
rect 6821 2304 6981 2356
rect 7033 2304 7192 2356
rect 7244 2304 7341 2356
rect 6329 2164 6365 2187
rect 6237 2125 6365 2164
rect 4728 1828 6012 2076
rect 4728 1772 4815 1828
rect 4871 1772 5025 1828
rect 5081 1772 5236 1828
rect 5292 1772 5448 1828
rect 5504 1772 5659 1828
rect 5715 1772 5869 1828
rect 5925 1772 6012 1828
rect 4728 1524 6012 1772
rect 4728 1472 4929 1524
rect 4981 1472 5140 1524
rect 5192 1472 5351 1524
rect 5403 1472 5562 1524
rect 5614 1472 5773 1524
rect 5825 1472 6012 1524
rect 4728 1064 6012 1472
rect 6237 1436 6365 1475
rect 6237 1380 6273 1436
rect 6329 1413 6365 1436
rect 6329 1380 6366 1413
rect 6237 1289 6366 1380
rect 6237 1237 6275 1289
rect 6327 1237 6366 1289
rect 6237 1196 6366 1237
rect 6461 1296 7341 2304
rect 7449 2590 7758 2631
rect 7449 2538 7488 2590
rect 7540 2538 7668 2590
rect 7720 2538 7758 2590
rect 7449 2451 7758 2538
rect 7449 2395 7486 2451
rect 7542 2395 7666 2451
rect 7722 2395 7758 2451
rect 7449 2116 7758 2395
rect 7449 2064 7488 2116
rect 7540 2064 7668 2116
rect 7720 2064 7758 2116
rect 7449 2023 7758 2064
rect 7866 1826 8461 2672
rect 7866 1774 7927 1826
rect 7979 1774 8138 1826
rect 8190 1774 8349 1826
rect 8401 1774 8461 1826
rect 6461 1244 6558 1296
rect 6610 1244 6769 1296
rect 6821 1244 6981 1296
rect 7033 1244 7192 1296
rect 7244 1244 7341 1296
rect 4728 1012 4929 1064
rect 4981 1012 5140 1064
rect 5192 1012 5351 1064
rect 5403 1012 5562 1064
rect 5614 1012 5773 1064
rect 5825 1012 6012 1064
rect 4728 788 6012 1012
rect 4728 736 4929 788
rect 4981 736 5140 788
rect 5192 736 5351 788
rect 5403 736 5562 788
rect 5614 736 5773 788
rect 5825 736 6012 788
rect 4728 328 6012 736
rect 4728 276 4929 328
rect 4981 276 5140 328
rect 5192 276 5351 328
rect 5403 276 5562 328
rect 5614 276 5773 328
rect 5825 276 6012 328
rect 6237 563 6366 604
rect 6237 511 6275 563
rect 6327 511 6366 563
rect 6237 420 6366 511
rect 6237 364 6273 420
rect 6329 387 6366 420
rect 6461 556 7341 1244
rect 7449 1536 7758 1577
rect 7449 1484 7488 1536
rect 7540 1484 7668 1536
rect 7720 1484 7758 1536
rect 7449 1205 7758 1484
rect 7449 1149 7486 1205
rect 7542 1149 7666 1205
rect 7722 1149 7758 1205
rect 7449 1062 7758 1149
rect 7449 1010 7488 1062
rect 7540 1010 7668 1062
rect 7720 1010 7758 1062
rect 7449 969 7758 1010
rect 7866 928 8461 1774
rect 7866 872 7925 928
rect 7981 872 8136 928
rect 8192 872 8347 928
rect 8403 872 8461 928
rect 6461 504 6558 556
rect 6610 504 6769 556
rect 6821 504 6981 556
rect 7033 504 7192 556
rect 7244 504 7341 556
rect 6329 364 6365 387
rect 6237 325 6365 364
rect 4728 28 6012 276
rect 4728 -28 4815 28
rect 4871 -28 5025 28
rect 5081 -28 5236 28
rect 5292 -28 5448 28
rect 5504 -28 5659 28
rect 5715 -28 5869 28
rect 5925 -28 6012 28
rect 4728 -151 6012 -28
rect 6461 -151 7341 504
rect 7449 790 7758 831
rect 7449 738 7488 790
rect 7540 738 7668 790
rect 7720 738 7758 790
rect 7449 651 7758 738
rect 7449 595 7486 651
rect 7542 595 7666 651
rect 7722 595 7758 651
rect 7449 316 7758 595
rect 7449 264 7488 316
rect 7540 264 7668 316
rect 7720 264 7758 316
rect 7449 223 7758 264
rect 7866 26 8461 872
rect 7866 -26 7927 26
rect 7979 -26 8138 26
rect 8190 -26 8349 26
rect 8401 -26 8461 26
rect 7866 -151 8461 -26
rect 8564 14428 9216 14551
rect 8564 14372 8647 14428
rect 8703 14372 8827 14428
rect 8883 14372 9216 14428
rect 8564 12628 9216 14372
rect 9812 14426 10121 14551
rect 9812 14374 9850 14426
rect 9902 14374 10030 14426
rect 10082 14374 10121 14426
rect 9333 14188 9462 14229
rect 9333 14136 9372 14188
rect 9424 14136 9462 14188
rect 9333 13805 9462 14136
rect 9333 13749 9370 13805
rect 9426 13749 9462 13805
rect 9333 13710 9462 13749
rect 9553 14036 9681 14075
rect 9553 13980 9589 14036
rect 9645 14014 9681 14036
rect 9645 13980 9682 14014
rect 9553 13973 9682 13980
rect 9553 13921 9591 13973
rect 9643 13921 9682 13973
rect 9553 13787 9682 13921
rect 9553 13735 9591 13787
rect 9643 13735 9682 13787
rect 9553 13694 9682 13735
rect 9812 13528 10121 14374
rect 9812 13472 9848 13528
rect 9904 13472 10028 13528
rect 10084 13472 10121 13528
rect 9333 13251 9462 13290
rect 9333 13195 9370 13251
rect 9426 13195 9462 13251
rect 9333 12864 9462 13195
rect 9553 13265 9682 13306
rect 9553 13213 9591 13265
rect 9643 13213 9682 13265
rect 9553 13079 9682 13213
rect 9553 13027 9591 13079
rect 9643 13027 9682 13079
rect 9553 13020 9682 13027
rect 9553 12964 9589 13020
rect 9645 12986 9682 13020
rect 9645 12964 9681 12986
rect 9553 12925 9681 12964
rect 9333 12812 9372 12864
rect 9424 12812 9462 12864
rect 9333 12771 9462 12812
rect 8564 12572 8647 12628
rect 8703 12572 8827 12628
rect 8883 12572 9216 12628
rect 8564 10828 9216 12572
rect 9812 12626 10121 13472
rect 9812 12574 9850 12626
rect 9902 12574 10030 12626
rect 10082 12574 10121 12626
rect 9333 12388 9462 12429
rect 9333 12336 9372 12388
rect 9424 12336 9462 12388
rect 9333 12005 9462 12336
rect 9333 11949 9370 12005
rect 9426 11949 9462 12005
rect 9333 11910 9462 11949
rect 9553 12236 9681 12275
rect 9553 12180 9589 12236
rect 9645 12214 9681 12236
rect 9645 12180 9682 12214
rect 9553 12173 9682 12180
rect 9553 12121 9591 12173
rect 9643 12121 9682 12173
rect 9553 11987 9682 12121
rect 9553 11935 9591 11987
rect 9643 11935 9682 11987
rect 9553 11894 9682 11935
rect 9812 11728 10121 12574
rect 9812 11672 9848 11728
rect 9904 11672 10028 11728
rect 10084 11672 10121 11728
rect 9333 11451 9462 11490
rect 9333 11395 9370 11451
rect 9426 11395 9462 11451
rect 9333 11064 9462 11395
rect 9553 11465 9682 11506
rect 9553 11413 9591 11465
rect 9643 11413 9682 11465
rect 9553 11279 9682 11413
rect 9553 11227 9591 11279
rect 9643 11227 9682 11279
rect 9553 11220 9682 11227
rect 9553 11164 9589 11220
rect 9645 11186 9682 11220
rect 9645 11164 9681 11186
rect 9553 11125 9681 11164
rect 9333 11012 9372 11064
rect 9424 11012 9462 11064
rect 9333 10971 9462 11012
rect 8564 10772 8647 10828
rect 8703 10772 8827 10828
rect 8883 10772 9216 10828
rect 8564 9028 9216 10772
rect 9812 10826 10121 11672
rect 9812 10774 9850 10826
rect 9902 10774 10030 10826
rect 10082 10774 10121 10826
rect 9333 10588 9462 10629
rect 9333 10536 9372 10588
rect 9424 10536 9462 10588
rect 9333 10205 9462 10536
rect 9333 10149 9370 10205
rect 9426 10149 9462 10205
rect 9333 10110 9462 10149
rect 9553 10436 9681 10475
rect 9553 10380 9589 10436
rect 9645 10414 9681 10436
rect 9645 10380 9682 10414
rect 9553 10373 9682 10380
rect 9553 10321 9591 10373
rect 9643 10321 9682 10373
rect 9553 10187 9682 10321
rect 9553 10135 9591 10187
rect 9643 10135 9682 10187
rect 9553 10094 9682 10135
rect 9812 9928 10121 10774
rect 9812 9872 9848 9928
rect 9904 9872 10028 9928
rect 10084 9872 10121 9928
rect 9333 9651 9462 9690
rect 9333 9595 9370 9651
rect 9426 9595 9462 9651
rect 9333 9264 9462 9595
rect 9553 9665 9682 9706
rect 9553 9613 9591 9665
rect 9643 9613 9682 9665
rect 9553 9479 9682 9613
rect 9553 9427 9591 9479
rect 9643 9427 9682 9479
rect 9553 9420 9682 9427
rect 9553 9364 9589 9420
rect 9645 9386 9682 9420
rect 9645 9364 9681 9386
rect 9553 9325 9681 9364
rect 9333 9212 9372 9264
rect 9424 9212 9462 9264
rect 9333 9171 9462 9212
rect 8564 8972 8647 9028
rect 8703 8972 8827 9028
rect 8883 8972 9216 9028
rect 8564 7228 9216 8972
rect 9812 9026 10121 9872
rect 9812 8974 9850 9026
rect 9902 8974 10030 9026
rect 10082 8974 10121 9026
rect 9333 8788 9462 8829
rect 9333 8736 9372 8788
rect 9424 8736 9462 8788
rect 9333 8405 9462 8736
rect 9333 8349 9370 8405
rect 9426 8349 9462 8405
rect 9333 8310 9462 8349
rect 9553 8636 9681 8675
rect 9553 8580 9589 8636
rect 9645 8614 9681 8636
rect 9645 8580 9682 8614
rect 9553 8573 9682 8580
rect 9553 8521 9591 8573
rect 9643 8521 9682 8573
rect 9553 8387 9682 8521
rect 9553 8335 9591 8387
rect 9643 8335 9682 8387
rect 9553 8294 9682 8335
rect 9812 8128 10121 8974
rect 9812 8072 9848 8128
rect 9904 8072 10028 8128
rect 10084 8072 10121 8128
rect 9333 7851 9462 7890
rect 9333 7795 9370 7851
rect 9426 7795 9462 7851
rect 9333 7464 9462 7795
rect 9553 7865 9682 7906
rect 9553 7813 9591 7865
rect 9643 7813 9682 7865
rect 9553 7679 9682 7813
rect 9553 7627 9591 7679
rect 9643 7627 9682 7679
rect 9553 7620 9682 7627
rect 9553 7564 9589 7620
rect 9645 7586 9682 7620
rect 9645 7564 9681 7586
rect 9553 7525 9681 7564
rect 9333 7412 9372 7464
rect 9424 7412 9462 7464
rect 9333 7371 9462 7412
rect 8564 7172 8647 7228
rect 8703 7172 8827 7228
rect 8883 7172 9216 7228
rect 8564 5428 9216 7172
rect 9812 7226 10121 8072
rect 9812 7174 9850 7226
rect 9902 7174 10030 7226
rect 10082 7174 10121 7226
rect 9333 6988 9462 7029
rect 9333 6936 9372 6988
rect 9424 6936 9462 6988
rect 9333 6605 9462 6936
rect 9333 6549 9370 6605
rect 9426 6549 9462 6605
rect 9333 6510 9462 6549
rect 9553 6836 9681 6875
rect 9553 6780 9589 6836
rect 9645 6814 9681 6836
rect 9645 6780 9682 6814
rect 9553 6773 9682 6780
rect 9553 6721 9591 6773
rect 9643 6721 9682 6773
rect 9553 6587 9682 6721
rect 9553 6535 9591 6587
rect 9643 6535 9682 6587
rect 9553 6494 9682 6535
rect 9812 6328 10121 7174
rect 9812 6272 9848 6328
rect 9904 6272 10028 6328
rect 10084 6272 10121 6328
rect 9333 6051 9462 6090
rect 9333 5995 9370 6051
rect 9426 5995 9462 6051
rect 9333 5664 9462 5995
rect 9553 6065 9682 6106
rect 9553 6013 9591 6065
rect 9643 6013 9682 6065
rect 9553 5879 9682 6013
rect 9553 5827 9591 5879
rect 9643 5827 9682 5879
rect 9553 5820 9682 5827
rect 9553 5764 9589 5820
rect 9645 5786 9682 5820
rect 9645 5764 9681 5786
rect 9553 5725 9681 5764
rect 9333 5612 9372 5664
rect 9424 5612 9462 5664
rect 9333 5571 9462 5612
rect 8564 5372 8647 5428
rect 8703 5372 8827 5428
rect 8883 5372 9216 5428
rect 8564 3628 9216 5372
rect 9812 5426 10121 6272
rect 9812 5374 9850 5426
rect 9902 5374 10030 5426
rect 10082 5374 10121 5426
rect 9333 5188 9462 5229
rect 9333 5136 9372 5188
rect 9424 5136 9462 5188
rect 9333 4805 9462 5136
rect 9333 4749 9370 4805
rect 9426 4749 9462 4805
rect 9333 4710 9462 4749
rect 9553 5036 9681 5075
rect 9553 4980 9589 5036
rect 9645 5014 9681 5036
rect 9645 4980 9682 5014
rect 9553 4973 9682 4980
rect 9553 4921 9591 4973
rect 9643 4921 9682 4973
rect 9553 4787 9682 4921
rect 9553 4735 9591 4787
rect 9643 4735 9682 4787
rect 9553 4694 9682 4735
rect 9812 4528 10121 5374
rect 9812 4472 9848 4528
rect 9904 4472 10028 4528
rect 10084 4472 10121 4528
rect 9333 4251 9462 4290
rect 9333 4195 9370 4251
rect 9426 4195 9462 4251
rect 9333 3864 9462 4195
rect 9553 4265 9682 4306
rect 9553 4213 9591 4265
rect 9643 4213 9682 4265
rect 9553 4079 9682 4213
rect 9553 4027 9591 4079
rect 9643 4027 9682 4079
rect 9553 4020 9682 4027
rect 9553 3964 9589 4020
rect 9645 3986 9682 4020
rect 9645 3964 9681 3986
rect 9553 3925 9681 3964
rect 9333 3812 9372 3864
rect 9424 3812 9462 3864
rect 9333 3771 9462 3812
rect 8564 3572 8647 3628
rect 8703 3572 8827 3628
rect 8883 3572 9216 3628
rect 8564 1828 9216 3572
rect 9812 3626 10121 4472
rect 9812 3574 9850 3626
rect 9902 3574 10030 3626
rect 10082 3574 10121 3626
rect 9333 3388 9462 3429
rect 9333 3336 9372 3388
rect 9424 3336 9462 3388
rect 9333 3005 9462 3336
rect 9333 2949 9370 3005
rect 9426 2949 9462 3005
rect 9333 2910 9462 2949
rect 9553 3236 9681 3275
rect 9553 3180 9589 3236
rect 9645 3214 9681 3236
rect 9645 3180 9682 3214
rect 9553 3173 9682 3180
rect 9553 3121 9591 3173
rect 9643 3121 9682 3173
rect 9553 2987 9682 3121
rect 9553 2935 9591 2987
rect 9643 2935 9682 2987
rect 9553 2894 9682 2935
rect 9812 2728 10121 3574
rect 9812 2672 9848 2728
rect 9904 2672 10028 2728
rect 10084 2672 10121 2728
rect 9333 2451 9462 2490
rect 9333 2395 9370 2451
rect 9426 2395 9462 2451
rect 9333 2064 9462 2395
rect 9553 2465 9682 2506
rect 9553 2413 9591 2465
rect 9643 2413 9682 2465
rect 9553 2279 9682 2413
rect 9553 2227 9591 2279
rect 9643 2227 9682 2279
rect 9553 2220 9682 2227
rect 9553 2164 9589 2220
rect 9645 2186 9682 2220
rect 9645 2164 9681 2186
rect 9553 2125 9681 2164
rect 9333 2012 9372 2064
rect 9424 2012 9462 2064
rect 9333 1971 9462 2012
rect 8564 1772 8647 1828
rect 8703 1772 8827 1828
rect 8883 1772 9216 1828
rect 8564 28 9216 1772
rect 9812 1826 10121 2672
rect 9812 1774 9850 1826
rect 9902 1774 10030 1826
rect 10082 1774 10121 1826
rect 9333 1588 9462 1629
rect 9333 1536 9372 1588
rect 9424 1536 9462 1588
rect 9333 1205 9462 1536
rect 9333 1149 9370 1205
rect 9426 1149 9462 1205
rect 9333 1110 9462 1149
rect 9553 1436 9681 1475
rect 9553 1380 9589 1436
rect 9645 1414 9681 1436
rect 9645 1380 9682 1414
rect 9553 1373 9682 1380
rect 9553 1321 9591 1373
rect 9643 1321 9682 1373
rect 9553 1187 9682 1321
rect 9553 1135 9591 1187
rect 9643 1135 9682 1187
rect 9553 1094 9682 1135
rect 9812 928 10121 1774
rect 9812 872 9848 928
rect 9904 872 10028 928
rect 10084 872 10121 928
rect 9333 651 9462 690
rect 9333 595 9370 651
rect 9426 595 9462 651
rect 9333 264 9462 595
rect 9553 665 9682 706
rect 9553 613 9591 665
rect 9643 613 9682 665
rect 9553 479 9682 613
rect 9553 427 9591 479
rect 9643 427 9682 479
rect 9553 420 9682 427
rect 9553 364 9589 420
rect 9645 386 9682 420
rect 9645 364 9681 386
rect 9553 325 9681 364
rect 9333 212 9372 264
rect 9424 212 9462 264
rect 9333 171 9462 212
rect 8564 -28 8647 28
rect 8703 -28 8827 28
rect 8883 -28 9216 28
rect 8564 -151 9216 -28
rect 9812 26 10121 872
rect 9812 -26 9850 26
rect 9902 -26 10030 26
rect 10082 -26 10121 26
rect 9812 -151 10121 -26
rect 10315 -151 10536 14551
rect 10692 -151 10914 14551
rect 11070 -164 11292 14564
rect 11448 14188 11669 14564
rect 11448 14136 11532 14188
rect 11584 14136 11669 14188
rect 11448 12864 11669 14136
rect 11448 12812 11532 12864
rect 11584 12812 11669 12864
rect 11448 12388 11669 12812
rect 11448 12336 11532 12388
rect 11584 12336 11669 12388
rect 11448 11064 11669 12336
rect 11448 11012 11532 11064
rect 11584 11012 11669 11064
rect 11448 10588 11669 11012
rect 11448 10536 11532 10588
rect 11584 10536 11669 10588
rect 11448 9264 11669 10536
rect 11448 9212 11532 9264
rect 11584 9212 11669 9264
rect 11448 8788 11669 9212
rect 11448 8736 11532 8788
rect 11584 8736 11669 8788
rect 11448 7464 11669 8736
rect 11448 7412 11532 7464
rect 11584 7412 11669 7464
rect 11448 6988 11669 7412
rect 11448 6936 11532 6988
rect 11584 6936 11669 6988
rect 11448 5664 11669 6936
rect 11448 5612 11532 5664
rect 11584 5612 11669 5664
rect 11448 5188 11669 5612
rect 11448 5136 11532 5188
rect 11584 5136 11669 5188
rect 11448 3864 11669 5136
rect 11448 3812 11532 3864
rect 11584 3812 11669 3864
rect 11448 3388 11669 3812
rect 11448 3336 11532 3388
rect 11584 3336 11669 3388
rect 11448 2064 11669 3336
rect 11448 2012 11532 2064
rect 11584 2012 11669 2064
rect 11448 1588 11669 2012
rect 11448 1536 11532 1588
rect 11584 1536 11669 1588
rect 11448 264 11669 1536
rect 11448 212 11532 264
rect 11584 212 11669 264
rect 11448 -164 11669 212
rect 11826 -164 12047 14564
rect 12203 -164 12425 14564
rect 12581 13957 12802 14564
rect 12581 13905 12665 13957
rect 12717 13905 12802 13957
rect 12581 13095 12802 13905
rect 12581 13043 12665 13095
rect 12717 13043 12802 13095
rect 12581 12157 12802 13043
rect 12581 12105 12665 12157
rect 12717 12105 12802 12157
rect 12581 11295 12802 12105
rect 12581 11243 12665 11295
rect 12717 11243 12802 11295
rect 12581 10357 12802 11243
rect 12581 10305 12665 10357
rect 12717 10305 12802 10357
rect 12581 9495 12802 10305
rect 12581 9443 12665 9495
rect 12717 9443 12802 9495
rect 12581 8557 12802 9443
rect 12581 8505 12665 8557
rect 12717 8505 12802 8557
rect 12581 7695 12802 8505
rect 12581 7643 12665 7695
rect 12717 7643 12802 7695
rect 12581 -164 12802 7643
rect 12959 6757 13180 14564
rect 12959 6705 13042 6757
rect 13094 6705 13180 6757
rect 12959 5895 13180 6705
rect 12959 5843 13042 5895
rect 13094 5843 13180 5895
rect 12959 4957 13180 5843
rect 12959 4905 13042 4957
rect 13094 4905 13180 4957
rect 12959 4095 13180 4905
rect 12959 4043 13042 4095
rect 13094 4043 13180 4095
rect 12959 3157 13180 4043
rect 12959 3105 13042 3157
rect 13094 3105 13180 3157
rect 12959 2295 13180 3105
rect 12959 2243 13042 2295
rect 13094 2243 13180 2295
rect 12959 1357 13180 2243
rect 12959 1305 13042 1357
rect 13094 1305 13180 1357
rect 12959 495 13180 1305
rect 12959 443 13042 495
rect 13094 443 13180 495
rect 12959 -164 13180 443
rect 13301 14426 14160 14551
rect 13301 14374 13387 14426
rect 13439 14374 13598 14426
rect 13650 14374 13810 14426
rect 13862 14374 14021 14426
rect 14073 14374 14160 14426
rect 13301 13528 14160 14374
rect 13301 13472 13385 13528
rect 13441 13472 13596 13528
rect 13652 13472 13808 13528
rect 13864 13472 14019 13528
rect 14075 13472 14160 13528
rect 13301 12626 14160 13472
rect 13301 12574 13387 12626
rect 13439 12574 13598 12626
rect 13650 12574 13810 12626
rect 13862 12574 14021 12626
rect 14073 12574 14160 12626
rect 13301 11728 14160 12574
rect 13301 11672 13385 11728
rect 13441 11672 13596 11728
rect 13652 11672 13808 11728
rect 13864 11672 14019 11728
rect 14075 11672 14160 11728
rect 13301 10826 14160 11672
rect 13301 10774 13387 10826
rect 13439 10774 13598 10826
rect 13650 10774 13810 10826
rect 13862 10774 14021 10826
rect 14073 10774 14160 10826
rect 13301 9928 14160 10774
rect 13301 9872 13385 9928
rect 13441 9872 13596 9928
rect 13652 9872 13808 9928
rect 13864 9872 14019 9928
rect 14075 9872 14160 9928
rect 13301 9026 14160 9872
rect 13301 8974 13387 9026
rect 13439 8974 13598 9026
rect 13650 8974 13810 9026
rect 13862 8974 14021 9026
rect 14073 8974 14160 9026
rect 13301 8128 14160 8974
rect 13301 8072 13385 8128
rect 13441 8072 13596 8128
rect 13652 8072 13808 8128
rect 13864 8072 14019 8128
rect 14075 8072 14160 8128
rect 13301 7226 14160 8072
rect 13301 7174 13387 7226
rect 13439 7174 13598 7226
rect 13650 7174 13810 7226
rect 13862 7174 14021 7226
rect 14073 7174 14160 7226
rect 13301 6328 14160 7174
rect 13301 6272 13385 6328
rect 13441 6272 13596 6328
rect 13652 6272 13808 6328
rect 13864 6272 14019 6328
rect 14075 6272 14160 6328
rect 13301 5426 14160 6272
rect 13301 5374 13387 5426
rect 13439 5374 13598 5426
rect 13650 5374 13810 5426
rect 13862 5374 14021 5426
rect 14073 5374 14160 5426
rect 13301 4528 14160 5374
rect 13301 4472 13385 4528
rect 13441 4472 13596 4528
rect 13652 4472 13808 4528
rect 13864 4472 14019 4528
rect 14075 4472 14160 4528
rect 13301 3626 14160 4472
rect 13301 3574 13387 3626
rect 13439 3574 13598 3626
rect 13650 3574 13810 3626
rect 13862 3574 14021 3626
rect 14073 3574 14160 3626
rect 13301 2728 14160 3574
rect 13301 2672 13385 2728
rect 13441 2672 13596 2728
rect 13652 2672 13808 2728
rect 13864 2672 14019 2728
rect 14075 2672 14160 2728
rect 13301 1826 14160 2672
rect 13301 1774 13387 1826
rect 13439 1774 13598 1826
rect 13650 1774 13810 1826
rect 13862 1774 14021 1826
rect 14073 1774 14160 1826
rect 13301 928 14160 1774
rect 13301 872 13385 928
rect 13441 872 13596 928
rect 13652 872 13808 928
rect 13864 872 14019 928
rect 14075 872 14160 928
rect 13301 26 14160 872
rect 13301 -26 13387 26
rect 13439 -26 13598 26
rect 13650 -26 13810 26
rect 13862 -26 14021 26
rect 14073 -26 14160 26
rect 13301 -151 14160 -26
rect 14355 14428 14981 14551
rect 14355 14372 14429 14428
rect 14485 14372 14640 14428
rect 14696 14372 14851 14428
rect 14907 14372 14981 14428
rect 14355 13964 14981 14372
rect 14355 13912 14536 13964
rect 14588 13912 14748 13964
rect 14800 13912 14981 13964
rect 14355 13088 14981 13912
rect 14355 13036 14536 13088
rect 14588 13036 14748 13088
rect 14800 13036 14981 13088
rect 14355 12628 14981 13036
rect 14355 12572 14429 12628
rect 14485 12572 14640 12628
rect 14696 12572 14851 12628
rect 14907 12572 14981 12628
rect 14355 12164 14981 12572
rect 14355 12112 14536 12164
rect 14588 12112 14748 12164
rect 14800 12112 14981 12164
rect 14355 11288 14981 12112
rect 14355 11236 14536 11288
rect 14588 11236 14748 11288
rect 14800 11236 14981 11288
rect 14355 10828 14981 11236
rect 14355 10772 14429 10828
rect 14485 10772 14640 10828
rect 14696 10772 14851 10828
rect 14907 10772 14981 10828
rect 14355 10364 14981 10772
rect 14355 10312 14536 10364
rect 14588 10312 14748 10364
rect 14800 10312 14981 10364
rect 14355 9488 14981 10312
rect 14355 9436 14536 9488
rect 14588 9436 14748 9488
rect 14800 9436 14981 9488
rect 14355 9028 14981 9436
rect 14355 8972 14429 9028
rect 14485 8972 14640 9028
rect 14696 8972 14851 9028
rect 14907 8972 14981 9028
rect 14355 8564 14981 8972
rect 14355 8512 14536 8564
rect 14588 8512 14748 8564
rect 14800 8512 14981 8564
rect 14355 7688 14981 8512
rect 14355 7636 14536 7688
rect 14588 7636 14748 7688
rect 14800 7636 14981 7688
rect 14355 7228 14981 7636
rect 14355 7172 14429 7228
rect 14485 7172 14640 7228
rect 14696 7172 14851 7228
rect 14907 7172 14981 7228
rect 14355 6764 14981 7172
rect 14355 6712 14536 6764
rect 14588 6712 14748 6764
rect 14800 6712 14981 6764
rect 14355 5888 14981 6712
rect 14355 5836 14536 5888
rect 14588 5836 14748 5888
rect 14800 5836 14981 5888
rect 14355 5428 14981 5836
rect 14355 5372 14429 5428
rect 14485 5372 14640 5428
rect 14696 5372 14851 5428
rect 14907 5372 14981 5428
rect 14355 4964 14981 5372
rect 14355 4912 14536 4964
rect 14588 4912 14748 4964
rect 14800 4912 14981 4964
rect 14355 4088 14981 4912
rect 14355 4036 14536 4088
rect 14588 4036 14748 4088
rect 14800 4036 14981 4088
rect 14355 3628 14981 4036
rect 14355 3572 14429 3628
rect 14485 3572 14640 3628
rect 14696 3572 14851 3628
rect 14907 3572 14981 3628
rect 14355 3164 14981 3572
rect 14355 3112 14536 3164
rect 14588 3112 14748 3164
rect 14800 3112 14981 3164
rect 14355 2288 14981 3112
rect 14355 2236 14536 2288
rect 14588 2236 14748 2288
rect 14800 2236 14981 2288
rect 14355 1828 14981 2236
rect 14355 1772 14429 1828
rect 14485 1772 14640 1828
rect 14696 1772 14851 1828
rect 14907 1772 14981 1828
rect 14355 1364 14981 1772
rect 14355 1312 14536 1364
rect 14588 1312 14748 1364
rect 14800 1312 14981 1364
rect 14355 488 14981 1312
rect 14355 436 14536 488
rect 14588 436 14748 488
rect 14800 436 14981 488
rect 14355 28 14981 436
rect 14355 -28 14429 28
rect 14485 -28 14640 28
rect 14696 -28 14851 28
rect 14907 -28 14981 28
rect 14355 -151 14981 -28
rect 15111 13848 15332 14564
rect 15111 13796 15194 13848
rect 15246 13796 15332 13848
rect 15111 6648 15332 13796
rect 15111 6596 15194 6648
rect 15246 6596 15332 6648
rect 15111 -164 15332 6596
rect 15488 13204 15710 14564
rect 15488 13152 15572 13204
rect 15624 13152 15710 13204
rect 15488 6004 15710 13152
rect 15488 5952 15572 6004
rect 15624 5952 15710 6004
rect 15488 -164 15710 5952
rect 15866 12048 16088 14564
rect 15866 11996 15950 12048
rect 16002 11996 16088 12048
rect 15866 4848 16088 11996
rect 15866 4796 15950 4848
rect 16002 4796 16088 4848
rect 15866 -164 16088 4796
rect 16244 11404 16465 14564
rect 16244 11352 16328 11404
rect 16380 11352 16465 11404
rect 16244 4204 16465 11352
rect 16244 4152 16328 4204
rect 16380 4152 16465 4204
rect 16244 -164 16465 4152
rect 16622 10248 16843 14564
rect 16622 10196 16705 10248
rect 16757 10196 16843 10248
rect 16622 3048 16843 10196
rect 16622 2996 16705 3048
rect 16757 2996 16843 3048
rect 16622 -164 16843 2996
rect 16999 9604 17221 14564
rect 16999 9552 17083 9604
rect 17135 9552 17221 9604
rect 16999 2404 17221 9552
rect 16999 2352 17083 2404
rect 17135 2352 17221 2404
rect 16999 -164 17221 2352
rect 17377 8448 17599 14564
rect 17377 8396 17461 8448
rect 17513 8396 17599 8448
rect 17377 1248 17599 8396
rect 17377 1196 17461 1248
rect 17513 1196 17599 1248
rect 17377 -164 17599 1196
rect 17755 7804 17976 14564
rect 18387 14428 19588 14551
rect 18387 14372 18433 14428
rect 18489 14372 18643 14428
rect 18699 14372 18854 14428
rect 18910 14372 19066 14428
rect 19122 14372 19277 14428
rect 19333 14372 19487 14428
rect 19543 14372 19588 14428
rect 18387 14127 19588 14372
rect 18387 14075 18540 14127
rect 18592 14075 18751 14127
rect 18803 14075 18962 14127
rect 19014 14075 19173 14127
rect 19225 14075 19384 14127
rect 19436 14075 19588 14127
rect 18154 14022 18284 14061
rect 18154 13966 18191 14022
rect 18247 13966 18284 14022
rect 18154 13804 18284 13966
rect 18154 13748 18191 13804
rect 18247 13748 18284 13804
rect 18154 13710 18284 13748
rect 18387 13664 19588 14075
rect 18387 13612 18540 13664
rect 18592 13612 18751 13664
rect 18803 13612 18962 13664
rect 19014 13612 19173 13664
rect 19225 13612 19384 13664
rect 19436 13612 19588 13664
rect 18387 13388 19588 13612
rect 18387 13336 18540 13388
rect 18592 13336 18751 13388
rect 18803 13336 18962 13388
rect 19014 13336 19173 13388
rect 19225 13336 19384 13388
rect 19436 13336 19588 13388
rect 18154 13252 18284 13290
rect 18154 13196 18191 13252
rect 18247 13196 18284 13252
rect 18154 13034 18284 13196
rect 18154 12978 18191 13034
rect 18247 12978 18284 13034
rect 18154 12939 18284 12978
rect 18387 12925 19588 13336
rect 18387 12873 18540 12925
rect 18592 12873 18751 12925
rect 18803 12873 18962 12925
rect 19014 12873 19173 12925
rect 19225 12873 19384 12925
rect 19436 12873 19588 12925
rect 18387 12628 19588 12873
rect 18387 12572 18433 12628
rect 18489 12572 18643 12628
rect 18699 12572 18854 12628
rect 18910 12572 19066 12628
rect 19122 12572 19277 12628
rect 19333 12572 19487 12628
rect 19543 12572 19588 12628
rect 18387 12327 19588 12572
rect 18387 12275 18540 12327
rect 18592 12275 18751 12327
rect 18803 12275 18962 12327
rect 19014 12275 19173 12327
rect 19225 12275 19384 12327
rect 19436 12275 19588 12327
rect 18154 12222 18284 12261
rect 18154 12166 18191 12222
rect 18247 12166 18284 12222
rect 18154 12004 18284 12166
rect 18154 11948 18191 12004
rect 18247 11948 18284 12004
rect 18154 11910 18284 11948
rect 18387 11864 19588 12275
rect 18387 11812 18540 11864
rect 18592 11812 18751 11864
rect 18803 11812 18962 11864
rect 19014 11812 19173 11864
rect 19225 11812 19384 11864
rect 19436 11812 19588 11864
rect 18387 11588 19588 11812
rect 18387 11536 18540 11588
rect 18592 11536 18751 11588
rect 18803 11536 18962 11588
rect 19014 11536 19173 11588
rect 19225 11536 19384 11588
rect 19436 11536 19588 11588
rect 18154 11452 18284 11490
rect 18154 11396 18191 11452
rect 18247 11396 18284 11452
rect 18154 11234 18284 11396
rect 18154 11178 18191 11234
rect 18247 11178 18284 11234
rect 18154 11139 18284 11178
rect 18387 11125 19588 11536
rect 18387 11073 18540 11125
rect 18592 11073 18751 11125
rect 18803 11073 18962 11125
rect 19014 11073 19173 11125
rect 19225 11073 19384 11125
rect 19436 11073 19588 11125
rect 18387 10828 19588 11073
rect 18387 10772 18433 10828
rect 18489 10772 18643 10828
rect 18699 10772 18854 10828
rect 18910 10772 19066 10828
rect 19122 10772 19277 10828
rect 19333 10772 19487 10828
rect 19543 10772 19588 10828
rect 18387 10527 19588 10772
rect 18387 10475 18540 10527
rect 18592 10475 18751 10527
rect 18803 10475 18962 10527
rect 19014 10475 19173 10527
rect 19225 10475 19384 10527
rect 19436 10475 19588 10527
rect 18154 10422 18284 10461
rect 18154 10366 18191 10422
rect 18247 10366 18284 10422
rect 18154 10204 18284 10366
rect 18154 10148 18191 10204
rect 18247 10148 18284 10204
rect 18154 10110 18284 10148
rect 18387 10064 19588 10475
rect 18387 10012 18540 10064
rect 18592 10012 18751 10064
rect 18803 10012 18962 10064
rect 19014 10012 19173 10064
rect 19225 10012 19384 10064
rect 19436 10012 19588 10064
rect 18387 9788 19588 10012
rect 18387 9736 18540 9788
rect 18592 9736 18751 9788
rect 18803 9736 18962 9788
rect 19014 9736 19173 9788
rect 19225 9736 19384 9788
rect 19436 9736 19588 9788
rect 18154 9652 18284 9690
rect 18154 9596 18191 9652
rect 18247 9596 18284 9652
rect 18154 9434 18284 9596
rect 18154 9378 18191 9434
rect 18247 9378 18284 9434
rect 18154 9339 18284 9378
rect 18387 9325 19588 9736
rect 18387 9273 18540 9325
rect 18592 9273 18751 9325
rect 18803 9273 18962 9325
rect 19014 9273 19173 9325
rect 19225 9273 19384 9325
rect 19436 9273 19588 9325
rect 18387 9028 19588 9273
rect 18387 8972 18433 9028
rect 18489 8972 18643 9028
rect 18699 8972 18854 9028
rect 18910 8972 19066 9028
rect 19122 8972 19277 9028
rect 19333 8972 19487 9028
rect 19543 8972 19588 9028
rect 18387 8727 19588 8972
rect 18387 8675 18540 8727
rect 18592 8675 18751 8727
rect 18803 8675 18962 8727
rect 19014 8675 19173 8727
rect 19225 8675 19384 8727
rect 19436 8675 19588 8727
rect 18154 8622 18284 8661
rect 18154 8566 18191 8622
rect 18247 8566 18284 8622
rect 18154 8404 18284 8566
rect 18154 8348 18191 8404
rect 18247 8348 18284 8404
rect 18154 8310 18284 8348
rect 18387 8264 19588 8675
rect 18387 8212 18540 8264
rect 18592 8212 18751 8264
rect 18803 8212 18962 8264
rect 19014 8212 19173 8264
rect 19225 8212 19384 8264
rect 19436 8212 19588 8264
rect 18387 7988 19588 8212
rect 18387 7936 18540 7988
rect 18592 7936 18751 7988
rect 18803 7936 18962 7988
rect 19014 7936 19173 7988
rect 19225 7936 19384 7988
rect 19436 7936 19588 7988
rect 17755 7752 17838 7804
rect 17890 7752 17976 7804
rect 17755 604 17976 7752
rect 18154 7852 18284 7890
rect 18154 7796 18191 7852
rect 18247 7796 18284 7852
rect 18154 7634 18284 7796
rect 18154 7578 18191 7634
rect 18247 7578 18284 7634
rect 18154 7539 18284 7578
rect 18387 7525 19588 7936
rect 18387 7473 18540 7525
rect 18592 7473 18751 7525
rect 18803 7473 18962 7525
rect 19014 7473 19173 7525
rect 19225 7473 19384 7525
rect 19436 7473 19588 7525
rect 18387 7228 19588 7473
rect 18387 7172 18433 7228
rect 18489 7172 18643 7228
rect 18699 7172 18854 7228
rect 18910 7172 19066 7228
rect 19122 7172 19277 7228
rect 19333 7172 19487 7228
rect 19543 7172 19588 7228
rect 18387 6927 19588 7172
rect 18387 6875 18540 6927
rect 18592 6875 18751 6927
rect 18803 6875 18962 6927
rect 19014 6875 19173 6927
rect 19225 6875 19384 6927
rect 19436 6875 19588 6927
rect 18154 6822 18284 6861
rect 18154 6766 18191 6822
rect 18247 6766 18284 6822
rect 18154 6604 18284 6766
rect 18154 6548 18191 6604
rect 18247 6548 18284 6604
rect 18154 6510 18284 6548
rect 18387 6464 19588 6875
rect 18387 6412 18540 6464
rect 18592 6412 18751 6464
rect 18803 6412 18962 6464
rect 19014 6412 19173 6464
rect 19225 6412 19384 6464
rect 19436 6412 19588 6464
rect 18387 6188 19588 6412
rect 18387 6136 18540 6188
rect 18592 6136 18751 6188
rect 18803 6136 18962 6188
rect 19014 6136 19173 6188
rect 19225 6136 19384 6188
rect 19436 6136 19588 6188
rect 18154 6052 18284 6090
rect 18154 5996 18191 6052
rect 18247 5996 18284 6052
rect 18154 5834 18284 5996
rect 18154 5778 18191 5834
rect 18247 5778 18284 5834
rect 18154 5739 18284 5778
rect 18387 5725 19588 6136
rect 18387 5673 18540 5725
rect 18592 5673 18751 5725
rect 18803 5673 18962 5725
rect 19014 5673 19173 5725
rect 19225 5673 19384 5725
rect 19436 5673 19588 5725
rect 18387 5428 19588 5673
rect 18387 5372 18433 5428
rect 18489 5372 18643 5428
rect 18699 5372 18854 5428
rect 18910 5372 19066 5428
rect 19122 5372 19277 5428
rect 19333 5372 19487 5428
rect 19543 5372 19588 5428
rect 18387 5127 19588 5372
rect 18387 5075 18540 5127
rect 18592 5075 18751 5127
rect 18803 5075 18962 5127
rect 19014 5075 19173 5127
rect 19225 5075 19384 5127
rect 19436 5075 19588 5127
rect 18154 5022 18284 5061
rect 18154 4966 18191 5022
rect 18247 4966 18284 5022
rect 18154 4804 18284 4966
rect 18154 4748 18191 4804
rect 18247 4748 18284 4804
rect 18154 4710 18284 4748
rect 18387 4664 19588 5075
rect 18387 4612 18540 4664
rect 18592 4612 18751 4664
rect 18803 4612 18962 4664
rect 19014 4612 19173 4664
rect 19225 4612 19384 4664
rect 19436 4612 19588 4664
rect 18387 4388 19588 4612
rect 18387 4336 18540 4388
rect 18592 4336 18751 4388
rect 18803 4336 18962 4388
rect 19014 4336 19173 4388
rect 19225 4336 19384 4388
rect 19436 4336 19588 4388
rect 18154 4252 18284 4290
rect 18154 4196 18191 4252
rect 18247 4196 18284 4252
rect 18154 4034 18284 4196
rect 18154 3978 18191 4034
rect 18247 3978 18284 4034
rect 18154 3939 18284 3978
rect 18387 3925 19588 4336
rect 18387 3873 18540 3925
rect 18592 3873 18751 3925
rect 18803 3873 18962 3925
rect 19014 3873 19173 3925
rect 19225 3873 19384 3925
rect 19436 3873 19588 3925
rect 18387 3628 19588 3873
rect 18387 3572 18433 3628
rect 18489 3572 18643 3628
rect 18699 3572 18854 3628
rect 18910 3572 19066 3628
rect 19122 3572 19277 3628
rect 19333 3572 19487 3628
rect 19543 3572 19588 3628
rect 18387 3327 19588 3572
rect 18387 3275 18540 3327
rect 18592 3275 18751 3327
rect 18803 3275 18962 3327
rect 19014 3275 19173 3327
rect 19225 3275 19384 3327
rect 19436 3275 19588 3327
rect 18154 3222 18284 3261
rect 18154 3166 18191 3222
rect 18247 3166 18284 3222
rect 18154 3004 18284 3166
rect 18154 2948 18191 3004
rect 18247 2948 18284 3004
rect 18154 2910 18284 2948
rect 18387 2864 19588 3275
rect 18387 2812 18540 2864
rect 18592 2812 18751 2864
rect 18803 2812 18962 2864
rect 19014 2812 19173 2864
rect 19225 2812 19384 2864
rect 19436 2812 19588 2864
rect 18387 2588 19588 2812
rect 18387 2536 18540 2588
rect 18592 2536 18751 2588
rect 18803 2536 18962 2588
rect 19014 2536 19173 2588
rect 19225 2536 19384 2588
rect 19436 2536 19588 2588
rect 18154 2452 18284 2490
rect 18154 2396 18191 2452
rect 18247 2396 18284 2452
rect 18154 2234 18284 2396
rect 18154 2178 18191 2234
rect 18247 2178 18284 2234
rect 18154 2139 18284 2178
rect 18387 2125 19588 2536
rect 18387 2073 18540 2125
rect 18592 2073 18751 2125
rect 18803 2073 18962 2125
rect 19014 2073 19173 2125
rect 19225 2073 19384 2125
rect 19436 2073 19588 2125
rect 18387 1828 19588 2073
rect 18387 1772 18433 1828
rect 18489 1772 18643 1828
rect 18699 1772 18854 1828
rect 18910 1772 19066 1828
rect 19122 1772 19277 1828
rect 19333 1772 19487 1828
rect 19543 1772 19588 1828
rect 18387 1527 19588 1772
rect 18387 1475 18540 1527
rect 18592 1475 18751 1527
rect 18803 1475 18962 1527
rect 19014 1475 19173 1527
rect 19225 1475 19384 1527
rect 19436 1475 19588 1527
rect 18154 1422 18284 1461
rect 18154 1366 18191 1422
rect 18247 1366 18284 1422
rect 18154 1204 18284 1366
rect 18154 1148 18191 1204
rect 18247 1148 18284 1204
rect 18154 1110 18284 1148
rect 18387 1064 19588 1475
rect 18387 1012 18540 1064
rect 18592 1012 18751 1064
rect 18803 1012 18962 1064
rect 19014 1012 19173 1064
rect 19225 1012 19384 1064
rect 19436 1012 19588 1064
rect 18387 788 19588 1012
rect 18387 736 18540 788
rect 18592 736 18751 788
rect 18803 736 18962 788
rect 19014 736 19173 788
rect 19225 736 19384 788
rect 19436 736 19588 788
rect 17755 552 17838 604
rect 17890 552 17976 604
rect 17755 -164 17976 552
rect 18154 652 18284 690
rect 18154 596 18191 652
rect 18247 596 18284 652
rect 18154 434 18284 596
rect 18154 378 18191 434
rect 18247 378 18284 434
rect 18154 339 18284 378
rect 18387 325 19588 736
rect 18387 273 18540 325
rect 18592 273 18751 325
rect 18803 273 18962 325
rect 19014 273 19173 325
rect 19225 273 19384 325
rect 19436 273 19588 325
rect 18387 28 19588 273
rect 18387 -28 18433 28
rect 18489 -28 18643 28
rect 18699 -28 18854 28
rect 18910 -28 19066 28
rect 19122 -28 19277 28
rect 19333 -28 19487 28
rect 19543 -28 19588 28
rect 18387 -151 19588 -28
rect 19696 14426 20510 14551
rect 19696 14374 19943 14426
rect 19995 14374 20154 14426
rect 20206 14374 20365 14426
rect 20417 14374 20510 14426
rect 19696 13964 20510 14374
rect 21824 14428 23952 14551
rect 21824 14372 21911 14428
rect 21967 14372 22122 14428
rect 22178 14372 22333 14428
rect 22389 14372 22543 14428
rect 22599 14372 22754 14428
rect 22810 14372 22966 14428
rect 23022 14372 23177 14428
rect 23233 14372 23387 14428
rect 23443 14372 23598 14428
rect 23654 14372 23809 14428
rect 23865 14372 23952 14428
rect 19696 13912 19897 13964
rect 19949 13912 20108 13964
rect 20160 13912 20319 13964
rect 20371 13912 20510 13964
rect 19696 13528 20510 13912
rect 20631 14202 20941 14243
rect 20631 14150 20670 14202
rect 20722 14150 20850 14202
rect 20902 14150 20941 14202
rect 20631 13988 20941 14150
rect 20631 13932 20668 13988
rect 20724 13932 20848 13988
rect 20904 13932 20941 13988
rect 20631 13859 20941 13932
rect 21393 14195 21703 14236
rect 21393 14143 21432 14195
rect 21484 14143 21612 14195
rect 21664 14143 21703 14195
rect 21393 13988 21703 14143
rect 21393 13932 21430 13988
rect 21486 13932 21610 13988
rect 21666 13932 21703 13988
rect 21393 13732 21703 13932
rect 21393 13680 21432 13732
rect 21484 13680 21612 13732
rect 21664 13680 21703 13732
rect 21393 13640 21703 13680
rect 19696 13526 19758 13528
rect 19814 13526 19969 13528
rect 19696 13474 19735 13526
rect 19814 13474 19915 13526
rect 19967 13474 19969 13526
rect 19696 13472 19758 13474
rect 19814 13472 19969 13474
rect 20025 13472 20181 13528
rect 20237 13472 20392 13528
rect 20448 13472 20510 13528
rect 19696 13088 20510 13472
rect 21824 13526 23952 14372
rect 21824 13474 21913 13526
rect 21965 13474 22124 13526
rect 22176 13474 22335 13526
rect 22387 13474 22545 13526
rect 22597 13474 22756 13526
rect 22808 13474 22968 13526
rect 23020 13474 23179 13526
rect 23231 13474 23389 13526
rect 23441 13474 23600 13526
rect 23652 13474 23811 13526
rect 23863 13474 23952 13526
rect 21393 13320 21703 13360
rect 21393 13268 21432 13320
rect 21484 13268 21612 13320
rect 21664 13268 21703 13320
rect 19696 13036 19897 13088
rect 19949 13036 20108 13088
rect 20160 13036 20319 13088
rect 20371 13036 20510 13088
rect 19696 12626 20510 13036
rect 20631 13068 20941 13141
rect 20631 13012 20668 13068
rect 20724 13012 20848 13068
rect 20904 13012 20941 13068
rect 20631 12850 20941 13012
rect 20631 12798 20670 12850
rect 20722 12798 20850 12850
rect 20902 12798 20941 12850
rect 20631 12757 20941 12798
rect 21393 13068 21703 13268
rect 21393 13012 21430 13068
rect 21486 13012 21610 13068
rect 21666 13012 21703 13068
rect 21393 12857 21703 13012
rect 21393 12805 21432 12857
rect 21484 12805 21612 12857
rect 21664 12805 21703 12857
rect 21393 12764 21703 12805
rect 19696 12574 19943 12626
rect 19995 12574 20154 12626
rect 20206 12574 20365 12626
rect 20417 12574 20510 12626
rect 19696 12164 20510 12574
rect 21824 12628 23952 13474
rect 21824 12572 21911 12628
rect 21967 12572 22122 12628
rect 22178 12572 22333 12628
rect 22389 12572 22543 12628
rect 22599 12572 22754 12628
rect 22810 12572 22966 12628
rect 23022 12572 23177 12628
rect 23233 12572 23387 12628
rect 23443 12572 23598 12628
rect 23654 12572 23809 12628
rect 23865 12572 23952 12628
rect 19696 12112 19897 12164
rect 19949 12112 20108 12164
rect 20160 12112 20319 12164
rect 20371 12112 20510 12164
rect 19696 11728 20510 12112
rect 20631 12402 20941 12443
rect 20631 12350 20670 12402
rect 20722 12350 20850 12402
rect 20902 12350 20941 12402
rect 20631 12188 20941 12350
rect 20631 12132 20668 12188
rect 20724 12132 20848 12188
rect 20904 12132 20941 12188
rect 20631 12059 20941 12132
rect 21393 12395 21703 12436
rect 21393 12343 21432 12395
rect 21484 12343 21612 12395
rect 21664 12343 21703 12395
rect 21393 12188 21703 12343
rect 21393 12132 21430 12188
rect 21486 12132 21610 12188
rect 21666 12132 21703 12188
rect 21393 11932 21703 12132
rect 21393 11880 21432 11932
rect 21484 11880 21612 11932
rect 21664 11880 21703 11932
rect 21393 11840 21703 11880
rect 19696 11726 19758 11728
rect 19814 11726 19969 11728
rect 19696 11674 19735 11726
rect 19814 11674 19915 11726
rect 19967 11674 19969 11726
rect 19696 11672 19758 11674
rect 19814 11672 19969 11674
rect 20025 11672 20181 11728
rect 20237 11672 20392 11728
rect 20448 11672 20510 11728
rect 19696 11288 20510 11672
rect 21824 11726 23952 12572
rect 21824 11674 21913 11726
rect 21965 11674 22124 11726
rect 22176 11674 22335 11726
rect 22387 11674 22545 11726
rect 22597 11674 22756 11726
rect 22808 11674 22968 11726
rect 23020 11674 23179 11726
rect 23231 11674 23389 11726
rect 23441 11674 23600 11726
rect 23652 11674 23811 11726
rect 23863 11674 23952 11726
rect 21393 11520 21703 11560
rect 21393 11468 21432 11520
rect 21484 11468 21612 11520
rect 21664 11468 21703 11520
rect 19696 11236 19897 11288
rect 19949 11236 20108 11288
rect 20160 11236 20319 11288
rect 20371 11236 20510 11288
rect 19696 10826 20510 11236
rect 20631 11268 20941 11341
rect 20631 11212 20668 11268
rect 20724 11212 20848 11268
rect 20904 11212 20941 11268
rect 20631 11050 20941 11212
rect 20631 10998 20670 11050
rect 20722 10998 20850 11050
rect 20902 10998 20941 11050
rect 20631 10957 20941 10998
rect 21393 11268 21703 11468
rect 21393 11212 21430 11268
rect 21486 11212 21610 11268
rect 21666 11212 21703 11268
rect 21393 11057 21703 11212
rect 21393 11005 21432 11057
rect 21484 11005 21612 11057
rect 21664 11005 21703 11057
rect 21393 10964 21703 11005
rect 19696 10774 19943 10826
rect 19995 10774 20154 10826
rect 20206 10774 20365 10826
rect 20417 10774 20510 10826
rect 19696 10364 20510 10774
rect 21824 10828 23952 11674
rect 21824 10772 21911 10828
rect 21967 10772 22122 10828
rect 22178 10772 22333 10828
rect 22389 10772 22543 10828
rect 22599 10772 22754 10828
rect 22810 10772 22966 10828
rect 23022 10772 23177 10828
rect 23233 10772 23387 10828
rect 23443 10772 23598 10828
rect 23654 10772 23809 10828
rect 23865 10772 23952 10828
rect 19696 10312 19897 10364
rect 19949 10312 20108 10364
rect 20160 10312 20319 10364
rect 20371 10312 20510 10364
rect 19696 9928 20510 10312
rect 20631 10602 20941 10643
rect 20631 10550 20670 10602
rect 20722 10550 20850 10602
rect 20902 10550 20941 10602
rect 20631 10388 20941 10550
rect 20631 10332 20668 10388
rect 20724 10332 20848 10388
rect 20904 10332 20941 10388
rect 20631 10259 20941 10332
rect 21393 10595 21703 10636
rect 21393 10543 21432 10595
rect 21484 10543 21612 10595
rect 21664 10543 21703 10595
rect 21393 10388 21703 10543
rect 21393 10332 21430 10388
rect 21486 10332 21610 10388
rect 21666 10332 21703 10388
rect 21393 10132 21703 10332
rect 21393 10080 21432 10132
rect 21484 10080 21612 10132
rect 21664 10080 21703 10132
rect 21393 10040 21703 10080
rect 19696 9926 19758 9928
rect 19814 9926 19969 9928
rect 19696 9874 19735 9926
rect 19814 9874 19915 9926
rect 19967 9874 19969 9926
rect 19696 9872 19758 9874
rect 19814 9872 19969 9874
rect 20025 9872 20181 9928
rect 20237 9872 20392 9928
rect 20448 9872 20510 9928
rect 19696 9488 20510 9872
rect 21824 9926 23952 10772
rect 21824 9874 21913 9926
rect 21965 9874 22124 9926
rect 22176 9874 22335 9926
rect 22387 9874 22545 9926
rect 22597 9874 22756 9926
rect 22808 9874 22968 9926
rect 23020 9874 23179 9926
rect 23231 9874 23389 9926
rect 23441 9874 23600 9926
rect 23652 9874 23811 9926
rect 23863 9874 23952 9926
rect 21393 9720 21703 9760
rect 21393 9668 21432 9720
rect 21484 9668 21612 9720
rect 21664 9668 21703 9720
rect 19696 9436 19897 9488
rect 19949 9436 20108 9488
rect 20160 9436 20319 9488
rect 20371 9436 20510 9488
rect 19696 9026 20510 9436
rect 20631 9468 20941 9541
rect 20631 9412 20668 9468
rect 20724 9412 20848 9468
rect 20904 9412 20941 9468
rect 20631 9250 20941 9412
rect 20631 9198 20670 9250
rect 20722 9198 20850 9250
rect 20902 9198 20941 9250
rect 20631 9157 20941 9198
rect 21393 9468 21703 9668
rect 21393 9412 21430 9468
rect 21486 9412 21610 9468
rect 21666 9412 21703 9468
rect 21393 9257 21703 9412
rect 21393 9205 21432 9257
rect 21484 9205 21612 9257
rect 21664 9205 21703 9257
rect 21393 9164 21703 9205
rect 19696 8974 19943 9026
rect 19995 8974 20154 9026
rect 20206 8974 20365 9026
rect 20417 8974 20510 9026
rect 19696 8564 20510 8974
rect 21824 9028 23952 9874
rect 21824 8972 21911 9028
rect 21967 8972 22122 9028
rect 22178 8972 22333 9028
rect 22389 8972 22543 9028
rect 22599 8972 22754 9028
rect 22810 8972 22966 9028
rect 23022 8972 23177 9028
rect 23233 8972 23387 9028
rect 23443 8972 23598 9028
rect 23654 8972 23809 9028
rect 23865 8972 23952 9028
rect 19696 8512 19897 8564
rect 19949 8512 20108 8564
rect 20160 8512 20319 8564
rect 20371 8512 20510 8564
rect 19696 8128 20510 8512
rect 20631 8802 20941 8843
rect 20631 8750 20670 8802
rect 20722 8750 20850 8802
rect 20902 8750 20941 8802
rect 20631 8588 20941 8750
rect 20631 8532 20668 8588
rect 20724 8532 20848 8588
rect 20904 8532 20941 8588
rect 20631 8459 20941 8532
rect 21393 8795 21703 8836
rect 21393 8743 21432 8795
rect 21484 8743 21612 8795
rect 21664 8743 21703 8795
rect 21393 8588 21703 8743
rect 21393 8532 21430 8588
rect 21486 8532 21610 8588
rect 21666 8532 21703 8588
rect 21393 8332 21703 8532
rect 21393 8280 21432 8332
rect 21484 8280 21612 8332
rect 21664 8280 21703 8332
rect 21393 8240 21703 8280
rect 19696 8126 19758 8128
rect 19814 8126 19969 8128
rect 19696 8074 19735 8126
rect 19814 8074 19915 8126
rect 19967 8074 19969 8126
rect 19696 8072 19758 8074
rect 19814 8072 19969 8074
rect 20025 8072 20181 8128
rect 20237 8072 20392 8128
rect 20448 8072 20510 8128
rect 19696 7688 20510 8072
rect 21824 8126 23952 8972
rect 21824 8074 21913 8126
rect 21965 8074 22124 8126
rect 22176 8074 22335 8126
rect 22387 8074 22545 8126
rect 22597 8074 22756 8126
rect 22808 8074 22968 8126
rect 23020 8074 23179 8126
rect 23231 8074 23389 8126
rect 23441 8074 23600 8126
rect 23652 8074 23811 8126
rect 23863 8074 23952 8126
rect 21393 7920 21703 7960
rect 21393 7868 21432 7920
rect 21484 7868 21612 7920
rect 21664 7868 21703 7920
rect 19696 7636 19897 7688
rect 19949 7636 20108 7688
rect 20160 7636 20319 7688
rect 20371 7636 20510 7688
rect 19696 7226 20510 7636
rect 20631 7668 20941 7741
rect 20631 7612 20668 7668
rect 20724 7612 20848 7668
rect 20904 7612 20941 7668
rect 20631 7450 20941 7612
rect 20631 7398 20670 7450
rect 20722 7398 20850 7450
rect 20902 7398 20941 7450
rect 20631 7357 20941 7398
rect 21393 7668 21703 7868
rect 21393 7612 21430 7668
rect 21486 7612 21610 7668
rect 21666 7612 21703 7668
rect 21393 7457 21703 7612
rect 21393 7405 21432 7457
rect 21484 7405 21612 7457
rect 21664 7405 21703 7457
rect 21393 7364 21703 7405
rect 19696 7174 19943 7226
rect 19995 7174 20154 7226
rect 20206 7174 20365 7226
rect 20417 7174 20510 7226
rect 19696 6764 20510 7174
rect 21824 7228 23952 8074
rect 21824 7172 21911 7228
rect 21967 7172 22122 7228
rect 22178 7172 22333 7228
rect 22389 7172 22543 7228
rect 22599 7172 22754 7228
rect 22810 7172 22966 7228
rect 23022 7172 23177 7228
rect 23233 7172 23387 7228
rect 23443 7172 23598 7228
rect 23654 7172 23809 7228
rect 23865 7172 23952 7228
rect 19696 6712 19897 6764
rect 19949 6712 20108 6764
rect 20160 6712 20319 6764
rect 20371 6712 20510 6764
rect 19696 6328 20510 6712
rect 20631 7002 20941 7043
rect 20631 6950 20670 7002
rect 20722 6950 20850 7002
rect 20902 6950 20941 7002
rect 20631 6788 20941 6950
rect 20631 6732 20668 6788
rect 20724 6732 20848 6788
rect 20904 6732 20941 6788
rect 20631 6659 20941 6732
rect 21393 6995 21703 7036
rect 21393 6943 21432 6995
rect 21484 6943 21612 6995
rect 21664 6943 21703 6995
rect 21393 6788 21703 6943
rect 21393 6732 21430 6788
rect 21486 6732 21610 6788
rect 21666 6732 21703 6788
rect 21393 6532 21703 6732
rect 21393 6480 21432 6532
rect 21484 6480 21612 6532
rect 21664 6480 21703 6532
rect 21393 6440 21703 6480
rect 19696 6326 19758 6328
rect 19814 6326 19969 6328
rect 19696 6274 19735 6326
rect 19814 6274 19915 6326
rect 19967 6274 19969 6326
rect 19696 6272 19758 6274
rect 19814 6272 19969 6274
rect 20025 6272 20181 6328
rect 20237 6272 20392 6328
rect 20448 6272 20510 6328
rect 19696 5888 20510 6272
rect 21824 6326 23952 7172
rect 21824 6274 21913 6326
rect 21965 6274 22124 6326
rect 22176 6274 22335 6326
rect 22387 6274 22545 6326
rect 22597 6274 22756 6326
rect 22808 6274 22968 6326
rect 23020 6274 23179 6326
rect 23231 6274 23389 6326
rect 23441 6274 23600 6326
rect 23652 6274 23811 6326
rect 23863 6274 23952 6326
rect 21393 6120 21703 6160
rect 21393 6068 21432 6120
rect 21484 6068 21612 6120
rect 21664 6068 21703 6120
rect 19696 5836 19897 5888
rect 19949 5836 20108 5888
rect 20160 5836 20319 5888
rect 20371 5836 20510 5888
rect 19696 5426 20510 5836
rect 20631 5868 20941 5941
rect 20631 5812 20668 5868
rect 20724 5812 20848 5868
rect 20904 5812 20941 5868
rect 20631 5650 20941 5812
rect 20631 5598 20670 5650
rect 20722 5598 20850 5650
rect 20902 5598 20941 5650
rect 20631 5557 20941 5598
rect 21393 5868 21703 6068
rect 21393 5812 21430 5868
rect 21486 5812 21610 5868
rect 21666 5812 21703 5868
rect 21393 5657 21703 5812
rect 21393 5605 21432 5657
rect 21484 5605 21612 5657
rect 21664 5605 21703 5657
rect 21393 5564 21703 5605
rect 19696 5374 19943 5426
rect 19995 5374 20154 5426
rect 20206 5374 20365 5426
rect 20417 5374 20510 5426
rect 19696 4964 20510 5374
rect 21824 5428 23952 6274
rect 21824 5372 21911 5428
rect 21967 5372 22122 5428
rect 22178 5372 22333 5428
rect 22389 5372 22543 5428
rect 22599 5372 22754 5428
rect 22810 5372 22966 5428
rect 23022 5372 23177 5428
rect 23233 5372 23387 5428
rect 23443 5372 23598 5428
rect 23654 5372 23809 5428
rect 23865 5372 23952 5428
rect 19696 4912 19897 4964
rect 19949 4912 20108 4964
rect 20160 4912 20319 4964
rect 20371 4912 20510 4964
rect 19696 4528 20510 4912
rect 20631 5202 20941 5243
rect 20631 5150 20670 5202
rect 20722 5150 20850 5202
rect 20902 5150 20941 5202
rect 20631 4988 20941 5150
rect 20631 4932 20668 4988
rect 20724 4932 20848 4988
rect 20904 4932 20941 4988
rect 20631 4859 20941 4932
rect 21393 5195 21703 5236
rect 21393 5143 21432 5195
rect 21484 5143 21612 5195
rect 21664 5143 21703 5195
rect 21393 4988 21703 5143
rect 21393 4932 21430 4988
rect 21486 4932 21610 4988
rect 21666 4932 21703 4988
rect 21393 4732 21703 4932
rect 21393 4680 21432 4732
rect 21484 4680 21612 4732
rect 21664 4680 21703 4732
rect 21393 4640 21703 4680
rect 19696 4526 19758 4528
rect 19814 4526 19969 4528
rect 19696 4474 19735 4526
rect 19814 4474 19915 4526
rect 19967 4474 19969 4526
rect 19696 4472 19758 4474
rect 19814 4472 19969 4474
rect 20025 4472 20181 4528
rect 20237 4472 20392 4528
rect 20448 4472 20510 4528
rect 19696 4088 20510 4472
rect 21824 4526 23952 5372
rect 21824 4474 21913 4526
rect 21965 4474 22124 4526
rect 22176 4474 22335 4526
rect 22387 4474 22545 4526
rect 22597 4474 22756 4526
rect 22808 4474 22968 4526
rect 23020 4474 23179 4526
rect 23231 4474 23389 4526
rect 23441 4474 23600 4526
rect 23652 4474 23811 4526
rect 23863 4474 23952 4526
rect 21393 4320 21703 4360
rect 21393 4268 21432 4320
rect 21484 4268 21612 4320
rect 21664 4268 21703 4320
rect 19696 4036 19897 4088
rect 19949 4036 20108 4088
rect 20160 4036 20319 4088
rect 20371 4036 20510 4088
rect 19696 3626 20510 4036
rect 20631 4068 20941 4141
rect 20631 4012 20668 4068
rect 20724 4012 20848 4068
rect 20904 4012 20941 4068
rect 20631 3850 20941 4012
rect 20631 3798 20670 3850
rect 20722 3798 20850 3850
rect 20902 3798 20941 3850
rect 20631 3757 20941 3798
rect 21393 4068 21703 4268
rect 21393 4012 21430 4068
rect 21486 4012 21610 4068
rect 21666 4012 21703 4068
rect 21393 3857 21703 4012
rect 21393 3805 21432 3857
rect 21484 3805 21612 3857
rect 21664 3805 21703 3857
rect 21393 3764 21703 3805
rect 19696 3574 19943 3626
rect 19995 3574 20154 3626
rect 20206 3574 20365 3626
rect 20417 3574 20510 3626
rect 19696 3164 20510 3574
rect 21824 3628 23952 4474
rect 21824 3572 21911 3628
rect 21967 3572 22122 3628
rect 22178 3572 22333 3628
rect 22389 3572 22543 3628
rect 22599 3572 22754 3628
rect 22810 3572 22966 3628
rect 23022 3572 23177 3628
rect 23233 3572 23387 3628
rect 23443 3572 23598 3628
rect 23654 3572 23809 3628
rect 23865 3572 23952 3628
rect 19696 3112 19897 3164
rect 19949 3112 20108 3164
rect 20160 3112 20319 3164
rect 20371 3112 20510 3164
rect 19696 2728 20510 3112
rect 20631 3402 20941 3443
rect 20631 3350 20670 3402
rect 20722 3350 20850 3402
rect 20902 3350 20941 3402
rect 20631 3188 20941 3350
rect 20631 3132 20668 3188
rect 20724 3132 20848 3188
rect 20904 3132 20941 3188
rect 20631 3059 20941 3132
rect 21393 3395 21703 3436
rect 21393 3343 21432 3395
rect 21484 3343 21612 3395
rect 21664 3343 21703 3395
rect 21393 3188 21703 3343
rect 21393 3132 21430 3188
rect 21486 3132 21610 3188
rect 21666 3132 21703 3188
rect 21393 2932 21703 3132
rect 21393 2880 21432 2932
rect 21484 2880 21612 2932
rect 21664 2880 21703 2932
rect 21393 2840 21703 2880
rect 19696 2726 19758 2728
rect 19814 2726 19969 2728
rect 19696 2674 19735 2726
rect 19814 2674 19915 2726
rect 19967 2674 19969 2726
rect 19696 2672 19758 2674
rect 19814 2672 19969 2674
rect 20025 2672 20181 2728
rect 20237 2672 20392 2728
rect 20448 2672 20510 2728
rect 19696 2288 20510 2672
rect 21824 2726 23952 3572
rect 21824 2674 21913 2726
rect 21965 2674 22124 2726
rect 22176 2674 22335 2726
rect 22387 2674 22545 2726
rect 22597 2674 22756 2726
rect 22808 2674 22968 2726
rect 23020 2674 23179 2726
rect 23231 2674 23389 2726
rect 23441 2674 23600 2726
rect 23652 2674 23811 2726
rect 23863 2674 23952 2726
rect 21393 2520 21703 2560
rect 21393 2468 21432 2520
rect 21484 2468 21612 2520
rect 21664 2468 21703 2520
rect 19696 2236 19897 2288
rect 19949 2236 20108 2288
rect 20160 2236 20319 2288
rect 20371 2236 20510 2288
rect 19696 1826 20510 2236
rect 20631 2268 20941 2341
rect 20631 2212 20668 2268
rect 20724 2212 20848 2268
rect 20904 2212 20941 2268
rect 20631 2050 20941 2212
rect 20631 1998 20670 2050
rect 20722 1998 20850 2050
rect 20902 1998 20941 2050
rect 20631 1957 20941 1998
rect 21393 2268 21703 2468
rect 21393 2212 21430 2268
rect 21486 2212 21610 2268
rect 21666 2212 21703 2268
rect 21393 2057 21703 2212
rect 21393 2005 21432 2057
rect 21484 2005 21612 2057
rect 21664 2005 21703 2057
rect 21393 1964 21703 2005
rect 19696 1774 19943 1826
rect 19995 1774 20154 1826
rect 20206 1774 20365 1826
rect 20417 1774 20510 1826
rect 19696 1364 20510 1774
rect 21824 1828 23952 2674
rect 21824 1772 21911 1828
rect 21967 1772 22122 1828
rect 22178 1772 22333 1828
rect 22389 1772 22543 1828
rect 22599 1772 22754 1828
rect 22810 1772 22966 1828
rect 23022 1772 23177 1828
rect 23233 1772 23387 1828
rect 23443 1772 23598 1828
rect 23654 1772 23809 1828
rect 23865 1772 23952 1828
rect 19696 1312 19897 1364
rect 19949 1312 20108 1364
rect 20160 1312 20319 1364
rect 20371 1312 20510 1364
rect 19696 928 20510 1312
rect 20631 1602 20941 1643
rect 20631 1550 20670 1602
rect 20722 1550 20850 1602
rect 20902 1550 20941 1602
rect 20631 1388 20941 1550
rect 20631 1332 20668 1388
rect 20724 1332 20848 1388
rect 20904 1332 20941 1388
rect 20631 1259 20941 1332
rect 21393 1595 21703 1636
rect 21393 1543 21432 1595
rect 21484 1543 21612 1595
rect 21664 1543 21703 1595
rect 21393 1388 21703 1543
rect 21393 1332 21430 1388
rect 21486 1332 21610 1388
rect 21666 1332 21703 1388
rect 21393 1132 21703 1332
rect 21393 1080 21432 1132
rect 21484 1080 21612 1132
rect 21664 1080 21703 1132
rect 21393 1040 21703 1080
rect 19696 926 19758 928
rect 19814 926 19969 928
rect 19696 874 19735 926
rect 19814 874 19915 926
rect 19967 874 19969 926
rect 19696 872 19758 874
rect 19814 872 19969 874
rect 20025 872 20181 928
rect 20237 872 20392 928
rect 20448 872 20510 928
rect 19696 488 20510 872
rect 21824 926 23952 1772
rect 21824 874 21913 926
rect 21965 874 22124 926
rect 22176 874 22335 926
rect 22387 874 22545 926
rect 22597 874 22756 926
rect 22808 874 22968 926
rect 23020 874 23179 926
rect 23231 874 23389 926
rect 23441 874 23600 926
rect 23652 874 23811 926
rect 23863 874 23952 926
rect 21393 720 21703 760
rect 21393 668 21432 720
rect 21484 668 21612 720
rect 21664 668 21703 720
rect 19696 436 19897 488
rect 19949 436 20108 488
rect 20160 436 20319 488
rect 20371 436 20510 488
rect 19696 26 20510 436
rect 20631 468 20941 541
rect 20631 412 20668 468
rect 20724 412 20848 468
rect 20904 412 20941 468
rect 20631 250 20941 412
rect 20631 198 20670 250
rect 20722 198 20850 250
rect 20902 198 20941 250
rect 20631 157 20941 198
rect 21393 468 21703 668
rect 21393 412 21430 468
rect 21486 412 21610 468
rect 21666 412 21703 468
rect 21393 257 21703 412
rect 21393 205 21432 257
rect 21484 205 21612 257
rect 21664 205 21703 257
rect 21393 164 21703 205
rect 19696 -26 19943 26
rect 19995 -26 20154 26
rect 20206 -26 20365 26
rect 20417 -26 20510 26
rect 19696 -151 20510 -26
rect 21824 28 23952 874
rect 21824 -28 21911 28
rect 21967 -28 22122 28
rect 22178 -28 22333 28
rect 22389 -28 22543 28
rect 22599 -28 22754 28
rect 22810 -28 22966 28
rect 23022 -28 23177 28
rect 23233 -28 23387 28
rect 23443 -28 23598 28
rect 23654 -28 23809 28
rect 23865 -28 23952 28
rect 21824 -151 23952 -28
<< via2 >>
rect 449 14426 505 14428
rect 449 14374 451 14426
rect 451 14374 503 14426
rect 503 14374 505 14426
rect 449 14372 505 14374
rect 660 14426 716 14428
rect 660 14374 662 14426
rect 662 14374 714 14426
rect 714 14374 716 14426
rect 660 14372 716 14374
rect 871 14426 927 14428
rect 871 14374 873 14426
rect 873 14374 925 14426
rect 925 14374 927 14426
rect 871 14372 927 14374
rect 1081 14426 1137 14428
rect 1081 14374 1083 14426
rect 1083 14374 1135 14426
rect 1135 14374 1137 14426
rect 1081 14372 1137 14374
rect 1292 14426 1348 14428
rect 1292 14374 1294 14426
rect 1294 14374 1346 14426
rect 1346 14374 1348 14426
rect 1292 14372 1348 14374
rect 1504 14426 1560 14428
rect 1504 14374 1506 14426
rect 1506 14374 1558 14426
rect 1558 14374 1560 14426
rect 1504 14372 1560 14374
rect 1715 14426 1771 14428
rect 1715 14374 1717 14426
rect 1717 14374 1769 14426
rect 1769 14374 1771 14426
rect 1715 14372 1771 14374
rect 1925 14426 1981 14428
rect 1925 14374 1927 14426
rect 1927 14374 1979 14426
rect 1979 14374 1981 14426
rect 1925 14372 1981 14374
rect 2136 14426 2192 14428
rect 2136 14374 2138 14426
rect 2138 14374 2190 14426
rect 2190 14374 2192 14426
rect 2136 14372 2192 14374
rect 2347 14426 2403 14428
rect 2347 14374 2349 14426
rect 2349 14374 2401 14426
rect 2401 14374 2403 14426
rect 2347 14372 2403 14374
rect 2652 13939 2708 13995
rect 2832 13939 2888 13995
rect 3414 13932 3470 13988
rect 3594 13932 3650 13988
rect 3879 13472 3935 13528
rect 4090 13472 4146 13528
rect 4302 13526 4358 13528
rect 4513 13526 4569 13528
rect 4302 13474 4352 13526
rect 4352 13474 4358 13526
rect 4513 13474 4532 13526
rect 4532 13474 4569 13526
rect 4302 13472 4358 13474
rect 4513 13472 4569 13474
rect 2652 13005 2708 13061
rect 2832 13005 2888 13061
rect 3414 13012 3470 13068
rect 3594 13012 3650 13068
rect 449 12626 505 12628
rect 449 12574 451 12626
rect 451 12574 503 12626
rect 503 12574 505 12626
rect 449 12572 505 12574
rect 660 12626 716 12628
rect 660 12574 662 12626
rect 662 12574 714 12626
rect 714 12574 716 12626
rect 660 12572 716 12574
rect 871 12626 927 12628
rect 871 12574 873 12626
rect 873 12574 925 12626
rect 925 12574 927 12626
rect 871 12572 927 12574
rect 1081 12626 1137 12628
rect 1081 12574 1083 12626
rect 1083 12574 1135 12626
rect 1135 12574 1137 12626
rect 1081 12572 1137 12574
rect 1292 12626 1348 12628
rect 1292 12574 1294 12626
rect 1294 12574 1346 12626
rect 1346 12574 1348 12626
rect 1292 12572 1348 12574
rect 1504 12626 1560 12628
rect 1504 12574 1506 12626
rect 1506 12574 1558 12626
rect 1558 12574 1560 12626
rect 1504 12572 1560 12574
rect 1715 12626 1771 12628
rect 1715 12574 1717 12626
rect 1717 12574 1769 12626
rect 1769 12574 1771 12626
rect 1715 12572 1771 12574
rect 1925 12626 1981 12628
rect 1925 12574 1927 12626
rect 1927 12574 1979 12626
rect 1979 12574 1981 12626
rect 1925 12572 1981 12574
rect 2136 12626 2192 12628
rect 2136 12574 2138 12626
rect 2138 12574 2190 12626
rect 2190 12574 2192 12626
rect 2136 12572 2192 12574
rect 2347 12626 2403 12628
rect 2347 12574 2349 12626
rect 2349 12574 2401 12626
rect 2401 12574 2403 12626
rect 2347 12572 2403 12574
rect 2652 12139 2708 12195
rect 2832 12139 2888 12195
rect 3414 12132 3470 12188
rect 3594 12132 3650 12188
rect 3879 11672 3935 11728
rect 4090 11672 4146 11728
rect 4302 11726 4358 11728
rect 4513 11726 4569 11728
rect 4302 11674 4352 11726
rect 4352 11674 4358 11726
rect 4513 11674 4532 11726
rect 4532 11674 4569 11726
rect 4302 11672 4358 11674
rect 4513 11672 4569 11674
rect 2652 11205 2708 11261
rect 2832 11205 2888 11261
rect 3414 11212 3470 11268
rect 3594 11212 3650 11268
rect 449 10826 505 10828
rect 449 10774 451 10826
rect 451 10774 503 10826
rect 503 10774 505 10826
rect 449 10772 505 10774
rect 660 10826 716 10828
rect 660 10774 662 10826
rect 662 10774 714 10826
rect 714 10774 716 10826
rect 660 10772 716 10774
rect 871 10826 927 10828
rect 871 10774 873 10826
rect 873 10774 925 10826
rect 925 10774 927 10826
rect 871 10772 927 10774
rect 1081 10826 1137 10828
rect 1081 10774 1083 10826
rect 1083 10774 1135 10826
rect 1135 10774 1137 10826
rect 1081 10772 1137 10774
rect 1292 10826 1348 10828
rect 1292 10774 1294 10826
rect 1294 10774 1346 10826
rect 1346 10774 1348 10826
rect 1292 10772 1348 10774
rect 1504 10826 1560 10828
rect 1504 10774 1506 10826
rect 1506 10774 1558 10826
rect 1558 10774 1560 10826
rect 1504 10772 1560 10774
rect 1715 10826 1771 10828
rect 1715 10774 1717 10826
rect 1717 10774 1769 10826
rect 1769 10774 1771 10826
rect 1715 10772 1771 10774
rect 1925 10826 1981 10828
rect 1925 10774 1927 10826
rect 1927 10774 1979 10826
rect 1979 10774 1981 10826
rect 1925 10772 1981 10774
rect 2136 10826 2192 10828
rect 2136 10774 2138 10826
rect 2138 10774 2190 10826
rect 2190 10774 2192 10826
rect 2136 10772 2192 10774
rect 2347 10826 2403 10828
rect 2347 10774 2349 10826
rect 2349 10774 2401 10826
rect 2401 10774 2403 10826
rect 2347 10772 2403 10774
rect 2652 10339 2708 10395
rect 2832 10339 2888 10395
rect 3414 10332 3470 10388
rect 3594 10332 3650 10388
rect 3879 9872 3935 9928
rect 4090 9872 4146 9928
rect 4302 9926 4358 9928
rect 4513 9926 4569 9928
rect 4302 9874 4352 9926
rect 4352 9874 4358 9926
rect 4513 9874 4532 9926
rect 4532 9874 4569 9926
rect 4302 9872 4358 9874
rect 4513 9872 4569 9874
rect 2652 9405 2708 9461
rect 2832 9405 2888 9461
rect 3414 9412 3470 9468
rect 3594 9412 3650 9468
rect 449 9026 505 9028
rect 449 8974 451 9026
rect 451 8974 503 9026
rect 503 8974 505 9026
rect 449 8972 505 8974
rect 660 9026 716 9028
rect 660 8974 662 9026
rect 662 8974 714 9026
rect 714 8974 716 9026
rect 660 8972 716 8974
rect 871 9026 927 9028
rect 871 8974 873 9026
rect 873 8974 925 9026
rect 925 8974 927 9026
rect 871 8972 927 8974
rect 1081 9026 1137 9028
rect 1081 8974 1083 9026
rect 1083 8974 1135 9026
rect 1135 8974 1137 9026
rect 1081 8972 1137 8974
rect 1292 9026 1348 9028
rect 1292 8974 1294 9026
rect 1294 8974 1346 9026
rect 1346 8974 1348 9026
rect 1292 8972 1348 8974
rect 1504 9026 1560 9028
rect 1504 8974 1506 9026
rect 1506 8974 1558 9026
rect 1558 8974 1560 9026
rect 1504 8972 1560 8974
rect 1715 9026 1771 9028
rect 1715 8974 1717 9026
rect 1717 8974 1769 9026
rect 1769 8974 1771 9026
rect 1715 8972 1771 8974
rect 1925 9026 1981 9028
rect 1925 8974 1927 9026
rect 1927 8974 1979 9026
rect 1979 8974 1981 9026
rect 1925 8972 1981 8974
rect 2136 9026 2192 9028
rect 2136 8974 2138 9026
rect 2138 8974 2190 9026
rect 2190 8974 2192 9026
rect 2136 8972 2192 8974
rect 2347 9026 2403 9028
rect 2347 8974 2349 9026
rect 2349 8974 2401 9026
rect 2401 8974 2403 9026
rect 2347 8972 2403 8974
rect 2652 8539 2708 8595
rect 2832 8539 2888 8595
rect 3414 8532 3470 8588
rect 3594 8532 3650 8588
rect 3879 8072 3935 8128
rect 4090 8072 4146 8128
rect 4302 8126 4358 8128
rect 4513 8126 4569 8128
rect 4302 8074 4352 8126
rect 4352 8074 4358 8126
rect 4513 8074 4532 8126
rect 4532 8074 4569 8126
rect 4302 8072 4358 8074
rect 4513 8072 4569 8074
rect 2652 7605 2708 7661
rect 2832 7605 2888 7661
rect 3414 7612 3470 7668
rect 3594 7612 3650 7668
rect 449 7226 505 7228
rect 449 7174 451 7226
rect 451 7174 503 7226
rect 503 7174 505 7226
rect 449 7172 505 7174
rect 660 7226 716 7228
rect 660 7174 662 7226
rect 662 7174 714 7226
rect 714 7174 716 7226
rect 660 7172 716 7174
rect 871 7226 927 7228
rect 871 7174 873 7226
rect 873 7174 925 7226
rect 925 7174 927 7226
rect 871 7172 927 7174
rect 1081 7226 1137 7228
rect 1081 7174 1083 7226
rect 1083 7174 1135 7226
rect 1135 7174 1137 7226
rect 1081 7172 1137 7174
rect 1292 7226 1348 7228
rect 1292 7174 1294 7226
rect 1294 7174 1346 7226
rect 1346 7174 1348 7226
rect 1292 7172 1348 7174
rect 1504 7226 1560 7228
rect 1504 7174 1506 7226
rect 1506 7174 1558 7226
rect 1558 7174 1560 7226
rect 1504 7172 1560 7174
rect 1715 7226 1771 7228
rect 1715 7174 1717 7226
rect 1717 7174 1769 7226
rect 1769 7174 1771 7226
rect 1715 7172 1771 7174
rect 1925 7226 1981 7228
rect 1925 7174 1927 7226
rect 1927 7174 1979 7226
rect 1979 7174 1981 7226
rect 1925 7172 1981 7174
rect 2136 7226 2192 7228
rect 2136 7174 2138 7226
rect 2138 7174 2190 7226
rect 2190 7174 2192 7226
rect 2136 7172 2192 7174
rect 2347 7226 2403 7228
rect 2347 7174 2349 7226
rect 2349 7174 2401 7226
rect 2401 7174 2403 7226
rect 2347 7172 2403 7174
rect 2652 6739 2708 6795
rect 2832 6739 2888 6795
rect 3414 6732 3470 6788
rect 3594 6732 3650 6788
rect 3879 6272 3935 6328
rect 4090 6272 4146 6328
rect 4302 6326 4358 6328
rect 4513 6326 4569 6328
rect 4302 6274 4352 6326
rect 4352 6274 4358 6326
rect 4513 6274 4532 6326
rect 4532 6274 4569 6326
rect 4302 6272 4358 6274
rect 4513 6272 4569 6274
rect 2652 5805 2708 5861
rect 2832 5805 2888 5861
rect 3414 5812 3470 5868
rect 3594 5812 3650 5868
rect 449 5426 505 5428
rect 449 5374 451 5426
rect 451 5374 503 5426
rect 503 5374 505 5426
rect 449 5372 505 5374
rect 660 5426 716 5428
rect 660 5374 662 5426
rect 662 5374 714 5426
rect 714 5374 716 5426
rect 660 5372 716 5374
rect 871 5426 927 5428
rect 871 5374 873 5426
rect 873 5374 925 5426
rect 925 5374 927 5426
rect 871 5372 927 5374
rect 1081 5426 1137 5428
rect 1081 5374 1083 5426
rect 1083 5374 1135 5426
rect 1135 5374 1137 5426
rect 1081 5372 1137 5374
rect 1292 5426 1348 5428
rect 1292 5374 1294 5426
rect 1294 5374 1346 5426
rect 1346 5374 1348 5426
rect 1292 5372 1348 5374
rect 1504 5426 1560 5428
rect 1504 5374 1506 5426
rect 1506 5374 1558 5426
rect 1558 5374 1560 5426
rect 1504 5372 1560 5374
rect 1715 5426 1771 5428
rect 1715 5374 1717 5426
rect 1717 5374 1769 5426
rect 1769 5374 1771 5426
rect 1715 5372 1771 5374
rect 1925 5426 1981 5428
rect 1925 5374 1927 5426
rect 1927 5374 1979 5426
rect 1979 5374 1981 5426
rect 1925 5372 1981 5374
rect 2136 5426 2192 5428
rect 2136 5374 2138 5426
rect 2138 5374 2190 5426
rect 2190 5374 2192 5426
rect 2136 5372 2192 5374
rect 2347 5426 2403 5428
rect 2347 5374 2349 5426
rect 2349 5374 2401 5426
rect 2401 5374 2403 5426
rect 2347 5372 2403 5374
rect 2652 4939 2708 4995
rect 2832 4939 2888 4995
rect 3414 4932 3470 4988
rect 3594 4932 3650 4988
rect 3879 4472 3935 4528
rect 4090 4472 4146 4528
rect 4302 4526 4358 4528
rect 4513 4526 4569 4528
rect 4302 4474 4352 4526
rect 4352 4474 4358 4526
rect 4513 4474 4532 4526
rect 4532 4474 4569 4526
rect 4302 4472 4358 4474
rect 4513 4472 4569 4474
rect 2652 4005 2708 4061
rect 2832 4005 2888 4061
rect 3414 4012 3470 4068
rect 3594 4012 3650 4068
rect 449 3626 505 3628
rect 449 3574 451 3626
rect 451 3574 503 3626
rect 503 3574 505 3626
rect 449 3572 505 3574
rect 660 3626 716 3628
rect 660 3574 662 3626
rect 662 3574 714 3626
rect 714 3574 716 3626
rect 660 3572 716 3574
rect 871 3626 927 3628
rect 871 3574 873 3626
rect 873 3574 925 3626
rect 925 3574 927 3626
rect 871 3572 927 3574
rect 1081 3626 1137 3628
rect 1081 3574 1083 3626
rect 1083 3574 1135 3626
rect 1135 3574 1137 3626
rect 1081 3572 1137 3574
rect 1292 3626 1348 3628
rect 1292 3574 1294 3626
rect 1294 3574 1346 3626
rect 1346 3574 1348 3626
rect 1292 3572 1348 3574
rect 1504 3626 1560 3628
rect 1504 3574 1506 3626
rect 1506 3574 1558 3626
rect 1558 3574 1560 3626
rect 1504 3572 1560 3574
rect 1715 3626 1771 3628
rect 1715 3574 1717 3626
rect 1717 3574 1769 3626
rect 1769 3574 1771 3626
rect 1715 3572 1771 3574
rect 1925 3626 1981 3628
rect 1925 3574 1927 3626
rect 1927 3574 1979 3626
rect 1979 3574 1981 3626
rect 1925 3572 1981 3574
rect 2136 3626 2192 3628
rect 2136 3574 2138 3626
rect 2138 3574 2190 3626
rect 2190 3574 2192 3626
rect 2136 3572 2192 3574
rect 2347 3626 2403 3628
rect 2347 3574 2349 3626
rect 2349 3574 2401 3626
rect 2401 3574 2403 3626
rect 2347 3572 2403 3574
rect 2652 3139 2708 3195
rect 2832 3139 2888 3195
rect 3414 3132 3470 3188
rect 3594 3132 3650 3188
rect 3879 2672 3935 2728
rect 4090 2672 4146 2728
rect 4302 2726 4358 2728
rect 4513 2726 4569 2728
rect 4302 2674 4352 2726
rect 4352 2674 4358 2726
rect 4513 2674 4532 2726
rect 4532 2674 4569 2726
rect 4302 2672 4358 2674
rect 4513 2672 4569 2674
rect 2652 2205 2708 2261
rect 2832 2205 2888 2261
rect 3414 2212 3470 2268
rect 3594 2212 3650 2268
rect 449 1826 505 1828
rect 449 1774 451 1826
rect 451 1774 503 1826
rect 503 1774 505 1826
rect 449 1772 505 1774
rect 660 1826 716 1828
rect 660 1774 662 1826
rect 662 1774 714 1826
rect 714 1774 716 1826
rect 660 1772 716 1774
rect 871 1826 927 1828
rect 871 1774 873 1826
rect 873 1774 925 1826
rect 925 1774 927 1826
rect 871 1772 927 1774
rect 1081 1826 1137 1828
rect 1081 1774 1083 1826
rect 1083 1774 1135 1826
rect 1135 1774 1137 1826
rect 1081 1772 1137 1774
rect 1292 1826 1348 1828
rect 1292 1774 1294 1826
rect 1294 1774 1346 1826
rect 1346 1774 1348 1826
rect 1292 1772 1348 1774
rect 1504 1826 1560 1828
rect 1504 1774 1506 1826
rect 1506 1774 1558 1826
rect 1558 1774 1560 1826
rect 1504 1772 1560 1774
rect 1715 1826 1771 1828
rect 1715 1774 1717 1826
rect 1717 1774 1769 1826
rect 1769 1774 1771 1826
rect 1715 1772 1771 1774
rect 1925 1826 1981 1828
rect 1925 1774 1927 1826
rect 1927 1774 1979 1826
rect 1979 1774 1981 1826
rect 1925 1772 1981 1774
rect 2136 1826 2192 1828
rect 2136 1774 2138 1826
rect 2138 1774 2190 1826
rect 2190 1774 2192 1826
rect 2136 1772 2192 1774
rect 2347 1826 2403 1828
rect 2347 1774 2349 1826
rect 2349 1774 2401 1826
rect 2401 1774 2403 1826
rect 2347 1772 2403 1774
rect 2652 1339 2708 1395
rect 2832 1339 2888 1395
rect 3414 1332 3470 1388
rect 3594 1332 3650 1388
rect 3879 872 3935 928
rect 4090 872 4146 928
rect 4302 926 4358 928
rect 4513 926 4569 928
rect 4302 874 4352 926
rect 4352 874 4358 926
rect 4513 874 4532 926
rect 4532 874 4569 926
rect 4302 872 4358 874
rect 4513 872 4569 874
rect 2652 405 2708 461
rect 2832 405 2888 461
rect 3414 412 3470 468
rect 3594 412 3650 468
rect 449 26 505 28
rect 449 -26 451 26
rect 451 -26 503 26
rect 503 -26 505 26
rect 449 -28 505 -26
rect 660 26 716 28
rect 660 -26 662 26
rect 662 -26 714 26
rect 714 -26 716 26
rect 660 -28 716 -26
rect 871 26 927 28
rect 871 -26 873 26
rect 873 -26 925 26
rect 925 -26 927 26
rect 871 -28 927 -26
rect 1081 26 1137 28
rect 1081 -26 1083 26
rect 1083 -26 1135 26
rect 1135 -26 1137 26
rect 1081 -28 1137 -26
rect 1292 26 1348 28
rect 1292 -26 1294 26
rect 1294 -26 1346 26
rect 1346 -26 1348 26
rect 1292 -28 1348 -26
rect 1504 26 1560 28
rect 1504 -26 1506 26
rect 1506 -26 1558 26
rect 1558 -26 1560 26
rect 1504 -28 1560 -26
rect 1715 26 1771 28
rect 1715 -26 1717 26
rect 1717 -26 1769 26
rect 1769 -26 1771 26
rect 1715 -28 1771 -26
rect 1925 26 1981 28
rect 1925 -26 1927 26
rect 1927 -26 1979 26
rect 1979 -26 1981 26
rect 1925 -28 1981 -26
rect 2136 26 2192 28
rect 2136 -26 2138 26
rect 2138 -26 2190 26
rect 2190 -26 2192 26
rect 2136 -28 2192 -26
rect 2347 26 2403 28
rect 2347 -26 2349 26
rect 2349 -26 2401 26
rect 2401 -26 2403 26
rect 2347 -28 2403 -26
rect 4815 14426 4871 14428
rect 4815 14374 4817 14426
rect 4817 14374 4869 14426
rect 4869 14374 4871 14426
rect 4815 14372 4871 14374
rect 5025 14426 5081 14428
rect 5025 14374 5027 14426
rect 5027 14374 5079 14426
rect 5079 14374 5081 14426
rect 5025 14372 5081 14374
rect 5236 14426 5292 14428
rect 5236 14374 5238 14426
rect 5238 14374 5290 14426
rect 5290 14374 5292 14426
rect 5236 14372 5292 14374
rect 5448 14426 5504 14428
rect 5448 14374 5450 14426
rect 5450 14374 5502 14426
rect 5502 14374 5504 14426
rect 5448 14372 5504 14374
rect 5659 14426 5715 14428
rect 5659 14374 5661 14426
rect 5661 14374 5713 14426
rect 5713 14374 5715 14426
rect 5659 14372 5715 14374
rect 5869 14426 5925 14428
rect 5869 14374 5871 14426
rect 5871 14374 5923 14426
rect 5923 14374 5925 14426
rect 5869 14372 5925 14374
rect 6273 13980 6329 14036
rect 6273 12964 6329 13020
rect 7486 13749 7542 13805
rect 7666 13749 7722 13805
rect 7925 13472 7981 13528
rect 8136 13472 8192 13528
rect 8347 13472 8403 13528
rect 4815 12626 4871 12628
rect 4815 12574 4817 12626
rect 4817 12574 4869 12626
rect 4869 12574 4871 12626
rect 4815 12572 4871 12574
rect 5025 12626 5081 12628
rect 5025 12574 5027 12626
rect 5027 12574 5079 12626
rect 5079 12574 5081 12626
rect 5025 12572 5081 12574
rect 5236 12626 5292 12628
rect 5236 12574 5238 12626
rect 5238 12574 5290 12626
rect 5290 12574 5292 12626
rect 5236 12572 5292 12574
rect 5448 12626 5504 12628
rect 5448 12574 5450 12626
rect 5450 12574 5502 12626
rect 5502 12574 5504 12626
rect 5448 12572 5504 12574
rect 5659 12626 5715 12628
rect 5659 12574 5661 12626
rect 5661 12574 5713 12626
rect 5713 12574 5715 12626
rect 5659 12572 5715 12574
rect 5869 12626 5925 12628
rect 5869 12574 5871 12626
rect 5871 12574 5923 12626
rect 5923 12574 5925 12626
rect 5869 12572 5925 12574
rect 6273 12180 6329 12236
rect 7486 13195 7542 13251
rect 7666 13195 7722 13251
rect 6273 11164 6329 11220
rect 7486 11949 7542 12005
rect 7666 11949 7722 12005
rect 7925 11672 7981 11728
rect 8136 11672 8192 11728
rect 8347 11672 8403 11728
rect 4815 10826 4871 10828
rect 4815 10774 4817 10826
rect 4817 10774 4869 10826
rect 4869 10774 4871 10826
rect 4815 10772 4871 10774
rect 5025 10826 5081 10828
rect 5025 10774 5027 10826
rect 5027 10774 5079 10826
rect 5079 10774 5081 10826
rect 5025 10772 5081 10774
rect 5236 10826 5292 10828
rect 5236 10774 5238 10826
rect 5238 10774 5290 10826
rect 5290 10774 5292 10826
rect 5236 10772 5292 10774
rect 5448 10826 5504 10828
rect 5448 10774 5450 10826
rect 5450 10774 5502 10826
rect 5502 10774 5504 10826
rect 5448 10772 5504 10774
rect 5659 10826 5715 10828
rect 5659 10774 5661 10826
rect 5661 10774 5713 10826
rect 5713 10774 5715 10826
rect 5659 10772 5715 10774
rect 5869 10826 5925 10828
rect 5869 10774 5871 10826
rect 5871 10774 5923 10826
rect 5923 10774 5925 10826
rect 5869 10772 5925 10774
rect 6273 10380 6329 10436
rect 7486 11395 7542 11451
rect 7666 11395 7722 11451
rect 6273 9364 6329 9420
rect 7486 10149 7542 10205
rect 7666 10149 7722 10205
rect 7925 9872 7981 9928
rect 8136 9872 8192 9928
rect 8347 9872 8403 9928
rect 4815 9026 4871 9028
rect 4815 8974 4817 9026
rect 4817 8974 4869 9026
rect 4869 8974 4871 9026
rect 4815 8972 4871 8974
rect 5025 9026 5081 9028
rect 5025 8974 5027 9026
rect 5027 8974 5079 9026
rect 5079 8974 5081 9026
rect 5025 8972 5081 8974
rect 5236 9026 5292 9028
rect 5236 8974 5238 9026
rect 5238 8974 5290 9026
rect 5290 8974 5292 9026
rect 5236 8972 5292 8974
rect 5448 9026 5504 9028
rect 5448 8974 5450 9026
rect 5450 8974 5502 9026
rect 5502 8974 5504 9026
rect 5448 8972 5504 8974
rect 5659 9026 5715 9028
rect 5659 8974 5661 9026
rect 5661 8974 5713 9026
rect 5713 8974 5715 9026
rect 5659 8972 5715 8974
rect 5869 9026 5925 9028
rect 5869 8974 5871 9026
rect 5871 8974 5923 9026
rect 5923 8974 5925 9026
rect 5869 8972 5925 8974
rect 6273 8580 6329 8636
rect 7486 9595 7542 9651
rect 7666 9595 7722 9651
rect 6273 7564 6329 7620
rect 7486 8349 7542 8405
rect 7666 8349 7722 8405
rect 7925 8072 7981 8128
rect 8136 8072 8192 8128
rect 8347 8072 8403 8128
rect 4815 7226 4871 7228
rect 4815 7174 4817 7226
rect 4817 7174 4869 7226
rect 4869 7174 4871 7226
rect 4815 7172 4871 7174
rect 5025 7226 5081 7228
rect 5025 7174 5027 7226
rect 5027 7174 5079 7226
rect 5079 7174 5081 7226
rect 5025 7172 5081 7174
rect 5236 7226 5292 7228
rect 5236 7174 5238 7226
rect 5238 7174 5290 7226
rect 5290 7174 5292 7226
rect 5236 7172 5292 7174
rect 5448 7226 5504 7228
rect 5448 7174 5450 7226
rect 5450 7174 5502 7226
rect 5502 7174 5504 7226
rect 5448 7172 5504 7174
rect 5659 7226 5715 7228
rect 5659 7174 5661 7226
rect 5661 7174 5713 7226
rect 5713 7174 5715 7226
rect 5659 7172 5715 7174
rect 5869 7226 5925 7228
rect 5869 7174 5871 7226
rect 5871 7174 5923 7226
rect 5923 7174 5925 7226
rect 5869 7172 5925 7174
rect 6273 6780 6329 6836
rect 7486 7795 7542 7851
rect 7666 7795 7722 7851
rect 6273 5764 6329 5820
rect 7486 6549 7542 6605
rect 7666 6549 7722 6605
rect 7925 6272 7981 6328
rect 8136 6272 8192 6328
rect 8347 6272 8403 6328
rect 4815 5426 4871 5428
rect 4815 5374 4817 5426
rect 4817 5374 4869 5426
rect 4869 5374 4871 5426
rect 4815 5372 4871 5374
rect 5025 5426 5081 5428
rect 5025 5374 5027 5426
rect 5027 5374 5079 5426
rect 5079 5374 5081 5426
rect 5025 5372 5081 5374
rect 5236 5426 5292 5428
rect 5236 5374 5238 5426
rect 5238 5374 5290 5426
rect 5290 5374 5292 5426
rect 5236 5372 5292 5374
rect 5448 5426 5504 5428
rect 5448 5374 5450 5426
rect 5450 5374 5502 5426
rect 5502 5374 5504 5426
rect 5448 5372 5504 5374
rect 5659 5426 5715 5428
rect 5659 5374 5661 5426
rect 5661 5374 5713 5426
rect 5713 5374 5715 5426
rect 5659 5372 5715 5374
rect 5869 5426 5925 5428
rect 5869 5374 5871 5426
rect 5871 5374 5923 5426
rect 5923 5374 5925 5426
rect 5869 5372 5925 5374
rect 6273 4980 6329 5036
rect 7486 5995 7542 6051
rect 7666 5995 7722 6051
rect 6273 3964 6329 4020
rect 7486 4749 7542 4805
rect 7666 4749 7722 4805
rect 7925 4472 7981 4528
rect 8136 4472 8192 4528
rect 8347 4472 8403 4528
rect 4815 3626 4871 3628
rect 4815 3574 4817 3626
rect 4817 3574 4869 3626
rect 4869 3574 4871 3626
rect 4815 3572 4871 3574
rect 5025 3626 5081 3628
rect 5025 3574 5027 3626
rect 5027 3574 5079 3626
rect 5079 3574 5081 3626
rect 5025 3572 5081 3574
rect 5236 3626 5292 3628
rect 5236 3574 5238 3626
rect 5238 3574 5290 3626
rect 5290 3574 5292 3626
rect 5236 3572 5292 3574
rect 5448 3626 5504 3628
rect 5448 3574 5450 3626
rect 5450 3574 5502 3626
rect 5502 3574 5504 3626
rect 5448 3572 5504 3574
rect 5659 3626 5715 3628
rect 5659 3574 5661 3626
rect 5661 3574 5713 3626
rect 5713 3574 5715 3626
rect 5659 3572 5715 3574
rect 5869 3626 5925 3628
rect 5869 3574 5871 3626
rect 5871 3574 5923 3626
rect 5923 3574 5925 3626
rect 5869 3572 5925 3574
rect 6273 3180 6329 3236
rect 7486 4195 7542 4251
rect 7666 4195 7722 4251
rect 6273 2164 6329 2220
rect 7486 2949 7542 3005
rect 7666 2949 7722 3005
rect 7925 2672 7981 2728
rect 8136 2672 8192 2728
rect 8347 2672 8403 2728
rect 4815 1826 4871 1828
rect 4815 1774 4817 1826
rect 4817 1774 4869 1826
rect 4869 1774 4871 1826
rect 4815 1772 4871 1774
rect 5025 1826 5081 1828
rect 5025 1774 5027 1826
rect 5027 1774 5079 1826
rect 5079 1774 5081 1826
rect 5025 1772 5081 1774
rect 5236 1826 5292 1828
rect 5236 1774 5238 1826
rect 5238 1774 5290 1826
rect 5290 1774 5292 1826
rect 5236 1772 5292 1774
rect 5448 1826 5504 1828
rect 5448 1774 5450 1826
rect 5450 1774 5502 1826
rect 5502 1774 5504 1826
rect 5448 1772 5504 1774
rect 5659 1826 5715 1828
rect 5659 1774 5661 1826
rect 5661 1774 5713 1826
rect 5713 1774 5715 1826
rect 5659 1772 5715 1774
rect 5869 1826 5925 1828
rect 5869 1774 5871 1826
rect 5871 1774 5923 1826
rect 5923 1774 5925 1826
rect 5869 1772 5925 1774
rect 6273 1380 6329 1436
rect 7486 2395 7542 2451
rect 7666 2395 7722 2451
rect 6273 364 6329 420
rect 7486 1149 7542 1205
rect 7666 1149 7722 1205
rect 7925 872 7981 928
rect 8136 872 8192 928
rect 8347 872 8403 928
rect 4815 26 4871 28
rect 4815 -26 4817 26
rect 4817 -26 4869 26
rect 4869 -26 4871 26
rect 4815 -28 4871 -26
rect 5025 26 5081 28
rect 5025 -26 5027 26
rect 5027 -26 5079 26
rect 5079 -26 5081 26
rect 5025 -28 5081 -26
rect 5236 26 5292 28
rect 5236 -26 5238 26
rect 5238 -26 5290 26
rect 5290 -26 5292 26
rect 5236 -28 5292 -26
rect 5448 26 5504 28
rect 5448 -26 5450 26
rect 5450 -26 5502 26
rect 5502 -26 5504 26
rect 5448 -28 5504 -26
rect 5659 26 5715 28
rect 5659 -26 5661 26
rect 5661 -26 5713 26
rect 5713 -26 5715 26
rect 5659 -28 5715 -26
rect 5869 26 5925 28
rect 5869 -26 5871 26
rect 5871 -26 5923 26
rect 5923 -26 5925 26
rect 5869 -28 5925 -26
rect 7486 595 7542 651
rect 7666 595 7722 651
rect 8647 14426 8703 14428
rect 8647 14374 8649 14426
rect 8649 14374 8701 14426
rect 8701 14374 8703 14426
rect 8647 14372 8703 14374
rect 8827 14426 8883 14428
rect 8827 14374 8829 14426
rect 8829 14374 8881 14426
rect 8881 14374 8883 14426
rect 8827 14372 8883 14374
rect 9370 13749 9426 13805
rect 9589 13980 9645 14036
rect 9848 13472 9904 13528
rect 10028 13472 10084 13528
rect 9370 13195 9426 13251
rect 9589 12964 9645 13020
rect 8647 12626 8703 12628
rect 8647 12574 8649 12626
rect 8649 12574 8701 12626
rect 8701 12574 8703 12626
rect 8647 12572 8703 12574
rect 8827 12626 8883 12628
rect 8827 12574 8829 12626
rect 8829 12574 8881 12626
rect 8881 12574 8883 12626
rect 8827 12572 8883 12574
rect 9370 11949 9426 12005
rect 9589 12180 9645 12236
rect 9848 11672 9904 11728
rect 10028 11672 10084 11728
rect 9370 11395 9426 11451
rect 9589 11164 9645 11220
rect 8647 10826 8703 10828
rect 8647 10774 8649 10826
rect 8649 10774 8701 10826
rect 8701 10774 8703 10826
rect 8647 10772 8703 10774
rect 8827 10826 8883 10828
rect 8827 10774 8829 10826
rect 8829 10774 8881 10826
rect 8881 10774 8883 10826
rect 8827 10772 8883 10774
rect 9370 10149 9426 10205
rect 9589 10380 9645 10436
rect 9848 9872 9904 9928
rect 10028 9872 10084 9928
rect 9370 9595 9426 9651
rect 9589 9364 9645 9420
rect 8647 9026 8703 9028
rect 8647 8974 8649 9026
rect 8649 8974 8701 9026
rect 8701 8974 8703 9026
rect 8647 8972 8703 8974
rect 8827 9026 8883 9028
rect 8827 8974 8829 9026
rect 8829 8974 8881 9026
rect 8881 8974 8883 9026
rect 8827 8972 8883 8974
rect 9370 8349 9426 8405
rect 9589 8580 9645 8636
rect 9848 8072 9904 8128
rect 10028 8072 10084 8128
rect 9370 7795 9426 7851
rect 9589 7564 9645 7620
rect 8647 7226 8703 7228
rect 8647 7174 8649 7226
rect 8649 7174 8701 7226
rect 8701 7174 8703 7226
rect 8647 7172 8703 7174
rect 8827 7226 8883 7228
rect 8827 7174 8829 7226
rect 8829 7174 8881 7226
rect 8881 7174 8883 7226
rect 8827 7172 8883 7174
rect 9370 6549 9426 6605
rect 9589 6780 9645 6836
rect 9848 6272 9904 6328
rect 10028 6272 10084 6328
rect 9370 5995 9426 6051
rect 9589 5764 9645 5820
rect 8647 5426 8703 5428
rect 8647 5374 8649 5426
rect 8649 5374 8701 5426
rect 8701 5374 8703 5426
rect 8647 5372 8703 5374
rect 8827 5426 8883 5428
rect 8827 5374 8829 5426
rect 8829 5374 8881 5426
rect 8881 5374 8883 5426
rect 8827 5372 8883 5374
rect 9370 4749 9426 4805
rect 9589 4980 9645 5036
rect 9848 4472 9904 4528
rect 10028 4472 10084 4528
rect 9370 4195 9426 4251
rect 9589 3964 9645 4020
rect 8647 3626 8703 3628
rect 8647 3574 8649 3626
rect 8649 3574 8701 3626
rect 8701 3574 8703 3626
rect 8647 3572 8703 3574
rect 8827 3626 8883 3628
rect 8827 3574 8829 3626
rect 8829 3574 8881 3626
rect 8881 3574 8883 3626
rect 8827 3572 8883 3574
rect 9370 2949 9426 3005
rect 9589 3180 9645 3236
rect 9848 2672 9904 2728
rect 10028 2672 10084 2728
rect 9370 2395 9426 2451
rect 9589 2164 9645 2220
rect 8647 1826 8703 1828
rect 8647 1774 8649 1826
rect 8649 1774 8701 1826
rect 8701 1774 8703 1826
rect 8647 1772 8703 1774
rect 8827 1826 8883 1828
rect 8827 1774 8829 1826
rect 8829 1774 8881 1826
rect 8881 1774 8883 1826
rect 8827 1772 8883 1774
rect 9370 1149 9426 1205
rect 9589 1380 9645 1436
rect 9848 872 9904 928
rect 10028 872 10084 928
rect 9370 595 9426 651
rect 9589 364 9645 420
rect 8647 26 8703 28
rect 8647 -26 8649 26
rect 8649 -26 8701 26
rect 8701 -26 8703 26
rect 8647 -28 8703 -26
rect 8827 26 8883 28
rect 8827 -26 8829 26
rect 8829 -26 8881 26
rect 8881 -26 8883 26
rect 8827 -28 8883 -26
rect 13385 13472 13441 13528
rect 13596 13472 13652 13528
rect 13808 13472 13864 13528
rect 14019 13472 14075 13528
rect 13385 11672 13441 11728
rect 13596 11672 13652 11728
rect 13808 11672 13864 11728
rect 14019 11672 14075 11728
rect 13385 9872 13441 9928
rect 13596 9872 13652 9928
rect 13808 9872 13864 9928
rect 14019 9872 14075 9928
rect 13385 8072 13441 8128
rect 13596 8072 13652 8128
rect 13808 8072 13864 8128
rect 14019 8072 14075 8128
rect 13385 6272 13441 6328
rect 13596 6272 13652 6328
rect 13808 6272 13864 6328
rect 14019 6272 14075 6328
rect 13385 4472 13441 4528
rect 13596 4472 13652 4528
rect 13808 4472 13864 4528
rect 14019 4472 14075 4528
rect 13385 2672 13441 2728
rect 13596 2672 13652 2728
rect 13808 2672 13864 2728
rect 14019 2672 14075 2728
rect 13385 872 13441 928
rect 13596 872 13652 928
rect 13808 872 13864 928
rect 14019 872 14075 928
rect 14429 14426 14485 14428
rect 14429 14374 14431 14426
rect 14431 14374 14483 14426
rect 14483 14374 14485 14426
rect 14429 14372 14485 14374
rect 14640 14426 14696 14428
rect 14640 14374 14642 14426
rect 14642 14374 14694 14426
rect 14694 14374 14696 14426
rect 14640 14372 14696 14374
rect 14851 14426 14907 14428
rect 14851 14374 14853 14426
rect 14853 14374 14905 14426
rect 14905 14374 14907 14426
rect 14851 14372 14907 14374
rect 14429 12626 14485 12628
rect 14429 12574 14431 12626
rect 14431 12574 14483 12626
rect 14483 12574 14485 12626
rect 14429 12572 14485 12574
rect 14640 12626 14696 12628
rect 14640 12574 14642 12626
rect 14642 12574 14694 12626
rect 14694 12574 14696 12626
rect 14640 12572 14696 12574
rect 14851 12626 14907 12628
rect 14851 12574 14853 12626
rect 14853 12574 14905 12626
rect 14905 12574 14907 12626
rect 14851 12572 14907 12574
rect 14429 10826 14485 10828
rect 14429 10774 14431 10826
rect 14431 10774 14483 10826
rect 14483 10774 14485 10826
rect 14429 10772 14485 10774
rect 14640 10826 14696 10828
rect 14640 10774 14642 10826
rect 14642 10774 14694 10826
rect 14694 10774 14696 10826
rect 14640 10772 14696 10774
rect 14851 10826 14907 10828
rect 14851 10774 14853 10826
rect 14853 10774 14905 10826
rect 14905 10774 14907 10826
rect 14851 10772 14907 10774
rect 14429 9026 14485 9028
rect 14429 8974 14431 9026
rect 14431 8974 14483 9026
rect 14483 8974 14485 9026
rect 14429 8972 14485 8974
rect 14640 9026 14696 9028
rect 14640 8974 14642 9026
rect 14642 8974 14694 9026
rect 14694 8974 14696 9026
rect 14640 8972 14696 8974
rect 14851 9026 14907 9028
rect 14851 8974 14853 9026
rect 14853 8974 14905 9026
rect 14905 8974 14907 9026
rect 14851 8972 14907 8974
rect 14429 7226 14485 7228
rect 14429 7174 14431 7226
rect 14431 7174 14483 7226
rect 14483 7174 14485 7226
rect 14429 7172 14485 7174
rect 14640 7226 14696 7228
rect 14640 7174 14642 7226
rect 14642 7174 14694 7226
rect 14694 7174 14696 7226
rect 14640 7172 14696 7174
rect 14851 7226 14907 7228
rect 14851 7174 14853 7226
rect 14853 7174 14905 7226
rect 14905 7174 14907 7226
rect 14851 7172 14907 7174
rect 14429 5426 14485 5428
rect 14429 5374 14431 5426
rect 14431 5374 14483 5426
rect 14483 5374 14485 5426
rect 14429 5372 14485 5374
rect 14640 5426 14696 5428
rect 14640 5374 14642 5426
rect 14642 5374 14694 5426
rect 14694 5374 14696 5426
rect 14640 5372 14696 5374
rect 14851 5426 14907 5428
rect 14851 5374 14853 5426
rect 14853 5374 14905 5426
rect 14905 5374 14907 5426
rect 14851 5372 14907 5374
rect 14429 3626 14485 3628
rect 14429 3574 14431 3626
rect 14431 3574 14483 3626
rect 14483 3574 14485 3626
rect 14429 3572 14485 3574
rect 14640 3626 14696 3628
rect 14640 3574 14642 3626
rect 14642 3574 14694 3626
rect 14694 3574 14696 3626
rect 14640 3572 14696 3574
rect 14851 3626 14907 3628
rect 14851 3574 14853 3626
rect 14853 3574 14905 3626
rect 14905 3574 14907 3626
rect 14851 3572 14907 3574
rect 14429 1826 14485 1828
rect 14429 1774 14431 1826
rect 14431 1774 14483 1826
rect 14483 1774 14485 1826
rect 14429 1772 14485 1774
rect 14640 1826 14696 1828
rect 14640 1774 14642 1826
rect 14642 1774 14694 1826
rect 14694 1774 14696 1826
rect 14640 1772 14696 1774
rect 14851 1826 14907 1828
rect 14851 1774 14853 1826
rect 14853 1774 14905 1826
rect 14905 1774 14907 1826
rect 14851 1772 14907 1774
rect 14429 26 14485 28
rect 14429 -26 14431 26
rect 14431 -26 14483 26
rect 14483 -26 14485 26
rect 14429 -28 14485 -26
rect 14640 26 14696 28
rect 14640 -26 14642 26
rect 14642 -26 14694 26
rect 14694 -26 14696 26
rect 14640 -28 14696 -26
rect 14851 26 14907 28
rect 14851 -26 14853 26
rect 14853 -26 14905 26
rect 14905 -26 14907 26
rect 14851 -28 14907 -26
rect 18433 14426 18489 14428
rect 18433 14374 18435 14426
rect 18435 14374 18487 14426
rect 18487 14374 18489 14426
rect 18433 14372 18489 14374
rect 18643 14426 18699 14428
rect 18643 14374 18645 14426
rect 18645 14374 18697 14426
rect 18697 14374 18699 14426
rect 18643 14372 18699 14374
rect 18854 14426 18910 14428
rect 18854 14374 18856 14426
rect 18856 14374 18908 14426
rect 18908 14374 18910 14426
rect 18854 14372 18910 14374
rect 19066 14426 19122 14428
rect 19066 14374 19068 14426
rect 19068 14374 19120 14426
rect 19120 14374 19122 14426
rect 19066 14372 19122 14374
rect 19277 14426 19333 14428
rect 19277 14374 19279 14426
rect 19279 14374 19331 14426
rect 19331 14374 19333 14426
rect 19277 14372 19333 14374
rect 19487 14426 19543 14428
rect 19487 14374 19489 14426
rect 19489 14374 19541 14426
rect 19541 14374 19543 14426
rect 19487 14372 19543 14374
rect 18191 14020 18247 14022
rect 18191 13968 18193 14020
rect 18193 13968 18245 14020
rect 18245 13968 18247 14020
rect 18191 13966 18247 13968
rect 18191 13802 18247 13804
rect 18191 13750 18193 13802
rect 18193 13750 18245 13802
rect 18245 13750 18247 13802
rect 18191 13748 18247 13750
rect 18191 13250 18247 13252
rect 18191 13198 18193 13250
rect 18193 13198 18245 13250
rect 18245 13198 18247 13250
rect 18191 13196 18247 13198
rect 18191 13032 18247 13034
rect 18191 12980 18193 13032
rect 18193 12980 18245 13032
rect 18245 12980 18247 13032
rect 18191 12978 18247 12980
rect 18433 12626 18489 12628
rect 18433 12574 18435 12626
rect 18435 12574 18487 12626
rect 18487 12574 18489 12626
rect 18433 12572 18489 12574
rect 18643 12626 18699 12628
rect 18643 12574 18645 12626
rect 18645 12574 18697 12626
rect 18697 12574 18699 12626
rect 18643 12572 18699 12574
rect 18854 12626 18910 12628
rect 18854 12574 18856 12626
rect 18856 12574 18908 12626
rect 18908 12574 18910 12626
rect 18854 12572 18910 12574
rect 19066 12626 19122 12628
rect 19066 12574 19068 12626
rect 19068 12574 19120 12626
rect 19120 12574 19122 12626
rect 19066 12572 19122 12574
rect 19277 12626 19333 12628
rect 19277 12574 19279 12626
rect 19279 12574 19331 12626
rect 19331 12574 19333 12626
rect 19277 12572 19333 12574
rect 19487 12626 19543 12628
rect 19487 12574 19489 12626
rect 19489 12574 19541 12626
rect 19541 12574 19543 12626
rect 19487 12572 19543 12574
rect 18191 12220 18247 12222
rect 18191 12168 18193 12220
rect 18193 12168 18245 12220
rect 18245 12168 18247 12220
rect 18191 12166 18247 12168
rect 18191 12002 18247 12004
rect 18191 11950 18193 12002
rect 18193 11950 18245 12002
rect 18245 11950 18247 12002
rect 18191 11948 18247 11950
rect 18191 11450 18247 11452
rect 18191 11398 18193 11450
rect 18193 11398 18245 11450
rect 18245 11398 18247 11450
rect 18191 11396 18247 11398
rect 18191 11232 18247 11234
rect 18191 11180 18193 11232
rect 18193 11180 18245 11232
rect 18245 11180 18247 11232
rect 18191 11178 18247 11180
rect 18433 10826 18489 10828
rect 18433 10774 18435 10826
rect 18435 10774 18487 10826
rect 18487 10774 18489 10826
rect 18433 10772 18489 10774
rect 18643 10826 18699 10828
rect 18643 10774 18645 10826
rect 18645 10774 18697 10826
rect 18697 10774 18699 10826
rect 18643 10772 18699 10774
rect 18854 10826 18910 10828
rect 18854 10774 18856 10826
rect 18856 10774 18908 10826
rect 18908 10774 18910 10826
rect 18854 10772 18910 10774
rect 19066 10826 19122 10828
rect 19066 10774 19068 10826
rect 19068 10774 19120 10826
rect 19120 10774 19122 10826
rect 19066 10772 19122 10774
rect 19277 10826 19333 10828
rect 19277 10774 19279 10826
rect 19279 10774 19331 10826
rect 19331 10774 19333 10826
rect 19277 10772 19333 10774
rect 19487 10826 19543 10828
rect 19487 10774 19489 10826
rect 19489 10774 19541 10826
rect 19541 10774 19543 10826
rect 19487 10772 19543 10774
rect 18191 10420 18247 10422
rect 18191 10368 18193 10420
rect 18193 10368 18245 10420
rect 18245 10368 18247 10420
rect 18191 10366 18247 10368
rect 18191 10202 18247 10204
rect 18191 10150 18193 10202
rect 18193 10150 18245 10202
rect 18245 10150 18247 10202
rect 18191 10148 18247 10150
rect 18191 9650 18247 9652
rect 18191 9598 18193 9650
rect 18193 9598 18245 9650
rect 18245 9598 18247 9650
rect 18191 9596 18247 9598
rect 18191 9432 18247 9434
rect 18191 9380 18193 9432
rect 18193 9380 18245 9432
rect 18245 9380 18247 9432
rect 18191 9378 18247 9380
rect 18433 9026 18489 9028
rect 18433 8974 18435 9026
rect 18435 8974 18487 9026
rect 18487 8974 18489 9026
rect 18433 8972 18489 8974
rect 18643 9026 18699 9028
rect 18643 8974 18645 9026
rect 18645 8974 18697 9026
rect 18697 8974 18699 9026
rect 18643 8972 18699 8974
rect 18854 9026 18910 9028
rect 18854 8974 18856 9026
rect 18856 8974 18908 9026
rect 18908 8974 18910 9026
rect 18854 8972 18910 8974
rect 19066 9026 19122 9028
rect 19066 8974 19068 9026
rect 19068 8974 19120 9026
rect 19120 8974 19122 9026
rect 19066 8972 19122 8974
rect 19277 9026 19333 9028
rect 19277 8974 19279 9026
rect 19279 8974 19331 9026
rect 19331 8974 19333 9026
rect 19277 8972 19333 8974
rect 19487 9026 19543 9028
rect 19487 8974 19489 9026
rect 19489 8974 19541 9026
rect 19541 8974 19543 9026
rect 19487 8972 19543 8974
rect 18191 8620 18247 8622
rect 18191 8568 18193 8620
rect 18193 8568 18245 8620
rect 18245 8568 18247 8620
rect 18191 8566 18247 8568
rect 18191 8402 18247 8404
rect 18191 8350 18193 8402
rect 18193 8350 18245 8402
rect 18245 8350 18247 8402
rect 18191 8348 18247 8350
rect 18191 7850 18247 7852
rect 18191 7798 18193 7850
rect 18193 7798 18245 7850
rect 18245 7798 18247 7850
rect 18191 7796 18247 7798
rect 18191 7632 18247 7634
rect 18191 7580 18193 7632
rect 18193 7580 18245 7632
rect 18245 7580 18247 7632
rect 18191 7578 18247 7580
rect 18433 7226 18489 7228
rect 18433 7174 18435 7226
rect 18435 7174 18487 7226
rect 18487 7174 18489 7226
rect 18433 7172 18489 7174
rect 18643 7226 18699 7228
rect 18643 7174 18645 7226
rect 18645 7174 18697 7226
rect 18697 7174 18699 7226
rect 18643 7172 18699 7174
rect 18854 7226 18910 7228
rect 18854 7174 18856 7226
rect 18856 7174 18908 7226
rect 18908 7174 18910 7226
rect 18854 7172 18910 7174
rect 19066 7226 19122 7228
rect 19066 7174 19068 7226
rect 19068 7174 19120 7226
rect 19120 7174 19122 7226
rect 19066 7172 19122 7174
rect 19277 7226 19333 7228
rect 19277 7174 19279 7226
rect 19279 7174 19331 7226
rect 19331 7174 19333 7226
rect 19277 7172 19333 7174
rect 19487 7226 19543 7228
rect 19487 7174 19489 7226
rect 19489 7174 19541 7226
rect 19541 7174 19543 7226
rect 19487 7172 19543 7174
rect 18191 6820 18247 6822
rect 18191 6768 18193 6820
rect 18193 6768 18245 6820
rect 18245 6768 18247 6820
rect 18191 6766 18247 6768
rect 18191 6602 18247 6604
rect 18191 6550 18193 6602
rect 18193 6550 18245 6602
rect 18245 6550 18247 6602
rect 18191 6548 18247 6550
rect 18191 6050 18247 6052
rect 18191 5998 18193 6050
rect 18193 5998 18245 6050
rect 18245 5998 18247 6050
rect 18191 5996 18247 5998
rect 18191 5832 18247 5834
rect 18191 5780 18193 5832
rect 18193 5780 18245 5832
rect 18245 5780 18247 5832
rect 18191 5778 18247 5780
rect 18433 5426 18489 5428
rect 18433 5374 18435 5426
rect 18435 5374 18487 5426
rect 18487 5374 18489 5426
rect 18433 5372 18489 5374
rect 18643 5426 18699 5428
rect 18643 5374 18645 5426
rect 18645 5374 18697 5426
rect 18697 5374 18699 5426
rect 18643 5372 18699 5374
rect 18854 5426 18910 5428
rect 18854 5374 18856 5426
rect 18856 5374 18908 5426
rect 18908 5374 18910 5426
rect 18854 5372 18910 5374
rect 19066 5426 19122 5428
rect 19066 5374 19068 5426
rect 19068 5374 19120 5426
rect 19120 5374 19122 5426
rect 19066 5372 19122 5374
rect 19277 5426 19333 5428
rect 19277 5374 19279 5426
rect 19279 5374 19331 5426
rect 19331 5374 19333 5426
rect 19277 5372 19333 5374
rect 19487 5426 19543 5428
rect 19487 5374 19489 5426
rect 19489 5374 19541 5426
rect 19541 5374 19543 5426
rect 19487 5372 19543 5374
rect 18191 5020 18247 5022
rect 18191 4968 18193 5020
rect 18193 4968 18245 5020
rect 18245 4968 18247 5020
rect 18191 4966 18247 4968
rect 18191 4802 18247 4804
rect 18191 4750 18193 4802
rect 18193 4750 18245 4802
rect 18245 4750 18247 4802
rect 18191 4748 18247 4750
rect 18191 4250 18247 4252
rect 18191 4198 18193 4250
rect 18193 4198 18245 4250
rect 18245 4198 18247 4250
rect 18191 4196 18247 4198
rect 18191 4032 18247 4034
rect 18191 3980 18193 4032
rect 18193 3980 18245 4032
rect 18245 3980 18247 4032
rect 18191 3978 18247 3980
rect 18433 3626 18489 3628
rect 18433 3574 18435 3626
rect 18435 3574 18487 3626
rect 18487 3574 18489 3626
rect 18433 3572 18489 3574
rect 18643 3626 18699 3628
rect 18643 3574 18645 3626
rect 18645 3574 18697 3626
rect 18697 3574 18699 3626
rect 18643 3572 18699 3574
rect 18854 3626 18910 3628
rect 18854 3574 18856 3626
rect 18856 3574 18908 3626
rect 18908 3574 18910 3626
rect 18854 3572 18910 3574
rect 19066 3626 19122 3628
rect 19066 3574 19068 3626
rect 19068 3574 19120 3626
rect 19120 3574 19122 3626
rect 19066 3572 19122 3574
rect 19277 3626 19333 3628
rect 19277 3574 19279 3626
rect 19279 3574 19331 3626
rect 19331 3574 19333 3626
rect 19277 3572 19333 3574
rect 19487 3626 19543 3628
rect 19487 3574 19489 3626
rect 19489 3574 19541 3626
rect 19541 3574 19543 3626
rect 19487 3572 19543 3574
rect 18191 3220 18247 3222
rect 18191 3168 18193 3220
rect 18193 3168 18245 3220
rect 18245 3168 18247 3220
rect 18191 3166 18247 3168
rect 18191 3002 18247 3004
rect 18191 2950 18193 3002
rect 18193 2950 18245 3002
rect 18245 2950 18247 3002
rect 18191 2948 18247 2950
rect 18191 2450 18247 2452
rect 18191 2398 18193 2450
rect 18193 2398 18245 2450
rect 18245 2398 18247 2450
rect 18191 2396 18247 2398
rect 18191 2232 18247 2234
rect 18191 2180 18193 2232
rect 18193 2180 18245 2232
rect 18245 2180 18247 2232
rect 18191 2178 18247 2180
rect 18433 1826 18489 1828
rect 18433 1774 18435 1826
rect 18435 1774 18487 1826
rect 18487 1774 18489 1826
rect 18433 1772 18489 1774
rect 18643 1826 18699 1828
rect 18643 1774 18645 1826
rect 18645 1774 18697 1826
rect 18697 1774 18699 1826
rect 18643 1772 18699 1774
rect 18854 1826 18910 1828
rect 18854 1774 18856 1826
rect 18856 1774 18908 1826
rect 18908 1774 18910 1826
rect 18854 1772 18910 1774
rect 19066 1826 19122 1828
rect 19066 1774 19068 1826
rect 19068 1774 19120 1826
rect 19120 1774 19122 1826
rect 19066 1772 19122 1774
rect 19277 1826 19333 1828
rect 19277 1774 19279 1826
rect 19279 1774 19331 1826
rect 19331 1774 19333 1826
rect 19277 1772 19333 1774
rect 19487 1826 19543 1828
rect 19487 1774 19489 1826
rect 19489 1774 19541 1826
rect 19541 1774 19543 1826
rect 19487 1772 19543 1774
rect 18191 1420 18247 1422
rect 18191 1368 18193 1420
rect 18193 1368 18245 1420
rect 18245 1368 18247 1420
rect 18191 1366 18247 1368
rect 18191 1202 18247 1204
rect 18191 1150 18193 1202
rect 18193 1150 18245 1202
rect 18245 1150 18247 1202
rect 18191 1148 18247 1150
rect 18191 650 18247 652
rect 18191 598 18193 650
rect 18193 598 18245 650
rect 18245 598 18247 650
rect 18191 596 18247 598
rect 18191 432 18247 434
rect 18191 380 18193 432
rect 18193 380 18245 432
rect 18245 380 18247 432
rect 18191 378 18247 380
rect 18433 26 18489 28
rect 18433 -26 18435 26
rect 18435 -26 18487 26
rect 18487 -26 18489 26
rect 18433 -28 18489 -26
rect 18643 26 18699 28
rect 18643 -26 18645 26
rect 18645 -26 18697 26
rect 18697 -26 18699 26
rect 18643 -28 18699 -26
rect 18854 26 18910 28
rect 18854 -26 18856 26
rect 18856 -26 18908 26
rect 18908 -26 18910 26
rect 18854 -28 18910 -26
rect 19066 26 19122 28
rect 19066 -26 19068 26
rect 19068 -26 19120 26
rect 19120 -26 19122 26
rect 19066 -28 19122 -26
rect 19277 26 19333 28
rect 19277 -26 19279 26
rect 19279 -26 19331 26
rect 19331 -26 19333 26
rect 19277 -28 19333 -26
rect 19487 26 19543 28
rect 19487 -26 19489 26
rect 19489 -26 19541 26
rect 19541 -26 19543 26
rect 19487 -28 19543 -26
rect 21911 14426 21967 14428
rect 21911 14374 21913 14426
rect 21913 14374 21965 14426
rect 21965 14374 21967 14426
rect 21911 14372 21967 14374
rect 22122 14426 22178 14428
rect 22122 14374 22124 14426
rect 22124 14374 22176 14426
rect 22176 14374 22178 14426
rect 22122 14372 22178 14374
rect 22333 14426 22389 14428
rect 22333 14374 22335 14426
rect 22335 14374 22387 14426
rect 22387 14374 22389 14426
rect 22333 14372 22389 14374
rect 22543 14426 22599 14428
rect 22543 14374 22545 14426
rect 22545 14374 22597 14426
rect 22597 14374 22599 14426
rect 22543 14372 22599 14374
rect 22754 14426 22810 14428
rect 22754 14374 22756 14426
rect 22756 14374 22808 14426
rect 22808 14374 22810 14426
rect 22754 14372 22810 14374
rect 22966 14426 23022 14428
rect 22966 14374 22968 14426
rect 22968 14374 23020 14426
rect 23020 14374 23022 14426
rect 22966 14372 23022 14374
rect 23177 14426 23233 14428
rect 23177 14374 23179 14426
rect 23179 14374 23231 14426
rect 23231 14374 23233 14426
rect 23177 14372 23233 14374
rect 23387 14426 23443 14428
rect 23387 14374 23389 14426
rect 23389 14374 23441 14426
rect 23441 14374 23443 14426
rect 23387 14372 23443 14374
rect 23598 14426 23654 14428
rect 23598 14374 23600 14426
rect 23600 14374 23652 14426
rect 23652 14374 23654 14426
rect 23598 14372 23654 14374
rect 23809 14426 23865 14428
rect 23809 14374 23811 14426
rect 23811 14374 23863 14426
rect 23863 14374 23865 14426
rect 23809 14372 23865 14374
rect 20668 13932 20724 13988
rect 20848 13932 20904 13988
rect 21430 13932 21486 13988
rect 21610 13932 21666 13988
rect 19758 13526 19814 13528
rect 19758 13474 19787 13526
rect 19787 13474 19814 13526
rect 19758 13472 19814 13474
rect 19969 13472 20025 13528
rect 20181 13472 20237 13528
rect 20392 13472 20448 13528
rect 20668 13012 20724 13068
rect 20848 13012 20904 13068
rect 21430 13012 21486 13068
rect 21610 13012 21666 13068
rect 21911 12626 21967 12628
rect 21911 12574 21913 12626
rect 21913 12574 21965 12626
rect 21965 12574 21967 12626
rect 21911 12572 21967 12574
rect 22122 12626 22178 12628
rect 22122 12574 22124 12626
rect 22124 12574 22176 12626
rect 22176 12574 22178 12626
rect 22122 12572 22178 12574
rect 22333 12626 22389 12628
rect 22333 12574 22335 12626
rect 22335 12574 22387 12626
rect 22387 12574 22389 12626
rect 22333 12572 22389 12574
rect 22543 12626 22599 12628
rect 22543 12574 22545 12626
rect 22545 12574 22597 12626
rect 22597 12574 22599 12626
rect 22543 12572 22599 12574
rect 22754 12626 22810 12628
rect 22754 12574 22756 12626
rect 22756 12574 22808 12626
rect 22808 12574 22810 12626
rect 22754 12572 22810 12574
rect 22966 12626 23022 12628
rect 22966 12574 22968 12626
rect 22968 12574 23020 12626
rect 23020 12574 23022 12626
rect 22966 12572 23022 12574
rect 23177 12626 23233 12628
rect 23177 12574 23179 12626
rect 23179 12574 23231 12626
rect 23231 12574 23233 12626
rect 23177 12572 23233 12574
rect 23387 12626 23443 12628
rect 23387 12574 23389 12626
rect 23389 12574 23441 12626
rect 23441 12574 23443 12626
rect 23387 12572 23443 12574
rect 23598 12626 23654 12628
rect 23598 12574 23600 12626
rect 23600 12574 23652 12626
rect 23652 12574 23654 12626
rect 23598 12572 23654 12574
rect 23809 12626 23865 12628
rect 23809 12574 23811 12626
rect 23811 12574 23863 12626
rect 23863 12574 23865 12626
rect 23809 12572 23865 12574
rect 20668 12132 20724 12188
rect 20848 12132 20904 12188
rect 21430 12132 21486 12188
rect 21610 12132 21666 12188
rect 19758 11726 19814 11728
rect 19758 11674 19787 11726
rect 19787 11674 19814 11726
rect 19758 11672 19814 11674
rect 19969 11672 20025 11728
rect 20181 11672 20237 11728
rect 20392 11672 20448 11728
rect 20668 11212 20724 11268
rect 20848 11212 20904 11268
rect 21430 11212 21486 11268
rect 21610 11212 21666 11268
rect 21911 10826 21967 10828
rect 21911 10774 21913 10826
rect 21913 10774 21965 10826
rect 21965 10774 21967 10826
rect 21911 10772 21967 10774
rect 22122 10826 22178 10828
rect 22122 10774 22124 10826
rect 22124 10774 22176 10826
rect 22176 10774 22178 10826
rect 22122 10772 22178 10774
rect 22333 10826 22389 10828
rect 22333 10774 22335 10826
rect 22335 10774 22387 10826
rect 22387 10774 22389 10826
rect 22333 10772 22389 10774
rect 22543 10826 22599 10828
rect 22543 10774 22545 10826
rect 22545 10774 22597 10826
rect 22597 10774 22599 10826
rect 22543 10772 22599 10774
rect 22754 10826 22810 10828
rect 22754 10774 22756 10826
rect 22756 10774 22808 10826
rect 22808 10774 22810 10826
rect 22754 10772 22810 10774
rect 22966 10826 23022 10828
rect 22966 10774 22968 10826
rect 22968 10774 23020 10826
rect 23020 10774 23022 10826
rect 22966 10772 23022 10774
rect 23177 10826 23233 10828
rect 23177 10774 23179 10826
rect 23179 10774 23231 10826
rect 23231 10774 23233 10826
rect 23177 10772 23233 10774
rect 23387 10826 23443 10828
rect 23387 10774 23389 10826
rect 23389 10774 23441 10826
rect 23441 10774 23443 10826
rect 23387 10772 23443 10774
rect 23598 10826 23654 10828
rect 23598 10774 23600 10826
rect 23600 10774 23652 10826
rect 23652 10774 23654 10826
rect 23598 10772 23654 10774
rect 23809 10826 23865 10828
rect 23809 10774 23811 10826
rect 23811 10774 23863 10826
rect 23863 10774 23865 10826
rect 23809 10772 23865 10774
rect 20668 10332 20724 10388
rect 20848 10332 20904 10388
rect 21430 10332 21486 10388
rect 21610 10332 21666 10388
rect 19758 9926 19814 9928
rect 19758 9874 19787 9926
rect 19787 9874 19814 9926
rect 19758 9872 19814 9874
rect 19969 9872 20025 9928
rect 20181 9872 20237 9928
rect 20392 9872 20448 9928
rect 20668 9412 20724 9468
rect 20848 9412 20904 9468
rect 21430 9412 21486 9468
rect 21610 9412 21666 9468
rect 21911 9026 21967 9028
rect 21911 8974 21913 9026
rect 21913 8974 21965 9026
rect 21965 8974 21967 9026
rect 21911 8972 21967 8974
rect 22122 9026 22178 9028
rect 22122 8974 22124 9026
rect 22124 8974 22176 9026
rect 22176 8974 22178 9026
rect 22122 8972 22178 8974
rect 22333 9026 22389 9028
rect 22333 8974 22335 9026
rect 22335 8974 22387 9026
rect 22387 8974 22389 9026
rect 22333 8972 22389 8974
rect 22543 9026 22599 9028
rect 22543 8974 22545 9026
rect 22545 8974 22597 9026
rect 22597 8974 22599 9026
rect 22543 8972 22599 8974
rect 22754 9026 22810 9028
rect 22754 8974 22756 9026
rect 22756 8974 22808 9026
rect 22808 8974 22810 9026
rect 22754 8972 22810 8974
rect 22966 9026 23022 9028
rect 22966 8974 22968 9026
rect 22968 8974 23020 9026
rect 23020 8974 23022 9026
rect 22966 8972 23022 8974
rect 23177 9026 23233 9028
rect 23177 8974 23179 9026
rect 23179 8974 23231 9026
rect 23231 8974 23233 9026
rect 23177 8972 23233 8974
rect 23387 9026 23443 9028
rect 23387 8974 23389 9026
rect 23389 8974 23441 9026
rect 23441 8974 23443 9026
rect 23387 8972 23443 8974
rect 23598 9026 23654 9028
rect 23598 8974 23600 9026
rect 23600 8974 23652 9026
rect 23652 8974 23654 9026
rect 23598 8972 23654 8974
rect 23809 9026 23865 9028
rect 23809 8974 23811 9026
rect 23811 8974 23863 9026
rect 23863 8974 23865 9026
rect 23809 8972 23865 8974
rect 20668 8532 20724 8588
rect 20848 8532 20904 8588
rect 21430 8532 21486 8588
rect 21610 8532 21666 8588
rect 19758 8126 19814 8128
rect 19758 8074 19787 8126
rect 19787 8074 19814 8126
rect 19758 8072 19814 8074
rect 19969 8072 20025 8128
rect 20181 8072 20237 8128
rect 20392 8072 20448 8128
rect 20668 7612 20724 7668
rect 20848 7612 20904 7668
rect 21430 7612 21486 7668
rect 21610 7612 21666 7668
rect 21911 7226 21967 7228
rect 21911 7174 21913 7226
rect 21913 7174 21965 7226
rect 21965 7174 21967 7226
rect 21911 7172 21967 7174
rect 22122 7226 22178 7228
rect 22122 7174 22124 7226
rect 22124 7174 22176 7226
rect 22176 7174 22178 7226
rect 22122 7172 22178 7174
rect 22333 7226 22389 7228
rect 22333 7174 22335 7226
rect 22335 7174 22387 7226
rect 22387 7174 22389 7226
rect 22333 7172 22389 7174
rect 22543 7226 22599 7228
rect 22543 7174 22545 7226
rect 22545 7174 22597 7226
rect 22597 7174 22599 7226
rect 22543 7172 22599 7174
rect 22754 7226 22810 7228
rect 22754 7174 22756 7226
rect 22756 7174 22808 7226
rect 22808 7174 22810 7226
rect 22754 7172 22810 7174
rect 22966 7226 23022 7228
rect 22966 7174 22968 7226
rect 22968 7174 23020 7226
rect 23020 7174 23022 7226
rect 22966 7172 23022 7174
rect 23177 7226 23233 7228
rect 23177 7174 23179 7226
rect 23179 7174 23231 7226
rect 23231 7174 23233 7226
rect 23177 7172 23233 7174
rect 23387 7226 23443 7228
rect 23387 7174 23389 7226
rect 23389 7174 23441 7226
rect 23441 7174 23443 7226
rect 23387 7172 23443 7174
rect 23598 7226 23654 7228
rect 23598 7174 23600 7226
rect 23600 7174 23652 7226
rect 23652 7174 23654 7226
rect 23598 7172 23654 7174
rect 23809 7226 23865 7228
rect 23809 7174 23811 7226
rect 23811 7174 23863 7226
rect 23863 7174 23865 7226
rect 23809 7172 23865 7174
rect 20668 6732 20724 6788
rect 20848 6732 20904 6788
rect 21430 6732 21486 6788
rect 21610 6732 21666 6788
rect 19758 6326 19814 6328
rect 19758 6274 19787 6326
rect 19787 6274 19814 6326
rect 19758 6272 19814 6274
rect 19969 6272 20025 6328
rect 20181 6272 20237 6328
rect 20392 6272 20448 6328
rect 20668 5812 20724 5868
rect 20848 5812 20904 5868
rect 21430 5812 21486 5868
rect 21610 5812 21666 5868
rect 21911 5426 21967 5428
rect 21911 5374 21913 5426
rect 21913 5374 21965 5426
rect 21965 5374 21967 5426
rect 21911 5372 21967 5374
rect 22122 5426 22178 5428
rect 22122 5374 22124 5426
rect 22124 5374 22176 5426
rect 22176 5374 22178 5426
rect 22122 5372 22178 5374
rect 22333 5426 22389 5428
rect 22333 5374 22335 5426
rect 22335 5374 22387 5426
rect 22387 5374 22389 5426
rect 22333 5372 22389 5374
rect 22543 5426 22599 5428
rect 22543 5374 22545 5426
rect 22545 5374 22597 5426
rect 22597 5374 22599 5426
rect 22543 5372 22599 5374
rect 22754 5426 22810 5428
rect 22754 5374 22756 5426
rect 22756 5374 22808 5426
rect 22808 5374 22810 5426
rect 22754 5372 22810 5374
rect 22966 5426 23022 5428
rect 22966 5374 22968 5426
rect 22968 5374 23020 5426
rect 23020 5374 23022 5426
rect 22966 5372 23022 5374
rect 23177 5426 23233 5428
rect 23177 5374 23179 5426
rect 23179 5374 23231 5426
rect 23231 5374 23233 5426
rect 23177 5372 23233 5374
rect 23387 5426 23443 5428
rect 23387 5374 23389 5426
rect 23389 5374 23441 5426
rect 23441 5374 23443 5426
rect 23387 5372 23443 5374
rect 23598 5426 23654 5428
rect 23598 5374 23600 5426
rect 23600 5374 23652 5426
rect 23652 5374 23654 5426
rect 23598 5372 23654 5374
rect 23809 5426 23865 5428
rect 23809 5374 23811 5426
rect 23811 5374 23863 5426
rect 23863 5374 23865 5426
rect 23809 5372 23865 5374
rect 20668 4932 20724 4988
rect 20848 4932 20904 4988
rect 21430 4932 21486 4988
rect 21610 4932 21666 4988
rect 19758 4526 19814 4528
rect 19758 4474 19787 4526
rect 19787 4474 19814 4526
rect 19758 4472 19814 4474
rect 19969 4472 20025 4528
rect 20181 4472 20237 4528
rect 20392 4472 20448 4528
rect 20668 4012 20724 4068
rect 20848 4012 20904 4068
rect 21430 4012 21486 4068
rect 21610 4012 21666 4068
rect 21911 3626 21967 3628
rect 21911 3574 21913 3626
rect 21913 3574 21965 3626
rect 21965 3574 21967 3626
rect 21911 3572 21967 3574
rect 22122 3626 22178 3628
rect 22122 3574 22124 3626
rect 22124 3574 22176 3626
rect 22176 3574 22178 3626
rect 22122 3572 22178 3574
rect 22333 3626 22389 3628
rect 22333 3574 22335 3626
rect 22335 3574 22387 3626
rect 22387 3574 22389 3626
rect 22333 3572 22389 3574
rect 22543 3626 22599 3628
rect 22543 3574 22545 3626
rect 22545 3574 22597 3626
rect 22597 3574 22599 3626
rect 22543 3572 22599 3574
rect 22754 3626 22810 3628
rect 22754 3574 22756 3626
rect 22756 3574 22808 3626
rect 22808 3574 22810 3626
rect 22754 3572 22810 3574
rect 22966 3626 23022 3628
rect 22966 3574 22968 3626
rect 22968 3574 23020 3626
rect 23020 3574 23022 3626
rect 22966 3572 23022 3574
rect 23177 3626 23233 3628
rect 23177 3574 23179 3626
rect 23179 3574 23231 3626
rect 23231 3574 23233 3626
rect 23177 3572 23233 3574
rect 23387 3626 23443 3628
rect 23387 3574 23389 3626
rect 23389 3574 23441 3626
rect 23441 3574 23443 3626
rect 23387 3572 23443 3574
rect 23598 3626 23654 3628
rect 23598 3574 23600 3626
rect 23600 3574 23652 3626
rect 23652 3574 23654 3626
rect 23598 3572 23654 3574
rect 23809 3626 23865 3628
rect 23809 3574 23811 3626
rect 23811 3574 23863 3626
rect 23863 3574 23865 3626
rect 23809 3572 23865 3574
rect 20668 3132 20724 3188
rect 20848 3132 20904 3188
rect 21430 3132 21486 3188
rect 21610 3132 21666 3188
rect 19758 2726 19814 2728
rect 19758 2674 19787 2726
rect 19787 2674 19814 2726
rect 19758 2672 19814 2674
rect 19969 2672 20025 2728
rect 20181 2672 20237 2728
rect 20392 2672 20448 2728
rect 20668 2212 20724 2268
rect 20848 2212 20904 2268
rect 21430 2212 21486 2268
rect 21610 2212 21666 2268
rect 21911 1826 21967 1828
rect 21911 1774 21913 1826
rect 21913 1774 21965 1826
rect 21965 1774 21967 1826
rect 21911 1772 21967 1774
rect 22122 1826 22178 1828
rect 22122 1774 22124 1826
rect 22124 1774 22176 1826
rect 22176 1774 22178 1826
rect 22122 1772 22178 1774
rect 22333 1826 22389 1828
rect 22333 1774 22335 1826
rect 22335 1774 22387 1826
rect 22387 1774 22389 1826
rect 22333 1772 22389 1774
rect 22543 1826 22599 1828
rect 22543 1774 22545 1826
rect 22545 1774 22597 1826
rect 22597 1774 22599 1826
rect 22543 1772 22599 1774
rect 22754 1826 22810 1828
rect 22754 1774 22756 1826
rect 22756 1774 22808 1826
rect 22808 1774 22810 1826
rect 22754 1772 22810 1774
rect 22966 1826 23022 1828
rect 22966 1774 22968 1826
rect 22968 1774 23020 1826
rect 23020 1774 23022 1826
rect 22966 1772 23022 1774
rect 23177 1826 23233 1828
rect 23177 1774 23179 1826
rect 23179 1774 23231 1826
rect 23231 1774 23233 1826
rect 23177 1772 23233 1774
rect 23387 1826 23443 1828
rect 23387 1774 23389 1826
rect 23389 1774 23441 1826
rect 23441 1774 23443 1826
rect 23387 1772 23443 1774
rect 23598 1826 23654 1828
rect 23598 1774 23600 1826
rect 23600 1774 23652 1826
rect 23652 1774 23654 1826
rect 23598 1772 23654 1774
rect 23809 1826 23865 1828
rect 23809 1774 23811 1826
rect 23811 1774 23863 1826
rect 23863 1774 23865 1826
rect 23809 1772 23865 1774
rect 20668 1332 20724 1388
rect 20848 1332 20904 1388
rect 21430 1332 21486 1388
rect 21610 1332 21666 1388
rect 19758 926 19814 928
rect 19758 874 19787 926
rect 19787 874 19814 926
rect 19758 872 19814 874
rect 19969 872 20025 928
rect 20181 872 20237 928
rect 20392 872 20448 928
rect 20668 412 20724 468
rect 20848 412 20904 468
rect 21430 412 21486 468
rect 21610 412 21666 468
rect 21911 26 21967 28
rect 21911 -26 21913 26
rect 21913 -26 21965 26
rect 21965 -26 21967 26
rect 21911 -28 21967 -26
rect 22122 26 22178 28
rect 22122 -26 22124 26
rect 22124 -26 22176 26
rect 22176 -26 22178 26
rect 22122 -28 22178 -26
rect 22333 26 22389 28
rect 22333 -26 22335 26
rect 22335 -26 22387 26
rect 22387 -26 22389 26
rect 22333 -28 22389 -26
rect 22543 26 22599 28
rect 22543 -26 22545 26
rect 22545 -26 22597 26
rect 22597 -26 22599 26
rect 22543 -28 22599 -26
rect 22754 26 22810 28
rect 22754 -26 22756 26
rect 22756 -26 22808 26
rect 22808 -26 22810 26
rect 22754 -28 22810 -26
rect 22966 26 23022 28
rect 22966 -26 22968 26
rect 22968 -26 23020 26
rect 23020 -26 23022 26
rect 22966 -28 23022 -26
rect 23177 26 23233 28
rect 23177 -26 23179 26
rect 23179 -26 23231 26
rect 23231 -26 23233 26
rect 23177 -28 23233 -26
rect 23387 26 23443 28
rect 23387 -26 23389 26
rect 23389 -26 23441 26
rect 23441 -26 23443 26
rect 23387 -28 23443 -26
rect 23598 26 23654 28
rect 23598 -26 23600 26
rect 23600 -26 23652 26
rect 23652 -26 23654 26
rect 23598 -28 23654 -26
rect 23809 26 23865 28
rect 23809 -26 23811 26
rect 23811 -26 23863 26
rect 23863 -26 23865 26
rect 23809 -28 23865 -26
<< metal3 >>
rect 0 14428 24219 14500
rect 0 14372 449 14428
rect 505 14372 660 14428
rect 716 14372 871 14428
rect 927 14372 1081 14428
rect 1137 14372 1292 14428
rect 1348 14372 1504 14428
rect 1560 14372 1715 14428
rect 1771 14372 1925 14428
rect 1981 14372 2136 14428
rect 2192 14372 2347 14428
rect 2403 14372 4815 14428
rect 4871 14372 5025 14428
rect 5081 14372 5236 14428
rect 5292 14372 5448 14428
rect 5504 14372 5659 14428
rect 5715 14372 5869 14428
rect 5925 14372 8647 14428
rect 8703 14372 8827 14428
rect 8883 14372 14429 14428
rect 14485 14372 14640 14428
rect 14696 14372 14851 14428
rect 14907 14372 18433 14428
rect 18489 14372 18643 14428
rect 18699 14372 18854 14428
rect 18910 14372 19066 14428
rect 19122 14372 19277 14428
rect 19333 14372 19487 14428
rect 19543 14372 21911 14428
rect 21967 14372 22122 14428
rect 22178 14372 22333 14428
rect 22389 14372 22543 14428
rect 22599 14372 22754 14428
rect 22810 14372 22966 14428
rect 23022 14372 23177 14428
rect 23233 14372 23387 14428
rect 23443 14372 23598 14428
rect 23654 14372 23809 14428
rect 23865 14372 24219 14428
rect 0 14300 24219 14372
rect 6245 14074 9638 14075
rect 0 13995 3687 14061
rect 0 13939 2652 13995
rect 2708 13939 2832 13995
rect 2888 13988 3687 13995
rect 2888 13939 3414 13988
rect 0 13932 3414 13939
rect 3470 13932 3594 13988
rect 3650 13932 3687 13988
rect 6237 14036 9682 14074
rect 6237 13980 6273 14036
rect 6329 13980 9589 14036
rect 9645 13980 9682 14036
rect 6237 13941 9682 13980
rect 18154 14022 18284 14061
rect 18154 13966 18191 14022
rect 18247 13966 18284 14022
rect 0 13859 3687 13932
rect 18154 13843 18284 13966
rect 20631 13988 24219 14061
rect 20631 13932 20668 13988
rect 20724 13932 20848 13988
rect 20904 13932 21430 13988
rect 21486 13932 21610 13988
rect 21666 13932 24219 13988
rect 20631 13859 24219 13932
rect 7449 13805 18284 13843
rect 7449 13749 7486 13805
rect 7542 13749 7666 13805
rect 7722 13749 9370 13805
rect 9426 13804 18284 13805
rect 9426 13749 18191 13804
rect 7449 13748 18191 13749
rect 18247 13748 18284 13804
rect 7449 13710 18284 13748
rect 0 13528 24219 13601
rect 0 13472 3879 13528
rect 3935 13472 4090 13528
rect 4146 13472 4302 13528
rect 4358 13472 4513 13528
rect 4569 13472 7925 13528
rect 7981 13472 8136 13528
rect 8192 13472 8347 13528
rect 8403 13472 9848 13528
rect 9904 13472 10028 13528
rect 10084 13472 13385 13528
rect 13441 13472 13596 13528
rect 13652 13472 13808 13528
rect 13864 13472 14019 13528
rect 14075 13472 19758 13528
rect 19814 13472 19969 13528
rect 20025 13472 20181 13528
rect 20237 13472 20392 13528
rect 20448 13472 24219 13528
rect 0 13399 24219 13472
rect 7449 13252 18284 13290
rect 7449 13251 18191 13252
rect 7449 13195 7486 13251
rect 7542 13195 7666 13251
rect 7722 13195 9370 13251
rect 9426 13196 18191 13251
rect 18247 13196 18284 13252
rect 9426 13195 18284 13196
rect 7449 13157 18284 13195
rect 0 13068 3687 13141
rect 0 13061 3414 13068
rect 0 13005 2652 13061
rect 2708 13005 2832 13061
rect 2888 13012 3414 13061
rect 3470 13012 3594 13068
rect 3650 13012 3687 13068
rect 2888 13005 3687 13012
rect 0 12939 3687 13005
rect 6237 13020 9682 13059
rect 6237 12964 6273 13020
rect 6329 12964 9589 13020
rect 9645 12964 9682 13020
rect 6237 12926 9682 12964
rect 18154 13034 18284 13157
rect 18154 12978 18191 13034
rect 18247 12978 18284 13034
rect 18154 12939 18284 12978
rect 20631 13068 24219 13141
rect 20631 13012 20668 13068
rect 20724 13012 20848 13068
rect 20904 13012 21430 13068
rect 21486 13012 21610 13068
rect 21666 13012 24219 13068
rect 20631 12939 24219 13012
rect 6245 12925 9638 12926
rect 0 12628 24219 12700
rect 0 12572 449 12628
rect 505 12572 660 12628
rect 716 12572 871 12628
rect 927 12572 1081 12628
rect 1137 12572 1292 12628
rect 1348 12572 1504 12628
rect 1560 12572 1715 12628
rect 1771 12572 1925 12628
rect 1981 12572 2136 12628
rect 2192 12572 2347 12628
rect 2403 12572 4815 12628
rect 4871 12572 5025 12628
rect 5081 12572 5236 12628
rect 5292 12572 5448 12628
rect 5504 12572 5659 12628
rect 5715 12572 5869 12628
rect 5925 12572 8647 12628
rect 8703 12572 8827 12628
rect 8883 12572 14429 12628
rect 14485 12572 14640 12628
rect 14696 12572 14851 12628
rect 14907 12572 18433 12628
rect 18489 12572 18643 12628
rect 18699 12572 18854 12628
rect 18910 12572 19066 12628
rect 19122 12572 19277 12628
rect 19333 12572 19487 12628
rect 19543 12572 21911 12628
rect 21967 12572 22122 12628
rect 22178 12572 22333 12628
rect 22389 12572 22543 12628
rect 22599 12572 22754 12628
rect 22810 12572 22966 12628
rect 23022 12572 23177 12628
rect 23233 12572 23387 12628
rect 23443 12572 23598 12628
rect 23654 12572 23809 12628
rect 23865 12572 24219 12628
rect 0 12500 24219 12572
rect 6245 12274 9638 12275
rect 0 12195 3687 12261
rect 0 12139 2652 12195
rect 2708 12139 2832 12195
rect 2888 12188 3687 12195
rect 2888 12139 3414 12188
rect 0 12132 3414 12139
rect 3470 12132 3594 12188
rect 3650 12132 3687 12188
rect 6237 12236 9682 12274
rect 6237 12180 6273 12236
rect 6329 12180 9589 12236
rect 9645 12180 9682 12236
rect 6237 12141 9682 12180
rect 18154 12222 18284 12261
rect 18154 12166 18191 12222
rect 18247 12166 18284 12222
rect 0 12059 3687 12132
rect 18154 12043 18284 12166
rect 20631 12188 24219 12261
rect 20631 12132 20668 12188
rect 20724 12132 20848 12188
rect 20904 12132 21430 12188
rect 21486 12132 21610 12188
rect 21666 12132 24219 12188
rect 20631 12059 24219 12132
rect 7449 12005 18284 12043
rect 7449 11949 7486 12005
rect 7542 11949 7666 12005
rect 7722 11949 9370 12005
rect 9426 12004 18284 12005
rect 9426 11949 18191 12004
rect 7449 11948 18191 11949
rect 18247 11948 18284 12004
rect 7449 11910 18284 11948
rect 0 11728 24219 11801
rect 0 11672 3879 11728
rect 3935 11672 4090 11728
rect 4146 11672 4302 11728
rect 4358 11672 4513 11728
rect 4569 11672 7925 11728
rect 7981 11672 8136 11728
rect 8192 11672 8347 11728
rect 8403 11672 9848 11728
rect 9904 11672 10028 11728
rect 10084 11672 13385 11728
rect 13441 11672 13596 11728
rect 13652 11672 13808 11728
rect 13864 11672 14019 11728
rect 14075 11672 19758 11728
rect 19814 11672 19969 11728
rect 20025 11672 20181 11728
rect 20237 11672 20392 11728
rect 20448 11672 24219 11728
rect 0 11599 24219 11672
rect 7449 11452 18284 11490
rect 7449 11451 18191 11452
rect 7449 11395 7486 11451
rect 7542 11395 7666 11451
rect 7722 11395 9370 11451
rect 9426 11396 18191 11451
rect 18247 11396 18284 11452
rect 9426 11395 18284 11396
rect 7449 11357 18284 11395
rect 0 11268 3687 11341
rect 0 11261 3414 11268
rect 0 11205 2652 11261
rect 2708 11205 2832 11261
rect 2888 11212 3414 11261
rect 3470 11212 3594 11268
rect 3650 11212 3687 11268
rect 2888 11205 3687 11212
rect 0 11139 3687 11205
rect 6237 11220 9682 11259
rect 6237 11164 6273 11220
rect 6329 11164 9589 11220
rect 9645 11164 9682 11220
rect 6237 11126 9682 11164
rect 18154 11234 18284 11357
rect 18154 11178 18191 11234
rect 18247 11178 18284 11234
rect 18154 11139 18284 11178
rect 20631 11268 24219 11341
rect 20631 11212 20668 11268
rect 20724 11212 20848 11268
rect 20904 11212 21430 11268
rect 21486 11212 21610 11268
rect 21666 11212 24219 11268
rect 20631 11139 24219 11212
rect 6245 11125 9638 11126
rect 0 10828 24219 10900
rect 0 10772 449 10828
rect 505 10772 660 10828
rect 716 10772 871 10828
rect 927 10772 1081 10828
rect 1137 10772 1292 10828
rect 1348 10772 1504 10828
rect 1560 10772 1715 10828
rect 1771 10772 1925 10828
rect 1981 10772 2136 10828
rect 2192 10772 2347 10828
rect 2403 10772 4815 10828
rect 4871 10772 5025 10828
rect 5081 10772 5236 10828
rect 5292 10772 5448 10828
rect 5504 10772 5659 10828
rect 5715 10772 5869 10828
rect 5925 10772 8647 10828
rect 8703 10772 8827 10828
rect 8883 10772 14429 10828
rect 14485 10772 14640 10828
rect 14696 10772 14851 10828
rect 14907 10772 18433 10828
rect 18489 10772 18643 10828
rect 18699 10772 18854 10828
rect 18910 10772 19066 10828
rect 19122 10772 19277 10828
rect 19333 10772 19487 10828
rect 19543 10772 21911 10828
rect 21967 10772 22122 10828
rect 22178 10772 22333 10828
rect 22389 10772 22543 10828
rect 22599 10772 22754 10828
rect 22810 10772 22966 10828
rect 23022 10772 23177 10828
rect 23233 10772 23387 10828
rect 23443 10772 23598 10828
rect 23654 10772 23809 10828
rect 23865 10772 24219 10828
rect 0 10700 24219 10772
rect 6245 10474 9638 10475
rect 0 10395 3687 10461
rect 0 10339 2652 10395
rect 2708 10339 2832 10395
rect 2888 10388 3687 10395
rect 2888 10339 3414 10388
rect 0 10332 3414 10339
rect 3470 10332 3594 10388
rect 3650 10332 3687 10388
rect 6237 10436 9682 10474
rect 6237 10380 6273 10436
rect 6329 10380 9589 10436
rect 9645 10380 9682 10436
rect 6237 10341 9682 10380
rect 18154 10422 18284 10461
rect 18154 10366 18191 10422
rect 18247 10366 18284 10422
rect 0 10259 3687 10332
rect 18154 10243 18284 10366
rect 20631 10388 24219 10461
rect 20631 10332 20668 10388
rect 20724 10332 20848 10388
rect 20904 10332 21430 10388
rect 21486 10332 21610 10388
rect 21666 10332 24219 10388
rect 20631 10259 24219 10332
rect 7449 10205 18284 10243
rect 7449 10149 7486 10205
rect 7542 10149 7666 10205
rect 7722 10149 9370 10205
rect 9426 10204 18284 10205
rect 9426 10149 18191 10204
rect 7449 10148 18191 10149
rect 18247 10148 18284 10204
rect 7449 10110 18284 10148
rect 0 9928 24219 10001
rect 0 9872 3879 9928
rect 3935 9872 4090 9928
rect 4146 9872 4302 9928
rect 4358 9872 4513 9928
rect 4569 9872 7925 9928
rect 7981 9872 8136 9928
rect 8192 9872 8347 9928
rect 8403 9872 9848 9928
rect 9904 9872 10028 9928
rect 10084 9872 13385 9928
rect 13441 9872 13596 9928
rect 13652 9872 13808 9928
rect 13864 9872 14019 9928
rect 14075 9872 19758 9928
rect 19814 9872 19969 9928
rect 20025 9872 20181 9928
rect 20237 9872 20392 9928
rect 20448 9872 24219 9928
rect 0 9799 24219 9872
rect 7449 9652 18284 9690
rect 7449 9651 18191 9652
rect 7449 9595 7486 9651
rect 7542 9595 7666 9651
rect 7722 9595 9370 9651
rect 9426 9596 18191 9651
rect 18247 9596 18284 9652
rect 9426 9595 18284 9596
rect 7449 9557 18284 9595
rect 0 9468 3687 9541
rect 0 9461 3414 9468
rect 0 9405 2652 9461
rect 2708 9405 2832 9461
rect 2888 9412 3414 9461
rect 3470 9412 3594 9468
rect 3650 9412 3687 9468
rect 2888 9405 3687 9412
rect 0 9339 3687 9405
rect 6237 9420 9682 9459
rect 6237 9364 6273 9420
rect 6329 9364 9589 9420
rect 9645 9364 9682 9420
rect 6237 9326 9682 9364
rect 18154 9434 18284 9557
rect 18154 9378 18191 9434
rect 18247 9378 18284 9434
rect 18154 9339 18284 9378
rect 20631 9468 24219 9541
rect 20631 9412 20668 9468
rect 20724 9412 20848 9468
rect 20904 9412 21430 9468
rect 21486 9412 21610 9468
rect 21666 9412 24219 9468
rect 20631 9339 24219 9412
rect 6245 9325 9638 9326
rect 0 9028 24219 9100
rect 0 8972 449 9028
rect 505 8972 660 9028
rect 716 8972 871 9028
rect 927 8972 1081 9028
rect 1137 8972 1292 9028
rect 1348 8972 1504 9028
rect 1560 8972 1715 9028
rect 1771 8972 1925 9028
rect 1981 8972 2136 9028
rect 2192 8972 2347 9028
rect 2403 8972 4815 9028
rect 4871 8972 5025 9028
rect 5081 8972 5236 9028
rect 5292 8972 5448 9028
rect 5504 8972 5659 9028
rect 5715 8972 5869 9028
rect 5925 8972 8647 9028
rect 8703 8972 8827 9028
rect 8883 8972 14429 9028
rect 14485 8972 14640 9028
rect 14696 8972 14851 9028
rect 14907 8972 18433 9028
rect 18489 8972 18643 9028
rect 18699 8972 18854 9028
rect 18910 8972 19066 9028
rect 19122 8972 19277 9028
rect 19333 8972 19487 9028
rect 19543 8972 21911 9028
rect 21967 8972 22122 9028
rect 22178 8972 22333 9028
rect 22389 8972 22543 9028
rect 22599 8972 22754 9028
rect 22810 8972 22966 9028
rect 23022 8972 23177 9028
rect 23233 8972 23387 9028
rect 23443 8972 23598 9028
rect 23654 8972 23809 9028
rect 23865 8972 24219 9028
rect 0 8900 24219 8972
rect 6245 8674 9638 8675
rect 0 8595 3687 8661
rect 0 8539 2652 8595
rect 2708 8539 2832 8595
rect 2888 8588 3687 8595
rect 2888 8539 3414 8588
rect 0 8532 3414 8539
rect 3470 8532 3594 8588
rect 3650 8532 3687 8588
rect 6237 8636 9682 8674
rect 6237 8580 6273 8636
rect 6329 8580 9589 8636
rect 9645 8580 9682 8636
rect 6237 8541 9682 8580
rect 18154 8622 18284 8661
rect 18154 8566 18191 8622
rect 18247 8566 18284 8622
rect 0 8459 3687 8532
rect 18154 8443 18284 8566
rect 20631 8588 24219 8661
rect 20631 8532 20668 8588
rect 20724 8532 20848 8588
rect 20904 8532 21430 8588
rect 21486 8532 21610 8588
rect 21666 8532 24219 8588
rect 20631 8459 24219 8532
rect 7449 8405 18284 8443
rect 7449 8349 7486 8405
rect 7542 8349 7666 8405
rect 7722 8349 9370 8405
rect 9426 8404 18284 8405
rect 9426 8349 18191 8404
rect 7449 8348 18191 8349
rect 18247 8348 18284 8404
rect 7449 8310 18284 8348
rect 0 8128 24219 8201
rect 0 8072 3879 8128
rect 3935 8072 4090 8128
rect 4146 8072 4302 8128
rect 4358 8072 4513 8128
rect 4569 8072 7925 8128
rect 7981 8072 8136 8128
rect 8192 8072 8347 8128
rect 8403 8072 9848 8128
rect 9904 8072 10028 8128
rect 10084 8072 13385 8128
rect 13441 8072 13596 8128
rect 13652 8072 13808 8128
rect 13864 8072 14019 8128
rect 14075 8072 19758 8128
rect 19814 8072 19969 8128
rect 20025 8072 20181 8128
rect 20237 8072 20392 8128
rect 20448 8072 24219 8128
rect 0 7999 24219 8072
rect 7449 7852 18284 7890
rect 7449 7851 18191 7852
rect 7449 7795 7486 7851
rect 7542 7795 7666 7851
rect 7722 7795 9370 7851
rect 9426 7796 18191 7851
rect 18247 7796 18284 7852
rect 9426 7795 18284 7796
rect 7449 7757 18284 7795
rect 0 7668 3687 7741
rect 0 7661 3414 7668
rect 0 7605 2652 7661
rect 2708 7605 2832 7661
rect 2888 7612 3414 7661
rect 3470 7612 3594 7668
rect 3650 7612 3687 7668
rect 2888 7605 3687 7612
rect 0 7539 3687 7605
rect 6237 7620 9682 7659
rect 6237 7564 6273 7620
rect 6329 7564 9589 7620
rect 9645 7564 9682 7620
rect 6237 7526 9682 7564
rect 18154 7634 18284 7757
rect 18154 7578 18191 7634
rect 18247 7578 18284 7634
rect 18154 7539 18284 7578
rect 20631 7668 24219 7741
rect 20631 7612 20668 7668
rect 20724 7612 20848 7668
rect 20904 7612 21430 7668
rect 21486 7612 21610 7668
rect 21666 7612 24219 7668
rect 20631 7539 24219 7612
rect 6245 7525 9638 7526
rect 0 7228 24219 7300
rect 0 7172 449 7228
rect 505 7172 660 7228
rect 716 7172 871 7228
rect 927 7172 1081 7228
rect 1137 7172 1292 7228
rect 1348 7172 1504 7228
rect 1560 7172 1715 7228
rect 1771 7172 1925 7228
rect 1981 7172 2136 7228
rect 2192 7172 2347 7228
rect 2403 7172 4815 7228
rect 4871 7172 5025 7228
rect 5081 7172 5236 7228
rect 5292 7172 5448 7228
rect 5504 7172 5659 7228
rect 5715 7172 5869 7228
rect 5925 7172 8647 7228
rect 8703 7172 8827 7228
rect 8883 7172 14429 7228
rect 14485 7172 14640 7228
rect 14696 7172 14851 7228
rect 14907 7172 18433 7228
rect 18489 7172 18643 7228
rect 18699 7172 18854 7228
rect 18910 7172 19066 7228
rect 19122 7172 19277 7228
rect 19333 7172 19487 7228
rect 19543 7172 21911 7228
rect 21967 7172 22122 7228
rect 22178 7172 22333 7228
rect 22389 7172 22543 7228
rect 22599 7172 22754 7228
rect 22810 7172 22966 7228
rect 23022 7172 23177 7228
rect 23233 7172 23387 7228
rect 23443 7172 23598 7228
rect 23654 7172 23809 7228
rect 23865 7172 24219 7228
rect 0 7100 24219 7172
rect 6245 6874 9638 6875
rect 0 6795 3687 6861
rect 0 6739 2652 6795
rect 2708 6739 2832 6795
rect 2888 6788 3687 6795
rect 2888 6739 3414 6788
rect 0 6732 3414 6739
rect 3470 6732 3594 6788
rect 3650 6732 3687 6788
rect 6237 6836 9682 6874
rect 6237 6780 6273 6836
rect 6329 6780 9589 6836
rect 9645 6780 9682 6836
rect 6237 6741 9682 6780
rect 18154 6822 18284 6861
rect 18154 6766 18191 6822
rect 18247 6766 18284 6822
rect 0 6659 3687 6732
rect 18154 6643 18284 6766
rect 20631 6788 24219 6861
rect 20631 6732 20668 6788
rect 20724 6732 20848 6788
rect 20904 6732 21430 6788
rect 21486 6732 21610 6788
rect 21666 6732 24219 6788
rect 20631 6659 24219 6732
rect 7449 6605 18284 6643
rect 7449 6549 7486 6605
rect 7542 6549 7666 6605
rect 7722 6549 9370 6605
rect 9426 6604 18284 6605
rect 9426 6549 18191 6604
rect 7449 6548 18191 6549
rect 18247 6548 18284 6604
rect 7449 6510 18284 6548
rect 0 6328 24219 6401
rect 0 6272 3879 6328
rect 3935 6272 4090 6328
rect 4146 6272 4302 6328
rect 4358 6272 4513 6328
rect 4569 6272 7925 6328
rect 7981 6272 8136 6328
rect 8192 6272 8347 6328
rect 8403 6272 9848 6328
rect 9904 6272 10028 6328
rect 10084 6272 13385 6328
rect 13441 6272 13596 6328
rect 13652 6272 13808 6328
rect 13864 6272 14019 6328
rect 14075 6272 19758 6328
rect 19814 6272 19969 6328
rect 20025 6272 20181 6328
rect 20237 6272 20392 6328
rect 20448 6272 24219 6328
rect 0 6199 24219 6272
rect 7449 6052 18284 6090
rect 7449 6051 18191 6052
rect 7449 5995 7486 6051
rect 7542 5995 7666 6051
rect 7722 5995 9370 6051
rect 9426 5996 18191 6051
rect 18247 5996 18284 6052
rect 9426 5995 18284 5996
rect 7449 5957 18284 5995
rect 0 5868 3687 5941
rect 0 5861 3414 5868
rect 0 5805 2652 5861
rect 2708 5805 2832 5861
rect 2888 5812 3414 5861
rect 3470 5812 3594 5868
rect 3650 5812 3687 5868
rect 2888 5805 3687 5812
rect 0 5739 3687 5805
rect 6237 5820 9682 5859
rect 6237 5764 6273 5820
rect 6329 5764 9589 5820
rect 9645 5764 9682 5820
rect 6237 5726 9682 5764
rect 18154 5834 18284 5957
rect 18154 5778 18191 5834
rect 18247 5778 18284 5834
rect 18154 5739 18284 5778
rect 20631 5868 24219 5941
rect 20631 5812 20668 5868
rect 20724 5812 20848 5868
rect 20904 5812 21430 5868
rect 21486 5812 21610 5868
rect 21666 5812 24219 5868
rect 20631 5739 24219 5812
rect 6245 5725 9638 5726
rect 0 5428 24219 5500
rect 0 5372 449 5428
rect 505 5372 660 5428
rect 716 5372 871 5428
rect 927 5372 1081 5428
rect 1137 5372 1292 5428
rect 1348 5372 1504 5428
rect 1560 5372 1715 5428
rect 1771 5372 1925 5428
rect 1981 5372 2136 5428
rect 2192 5372 2347 5428
rect 2403 5372 4815 5428
rect 4871 5372 5025 5428
rect 5081 5372 5236 5428
rect 5292 5372 5448 5428
rect 5504 5372 5659 5428
rect 5715 5372 5869 5428
rect 5925 5372 8647 5428
rect 8703 5372 8827 5428
rect 8883 5372 14429 5428
rect 14485 5372 14640 5428
rect 14696 5372 14851 5428
rect 14907 5372 18433 5428
rect 18489 5372 18643 5428
rect 18699 5372 18854 5428
rect 18910 5372 19066 5428
rect 19122 5372 19277 5428
rect 19333 5372 19487 5428
rect 19543 5372 21911 5428
rect 21967 5372 22122 5428
rect 22178 5372 22333 5428
rect 22389 5372 22543 5428
rect 22599 5372 22754 5428
rect 22810 5372 22966 5428
rect 23022 5372 23177 5428
rect 23233 5372 23387 5428
rect 23443 5372 23598 5428
rect 23654 5372 23809 5428
rect 23865 5372 24219 5428
rect 0 5300 24219 5372
rect 6245 5074 9638 5075
rect 0 4995 3687 5061
rect 0 4939 2652 4995
rect 2708 4939 2832 4995
rect 2888 4988 3687 4995
rect 2888 4939 3414 4988
rect 0 4932 3414 4939
rect 3470 4932 3594 4988
rect 3650 4932 3687 4988
rect 6237 5036 9682 5074
rect 6237 4980 6273 5036
rect 6329 4980 9589 5036
rect 9645 4980 9682 5036
rect 6237 4941 9682 4980
rect 18154 5022 18284 5061
rect 18154 4966 18191 5022
rect 18247 4966 18284 5022
rect 0 4859 3687 4932
rect 18154 4843 18284 4966
rect 20631 4988 24219 5061
rect 20631 4932 20668 4988
rect 20724 4932 20848 4988
rect 20904 4932 21430 4988
rect 21486 4932 21610 4988
rect 21666 4932 24219 4988
rect 20631 4859 24219 4932
rect 7449 4805 18284 4843
rect 7449 4749 7486 4805
rect 7542 4749 7666 4805
rect 7722 4749 9370 4805
rect 9426 4804 18284 4805
rect 9426 4749 18191 4804
rect 7449 4748 18191 4749
rect 18247 4748 18284 4804
rect 7449 4710 18284 4748
rect 0 4528 24219 4601
rect 0 4472 3879 4528
rect 3935 4472 4090 4528
rect 4146 4472 4302 4528
rect 4358 4472 4513 4528
rect 4569 4472 7925 4528
rect 7981 4472 8136 4528
rect 8192 4472 8347 4528
rect 8403 4472 9848 4528
rect 9904 4472 10028 4528
rect 10084 4472 13385 4528
rect 13441 4472 13596 4528
rect 13652 4472 13808 4528
rect 13864 4472 14019 4528
rect 14075 4472 19758 4528
rect 19814 4472 19969 4528
rect 20025 4472 20181 4528
rect 20237 4472 20392 4528
rect 20448 4472 24219 4528
rect 0 4399 24219 4472
rect 7449 4252 18284 4290
rect 7449 4251 18191 4252
rect 7449 4195 7486 4251
rect 7542 4195 7666 4251
rect 7722 4195 9370 4251
rect 9426 4196 18191 4251
rect 18247 4196 18284 4252
rect 9426 4195 18284 4196
rect 7449 4157 18284 4195
rect 0 4068 3687 4141
rect 0 4061 3414 4068
rect 0 4005 2652 4061
rect 2708 4005 2832 4061
rect 2888 4012 3414 4061
rect 3470 4012 3594 4068
rect 3650 4012 3687 4068
rect 2888 4005 3687 4012
rect 0 3939 3687 4005
rect 6237 4020 9682 4059
rect 6237 3964 6273 4020
rect 6329 3964 9589 4020
rect 9645 3964 9682 4020
rect 6237 3926 9682 3964
rect 18154 4034 18284 4157
rect 18154 3978 18191 4034
rect 18247 3978 18284 4034
rect 18154 3939 18284 3978
rect 20631 4068 24219 4141
rect 20631 4012 20668 4068
rect 20724 4012 20848 4068
rect 20904 4012 21430 4068
rect 21486 4012 21610 4068
rect 21666 4012 24219 4068
rect 20631 3939 24219 4012
rect 6245 3925 9638 3926
rect 0 3628 24219 3700
rect 0 3572 449 3628
rect 505 3572 660 3628
rect 716 3572 871 3628
rect 927 3572 1081 3628
rect 1137 3572 1292 3628
rect 1348 3572 1504 3628
rect 1560 3572 1715 3628
rect 1771 3572 1925 3628
rect 1981 3572 2136 3628
rect 2192 3572 2347 3628
rect 2403 3572 4815 3628
rect 4871 3572 5025 3628
rect 5081 3572 5236 3628
rect 5292 3572 5448 3628
rect 5504 3572 5659 3628
rect 5715 3572 5869 3628
rect 5925 3572 8647 3628
rect 8703 3572 8827 3628
rect 8883 3572 14429 3628
rect 14485 3572 14640 3628
rect 14696 3572 14851 3628
rect 14907 3572 18433 3628
rect 18489 3572 18643 3628
rect 18699 3572 18854 3628
rect 18910 3572 19066 3628
rect 19122 3572 19277 3628
rect 19333 3572 19487 3628
rect 19543 3572 21911 3628
rect 21967 3572 22122 3628
rect 22178 3572 22333 3628
rect 22389 3572 22543 3628
rect 22599 3572 22754 3628
rect 22810 3572 22966 3628
rect 23022 3572 23177 3628
rect 23233 3572 23387 3628
rect 23443 3572 23598 3628
rect 23654 3572 23809 3628
rect 23865 3572 24219 3628
rect 0 3500 24219 3572
rect 6245 3274 9638 3275
rect 0 3195 3687 3261
rect 0 3139 2652 3195
rect 2708 3139 2832 3195
rect 2888 3188 3687 3195
rect 2888 3139 3414 3188
rect 0 3132 3414 3139
rect 3470 3132 3594 3188
rect 3650 3132 3687 3188
rect 6237 3236 9682 3274
rect 6237 3180 6273 3236
rect 6329 3180 9589 3236
rect 9645 3180 9682 3236
rect 6237 3141 9682 3180
rect 18154 3222 18284 3261
rect 18154 3166 18191 3222
rect 18247 3166 18284 3222
rect 0 3059 3687 3132
rect 18154 3043 18284 3166
rect 20631 3188 24219 3261
rect 20631 3132 20668 3188
rect 20724 3132 20848 3188
rect 20904 3132 21430 3188
rect 21486 3132 21610 3188
rect 21666 3132 24219 3188
rect 20631 3059 24219 3132
rect 7449 3005 18284 3043
rect 7449 2949 7486 3005
rect 7542 2949 7666 3005
rect 7722 2949 9370 3005
rect 9426 3004 18284 3005
rect 9426 2949 18191 3004
rect 7449 2948 18191 2949
rect 18247 2948 18284 3004
rect 7449 2910 18284 2948
rect 0 2728 24219 2801
rect 0 2672 3879 2728
rect 3935 2672 4090 2728
rect 4146 2672 4302 2728
rect 4358 2672 4513 2728
rect 4569 2672 7925 2728
rect 7981 2672 8136 2728
rect 8192 2672 8347 2728
rect 8403 2672 9848 2728
rect 9904 2672 10028 2728
rect 10084 2672 13385 2728
rect 13441 2672 13596 2728
rect 13652 2672 13808 2728
rect 13864 2672 14019 2728
rect 14075 2672 19758 2728
rect 19814 2672 19969 2728
rect 20025 2672 20181 2728
rect 20237 2672 20392 2728
rect 20448 2672 24219 2728
rect 0 2599 24219 2672
rect 7449 2452 18284 2490
rect 7449 2451 18191 2452
rect 7449 2395 7486 2451
rect 7542 2395 7666 2451
rect 7722 2395 9370 2451
rect 9426 2396 18191 2451
rect 18247 2396 18284 2452
rect 9426 2395 18284 2396
rect 7449 2357 18284 2395
rect 0 2268 3687 2341
rect 0 2261 3414 2268
rect 0 2205 2652 2261
rect 2708 2205 2832 2261
rect 2888 2212 3414 2261
rect 3470 2212 3594 2268
rect 3650 2212 3687 2268
rect 2888 2205 3687 2212
rect 0 2139 3687 2205
rect 6237 2220 9682 2259
rect 6237 2164 6273 2220
rect 6329 2164 9589 2220
rect 9645 2164 9682 2220
rect 6237 2126 9682 2164
rect 18154 2234 18284 2357
rect 18154 2178 18191 2234
rect 18247 2178 18284 2234
rect 18154 2139 18284 2178
rect 20631 2268 24219 2341
rect 20631 2212 20668 2268
rect 20724 2212 20848 2268
rect 20904 2212 21430 2268
rect 21486 2212 21610 2268
rect 21666 2212 24219 2268
rect 20631 2139 24219 2212
rect 6245 2125 9638 2126
rect 0 1828 24219 1900
rect 0 1772 449 1828
rect 505 1772 660 1828
rect 716 1772 871 1828
rect 927 1772 1081 1828
rect 1137 1772 1292 1828
rect 1348 1772 1504 1828
rect 1560 1772 1715 1828
rect 1771 1772 1925 1828
rect 1981 1772 2136 1828
rect 2192 1772 2347 1828
rect 2403 1772 4815 1828
rect 4871 1772 5025 1828
rect 5081 1772 5236 1828
rect 5292 1772 5448 1828
rect 5504 1772 5659 1828
rect 5715 1772 5869 1828
rect 5925 1772 8647 1828
rect 8703 1772 8827 1828
rect 8883 1772 14429 1828
rect 14485 1772 14640 1828
rect 14696 1772 14851 1828
rect 14907 1772 18433 1828
rect 18489 1772 18643 1828
rect 18699 1772 18854 1828
rect 18910 1772 19066 1828
rect 19122 1772 19277 1828
rect 19333 1772 19487 1828
rect 19543 1772 21911 1828
rect 21967 1772 22122 1828
rect 22178 1772 22333 1828
rect 22389 1772 22543 1828
rect 22599 1772 22754 1828
rect 22810 1772 22966 1828
rect 23022 1772 23177 1828
rect 23233 1772 23387 1828
rect 23443 1772 23598 1828
rect 23654 1772 23809 1828
rect 23865 1772 24219 1828
rect 0 1700 24219 1772
rect 6245 1474 9638 1475
rect 0 1395 3687 1461
rect 0 1339 2652 1395
rect 2708 1339 2832 1395
rect 2888 1388 3687 1395
rect 2888 1339 3414 1388
rect 0 1332 3414 1339
rect 3470 1332 3594 1388
rect 3650 1332 3687 1388
rect 6237 1436 9682 1474
rect 6237 1380 6273 1436
rect 6329 1380 9589 1436
rect 9645 1380 9682 1436
rect 6237 1341 9682 1380
rect 18154 1422 18284 1461
rect 18154 1366 18191 1422
rect 18247 1366 18284 1422
rect 0 1259 3687 1332
rect 18154 1243 18284 1366
rect 20631 1388 24219 1461
rect 20631 1332 20668 1388
rect 20724 1332 20848 1388
rect 20904 1332 21430 1388
rect 21486 1332 21610 1388
rect 21666 1332 24219 1388
rect 20631 1259 24219 1332
rect 7449 1205 18284 1243
rect 7449 1149 7486 1205
rect 7542 1149 7666 1205
rect 7722 1149 9370 1205
rect 9426 1204 18284 1205
rect 9426 1149 18191 1204
rect 7449 1148 18191 1149
rect 18247 1148 18284 1204
rect 7449 1110 18284 1148
rect 0 928 24219 1001
rect 0 872 3879 928
rect 3935 872 4090 928
rect 4146 872 4302 928
rect 4358 872 4513 928
rect 4569 872 7925 928
rect 7981 872 8136 928
rect 8192 872 8347 928
rect 8403 872 9848 928
rect 9904 872 10028 928
rect 10084 872 13385 928
rect 13441 872 13596 928
rect 13652 872 13808 928
rect 13864 872 14019 928
rect 14075 872 19758 928
rect 19814 872 19969 928
rect 20025 872 20181 928
rect 20237 872 20392 928
rect 20448 872 24219 928
rect 0 799 24219 872
rect 7449 652 18284 690
rect 7449 651 18191 652
rect 7449 595 7486 651
rect 7542 595 7666 651
rect 7722 595 9370 651
rect 9426 596 18191 651
rect 18247 596 18284 652
rect 9426 595 18284 596
rect 7449 557 18284 595
rect 0 468 3687 541
rect 0 461 3414 468
rect 0 405 2652 461
rect 2708 405 2832 461
rect 2888 412 3414 461
rect 3470 412 3594 468
rect 3650 412 3687 468
rect 2888 405 3687 412
rect 0 339 3687 405
rect 6237 420 9682 459
rect 6237 364 6273 420
rect 6329 364 9589 420
rect 9645 364 9682 420
rect 6237 326 9682 364
rect 18154 434 18284 557
rect 18154 378 18191 434
rect 18247 378 18284 434
rect 18154 339 18284 378
rect 20631 468 24219 541
rect 20631 412 20668 468
rect 20724 412 20848 468
rect 20904 412 21430 468
rect 21486 412 21610 468
rect 21666 412 24219 468
rect 20631 339 24219 412
rect 6245 325 9638 326
rect 0 28 24219 100
rect 0 -28 449 28
rect 505 -28 660 28
rect 716 -28 871 28
rect 927 -28 1081 28
rect 1137 -28 1292 28
rect 1348 -28 1504 28
rect 1560 -28 1715 28
rect 1771 -28 1925 28
rect 1981 -28 2136 28
rect 2192 -28 2347 28
rect 2403 -28 4815 28
rect 4871 -28 5025 28
rect 5081 -28 5236 28
rect 5292 -28 5448 28
rect 5504 -28 5659 28
rect 5715 -28 5869 28
rect 5925 -28 8647 28
rect 8703 -28 8827 28
rect 8883 -28 14429 28
rect 14485 -28 14640 28
rect 14696 -28 14851 28
rect 14907 -28 18433 28
rect 18489 -28 18643 28
rect 18699 -28 18854 28
rect 18910 -28 19066 28
rect 19122 -28 19277 28
rect 19333 -28 19487 28
rect 19543 -28 21911 28
rect 21967 -28 22122 28
rect 22178 -28 22333 28
rect 22389 -28 22543 28
rect 22599 -28 22754 28
rect 22810 -28 22966 28
rect 23022 -28 23177 28
rect 23233 -28 23387 28
rect 23443 -28 23598 28
rect 23654 -28 23809 28
rect 23865 -28 24219 28
rect 0 -100 24219 -28
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_0
timestamp 1698431365
transform 1 0 11558 0 1 1562
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_1
timestamp 1698431365
transform 1 0 11558 0 1 2038
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_2
timestamp 1698431365
transform 1 0 12691 0 1 7669
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_3
timestamp 1698431365
transform 1 0 12691 0 1 8531
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_4
timestamp 1698431365
transform 1 0 12691 0 1 9469
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_5
timestamp 1698431365
transform 1 0 12691 0 1 10331
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_6
timestamp 1698431365
transform 1 0 12691 0 1 11269
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_7
timestamp 1698431365
transform 1 0 12691 0 1 12131
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_8
timestamp 1698431365
transform 1 0 11558 0 1 14162
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_9
timestamp 1698431365
transform 1 0 11558 0 1 12362
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_10
timestamp 1698431365
transform 1 0 11558 0 1 10562
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_11
timestamp 1698431365
transform 1 0 11558 0 1 8762
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_12
timestamp 1698431365
transform 1 0 11558 0 1 6962
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_13
timestamp 1698431365
transform 1 0 11558 0 1 5162
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_14
timestamp 1698431365
transform 1 0 11558 0 1 3362
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_15
timestamp 1698431365
transform 1 0 13068 0 1 6731
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_16
timestamp 1698431365
transform 1 0 12691 0 1 13931
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_17
timestamp 1698431365
transform 1 0 12691 0 1 13069
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_18
timestamp 1698431365
transform 1 0 13068 0 1 469
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_19
timestamp 1698431365
transform 1 0 13068 0 1 1331
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_20
timestamp 1698431365
transform 1 0 13068 0 1 2269
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_21
timestamp 1698431365
transform 1 0 13068 0 1 3131
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_22
timestamp 1698431365
transform 1 0 13068 0 1 4069
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_23
timestamp 1698431365
transform 1 0 13068 0 1 4931
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_24
timestamp 1698431365
transform 1 0 13068 0 1 5869
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_25
timestamp 1698431365
transform 1 0 11558 0 1 12838
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_26
timestamp 1698431365
transform 1 0 11558 0 1 11038
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_27
timestamp 1698431365
transform 1 0 11558 0 1 9238
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_28
timestamp 1698431365
transform 1 0 11558 0 1 7438
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_29
timestamp 1698431365
transform 1 0 11558 0 1 5638
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_30
timestamp 1698431365
transform 1 0 11558 0 1 3838
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_31
timestamp 1698431365
transform 1 0 17864 0 1 578
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_32
timestamp 1698431365
transform 1 0 17487 0 1 1222
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_33
timestamp 1698431365
transform 1 0 17109 0 1 2378
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_34
timestamp 1698431365
transform 1 0 16731 0 1 3022
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_35
timestamp 1698431365
transform 1 0 16354 0 1 4178
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_36
timestamp 1698431365
transform 1 0 15976 0 1 4822
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_37
timestamp 1698431365
transform 1 0 15598 0 1 5978
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_38
timestamp 1698431365
transform 1 0 15220 0 1 6622
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_39
timestamp 1698431365
transform 1 0 15220 0 1 13822
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_40
timestamp 1698431365
transform 1 0 15598 0 1 13178
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_41
timestamp 1698431365
transform 1 0 15976 0 1 12022
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_42
timestamp 1698431365
transform 1 0 16354 0 1 11378
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_43
timestamp 1698431365
transform 1 0 16731 0 1 10222
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_44
timestamp 1698431365
transform 1 0 17109 0 1 9578
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_45
timestamp 1698431365
transform 1 0 17487 0 1 8422
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_46
timestamp 1698431365
transform 1 0 17864 0 1 7778
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_47
timestamp 1698431365
transform 1 0 11558 0 1 238
box 0 0 1 1
use xdec8_128x8m81  xdec8_128x8m81_0
timestamp 1698431365
transform 1 0 0 0 1 7200
box 1426 -1 22889 7201
use xdec8_128x8m81  xdec8_128x8m81_1
timestamp 1698431365
transform 1 0 0 0 1 0
box 1426 -1 22889 7201
<< labels >>
rlabel metal3 s 830 5840 830 5840 4 LWL[6]
port 1 nsew
rlabel metal3 s 830 6760 830 6760 4 LWL[7]
port 2 nsew
rlabel metal3 s 23423 13960 23423 13960 4 RWL[15]
port 3 nsew
rlabel metal3 s 23423 13040 23423 13040 4 RWL[14]
port 4 nsew
rlabel metal3 s 23423 12160 23423 12160 4 RWL[13]
port 5 nsew
rlabel metal3 s 23423 11240 23423 11240 4 RWL[12]
port 6 nsew
rlabel metal3 s 830 8560 830 8560 4 LWL[9]
port 7 nsew
rlabel metal3 s 830 7640 830 7640 4 LWL[8]
port 8 nsew
rlabel metal3 s 830 440 830 440 4 LWL[0]
port 9 nsew
rlabel metal3 s 830 1360 830 1360 4 LWL[1]
port 10 nsew
rlabel metal3 s 830 2240 830 2240 4 LWL[2]
port 11 nsew
rlabel metal3 s 830 3160 830 3160 4 LWL[3]
port 12 nsew
rlabel metal3 s 830 4040 830 4040 4 LWL[4]
port 13 nsew
rlabel metal3 s 830 4960 830 4960 4 LWL[5]
port 14 nsew
rlabel metal3 s 23423 10360 23423 10360 4 RWL[11]
port 15 nsew
rlabel metal3 s 23423 9440 23423 9440 4 RWL[10]
port 16 nsew
rlabel metal3 s 23423 8560 23423 8560 4 RWL[9]
port 17 nsew
rlabel metal3 s 23423 7640 23423 7640 4 RWL[8]
port 18 nsew
rlabel metal3 s 23423 6760 23423 6760 4 RWL[7]
port 19 nsew
rlabel metal3 s 23423 4960 23423 4960 4 RWL[5]
port 20 nsew
rlabel metal3 s 23423 3160 23423 3160 4 RWL[3]
port 21 nsew
rlabel metal3 s 23423 1360 23423 1360 4 RWL[1]
port 22 nsew
rlabel metal3 s 23423 440 23423 440 4 RWL[0]
port 23 nsew
rlabel metal3 s 23423 2240 23423 2240 4 RWL[2]
port 24 nsew
rlabel metal3 s 830 13960 830 13960 4 LWL[15]
port 25 nsew
rlabel metal3 s 830 13040 830 13040 4 LWL[14]
port 26 nsew
rlabel metal3 s 830 12160 830 12160 4 LWL[13]
port 27 nsew
rlabel metal3 s 830 11240 830 11240 4 LWL[12]
port 28 nsew
rlabel metal3 s 830 10360 830 10360 4 LWL[11]
port 29 nsew
rlabel metal3 s 830 9440 830 9440 4 LWL[10]
port 30 nsew
rlabel metal3 s 23423 4040 23423 4040 4 RWL[4]
port 31 nsew
rlabel metal3 s 23423 5840 23423 5840 4 RWL[6]
port 32 nsew
rlabel metal2 s 17109 238 17109 238 4 xa[2]
port 33 nsew
rlabel metal2 s 6900 45 6900 45 4 men
port 34 nsew
rlabel metal2 s 17864 238 17864 238 4 xa[0]
port 35 nsew
rlabel metal2 s 16731 238 16731 238 4 xa[3]
port 36 nsew
rlabel metal2 s 16354 238 16354 238 4 xa[4]
port 37 nsew
rlabel metal2 s 15976 238 15976 238 4 xa[5]
port 38 nsew
rlabel metal2 s 15598 238 15598 238 4 xa[6]
port 39 nsew
rlabel metal2 s 15220 238 15220 238 4 xa[7]
port 40 nsew
rlabel metal2 s 11935 238 11935 238 4 xb[3]
port 41 nsew
rlabel metal2 s 12313 238 12313 238 4 xb[2]
port 42 nsew
rlabel metal2 s 12691 238 12691 238 4 xb[1]
port 43 nsew
rlabel metal2 s 13068 238 13068 238 4 xb[0]
port 44 nsew
rlabel metal2 s 11558 238 11558 238 4 xc
port 45 nsew
rlabel metal2 s 17487 238 17487 238 4 xa[1]
port 46 nsew
<< properties >>
string GDS_END 1698910
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 1691600
<< end >>
