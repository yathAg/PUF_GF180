magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< nwell >>
rect 2209 5116 4648 6727
rect 2137 5115 4648 5116
rect 2101 4660 4696 5115
rect 2780 736 4529 1473
rect 2815 373 4520 736
<< mvnmos >>
rect 2332 3317 2452 3999
rect 2556 3317 2676 3999
rect 2780 3317 2900 3999
rect 3004 3317 3124 3999
rect 3228 3317 3348 3999
rect 3452 3317 3572 3999
rect 3676 3317 3796 3999
rect 3900 3317 4020 3999
rect 4124 3317 4244 3999
rect 4348 3317 4468 3999
rect 2589 2510 2709 3078
rect 2813 2510 2933 3078
rect 3037 2510 3157 3078
rect 3261 2510 3381 3078
rect 3485 2510 3605 3078
rect 3709 2510 3829 3078
rect 3933 2510 4053 3078
rect 4157 2510 4277 3078
rect 3034 1702 3154 2156
rect 3482 1702 3602 2156
rect 3706 1702 3826 2156
rect 3930 1702 4050 2156
rect 4154 1702 4274 2156
<< mvpmos >>
rect 2464 6132 2584 6586
rect 2688 6132 2808 6586
rect 3151 6132 3271 6586
rect 3375 6132 3495 6586
rect 3599 6132 3719 6586
rect 4049 6132 4169 6586
rect 4273 6132 4393 6586
rect 2464 5266 2584 5720
rect 2688 5266 2808 5720
rect 3375 5266 3495 5720
rect 4049 5266 4169 5720
rect 4273 5266 4393 5720
rect 2797 4802 2917 4984
rect 3021 4802 3141 4984
rect 3245 4802 3365 4984
rect 3469 4802 3589 4984
rect 3693 4802 3813 4984
rect 3917 4802 4037 4984
rect 3034 877 3154 1331
rect 3258 877 3378 1331
rect 3482 877 3602 1331
rect 3706 877 3826 1331
rect 3930 877 4050 1331
rect 4154 877 4274 1331
<< mvndiff >>
rect 2244 3986 2332 3999
rect 2244 3330 2257 3986
rect 2303 3330 2332 3986
rect 2244 3317 2332 3330
rect 2452 3986 2556 3999
rect 2452 3330 2481 3986
rect 2527 3330 2556 3986
rect 2452 3317 2556 3330
rect 2676 3986 2780 3999
rect 2676 3330 2705 3986
rect 2751 3330 2780 3986
rect 2676 3317 2780 3330
rect 2900 3986 3004 3999
rect 2900 3330 2929 3986
rect 2975 3330 3004 3986
rect 2900 3317 3004 3330
rect 3124 3986 3228 3999
rect 3124 3330 3153 3986
rect 3199 3330 3228 3986
rect 3124 3317 3228 3330
rect 3348 3986 3452 3999
rect 3348 3330 3377 3986
rect 3423 3330 3452 3986
rect 3348 3317 3452 3330
rect 3572 3986 3676 3999
rect 3572 3330 3601 3986
rect 3647 3330 3676 3986
rect 3572 3317 3676 3330
rect 3796 3986 3900 3999
rect 3796 3330 3825 3986
rect 3871 3330 3900 3986
rect 3796 3317 3900 3330
rect 4020 3986 4124 3999
rect 4020 3330 4049 3986
rect 4095 3330 4124 3986
rect 4020 3317 4124 3330
rect 4244 3986 4348 3999
rect 4244 3330 4273 3986
rect 4319 3330 4348 3986
rect 4244 3317 4348 3330
rect 4468 3986 4556 3999
rect 4468 3330 4497 3986
rect 4543 3330 4556 3986
rect 4468 3317 4556 3330
rect 2501 3065 2589 3078
rect 2501 3019 2514 3065
rect 2560 3019 2589 3065
rect 2501 2941 2589 3019
rect 2501 2895 2514 2941
rect 2560 2895 2589 2941
rect 2501 2817 2589 2895
rect 2501 2771 2514 2817
rect 2560 2771 2589 2817
rect 2501 2693 2589 2771
rect 2501 2647 2514 2693
rect 2560 2647 2589 2693
rect 2501 2569 2589 2647
rect 2501 2523 2514 2569
rect 2560 2523 2589 2569
rect 2501 2510 2589 2523
rect 2709 3065 2813 3078
rect 2709 3019 2738 3065
rect 2784 3019 2813 3065
rect 2709 2941 2813 3019
rect 2709 2895 2738 2941
rect 2784 2895 2813 2941
rect 2709 2817 2813 2895
rect 2709 2771 2738 2817
rect 2784 2771 2813 2817
rect 2709 2693 2813 2771
rect 2709 2647 2738 2693
rect 2784 2647 2813 2693
rect 2709 2569 2813 2647
rect 2709 2523 2738 2569
rect 2784 2523 2813 2569
rect 2709 2510 2813 2523
rect 2933 3065 3037 3078
rect 2933 3019 2962 3065
rect 3008 3019 3037 3065
rect 2933 2941 3037 3019
rect 2933 2895 2962 2941
rect 3008 2895 3037 2941
rect 2933 2817 3037 2895
rect 2933 2771 2962 2817
rect 3008 2771 3037 2817
rect 2933 2693 3037 2771
rect 2933 2647 2962 2693
rect 3008 2647 3037 2693
rect 2933 2569 3037 2647
rect 2933 2523 2962 2569
rect 3008 2523 3037 2569
rect 2933 2510 3037 2523
rect 3157 3065 3261 3078
rect 3157 3019 3186 3065
rect 3232 3019 3261 3065
rect 3157 2941 3261 3019
rect 3157 2895 3186 2941
rect 3232 2895 3261 2941
rect 3157 2817 3261 2895
rect 3157 2771 3186 2817
rect 3232 2771 3261 2817
rect 3157 2693 3261 2771
rect 3157 2647 3186 2693
rect 3232 2647 3261 2693
rect 3157 2569 3261 2647
rect 3157 2523 3186 2569
rect 3232 2523 3261 2569
rect 3157 2510 3261 2523
rect 3381 3065 3485 3078
rect 3381 3019 3410 3065
rect 3456 3019 3485 3065
rect 3381 2941 3485 3019
rect 3381 2895 3410 2941
rect 3456 2895 3485 2941
rect 3381 2817 3485 2895
rect 3381 2771 3410 2817
rect 3456 2771 3485 2817
rect 3381 2693 3485 2771
rect 3381 2647 3410 2693
rect 3456 2647 3485 2693
rect 3381 2569 3485 2647
rect 3381 2523 3410 2569
rect 3456 2523 3485 2569
rect 3381 2510 3485 2523
rect 3605 3065 3709 3078
rect 3605 3019 3634 3065
rect 3680 3019 3709 3065
rect 3605 2941 3709 3019
rect 3605 2895 3634 2941
rect 3680 2895 3709 2941
rect 3605 2817 3709 2895
rect 3605 2771 3634 2817
rect 3680 2771 3709 2817
rect 3605 2693 3709 2771
rect 3605 2647 3634 2693
rect 3680 2647 3709 2693
rect 3605 2569 3709 2647
rect 3605 2523 3634 2569
rect 3680 2523 3709 2569
rect 3605 2510 3709 2523
rect 3829 3065 3933 3078
rect 3829 3019 3858 3065
rect 3904 3019 3933 3065
rect 3829 2941 3933 3019
rect 3829 2895 3858 2941
rect 3904 2895 3933 2941
rect 3829 2817 3933 2895
rect 3829 2771 3858 2817
rect 3904 2771 3933 2817
rect 3829 2693 3933 2771
rect 3829 2647 3858 2693
rect 3904 2647 3933 2693
rect 3829 2569 3933 2647
rect 3829 2523 3858 2569
rect 3904 2523 3933 2569
rect 3829 2510 3933 2523
rect 4053 3065 4157 3078
rect 4053 3019 4082 3065
rect 4128 3019 4157 3065
rect 4053 2941 4157 3019
rect 4053 2895 4082 2941
rect 4128 2895 4157 2941
rect 4053 2817 4157 2895
rect 4053 2771 4082 2817
rect 4128 2771 4157 2817
rect 4053 2693 4157 2771
rect 4053 2647 4082 2693
rect 4128 2647 4157 2693
rect 4053 2569 4157 2647
rect 4053 2523 4082 2569
rect 4128 2523 4157 2569
rect 4053 2510 4157 2523
rect 4277 3065 4365 3078
rect 4277 3019 4306 3065
rect 4352 3019 4365 3065
rect 4277 2941 4365 3019
rect 4277 2895 4306 2941
rect 4352 2895 4365 2941
rect 4277 2817 4365 2895
rect 4277 2771 4306 2817
rect 4352 2771 4365 2817
rect 4277 2693 4365 2771
rect 4277 2647 4306 2693
rect 4352 2647 4365 2693
rect 4277 2569 4365 2647
rect 4277 2523 4306 2569
rect 4352 2523 4365 2569
rect 4277 2510 4365 2523
rect 2946 2143 3034 2156
rect 2946 2097 2959 2143
rect 3005 2097 3034 2143
rect 2946 2015 3034 2097
rect 2946 1969 2959 2015
rect 3005 1969 3034 2015
rect 2946 1888 3034 1969
rect 2946 1842 2959 1888
rect 3005 1842 3034 1888
rect 2946 1761 3034 1842
rect 2946 1715 2959 1761
rect 3005 1715 3034 1761
rect 2946 1702 3034 1715
rect 3154 2143 3242 2156
rect 3154 2097 3183 2143
rect 3229 2097 3242 2143
rect 3154 2015 3242 2097
rect 3154 1969 3183 2015
rect 3229 1969 3242 2015
rect 3154 1888 3242 1969
rect 3154 1842 3183 1888
rect 3229 1842 3242 1888
rect 3154 1761 3242 1842
rect 3154 1715 3183 1761
rect 3229 1715 3242 1761
rect 3154 1702 3242 1715
rect 3394 2143 3482 2156
rect 3394 2097 3407 2143
rect 3453 2097 3482 2143
rect 3394 2015 3482 2097
rect 3394 1969 3407 2015
rect 3453 1969 3482 2015
rect 3394 1888 3482 1969
rect 3394 1842 3407 1888
rect 3453 1842 3482 1888
rect 3394 1761 3482 1842
rect 3394 1715 3407 1761
rect 3453 1715 3482 1761
rect 3394 1702 3482 1715
rect 3602 2143 3706 2156
rect 3602 2097 3631 2143
rect 3677 2097 3706 2143
rect 3602 2015 3706 2097
rect 3602 1969 3631 2015
rect 3677 1969 3706 2015
rect 3602 1888 3706 1969
rect 3602 1842 3631 1888
rect 3677 1842 3706 1888
rect 3602 1761 3706 1842
rect 3602 1715 3631 1761
rect 3677 1715 3706 1761
rect 3602 1702 3706 1715
rect 3826 2143 3930 2156
rect 3826 2097 3855 2143
rect 3901 2097 3930 2143
rect 3826 2015 3930 2097
rect 3826 1969 3855 2015
rect 3901 1969 3930 2015
rect 3826 1888 3930 1969
rect 3826 1842 3855 1888
rect 3901 1842 3930 1888
rect 3826 1761 3930 1842
rect 3826 1715 3855 1761
rect 3901 1715 3930 1761
rect 3826 1702 3930 1715
rect 4050 2143 4154 2156
rect 4050 2097 4079 2143
rect 4125 2097 4154 2143
rect 4050 2015 4154 2097
rect 4050 1969 4079 2015
rect 4125 1969 4154 2015
rect 4050 1888 4154 1969
rect 4050 1842 4079 1888
rect 4125 1842 4154 1888
rect 4050 1761 4154 1842
rect 4050 1715 4079 1761
rect 4125 1715 4154 1761
rect 4050 1702 4154 1715
rect 4274 2143 4362 2156
rect 4274 2097 4303 2143
rect 4349 2097 4362 2143
rect 4274 2015 4362 2097
rect 4274 1969 4303 2015
rect 4349 1969 4362 2015
rect 4274 1888 4362 1969
rect 4274 1842 4303 1888
rect 4349 1842 4362 1888
rect 4274 1761 4362 1842
rect 4274 1715 4303 1761
rect 4349 1715 4362 1761
rect 4274 1702 4362 1715
<< mvpdiff >>
rect 2376 6573 2464 6586
rect 2376 6527 2389 6573
rect 2435 6527 2464 6573
rect 2376 6446 2464 6527
rect 2376 6400 2389 6446
rect 2435 6400 2464 6446
rect 2376 6319 2464 6400
rect 2376 6273 2389 6319
rect 2435 6273 2464 6319
rect 2376 6191 2464 6273
rect 2376 6145 2389 6191
rect 2435 6145 2464 6191
rect 2376 6132 2464 6145
rect 2584 6573 2688 6586
rect 2584 6527 2613 6573
rect 2659 6527 2688 6573
rect 2584 6446 2688 6527
rect 2584 6400 2613 6446
rect 2659 6400 2688 6446
rect 2584 6319 2688 6400
rect 2584 6273 2613 6319
rect 2659 6273 2688 6319
rect 2584 6191 2688 6273
rect 2584 6145 2613 6191
rect 2659 6145 2688 6191
rect 2584 6132 2688 6145
rect 2808 6573 2896 6586
rect 2808 6527 2837 6573
rect 2883 6527 2896 6573
rect 2808 6446 2896 6527
rect 2808 6400 2837 6446
rect 2883 6400 2896 6446
rect 2808 6319 2896 6400
rect 2808 6273 2837 6319
rect 2883 6273 2896 6319
rect 2808 6191 2896 6273
rect 2808 6145 2837 6191
rect 2883 6145 2896 6191
rect 2808 6132 2896 6145
rect 3063 6573 3151 6586
rect 3063 6527 3076 6573
rect 3122 6527 3151 6573
rect 3063 6446 3151 6527
rect 3063 6400 3076 6446
rect 3122 6400 3151 6446
rect 3063 6319 3151 6400
rect 3063 6273 3076 6319
rect 3122 6273 3151 6319
rect 3063 6191 3151 6273
rect 3063 6145 3076 6191
rect 3122 6145 3151 6191
rect 3063 6132 3151 6145
rect 3271 6573 3375 6586
rect 3271 6527 3300 6573
rect 3346 6527 3375 6573
rect 3271 6446 3375 6527
rect 3271 6400 3300 6446
rect 3346 6400 3375 6446
rect 3271 6319 3375 6400
rect 3271 6273 3300 6319
rect 3346 6273 3375 6319
rect 3271 6191 3375 6273
rect 3271 6145 3300 6191
rect 3346 6145 3375 6191
rect 3271 6132 3375 6145
rect 3495 6573 3599 6586
rect 3495 6527 3524 6573
rect 3570 6527 3599 6573
rect 3495 6446 3599 6527
rect 3495 6400 3524 6446
rect 3570 6400 3599 6446
rect 3495 6319 3599 6400
rect 3495 6273 3524 6319
rect 3570 6273 3599 6319
rect 3495 6191 3599 6273
rect 3495 6145 3524 6191
rect 3570 6145 3599 6191
rect 3495 6132 3599 6145
rect 3719 6573 3807 6586
rect 3719 6527 3748 6573
rect 3794 6527 3807 6573
rect 3719 6446 3807 6527
rect 3719 6400 3748 6446
rect 3794 6400 3807 6446
rect 3719 6319 3807 6400
rect 3719 6273 3748 6319
rect 3794 6273 3807 6319
rect 3719 6191 3807 6273
rect 3719 6145 3748 6191
rect 3794 6145 3807 6191
rect 3719 6132 3807 6145
rect 3961 6573 4049 6586
rect 3961 6527 3974 6573
rect 4020 6527 4049 6573
rect 3961 6446 4049 6527
rect 3961 6400 3974 6446
rect 4020 6400 4049 6446
rect 3961 6319 4049 6400
rect 3961 6273 3974 6319
rect 4020 6273 4049 6319
rect 3961 6191 4049 6273
rect 3961 6145 3974 6191
rect 4020 6145 4049 6191
rect 3961 6132 4049 6145
rect 4169 6573 4273 6586
rect 4169 6527 4198 6573
rect 4244 6527 4273 6573
rect 4169 6446 4273 6527
rect 4169 6400 4198 6446
rect 4244 6400 4273 6446
rect 4169 6319 4273 6400
rect 4169 6273 4198 6319
rect 4244 6273 4273 6319
rect 4169 6191 4273 6273
rect 4169 6145 4198 6191
rect 4244 6145 4273 6191
rect 4169 6132 4273 6145
rect 4393 6573 4481 6586
rect 4393 6527 4422 6573
rect 4468 6527 4481 6573
rect 4393 6446 4481 6527
rect 4393 6400 4422 6446
rect 4468 6400 4481 6446
rect 4393 6319 4481 6400
rect 4393 6273 4422 6319
rect 4468 6273 4481 6319
rect 4393 6191 4481 6273
rect 4393 6145 4422 6191
rect 4468 6145 4481 6191
rect 4393 6132 4481 6145
rect 2376 5707 2464 5720
rect 2376 5661 2389 5707
rect 2435 5661 2464 5707
rect 2376 5580 2464 5661
rect 2376 5534 2389 5580
rect 2435 5534 2464 5580
rect 2376 5453 2464 5534
rect 2376 5407 2389 5453
rect 2435 5407 2464 5453
rect 2376 5325 2464 5407
rect 2376 5279 2389 5325
rect 2435 5279 2464 5325
rect 2376 5266 2464 5279
rect 2584 5707 2688 5720
rect 2584 5661 2613 5707
rect 2659 5661 2688 5707
rect 2584 5580 2688 5661
rect 2584 5534 2613 5580
rect 2659 5534 2688 5580
rect 2584 5453 2688 5534
rect 2584 5407 2613 5453
rect 2659 5407 2688 5453
rect 2584 5325 2688 5407
rect 2584 5279 2613 5325
rect 2659 5279 2688 5325
rect 2584 5266 2688 5279
rect 2808 5707 2896 5720
rect 2808 5661 2837 5707
rect 2883 5661 2896 5707
rect 2808 5580 2896 5661
rect 2808 5534 2837 5580
rect 2883 5534 2896 5580
rect 2808 5453 2896 5534
rect 2808 5407 2837 5453
rect 2883 5407 2896 5453
rect 2808 5325 2896 5407
rect 2808 5279 2837 5325
rect 2883 5279 2896 5325
rect 2808 5266 2896 5279
rect 3287 5707 3375 5720
rect 3287 5661 3300 5707
rect 3346 5661 3375 5707
rect 3287 5580 3375 5661
rect 3287 5534 3300 5580
rect 3346 5534 3375 5580
rect 3287 5453 3375 5534
rect 3287 5407 3300 5453
rect 3346 5407 3375 5453
rect 3287 5325 3375 5407
rect 3287 5279 3300 5325
rect 3346 5279 3375 5325
rect 3287 5266 3375 5279
rect 3495 5707 3583 5720
rect 3495 5661 3524 5707
rect 3570 5661 3583 5707
rect 3495 5580 3583 5661
rect 3495 5534 3524 5580
rect 3570 5534 3583 5580
rect 3495 5453 3583 5534
rect 3495 5407 3524 5453
rect 3570 5407 3583 5453
rect 3495 5325 3583 5407
rect 3495 5279 3524 5325
rect 3570 5279 3583 5325
rect 3495 5266 3583 5279
rect 3961 5707 4049 5720
rect 3961 5661 3974 5707
rect 4020 5661 4049 5707
rect 3961 5580 4049 5661
rect 3961 5534 3974 5580
rect 4020 5534 4049 5580
rect 3961 5453 4049 5534
rect 3961 5407 3974 5453
rect 4020 5407 4049 5453
rect 3961 5325 4049 5407
rect 3961 5279 3974 5325
rect 4020 5279 4049 5325
rect 3961 5266 4049 5279
rect 4169 5707 4273 5720
rect 4169 5661 4198 5707
rect 4244 5661 4273 5707
rect 4169 5580 4273 5661
rect 4169 5534 4198 5580
rect 4244 5534 4273 5580
rect 4169 5453 4273 5534
rect 4169 5407 4198 5453
rect 4244 5407 4273 5453
rect 4169 5325 4273 5407
rect 4169 5279 4198 5325
rect 4244 5279 4273 5325
rect 4169 5266 4273 5279
rect 4393 5707 4481 5720
rect 4393 5661 4422 5707
rect 4468 5661 4481 5707
rect 4393 5580 4481 5661
rect 4393 5534 4422 5580
rect 4468 5534 4481 5580
rect 4393 5453 4481 5534
rect 4393 5407 4422 5453
rect 4468 5407 4481 5453
rect 4393 5325 4481 5407
rect 4393 5279 4422 5325
rect 4468 5279 4481 5325
rect 4393 5266 4481 5279
rect 2709 4971 2797 4984
rect 2709 4925 2722 4971
rect 2768 4925 2797 4971
rect 2709 4861 2797 4925
rect 2709 4815 2722 4861
rect 2768 4815 2797 4861
rect 2709 4802 2797 4815
rect 2917 4971 3021 4984
rect 2917 4925 2946 4971
rect 2992 4925 3021 4971
rect 2917 4861 3021 4925
rect 2917 4815 2946 4861
rect 2992 4815 3021 4861
rect 2917 4802 3021 4815
rect 3141 4971 3245 4984
rect 3141 4925 3170 4971
rect 3216 4925 3245 4971
rect 3141 4861 3245 4925
rect 3141 4815 3170 4861
rect 3216 4815 3245 4861
rect 3141 4802 3245 4815
rect 3365 4971 3469 4984
rect 3365 4925 3394 4971
rect 3440 4925 3469 4971
rect 3365 4861 3469 4925
rect 3365 4815 3394 4861
rect 3440 4815 3469 4861
rect 3365 4802 3469 4815
rect 3589 4971 3693 4984
rect 3589 4925 3618 4971
rect 3664 4925 3693 4971
rect 3589 4861 3693 4925
rect 3589 4815 3618 4861
rect 3664 4815 3693 4861
rect 3589 4802 3693 4815
rect 3813 4971 3917 4984
rect 3813 4925 3842 4971
rect 3888 4925 3917 4971
rect 3813 4861 3917 4925
rect 3813 4815 3842 4861
rect 3888 4815 3917 4861
rect 3813 4802 3917 4815
rect 4037 4971 4125 4984
rect 4037 4925 4066 4971
rect 4112 4925 4125 4971
rect 4037 4861 4125 4925
rect 4037 4815 4066 4861
rect 4112 4815 4125 4861
rect 4037 4802 4125 4815
rect 2946 1318 3034 1331
rect 2946 1272 2959 1318
rect 3005 1272 3034 1318
rect 2946 1190 3034 1272
rect 2946 1144 2959 1190
rect 3005 1144 3034 1190
rect 2946 1063 3034 1144
rect 2946 1017 2959 1063
rect 3005 1017 3034 1063
rect 2946 936 3034 1017
rect 2946 890 2959 936
rect 3005 890 3034 936
rect 2946 877 3034 890
rect 3154 1318 3258 1331
rect 3154 1272 3183 1318
rect 3229 1272 3258 1318
rect 3154 1190 3258 1272
rect 3154 1144 3183 1190
rect 3229 1144 3258 1190
rect 3154 1063 3258 1144
rect 3154 1017 3183 1063
rect 3229 1017 3258 1063
rect 3154 936 3258 1017
rect 3154 890 3183 936
rect 3229 890 3258 936
rect 3154 877 3258 890
rect 3378 1318 3482 1331
rect 3378 1272 3407 1318
rect 3453 1272 3482 1318
rect 3378 1190 3482 1272
rect 3378 1144 3407 1190
rect 3453 1144 3482 1190
rect 3378 1063 3482 1144
rect 3378 1017 3407 1063
rect 3453 1017 3482 1063
rect 3378 936 3482 1017
rect 3378 890 3407 936
rect 3453 890 3482 936
rect 3378 877 3482 890
rect 3602 1318 3706 1331
rect 3602 1272 3631 1318
rect 3677 1272 3706 1318
rect 3602 1190 3706 1272
rect 3602 1144 3631 1190
rect 3677 1144 3706 1190
rect 3602 1063 3706 1144
rect 3602 1017 3631 1063
rect 3677 1017 3706 1063
rect 3602 936 3706 1017
rect 3602 890 3631 936
rect 3677 890 3706 936
rect 3602 877 3706 890
rect 3826 1318 3930 1331
rect 3826 1272 3855 1318
rect 3901 1272 3930 1318
rect 3826 1190 3930 1272
rect 3826 1144 3855 1190
rect 3901 1144 3930 1190
rect 3826 1063 3930 1144
rect 3826 1017 3855 1063
rect 3901 1017 3930 1063
rect 3826 936 3930 1017
rect 3826 890 3855 936
rect 3901 890 3930 936
rect 3826 877 3930 890
rect 4050 1318 4154 1331
rect 4050 1272 4079 1318
rect 4125 1272 4154 1318
rect 4050 1190 4154 1272
rect 4050 1144 4079 1190
rect 4125 1144 4154 1190
rect 4050 1063 4154 1144
rect 4050 1017 4079 1063
rect 4125 1017 4154 1063
rect 4050 936 4154 1017
rect 4050 890 4079 936
rect 4125 890 4154 936
rect 4050 877 4154 890
rect 4274 1318 4362 1331
rect 4274 1272 4303 1318
rect 4349 1272 4362 1318
rect 4274 1190 4362 1272
rect 4274 1144 4303 1190
rect 4349 1144 4362 1190
rect 4274 1063 4362 1144
rect 4274 1017 4303 1063
rect 4349 1017 4362 1063
rect 4274 936 4362 1017
rect 4274 890 4303 936
rect 4349 890 4362 936
rect 4274 877 4362 890
<< mvndiffc >>
rect 2257 3330 2303 3986
rect 2481 3330 2527 3986
rect 2705 3330 2751 3986
rect 2929 3330 2975 3986
rect 3153 3330 3199 3986
rect 3377 3330 3423 3986
rect 3601 3330 3647 3986
rect 3825 3330 3871 3986
rect 4049 3330 4095 3986
rect 4273 3330 4319 3986
rect 4497 3330 4543 3986
rect 2514 3019 2560 3065
rect 2514 2895 2560 2941
rect 2514 2771 2560 2817
rect 2514 2647 2560 2693
rect 2514 2523 2560 2569
rect 2738 3019 2784 3065
rect 2738 2895 2784 2941
rect 2738 2771 2784 2817
rect 2738 2647 2784 2693
rect 2738 2523 2784 2569
rect 2962 3019 3008 3065
rect 2962 2895 3008 2941
rect 2962 2771 3008 2817
rect 2962 2647 3008 2693
rect 2962 2523 3008 2569
rect 3186 3019 3232 3065
rect 3186 2895 3232 2941
rect 3186 2771 3232 2817
rect 3186 2647 3232 2693
rect 3186 2523 3232 2569
rect 3410 3019 3456 3065
rect 3410 2895 3456 2941
rect 3410 2771 3456 2817
rect 3410 2647 3456 2693
rect 3410 2523 3456 2569
rect 3634 3019 3680 3065
rect 3634 2895 3680 2941
rect 3634 2771 3680 2817
rect 3634 2647 3680 2693
rect 3634 2523 3680 2569
rect 3858 3019 3904 3065
rect 3858 2895 3904 2941
rect 3858 2771 3904 2817
rect 3858 2647 3904 2693
rect 3858 2523 3904 2569
rect 4082 3019 4128 3065
rect 4082 2895 4128 2941
rect 4082 2771 4128 2817
rect 4082 2647 4128 2693
rect 4082 2523 4128 2569
rect 4306 3019 4352 3065
rect 4306 2895 4352 2941
rect 4306 2771 4352 2817
rect 4306 2647 4352 2693
rect 4306 2523 4352 2569
rect 2959 2097 3005 2143
rect 2959 1969 3005 2015
rect 2959 1842 3005 1888
rect 2959 1715 3005 1761
rect 3183 2097 3229 2143
rect 3183 1969 3229 2015
rect 3183 1842 3229 1888
rect 3183 1715 3229 1761
rect 3407 2097 3453 2143
rect 3407 1969 3453 2015
rect 3407 1842 3453 1888
rect 3407 1715 3453 1761
rect 3631 2097 3677 2143
rect 3631 1969 3677 2015
rect 3631 1842 3677 1888
rect 3631 1715 3677 1761
rect 3855 2097 3901 2143
rect 3855 1969 3901 2015
rect 3855 1842 3901 1888
rect 3855 1715 3901 1761
rect 4079 2097 4125 2143
rect 4079 1969 4125 2015
rect 4079 1842 4125 1888
rect 4079 1715 4125 1761
rect 4303 2097 4349 2143
rect 4303 1969 4349 2015
rect 4303 1842 4349 1888
rect 4303 1715 4349 1761
<< mvpdiffc >>
rect 2389 6527 2435 6573
rect 2389 6400 2435 6446
rect 2389 6273 2435 6319
rect 2389 6145 2435 6191
rect 2613 6527 2659 6573
rect 2613 6400 2659 6446
rect 2613 6273 2659 6319
rect 2613 6145 2659 6191
rect 2837 6527 2883 6573
rect 2837 6400 2883 6446
rect 2837 6273 2883 6319
rect 2837 6145 2883 6191
rect 3076 6527 3122 6573
rect 3076 6400 3122 6446
rect 3076 6273 3122 6319
rect 3076 6145 3122 6191
rect 3300 6527 3346 6573
rect 3300 6400 3346 6446
rect 3300 6273 3346 6319
rect 3300 6145 3346 6191
rect 3524 6527 3570 6573
rect 3524 6400 3570 6446
rect 3524 6273 3570 6319
rect 3524 6145 3570 6191
rect 3748 6527 3794 6573
rect 3748 6400 3794 6446
rect 3748 6273 3794 6319
rect 3748 6145 3794 6191
rect 3974 6527 4020 6573
rect 3974 6400 4020 6446
rect 3974 6273 4020 6319
rect 3974 6145 4020 6191
rect 4198 6527 4244 6573
rect 4198 6400 4244 6446
rect 4198 6273 4244 6319
rect 4198 6145 4244 6191
rect 4422 6527 4468 6573
rect 4422 6400 4468 6446
rect 4422 6273 4468 6319
rect 4422 6145 4468 6191
rect 2389 5661 2435 5707
rect 2389 5534 2435 5580
rect 2389 5407 2435 5453
rect 2389 5279 2435 5325
rect 2613 5661 2659 5707
rect 2613 5534 2659 5580
rect 2613 5407 2659 5453
rect 2613 5279 2659 5325
rect 2837 5661 2883 5707
rect 2837 5534 2883 5580
rect 2837 5407 2883 5453
rect 2837 5279 2883 5325
rect 3300 5661 3346 5707
rect 3300 5534 3346 5580
rect 3300 5407 3346 5453
rect 3300 5279 3346 5325
rect 3524 5661 3570 5707
rect 3524 5534 3570 5580
rect 3524 5407 3570 5453
rect 3524 5279 3570 5325
rect 3974 5661 4020 5707
rect 3974 5534 4020 5580
rect 3974 5407 4020 5453
rect 3974 5279 4020 5325
rect 4198 5661 4244 5707
rect 4198 5534 4244 5580
rect 4198 5407 4244 5453
rect 4198 5279 4244 5325
rect 4422 5661 4468 5707
rect 4422 5534 4468 5580
rect 4422 5407 4468 5453
rect 4422 5279 4468 5325
rect 2722 4925 2768 4971
rect 2722 4815 2768 4861
rect 2946 4925 2992 4971
rect 2946 4815 2992 4861
rect 3170 4925 3216 4971
rect 3170 4815 3216 4861
rect 3394 4925 3440 4971
rect 3394 4815 3440 4861
rect 3618 4925 3664 4971
rect 3618 4815 3664 4861
rect 3842 4925 3888 4971
rect 3842 4815 3888 4861
rect 4066 4925 4112 4971
rect 4066 4815 4112 4861
rect 2959 1272 3005 1318
rect 2959 1144 3005 1190
rect 2959 1017 3005 1063
rect 2959 890 3005 936
rect 3183 1272 3229 1318
rect 3183 1144 3229 1190
rect 3183 1017 3229 1063
rect 3183 890 3229 936
rect 3407 1272 3453 1318
rect 3407 1144 3453 1190
rect 3407 1017 3453 1063
rect 3407 890 3453 936
rect 3631 1272 3677 1318
rect 3631 1144 3677 1190
rect 3631 1017 3677 1063
rect 3631 890 3677 936
rect 3855 1272 3901 1318
rect 3855 1144 3901 1190
rect 3855 1017 3901 1063
rect 3855 890 3901 936
rect 4079 1272 4125 1318
rect 4079 1144 4125 1190
rect 4079 1017 4125 1063
rect 4079 890 4125 936
rect 4303 1272 4349 1318
rect 4303 1144 4349 1190
rect 4303 1017 4349 1063
rect 4303 890 4349 936
<< psubdiff >>
rect 1835 7103 5034 7162
rect 1835 7057 1892 7103
rect 1938 7057 2072 7103
rect 2118 7057 2230 7103
rect 2276 7057 2388 7103
rect 2434 7057 2546 7103
rect 2592 7057 2704 7103
rect 2750 7057 2862 7103
rect 2908 7057 3021 7103
rect 3067 7057 3179 7103
rect 3225 7057 3337 7103
rect 3383 7057 3495 7103
rect 3541 7057 3653 7103
rect 3699 7057 3811 7103
rect 3857 7057 3970 7103
rect 4016 7057 4128 7103
rect 4174 7057 4286 7103
rect 4332 7057 4444 7103
rect 4490 7057 4602 7103
rect 4648 7057 4760 7103
rect 4806 7057 5034 7103
rect 1835 6997 5034 7057
rect 1835 6940 1995 6997
rect 1835 6894 1892 6940
rect 1938 6894 1995 6940
rect 1835 6777 1995 6894
rect 1835 6731 1892 6777
rect 1938 6731 1995 6777
rect 1835 6614 1995 6731
rect 1835 6568 1892 6614
rect 1938 6568 1995 6614
rect 1835 6450 1995 6568
rect 1835 6404 1892 6450
rect 1938 6404 1995 6450
rect 1835 6287 1995 6404
rect 1835 6241 1892 6287
rect 1938 6241 1995 6287
rect 1835 6124 1995 6241
rect 1835 6078 1892 6124
rect 1938 6078 1995 6124
rect 1835 5961 1995 6078
rect 1835 5915 1892 5961
rect 1938 5915 1995 5961
rect 1835 5797 1995 5915
rect 1835 5751 1892 5797
rect 1938 5751 1995 5797
rect 1835 5634 1995 5751
rect 1835 5588 1892 5634
rect 1938 5588 1995 5634
rect 1835 5471 1995 5588
rect 1835 5425 1892 5471
rect 1938 5425 1995 5471
rect 1835 5308 1995 5425
rect 1835 5262 1892 5308
rect 1938 5262 1995 5308
rect 1835 5145 1995 5262
rect 1835 5099 1892 5145
rect 1938 5099 1995 5145
rect 1835 4981 1995 5099
rect 1835 4935 1892 4981
rect 1938 4935 1995 4981
rect 1835 4818 1995 4935
rect 1835 4772 1892 4818
rect 1938 4772 1995 4818
rect 1835 4655 1995 4772
rect 1835 4609 1892 4655
rect 1938 4609 1995 4655
rect 1835 4491 1995 4609
rect 1835 4445 1892 4491
rect 1938 4445 1995 4491
rect 1835 4328 1995 4445
rect 1835 4282 1892 4328
rect 1938 4282 1995 4328
rect 1835 4165 1995 4282
rect 1835 4119 1892 4165
rect 1938 4119 1995 4165
rect 1835 4001 1995 4119
rect 1835 3955 1892 4001
rect 1938 3955 1995 4001
rect 1835 3838 1995 3955
rect 1835 3792 1892 3838
rect 1938 3792 1995 3838
rect 1835 3675 1995 3792
rect 1835 3629 1892 3675
rect 1938 3629 1995 3675
rect 1835 3512 1995 3629
rect 1835 3466 1892 3512
rect 1938 3466 1995 3512
rect 1835 3349 1995 3466
rect 1835 3303 1892 3349
rect 1938 3303 1995 3349
rect 1835 3185 1995 3303
rect 1835 3139 1892 3185
rect 1938 3139 1995 3185
rect 1835 3022 1995 3139
rect 1835 2976 1892 3022
rect 1938 2976 1995 3022
rect 1835 2859 1995 2976
rect 1835 2813 1892 2859
rect 1938 2813 1995 2859
rect 1835 2696 1995 2813
rect 1835 2650 1892 2696
rect 1938 2650 1995 2696
rect 1835 2532 1995 2650
rect 1835 2486 1892 2532
rect 1938 2486 1995 2532
rect 1835 2369 1995 2486
rect 1835 2323 1892 2369
rect 1938 2323 1995 2369
rect 1835 2206 1995 2323
rect 1835 2160 1892 2206
rect 1938 2160 1995 2206
rect 1835 2102 1995 2160
rect 1835 2043 2627 2102
rect 1835 1997 1892 2043
rect 1938 1997 2050 2043
rect 2096 1997 2208 2043
rect 2254 1997 2366 2043
rect 2412 1997 2524 2043
rect 2570 1997 2627 2043
rect 1835 1937 2627 1997
rect 2468 1789 2627 1937
rect 2468 1743 2524 1789
rect 2570 1743 2627 1789
rect 2468 1626 2627 1743
rect 2468 1580 2524 1626
rect 2570 1580 2627 1626
rect 2468 1462 2627 1580
rect 2468 1416 2524 1462
rect 2570 1416 2627 1462
rect 2468 1299 2627 1416
rect 2468 1253 2524 1299
rect 2570 1253 2627 1299
rect 2468 1136 2627 1253
rect 2468 1090 2524 1136
rect 2570 1090 2627 1136
rect 2468 972 2627 1090
rect 2468 926 2524 972
rect 2570 926 2627 972
rect 2468 809 2627 926
rect 4875 1055 5034 6997
rect 4875 1009 4932 1055
rect 4978 1009 5034 1055
rect 4875 892 5034 1009
rect 2468 763 2524 809
rect 2570 763 2627 809
rect 4875 846 4932 892
rect 4978 846 5034 892
rect 2468 646 2627 763
rect 4875 728 5034 846
rect 4875 682 4932 728
rect 4978 682 5034 728
rect 2468 600 2524 646
rect 2570 600 2627 646
rect 2468 482 2627 600
rect 4875 565 5034 682
rect 2468 436 2524 482
rect 2570 436 2627 482
rect 2468 319 2627 436
rect 2468 273 2524 319
rect 2570 273 2627 319
rect 2468 235 2627 273
rect 4875 519 4932 565
rect 4978 519 5034 565
rect 4875 402 5034 519
rect 4875 356 4932 402
rect 4978 356 5034 402
rect 2468 234 2628 235
rect 4875 234 5034 356
rect 2468 175 5034 234
rect 2468 129 2781 175
rect 2827 129 2939 175
rect 2985 129 3097 175
rect 3143 129 3256 175
rect 3302 129 3414 175
rect 3460 129 3572 175
rect 3618 129 3730 175
rect 3776 129 3888 175
rect 3934 129 4046 175
rect 4092 129 4205 175
rect 4251 129 4363 175
rect 4409 129 4521 175
rect 4567 129 5034 175
rect 2468 69 5034 129
<< nsubdiff >>
rect 2245 4911 2400 4968
rect 2245 4865 2299 4911
rect 2345 4865 2400 4911
rect 2245 4808 2400 4865
rect 4398 4911 4553 4968
rect 4398 4865 4452 4911
rect 4498 4865 4553 4911
rect 4398 4808 4553 4865
rect 2957 624 4377 681
rect 2957 578 3011 624
rect 3057 578 3170 624
rect 3216 578 3328 624
rect 3374 578 3486 624
rect 3532 578 3644 624
rect 3690 578 3802 624
rect 3848 578 3960 624
rect 4006 578 4118 624
rect 4164 578 4277 624
rect 4323 578 4377 624
rect 2957 521 4377 578
<< psubdiffcont >>
rect 1892 7057 1938 7103
rect 2072 7057 2118 7103
rect 2230 7057 2276 7103
rect 2388 7057 2434 7103
rect 2546 7057 2592 7103
rect 2704 7057 2750 7103
rect 2862 7057 2908 7103
rect 3021 7057 3067 7103
rect 3179 7057 3225 7103
rect 3337 7057 3383 7103
rect 3495 7057 3541 7103
rect 3653 7057 3699 7103
rect 3811 7057 3857 7103
rect 3970 7057 4016 7103
rect 4128 7057 4174 7103
rect 4286 7057 4332 7103
rect 4444 7057 4490 7103
rect 4602 7057 4648 7103
rect 4760 7057 4806 7103
rect 1892 6894 1938 6940
rect 1892 6731 1938 6777
rect 1892 6568 1938 6614
rect 1892 6404 1938 6450
rect 1892 6241 1938 6287
rect 1892 6078 1938 6124
rect 1892 5915 1938 5961
rect 1892 5751 1938 5797
rect 1892 5588 1938 5634
rect 1892 5425 1938 5471
rect 1892 5262 1938 5308
rect 1892 5099 1938 5145
rect 1892 4935 1938 4981
rect 1892 4772 1938 4818
rect 1892 4609 1938 4655
rect 1892 4445 1938 4491
rect 1892 4282 1938 4328
rect 1892 4119 1938 4165
rect 1892 3955 1938 4001
rect 1892 3792 1938 3838
rect 1892 3629 1938 3675
rect 1892 3466 1938 3512
rect 1892 3303 1938 3349
rect 1892 3139 1938 3185
rect 1892 2976 1938 3022
rect 1892 2813 1938 2859
rect 1892 2650 1938 2696
rect 1892 2486 1938 2532
rect 1892 2323 1938 2369
rect 1892 2160 1938 2206
rect 1892 1997 1938 2043
rect 2050 1997 2096 2043
rect 2208 1997 2254 2043
rect 2366 1997 2412 2043
rect 2524 1997 2570 2043
rect 2524 1743 2570 1789
rect 2524 1580 2570 1626
rect 2524 1416 2570 1462
rect 2524 1253 2570 1299
rect 2524 1090 2570 1136
rect 2524 926 2570 972
rect 4932 1009 4978 1055
rect 2524 763 2570 809
rect 4932 846 4978 892
rect 4932 682 4978 728
rect 2524 600 2570 646
rect 2524 436 2570 482
rect 2524 273 2570 319
rect 4932 519 4978 565
rect 4932 356 4978 402
rect 2781 129 2827 175
rect 2939 129 2985 175
rect 3097 129 3143 175
rect 3256 129 3302 175
rect 3414 129 3460 175
rect 3572 129 3618 175
rect 3730 129 3776 175
rect 3888 129 3934 175
rect 4046 129 4092 175
rect 4205 129 4251 175
rect 4363 129 4409 175
rect 4521 129 4567 175
<< nsubdiffcont >>
rect 2299 4865 2345 4911
rect 4452 4865 4498 4911
rect 3011 578 3057 624
rect 3170 578 3216 624
rect 3328 578 3374 624
rect 3486 578 3532 624
rect 3644 578 3690 624
rect 3802 578 3848 624
rect 3960 578 4006 624
rect 4118 578 4164 624
rect 4277 578 4323 624
<< polysilicon >>
rect 3151 6740 3719 6759
rect 3151 6694 3412 6740
rect 3458 6694 3719 6740
rect 3151 6659 3719 6694
rect 2464 6586 2584 6659
rect 2688 6586 2808 6659
rect 3151 6586 3271 6659
rect 3375 6586 3495 6659
rect 3599 6586 3719 6659
rect 4049 6586 4169 6659
rect 4273 6586 4393 6659
rect 2464 5720 2584 6132
rect 2688 5720 2808 6132
rect 3151 6059 3271 6132
rect 3375 6059 3495 6132
rect 3599 6059 3719 6132
rect 3375 5793 3494 6059
rect 3375 5720 3495 5793
rect 4049 5720 4169 6132
rect 4273 5720 4393 6132
rect 2095 5216 2179 5235
rect 2095 5170 2114 5216
rect 2160 5206 2179 5216
rect 2464 5206 2584 5266
rect 2688 5206 2808 5266
rect 2160 5170 2808 5206
rect 3375 5193 3495 5266
rect 4049 5206 4169 5266
rect 4273 5206 4393 5266
rect 4635 5216 4719 5235
rect 4635 5206 4654 5216
rect 2095 5151 2808 5170
rect 4049 5170 4654 5206
rect 4700 5170 4719 5216
rect 4049 5151 4719 5170
rect 2797 4984 2917 5056
rect 3021 4984 3141 5056
rect 3245 4984 3365 5056
rect 3469 4984 3589 5056
rect 3693 4984 3813 5056
rect 3917 4984 4037 5056
rect 2797 4740 2917 4802
rect 2699 4721 2917 4740
rect 2699 4675 2718 4721
rect 2764 4675 2917 4721
rect 2699 4656 2917 4675
rect 3021 4621 3141 4802
rect 2556 4507 2760 4526
rect 2556 4461 2695 4507
rect 2741 4461 2760 4507
rect 2556 4442 2760 4461
rect 2332 3999 2452 4070
rect 2556 3999 2676 4442
rect 3021 4310 3124 4621
rect 3245 4507 3365 4802
rect 3469 4728 3589 4802
rect 3693 4758 3813 4802
rect 3245 4461 3264 4507
rect 3310 4461 3365 4507
rect 3021 4291 3159 4310
rect 3021 4267 3094 4291
rect 2780 4245 3094 4267
rect 3140 4245 3159 4291
rect 2780 4226 3159 4245
rect 2780 4197 3124 4226
rect 2780 3999 2900 4197
rect 3004 3999 3124 4197
rect 3245 4105 3365 4461
rect 3487 4619 3589 4728
rect 3720 4623 3813 4758
rect 3917 4742 4037 4802
rect 3917 4723 4121 4742
rect 3917 4677 4056 4723
rect 4102 4677 4121 4723
rect 3917 4658 4121 4677
rect 3487 4507 3615 4619
rect 3487 4461 3550 4507
rect 3596 4461 3615 4507
rect 3487 4108 3615 4461
rect 3720 4291 3848 4623
rect 3720 4245 3739 4291
rect 3785 4267 3848 4291
rect 4124 4507 4244 4526
rect 4124 4461 4143 4507
rect 4189 4461 4244 4507
rect 3785 4245 4020 4267
rect 3720 4197 4020 4245
rect 3245 4071 3348 4105
rect 3487 4071 3572 4108
rect 3720 4101 3848 4197
rect 3720 4071 3796 4101
rect 3228 3999 3348 4071
rect 3452 3999 3572 4071
rect 3676 3999 3796 4071
rect 3900 3999 4020 4197
rect 4124 3999 4244 4461
rect 4348 3999 4468 4070
rect 2332 3253 2452 3317
rect 2257 3243 2452 3253
rect 2556 3243 2676 3317
rect 2780 3243 2900 3317
rect 3004 3243 3124 3317
rect 3228 3243 3348 3317
rect 3452 3243 3572 3317
rect 3676 3243 3796 3317
rect 3900 3243 4020 3317
rect 4124 3243 4244 3317
rect 4348 3253 4468 3317
rect 4348 3243 4611 3253
rect 2257 3208 2450 3243
rect 2257 3162 2331 3208
rect 2377 3162 2450 3208
rect 2257 3116 2450 3162
rect 4418 3208 4611 3243
rect 4418 3162 4492 3208
rect 4538 3162 4611 3208
rect 2589 3078 2709 3150
rect 2813 3078 2933 3150
rect 3037 3078 3157 3150
rect 3261 3078 3381 3150
rect 3485 3078 3605 3150
rect 3709 3078 3829 3150
rect 3933 3078 4053 3150
rect 4157 3078 4277 3150
rect 4418 3116 4611 3162
rect 2589 2447 2709 2510
rect 2813 2447 2933 2510
rect 3037 2447 3157 2510
rect 3261 2447 3381 2510
rect 3485 2447 3605 2510
rect 3709 2447 3829 2510
rect 3933 2447 4053 2510
rect 4157 2447 4277 2510
rect 2589 2401 4277 2447
rect 2589 2355 2663 2401
rect 2709 2355 2966 2401
rect 3012 2355 3412 2401
rect 3458 2355 3864 2401
rect 3910 2355 4156 2401
rect 4202 2355 4277 2401
rect 2589 2309 4277 2355
rect 3034 2156 3154 2229
rect 3482 2156 3602 2229
rect 3706 2156 3826 2229
rect 3930 2156 4050 2229
rect 4154 2156 4274 2229
rect 3034 1595 3154 1702
rect 3034 1593 3378 1595
rect 2870 1574 3378 1593
rect 2870 1528 2889 1574
rect 3029 1534 3378 1574
rect 3029 1528 3154 1534
rect 2870 1509 3154 1528
rect 3034 1331 3154 1509
rect 3258 1331 3378 1534
rect 3482 1593 3602 1702
rect 3706 1642 3826 1702
rect 3930 1642 4050 1702
rect 3706 1593 4050 1642
rect 3482 1588 4050 1593
rect 3482 1574 3826 1588
rect 3482 1528 3549 1574
rect 3689 1528 3826 1574
rect 3482 1509 3826 1528
rect 3482 1331 3602 1509
rect 3706 1331 3826 1509
rect 4154 1581 4274 1702
rect 4154 1562 4449 1581
rect 4154 1516 4290 1562
rect 4430 1516 4449 1562
rect 4154 1497 4449 1516
rect 4154 1452 4274 1497
rect 3930 1391 4274 1452
rect 3930 1331 4050 1391
rect 4154 1331 4274 1391
rect 3034 804 3154 877
rect 3258 804 3378 877
rect 3482 804 3602 877
rect 3706 804 3826 877
rect 3930 804 4050 877
rect 4154 804 4274 877
<< polycontact >>
rect 3412 6694 3458 6740
rect 2114 5170 2160 5216
rect 4654 5170 4700 5216
rect 2718 4675 2764 4721
rect 2695 4461 2741 4507
rect 3264 4461 3310 4507
rect 3094 4245 3140 4291
rect 4056 4677 4102 4723
rect 3550 4461 3596 4507
rect 3739 4245 3785 4291
rect 4143 4461 4189 4507
rect 2331 3162 2377 3208
rect 4492 3162 4538 3208
rect 2663 2355 2709 2401
rect 2966 2355 3012 2401
rect 3412 2355 3458 2401
rect 3864 2355 3910 2401
rect 4156 2355 4202 2401
rect 2889 1528 3029 1574
rect 3549 1528 3689 1574
rect 4290 1516 4430 1562
<< metal1 >>
rect 1756 8029 2524 8033
rect 3076 8029 4501 8033
rect 1756 8009 2633 8029
rect 1756 7957 2355 8009
rect 2407 7957 2541 8009
rect 2593 7957 2633 8009
rect 1756 7937 2633 7957
rect 2951 8009 4501 8029
rect 2951 7957 2981 8009
rect 3033 7957 3167 8009
rect 3219 7957 4219 8009
rect 4271 7957 4405 8009
rect 4457 7957 4501 8009
rect 2951 7937 4501 7957
rect 1756 7936 2524 7937
rect 3076 7936 4501 7937
rect 2430 7824 2524 7936
rect 2430 7800 4501 7824
rect 2430 7748 2737 7800
rect 2789 7748 2923 7800
rect 2975 7748 3541 7800
rect 3593 7748 3727 7800
rect 3779 7748 4501 7800
rect 2430 7727 4501 7748
rect 1756 7478 4885 7616
rect 1251 7339 4501 7362
rect 1251 7287 3410 7339
rect 3462 7287 4501 7339
rect 1251 7265 4501 7287
rect 1844 7103 5025 7153
rect 1844 7057 1892 7103
rect 1938 7057 2072 7103
rect 2118 7057 2230 7103
rect 2276 7057 2388 7103
rect 2434 7057 2546 7103
rect 2592 7057 2704 7103
rect 2750 7057 2862 7103
rect 2908 7057 3021 7103
rect 3067 7057 3179 7103
rect 3225 7057 3337 7103
rect 3383 7057 3495 7103
rect 3541 7057 3653 7103
rect 3699 7057 3811 7103
rect 3857 7057 3970 7103
rect 4016 7057 4128 7103
rect 4174 7057 4286 7103
rect 4332 7057 4444 7103
rect 4490 7057 4602 7103
rect 4648 7057 4760 7103
rect 4806 7057 5025 7103
rect 1844 7006 5025 7057
rect 1844 6940 1986 7006
rect 1844 6894 1892 6940
rect 1938 6894 1986 6940
rect 1844 6777 1986 6894
rect 3271 6823 3609 6899
rect 3387 6822 3482 6823
rect 1844 6731 1892 6777
rect 1938 6731 1986 6777
rect 2797 6741 2925 6763
rect 3388 6750 3482 6822
rect 1844 6614 1986 6731
rect 1844 6568 1892 6614
rect 1938 6568 1986 6614
rect 2387 6740 3310 6741
rect 2387 6688 2835 6740
rect 2887 6688 3310 6740
rect 2387 6666 3310 6688
rect 2387 6577 2458 6666
rect 1844 6450 1986 6568
rect 1844 6404 1892 6450
rect 1938 6404 1986 6450
rect 1844 6287 1986 6404
rect 1844 6241 1892 6287
rect 1938 6241 1986 6287
rect 1844 6124 1986 6241
rect 2386 6573 2458 6577
rect 2386 6527 2389 6573
rect 2435 6527 2458 6573
rect 2386 6446 2458 6527
rect 2613 6573 2659 6586
rect 2613 6464 2659 6527
rect 2837 6573 2883 6666
rect 3239 6586 3310 6666
rect 3388 6698 3408 6750
rect 3460 6698 3482 6750
rect 3388 6694 3412 6698
rect 3458 6694 3482 6698
rect 3388 6657 3482 6694
rect 3559 6718 4483 6741
rect 3559 6666 3970 6718
rect 4022 6666 4483 6718
rect 3559 6586 3631 6666
rect 3932 6644 4060 6666
rect 3076 6573 3122 6586
rect 2386 6400 2389 6446
rect 2435 6400 2458 6446
rect 2386 6319 2458 6400
rect 2386 6273 2389 6319
rect 2435 6273 2458 6319
rect 2386 6191 2458 6273
rect 2386 6145 2389 6191
rect 2435 6145 2458 6191
rect 2596 6446 2688 6464
rect 2596 6400 2613 6446
rect 2659 6424 2688 6446
rect 2596 6372 2616 6400
rect 2668 6372 2688 6424
rect 2596 6319 2688 6372
rect 2596 6273 2613 6319
rect 2659 6273 2688 6319
rect 2596 6238 2688 6273
rect 2596 6191 2616 6238
rect 2596 6145 2613 6191
rect 2668 6186 2688 6238
rect 2659 6145 2688 6186
rect 2837 6446 2883 6527
rect 2837 6319 2883 6400
rect 2837 6191 2883 6273
rect 3050 6527 3076 6533
rect 3239 6573 3346 6586
rect 3122 6527 3142 6533
rect 3050 6503 3142 6527
rect 3050 6451 3070 6503
rect 3122 6451 3142 6503
rect 3050 6446 3142 6451
rect 3050 6400 3076 6446
rect 3122 6400 3142 6446
rect 3050 6319 3142 6400
rect 3050 6317 3076 6319
rect 3050 6265 3070 6317
rect 3122 6265 3142 6319
rect 3050 6225 3142 6265
rect 3239 6527 3300 6573
rect 3239 6464 3346 6527
rect 3524 6573 3631 6586
rect 3570 6527 3631 6573
rect 3748 6573 3794 6586
rect 3524 6464 3631 6527
rect 3239 6446 3369 6464
rect 3239 6424 3300 6446
rect 3346 6424 3369 6446
rect 3239 6372 3297 6424
rect 3349 6372 3369 6424
rect 3239 6319 3369 6372
rect 3239 6273 3300 6319
rect 3346 6273 3369 6319
rect 3239 6238 3369 6273
rect 2386 6132 2458 6145
rect 2613 6132 2659 6145
rect 2837 6132 2883 6145
rect 3076 6191 3122 6225
rect 3076 6132 3122 6145
rect 3239 6186 3297 6238
rect 3349 6186 3369 6238
rect 3239 6145 3300 6186
rect 3346 6145 3369 6186
rect 3503 6446 3631 6464
rect 3503 6424 3524 6446
rect 3570 6424 3631 6446
rect 3503 6372 3523 6424
rect 3575 6372 3631 6424
rect 3503 6319 3631 6372
rect 3503 6273 3524 6319
rect 3570 6273 3631 6319
rect 3503 6238 3631 6273
rect 3503 6186 3523 6238
rect 3575 6186 3631 6238
rect 3722 6527 3748 6533
rect 3939 6573 4055 6644
rect 3794 6527 3814 6533
rect 3722 6503 3814 6527
rect 3722 6451 3742 6503
rect 3794 6451 3814 6503
rect 3722 6446 3814 6451
rect 3722 6400 3748 6446
rect 3794 6400 3814 6446
rect 3722 6319 3814 6400
rect 3722 6317 3748 6319
rect 3722 6265 3742 6317
rect 3794 6265 3814 6319
rect 3722 6225 3814 6265
rect 3939 6527 3974 6573
rect 4020 6527 4055 6573
rect 3939 6446 4055 6527
rect 4198 6573 4244 6586
rect 4198 6464 4244 6527
rect 4411 6573 4483 6666
rect 4411 6527 4422 6573
rect 4468 6527 4483 6573
rect 3939 6400 3974 6446
rect 4020 6400 4055 6446
rect 3939 6319 4055 6400
rect 3939 6273 3974 6319
rect 4020 6273 4055 6319
rect 3503 6145 3524 6186
rect 3570 6145 3631 6186
rect 3239 6140 3346 6145
rect 3300 6132 3346 6140
rect 3524 6140 3631 6145
rect 3748 6191 3794 6225
rect 3524 6132 3570 6140
rect 3748 6132 3794 6145
rect 3939 6191 4055 6273
rect 3939 6145 3974 6191
rect 4020 6145 4055 6191
rect 4181 6446 4273 6464
rect 4181 6400 4198 6446
rect 4244 6424 4273 6446
rect 4181 6372 4201 6400
rect 4253 6372 4273 6424
rect 4181 6319 4273 6372
rect 4181 6273 4198 6319
rect 4244 6273 4273 6319
rect 4181 6238 4273 6273
rect 4181 6191 4201 6238
rect 4181 6145 4198 6191
rect 4253 6186 4273 6238
rect 4244 6145 4273 6186
rect 4411 6446 4483 6527
rect 4411 6400 4422 6446
rect 4468 6400 4483 6446
rect 4411 6319 4483 6400
rect 4411 6273 4422 6319
rect 4468 6273 4483 6319
rect 4411 6191 4483 6273
rect 4411 6145 4422 6191
rect 4468 6145 4483 6191
rect 3939 6140 4055 6145
rect 3974 6132 4020 6140
rect 4198 6132 4244 6145
rect 4411 6140 4483 6145
rect 4422 6132 4468 6140
rect 1844 6078 1892 6124
rect 1938 6078 1986 6124
rect 1844 5961 1986 6078
rect 1844 5915 1892 5961
rect 1938 5915 1986 5961
rect 1844 5797 1986 5915
rect 1844 5751 1892 5797
rect 1938 5751 1986 5797
rect 1844 5634 1986 5751
rect 2378 5884 2467 6061
rect 2843 5884 2933 6061
rect 3278 6057 4468 6061
rect 3276 6036 4468 6057
rect 3276 5984 3316 6036
rect 3368 5984 4468 6036
rect 3276 5968 4468 5984
rect 3276 5964 3404 5968
rect 3467 5884 3595 5885
rect 2378 5864 3595 5884
rect 2378 5812 3503 5864
rect 3555 5812 3595 5864
rect 2378 5792 3595 5812
rect 2378 5791 3591 5792
rect 2378 5711 2467 5791
rect 1844 5588 1892 5634
rect 1938 5588 1986 5634
rect 1844 5471 1986 5588
rect 1844 5425 1892 5471
rect 1938 5425 1986 5471
rect 1844 5308 1986 5425
rect 1844 5262 1892 5308
rect 1938 5262 1986 5308
rect 2377 5707 2467 5711
rect 2377 5661 2389 5707
rect 2435 5661 2467 5707
rect 2377 5580 2467 5661
rect 2377 5534 2389 5580
rect 2435 5534 2467 5580
rect 2377 5453 2467 5534
rect 2377 5407 2389 5453
rect 2435 5407 2467 5453
rect 2377 5325 2467 5407
rect 2377 5304 2389 5325
rect 2435 5304 2467 5325
rect 2613 5707 2659 5720
rect 2613 5580 2659 5661
rect 2613 5453 2659 5534
rect 2613 5325 2659 5407
rect 2389 5266 2435 5279
rect 1844 5145 1986 5262
rect 1844 5099 1892 5145
rect 1938 5099 1986 5145
rect 1844 4981 1986 5099
rect 1844 4935 1892 4981
rect 1938 4935 1986 4981
rect 1844 4818 1986 4935
rect 1844 4772 1892 4818
rect 1938 4772 1986 4818
rect 1844 4655 1986 4772
rect 1844 4609 1892 4655
rect 1938 4609 1986 4655
rect 1844 4491 1986 4609
rect 1844 4445 1892 4491
rect 1938 4445 1986 4491
rect 1844 4328 1986 4445
rect 1844 4282 1892 4328
rect 1938 4282 1986 4328
rect 1844 4165 1986 4282
rect 1844 4119 1892 4165
rect 1938 4119 1986 4165
rect 1844 4001 1986 4119
rect 1844 3955 1892 4001
rect 1938 3955 1986 4001
rect 1844 3838 1986 3955
rect 1844 3792 1892 3838
rect 1938 3792 1986 3838
rect 1844 3675 1986 3792
rect 1844 3629 1892 3675
rect 1938 3629 1986 3675
rect 1844 3512 1986 3629
rect 1844 3466 1892 3512
rect 1938 3466 1986 3512
rect 1844 3349 1986 3466
rect 1844 3303 1892 3349
rect 1938 3303 1986 3349
rect 1844 3185 1986 3303
rect 1844 3139 1892 3185
rect 1938 3139 1986 3185
rect 1844 3022 1986 3139
rect 1844 2976 1892 3022
rect 1938 2976 1986 3022
rect 1844 2859 1986 2976
rect 1844 2813 1892 2859
rect 1938 2813 1986 2859
rect 1844 2696 1986 2813
rect 1844 2650 1892 2696
rect 1938 2650 1986 2696
rect 1844 2532 1986 2650
rect 1844 2486 1892 2532
rect 1938 2486 1986 2532
rect 1844 2369 1986 2486
rect 1844 2323 1892 2369
rect 1938 2323 1986 2369
rect 1844 2206 1986 2323
rect 2064 5216 2171 5227
rect 2064 5170 2114 5216
rect 2160 5170 2171 5216
rect 2613 5195 2659 5279
rect 2837 5707 2883 5791
rect 2837 5580 2883 5661
rect 2837 5453 2883 5534
rect 2837 5325 2883 5407
rect 2837 5266 2883 5279
rect 3300 5707 3346 5720
rect 3300 5580 3346 5661
rect 3300 5453 3346 5534
rect 3300 5325 3346 5407
rect 3300 5195 3346 5279
rect 2064 5159 2171 5170
rect 2064 2438 2136 5159
rect 2448 5120 3346 5195
rect 3524 5707 3570 5720
rect 3524 5580 3570 5661
rect 3524 5453 3570 5534
rect 3524 5325 3570 5407
rect 3524 5195 3570 5279
rect 3974 5707 4020 5968
rect 3974 5580 4020 5661
rect 3974 5453 4020 5534
rect 3974 5325 4020 5407
rect 3974 5266 4020 5279
rect 4198 5707 4244 5720
rect 4198 5580 4244 5661
rect 4198 5453 4244 5534
rect 4198 5325 4244 5407
rect 4198 5195 4244 5279
rect 4422 5707 4468 5968
rect 4422 5580 4468 5661
rect 4422 5453 4468 5534
rect 4422 5325 4468 5407
rect 4422 5266 4468 5279
rect 4643 5216 4916 5227
rect 3524 5120 4340 5195
rect 4643 5170 4654 5216
rect 4700 5170 4916 5216
rect 4643 5159 4916 5170
rect 2287 5025 2379 5030
rect 2286 5024 2380 5025
rect 2264 5000 2380 5024
rect 2264 4948 2307 5000
rect 2359 4948 2380 5000
rect 2264 4911 2380 4948
rect 2264 4865 2299 4911
rect 2345 4865 2380 4911
rect 2264 4814 2380 4865
rect 2264 4762 2307 4814
rect 2359 4762 2380 4814
rect 2264 4719 2380 4762
rect 2448 4319 2520 5120
rect 3151 5025 3243 5030
rect 3623 5025 3715 5030
rect 3151 5024 3245 5025
rect 3623 5024 3717 5025
rect 3144 5000 3260 5024
rect 2722 4975 2768 4984
rect 2679 4971 2794 4975
rect 2679 4943 2722 4971
rect 2768 4943 2794 4971
rect 2679 4891 2721 4943
rect 2773 4891 2794 4943
rect 2679 4861 2794 4891
rect 2679 4815 2722 4861
rect 2768 4815 2794 4861
rect 2679 4757 2794 4815
rect 2679 4721 2721 4757
rect 2679 4675 2718 4721
rect 2773 4705 2794 4757
rect 2764 4675 2794 4705
rect 2679 4664 2794 4675
rect 2911 4971 2992 4984
rect 2911 4925 2946 4971
rect 2911 4861 2992 4925
rect 2911 4815 2946 4861
rect 2911 4802 2992 4815
rect 3144 4971 3171 5000
rect 3144 4925 3170 4971
rect 3223 4948 3260 5000
rect 3610 5000 3725 5024
rect 3216 4925 3260 4948
rect 3144 4861 3260 4925
rect 3144 4815 3170 4861
rect 3216 4815 3260 4861
rect 3144 4814 3260 4815
rect 2911 4532 2975 4802
rect 3144 4762 3171 4814
rect 3223 4762 3260 4814
rect 3394 4975 3440 4984
rect 3394 4971 3471 4975
rect 3440 4925 3471 4971
rect 3394 4861 3471 4925
rect 3440 4815 3471 4861
rect 3394 4802 3471 4815
rect 3144 4719 3260 4762
rect 2684 4510 2992 4532
rect 2684 4507 2722 4510
rect 2684 4461 2695 4507
rect 2684 4458 2722 4461
rect 2774 4458 2902 4510
rect 2954 4458 2992 4510
rect 2684 4436 2992 4458
rect 3083 4510 3329 4544
rect 3083 4458 3231 4510
rect 3283 4507 3329 4510
rect 3310 4461 3329 4507
rect 3283 4458 3329 4461
rect 2332 4298 2520 4319
rect 2332 4246 2428 4298
rect 2480 4246 2520 4298
rect 2332 4226 2520 4246
rect 2332 4145 2403 4226
rect 2332 4071 2518 4145
rect 2446 3999 2518 4071
rect 2257 3988 2303 3999
rect 2213 3986 2329 3988
rect 2213 3330 2257 3986
rect 2303 3330 2329 3986
rect 2446 3986 2527 3999
rect 2446 3910 2481 3986
rect 2213 3244 2329 3330
rect 2705 3986 2751 3999
rect 2481 3317 2527 3330
rect 2679 3330 2705 3411
rect 2911 3986 2975 4436
rect 3083 4424 3329 4458
rect 3083 4299 3293 4326
rect 3399 4322 3471 4802
rect 3610 4971 3643 5000
rect 3610 4925 3618 4971
rect 3695 4948 3725 5000
rect 3664 4925 3725 4948
rect 3610 4861 3725 4925
rect 3610 4815 3618 4861
rect 3664 4815 3725 4861
rect 3610 4814 3725 4815
rect 3610 4762 3643 4814
rect 3695 4762 3725 4814
rect 3842 4973 3888 4984
rect 3842 4971 3958 4973
rect 3888 4925 3958 4971
rect 3842 4861 3958 4925
rect 3888 4815 3958 4861
rect 3842 4802 3958 4815
rect 3610 4719 3725 4762
rect 3539 4510 3758 4544
rect 3886 4532 3958 4802
rect 4039 4971 4155 4984
rect 4039 4943 4066 4971
rect 4039 4891 4060 4943
rect 4112 4891 4155 4971
rect 4039 4861 4155 4891
rect 4039 4815 4066 4861
rect 4112 4815 4155 4861
rect 4039 4757 4155 4815
rect 4039 4723 4060 4757
rect 4039 4677 4056 4723
rect 4112 4705 4155 4757
rect 4102 4677 4155 4705
rect 4039 4664 4155 4677
rect 3539 4507 3587 4510
rect 3539 4461 3550 4507
rect 3539 4458 3587 4461
rect 3639 4458 3758 4510
rect 3539 4424 3758 4458
rect 3883 4510 4200 4532
rect 3883 4458 3921 4510
rect 3973 4458 4101 4510
rect 4153 4507 4200 4510
rect 4189 4461 4200 4507
rect 4153 4458 4200 4461
rect 3883 4436 4200 4458
rect 4268 4530 4340 5120
rect 4418 5025 4510 5030
rect 4418 5024 4512 5025
rect 4418 5000 4534 5024
rect 4418 4948 4438 5000
rect 4490 4948 4534 5000
rect 4418 4911 4534 4948
rect 4418 4865 4452 4911
rect 4498 4865 4534 4911
rect 4418 4814 4534 4865
rect 4418 4762 4438 4814
rect 4490 4762 4534 4814
rect 4418 4719 4534 4762
rect 4268 4509 4396 4530
rect 4268 4457 4304 4509
rect 4356 4457 4396 4509
rect 4268 4437 4396 4457
rect 3083 4291 3121 4299
rect 3083 4245 3094 4291
rect 3173 4247 3293 4299
rect 3140 4245 3293 4247
rect 3083 4202 3293 4245
rect 3371 4299 3499 4322
rect 3371 4247 3409 4299
rect 3461 4247 3499 4299
rect 3371 4225 3499 4247
rect 3577 4299 3796 4326
rect 3577 4247 3697 4299
rect 3749 4291 3796 4299
rect 3577 4245 3739 4247
rect 3785 4245 3796 4291
rect 3399 3999 3471 4225
rect 3577 4202 3796 4245
rect 3886 3999 3958 4436
rect 4268 4227 4340 4437
rect 4475 4322 4547 4533
rect 4474 4319 4547 4322
rect 4440 4298 4568 4319
rect 4440 4246 4476 4298
rect 4528 4246 4568 4298
rect 4440 4226 4568 4246
rect 4474 4225 4547 4226
rect 4475 4145 4547 4225
rect 4273 4071 4547 4145
rect 2911 3891 2929 3986
rect 2751 3330 2794 3411
rect 2679 3245 2794 3330
rect 3153 3986 3199 3999
rect 2929 3317 2975 3330
rect 3144 3330 3153 3411
rect 3377 3986 3471 3999
rect 3199 3330 3260 3411
rect 3144 3245 3260 3330
rect 3423 3855 3471 3986
rect 3601 3986 3647 3999
rect 3377 3317 3423 3330
rect 3825 3986 3958 3999
rect 3647 3330 3725 3411
rect 3601 3317 3725 3330
rect 3871 3891 3958 3986
rect 4049 3986 4095 3999
rect 3825 3317 3871 3330
rect 3610 3245 3725 3317
rect 4049 3245 4095 3330
rect 4273 3986 4319 4071
rect 4273 3317 4319 3330
rect 4497 3988 4543 3999
rect 4497 3986 4657 3988
rect 4543 3330 4657 3986
rect 4497 3317 4657 3330
rect 4541 3245 4657 3317
rect 2213 3242 2411 3244
rect 2213 3221 2486 3242
rect 2213 3208 2394 3221
rect 2213 3162 2331 3208
rect 2377 3169 2394 3208
rect 2446 3169 2486 3221
rect 2377 3162 2486 3169
rect 2213 3149 2486 3162
rect 2679 3152 4095 3245
rect 4540 3244 4657 3245
rect 4457 3242 4657 3244
rect 4378 3221 4657 3242
rect 4378 3169 4414 3221
rect 4466 3208 4657 3221
rect 4466 3169 4492 3208
rect 4378 3162 4492 3169
rect 4538 3162 4657 3208
rect 2213 3125 2411 3149
rect 2514 3065 2560 3078
rect 2514 2941 2560 3019
rect 2501 2895 2514 2929
rect 2703 3065 2818 3152
rect 2703 3019 2738 3065
rect 2784 3019 2818 3065
rect 2703 2941 2818 3019
rect 2560 2899 2593 2929
rect 2501 2847 2521 2895
rect 2573 2847 2593 2899
rect 2501 2817 2593 2847
rect 2501 2771 2514 2817
rect 2560 2771 2593 2817
rect 2501 2713 2593 2771
rect 2501 2693 2521 2713
rect 2501 2647 2514 2693
rect 2573 2661 2593 2713
rect 2560 2647 2593 2661
rect 2501 2621 2593 2647
rect 2703 2895 2738 2941
rect 2784 2895 2818 2941
rect 2962 3065 3008 3078
rect 2962 2941 3008 3019
rect 2703 2817 2818 2895
rect 2703 2771 2738 2817
rect 2784 2771 2818 2817
rect 2703 2693 2818 2771
rect 2703 2647 2738 2693
rect 2784 2647 2818 2693
rect 2514 2569 2560 2621
rect 2514 2510 2560 2523
rect 2703 2569 2818 2647
rect 2938 2899 2962 2929
rect 3151 3065 3266 3152
rect 3151 3019 3186 3065
rect 3232 3019 3266 3065
rect 3151 2941 3266 3019
rect 3008 2899 3030 2929
rect 2938 2847 2958 2899
rect 3010 2847 3030 2899
rect 2938 2817 3030 2847
rect 2938 2771 2962 2817
rect 3008 2771 3030 2817
rect 2938 2713 3030 2771
rect 2938 2661 2958 2713
rect 3010 2661 3030 2713
rect 2938 2647 2962 2661
rect 3008 2647 3030 2661
rect 2938 2621 3030 2647
rect 3151 2895 3186 2941
rect 3232 2895 3266 2941
rect 3410 3065 3456 3078
rect 3410 2941 3456 3019
rect 3151 2817 3266 2895
rect 3151 2771 3186 2817
rect 3232 2771 3266 2817
rect 3151 2693 3266 2771
rect 3151 2647 3186 2693
rect 3232 2647 3266 2693
rect 2703 2523 2738 2569
rect 2784 2523 2818 2569
rect 2703 2518 2818 2523
rect 2962 2569 3008 2621
rect 2738 2510 2784 2518
rect 2962 2510 3008 2523
rect 3151 2569 3266 2647
rect 3386 2899 3410 2929
rect 3599 3065 3714 3152
rect 3599 3019 3634 3065
rect 3680 3019 3714 3065
rect 3599 2941 3714 3019
rect 3456 2899 3478 2929
rect 3386 2847 3406 2899
rect 3458 2847 3478 2899
rect 3386 2817 3478 2847
rect 3386 2771 3410 2817
rect 3456 2771 3478 2817
rect 3386 2713 3478 2771
rect 3386 2661 3406 2713
rect 3458 2661 3478 2713
rect 3386 2647 3410 2661
rect 3456 2647 3478 2661
rect 3386 2621 3478 2647
rect 3599 2895 3634 2941
rect 3680 2895 3714 2941
rect 3858 3065 3904 3078
rect 3858 2941 3904 3019
rect 3599 2817 3714 2895
rect 3599 2771 3634 2817
rect 3680 2771 3714 2817
rect 3599 2693 3714 2771
rect 3599 2647 3634 2693
rect 3680 2647 3714 2693
rect 3151 2523 3186 2569
rect 3232 2523 3266 2569
rect 3151 2518 3266 2523
rect 3410 2569 3456 2621
rect 3186 2510 3232 2518
rect 3410 2510 3456 2523
rect 3599 2569 3714 2647
rect 3834 2899 3858 2929
rect 4047 3065 4162 3152
rect 4378 3149 4657 3162
rect 4457 3125 4657 3149
rect 4047 3019 4082 3065
rect 4128 3019 4162 3065
rect 4047 2941 4162 3019
rect 3904 2899 3926 2929
rect 3834 2847 3854 2899
rect 3906 2847 3926 2899
rect 3834 2817 3926 2847
rect 3834 2771 3858 2817
rect 3904 2771 3926 2817
rect 3834 2713 3926 2771
rect 3834 2661 3854 2713
rect 3906 2661 3926 2713
rect 3834 2647 3858 2661
rect 3904 2647 3926 2661
rect 3834 2621 3926 2647
rect 4047 2895 4082 2941
rect 4128 2895 4162 2941
rect 4306 3065 4352 3078
rect 4306 2941 4352 3019
rect 4047 2817 4162 2895
rect 4047 2771 4082 2817
rect 4128 2771 4162 2817
rect 4047 2693 4162 2771
rect 4047 2647 4082 2693
rect 4128 2647 4162 2693
rect 3599 2523 3634 2569
rect 3680 2523 3714 2569
rect 3599 2518 3714 2523
rect 3858 2569 3904 2621
rect 3634 2510 3680 2518
rect 3858 2510 3904 2523
rect 4047 2569 4162 2647
rect 4271 2899 4306 2929
rect 4271 2847 4291 2899
rect 4352 2895 4363 2929
rect 4343 2847 4363 2895
rect 4271 2817 4363 2847
rect 4271 2771 4306 2817
rect 4352 2771 4363 2817
rect 4271 2713 4363 2771
rect 4271 2661 4291 2713
rect 4343 2693 4363 2713
rect 4271 2647 4306 2661
rect 4352 2647 4363 2693
rect 4271 2621 4363 2647
rect 4047 2523 4082 2569
rect 4128 2523 4162 2569
rect 4047 2518 4162 2523
rect 4306 2569 4352 2621
rect 4082 2510 4128 2518
rect 4306 2510 4352 2523
rect 4844 2438 4916 5159
rect 2064 2401 4916 2438
rect 2064 2355 2663 2401
rect 2709 2355 2966 2401
rect 3012 2355 3412 2401
rect 3458 2355 3864 2401
rect 3910 2355 4156 2401
rect 4202 2355 4916 2401
rect 2064 2318 4916 2355
rect 1844 2160 1892 2206
rect 1938 2160 1986 2206
rect 1844 2094 1986 2160
rect 3608 2161 3700 2201
rect 2959 2143 3005 2156
rect 1844 2093 1987 2094
rect 1844 2043 2619 2093
rect 1844 1997 1892 2043
rect 1938 1997 2050 2043
rect 2096 1997 2208 2043
rect 2254 1997 2366 2043
rect 2412 1997 2524 2043
rect 2570 1997 2619 2043
rect 2959 2029 3005 2097
rect 3183 2143 3229 2156
rect 1844 1946 2619 1997
rect 2477 1908 2619 1946
rect 2477 1856 2543 1908
rect 2595 1856 2619 1908
rect 2477 1789 2619 1856
rect 2477 1743 2524 1789
rect 2570 1743 2619 1789
rect 2477 1722 2619 1743
rect 2477 1670 2543 1722
rect 2595 1670 2619 1722
rect 2941 2015 3033 2029
rect 2941 1969 2959 2015
rect 3005 1989 3033 2015
rect 2941 1937 2961 1969
rect 3013 1937 3033 1989
rect 2941 1888 3033 1937
rect 2941 1842 2959 1888
rect 3005 1842 3033 1888
rect 2941 1803 3033 1842
rect 2941 1761 2961 1803
rect 2941 1721 2959 1761
rect 3013 1751 3033 1803
rect 3005 1721 3033 1751
rect 3183 2015 3229 2097
rect 3407 2143 3453 2156
rect 3407 2030 3453 2097
rect 3608 2109 3628 2161
rect 3680 2109 3700 2161
rect 4054 2161 4146 2201
rect 3608 2097 3631 2109
rect 3677 2097 3700 2109
rect 3183 1888 3229 1969
rect 3183 1761 3229 1842
rect 2959 1702 3005 1715
rect 2477 1626 2619 1670
rect 2477 1580 2524 1626
rect 2570 1580 2619 1626
rect 2477 1462 2619 1580
rect 2749 1577 3057 1597
rect 2749 1525 2779 1577
rect 2831 1574 2965 1577
rect 3017 1574 3057 1577
rect 2831 1528 2889 1574
rect 3029 1528 3057 1574
rect 2831 1525 2965 1528
rect 3017 1525 3057 1528
rect 2749 1505 3057 1525
rect 3183 1585 3229 1715
rect 3386 2015 3478 2030
rect 3386 1990 3407 2015
rect 3453 1990 3478 2015
rect 3386 1938 3406 1990
rect 3458 1938 3478 1990
rect 3386 1888 3478 1938
rect 3608 2015 3700 2097
rect 3855 2143 3901 2156
rect 3855 2030 3901 2097
rect 4054 2109 4074 2161
rect 4126 2109 4146 2161
rect 4054 2097 4079 2109
rect 4125 2097 4146 2109
rect 3608 1975 3631 2015
rect 3677 1975 3700 2015
rect 3608 1923 3628 1975
rect 3680 1923 3700 1975
rect 3608 1893 3700 1923
rect 3828 2015 3920 2030
rect 3828 1990 3855 2015
rect 3828 1938 3848 1990
rect 3901 1969 3920 2015
rect 3900 1938 3920 1969
rect 3386 1842 3407 1888
rect 3453 1842 3478 1888
rect 3386 1804 3478 1842
rect 3386 1752 3406 1804
rect 3458 1752 3478 1804
rect 3386 1715 3407 1752
rect 3453 1715 3478 1752
rect 3386 1711 3478 1715
rect 3631 1888 3677 1893
rect 3631 1761 3677 1842
rect 3407 1702 3453 1711
rect 3631 1702 3677 1715
rect 3828 1888 3920 1938
rect 4054 2015 4146 2097
rect 4303 2143 4349 2156
rect 4303 2030 4349 2097
rect 4054 1975 4079 2015
rect 4125 1975 4146 2015
rect 4054 1923 4074 1975
rect 4126 1923 4146 1975
rect 4054 1893 4146 1923
rect 4276 2015 4368 2030
rect 4276 1990 4303 2015
rect 4276 1938 4296 1990
rect 4349 1969 4368 2015
rect 4348 1938 4368 1969
rect 3828 1842 3855 1888
rect 3901 1842 3920 1888
rect 3828 1804 3920 1842
rect 3828 1752 3848 1804
rect 3900 1761 3920 1804
rect 3828 1715 3855 1752
rect 3901 1715 3920 1761
rect 3828 1711 3920 1715
rect 4079 1888 4125 1893
rect 4079 1761 4125 1842
rect 3855 1702 3901 1711
rect 4079 1702 4125 1715
rect 4276 1888 4368 1938
rect 4276 1842 4303 1888
rect 4349 1842 4368 1888
rect 4276 1804 4368 1842
rect 4276 1752 4296 1804
rect 4348 1761 4368 1804
rect 4276 1715 4303 1752
rect 4349 1715 4368 1761
rect 4276 1711 4368 1715
rect 4303 1702 4349 1711
rect 3183 1574 3700 1585
rect 3183 1528 3549 1574
rect 3689 1528 3700 1574
rect 3183 1517 3700 1528
rect 4251 1566 4559 1586
rect 2477 1416 2524 1462
rect 2570 1416 2619 1462
rect 2477 1299 2619 1416
rect 2477 1253 2524 1299
rect 2570 1253 2619 1299
rect 2477 1136 2619 1253
rect 2477 1090 2524 1136
rect 2570 1105 2619 1136
rect 2477 1053 2543 1090
rect 2595 1053 2619 1105
rect 2477 972 2619 1053
rect 2477 926 2524 972
rect 2570 926 2619 972
rect 2477 919 2619 926
rect 2477 867 2543 919
rect 2595 867 2619 919
rect 2477 809 2619 867
rect 2477 763 2524 809
rect 2570 763 2619 809
rect 2477 646 2619 763
rect 2477 600 2524 646
rect 2570 600 2619 646
rect 2477 482 2619 600
rect 2925 1318 3040 1331
rect 2925 1272 2959 1318
rect 3005 1272 3040 1318
rect 2925 1190 3040 1272
rect 2925 1144 2959 1190
rect 3005 1144 3040 1190
rect 2925 1063 3040 1144
rect 2925 1017 2959 1063
rect 3005 1017 3040 1063
rect 2925 936 3040 1017
rect 2925 890 2959 936
rect 3005 890 3040 936
rect 2925 661 3040 890
rect 3183 1318 3229 1517
rect 4251 1514 4281 1566
rect 4333 1562 4467 1566
rect 4430 1516 4467 1562
rect 4333 1514 4467 1516
rect 4519 1514 4559 1566
rect 4251 1494 4559 1514
rect 3183 1190 3229 1272
rect 3183 1063 3229 1144
rect 3183 936 3229 1017
rect 3183 877 3229 890
rect 3373 1318 3488 1331
rect 3373 1272 3407 1318
rect 3453 1272 3488 1318
rect 3373 1190 3488 1272
rect 3373 1144 3407 1190
rect 3453 1144 3488 1190
rect 3373 1063 3488 1144
rect 3373 1017 3407 1063
rect 3453 1017 3488 1063
rect 3601 1318 3693 1336
rect 3601 1296 3631 1318
rect 3601 1244 3621 1296
rect 3677 1272 3693 1318
rect 3673 1244 3693 1272
rect 3601 1190 3693 1244
rect 3601 1144 3631 1190
rect 3677 1144 3693 1190
rect 3601 1110 3693 1144
rect 3601 1058 3621 1110
rect 3673 1063 3693 1110
rect 3601 1017 3631 1058
rect 3677 1017 3693 1063
rect 3820 1318 3936 1331
rect 3820 1272 3855 1318
rect 3901 1272 3936 1318
rect 3820 1190 3936 1272
rect 3820 1144 3855 1190
rect 3901 1144 3936 1190
rect 3820 1063 3936 1144
rect 3820 1017 3855 1063
rect 3901 1017 3936 1063
rect 4061 1318 4153 1336
rect 4061 1272 4079 1318
rect 4125 1296 4153 1318
rect 4061 1244 4081 1272
rect 4133 1244 4153 1296
rect 4061 1190 4153 1244
rect 4061 1144 4079 1190
rect 4125 1144 4153 1190
rect 4061 1110 4153 1144
rect 4061 1063 4081 1110
rect 4061 1017 4079 1063
rect 4133 1058 4153 1110
rect 4125 1017 4153 1058
rect 4268 1318 4384 1331
rect 4268 1272 4303 1318
rect 4349 1272 4384 1318
rect 4268 1190 4384 1272
rect 4268 1144 4303 1190
rect 4349 1144 4384 1190
rect 4268 1063 4384 1144
rect 4268 1017 4303 1063
rect 4349 1017 4384 1063
rect 3373 936 3488 1017
rect 3373 890 3407 936
rect 3453 890 3488 936
rect 3373 661 3488 890
rect 3631 936 3677 1017
rect 3631 877 3677 890
rect 3820 936 3936 1017
rect 3820 890 3855 936
rect 3901 890 3936 936
rect 3820 661 3936 890
rect 4079 936 4125 1017
rect 4079 877 4125 890
rect 4268 936 4384 1017
rect 4268 890 4303 936
rect 4349 890 4384 936
rect 4268 661 4384 890
rect 2925 624 4384 661
rect 2925 578 3011 624
rect 3057 578 3170 624
rect 3216 578 3328 624
rect 3374 578 3486 624
rect 3532 578 3644 624
rect 3690 578 3802 624
rect 3848 578 3960 624
rect 4006 578 4118 624
rect 4164 578 4277 624
rect 4323 578 4384 624
rect 2925 545 4384 578
rect 2924 544 4384 545
rect 4883 1105 5025 1155
rect 4883 1053 4929 1105
rect 4981 1053 5025 1105
rect 4883 1009 4932 1053
rect 4978 1009 5025 1053
rect 4883 919 5025 1009
rect 4883 867 4929 919
rect 4981 867 5025 919
rect 4883 846 4932 867
rect 4978 846 5025 867
rect 4883 728 5025 846
rect 4883 682 4932 728
rect 4978 682 5025 728
rect 4883 565 5025 682
rect 2477 436 2524 482
rect 2570 436 2619 482
rect 2723 541 4570 544
rect 2723 522 3031 541
rect 2723 470 2761 522
rect 2813 470 2941 522
rect 2993 470 3031 522
rect 2723 448 3031 470
rect 3182 522 3490 541
rect 3182 470 3220 522
rect 3272 470 3400 522
rect 3452 470 3490 522
rect 3182 448 3490 470
rect 4262 522 4570 541
rect 4262 470 4300 522
rect 4352 470 4480 522
rect 4532 470 4570 522
rect 4262 448 4570 470
rect 4883 519 4932 565
rect 4978 519 5025 565
rect 2477 319 2619 436
rect 2477 273 2524 319
rect 2570 273 2619 319
rect 2477 225 2619 273
rect 4883 402 5025 519
rect 4883 356 4932 402
rect 4978 356 5025 402
rect 4883 225 5025 356
rect 2477 175 5025 225
rect 2477 129 2781 175
rect 2827 129 2939 175
rect 2985 129 3097 175
rect 3143 129 3256 175
rect 3302 129 3414 175
rect 3460 129 3572 175
rect 3618 129 3730 175
rect 3776 129 3888 175
rect 3934 129 4046 175
rect 4092 129 4205 175
rect 4251 129 4363 175
rect 4409 129 4521 175
rect 4567 129 5025 175
rect 2477 78 5025 129
<< via1 >>
rect 2355 7957 2407 8009
rect 2541 7957 2593 8009
rect 2981 7957 3033 8009
rect 3167 7957 3219 8009
rect 4219 7957 4271 8009
rect 4405 7957 4457 8009
rect 2737 7748 2789 7800
rect 2923 7748 2975 7800
rect 3541 7748 3593 7800
rect 3727 7748 3779 7800
rect 3410 7287 3462 7339
rect 2835 6688 2887 6740
rect 3408 6740 3460 6750
rect 3408 6698 3412 6740
rect 3412 6698 3458 6740
rect 3458 6698 3460 6740
rect 3970 6666 4022 6718
rect 2616 6400 2659 6424
rect 2659 6400 2668 6424
rect 2616 6372 2668 6400
rect 2616 6191 2668 6238
rect 2616 6186 2659 6191
rect 2659 6186 2668 6191
rect 3070 6451 3122 6503
rect 3070 6273 3076 6317
rect 3076 6273 3122 6317
rect 3070 6265 3122 6273
rect 3297 6400 3300 6424
rect 3300 6400 3346 6424
rect 3346 6400 3349 6424
rect 3297 6372 3349 6400
rect 3297 6191 3349 6238
rect 3297 6186 3300 6191
rect 3300 6186 3346 6191
rect 3346 6186 3349 6191
rect 3523 6400 3524 6424
rect 3524 6400 3570 6424
rect 3570 6400 3575 6424
rect 3523 6372 3575 6400
rect 3523 6191 3575 6238
rect 3523 6186 3524 6191
rect 3524 6186 3570 6191
rect 3570 6186 3575 6191
rect 3742 6451 3794 6503
rect 3742 6273 3748 6317
rect 3748 6273 3794 6317
rect 3742 6265 3794 6273
rect 4201 6400 4244 6424
rect 4244 6400 4253 6424
rect 4201 6372 4253 6400
rect 4201 6191 4253 6238
rect 4201 6186 4244 6191
rect 4244 6186 4253 6191
rect 3316 5984 3368 6036
rect 3503 5812 3555 5864
rect 2307 4948 2359 5000
rect 2307 4762 2359 4814
rect 2721 4925 2722 4943
rect 2722 4925 2768 4943
rect 2768 4925 2773 4943
rect 2721 4891 2773 4925
rect 2721 4721 2773 4757
rect 2721 4705 2764 4721
rect 2764 4705 2773 4721
rect 3171 4971 3223 5000
rect 3171 4948 3216 4971
rect 3216 4948 3223 4971
rect 3171 4762 3223 4814
rect 2722 4507 2774 4510
rect 2722 4461 2741 4507
rect 2741 4461 2774 4507
rect 2722 4458 2774 4461
rect 2902 4458 2954 4510
rect 3231 4507 3283 4510
rect 3231 4461 3264 4507
rect 3264 4461 3283 4507
rect 3231 4458 3283 4461
rect 2428 4246 2480 4298
rect 3643 4971 3695 5000
rect 3643 4948 3664 4971
rect 3664 4948 3695 4971
rect 3643 4762 3695 4814
rect 4060 4925 4066 4943
rect 4066 4925 4112 4943
rect 4060 4891 4112 4925
rect 4060 4723 4112 4757
rect 4060 4705 4102 4723
rect 4102 4705 4112 4723
rect 3587 4507 3639 4510
rect 3587 4461 3596 4507
rect 3596 4461 3639 4507
rect 3587 4458 3639 4461
rect 3921 4458 3973 4510
rect 4101 4507 4153 4510
rect 4101 4461 4143 4507
rect 4143 4461 4153 4507
rect 4101 4458 4153 4461
rect 4438 4948 4490 5000
rect 4438 4762 4490 4814
rect 4304 4457 4356 4509
rect 3121 4291 3173 4299
rect 3121 4247 3140 4291
rect 3140 4247 3173 4291
rect 3409 4247 3461 4299
rect 3697 4291 3749 4299
rect 3697 4247 3739 4291
rect 3739 4247 3749 4291
rect 4476 4246 4528 4298
rect 2394 3169 2446 3221
rect 4414 3169 4466 3221
rect 2521 2895 2560 2899
rect 2560 2895 2573 2899
rect 2521 2847 2573 2895
rect 2521 2693 2573 2713
rect 2521 2661 2560 2693
rect 2560 2661 2573 2693
rect 2958 2895 2962 2899
rect 2962 2895 3008 2899
rect 3008 2895 3010 2899
rect 2958 2847 3010 2895
rect 2958 2693 3010 2713
rect 2958 2661 2962 2693
rect 2962 2661 3008 2693
rect 3008 2661 3010 2693
rect 3406 2895 3410 2899
rect 3410 2895 3456 2899
rect 3456 2895 3458 2899
rect 3406 2847 3458 2895
rect 3406 2693 3458 2713
rect 3406 2661 3410 2693
rect 3410 2661 3456 2693
rect 3456 2661 3458 2693
rect 3854 2895 3858 2899
rect 3858 2895 3904 2899
rect 3904 2895 3906 2899
rect 3854 2847 3906 2895
rect 3854 2693 3906 2713
rect 3854 2661 3858 2693
rect 3858 2661 3904 2693
rect 3904 2661 3906 2693
rect 4291 2895 4306 2899
rect 4306 2895 4343 2899
rect 4291 2847 4343 2895
rect 4291 2693 4343 2713
rect 4291 2661 4306 2693
rect 4306 2661 4343 2693
rect 2543 1856 2595 1908
rect 2543 1670 2595 1722
rect 2961 1969 3005 1989
rect 3005 1969 3013 1989
rect 2961 1937 3013 1969
rect 2961 1761 3013 1803
rect 2961 1751 3005 1761
rect 3005 1751 3013 1761
rect 3628 2143 3680 2161
rect 3628 2109 3631 2143
rect 3631 2109 3677 2143
rect 3677 2109 3680 2143
rect 2779 1525 2831 1577
rect 2965 1574 3017 1577
rect 2965 1528 3017 1574
rect 2965 1525 3017 1528
rect 3406 1969 3407 1990
rect 3407 1969 3453 1990
rect 3453 1969 3458 1990
rect 3406 1938 3458 1969
rect 4074 2143 4126 2161
rect 4074 2109 4079 2143
rect 4079 2109 4125 2143
rect 4125 2109 4126 2143
rect 3628 1969 3631 1975
rect 3631 1969 3677 1975
rect 3677 1969 3680 1975
rect 3628 1923 3680 1969
rect 3848 1969 3855 1990
rect 3855 1969 3900 1990
rect 3848 1938 3900 1969
rect 3406 1761 3458 1804
rect 3406 1752 3407 1761
rect 3407 1752 3453 1761
rect 3453 1752 3458 1761
rect 4074 1969 4079 1975
rect 4079 1969 4125 1975
rect 4125 1969 4126 1975
rect 4074 1923 4126 1969
rect 4296 1969 4303 1990
rect 4303 1969 4348 1990
rect 4296 1938 4348 1969
rect 3848 1761 3900 1804
rect 3848 1752 3855 1761
rect 3855 1752 3900 1761
rect 4296 1761 4348 1804
rect 4296 1752 4303 1761
rect 4303 1752 4348 1761
rect 2543 1090 2570 1105
rect 2570 1090 2595 1105
rect 2543 1053 2595 1090
rect 2543 867 2595 919
rect 4281 1562 4333 1566
rect 4281 1516 4290 1562
rect 4290 1516 4333 1562
rect 4281 1514 4333 1516
rect 4467 1514 4519 1566
rect 3621 1272 3631 1296
rect 3631 1272 3673 1296
rect 3621 1244 3673 1272
rect 3621 1063 3673 1110
rect 3621 1058 3631 1063
rect 3631 1058 3673 1063
rect 4081 1272 4125 1296
rect 4125 1272 4133 1296
rect 4081 1244 4133 1272
rect 4081 1063 4133 1110
rect 4081 1058 4125 1063
rect 4125 1058 4133 1063
rect 4929 1055 4981 1105
rect 4929 1053 4932 1055
rect 4932 1053 4978 1055
rect 4978 1053 4981 1055
rect 4929 892 4981 919
rect 4929 867 4932 892
rect 4932 867 4978 892
rect 4978 867 4981 892
rect 2761 470 2813 522
rect 2941 470 2993 522
rect 3220 470 3272 522
rect 3400 470 3452 522
rect 4300 470 4352 522
rect 4480 470 4532 522
<< metal2 >>
rect 2433 8033 2522 8146
rect 3052 8033 3141 8146
rect 2432 8029 2522 8033
rect 3051 8029 3141 8033
rect 2325 8009 2633 8029
rect 2325 7957 2355 8009
rect 2407 7957 2541 8009
rect 2593 7957 2633 8009
rect 2325 7937 2633 7957
rect 2951 8011 3259 8029
rect 2951 7955 2979 8011
rect 3035 7955 3165 8011
rect 3221 7955 3259 8011
rect 2951 7937 3259 7955
rect 2432 7936 2522 7937
rect 3051 7936 3141 7937
rect 2812 7820 2906 7824
rect 3671 7820 3761 8146
rect 4290 8033 4380 8146
rect 3950 8029 4380 8033
rect 3950 8009 4497 8029
rect 3950 7957 4219 8009
rect 4271 7957 4405 8009
rect 4457 7957 4497 8009
rect 3950 7937 4497 7957
rect 3950 7936 4380 7937
rect 1684 7802 1992 7820
rect 1684 7746 1712 7802
rect 1768 7746 1898 7802
rect 1954 7746 1992 7802
rect 1684 7728 1992 7746
rect 2707 7800 3015 7820
rect 2707 7748 2737 7800
rect 2789 7748 2923 7800
rect 2975 7748 3015 7800
rect 2707 7728 3015 7748
rect 3511 7800 3819 7820
rect 3511 7748 3541 7800
rect 3593 7748 3727 7800
rect 3779 7748 3819 7800
rect 3511 7728 3819 7748
rect 2812 7727 2906 7728
rect 3671 7727 3761 7728
rect 2813 6763 2906 7727
rect 3373 7339 3501 7362
rect 3373 7287 3410 7339
rect 3462 7287 3501 7339
rect 3373 7265 3501 7287
rect 2798 6740 2926 6763
rect 2798 6688 2835 6740
rect 2887 6688 2926 6740
rect 2798 6666 2926 6688
rect 3388 6750 3482 7265
rect 3388 6698 3408 6750
rect 3460 6698 3482 6750
rect 3950 6741 4044 7936
rect 3388 6657 3482 6698
rect 3933 6718 4061 6741
rect 3933 6666 3970 6718
rect 4022 6666 4061 6718
rect 3933 6644 4061 6666
rect 3050 6505 3142 6533
rect 2595 6424 2688 6464
rect 2595 6372 2616 6424
rect 2668 6372 2688 6424
rect 2595 6238 2688 6372
rect 2595 6186 2616 6238
rect 2668 6186 2688 6238
rect 3050 6449 3068 6505
rect 3124 6449 3142 6505
rect 3722 6505 3814 6533
rect 3050 6319 3142 6449
rect 3050 6263 3068 6319
rect 3124 6263 3142 6319
rect 3050 6225 3142 6263
rect 3277 6424 3369 6464
rect 3277 6372 3297 6424
rect 3349 6372 3369 6424
rect 3277 6238 3369 6372
rect 2595 6146 2688 6186
rect 3277 6186 3297 6238
rect 3349 6186 3369 6238
rect 3277 6172 3369 6186
rect 3503 6424 3595 6464
rect 3503 6372 3523 6424
rect 3575 6372 3595 6424
rect 3503 6238 3595 6372
rect 3503 6186 3523 6238
rect 3575 6186 3595 6238
rect 3722 6449 3740 6505
rect 3796 6449 3814 6505
rect 3722 6319 3814 6449
rect 3722 6263 3740 6319
rect 3796 6263 3814 6319
rect 3722 6225 3814 6263
rect 4181 6424 4274 6464
rect 4181 6372 4201 6424
rect 4253 6372 4274 6424
rect 4181 6238 4274 6372
rect 3503 6172 3595 6186
rect 4181 6186 4201 6238
rect 4253 6186 4274 6238
rect 2595 6061 2685 6146
rect 2071 5968 2685 6061
rect 3276 6057 3370 6172
rect 3276 6036 3403 6057
rect 3276 5984 3316 6036
rect 3368 5984 3403 6036
rect 2071 4533 2160 5968
rect 3276 5964 3403 5984
rect 3276 5791 3370 5964
rect 3502 5885 3596 6172
rect 4181 6063 4274 6186
rect 4181 5966 4696 6063
rect 3468 5864 3596 5885
rect 3468 5812 3503 5864
rect 3555 5812 3596 5864
rect 3468 5792 3596 5812
rect 3502 5791 3596 5792
rect 2287 5002 2379 5030
rect 2287 4946 2305 5002
rect 2361 4946 2379 5002
rect 3151 5002 3243 5030
rect 2287 4816 2379 4946
rect 2287 4760 2305 4816
rect 2361 4760 2379 4816
rect 2287 4722 2379 4760
rect 2701 4945 2793 4973
rect 2701 4889 2719 4945
rect 2775 4889 2793 4945
rect 2701 4759 2793 4889
rect 2701 4703 2719 4759
rect 2775 4703 2793 4759
rect 3151 4946 3169 5002
rect 3225 4946 3243 5002
rect 3151 4816 3243 4946
rect 3151 4760 3169 4816
rect 3225 4760 3243 4816
rect 3151 4722 3243 4760
rect 3623 5002 3715 5030
rect 3623 4946 3641 5002
rect 3697 4946 3715 5002
rect 4418 5002 4510 5030
rect 3623 4816 3715 4946
rect 3623 4760 3641 4816
rect 3697 4760 3715 4816
rect 3623 4722 3715 4760
rect 4040 4945 4132 4973
rect 4040 4889 4058 4945
rect 4114 4889 4132 4945
rect 4040 4759 4132 4889
rect 2701 4665 2793 4703
rect 4040 4703 4058 4759
rect 4114 4703 4132 4759
rect 4418 4946 4436 5002
rect 4492 4946 4510 5002
rect 4418 4816 4510 4946
rect 4418 4760 4436 4816
rect 4492 4760 4510 4816
rect 4418 4722 4510 4760
rect 4040 4665 4132 4703
rect 2071 4510 4461 4533
rect 2071 4458 2722 4510
rect 2774 4458 2902 4510
rect 2954 4458 3231 4510
rect 3283 4458 3587 4510
rect 3639 4458 3921 4510
rect 3973 4458 4101 4510
rect 4153 4509 4461 4510
rect 4153 4458 4304 4509
rect 2071 4457 4304 4458
rect 4356 4457 4461 4509
rect 2071 4436 4461 4457
rect 2071 2309 2160 4436
rect 4602 4322 4696 5966
rect 2388 4299 4696 4322
rect 2388 4298 3121 4299
rect 2388 4246 2428 4298
rect 2480 4247 3121 4298
rect 3173 4247 3409 4299
rect 3461 4247 3697 4299
rect 3749 4298 4696 4299
rect 3749 4247 4476 4298
rect 2480 4246 4476 4247
rect 4528 4246 4696 4298
rect 2388 4225 4696 4246
rect 2358 3221 2698 3245
rect 2358 3150 2394 3221
rect 2446 3206 2698 3221
rect 2450 3150 2606 3206
rect 2662 3150 2698 3206
rect 2358 3111 2698 3150
rect 4167 3221 4507 3245
rect 4167 3206 4414 3221
rect 4466 3206 4507 3221
rect 4167 3150 4203 3206
rect 4259 3169 4414 3206
rect 4259 3150 4415 3169
rect 4471 3150 4507 3206
rect 4167 3111 4507 3150
rect 2501 2901 2593 2929
rect 2501 2845 2519 2901
rect 2575 2845 2593 2901
rect 2501 2715 2593 2845
rect 2501 2659 2519 2715
rect 2575 2659 2593 2715
rect 2501 2621 2593 2659
rect 2938 2901 3030 2929
rect 2938 2845 2956 2901
rect 3012 2845 3030 2901
rect 2938 2715 3030 2845
rect 2938 2659 2956 2715
rect 3012 2659 3030 2715
rect 2938 2621 3030 2659
rect 3386 2901 3478 2929
rect 3386 2845 3404 2901
rect 3460 2845 3478 2901
rect 3386 2715 3478 2845
rect 3386 2659 3404 2715
rect 3460 2659 3478 2715
rect 3386 2621 3478 2659
rect 3834 2901 3926 2929
rect 3834 2845 3852 2901
rect 3908 2845 3926 2901
rect 3834 2715 3926 2845
rect 3834 2659 3852 2715
rect 3908 2659 3926 2715
rect 3834 2621 3926 2659
rect 4271 2901 4363 2929
rect 4271 2845 4289 2901
rect 4345 2845 4363 2901
rect 4271 2715 4363 2845
rect 4271 2659 4289 2715
rect 4345 2659 4363 2715
rect 4271 2621 4363 2659
rect 4602 2311 4696 4225
rect 2071 2216 2838 2309
rect 2523 1910 2615 1938
rect 2523 1854 2541 1910
rect 2597 1854 2615 1910
rect 2523 1724 2615 1854
rect 2523 1668 2541 1724
rect 2597 1668 2615 1724
rect 2523 1630 2615 1668
rect 2749 1597 2838 2216
rect 4279 2214 4907 2311
rect 3608 2163 3700 2201
rect 3608 2107 3626 2163
rect 3682 2107 3700 2163
rect 2941 1991 3033 2029
rect 2941 1935 2959 1991
rect 3015 1935 3033 1991
rect 2941 1805 3033 1935
rect 2941 1749 2959 1805
rect 3015 1749 3033 1805
rect 2941 1721 3033 1749
rect 3386 1990 3479 2030
rect 3386 1938 3406 1990
rect 3458 1938 3479 1990
rect 3386 1804 3479 1938
rect 3608 1977 3700 2107
rect 4054 2163 4146 2201
rect 4054 2107 4072 2163
rect 4128 2107 4146 2163
rect 3608 1921 3626 1977
rect 3682 1921 3700 1977
rect 3608 1893 3700 1921
rect 3827 1990 3921 2030
rect 3827 1938 3848 1990
rect 3900 1938 3921 1990
rect 3386 1752 3406 1804
rect 3458 1781 3479 1804
rect 3827 1804 3921 1938
rect 4054 1977 4146 2107
rect 4054 1921 4072 1977
rect 4128 1921 4146 1977
rect 4054 1893 4146 1921
rect 4275 1990 4369 2030
rect 4275 1938 4296 1990
rect 4348 1938 4369 1990
rect 3458 1780 3480 1781
rect 3827 1780 3848 1804
rect 3458 1752 3848 1780
rect 3900 1752 3921 1804
rect 4275 1804 4369 1938
rect 4275 1780 4296 1804
rect 3386 1683 3921 1752
rect 4060 1752 4296 1780
rect 4348 1752 4369 1804
rect 4060 1683 4369 1752
rect 2749 1577 3057 1597
rect 2749 1525 2779 1577
rect 2831 1525 2965 1577
rect 3017 1525 3057 1577
rect 2749 1505 3057 1525
rect 2749 1504 2838 1505
rect 3601 1296 3695 1683
rect 3601 1244 3621 1296
rect 3673 1244 3695 1296
rect 2523 1107 2615 1135
rect 2523 1051 2541 1107
rect 2597 1051 2615 1107
rect 2523 921 2615 1051
rect 2523 865 2541 921
rect 2597 865 2615 921
rect 2523 827 2615 865
rect 3601 1110 3695 1244
rect 3601 1058 3621 1110
rect 3673 1058 3695 1110
rect 2723 524 3031 545
rect 2723 468 2759 524
rect 2815 468 2939 524
rect 2995 468 3031 524
rect 2723 448 3031 468
rect 3182 524 3490 545
rect 3182 468 3218 524
rect 3274 468 3398 524
rect 3454 468 3490 524
rect 3182 448 3490 468
rect 3601 -196 3695 1058
rect 4060 1296 4154 1683
rect 4466 1586 4560 2214
rect 4251 1566 4560 1586
rect 4251 1514 4281 1566
rect 4333 1514 4467 1566
rect 4519 1514 4560 1566
rect 4251 1504 4560 1514
rect 4251 1494 4559 1504
rect 4060 1244 4081 1296
rect 4133 1244 4154 1296
rect 4060 1110 4154 1244
rect 4060 1058 4081 1110
rect 4133 1058 4154 1110
rect 4060 -196 4154 1058
rect 4909 1107 5001 1135
rect 4909 1051 4927 1107
rect 4983 1051 5001 1107
rect 4909 921 5001 1051
rect 4909 865 4927 921
rect 4983 865 5001 921
rect 4909 827 5001 865
rect 4262 524 4570 545
rect 4262 468 4298 524
rect 4354 468 4478 524
rect 4534 468 4570 524
rect 4262 448 4570 468
<< via2 >>
rect 2979 8009 3035 8011
rect 2979 7957 2981 8009
rect 2981 7957 3033 8009
rect 3033 7957 3035 8009
rect 2979 7955 3035 7957
rect 3165 8009 3221 8011
rect 3165 7957 3167 8009
rect 3167 7957 3219 8009
rect 3219 7957 3221 8009
rect 3165 7955 3221 7957
rect 1712 7746 1768 7802
rect 1898 7746 1954 7802
rect 3068 6503 3124 6505
rect 3068 6451 3070 6503
rect 3070 6451 3122 6503
rect 3122 6451 3124 6503
rect 3068 6449 3124 6451
rect 3068 6317 3124 6319
rect 3068 6265 3070 6317
rect 3070 6265 3122 6317
rect 3122 6265 3124 6317
rect 3068 6263 3124 6265
rect 3740 6503 3796 6505
rect 3740 6451 3742 6503
rect 3742 6451 3794 6503
rect 3794 6451 3796 6503
rect 3740 6449 3796 6451
rect 3740 6317 3796 6319
rect 3740 6265 3742 6317
rect 3742 6265 3794 6317
rect 3794 6265 3796 6317
rect 3740 6263 3796 6265
rect 2305 5000 2361 5002
rect 2305 4948 2307 5000
rect 2307 4948 2359 5000
rect 2359 4948 2361 5000
rect 2305 4946 2361 4948
rect 2305 4814 2361 4816
rect 2305 4762 2307 4814
rect 2307 4762 2359 4814
rect 2359 4762 2361 4814
rect 2305 4760 2361 4762
rect 2719 4943 2775 4945
rect 2719 4891 2721 4943
rect 2721 4891 2773 4943
rect 2773 4891 2775 4943
rect 2719 4889 2775 4891
rect 2719 4757 2775 4759
rect 2719 4705 2721 4757
rect 2721 4705 2773 4757
rect 2773 4705 2775 4757
rect 2719 4703 2775 4705
rect 3169 5000 3225 5002
rect 3169 4948 3171 5000
rect 3171 4948 3223 5000
rect 3223 4948 3225 5000
rect 3169 4946 3225 4948
rect 3169 4814 3225 4816
rect 3169 4762 3171 4814
rect 3171 4762 3223 4814
rect 3223 4762 3225 4814
rect 3169 4760 3225 4762
rect 3641 5000 3697 5002
rect 3641 4948 3643 5000
rect 3643 4948 3695 5000
rect 3695 4948 3697 5000
rect 3641 4946 3697 4948
rect 3641 4814 3697 4816
rect 3641 4762 3643 4814
rect 3643 4762 3695 4814
rect 3695 4762 3697 4814
rect 3641 4760 3697 4762
rect 4058 4943 4114 4945
rect 4058 4891 4060 4943
rect 4060 4891 4112 4943
rect 4112 4891 4114 4943
rect 4058 4889 4114 4891
rect 4058 4757 4114 4759
rect 4058 4705 4060 4757
rect 4060 4705 4112 4757
rect 4112 4705 4114 4757
rect 4058 4703 4114 4705
rect 4436 5000 4492 5002
rect 4436 4948 4438 5000
rect 4438 4948 4490 5000
rect 4490 4948 4492 5000
rect 4436 4946 4492 4948
rect 4436 4814 4492 4816
rect 4436 4762 4438 4814
rect 4438 4762 4490 4814
rect 4490 4762 4492 4814
rect 4436 4760 4492 4762
rect 2394 3169 2446 3206
rect 2446 3169 2450 3206
rect 2394 3150 2450 3169
rect 2606 3150 2662 3206
rect 4203 3150 4259 3206
rect 4415 3169 4466 3206
rect 4466 3169 4471 3206
rect 4415 3150 4471 3169
rect 2519 2899 2575 2901
rect 2519 2847 2521 2899
rect 2521 2847 2573 2899
rect 2573 2847 2575 2899
rect 2519 2845 2575 2847
rect 2519 2713 2575 2715
rect 2519 2661 2521 2713
rect 2521 2661 2573 2713
rect 2573 2661 2575 2713
rect 2519 2659 2575 2661
rect 2956 2899 3012 2901
rect 2956 2847 2958 2899
rect 2958 2847 3010 2899
rect 3010 2847 3012 2899
rect 2956 2845 3012 2847
rect 2956 2713 3012 2715
rect 2956 2661 2958 2713
rect 2958 2661 3010 2713
rect 3010 2661 3012 2713
rect 2956 2659 3012 2661
rect 3404 2899 3460 2901
rect 3404 2847 3406 2899
rect 3406 2847 3458 2899
rect 3458 2847 3460 2899
rect 3404 2845 3460 2847
rect 3404 2713 3460 2715
rect 3404 2661 3406 2713
rect 3406 2661 3458 2713
rect 3458 2661 3460 2713
rect 3404 2659 3460 2661
rect 3852 2899 3908 2901
rect 3852 2847 3854 2899
rect 3854 2847 3906 2899
rect 3906 2847 3908 2899
rect 3852 2845 3908 2847
rect 3852 2713 3908 2715
rect 3852 2661 3854 2713
rect 3854 2661 3906 2713
rect 3906 2661 3908 2713
rect 3852 2659 3908 2661
rect 4289 2899 4345 2901
rect 4289 2847 4291 2899
rect 4291 2847 4343 2899
rect 4343 2847 4345 2899
rect 4289 2845 4345 2847
rect 4289 2713 4345 2715
rect 4289 2661 4291 2713
rect 4291 2661 4343 2713
rect 4343 2661 4345 2713
rect 4289 2659 4345 2661
rect 2541 1908 2597 1910
rect 2541 1856 2543 1908
rect 2543 1856 2595 1908
rect 2595 1856 2597 1908
rect 2541 1854 2597 1856
rect 2541 1722 2597 1724
rect 2541 1670 2543 1722
rect 2543 1670 2595 1722
rect 2595 1670 2597 1722
rect 2541 1668 2597 1670
rect 3626 2161 3682 2163
rect 3626 2109 3628 2161
rect 3628 2109 3680 2161
rect 3680 2109 3682 2161
rect 3626 2107 3682 2109
rect 2959 1989 3015 1991
rect 2959 1937 2961 1989
rect 2961 1937 3013 1989
rect 3013 1937 3015 1989
rect 2959 1935 3015 1937
rect 2959 1803 3015 1805
rect 2959 1751 2961 1803
rect 2961 1751 3013 1803
rect 3013 1751 3015 1803
rect 2959 1749 3015 1751
rect 4072 2161 4128 2163
rect 4072 2109 4074 2161
rect 4074 2109 4126 2161
rect 4126 2109 4128 2161
rect 4072 2107 4128 2109
rect 3626 1975 3682 1977
rect 3626 1923 3628 1975
rect 3628 1923 3680 1975
rect 3680 1923 3682 1975
rect 3626 1921 3682 1923
rect 4072 1975 4128 1977
rect 4072 1923 4074 1975
rect 4074 1923 4126 1975
rect 4126 1923 4128 1975
rect 4072 1921 4128 1923
rect 2541 1105 2597 1107
rect 2541 1053 2543 1105
rect 2543 1053 2595 1105
rect 2595 1053 2597 1105
rect 2541 1051 2597 1053
rect 2541 919 2597 921
rect 2541 867 2543 919
rect 2543 867 2595 919
rect 2595 867 2597 919
rect 2541 865 2597 867
rect 2759 522 2815 524
rect 2759 470 2761 522
rect 2761 470 2813 522
rect 2813 470 2815 522
rect 2759 468 2815 470
rect 2939 522 2995 524
rect 2939 470 2941 522
rect 2941 470 2993 522
rect 2993 470 2995 522
rect 2939 468 2995 470
rect 3218 522 3274 524
rect 3218 470 3220 522
rect 3220 470 3272 522
rect 3272 470 3274 522
rect 3218 468 3274 470
rect 3398 522 3454 524
rect 3398 470 3400 522
rect 3400 470 3452 522
rect 3452 470 3454 522
rect 3398 468 3454 470
rect 4927 1105 4983 1107
rect 4927 1053 4929 1105
rect 4929 1053 4981 1105
rect 4981 1053 4983 1105
rect 4927 1051 4983 1053
rect 4927 919 4983 921
rect 4927 867 4929 919
rect 4929 867 4981 919
rect 4981 867 4983 919
rect 4927 865 4983 867
rect 4298 522 4354 524
rect 4298 470 4300 522
rect 4300 470 4352 522
rect 4352 470 4354 522
rect 4298 468 4354 470
rect 4478 522 4534 524
rect 4478 470 4480 522
rect 4480 470 4532 522
rect 4532 470 4534 522
rect 4478 468 4534 470
<< metal3 >>
rect 2430 8030 3130 8033
rect 2430 8011 3260 8030
rect 2430 7955 2979 8011
rect 3035 7955 3165 8011
rect 3221 7955 3260 8011
rect 2430 7937 3260 7955
rect 2430 7936 3130 7937
rect 2430 7824 2524 7936
rect 1684 7802 2524 7824
rect 1684 7746 1712 7802
rect 1768 7746 1898 7802
rect 1954 7746 2524 7802
rect 1684 7727 2524 7746
rect -356 6505 4955 7106
rect -356 6449 3068 6505
rect 3124 6449 3740 6505
rect 3796 6449 4955 6505
rect -356 6319 4955 6449
rect -356 6263 3068 6319
rect 3124 6263 3740 6319
rect 3796 6263 4955 6319
rect -356 5002 4955 6263
rect -356 4946 2305 5002
rect 2361 4946 3169 5002
rect 3225 4946 3641 5002
rect 3697 4946 4436 5002
rect 4492 4946 4955 5002
rect -356 4945 4955 4946
rect -356 4889 2719 4945
rect 2775 4889 4058 4945
rect 4114 4889 4955 4945
rect -356 4816 4955 4889
rect -356 4760 2305 4816
rect 2361 4760 3169 4816
rect 3225 4760 3641 4816
rect 3697 4760 4436 4816
rect 4492 4760 4955 4816
rect -356 4759 4955 4760
rect -356 4703 2719 4759
rect 2775 4703 4058 4759
rect 4114 4703 4955 4759
rect -356 4383 4955 4703
rect -356 3206 5006 4097
rect -356 3150 2394 3206
rect 2450 3150 2606 3206
rect 2662 3150 4203 3206
rect 4259 3150 4415 3206
rect 4471 3150 5006 3206
rect -356 2901 5006 3150
rect -356 2845 2519 2901
rect 2575 2845 2956 2901
rect 3012 2845 3404 2901
rect 3460 2845 3852 2901
rect 3908 2845 4289 2901
rect 4345 2845 5006 2901
rect -356 2715 5006 2845
rect -356 2659 2519 2715
rect 2575 2659 2956 2715
rect 3012 2659 3404 2715
rect 3460 2659 3852 2715
rect 3908 2659 4289 2715
rect 4345 2659 5006 2715
rect -356 2163 5006 2659
rect -356 2107 3626 2163
rect 3682 2107 4072 2163
rect 4128 2107 5006 2163
rect -356 1991 5006 2107
rect -356 1935 2959 1991
rect 3015 1977 5006 1991
rect 3015 1935 3626 1977
rect -356 1921 3626 1935
rect 3682 1921 4072 1977
rect 4128 1921 5006 1977
rect -356 1910 5006 1921
rect -356 1854 2541 1910
rect 2597 1854 5006 1910
rect -356 1805 5006 1854
rect -356 1749 2959 1805
rect 3015 1749 5006 1805
rect -356 1724 5006 1749
rect -356 1668 2541 1724
rect 2597 1668 5006 1724
rect -356 1107 5006 1668
rect -356 1051 2541 1107
rect 2597 1051 4927 1107
rect 4983 1051 5006 1107
rect -356 951 5006 1051
rect -357 921 5006 951
rect -357 865 2541 921
rect 2597 865 4927 921
rect 4983 865 5006 921
rect -357 817 5006 865
rect -356 695 5006 817
rect -356 524 5006 545
rect -356 468 2759 524
rect 2815 468 2939 524
rect 2995 468 3218 524
rect 3274 468 3398 524
rect 3454 468 4298 524
rect 4354 468 4478 524
rect 4534 468 5006 524
rect -356 -172 5006 468
use M1_NWELL$$44998700_R90_256x8m81  M1_NWELL$$44998700_R90_256x8m81_0
timestamp 1698431365
transform 0 -1 2322 1 0 4888
box 0 0 1 1
use M1_NWELL$$44998700_R90_256x8m81  M1_NWELL$$44998700_R90_256x8m81_1
timestamp 1698431365
transform 0 -1 4475 1 0 4888
box 0 0 1 1
use M1_NWELL$$46278700_256x8m81  M1_NWELL$$46278700_256x8m81_0
timestamp 1698431365
transform 1 0 3667 0 1 601
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_0
timestamp 1698431365
transform -1 0 3887 0 1 2378
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_1
timestamp 1698431365
transform -1 0 4179 0 1 2378
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_2
timestamp 1698431365
transform 1 0 4515 0 1 3185
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_3
timestamp 1698431365
transform -1 0 2989 0 1 2378
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_4
timestamp 1698431365
transform 1 0 2354 0 1 3185
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_5
timestamp 1698431365
transform 1 0 2686 0 1 2378
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_6
timestamp 1698431365
transform -1 0 3435 0 1 2378
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_0
timestamp 1698431365
transform 1 0 3287 0 1 4484
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_1
timestamp 1698431365
transform 1 0 3117 0 1 4268
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_2
timestamp 1698431365
transform 1 0 2741 0 1 4698
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_3
timestamp 1698431365
transform 1 0 2137 0 1 5193
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_4
timestamp 1698431365
transform 1 0 2718 0 1 4484
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_5
timestamp 1698431365
transform 1 0 4677 0 1 5193
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_6
timestamp 1698431365
transform 1 0 3435 0 1 6717
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_7
timestamp 1698431365
transform 1 0 3762 0 1 4268
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_8
timestamp 1698431365
transform 1 0 3573 0 1 4484
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_9
timestamp 1698431365
transform 1 0 4166 0 1 4484
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_10
timestamp 1698431365
transform 1 0 4079 0 1 4700
box 0 0 1 1
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_0
timestamp 1698431365
transform 1 0 3619 0 1 1551
box 0 0 1 1
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_1
timestamp 1698431365
transform 1 0 4360 0 1 1539
box 0 0 1 1
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_2
timestamp 1698431365
transform 1 0 2959 0 1 1551
box 0 0 1 1
use M1_PSUB$$46554156_R90_256x8m81  M1_PSUB$$46554156_R90_256x8m81_0
timestamp 1698431365
transform 0 -1 2547 1 0 1031
box 0 0 1 1
use M1_PSUB$$46555180_256x8m81  M1_PSUB$$46555180_256x8m81_0
timestamp 1698431365
transform 1 0 3439 0 1 7080
box 0 0 1 1
use M1_PSUB$$46556204_256x8m81  M1_PSUB$$46556204_256x8m81_0
timestamp 1698431365
transform 1 0 1915 0 1 4550
box 0 0 1 1
use M1_PSUB$$46557228_256x8m81  M1_PSUB$$46557228_256x8m81_0
timestamp 1698431365
transform 1 0 2231 0 1 2020
box 0 0 1 1
use M1_PSUB$$46558252_256x8m81  M1_PSUB$$46558252_256x8m81_0
timestamp 1698431365
transform 1 0 3674 0 1 152
box 0 0 1 1
use M3_M2$$43371564_256x8m81  M3_M2$$43371564_256x8m81_0
timestamp 1698431365
transform 1 0 4337 0 1 3178
box 0 0 1 1
use M3_M2$$43371564_256x8m81  M3_M2$$43371564_256x8m81_1
timestamp 1698431365
transform 1 0 2528 0 1 3178
box 0 0 1 1
use nmos_1p2$$45107244_256x8m81  nmos_1p2$$45107244_256x8m81_0
timestamp 1698431365
transform -1 0 4243 0 -1 2156
box -31 0 -30 1
use nmos_1p2$$46550060_256x8m81  nmos_1p2$$46550060_256x8m81_0
timestamp 1698431365
transform 1 0 2620 0 1 2510
box -31 0 -30 1
use nmos_1p2$$46551084_256x8m81  nmos_1p2$$46551084_256x8m81_0
timestamp 1698431365
transform -1 0 3123 0 -1 2156
box -31 0 -30 1
use nmos_1p2$$46552108_256x8m81  nmos_1p2$$46552108_256x8m81_0
timestamp 1698431365
transform 1 0 2587 0 1 3317
box -31 0 -30 1
use nmos_1p2$$46553132_256x8m81  nmos_1p2$$46553132_256x8m81_0
timestamp 1698431365
transform 1 0 4379 0 1 3317
box -31 0 -30 1
use nmos_1p2$$46553132_256x8m81  nmos_1p2$$46553132_256x8m81_1
timestamp 1698431365
transform 1 0 2363 0 1 3317
box -31 0 -30 1
use pmos_1p2$$46285868_256x8m81  pmos_1p2$$46285868_256x8m81_0
timestamp 1698431365
transform 1 0 3406 0 1 5266
box -31 0 -30 1
use pmos_1p2$$46286892_256x8m81  pmos_1p2$$46286892_256x8m81_0
timestamp 1698431365
transform 1 0 3182 0 1 6132
box -31 0 -30 1
use pmos_1p2$$46549036_256x8m81  pmos_1p2$$46549036_256x8m81_0
timestamp 1698431365
transform -1 0 4243 0 -1 1331
box -31 0 -30 1
use pmos_1p2$$46896172_256x8m81  pmos_1p2$$46896172_256x8m81_0
timestamp 1698431365
transform 1 0 3052 0 1 4802
box -31 0 -30 1
use pmos_1p2$$46897196_256x8m81  pmos_1p2$$46897196_256x8m81_0
timestamp 1698431365
transform 1 0 2495 0 1 6132
box -31 0 -30 1
use pmos_1p2$$46897196_256x8m81  pmos_1p2$$46897196_256x8m81_1
timestamp 1698431365
transform 1 0 2495 0 1 5266
box -31 0 -30 1
use pmos_1p2$$46897196_256x8m81  pmos_1p2$$46897196_256x8m81_2
timestamp 1698431365
transform 1 0 4080 0 1 6132
box -31 0 -30 1
use pmos_1p2$$46897196_256x8m81  pmos_1p2$$46897196_256x8m81_3
timestamp 1698431365
transform 1 0 4080 0 1 5266
box -31 0 -30 1
use pmos_1p2$$46898220_256x8m81  pmos_1p2$$46898220_256x8m81_0
timestamp 1698431365
transform 1 0 2828 0 1 4802
box -31 0 -30 1
use pmos_1p2$$46898220_256x8m81  pmos_1p2$$46898220_256x8m81_1
timestamp 1698431365
transform 1 0 3948 0 1 4802
box -31 0 -30 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_0
timestamp 1698431365
transform 1 0 3386 0 1 2621
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_1
timestamp 1698431365
transform 1 0 4909 0 1 827
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_2
timestamp 1698431365
transform 1 0 3834 0 1 2621
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_3
timestamp 1698431365
transform -1 0 3700 0 -1 2201
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_4
timestamp 1698431365
transform -1 0 4146 0 -1 2201
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_5
timestamp 1698431365
transform 1 0 4271 0 1 2621
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_6
timestamp 1698431365
transform 1 0 2938 0 1 2621
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_7
timestamp 1698431365
transform -1 0 3033 0 -1 2029
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_8
timestamp 1698431365
transform 1 0 2523 0 1 827
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_9
timestamp 1698431365
transform 1 0 2523 0 1 1630
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_10
timestamp 1698431365
transform 1 0 2501 0 1 2621
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_11
timestamp 1698431365
transform 1 0 3050 0 1 6225
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_12
timestamp 1698431365
transform 1 0 2701 0 1 4665
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_13
timestamp 1698431365
transform 1 0 3151 0 1 4722
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_14
timestamp 1698431365
transform 1 0 2287 0 1 4722
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_15
timestamp 1698431365
transform 1 0 3623 0 1 4722
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_16
timestamp 1698431365
transform 1 0 3722 0 1 6225
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_17
timestamp 1698431365
transform 1 0 4040 0 1 4665
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_18
timestamp 1698431365
transform 1 0 4418 0 1 4722
box 0 0 1 1
use via1_2_x2_R90_256x8m81  via1_2_x2_R90_256x8m81_0
timestamp 1698431365
transform 0 -1 3259 1 0 7937
box 0 0 1 1
use via1_2_x2_R270_256x8m81  via1_2_x2_R270_256x8m81_0
timestamp 1698431365
transform 0 1 4262 -1 0 544
box 0 0 1 1
use via1_2_x2_R270_256x8m81  via1_2_x2_R270_256x8m81_1
timestamp 1698431365
transform 0 1 2723 -1 0 544
box 0 0 1 1
use via1_2_x2_R270_256x8m81  via1_2_x2_R270_256x8m81_2
timestamp 1698431365
transform 0 1 3182 -1 0 544
box 0 0 1 1
use via1_256x8m81  via1_256x8m81_0
timestamp 1698431365
transform 1 0 3388 0 -1 6790
box 0 0 1 1
use via1_R90_256x8m81  via1_R90_256x8m81_0
timestamp 1698431365
transform 0 -1 4506 1 0 3149
box 0 0 1 1
use via1_R90_256x8m81  via1_R90_256x8m81_1
timestamp 1698431365
transform 0 -1 2486 1 0 3149
box 0 0 1 1
use via1_R90_256x8m81  via1_R90_256x8m81_2
timestamp 1698431365
transform 0 -1 2520 1 0 4226
box 0 0 1 1
use via1_R90_256x8m81  via1_R90_256x8m81_3
timestamp 1698431365
transform 0 -1 4396 1 0 4437
box 0 0 1 1
use via1_R90_256x8m81  via1_R90_256x8m81_4
timestamp 1698431365
transform 0 -1 4568 1 0 4226
box 0 0 1 1
use via1_R90_256x8m81  via1_R90_256x8m81_5
timestamp 1698431365
transform 0 -1 3595 1 0 5792
box 0 0 1 1
use via1_R90_256x8m81  via1_R90_256x8m81_6
timestamp 1698431365
transform 0 1 3276 1 0 5964
box 0 0 1 1
use via1_R270_256x8m81  via1_R270_256x8m81_0
timestamp 1698431365
transform 0 -1 2925 -1 0 6762
box 0 0 1 1
use via1_R270_256x8m81  via1_R270_256x8m81_1
timestamp 1698431365
transform 0 1 3083 -1 0 4321
box 0 0 1 1
use via1_R270_256x8m81  via1_R270_256x8m81_2
timestamp 1698431365
transform 0 1 3193 -1 0 4532
box 0 0 1 1
use via1_R270_256x8m81  via1_R270_256x8m81_3
timestamp 1698431365
transform 0 -1 3500 -1 0 7361
box 0 0 1 1
use via1_R270_256x8m81  via1_R270_256x8m81_4
timestamp 1698431365
transform 0 -1 4060 -1 0 6740
box 0 0 1 1
use via1_R270_256x8m81  via1_R270_256x8m81_5
timestamp 1698431365
transform 0 1 3659 -1 0 4321
box 0 0 1 1
use via1_R270_256x8m81  via1_R270_256x8m81_6
timestamp 1698431365
transform 0 1 3371 -1 0 4321
box 0 0 1 1
use via1_R270_256x8m81  via1_R270_256x8m81_7
timestamp 1698431365
transform 0 1 3549 -1 0 4532
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_0
timestamp 1698431365
transform -1 0 4153 0 1 1018
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_1
timestamp 1698431365
transform 1 0 4276 0 1 1712
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_2
timestamp 1698431365
transform 1 0 3601 0 1 1018
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_3
timestamp 1698431365
transform -1 0 3920 0 1 1712
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_4
timestamp 1698431365
transform -1 0 3478 0 1 1712
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_5
timestamp 1698431365
transform 1 0 2596 0 1 6146
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_6
timestamp 1698431365
transform 1 0 4181 0 1 6146
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_7
timestamp 1698431365
transform 1 0 3503 0 1 6146
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_8
timestamp 1698431365
transform -1 0 3369 0 1 6146
box 0 0 1 1
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_0
timestamp 1698431365
transform 0 -1 4559 1 0 1494
box 0 0 1 1
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_1
timestamp 1698431365
transform 0 -1 3057 1 0 1505
box 0 0 1 1
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_2
timestamp 1698431365
transform 0 -1 2633 1 0 7937
box 0 0 1 1
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_3
timestamp 1698431365
transform 0 -1 3015 1 0 7728
box 0 0 1 1
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_4
timestamp 1698431365
transform 0 -1 3819 1 0 7728
box 0 0 1 1
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_5
timestamp 1698431365
transform 0 -1 4497 1 0 7937
box 0 0 1 1
use via1_x2_R270_256x8m81  via1_x2_R270_256x8m81_0
timestamp 1698431365
transform 0 1 2684 -1 0 4532
box 0 0 1 1
use via1_x2_R270_256x8m81  via1_x2_R270_256x8m81_1
timestamp 1698431365
transform 0 1 3883 -1 0 4532
box 0 0 1 1
use via2_x2_R90_256x8m81  via2_x2_R90_256x8m81_0
timestamp 1698431365
transform 0 -1 1992 1 0 7728
box 0 0 1 1
<< labels >>
rlabel metal1 s 3452 7551 3452 7551 4 wep
port 1 nsew
rlabel metal1 s 3437 7996 3437 7996 4 db
port 2 nsew
rlabel metal1 s 4471 2403 4471 2403 4 se
port 3 nsew
rlabel metal1 s 2040 7295 2040 7295 4 pcb
port 4 nsew
rlabel metal1 s 3432 7780 3432 7780 4 d
port 5 nsew
rlabel metal3 s 1179 5153 1179 5153 4 vdd
port 6 nsew
rlabel metal3 s 1247 2410 1247 2410 4 vss
port 7 nsew
rlabel metal3 s 1032 116 1032 116 4 vdd
port 6 nsew
rlabel metal2 s 3648 -136 3648 -136 4 qp
port 8 nsew
rlabel metal2 s 3995 7030 3995 7030 4 db
port 2 nsew
rlabel metal2 s 2868 7030 2868 7030 4 d
port 5 nsew
rlabel metal2 s 4111 -136 4111 -136 4 qn
port 9 nsew
<< properties >>
string GDS_END 476260
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 462254
<< end >>
