magic
tech gf180mcuD
magscale 1 10
timestamp 1698431365
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_0
timestamp 1698431365
transform -1 0 600 0 1 11700
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1
timestamp 1698431365
transform -1 0 600 0 1 4500
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_2
timestamp 1698431365
transform -1 0 600 0 1 8100
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_3
timestamp 1698431365
transform -1 0 600 0 1 15300
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_4
timestamp 1698431365
transform -1 0 600 0 1 9900
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_5
timestamp 1698431365
transform -1 0 600 0 1 13500
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_6
timestamp 1698431365
transform -1 0 600 0 1 2700
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_7
timestamp 1698431365
transform -1 0 600 0 1 6300
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_8
timestamp 1698431365
transform -1 0 600 0 1 900
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_9
timestamp 1698431365
transform -1 0 600 0 1 29700
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_10
timestamp 1698431365
transform -1 0 600 0 1 35100
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_11
timestamp 1698431365
transform -1 0 600 0 1 33300
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_12
timestamp 1698431365
transform -1 0 600 0 1 36900
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_13
timestamp 1698431365
transform -1 0 600 0 1 31500
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_14
timestamp 1698431365
transform -1 0 600 0 1 18900
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_15
timestamp 1698431365
transform -1 0 600 0 1 26100
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_16
timestamp 1698431365
transform -1 0 600 0 1 22500
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_17
timestamp 1698431365
transform -1 0 600 0 1 24300
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_18
timestamp 1698431365
transform -1 0 600 0 1 27900
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_19
timestamp 1698431365
transform -1 0 600 0 1 20700
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_20
timestamp 1698431365
transform -1 0 600 0 1 42300
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_21
timestamp 1698431365
transform -1 0 600 0 1 45900
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_22
timestamp 1698431365
transform -1 0 600 0 1 49500
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_23
timestamp 1698431365
transform -1 0 600 0 1 56700
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_24
timestamp 1698431365
transform -1 0 600 0 1 53100
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_25
timestamp 1698431365
transform -1 0 600 0 1 40500
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_26
timestamp 1698431365
transform -1 0 600 0 1 44100
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_27
timestamp 1698431365
transform -1 0 600 0 1 47700
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_28
timestamp 1698431365
transform -1 0 600 0 1 54900
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_29
timestamp 1698431365
transform -1 0 600 0 1 51300
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_30
timestamp 1698431365
transform -1 0 600 0 1 38700
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_31
timestamp 1698431365
transform -1 0 600 0 1 17100
box -68 -68 668 1868
use 018SRAM_cell1_512x8m81  018SRAM_cell1_512x8m81_0
timestamp 1698431365
transform -1 0 600 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_512x8m81  018SRAM_cell1_512x8m81_1
timestamp 1698431365
transform -1 0 600 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_0
timestamp 1698431365
transform -1 0 16800 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_1
timestamp 1698431365
transform -1 0 16200 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_2
timestamp 1698431365
transform -1 0 15600 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_3
timestamp 1698431365
transform -1 0 15000 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_4
timestamp 1698431365
transform -1 0 13800 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_5
timestamp 1698431365
transform -1 0 14400 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_6
timestamp 1698431365
transform -1 0 13200 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_7
timestamp 1698431365
transform -1 0 12600 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_8
timestamp 1698431365
transform -1 0 18000 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_9
timestamp 1698431365
transform -1 0 18600 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_10
timestamp 1698431365
transform -1 0 19800 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_11
timestamp 1698431365
transform -1 0 19200 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_12
timestamp 1698431365
transform -1 0 20400 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_13
timestamp 1698431365
transform -1 0 21000 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_14
timestamp 1698431365
transform -1 0 21600 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_15
timestamp 1698431365
transform -1 0 22200 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_16
timestamp 1698431365
transform -1 0 7800 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_17
timestamp 1698431365
transform -1 0 9000 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_18
timestamp 1698431365
transform -1 0 8400 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_19
timestamp 1698431365
transform -1 0 9600 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_20
timestamp 1698431365
transform -1 0 10200 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_21
timestamp 1698431365
transform -1 0 10800 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_22
timestamp 1698431365
transform -1 0 11400 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_23
timestamp 1698431365
transform -1 0 6000 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_24
timestamp 1698431365
transform -1 0 5400 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_25
timestamp 1698431365
transform -1 0 4800 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_26
timestamp 1698431365
transform -1 0 4200 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_27
timestamp 1698431365
transform -1 0 3000 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_28
timestamp 1698431365
transform -1 0 3600 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_29
timestamp 1698431365
transform -1 0 2400 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_30
timestamp 1698431365
transform -1 0 1800 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_31
timestamp 1698431365
transform -1 0 7200 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_32
timestamp 1698431365
transform -1 0 4200 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_33
timestamp 1698431365
transform -1 0 3000 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_34
timestamp 1698431365
transform -1 0 3600 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_35
timestamp 1698431365
transform -1 0 2400 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_36
timestamp 1698431365
transform -1 0 1800 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_37
timestamp 1698431365
transform -1 0 5400 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_38
timestamp 1698431365
transform -1 0 4800 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_39
timestamp 1698431365
transform -1 0 10800 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_40
timestamp 1698431365
transform -1 0 7200 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_41
timestamp 1698431365
transform -1 0 11400 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_42
timestamp 1698431365
transform -1 0 7800 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_43
timestamp 1698431365
transform -1 0 9000 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_44
timestamp 1698431365
transform -1 0 8400 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_45
timestamp 1698431365
transform -1 0 9600 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_46
timestamp 1698431365
transform -1 0 10200 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_47
timestamp 1698431365
transform -1 0 6000 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_48
timestamp 1698431365
transform -1 0 13800 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_49
timestamp 1698431365
transform -1 0 16200 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_50
timestamp 1698431365
transform -1 0 12600 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_51
timestamp 1698431365
transform -1 0 13200 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_52
timestamp 1698431365
transform -1 0 16800 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_53
timestamp 1698431365
transform -1 0 14400 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_54
timestamp 1698431365
transform -1 0 15000 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_55
timestamp 1698431365
transform -1 0 15600 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_56
timestamp 1698431365
transform -1 0 19200 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_57
timestamp 1698431365
transform -1 0 18600 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_58
timestamp 1698431365
transform -1 0 21000 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_59
timestamp 1698431365
transform -1 0 20400 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_60
timestamp 1698431365
transform -1 0 21600 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_61
timestamp 1698431365
transform -1 0 19800 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_62
timestamp 1698431365
transform -1 0 22200 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_63
timestamp 1698431365
transform -1 0 18000 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_0
timestamp 1698431365
transform 1 0 22800 0 -1 7200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_1
timestamp 1698431365
transform 1 0 22800 0 -1 9000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_2
timestamp 1698431365
transform 1 0 22800 0 -1 5400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_3
timestamp 1698431365
transform 1 0 22800 0 -1 3600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_4
timestamp 1698431365
transform 1 0 22800 0 -1 10800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_5
timestamp 1698431365
transform 1 0 22800 0 -1 18000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_6
timestamp 1698431365
transform 1 0 22800 0 -1 16200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_7
timestamp 1698431365
transform 1 0 22800 0 -1 14400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_8
timestamp 1698431365
transform 1 0 22800 0 -1 12600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_9
timestamp 1698431365
transform 1 0 22800 0 -1 1800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_10
timestamp 1698431365
transform 1 0 22800 0 1 5400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_11
timestamp 1698431365
transform 1 0 22800 0 1 7200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_12
timestamp 1698431365
transform 1 0 22800 0 1 10800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_13
timestamp 1698431365
transform 1 0 22800 0 1 14400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_14
timestamp 1698431365
transform 1 0 22800 0 1 3600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_15
timestamp 1698431365
transform 1 0 22800 0 1 9000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_16
timestamp 1698431365
transform 1 0 22800 0 1 12600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_17
timestamp 1698431365
transform 1 0 22800 0 1 16200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_18
timestamp 1698431365
transform 1 0 22800 0 1 1800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_19
timestamp 1698431365
transform 1 0 22800 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_20
timestamp 1698431365
transform 1 0 22800 0 -1 37800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_21
timestamp 1698431365
transform 1 0 22800 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_22
timestamp 1698431365
transform 1 0 22800 0 -1 36000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_23
timestamp 1698431365
transform 1 0 22800 0 -1 34200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_24
timestamp 1698431365
transform 1 0 22800 0 -1 32400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_25
timestamp 1698431365
transform 1 0 22800 0 -1 23400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_26
timestamp 1698431365
transform 1 0 22800 0 -1 19800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_27
timestamp 1698431365
transform 1 0 22800 0 -1 21600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_28
timestamp 1698431365
transform 1 0 22800 0 -1 28800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_29
timestamp 1698431365
transform 1 0 22800 0 -1 27000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_30
timestamp 1698431365
transform 1 0 22800 0 -1 25200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_31
timestamp 1698431365
transform 1 0 22800 0 1 36000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_32
timestamp 1698431365
transform 1 0 22800 0 1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_33
timestamp 1698431365
transform 1 0 22800 0 1 21600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_34
timestamp 1698431365
transform 1 0 22800 0 1 25200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_35
timestamp 1698431365
transform 1 0 22800 0 1 28800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_36
timestamp 1698431365
transform 1 0 22800 0 1 32400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_37
timestamp 1698431365
transform 1 0 22800 0 1 34200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_38
timestamp 1698431365
transform 1 0 22800 0 1 19800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_39
timestamp 1698431365
transform 1 0 22800 0 1 23400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_40
timestamp 1698431365
transform 1 0 22800 0 1 27000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_41
timestamp 1698431365
transform 1 0 22800 0 1 37800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_42
timestamp 1698431365
transform 1 0 22800 0 -1 55800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_43
timestamp 1698431365
transform 1 0 22800 0 -1 52200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_44
timestamp 1698431365
transform 1 0 22800 0 -1 48600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_45
timestamp 1698431365
transform 1 0 22800 0 -1 43200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_46
timestamp 1698431365
transform 1 0 22800 0 -1 41400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_47
timestamp 1698431365
transform 1 0 22800 0 -1 57600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_48
timestamp 1698431365
transform 1 0 22800 0 -1 54000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_49
timestamp 1698431365
transform 1 0 22800 0 -1 50400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_50
timestamp 1698431365
transform 1 0 22800 0 -1 46800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_51
timestamp 1698431365
transform 1 0 22800 0 -1 45000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_52
timestamp 1698431365
transform 1 0 22800 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_53
timestamp 1698431365
transform 1 0 22800 0 1 54000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_54
timestamp 1698431365
transform 1 0 22800 0 1 39600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_55
timestamp 1698431365
transform 1 0 22800 0 1 46800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_56
timestamp 1698431365
transform 1 0 22800 0 1 55800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_57
timestamp 1698431365
transform 1 0 22800 0 1 50400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_58
timestamp 1698431365
transform 1 0 22800 0 1 43200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_59
timestamp 1698431365
transform 1 0 22800 0 1 57600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_60
timestamp 1698431365
transform 1 0 22800 0 1 45000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_61
timestamp 1698431365
transform 1 0 22800 0 1 52200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_62
timestamp 1698431365
transform 1 0 22800 0 1 41400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_63
timestamp 1698431365
transform 1 0 22800 0 1 48600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_64
timestamp 1698431365
transform 1 0 22800 0 -1 39600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_65
timestamp 1698431365
transform 1 0 22800 0 1 18000
box -68 -68 668 968
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_0
timestamp 1698431365
transform -1 0 17400 0 1 0
box -68 -68 668 968
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_1
timestamp 1698431365
transform -1 0 6600 0 1 0
box -68 -68 668 968
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_2
timestamp 1698431365
transform -1 0 1200 0 1 0
box -68 -68 668 968
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_3
timestamp 1698431365
transform -1 0 6600 0 -1 59400
box -68 -68 668 968
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_4
timestamp 1698431365
transform -1 0 17400 0 -1 59400
box -68 -68 668 968
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_5
timestamp 1698431365
transform 1 0 22200 0 -1 59400
box -68 -68 668 968
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_6
timestamp 1698431365
transform -1 0 12000 0 1 0
box -68 -68 668 968
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_7
timestamp 1698431365
transform -1 0 12000 0 -1 59400
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_0
timestamp 1698431365
transform 1 0 22200 0 1 0
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_1
timestamp 1698431365
transform -1 0 1200 0 -1 3600
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_2
timestamp 1698431365
transform -1 0 1200 0 -1 5400
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_3
timestamp 1698431365
transform -1 0 1200 0 1 1800
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_4
timestamp 1698431365
transform -1 0 1200 0 1 3600
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_5
timestamp 1698431365
transform -1 0 1200 0 -1 16200
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_6
timestamp 1698431365
transform -1 0 1200 0 1 5400
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_7
timestamp 1698431365
transform -1 0 1200 0 1 9000
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_8
timestamp 1698431365
transform -1 0 1200 0 1 7200
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_9
timestamp 1698431365
transform -1 0 1200 0 1 10800
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_10
timestamp 1698431365
transform -1 0 1200 0 1 12600
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_11
timestamp 1698431365
transform -1 0 1200 0 -1 1800
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_12
timestamp 1698431365
transform -1 0 1200 0 -1 14400
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_13
timestamp 1698431365
transform -1 0 1200 0 -1 18000
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_14
timestamp 1698431365
transform -1 0 1200 0 -1 7200
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_15
timestamp 1698431365
transform -1 0 1200 0 -1 10800
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_16
timestamp 1698431365
transform -1 0 1200 0 1 14400
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_17
timestamp 1698431365
transform -1 0 1200 0 -1 12600
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_18
timestamp 1698431365
transform -1 0 1200 0 -1 9000
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_19
timestamp 1698431365
transform -1 0 1200 0 1 16200
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_20
timestamp 1698431365
transform -1 0 1200 0 1 34200
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_21
timestamp 1698431365
transform -1 0 1200 0 1 36000
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_22
timestamp 1698431365
transform -1 0 1200 0 1 37800
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_23
timestamp 1698431365
transform -1 0 1200 0 -1 23400
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_24
timestamp 1698431365
transform -1 0 1200 0 -1 30600
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_25
timestamp 1698431365
transform -1 0 1200 0 -1 36000
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_26
timestamp 1698431365
transform -1 0 1200 0 -1 27000
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_27
timestamp 1698431365
transform -1 0 1200 0 1 30600
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_28
timestamp 1698431365
transform -1 0 1200 0 -1 28800
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_29
timestamp 1698431365
transform -1 0 1200 0 -1 34200
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_30
timestamp 1698431365
transform -1 0 1200 0 -1 32400
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_31
timestamp 1698431365
transform -1 0 1200 0 1 27000
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_32
timestamp 1698431365
transform -1 0 1200 0 -1 37800
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_33
timestamp 1698431365
transform -1 0 1200 0 1 28800
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_34
timestamp 1698431365
transform -1 0 1200 0 -1 19800
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_35
timestamp 1698431365
transform -1 0 1200 0 1 23400
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_36
timestamp 1698431365
transform -1 0 1200 0 1 25200
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_37
timestamp 1698431365
transform -1 0 1200 0 1 21600
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_38
timestamp 1698431365
transform -1 0 1200 0 1 19800
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_39
timestamp 1698431365
transform -1 0 1200 0 -1 25200
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_40
timestamp 1698431365
transform -1 0 1200 0 1 32400
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_41
timestamp 1698431365
transform -1 0 1200 0 -1 21600
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_42
timestamp 1698431365
transform -1 0 1200 0 -1 50400
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_43
timestamp 1698431365
transform -1 0 1200 0 1 57600
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_44
timestamp 1698431365
transform -1 0 1200 0 1 54000
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_45
timestamp 1698431365
transform -1 0 1200 0 1 46800
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_46
timestamp 1698431365
transform -1 0 1200 0 1 41400
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_47
timestamp 1698431365
transform -1 0 1200 0 1 39600
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_48
timestamp 1698431365
transform -1 0 1200 0 1 43200
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_49
timestamp 1698431365
transform -1 0 1200 0 1 45000
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_50
timestamp 1698431365
transform -1 0 1200 0 1 55800
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_51
timestamp 1698431365
transform -1 0 1200 0 1 52200
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_52
timestamp 1698431365
transform -1 0 1200 0 1 50400
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_53
timestamp 1698431365
transform -1 0 1200 0 1 48600
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_54
timestamp 1698431365
transform -1 0 1200 0 -1 59400
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_55
timestamp 1698431365
transform -1 0 1200 0 -1 46800
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_56
timestamp 1698431365
transform -1 0 1200 0 -1 57600
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_57
timestamp 1698431365
transform -1 0 1200 0 -1 45000
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_58
timestamp 1698431365
transform -1 0 1200 0 -1 52200
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_59
timestamp 1698431365
transform -1 0 1200 0 -1 48600
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_60
timestamp 1698431365
transform -1 0 1200 0 -1 54000
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_61
timestamp 1698431365
transform -1 0 1200 0 -1 41400
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_62
timestamp 1698431365
transform -1 0 1200 0 -1 43200
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_63
timestamp 1698431365
transform -1 0 1200 0 -1 55800
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_64
timestamp 1698431365
transform -1 0 1200 0 -1 39600
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_65
timestamp 1698431365
transform -1 0 1200 0 1 18000
box -68 -68 668 968
use M1_NWELL$$44998700_512x8m81  M1_NWELL$$44998700_512x8m81_0
timestamp 1698431365
transform 1 0 23318 0 1 -22942
box 0 0 1 1
use M1_NWELL$$44998700_512x8m81  M1_NWELL$$44998700_512x8m81_1
timestamp 1698431365
transform 1 0 22774 0 1 -22942
box 0 0 1 1
use M1_NWELL$$46277676_512x8m81  M1_NWELL$$46277676_512x8m81_0
timestamp 1698431365
transform 1 0 23050 0 1 -14622
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_0
timestamp 1698431365
transform 1 0 23615 0 -1 7200
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_1
timestamp 1698431365
transform 1 0 23615 0 -1 5400
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_2
timestamp 1698431365
transform 1 0 23615 0 -1 1800
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_3
timestamp 1698431365
transform 1 0 23615 0 -1 240
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_4
timestamp 1698431365
transform 1 0 23615 0 -1 16200
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_5
timestamp 1698431365
transform 1 0 23615 0 -1 12600
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_6
timestamp 1698431365
transform 1 0 23615 0 -1 9000
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_7
timestamp 1698431365
transform 1 0 23615 0 -1 14400
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_8
timestamp 1698431365
transform 1 0 23615 0 -1 10800
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_9
timestamp 1698431365
transform 1 0 23615 0 -1 3600
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_10
timestamp 1698431365
transform 1 0 23615 0 -1 21600
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_11
timestamp 1698431365
transform 1 0 23615 0 -1 37800
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_12
timestamp 1698431365
transform 1 0 23615 0 -1 36000
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_13
timestamp 1698431365
transform 1 0 23615 0 -1 34200
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_14
timestamp 1698431365
transform 1 0 23615 0 -1 32400
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_15
timestamp 1698431365
transform 1 0 23615 0 -1 30600
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_16
timestamp 1698431365
transform 1 0 23615 0 -1 27000
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_17
timestamp 1698431365
transform 1 0 23615 0 -1 23400
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_18
timestamp 1698431365
transform 1 0 23615 0 -1 19800
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_19
timestamp 1698431365
transform 1 0 23615 0 -1 28800
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_20
timestamp 1698431365
transform 1 0 23615 0 -1 25200
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_21
timestamp 1698431365
transform 1 0 23615 0 -1 55800
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_22
timestamp 1698431365
transform 1 0 23615 0 -1 54000
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_23
timestamp 1698431365
transform 1 0 23615 0 -1 52200
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_24
timestamp 1698431365
transform 1 0 23615 0 -1 50400
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_25
timestamp 1698431365
transform 1 0 23615 0 -1 48600
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_26
timestamp 1698431365
transform 1 0 23615 0 -1 46800
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_27
timestamp 1698431365
transform 1 0 23615 0 -1 45000
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_28
timestamp 1698431365
transform 1 0 23615 0 -1 43200
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_29
timestamp 1698431365
transform 1 0 23615 0 -1 41400
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_30
timestamp 1698431365
transform 1 0 23615 0 -1 39600
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_31
timestamp 1698431365
transform 1 0 23615 0 -1 57600
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_32
timestamp 1698431365
transform 1 0 23615 0 -1 59160
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_33
timestamp 1698431365
transform 1 0 23615 0 -1 18000
box 0 0 1 1
use M1_POLY2$$46559276_512x8m81_0  M1_POLY2$$46559276_512x8m81_0_0
timestamp 1698431365
transform -1 0 22809 0 1 -19544
box 0 0 1 1
use M1_POLY2$$46559276_512x8m81_0  M1_POLY2$$46559276_512x8m81_0_1
timestamp 1698431365
transform 1 0 23393 0 1 -15883
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_0
timestamp 1698431365
transform 1 0 -215 0 1 141
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_1
timestamp 1698431365
transform 1 0 -215 0 1 1800
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_2
timestamp 1698431365
transform 1 0 -215 0 1 3600
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_3
timestamp 1698431365
transform 1 0 -215 0 1 7200
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_4
timestamp 1698431365
transform 1 0 -215 0 1 5400
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_5
timestamp 1698431365
transform 1 0 -215 0 1 14400
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_6
timestamp 1698431365
transform 1 0 -215 0 1 12600
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_7
timestamp 1698431365
transform 1 0 -215 0 1 16200
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_8
timestamp 1698431365
transform 1 0 -215 0 1 18000
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_9
timestamp 1698431365
transform 1 0 -215 0 1 10800
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_10
timestamp 1698431365
transform 1 0 -215 0 1 9000
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_11
timestamp 1698431365
transform 1 0 -215 0 1 21600
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_12
timestamp 1698431365
transform 1 0 -215 0 1 19800
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_13
timestamp 1698431365
transform 1 0 -215 0 1 23400
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_14
timestamp 1698431365
transform 1 0 -215 0 1 25200
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_15
timestamp 1698431365
transform 1 0 -215 0 1 28800
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_16
timestamp 1698431365
transform 1 0 -215 0 1 27000
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_17
timestamp 1698431365
transform 1 0 -215 0 1 30600
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_18
timestamp 1698431365
transform 1 0 -215 0 1 32400
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_19
timestamp 1698431365
transform 1 0 -215 0 1 36000
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_20
timestamp 1698431365
transform 1 0 -215 0 1 34200
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_21
timestamp 1698431365
transform 1 0 -215 0 1 37800
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_22
timestamp 1698431365
transform 1 0 -215 0 1 39600
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_23
timestamp 1698431365
transform 1 0 -215 0 1 43200
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_24
timestamp 1698431365
transform 1 0 -215 0 1 41400
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_25
timestamp 1698431365
transform 1 0 -215 0 1 45000
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_26
timestamp 1698431365
transform 1 0 -215 0 1 46800
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_27
timestamp 1698431365
transform 1 0 -215 0 1 50400
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_28
timestamp 1698431365
transform 1 0 -215 0 1 48600
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_29
timestamp 1698431365
transform 1 0 -215 0 1 52200
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_30
timestamp 1698431365
transform 1 0 -215 0 1 54000
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_31
timestamp 1698431365
transform 1 0 -215 0 1 57600
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_32
timestamp 1698431365
transform 1 0 -215 0 1 55800
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_33
timestamp 1698431365
transform 1 0 -215 0 1 59259
box 0 0 1 1
use M1_PSUB$$46274604_512x8m81  M1_PSUB$$46274604_512x8m81_0
timestamp 1698431365
transform 1 0 23107 0 1 -16617
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_0
timestamp 1698431365
transform 1 0 23613 0 -1 16198
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_1
timestamp 1698431365
transform 1 0 23613 0 -1 12598
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_2
timestamp 1698431365
transform 1 0 23613 0 -1 8998
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_3
timestamp 1698431365
transform 1 0 23613 0 -1 5398
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_4
timestamp 1698431365
transform 1 0 23613 0 -1 1798
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_5
timestamp 1698431365
transform 1 0 23613 0 -1 10802
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_6
timestamp 1698431365
transform 1 0 23613 0 -1 3602
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_7
timestamp 1698431365
transform 1 0 23613 0 -1 265
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_8
timestamp 1698431365
transform 1 0 23613 0 -1 14402
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_9
timestamp 1698431365
transform 1 0 23613 0 -1 7202
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_10
timestamp 1698431365
transform 1 0 23613 0 -1 32398
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_11
timestamp 1698431365
transform 1 0 23613 0 -1 30598
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_12
timestamp 1698431365
transform 1 0 23613 0 -1 26998
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_13
timestamp 1698431365
transform 1 0 23613 0 -1 23398
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_14
timestamp 1698431365
transform 1 0 23613 0 -1 19798
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_15
timestamp 1698431365
transform 1 0 23613 0 -1 25202
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_16
timestamp 1698431365
transform 1 0 23613 0 -1 28798
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_17
timestamp 1698431365
transform 1 0 23613 0 -1 37798
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_18
timestamp 1698431365
transform 1 0 23613 0 -1 21602
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_19
timestamp 1698431365
transform 1 0 23613 0 -1 35998
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_20
timestamp 1698431365
transform 1 0 23613 0 -1 34198
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_21
timestamp 1698431365
transform 1 0 23613 0 -1 55798
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_22
timestamp 1698431365
transform 1 0 23613 0 -1 53998
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_23
timestamp 1698431365
transform 1 0 23613 0 -1 52198
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_24
timestamp 1698431365
transform 1 0 23613 0 -1 50398
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_25
timestamp 1698431365
transform 1 0 23613 0 -1 48598
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_26
timestamp 1698431365
transform 1 0 23613 0 -1 46798
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_27
timestamp 1698431365
transform 1 0 23613 0 -1 44998
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_28
timestamp 1698431365
transform 1 0 23613 0 -1 43198
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_29
timestamp 1698431365
transform 1 0 23613 0 -1 41398
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_30
timestamp 1698431365
transform 1 0 23613 0 -1 39598
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_31
timestamp 1698431365
transform 1 0 23613 0 -1 59135
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_32
timestamp 1698431365
transform 1 0 23613 0 -1 57598
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_33
timestamp 1698431365
transform 1 0 23613 0 -1 18002
box 0 0 1 1
use M2_M1$$47117356_512x8m81  M2_M1$$47117356_512x8m81_0
timestamp 1698431365
transform 1 0 23114 0 1 -20269
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_0
timestamp 1698431365
transform 1 0 -215 0 1 1800
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_1
timestamp 1698431365
transform 1 0 -215 0 1 3600
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_2
timestamp 1698431365
transform 1 0 -215 0 1 5400
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_3
timestamp 1698431365
transform 1 0 -215 0 1 7200
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_4
timestamp 1698431365
transform 1 0 -215 0 1 9000
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_5
timestamp 1698431365
transform 1 0 -215 0 1 10800
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_6
timestamp 1698431365
transform 1 0 -215 0 1 12600
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_7
timestamp 1698431365
transform 1 0 -215 0 1 14400
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_8
timestamp 1698431365
transform 1 0 -215 0 1 16200
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_9
timestamp 1698431365
transform 1 0 -215 0 1 18000
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_10
timestamp 1698431365
transform 1 0 -215 0 1 37800
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_11
timestamp 1698431365
transform 1 0 -215 0 1 36000
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_12
timestamp 1698431365
transform 1 0 -215 0 1 34200
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_13
timestamp 1698431365
transform 1 0 -215 0 1 32400
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_14
timestamp 1698431365
transform 1 0 -215 0 1 30600
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_15
timestamp 1698431365
transform 1 0 -215 0 1 28800
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_16
timestamp 1698431365
transform 1 0 -215 0 1 27000
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_17
timestamp 1698431365
transform 1 0 -215 0 1 25200
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_18
timestamp 1698431365
transform 1 0 -215 0 1 19800
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_19
timestamp 1698431365
transform 1 0 -215 0 1 21600
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_20
timestamp 1698431365
transform 1 0 -219 0 1 23400
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_21
timestamp 1698431365
transform 1 0 -215 0 1 57599
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_22
timestamp 1698431365
transform 1 0 -215 0 1 55800
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_23
timestamp 1698431365
transform 1 0 -215 0 1 54000
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_24
timestamp 1698431365
transform 1 0 -215 0 1 52200
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_25
timestamp 1698431365
transform 1 0 -215 0 1 50399
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_26
timestamp 1698431365
transform 1 0 -215 0 1 48600
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_27
timestamp 1698431365
transform 1 0 -215 0 1 46801
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_28
timestamp 1698431365
transform 1 0 -215 0 1 45000
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_29
timestamp 1698431365
transform 1 0 -215 0 1 43200
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_30
timestamp 1698431365
transform 1 0 -215 0 1 41400
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_31
timestamp 1698431365
transform 1 0 -215 0 1 39600
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_32
timestamp 1698431365
transform 1 0 -215 0 1 59198
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_0
timestamp 1698431365
transform 0 -1 -216 1 0 -4
box 0 0 1 1
use nmos_5p04310591302096_512x8m81  nmos_5p04310591302096_512x8m81_0
timestamp 1698431365
transform 1 0 22940 0 1 -19403
box 0 0 1 1
use nmos_5p04310591302098_512x8m81  nmos_5p04310591302098_512x8m81_0
timestamp 1698431365
transform 1 0 22936 0 1 -16318
box 0 0 1 1
use pmos_5p04310591302095_512x8m81  pmos_5p04310591302095_512x8m81_0
timestamp 1698431365
transform 1 0 22936 0 1 -15738
box 0 0 1 1
use pmos_5p04310591302097_512x8m81  pmos_5p04310591302097_512x8m81_0
timestamp 1698431365
transform 1 0 22940 0 -1 -19684
box 0 0 1 1
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_0
timestamp 1698431365
transform 1 0 23283 0 1 -18447
box 0 0 1 1
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_1
timestamp 1698431365
transform 1 0 23285 0 1 -15470
box 0 0 1 1
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_2
timestamp 1698431365
transform 1 0 23288 0 1 -22897
box 0 0 1 1
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_3
timestamp 1698431365
transform 1 0 22846 0 1 -22711
box 0 0 1 1
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_4
timestamp 1698431365
transform 1 0 22842 0 1 -17909
box 0 0 1 1
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_5
timestamp 1698431365
transform 1 0 22842 0 1 -19052
box 0 0 1 1
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_6
timestamp 1698431365
transform 1 0 22837 0 1 -15470
box 0 0 1 1
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_7
timestamp 1698431365
transform 1 0 23288 0 1 -22711
box 0 0 1 1
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_8
timestamp 1698431365
transform 1 0 22842 0 1 -18447
box 0 0 1 1
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_9
timestamp 1698431365
transform 1 0 22846 0 1 -22897
box 0 0 1 1
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_10
timestamp 1698431365
transform 1 0 23283 0 1 -17909
box 0 0 1 1
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_11
timestamp 1698431365
transform 1 0 23283 0 1 -19052
box 0 0 1 1
use via1_2_x2_R90_512x8m81_0  via1_2_x2_R90_512x8m81_0_0
timestamp 1698431365
transform 0 -1 23187 1 0 -14670
box 0 0 1 1
use via1_2_x2_R270_512x8m81_0  via1_2_x2_R270_512x8m81_0_0
timestamp 1698431365
transform 0 1 22794 -1 0 -12002
box 0 0 1 1
use ypass_gate_512x8m81_0  ypass_gate_512x8m81_0_0
timestamp 1698431365
transform -1 0 23395 0 1 -13448
box -154 88 521 12143
<< properties >>
string GDS_END 2520180
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 2481608
<< end >>
