magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 377 6022 870
rect -86 352 1193 377
rect 4269 352 6022 377
<< pwell >>
rect 1193 352 4269 377
rect -86 -86 6022 352
<< mvnmos >>
rect 124 156 244 232
rect 348 156 468 232
rect 516 156 636 232
rect 740 156 860 232
rect 908 156 1028 232
rect 1432 144 1552 237
rect 1750 144 1870 237
rect 2208 124 2328 219
rect 2432 124 2552 219
rect 2600 124 2720 219
rect 2900 185 3020 257
rect 3068 185 3188 257
rect 3292 185 3412 257
rect 3516 185 3636 257
rect 4029 158 4149 232
rect 4197 158 4317 232
rect 4465 69 4585 232
rect 4689 69 4809 232
rect 4913 69 5033 232
rect 5137 69 5257 232
rect 5361 69 5481 232
rect 5585 69 5705 232
<< mvpmos >>
rect 124 556 224 628
rect 348 556 448 628
rect 496 556 596 628
rect 740 556 840 628
rect 888 556 988 628
rect 1432 497 1532 660
rect 1750 497 1850 660
rect 2188 518 2288 590
rect 2392 518 2492 590
rect 2540 518 2640 590
rect 2864 497 2964 660
rect 3068 497 3168 660
rect 3520 497 3620 580
rect 3724 497 3824 580
rect 4072 497 4172 591
rect 4276 497 4376 591
rect 4532 472 4632 716
rect 4736 472 4836 716
rect 4940 472 5040 716
rect 5147 472 5247 716
rect 5353 472 5453 716
rect 5585 472 5685 716
<< mvndiff >>
rect 1300 244 1372 257
rect 36 219 124 232
rect 36 173 49 219
rect 95 173 124 219
rect 36 156 124 173
rect 244 215 348 232
rect 244 169 273 215
rect 319 169 348 215
rect 244 156 348 169
rect 468 156 516 232
rect 636 219 740 232
rect 636 173 665 219
rect 711 173 740 219
rect 636 156 740 173
rect 860 156 908 232
rect 1028 156 1160 232
rect 1088 95 1160 156
rect 1300 198 1313 244
rect 1359 237 1372 244
rect 1940 244 2012 257
rect 1940 237 1953 244
rect 1359 198 1432 237
rect 1300 144 1432 198
rect 1552 144 1750 237
rect 1870 198 1953 237
rect 1999 198 2012 244
rect 2780 219 2900 257
rect 1870 144 2012 198
rect 2120 183 2208 219
rect 1088 49 1101 95
rect 1147 49 1160 95
rect 1088 36 1160 49
rect 1612 95 1684 144
rect 1612 49 1625 95
rect 1671 49 1684 95
rect 1612 36 1684 49
rect 2120 137 2133 183
rect 2179 137 2208 183
rect 2120 124 2208 137
rect 2328 193 2432 219
rect 2328 147 2357 193
rect 2403 147 2432 193
rect 2328 124 2432 147
rect 2552 124 2600 219
rect 2720 185 2900 219
rect 3020 185 3068 257
rect 3188 244 3292 257
rect 3188 198 3217 244
rect 3263 198 3292 244
rect 3188 185 3292 198
rect 3412 244 3516 257
rect 3412 198 3441 244
rect 3487 198 3516 244
rect 3412 185 3516 198
rect 3636 244 3724 257
rect 3636 198 3665 244
rect 3711 198 3724 244
rect 3636 185 3724 198
rect 2720 183 2840 185
rect 2720 137 2781 183
rect 2827 137 2840 183
rect 2720 124 2840 137
rect 3884 244 3956 257
rect 3884 198 3897 244
rect 3943 232 3956 244
rect 3943 198 4029 232
rect 3884 158 4029 198
rect 4149 158 4197 232
rect 4317 193 4465 232
rect 4317 158 4390 193
rect 4377 147 4390 158
rect 4436 147 4465 193
rect 4377 69 4465 147
rect 4585 218 4689 232
rect 4585 172 4614 218
rect 4660 172 4689 218
rect 4585 69 4689 172
rect 4809 218 4913 232
rect 4809 172 4838 218
rect 4884 172 4913 218
rect 4809 69 4913 172
rect 5033 218 5137 232
rect 5033 172 5062 218
rect 5108 172 5137 218
rect 5033 69 5137 172
rect 5257 149 5361 232
rect 5257 103 5286 149
rect 5332 103 5361 149
rect 5257 69 5361 103
rect 5481 218 5585 232
rect 5481 172 5510 218
rect 5556 172 5585 218
rect 5481 69 5585 172
rect 5705 218 5793 232
rect 5705 172 5734 218
rect 5780 172 5793 218
rect 5705 69 5793 172
<< mvpdiff >>
rect 1048 707 1120 720
rect 1048 661 1061 707
rect 1107 661 1120 707
rect 1048 628 1120 661
rect 1618 716 1690 729
rect 1618 670 1631 716
rect 1677 670 1690 716
rect 1618 660 1690 670
rect 36 615 124 628
rect 36 569 49 615
rect 95 569 124 615
rect 36 556 124 569
rect 224 615 348 628
rect 224 569 263 615
rect 309 569 348 615
rect 224 556 348 569
rect 448 556 496 628
rect 596 615 740 628
rect 596 569 665 615
rect 711 569 740 615
rect 596 556 740 569
rect 840 556 888 628
rect 988 556 1120 628
rect 1344 556 1432 660
rect 1344 510 1357 556
rect 1403 510 1432 556
rect 1344 497 1432 510
rect 1532 497 1750 660
rect 1850 556 1938 660
rect 2700 718 2772 731
rect 2700 672 2713 718
rect 2759 672 2772 718
rect 2700 660 2772 672
rect 2700 590 2864 660
rect 1850 510 1879 556
rect 1925 510 1938 556
rect 2100 577 2188 590
rect 2100 531 2113 577
rect 2159 531 2188 577
rect 2100 518 2188 531
rect 2288 577 2392 590
rect 2288 531 2317 577
rect 2363 531 2392 577
rect 2288 518 2392 531
rect 2492 518 2540 590
rect 2640 518 2864 590
rect 1850 497 1938 510
rect 2700 497 2864 518
rect 2964 556 3068 660
rect 2964 510 2993 556
rect 3039 510 3068 556
rect 2964 497 3068 510
rect 3168 647 3256 660
rect 3168 601 3197 647
rect 3243 601 3256 647
rect 3168 497 3256 601
rect 4444 665 4532 716
rect 4444 591 4457 665
rect 3432 562 3520 580
rect 3432 516 3445 562
rect 3491 516 3520 562
rect 3432 497 3520 516
rect 3620 562 3724 580
rect 3620 516 3649 562
rect 3695 516 3724 562
rect 3620 497 3724 516
rect 3824 562 3912 580
rect 3824 516 3853 562
rect 3899 516 3912 562
rect 3824 497 3912 516
rect 3984 578 4072 591
rect 3984 532 3997 578
rect 4043 532 4072 578
rect 3984 497 4072 532
rect 4172 556 4276 591
rect 4172 510 4201 556
rect 4247 510 4276 556
rect 4172 497 4276 510
rect 4376 525 4457 591
rect 4503 525 4532 665
rect 4376 497 4532 525
rect 4436 472 4532 497
rect 4632 665 4736 716
rect 4632 525 4661 665
rect 4707 525 4736 665
rect 4632 472 4736 525
rect 4836 665 4940 716
rect 4836 525 4865 665
rect 4911 525 4940 665
rect 4836 472 4940 525
rect 5040 665 5147 716
rect 5040 525 5072 665
rect 5118 525 5147 665
rect 5040 472 5147 525
rect 5247 665 5353 716
rect 5247 525 5276 665
rect 5322 525 5353 665
rect 5247 472 5353 525
rect 5453 665 5585 716
rect 5453 525 5495 665
rect 5541 525 5585 665
rect 5453 472 5585 525
rect 5685 665 5773 716
rect 5685 525 5714 665
rect 5760 525 5773 665
rect 5685 472 5773 525
<< mvndiffc >>
rect 49 173 95 219
rect 273 169 319 215
rect 665 173 711 219
rect 1313 198 1359 244
rect 1953 198 1999 244
rect 1101 49 1147 95
rect 1625 49 1671 95
rect 2133 137 2179 183
rect 2357 147 2403 193
rect 3217 198 3263 244
rect 3441 198 3487 244
rect 3665 198 3711 244
rect 2781 137 2827 183
rect 3897 198 3943 244
rect 4390 147 4436 193
rect 4614 172 4660 218
rect 4838 172 4884 218
rect 5062 172 5108 218
rect 5286 103 5332 149
rect 5510 172 5556 218
rect 5734 172 5780 218
<< mvpdiffc >>
rect 1061 661 1107 707
rect 1631 670 1677 716
rect 49 569 95 615
rect 263 569 309 615
rect 665 569 711 615
rect 1357 510 1403 556
rect 2713 672 2759 718
rect 1879 510 1925 556
rect 2113 531 2159 577
rect 2317 531 2363 577
rect 2993 510 3039 556
rect 3197 601 3243 647
rect 3445 516 3491 562
rect 3649 516 3695 562
rect 3853 516 3899 562
rect 3997 532 4043 578
rect 4201 510 4247 556
rect 4457 525 4503 665
rect 4661 525 4707 665
rect 4865 525 4911 665
rect 5072 525 5118 665
rect 5276 525 5322 665
rect 5495 525 5541 665
rect 5714 525 5760 665
<< polysilicon >>
rect 124 720 988 760
rect 124 628 224 720
rect 348 628 448 672
rect 496 628 596 672
rect 740 628 840 672
rect 888 628 988 720
rect 1432 660 1532 717
rect 1750 720 2492 760
rect 1750 660 1850 720
rect 2392 671 2492 720
rect 124 486 224 556
rect 124 351 244 486
rect 124 305 150 351
rect 196 305 244 351
rect 124 232 244 305
rect 348 351 448 556
rect 496 480 596 556
rect 496 434 520 480
rect 566 434 596 480
rect 496 421 596 434
rect 348 305 375 351
rect 421 305 448 351
rect 348 276 448 305
rect 740 419 840 556
rect 888 512 988 556
rect 2188 590 2288 634
rect 2392 625 2433 671
rect 2479 625 2492 671
rect 3068 720 4172 760
rect 2864 660 2964 704
rect 3068 660 3168 720
rect 2392 590 2492 625
rect 2540 590 2640 634
rect 740 373 753 419
rect 799 373 840 419
rect 740 276 840 373
rect 1432 415 1532 497
rect 1432 369 1455 415
rect 1501 369 1532 415
rect 908 337 1028 350
rect 908 291 956 337
rect 1002 291 1028 337
rect 348 232 468 276
rect 516 232 636 276
rect 740 232 860 276
rect 908 232 1028 291
rect 1432 281 1532 369
rect 1750 363 1850 497
rect 1750 317 1763 363
rect 1809 317 1850 363
rect 2188 456 2288 518
rect 2188 410 2201 456
rect 2247 410 2288 456
rect 2392 454 2492 518
rect 2540 485 2640 518
rect 3520 659 3620 672
rect 3520 613 3537 659
rect 3583 613 3620 659
rect 3520 580 3620 613
rect 3724 580 3824 624
rect 4072 591 4172 720
rect 4532 716 4632 760
rect 4736 716 4836 760
rect 4940 716 5040 760
rect 5147 716 5247 760
rect 5353 716 5453 760
rect 5585 716 5685 760
rect 4276 591 4376 635
rect 2540 439 2581 485
rect 2627 439 2640 485
rect 2540 426 2640 439
rect 2188 378 2288 410
rect 2188 338 2552 378
rect 1750 281 1850 317
rect 2432 298 2552 338
rect 124 64 244 156
rect 348 112 468 156
rect 516 64 636 156
rect 740 112 860 156
rect 908 112 1028 156
rect 124 24 636 64
rect 1432 237 1552 281
rect 1750 237 1870 281
rect 2208 219 2328 263
rect 2432 252 2473 298
rect 2519 252 2552 298
rect 2432 219 2552 252
rect 2600 263 2640 426
rect 2864 412 2964 497
rect 2864 392 3020 412
rect 2864 346 2877 392
rect 2923 346 3020 392
rect 2864 333 3020 346
rect 2600 219 2720 263
rect 2900 257 3020 333
rect 3068 304 3168 497
rect 3520 304 3620 497
rect 3724 423 3824 497
rect 3068 257 3188 304
rect 3292 257 3412 304
rect 3520 301 3636 304
rect 3516 257 3636 301
rect 1432 100 1552 144
rect 1750 64 1870 144
rect 2900 141 3020 185
rect 3068 141 3188 185
rect 3292 152 3412 185
rect 2208 64 2328 124
rect 2432 80 2552 124
rect 2600 80 2720 124
rect 3292 106 3305 152
rect 3351 106 3412 152
rect 3516 141 3636 185
rect 1750 24 2328 64
rect 3292 64 3412 106
rect 3784 64 3824 423
rect 4072 453 4172 497
rect 4072 324 4149 453
rect 4029 311 4149 324
rect 4029 265 4042 311
rect 4088 265 4149 311
rect 4276 439 4376 497
rect 4276 393 4317 439
rect 4363 393 4376 439
rect 4276 380 4376 393
rect 4276 287 4317 380
rect 4532 351 4632 472
rect 4736 417 4836 472
rect 4736 351 4809 417
rect 4940 380 5040 472
rect 5147 380 5247 472
rect 5353 380 5453 472
rect 5585 380 5685 472
rect 4532 350 4809 351
rect 4029 232 4149 265
rect 4197 232 4317 287
rect 4465 337 4809 350
rect 4465 291 4498 337
rect 4544 311 4809 337
rect 4544 291 4585 311
rect 4465 232 4585 291
rect 4689 232 4809 311
rect 4913 361 5705 380
rect 4913 315 4964 361
rect 5386 315 5705 361
rect 4913 296 5705 315
rect 4913 232 5033 296
rect 5137 232 5257 296
rect 5361 232 5481 296
rect 5585 232 5705 296
rect 4029 114 4149 158
rect 4197 114 4317 158
rect 3292 24 3824 64
rect 4465 24 4585 69
rect 4689 24 4809 69
rect 4913 24 5033 69
rect 5137 24 5257 69
rect 5361 24 5481 69
rect 5585 24 5705 69
<< polycontact >>
rect 150 305 196 351
rect 520 434 566 480
rect 375 305 421 351
rect 2433 625 2479 671
rect 753 373 799 419
rect 1455 369 1501 415
rect 956 291 1002 337
rect 1763 317 1809 363
rect 2201 410 2247 456
rect 3537 613 3583 659
rect 2581 439 2627 485
rect 2473 252 2519 298
rect 2877 346 2923 392
rect 3305 106 3351 152
rect 4042 265 4088 311
rect 4317 393 4363 439
rect 4498 291 4544 337
rect 4964 315 5386 361
<< metal1 >>
rect 0 724 5936 844
rect 49 615 95 628
rect 252 615 320 724
rect 1050 707 1118 724
rect 1050 661 1061 707
rect 1107 661 1118 707
rect 1620 716 1688 724
rect 1164 632 1558 678
rect 1620 670 1631 716
rect 1677 670 1688 716
rect 2702 718 2770 724
rect 2702 672 2713 718
rect 2759 672 2770 718
rect 1164 615 1210 632
rect 252 569 263 615
rect 309 569 320 615
rect 654 569 665 615
rect 711 569 1210 615
rect 1512 624 1558 632
rect 1773 624 2170 659
rect 1512 613 2170 624
rect 1512 578 1819 613
rect 2102 577 2170 613
rect 2422 625 2433 671
rect 2479 626 2490 671
rect 2864 632 3142 678
rect 2864 626 2910 632
rect 2479 625 2910 626
rect 49 523 95 569
rect 1357 556 1414 567
rect 49 480 1013 523
rect 1403 532 1414 556
rect 1879 556 1999 567
rect 1403 510 1809 532
rect 1357 486 1809 510
rect 1925 510 1999 556
rect 2102 531 2113 577
rect 2159 531 2170 577
rect 2317 577 2363 603
rect 2422 580 2910 625
rect 1879 499 1999 510
rect 49 477 520 480
rect 49 219 95 477
rect 566 477 1013 480
rect 49 156 95 173
rect 141 351 206 430
rect 141 305 150 351
rect 196 305 206 351
rect 141 119 206 305
rect 365 351 430 430
rect 520 421 566 434
rect 682 419 886 430
rect 682 373 753 419
rect 799 373 886 419
rect 682 354 886 373
rect 365 305 375 351
rect 421 305 430 351
rect 273 215 319 232
rect 273 60 319 169
rect 365 119 430 305
rect 945 337 1013 477
rect 1242 415 1558 430
rect 1242 369 1455 415
rect 1501 369 1558 415
rect 1242 354 1558 369
rect 1763 363 1809 486
rect 945 291 956 337
rect 1002 291 1013 337
rect 1763 279 1809 317
rect 1302 244 1809 279
rect 654 173 665 219
rect 711 187 722 219
rect 1302 198 1313 244
rect 1359 233 1809 244
rect 1942 456 1999 499
rect 1942 410 2201 456
rect 2247 410 2258 456
rect 1942 409 2258 410
rect 1942 244 2010 409
rect 2317 392 2363 531
rect 2982 510 2993 556
rect 3039 510 3050 556
rect 2982 485 3050 510
rect 3096 540 3142 632
rect 3197 647 3243 724
rect 3197 586 3243 601
rect 3340 659 3598 662
rect 3340 613 3537 659
rect 3583 613 3598 659
rect 3340 608 3598 613
rect 3340 540 3386 608
rect 3986 578 4054 724
rect 3649 562 3695 578
rect 3096 493 3386 540
rect 3434 516 3445 562
rect 3491 516 3502 562
rect 2570 439 2581 485
rect 2627 439 3050 485
rect 2570 438 3050 439
rect 2993 408 3050 438
rect 3434 408 3502 516
rect 3649 421 3695 516
rect 2317 346 2877 392
rect 2923 346 2934 392
rect 2993 361 3502 408
rect 3562 375 3695 421
rect 3853 562 3899 578
rect 3986 532 3997 578
rect 4043 532 4054 578
rect 4457 665 4503 724
rect 4201 556 4247 567
rect 3853 486 3899 516
rect 4201 486 4247 510
rect 4457 506 4503 525
rect 4661 665 4707 676
rect 3853 440 4247 486
rect 2317 345 2934 346
rect 1359 198 1370 233
rect 1942 198 1953 244
rect 1999 198 2010 244
rect 711 173 1250 187
rect 654 152 1250 173
rect 1522 152 1863 187
rect 2133 183 2179 194
rect 654 141 2133 152
rect 1204 106 1568 141
rect 1817 137 2133 141
rect 1817 106 2179 137
rect 2357 193 2403 345
rect 2462 298 2995 299
rect 2462 252 2473 298
rect 2519 252 2995 298
rect 2357 136 2403 147
rect 2770 137 2781 183
rect 2827 137 2838 183
rect 1090 60 1101 95
rect 0 49 1101 60
rect 1147 60 1158 95
rect 1614 60 1625 95
rect 1147 49 1625 60
rect 1671 60 1682 95
rect 2770 60 2838 137
rect 2949 152 2995 252
rect 3206 244 3274 361
rect 3562 244 3608 375
rect 3853 244 3899 440
rect 4661 439 4707 525
rect 4865 665 4911 724
rect 4865 506 4911 525
rect 5062 665 5128 676
rect 5062 525 5072 665
rect 5118 525 5128 665
rect 4306 393 4317 439
rect 4363 393 4707 439
rect 5062 458 5128 525
rect 5276 665 5322 724
rect 5276 506 5322 525
rect 5488 665 5582 676
rect 5488 525 5495 665
rect 5541 525 5582 665
rect 5488 458 5582 525
rect 5714 665 5760 724
rect 5714 506 5760 525
rect 5062 411 5582 458
rect 4614 361 4707 393
rect 4015 311 4246 318
rect 4015 265 4042 311
rect 4088 265 4246 311
rect 3206 198 3217 244
rect 3263 198 3274 244
rect 3430 198 3441 244
rect 3487 198 3608 244
rect 3654 198 3665 244
rect 3711 198 3897 244
rect 3943 198 3954 244
rect 4015 242 4246 265
rect 4298 291 4498 337
rect 4544 291 4555 337
rect 4298 290 4555 291
rect 4614 315 4964 361
rect 5386 315 5421 361
rect 3562 152 3608 198
rect 4298 152 4344 290
rect 4614 218 4660 315
rect 5488 269 5582 411
rect 2949 106 3305 152
rect 3351 106 3362 152
rect 3562 106 4344 152
rect 4390 193 4436 204
rect 4614 161 4660 172
rect 4838 218 4884 229
rect 4390 60 4436 147
rect 4838 60 4884 172
rect 5062 223 5582 269
rect 5062 218 5108 223
rect 5062 161 5108 172
rect 5488 218 5582 223
rect 5488 172 5510 218
rect 5556 172 5582 218
rect 5275 149 5343 150
rect 5275 103 5286 149
rect 5332 103 5343 149
rect 5488 119 5582 172
rect 5734 218 5780 229
rect 5275 60 5343 103
rect 5734 60 5780 172
rect 1671 49 5936 60
rect 0 -60 5936 49
<< labels >>
flabel metal1 s 682 354 886 430 0 FreeSans 600 0 0 0 D
port 1 nsew default input
flabel metal1 s 5488 458 5582 676 0 FreeSans 600 0 0 0 Q
port 6 nsew default output
flabel metal1 s 141 119 206 430 0 FreeSans 600 0 0 0 SE
port 2 nsew default input
flabel metal1 s 4015 242 4246 318 0 FreeSans 600 0 0 0 SETN
port 3 nsew default input
flabel metal1 s 365 119 430 430 0 FreeSans 600 0 0 0 SI
port 4 nsew default input
flabel metal1 s 0 724 5936 844 0 FreeSans 600 0 0 0 VDD
port 7 nsew power bidirectional abutment
flabel metal1 s 273 229 319 232 0 FreeSans 600 0 0 0 VSS
port 10 nsew ground bidirectional abutment
flabel metal1 s 1242 354 1558 430 0 FreeSans 600 0 0 0 CLK
port 5 nsew clock input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 8 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 9 nsew ground bidirectional
rlabel metal1 s 5062 458 5128 676 1 Q
port 6 nsew default output
rlabel metal1 s 5062 411 5582 458 1 Q
port 6 nsew default output
rlabel metal1 s 5488 269 5582 411 1 Q
port 6 nsew default output
rlabel metal1 s 5062 223 5582 269 1 Q
port 6 nsew default output
rlabel metal1 s 5488 161 5582 223 1 Q
port 6 nsew default output
rlabel metal1 s 5062 161 5108 223 1 Q
port 6 nsew default output
rlabel metal1 s 5488 119 5582 161 1 Q
port 6 nsew default output
rlabel metal1 s 5714 672 5760 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5276 672 5322 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4865 672 4911 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4457 672 4503 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3986 672 4054 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3197 672 3243 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2702 672 2770 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1620 672 1688 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1050 672 1118 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 252 672 320 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5714 670 5760 672 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5276 670 5322 672 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4865 670 4911 672 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4457 670 4503 672 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3986 670 4054 672 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3197 670 3243 672 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1620 670 1688 672 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1050 670 1118 672 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 252 670 320 672 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5714 661 5760 670 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5276 661 5322 670 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4865 661 4911 670 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4457 661 4503 670 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3986 661 4054 670 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3197 661 3243 670 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1050 661 1118 670 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 252 661 320 670 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5714 586 5760 661 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5276 586 5322 661 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4865 586 4911 661 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4457 586 4503 661 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3986 586 4054 661 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3197 586 3243 661 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 252 586 320 661 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5714 569 5760 586 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5276 569 5322 586 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4865 569 4911 586 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4457 569 4503 586 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3986 569 4054 586 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 252 569 320 586 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5714 532 5760 569 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5276 532 5322 569 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4865 532 4911 569 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4457 532 4503 569 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3986 532 4054 569 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5714 506 5760 532 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5276 506 5322 532 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4865 506 4911 532 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4457 506 4503 532 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5734 204 5780 229 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 4838 204 4884 229 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 273 204 319 229 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 5734 183 5780 204 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 4838 183 4884 204 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 4390 183 4436 204 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 273 183 319 204 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 5734 150 5780 183 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 4838 150 4884 183 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 4390 150 4436 183 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 2770 150 2838 183 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 273 150 319 183 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 5734 95 5780 150 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 5275 95 5343 150 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 4838 95 4884 150 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 4390 95 4436 150 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 2770 95 2838 150 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 273 95 319 150 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 5734 60 5780 95 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 5275 60 5343 95 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 4838 60 4884 95 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 4390 60 4436 95 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 2770 60 2838 95 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 1614 60 1682 95 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 1090 60 1158 95 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 273 60 319 95 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 5936 60 1 VSS
port 10 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 5936 784
string GDS_END 316014
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 304126
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
