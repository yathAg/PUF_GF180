magic
tech gf180mcuB
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 352 4342 870
<< pwell >>
rect -86 -86 4342 352
<< metal1 >>
rect 0 724 4256 844
rect 49 515 95 724
rect 49 60 95 226
rect 141 205 202 567
rect 451 360 740 450
rect 660 248 740 360
rect 1024 569 1092 724
rect 1246 430 1323 585
rect 1470 569 1538 724
rect 1685 430 1768 585
rect 1906 569 1974 724
rect 901 360 1151 430
rect 1246 360 1768 430
rect 901 110 987 360
rect 1033 60 1079 232
rect 1246 120 1320 360
rect 1481 60 1527 232
rect 1685 120 1768 360
rect 1929 60 1975 232
rect 2481 430 2555 664
rect 2282 354 2555 430
rect 2282 261 2355 354
rect 3029 569 3098 724
rect 2815 356 3195 426
rect 3021 60 3067 229
rect 3886 563 3954 724
rect 3745 356 4083 424
rect 3917 60 3963 229
rect 0 -60 4256 60
<< obsm1 >>
rect 542 620 947 666
rect 542 594 610 620
rect 252 215 299 590
rect 345 548 610 594
rect 345 314 391 548
rect 345 268 458 314
rect 408 215 458 268
rect 252 169 330 215
rect 408 169 582 215
rect 786 156 855 574
rect 901 523 947 620
rect 1151 632 1424 678
rect 1151 523 1197 632
rect 901 476 1197 523
rect 1378 523 1424 632
rect 1584 631 1860 678
rect 1584 523 1630 631
rect 1378 476 1630 523
rect 1814 523 1860 631
rect 2098 523 2144 601
rect 1814 476 2144 523
rect 2190 544 2424 590
rect 2021 226 2067 476
rect 2190 364 2236 544
rect 2113 292 2236 364
rect 2021 158 2144 226
rect 2190 215 2236 292
rect 2625 632 2966 678
rect 2190 169 2438 215
rect 2625 156 2671 632
rect 2717 515 2863 585
rect 2920 523 2966 632
rect 3148 632 3515 678
rect 3148 523 3194 632
rect 2717 229 2767 515
rect 2920 476 3194 523
rect 2717 159 2863 229
rect 3245 156 3291 585
rect 3449 156 3515 632
rect 3561 563 3733 609
rect 3561 216 3607 563
rect 4120 517 4187 628
rect 3653 471 4187 517
rect 3653 335 3699 471
rect 3561 170 3750 216
rect 4141 156 4187 471
<< labels >>
rlabel metal1 s 3745 356 4083 424 6 I0
port 1 nsew default input
rlabel metal1 s 2815 356 3195 426 6 I1
port 2 nsew default input
rlabel metal1 s 141 205 202 567 6 I2
port 3 nsew default input
rlabel metal1 s 901 110 987 360 6 I3
port 4 nsew default input
rlabel metal1 s 901 360 1151 430 6 I3
port 4 nsew default input
rlabel metal1 s 660 248 740 360 6 S0
port 5 nsew default input
rlabel metal1 s 451 360 740 450 6 S0
port 5 nsew default input
rlabel metal1 s 2282 261 2355 354 6 S1
port 6 nsew default input
rlabel metal1 s 2282 354 2555 430 6 S1
port 6 nsew default input
rlabel metal1 s 2481 430 2555 664 6 S1
port 6 nsew default input
rlabel metal1 s 1685 120 1768 360 6 Z
port 7 nsew default output
rlabel metal1 s 1246 120 1320 360 6 Z
port 7 nsew default output
rlabel metal1 s 1246 360 1768 430 6 Z
port 7 nsew default output
rlabel metal1 s 1685 430 1768 585 6 Z
port 7 nsew default output
rlabel metal1 s 1246 430 1323 585 6 Z
port 7 nsew default output
rlabel metal1 s 3886 563 3954 724 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3029 569 3098 724 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1906 569 1974 724 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1470 569 1538 724 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1024 569 1092 724 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 49 515 95 724 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 724 4256 844 6 VDD
port 8 nsew power bidirectional abutment
rlabel nwell s -86 352 4342 870 6 VNW
port 9 nsew power bidirectional
rlabel pwell s -86 -86 4342 352 6 VPW
port 10 nsew ground bidirectional
rlabel metal1 s 0 -60 4256 60 8 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 3917 60 3963 229 6 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 3021 60 3067 229 6 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 1929 60 1975 232 6 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 1481 60 1527 232 6 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 1033 60 1079 232 6 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 226 6 VSS
port 11 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4256 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 698698
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 690048
<< end >>
