magic
tech gf180mcuB
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 352 1206 870
<< pwell >>
rect -86 -86 1206 352
<< metal1 >>
rect 0 724 1120 844
rect 130 232 200 438
rect 248 200 308 545
rect 584 570 802 662
rect 354 354 538 430
rect 354 246 430 354
rect 584 346 644 570
rect 906 506 952 724
rect 690 354 990 430
rect 610 209 972 255
rect 610 200 656 209
rect 50 60 96 174
rect 248 112 656 200
rect 702 60 748 163
rect 926 113 972 209
rect 0 -60 1120 60
<< obsm1 >>
rect 50 630 504 676
rect 50 506 96 630
rect 458 506 504 630
<< labels >>
rlabel metal1 s 354 246 430 354 6 A1
port 1 nsew default input
rlabel metal1 s 354 354 538 430 6 A1
port 1 nsew default input
rlabel metal1 s 130 232 200 438 6 A2
port 2 nsew default input
rlabel metal1 s 584 346 644 570 6 B
port 3 nsew default input
rlabel metal1 s 584 570 802 662 6 B
port 3 nsew default input
rlabel metal1 s 690 354 990 430 6 C
port 4 nsew default input
rlabel metal1 s 926 113 972 209 6 ZN
port 5 nsew default output
rlabel metal1 s 248 112 656 200 6 ZN
port 5 nsew default output
rlabel metal1 s 610 200 656 209 6 ZN
port 5 nsew default output
rlabel metal1 s 610 209 972 255 6 ZN
port 5 nsew default output
rlabel metal1 s 248 200 308 545 6 ZN
port 5 nsew default output
rlabel metal1 s 906 506 952 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 724 1120 844 6 VDD
port 6 nsew power bidirectional abutment
rlabel nwell s -86 352 1206 870 6 VNW
port 7 nsew power bidirectional
rlabel pwell s -86 -86 1206 352 6 VPW
port 8 nsew ground bidirectional
rlabel metal1 s 0 -60 1120 60 8 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 702 60 748 163 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 50 60 96 174 6 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1120 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1280044
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1276526
<< end >>
