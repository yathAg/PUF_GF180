magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 453 4230 1094
<< pwell >>
rect -86 -86 4230 453
<< mvnmos >>
rect 124 175 244 333
rect 348 175 468 333
rect 716 194 836 312
rect 940 194 1060 312
rect 1176 194 1296 312
rect 1346 194 1466 312
rect 1614 215 1734 333
rect 1782 215 1902 333
rect 2006 215 2126 333
rect 2230 215 2350 333
rect 2862 215 2982 333
rect 3030 215 3150 333
rect 3298 69 3418 333
rect 3676 69 3796 333
rect 3900 69 4020 333
<< mvpmos >>
rect 144 573 244 849
rect 348 573 448 849
rect 736 593 836 793
rect 989 593 1089 793
rect 1193 593 1293 793
rect 1366 593 1466 793
rect 1586 593 1686 793
rect 1802 593 1902 793
rect 2230 573 2330 773
rect 2498 573 2598 773
rect 2846 573 2946 773
rect 3050 573 3150 773
rect 3298 573 3398 939
rect 3696 573 3796 939
rect 3900 573 4000 939
<< mvndiff >>
rect 36 320 124 333
rect 36 274 49 320
rect 95 274 124 320
rect 36 175 124 274
rect 244 234 348 333
rect 244 188 273 234
rect 319 188 348 234
rect 244 175 348 188
rect 468 320 556 333
rect 468 274 497 320
rect 543 274 556 320
rect 1534 312 1614 333
rect 468 175 556 274
rect 628 253 716 312
rect 628 207 641 253
rect 687 207 716 253
rect 628 194 716 207
rect 836 299 940 312
rect 836 253 865 299
rect 911 253 940 299
rect 836 194 940 253
rect 1060 299 1176 312
rect 1060 253 1089 299
rect 1135 253 1176 299
rect 1060 194 1176 253
rect 1296 194 1346 312
rect 1466 253 1614 312
rect 1466 207 1495 253
rect 1541 215 1614 253
rect 1734 215 1782 333
rect 1902 320 2006 333
rect 1902 274 1931 320
rect 1977 274 2006 320
rect 1902 215 2006 274
rect 2126 274 2230 333
rect 2126 228 2155 274
rect 2201 228 2230 274
rect 2126 215 2230 228
rect 2350 320 2438 333
rect 2350 274 2379 320
rect 2425 274 2438 320
rect 2350 215 2438 274
rect 1541 207 1554 215
rect 1466 194 1554 207
rect 2774 299 2862 333
rect 2774 253 2787 299
rect 2833 253 2862 299
rect 2774 215 2862 253
rect 2982 215 3030 333
rect 3150 222 3298 333
rect 3150 215 3223 222
rect 3210 82 3223 215
rect 3269 82 3298 222
rect 3210 69 3298 82
rect 3418 320 3506 333
rect 3418 180 3447 320
rect 3493 180 3506 320
rect 3418 69 3506 180
rect 3588 222 3676 333
rect 3588 82 3601 222
rect 3647 82 3676 222
rect 3588 69 3676 82
rect 3796 320 3900 333
rect 3796 180 3825 320
rect 3871 180 3900 320
rect 3796 69 3900 180
rect 4020 222 4108 333
rect 4020 82 4049 222
rect 4095 82 4108 222
rect 4020 69 4108 82
<< mvpdiff >>
rect 56 637 144 849
rect 56 591 69 637
rect 115 591 144 637
rect 56 573 144 591
rect 244 836 348 849
rect 244 790 273 836
rect 319 790 348 836
rect 244 573 348 790
rect 448 632 536 849
rect 1962 823 2034 836
rect 1962 793 1975 823
rect 448 586 477 632
rect 523 586 536 632
rect 648 780 736 793
rect 648 734 661 780
rect 707 734 736 780
rect 648 593 736 734
rect 836 746 989 793
rect 836 606 865 746
rect 911 606 989 746
rect 836 593 989 606
rect 1089 746 1193 793
rect 1089 606 1118 746
rect 1164 606 1193 746
rect 1089 593 1193 606
rect 1293 593 1366 793
rect 1466 780 1586 793
rect 1466 734 1495 780
rect 1541 734 1586 780
rect 1466 593 1586 734
rect 1686 652 1802 793
rect 1686 606 1715 652
rect 1761 606 1802 652
rect 1686 593 1802 606
rect 1902 777 1975 793
rect 2021 777 2034 823
rect 1902 593 2034 777
rect 3218 773 3298 939
rect 2142 632 2230 773
rect 448 573 536 586
rect 2142 586 2155 632
rect 2201 586 2230 632
rect 2142 573 2230 586
rect 2330 726 2498 773
rect 2330 586 2359 726
rect 2405 586 2498 726
rect 2330 573 2498 586
rect 2598 632 2686 773
rect 2598 586 2627 632
rect 2673 586 2686 632
rect 2598 573 2686 586
rect 2758 760 2846 773
rect 2758 714 2771 760
rect 2817 714 2846 760
rect 2758 573 2846 714
rect 2946 748 3050 773
rect 2946 608 2975 748
rect 3021 608 3050 748
rect 2946 573 3050 608
rect 3150 760 3298 773
rect 3150 620 3179 760
rect 3225 620 3298 760
rect 3150 573 3298 620
rect 3398 726 3486 939
rect 3398 586 3427 726
rect 3473 586 3486 726
rect 3398 573 3486 586
rect 3608 926 3696 939
rect 3608 786 3621 926
rect 3667 786 3696 926
rect 3608 573 3696 786
rect 3796 726 3900 939
rect 3796 586 3825 726
rect 3871 586 3900 726
rect 3796 573 3900 586
rect 4000 926 4088 939
rect 4000 786 4029 926
rect 4075 786 4088 926
rect 4000 573 4088 786
<< mvndiffc >>
rect 49 274 95 320
rect 273 188 319 234
rect 497 274 543 320
rect 641 207 687 253
rect 865 253 911 299
rect 1089 253 1135 299
rect 1495 207 1541 253
rect 1931 274 1977 320
rect 2155 228 2201 274
rect 2379 274 2425 320
rect 2787 253 2833 299
rect 3223 82 3269 222
rect 3447 180 3493 320
rect 3601 82 3647 222
rect 3825 180 3871 320
rect 4049 82 4095 222
<< mvpdiffc >>
rect 69 591 115 637
rect 273 790 319 836
rect 477 586 523 632
rect 661 734 707 780
rect 865 606 911 746
rect 1118 606 1164 746
rect 1495 734 1541 780
rect 1715 606 1761 652
rect 1975 777 2021 823
rect 2155 586 2201 632
rect 2359 586 2405 726
rect 2627 586 2673 632
rect 2771 714 2817 760
rect 2975 608 3021 748
rect 3179 620 3225 760
rect 3427 586 3473 726
rect 3621 786 3667 926
rect 3825 586 3871 726
rect 4029 786 4075 926
<< polysilicon >>
rect 348 933 1293 973
rect 144 849 244 893
rect 348 849 448 933
rect 989 872 1089 885
rect 736 793 836 837
rect 989 826 1002 872
rect 1048 826 1089 872
rect 989 793 1089 826
rect 1193 872 1293 933
rect 1193 826 1234 872
rect 1280 826 1293 872
rect 1802 913 2946 953
rect 3298 939 3398 983
rect 3696 939 3796 983
rect 3900 939 4000 983
rect 1193 793 1293 826
rect 1366 793 1466 837
rect 1586 793 1686 837
rect 1802 793 1902 913
rect 2230 852 2330 865
rect 2230 806 2243 852
rect 2289 806 2330 852
rect 2230 773 2330 806
rect 2498 773 2598 817
rect 2846 773 2946 913
rect 3050 773 3150 817
rect 144 494 244 573
rect 144 448 157 494
rect 203 448 244 494
rect 144 377 244 448
rect 124 333 244 377
rect 348 412 448 573
rect 348 366 361 412
rect 407 377 448 412
rect 736 411 836 593
rect 989 533 1089 593
rect 1193 549 1293 593
rect 1366 560 1466 593
rect 989 493 1147 533
rect 407 366 468 377
rect 348 333 468 366
rect 736 365 749 411
rect 795 365 836 411
rect 1107 412 1147 493
rect 1366 514 1407 560
rect 1453 514 1466 560
rect 1586 549 1686 593
rect 1107 391 1296 412
rect 1107 372 1237 391
rect 736 356 836 365
rect 716 312 836 356
rect 940 312 1060 356
rect 1176 345 1237 372
rect 1283 345 1296 391
rect 1366 356 1466 514
rect 1176 312 1296 345
rect 1346 312 1466 356
rect 1614 468 1686 549
rect 1614 422 1627 468
rect 1673 422 1686 468
rect 1614 377 1686 422
rect 1802 377 1902 593
rect 2230 377 2330 573
rect 2498 529 2598 573
rect 1614 333 1734 377
rect 1782 333 1902 377
rect 2006 333 2126 377
rect 2230 333 2350 377
rect 124 131 244 175
rect 348 102 468 175
rect 716 150 836 194
rect 940 102 1060 194
rect 1176 150 1296 194
rect 1346 150 1466 194
rect 1614 171 1734 215
rect 1782 171 1902 215
rect 2006 182 2126 215
rect 348 62 1060 102
rect 2006 136 2019 182
rect 2065 136 2126 182
rect 2230 171 2350 215
rect 2006 123 2126 136
rect 2498 123 2597 529
rect 2846 412 2946 573
rect 2846 393 2887 412
rect 2862 366 2887 393
rect 2933 393 2946 412
rect 3050 515 3150 573
rect 3050 469 3091 515
rect 3137 469 3150 515
rect 2933 366 2982 393
rect 3050 377 3150 469
rect 2862 333 2982 366
rect 3030 333 3150 377
rect 3298 412 3398 573
rect 3298 366 3311 412
rect 3357 377 3398 412
rect 3696 471 3796 573
rect 3900 471 4000 573
rect 3696 412 4000 471
rect 3696 377 3709 412
rect 3357 366 3418 377
rect 3298 333 3418 366
rect 3676 366 3709 377
rect 3755 393 4000 412
rect 3755 366 3796 393
rect 3676 333 3796 366
rect 3900 377 4000 393
rect 3900 333 4020 377
rect 2862 171 2982 215
rect 3030 171 3150 215
rect 2006 83 2597 123
rect 3298 25 3418 69
rect 3676 25 3796 69
rect 3900 25 4020 69
<< polycontact >>
rect 1002 826 1048 872
rect 1234 826 1280 872
rect 2243 806 2289 852
rect 157 448 203 494
rect 361 366 407 412
rect 749 365 795 411
rect 1407 514 1453 560
rect 1237 345 1283 391
rect 1627 422 1673 468
rect 2019 136 2065 182
rect 2887 366 2933 412
rect 3091 469 3137 515
rect 3311 366 3357 412
rect 3709 366 3755 412
<< metal1 >>
rect 0 926 4144 1098
rect 0 918 3621 926
rect 273 836 319 918
rect 273 779 319 790
rect 661 780 707 918
rect 661 723 707 734
rect 753 826 1002 872
rect 1048 826 1059 872
rect 1223 826 1234 872
rect 1280 826 1291 872
rect 69 637 407 648
rect 753 643 799 826
rect 115 602 407 637
rect 69 580 115 591
rect 142 494 278 542
rect 142 448 157 494
rect 203 448 278 494
rect 361 412 407 602
rect 361 348 407 366
rect 49 320 407 348
rect 95 302 407 320
rect 477 632 799 643
rect 523 597 799 632
rect 865 746 911 757
rect 523 586 543 597
rect 477 320 543 586
rect 615 411 795 430
rect 615 365 749 411
rect 615 354 795 365
rect 49 263 95 274
rect 477 274 497 320
rect 477 263 543 274
rect 865 299 911 606
rect 641 253 687 264
rect 273 234 319 245
rect 273 90 319 188
rect 865 242 911 253
rect 1089 746 1164 757
rect 1089 606 1118 746
rect 1223 677 1291 826
rect 1495 780 1541 918
rect 1975 823 2021 918
rect 1975 766 2021 777
rect 2243 852 2289 863
rect 1495 723 1541 734
rect 1587 720 1930 755
rect 2243 735 2289 806
rect 2771 760 2817 918
rect 2055 720 2289 735
rect 1587 709 2289 720
rect 1587 677 1633 709
rect 1223 631 1633 677
rect 1885 689 2289 709
rect 2359 726 2405 737
rect 1885 674 2089 689
rect 1715 652 1761 663
rect 1089 483 1164 606
rect 1715 560 1761 606
rect 2155 632 2201 643
rect 2155 560 2201 586
rect 1396 514 1407 560
rect 1453 514 2201 560
rect 3179 760 3225 918
rect 3667 918 4029 926
rect 3621 775 3667 786
rect 4075 918 4144 926
rect 4029 775 4075 786
rect 2771 703 2817 714
rect 2975 748 3021 759
rect 1089 468 1362 483
rect 1089 437 1627 468
rect 1089 299 1135 437
rect 1328 422 1627 437
rect 1673 422 1684 468
rect 1226 345 1237 391
rect 1283 376 1294 391
rect 1283 345 1633 376
rect 1226 330 1633 345
rect 1089 242 1135 253
rect 1495 253 1541 264
rect 641 90 687 207
rect 1495 90 1541 207
rect 1587 182 1633 330
rect 1931 320 1977 514
rect 2359 423 2405 586
rect 2287 377 2405 423
rect 2627 632 2975 643
rect 2673 608 2975 632
rect 3179 609 3225 620
rect 3427 726 3489 737
rect 2673 597 3021 608
rect 1931 263 1977 274
rect 2155 274 2201 285
rect 2155 196 2201 228
rect 2287 196 2333 377
rect 2627 331 2673 586
rect 3473 586 3489 726
rect 3427 526 3489 586
rect 3091 515 3489 526
rect 3137 469 3489 515
rect 3091 458 3489 469
rect 3443 423 3489 458
rect 3825 726 3890 737
rect 3871 586 3890 726
rect 2379 320 2673 331
rect 2425 310 2673 320
rect 2887 412 2933 423
rect 3443 412 3755 423
rect 2887 318 2933 366
rect 3040 366 3311 412
rect 3357 366 3368 412
rect 3443 366 3709 412
rect 2425 299 2833 310
rect 2425 274 2787 299
rect 2379 253 2787 274
rect 2379 242 2833 253
rect 2887 242 2994 318
rect 3040 196 3086 366
rect 3443 355 3755 366
rect 3443 320 3493 355
rect 1587 136 2019 182
rect 2065 136 2076 182
rect 2155 150 3086 196
rect 3223 222 3269 233
rect 0 82 3223 90
rect 3443 180 3447 320
rect 3825 320 3890 586
rect 3443 169 3493 180
rect 3601 222 3647 233
rect 3269 82 3601 90
rect 3871 180 3890 320
rect 3825 169 3890 180
rect 4049 222 4095 233
rect 3647 82 4049 90
rect 4095 82 4144 90
rect 0 -90 4144 82
<< labels >>
flabel metal1 s 142 448 278 542 0 FreeSans 200 0 0 0 CLK
port 3 nsew clock input
flabel metal1 s 615 354 795 430 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 3825 169 3890 737 0 FreeSans 200 0 0 0 Q
port 4 nsew default output
flabel metal1 s 2887 318 2933 423 0 FreeSans 200 0 0 0 SETN
port 2 nsew default input
flabel metal1 s 0 918 4144 1098 0 FreeSans 200 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 1495 245 1541 264 0 FreeSans 200 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 6 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 2887 242 2994 318 1 SETN
port 2 nsew default input
rlabel metal1 s 4029 779 4075 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3621 779 3667 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3179 779 3225 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2771 779 2817 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1975 779 2021 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1495 779 1541 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 661 779 707 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 779 319 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4029 775 4075 779 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3621 775 3667 779 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3179 775 3225 779 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2771 775 2817 779 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1975 775 2021 779 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1495 775 1541 779 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 661 775 707 779 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3179 766 3225 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2771 766 2817 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1975 766 2021 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1495 766 1541 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 661 766 707 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3179 723 3225 766 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2771 723 2817 766 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1495 723 1541 766 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 661 723 707 766 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3179 703 3225 723 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2771 703 2817 723 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3179 609 3225 703 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 641 245 687 264 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1495 233 1541 245 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 641 233 687 245 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 233 319 245 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4049 90 4095 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3601 90 3647 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3223 90 3269 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1495 90 1541 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 641 90 687 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 4144 90 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4144 1008
string GDS_END 683066
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 673668
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
