magic
tech gf180mcuB
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 352 7030 870
<< pwell >>
rect -86 -86 7030 352
<< mvnmos >>
rect 348 138 468 214
rect 572 138 692 214
rect 796 138 916 214
rect 1020 138 1140 214
rect 1244 138 1364 214
rect 1468 138 1588 214
rect 1692 138 1812 214
rect 1916 138 2036 214
rect 2400 138 2520 232
rect 2624 138 2744 232
rect 2848 138 2968 232
rect 3072 138 3192 232
rect 3296 138 3416 232
rect 3520 138 3640 232
rect 3744 138 3864 232
rect 3968 138 4088 232
rect 4192 138 4312 232
rect 4416 138 4536 232
rect 4640 138 4760 232
rect 4864 138 4984 232
rect 5088 138 5208 232
rect 5312 138 5432 232
rect 5536 138 5656 232
rect 5760 138 5880 232
rect 5984 138 6104 232
rect 6208 138 6328 232
rect 6432 138 6552 232
rect 6656 138 6776 232
<< mvpmos >>
rect 124 552 224 716
rect 348 552 448 716
rect 572 552 672 716
rect 796 552 896 716
rect 1020 552 1120 716
rect 1244 552 1344 716
rect 1468 552 1568 716
rect 1692 552 1792 716
rect 1916 552 2016 716
rect 2160 552 2260 716
rect 2400 472 2500 716
rect 2624 472 2724 716
rect 2848 472 2948 716
rect 3072 472 3172 716
rect 3296 472 3396 716
rect 3520 472 3620 716
rect 3744 472 3844 716
rect 3968 472 4068 716
rect 4192 472 4292 716
rect 4416 472 4516 716
rect 4640 472 4740 716
rect 4864 472 4964 716
rect 5088 472 5188 716
rect 5312 472 5412 716
rect 5536 472 5636 716
rect 5760 472 5860 716
rect 5984 472 6084 716
rect 6208 472 6308 716
rect 6432 472 6532 716
rect 6676 472 6776 716
<< mvndiff >>
rect 260 197 348 214
rect 260 151 273 197
rect 319 151 348 197
rect 260 138 348 151
rect 468 197 572 214
rect 468 151 497 197
rect 543 151 572 197
rect 468 138 572 151
rect 692 197 796 214
rect 692 151 721 197
rect 767 151 796 197
rect 692 138 796 151
rect 916 197 1020 214
rect 916 151 945 197
rect 991 151 1020 197
rect 916 138 1020 151
rect 1140 197 1244 214
rect 1140 151 1169 197
rect 1215 151 1244 197
rect 1140 138 1244 151
rect 1364 197 1468 214
rect 1364 151 1393 197
rect 1439 151 1468 197
rect 1364 138 1468 151
rect 1588 197 1692 214
rect 1588 151 1617 197
rect 1663 151 1692 197
rect 1588 138 1692 151
rect 1812 197 1916 214
rect 1812 151 1841 197
rect 1887 151 1916 197
rect 1812 138 1916 151
rect 2036 197 2124 214
rect 2036 151 2065 197
rect 2111 151 2124 197
rect 2036 138 2124 151
rect 2276 197 2400 232
rect 2276 151 2289 197
rect 2335 151 2400 197
rect 2276 138 2400 151
rect 2520 197 2624 232
rect 2520 151 2549 197
rect 2595 151 2624 197
rect 2520 138 2624 151
rect 2744 197 2848 232
rect 2744 151 2773 197
rect 2819 151 2848 197
rect 2744 138 2848 151
rect 2968 197 3072 232
rect 2968 151 2997 197
rect 3043 151 3072 197
rect 2968 138 3072 151
rect 3192 197 3296 232
rect 3192 151 3221 197
rect 3267 151 3296 197
rect 3192 138 3296 151
rect 3416 197 3520 232
rect 3416 151 3445 197
rect 3491 151 3520 197
rect 3416 138 3520 151
rect 3640 197 3744 232
rect 3640 151 3669 197
rect 3715 151 3744 197
rect 3640 138 3744 151
rect 3864 197 3968 232
rect 3864 151 3893 197
rect 3939 151 3968 197
rect 3864 138 3968 151
rect 4088 197 4192 232
rect 4088 151 4117 197
rect 4163 151 4192 197
rect 4088 138 4192 151
rect 4312 197 4416 232
rect 4312 151 4341 197
rect 4387 151 4416 197
rect 4312 138 4416 151
rect 4536 197 4640 232
rect 4536 151 4565 197
rect 4611 151 4640 197
rect 4536 138 4640 151
rect 4760 197 4864 232
rect 4760 151 4789 197
rect 4835 151 4864 197
rect 4760 138 4864 151
rect 4984 197 5088 232
rect 4984 151 5013 197
rect 5059 151 5088 197
rect 4984 138 5088 151
rect 5208 197 5312 232
rect 5208 151 5237 197
rect 5283 151 5312 197
rect 5208 138 5312 151
rect 5432 197 5536 232
rect 5432 151 5461 197
rect 5507 151 5536 197
rect 5432 138 5536 151
rect 5656 197 5760 232
rect 5656 151 5685 197
rect 5731 151 5760 197
rect 5656 138 5760 151
rect 5880 197 5984 232
rect 5880 151 5909 197
rect 5955 151 5984 197
rect 5880 138 5984 151
rect 6104 197 6208 232
rect 6104 151 6133 197
rect 6179 151 6208 197
rect 6104 138 6208 151
rect 6328 197 6432 232
rect 6328 151 6357 197
rect 6403 151 6432 197
rect 6328 138 6432 151
rect 6552 197 6656 232
rect 6552 151 6581 197
rect 6627 151 6656 197
rect 6552 138 6656 151
rect 6776 197 6864 232
rect 6776 151 6805 197
rect 6851 151 6864 197
rect 6776 138 6864 151
<< mvpdiff >>
rect 36 703 124 716
rect 36 657 49 703
rect 95 657 124 703
rect 36 552 124 657
rect 224 665 348 716
rect 224 619 273 665
rect 319 619 348 665
rect 224 552 348 619
rect 448 667 572 716
rect 448 621 477 667
rect 523 621 572 667
rect 448 552 572 621
rect 672 665 796 716
rect 672 619 701 665
rect 747 619 796 665
rect 672 552 796 619
rect 896 667 1020 716
rect 896 621 925 667
rect 971 621 1020 667
rect 896 552 1020 621
rect 1120 665 1244 716
rect 1120 619 1149 665
rect 1195 619 1244 665
rect 1120 552 1244 619
rect 1344 667 1468 716
rect 1344 621 1373 667
rect 1419 621 1468 667
rect 1344 552 1468 621
rect 1568 665 1692 716
rect 1568 619 1597 665
rect 1643 619 1692 665
rect 1568 552 1692 619
rect 1792 667 1916 716
rect 1792 621 1821 667
rect 1867 621 1916 667
rect 1792 552 1916 621
rect 2016 665 2160 716
rect 2016 619 2065 665
rect 2111 619 2160 665
rect 2016 552 2160 619
rect 2260 703 2400 716
rect 2260 657 2325 703
rect 2371 657 2400 703
rect 2260 552 2400 657
rect 2320 472 2400 552
rect 2500 665 2624 716
rect 2500 525 2549 665
rect 2595 525 2624 665
rect 2500 472 2624 525
rect 2724 703 2848 716
rect 2724 657 2753 703
rect 2799 657 2848 703
rect 2724 472 2848 657
rect 2948 665 3072 716
rect 2948 525 2977 665
rect 3023 525 3072 665
rect 2948 472 3072 525
rect 3172 703 3296 716
rect 3172 657 3201 703
rect 3247 657 3296 703
rect 3172 472 3296 657
rect 3396 665 3520 716
rect 3396 525 3425 665
rect 3471 525 3520 665
rect 3396 472 3520 525
rect 3620 703 3744 716
rect 3620 657 3649 703
rect 3695 657 3744 703
rect 3620 472 3744 657
rect 3844 665 3968 716
rect 3844 525 3873 665
rect 3919 525 3968 665
rect 3844 472 3968 525
rect 4068 703 4192 716
rect 4068 657 4097 703
rect 4143 657 4192 703
rect 4068 472 4192 657
rect 4292 665 4416 716
rect 4292 525 4321 665
rect 4367 525 4416 665
rect 4292 472 4416 525
rect 4516 703 4640 716
rect 4516 657 4545 703
rect 4591 657 4640 703
rect 4516 472 4640 657
rect 4740 665 4864 716
rect 4740 525 4769 665
rect 4815 525 4864 665
rect 4740 472 4864 525
rect 4964 703 5088 716
rect 4964 657 4993 703
rect 5039 657 5088 703
rect 4964 472 5088 657
rect 5188 665 5312 716
rect 5188 525 5217 665
rect 5263 525 5312 665
rect 5188 472 5312 525
rect 5412 703 5536 716
rect 5412 657 5441 703
rect 5487 657 5536 703
rect 5412 472 5536 657
rect 5636 665 5760 716
rect 5636 525 5665 665
rect 5711 525 5760 665
rect 5636 472 5760 525
rect 5860 703 5984 716
rect 5860 657 5889 703
rect 5935 657 5984 703
rect 5860 472 5984 657
rect 6084 665 6208 716
rect 6084 525 6113 665
rect 6159 525 6208 665
rect 6084 472 6208 525
rect 6308 703 6432 716
rect 6308 657 6337 703
rect 6383 657 6432 703
rect 6308 472 6432 657
rect 6532 665 6676 716
rect 6532 525 6581 665
rect 6627 525 6676 665
rect 6532 472 6676 525
rect 6776 693 6864 716
rect 6776 553 6805 693
rect 6851 553 6864 693
rect 6776 472 6864 553
<< mvndiffc >>
rect 273 151 319 197
rect 497 151 543 197
rect 721 151 767 197
rect 945 151 991 197
rect 1169 151 1215 197
rect 1393 151 1439 197
rect 1617 151 1663 197
rect 1841 151 1887 197
rect 2065 151 2111 197
rect 2289 151 2335 197
rect 2549 151 2595 197
rect 2773 151 2819 197
rect 2997 151 3043 197
rect 3221 151 3267 197
rect 3445 151 3491 197
rect 3669 151 3715 197
rect 3893 151 3939 197
rect 4117 151 4163 197
rect 4341 151 4387 197
rect 4565 151 4611 197
rect 4789 151 4835 197
rect 5013 151 5059 197
rect 5237 151 5283 197
rect 5461 151 5507 197
rect 5685 151 5731 197
rect 5909 151 5955 197
rect 6133 151 6179 197
rect 6357 151 6403 197
rect 6581 151 6627 197
rect 6805 151 6851 197
<< mvpdiffc >>
rect 49 657 95 703
rect 273 619 319 665
rect 477 621 523 667
rect 701 619 747 665
rect 925 621 971 667
rect 1149 619 1195 665
rect 1373 621 1419 667
rect 1597 619 1643 665
rect 1821 621 1867 667
rect 2065 619 2111 665
rect 2325 657 2371 703
rect 2549 525 2595 665
rect 2753 657 2799 703
rect 2977 525 3023 665
rect 3201 657 3247 703
rect 3425 525 3471 665
rect 3649 657 3695 703
rect 3873 525 3919 665
rect 4097 657 4143 703
rect 4321 525 4367 665
rect 4545 657 4591 703
rect 4769 525 4815 665
rect 4993 657 5039 703
rect 5217 525 5263 665
rect 5441 657 5487 703
rect 5665 525 5711 665
rect 5889 657 5935 703
rect 6113 525 6159 665
rect 6337 657 6383 703
rect 6581 525 6627 665
rect 6805 553 6851 693
<< polysilicon >>
rect 124 716 224 760
rect 348 716 448 760
rect 572 716 672 760
rect 796 716 896 760
rect 1020 716 1120 760
rect 1244 716 1344 760
rect 1468 716 1568 760
rect 1692 716 1792 760
rect 1916 716 2016 760
rect 2160 716 2260 760
rect 2400 716 2500 760
rect 2624 716 2724 760
rect 2848 716 2948 760
rect 3072 716 3172 760
rect 3296 716 3396 760
rect 3520 716 3620 760
rect 3744 716 3844 760
rect 3968 716 4068 760
rect 4192 716 4292 760
rect 4416 716 4516 760
rect 4640 716 4740 760
rect 4864 716 4964 760
rect 5088 716 5188 760
rect 5312 716 5412 760
rect 5536 716 5636 760
rect 5760 716 5860 760
rect 5984 716 6084 760
rect 6208 716 6308 760
rect 6432 716 6532 760
rect 6676 716 6776 760
rect 124 407 224 552
rect 348 407 448 552
rect 572 407 672 552
rect 796 407 896 552
rect 1020 407 1120 552
rect 1244 407 1344 552
rect 1468 407 1568 552
rect 1692 407 1792 552
rect 1916 407 2016 552
rect 2160 407 2260 552
rect 124 394 2260 407
rect 124 348 137 394
rect 1969 348 2260 394
rect 124 335 2260 348
rect 2400 412 2500 472
rect 2624 412 2724 472
rect 2848 412 2948 472
rect 3072 412 3172 472
rect 3296 412 3396 472
rect 3520 412 3620 472
rect 3744 412 3844 472
rect 3968 412 4068 472
rect 4192 412 4292 472
rect 4416 412 4516 472
rect 4640 412 4740 472
rect 4864 412 4964 472
rect 5088 412 5188 472
rect 5312 412 5412 472
rect 5536 412 5636 472
rect 5760 412 5860 472
rect 5984 412 6084 472
rect 6208 412 6308 472
rect 6432 412 6532 472
rect 6676 412 6776 472
rect 2400 399 6776 412
rect 2400 353 2413 399
rect 4245 353 4783 399
rect 6521 353 6776 399
rect 2400 340 6776 353
rect 348 214 468 335
rect 572 214 692 335
rect 796 214 916 335
rect 1020 214 1140 335
rect 1244 214 1364 335
rect 1468 214 1588 335
rect 1692 214 1812 335
rect 1916 214 2036 335
rect 2400 232 2520 340
rect 2624 232 2744 340
rect 2848 232 2968 340
rect 3072 232 3192 340
rect 3296 232 3416 340
rect 3520 232 3640 340
rect 3744 232 3864 340
rect 3968 232 4088 340
rect 4192 232 4312 340
rect 4416 232 4536 340
rect 4640 232 4760 340
rect 4864 232 4984 340
rect 5088 232 5208 340
rect 5312 232 5432 340
rect 5536 232 5656 340
rect 5760 232 5880 340
rect 5984 232 6104 340
rect 6208 232 6328 340
rect 6432 232 6552 340
rect 6656 232 6776 340
rect 348 94 468 138
rect 572 94 692 138
rect 796 94 916 138
rect 1020 94 1140 138
rect 1244 94 1364 138
rect 1468 94 1588 138
rect 1692 94 1812 138
rect 1916 94 2036 138
rect 2400 94 2520 138
rect 2624 94 2744 138
rect 2848 94 2968 138
rect 3072 94 3192 138
rect 3296 94 3416 138
rect 3520 94 3640 138
rect 3744 94 3864 138
rect 3968 94 4088 138
rect 4192 94 4312 138
rect 4416 94 4536 138
rect 4640 94 4760 138
rect 4864 94 4984 138
rect 5088 94 5208 138
rect 5312 94 5432 138
rect 5536 94 5656 138
rect 5760 94 5880 138
rect 5984 94 6104 138
rect 6208 94 6328 138
rect 6432 94 6552 138
rect 6656 94 6776 138
<< polycontact >>
rect 137 348 1969 394
rect 2413 353 4245 399
rect 4783 353 6521 399
<< metal1 >>
rect 0 724 6944 844
rect 49 703 95 724
rect 49 646 95 657
rect 273 665 319 678
rect 273 552 319 619
rect 477 667 523 724
rect 477 610 523 621
rect 701 665 747 678
rect 701 552 747 619
rect 925 667 971 724
rect 925 610 971 621
rect 1149 665 1195 678
rect 1149 552 1195 619
rect 1373 667 1419 724
rect 1373 610 1419 621
rect 1597 665 1643 678
rect 1597 564 1643 619
rect 1821 667 1867 724
rect 2325 703 2371 724
rect 1821 610 1867 621
rect 2065 665 2111 678
rect 2753 703 2799 724
rect 2325 646 2371 657
rect 2549 665 2595 678
rect 2065 564 2111 619
rect 1597 552 2111 564
rect 273 506 2111 552
rect 126 394 1980 424
rect 126 348 137 394
rect 1969 348 1980 394
rect 2065 399 2111 506
rect 3201 703 3247 724
rect 2753 646 2799 657
rect 2977 665 3023 678
rect 2595 525 2977 600
rect 3649 703 3695 724
rect 3201 646 3247 657
rect 3425 665 3471 678
rect 3023 525 3425 600
rect 4097 703 4143 724
rect 3649 646 3695 657
rect 3873 665 3919 678
rect 3471 525 3873 600
rect 4545 703 4591 724
rect 4097 646 4143 657
rect 4321 665 4367 678
rect 3919 525 4321 600
rect 4993 703 5039 724
rect 4545 646 4591 657
rect 4769 665 4815 678
rect 4367 525 4769 600
rect 5441 703 5487 724
rect 4993 646 5039 657
rect 5217 665 5263 678
rect 4815 525 5217 600
rect 5889 703 5935 724
rect 5441 646 5487 657
rect 5665 665 5711 678
rect 5263 525 5665 600
rect 6337 703 6383 724
rect 5889 646 5935 657
rect 6113 665 6159 678
rect 5711 525 6113 600
rect 6805 693 6851 724
rect 6337 646 6383 657
rect 6581 665 6627 678
rect 6159 525 6581 600
rect 6805 542 6851 553
rect 2549 454 6627 525
rect 2065 353 2413 399
rect 4245 353 4256 399
rect 2065 301 2111 353
rect 4446 307 4626 454
rect 4772 353 4783 399
rect 6521 353 6532 399
rect 273 254 2111 301
rect 273 197 319 254
rect 273 137 319 151
rect 497 197 543 208
rect 497 60 543 151
rect 721 197 767 254
rect 721 137 767 151
rect 945 197 991 208
rect 945 60 991 151
rect 1169 197 1215 254
rect 1169 137 1215 151
rect 1393 197 1439 208
rect 1393 60 1439 151
rect 1617 197 1663 254
rect 1617 137 1663 151
rect 1841 197 1887 208
rect 1841 60 1887 151
rect 2065 197 2111 254
rect 2549 243 6627 307
rect 2065 137 2111 151
rect 2289 197 2335 208
rect 2289 60 2335 151
rect 2549 197 2601 243
rect 2997 197 3043 243
rect 3445 197 3491 243
rect 3893 197 3939 243
rect 4341 197 4387 243
rect 4789 197 4835 243
rect 5237 197 5283 243
rect 5685 197 5731 243
rect 6133 197 6179 243
rect 6581 197 6627 243
rect 2595 151 2601 197
rect 2549 137 2601 151
rect 2762 151 2773 197
rect 2819 151 2830 197
rect 2762 60 2830 151
rect 2997 137 3043 151
rect 3210 151 3221 197
rect 3267 151 3278 197
rect 3210 60 3278 151
rect 3445 137 3491 151
rect 3658 151 3669 197
rect 3715 151 3726 197
rect 3658 60 3726 151
rect 3893 137 3939 151
rect 4106 151 4117 197
rect 4163 151 4174 197
rect 4106 60 4174 151
rect 4341 137 4387 151
rect 4554 151 4565 197
rect 4611 151 4622 197
rect 4554 60 4622 151
rect 4789 137 4835 151
rect 5002 151 5013 197
rect 5059 151 5070 197
rect 5002 60 5070 151
rect 5237 137 5283 151
rect 5450 151 5461 197
rect 5507 151 5518 197
rect 5450 60 5518 151
rect 5685 137 5731 151
rect 5898 151 5909 197
rect 5955 151 5966 197
rect 5898 60 5966 151
rect 6133 137 6179 151
rect 6346 151 6357 197
rect 6403 151 6414 197
rect 6346 60 6414 151
rect 6581 137 6627 151
rect 6805 197 6851 210
rect 6805 60 6851 151
rect 0 -60 6944 60
<< labels >>
flabel metal1 s 0 724 6944 844 0 FreeSans 600 0 0 0 VDD
port 3 nsew power bidirectional abutment
flabel metal1 s 6805 208 6851 210 0 FreeSans 600 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel metal1 s 6581 600 6627 678 0 FreeSans 600 0 0 0 Z
port 2 nsew default output
flabel metal1 s 126 348 1980 424 0 FreeSans 600 0 0 0 I
port 1 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 4 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 6113 600 6159 678 1 Z
port 2 nsew default output
rlabel metal1 s 5665 600 5711 678 1 Z
port 2 nsew default output
rlabel metal1 s 5217 600 5263 678 1 Z
port 2 nsew default output
rlabel metal1 s 4769 600 4815 678 1 Z
port 2 nsew default output
rlabel metal1 s 4321 600 4367 678 1 Z
port 2 nsew default output
rlabel metal1 s 3873 600 3919 678 1 Z
port 2 nsew default output
rlabel metal1 s 3425 600 3471 678 1 Z
port 2 nsew default output
rlabel metal1 s 2977 600 3023 678 1 Z
port 2 nsew default output
rlabel metal1 s 2549 600 2595 678 1 Z
port 2 nsew default output
rlabel metal1 s 2549 454 6627 600 1 Z
port 2 nsew default output
rlabel metal1 s 4446 307 4626 454 1 Z
port 2 nsew default output
rlabel metal1 s 2549 243 6627 307 1 Z
port 2 nsew default output
rlabel metal1 s 6581 137 6627 243 1 Z
port 2 nsew default output
rlabel metal1 s 6133 137 6179 243 1 Z
port 2 nsew default output
rlabel metal1 s 5685 137 5731 243 1 Z
port 2 nsew default output
rlabel metal1 s 5237 137 5283 243 1 Z
port 2 nsew default output
rlabel metal1 s 4789 137 4835 243 1 Z
port 2 nsew default output
rlabel metal1 s 4341 137 4387 243 1 Z
port 2 nsew default output
rlabel metal1 s 3893 137 3939 243 1 Z
port 2 nsew default output
rlabel metal1 s 3445 137 3491 243 1 Z
port 2 nsew default output
rlabel metal1 s 2997 137 3043 243 1 Z
port 2 nsew default output
rlabel metal1 s 2549 137 2601 243 1 Z
port 2 nsew default output
rlabel metal1 s 6805 646 6851 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 6337 646 6383 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 5889 646 5935 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 5441 646 5487 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4993 646 5039 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4545 646 4591 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4097 646 4143 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3649 646 3695 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3201 646 3247 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2753 646 2799 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2325 646 2371 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1821 646 1867 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1373 646 1419 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 925 646 971 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 477 646 523 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 646 95 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 6805 610 6851 646 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1821 610 1867 646 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1373 610 1419 646 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 925 610 971 646 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 477 610 523 646 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 6805 542 6851 610 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 6805 197 6851 208 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2289 197 2335 208 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1841 197 1887 208 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1393 197 1439 208 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 945 197 991 208 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 497 197 543 208 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 6805 60 6851 197 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 6346 60 6414 197 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 5898 60 5966 197 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 5450 60 5518 197 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 5002 60 5070 197 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 4554 60 4622 197 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 4106 60 4174 197 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3658 60 3726 197 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3210 60 3278 197 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2762 60 2830 197 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2289 60 2335 197 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1841 60 1887 197 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1393 60 1439 197 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 945 60 991 197 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 497 60 543 197 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 6944 60 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 6944 784
string GDS_END 815162
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 801190
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
