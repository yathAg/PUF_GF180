magic
tech gf180mcuA
magscale 1 10
timestamp 1698431365
<< obsm1 >>
rect -32 13108 15032 69957
<< metal2 >>
rect 672 65679 748 70000
rect 1193 66054 1269 70000
rect 2066 65990 2142 70000
rect 2277 66954 2353 70000
rect 13734 52998 13810 70000
rect 13880 52862 13956 70000
rect 14026 53238 14102 70000
rect 14172 63950 14248 70000
<< obsm2 >>
rect 0 65619 612 69645
rect 808 65994 1133 69645
rect 1329 65994 2006 69645
rect 808 65930 2006 65994
rect 2202 66894 2217 69645
rect 2413 66894 13674 69645
rect 2202 65930 13674 66894
rect 808 65619 13674 65930
rect 0 52938 13674 65619
rect 0 52802 13820 52938
rect 14308 63890 15000 69645
rect 14162 53178 15000 63890
rect 14016 52802 15000 53178
rect 0 0 15000 52802
<< metal3 >>
rect 0 68400 1864 69678
rect 0 66800 4736 68200
rect 13600 68400 15000 69678
rect 0 65200 1864 66600
rect 14718 66800 15000 68200
rect 0 63600 200 65000
rect 12712 65200 15000 66600
rect 0 62000 200 63400
rect 14800 63600 15000 65000
rect 0 60400 3956 61800
rect 0 58800 3586 60200
rect 14258 62000 15000 63400
rect 10816 60400 15000 61800
rect 0 57200 3947 58600
rect 0 55600 3586 57000
rect 11035 58800 15000 60200
rect 10424 57200 15000 58600
rect 0 54000 3586 55400
rect 0 52400 1814 53800
rect 14718 55600 15000 57000
rect 14718 54000 15000 55400
rect 0 50800 200 52200
rect 14718 52400 15000 53800
rect 0 49200 200 50600
rect 11234 50800 15000 52200
rect 0 46000 200 49000
rect 14800 49200 15000 50600
rect 0 42800 464 45800
rect 11930 46000 15000 49000
rect 0 41200 1963 42600
rect 14718 42800 15000 45800
rect 0 39600 200 41000
rect 14718 41200 15000 42600
rect 0 36400 1808 39400
rect 13273 39600 15000 41000
rect 0 33200 1808 36200
rect 0 30000 1808 33000
rect 0 26800 1808 29800
rect 14718 36400 15000 39400
rect 14718 33200 15000 36200
rect 14718 30000 15000 33000
rect 0 25200 597 26600
rect 14718 26800 15000 29800
rect 0 23600 462 25000
rect 14391 25200 15000 26600
rect 0 20400 200 23400
rect 14487 23600 15000 25000
rect 0 17200 200 20200
rect 0 14000 200 17000
rect 12167 20400 15000 23400
rect 12167 17200 15000 20200
rect 12167 14000 15000 17000
rect 5000 4000 10000 9000
<< obsm3 >>
rect 2224 68560 13240 69678
rect 5096 68040 13240 68560
rect 5096 66960 14358 68040
rect 5096 66440 12352 66960
rect 2224 64840 12352 66440
rect 560 63760 14440 64840
rect 560 62160 13898 63760
rect 4316 60040 10456 62160
rect 3946 58960 10675 60040
rect 4307 56840 10064 58960
rect 3946 53640 14358 56840
rect 2174 52560 14358 53640
rect 2174 52040 10874 52560
rect 560 50440 10874 52040
rect 560 49360 14440 50440
rect 560 46160 11570 49360
rect 824 45640 11570 46160
rect 824 42960 14358 45640
rect 2323 41360 14358 42960
rect 2323 40840 12913 41360
rect 560 39760 12913 40840
rect 2168 39240 12913 39760
rect 2168 26960 14358 39240
rect 2168 26440 14031 26960
rect 957 24840 14031 26440
rect 822 23760 14127 24840
rect 822 23240 11807 23760
rect 560 13640 11807 23240
rect 200 9360 14800 13640
rect 200 3640 4640 9360
rect 10360 3640 14800 9360
rect 200 0 14800 3640
<< labels >>
rlabel metal2 s 13880 52862 13956 70000 6 A
port 1 nsew signal input
rlabel metal2 s 672 65679 748 70000 6 CS
port 2 nsew signal input
rlabel metal3 s 14487 23600 15000 25000 6 DVDD
port 3 nsew power bidirectional
rlabel metal3 s 14718 36400 15000 39400 6 DVDD
port 3 nsew power bidirectional
rlabel metal3 s 14718 33200 15000 36200 6 DVDD
port 3 nsew power bidirectional
rlabel metal3 s 14718 30000 15000 33000 6 DVDD
port 3 nsew power bidirectional
rlabel metal3 s 14718 26800 15000 29800 6 DVDD
port 3 nsew power bidirectional
rlabel metal3 s 14718 42800 15000 45800 6 DVDD
port 3 nsew power bidirectional
rlabel metal3 s 14718 41200 15000 42600 6 DVDD
port 3 nsew power bidirectional
rlabel metal3 s 14718 55600 15000 57000 6 DVDD
port 3 nsew power bidirectional
rlabel metal3 s 14718 54000 15000 55400 6 DVDD
port 3 nsew power bidirectional
rlabel metal3 s 14718 52400 15000 53800 6 DVDD
port 3 nsew power bidirectional
rlabel metal3 s 11035 58800 15000 60200 6 DVDD
port 3 nsew power bidirectional
rlabel metal3 s 14718 66800 15000 68200 6 DVDD
port 3 nsew power bidirectional
rlabel metal3 s 0 66800 4736 68200 6 DVDD
port 3 nsew power bidirectional
rlabel metal3 s 0 58800 3586 60200 6 DVDD
port 3 nsew power bidirectional
rlabel metal3 s 0 52400 1814 53800 6 DVDD
port 3 nsew power bidirectional
rlabel metal3 s 0 54000 3586 55400 6 DVDD
port 3 nsew power bidirectional
rlabel metal3 s 0 55600 3586 57000 6 DVDD
port 3 nsew power bidirectional
rlabel metal3 s 0 41200 1963 42600 6 DVDD
port 3 nsew power bidirectional
rlabel metal3 s 0 42800 464 45800 6 DVDD
port 3 nsew power bidirectional
rlabel metal3 s 0 26800 1808 29800 6 DVDD
port 3 nsew power bidirectional
rlabel metal3 s 0 30000 1808 33000 6 DVDD
port 3 nsew power bidirectional
rlabel metal3 s 0 33200 1808 36200 6 DVDD
port 3 nsew power bidirectional
rlabel metal3 s 0 36400 1808 39400 6 DVDD
port 3 nsew power bidirectional
rlabel metal3 s 0 23600 462 25000 6 DVDD
port 3 nsew power bidirectional
rlabel metal3 s 12167 20400 15000 23400 6 DVSS
port 4 nsew ground bidirectional
rlabel metal3 s 12167 17200 15000 20200 6 DVSS
port 4 nsew ground bidirectional
rlabel metal3 s 12167 14000 15000 17000 6 DVSS
port 4 nsew ground bidirectional
rlabel metal3 s 14391 25200 15000 26600 6 DVSS
port 4 nsew ground bidirectional
rlabel metal3 s 13273 39600 15000 41000 6 DVSS
port 4 nsew ground bidirectional
rlabel metal3 s 11930 46000 15000 49000 6 DVSS
port 4 nsew ground bidirectional
rlabel metal3 s 10424 57200 15000 58600 6 DVSS
port 4 nsew ground bidirectional
rlabel metal3 s 10816 60400 15000 61800 6 DVSS
port 4 nsew ground bidirectional
rlabel metal3 s 12712 65200 15000 66600 6 DVSS
port 4 nsew ground bidirectional
rlabel metal3 s 13600 68400 15000 69678 6 DVSS
port 4 nsew ground bidirectional
rlabel metal3 s 0 68400 1864 69678 6 DVSS
port 4 nsew ground bidirectional
rlabel metal3 s 0 65200 1864 66600 6 DVSS
port 4 nsew ground bidirectional
rlabel metal3 s 0 60400 3956 61800 6 DVSS
port 4 nsew ground bidirectional
rlabel metal3 s 0 57200 3947 58600 6 DVSS
port 4 nsew ground bidirectional
rlabel metal3 s 0 46000 200 49000 6 DVSS
port 4 nsew ground bidirectional
rlabel metal3 s 0 39600 200 41000 6 DVSS
port 4 nsew ground bidirectional
rlabel metal3 s 0 25200 597 26600 6 DVSS
port 4 nsew ground bidirectional
rlabel metal3 s 0 14000 200 17000 6 DVSS
port 4 nsew ground bidirectional
rlabel metal3 s 0 17200 200 20200 6 DVSS
port 4 nsew ground bidirectional
rlabel metal3 s 0 20400 200 23400 6 DVSS
port 4 nsew ground bidirectional
rlabel metal2 s 2277 66954 2353 70000 6 IE
port 5 nsew signal input
rlabel metal2 s 14026 53238 14102 70000 6 OE
port 6 nsew signal input
rlabel metal3 s 5000 4000 10000 9000 6 PAD
port 7 nsew signal bidirectional
rlabel metal2 s 2066 65990 2142 70000 6 PD
port 8 nsew signal input
rlabel metal2 s 1193 66054 1269 70000 6 PU
port 9 nsew signal input
rlabel metal2 s 13734 52998 13810 70000 6 SL
port 10 nsew signal input
rlabel metal3 s 11234 50800 15000 52200 6 VDD
port 11 nsew power bidirectional
rlabel metal3 s 14258 62000 15000 63400 6 VDD
port 11 nsew power bidirectional
rlabel metal3 s 0 62000 200 63400 6 VDD
port 11 nsew power bidirectional
rlabel metal3 s 0 50800 200 52200 6 VDD
port 11 nsew power bidirectional
rlabel metal3 s 14800 49200 15000 50600 6 VSS
port 12 nsew ground bidirectional
rlabel metal3 s 14800 63600 15000 65000 6 VSS
port 12 nsew ground bidirectional
rlabel metal3 s 0 63600 200 65000 6 VSS
port 12 nsew ground bidirectional
rlabel metal3 s 0 49200 200 50600 6 VSS
port 12 nsew ground bidirectional
rlabel metal2 s 14172 63950 14248 70000 6 Y
port 13 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 15000 70000
string LEFclass PAD INOUT
string LEFsite GF_IO_Site
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2011524
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 2009750
<< end >>
