magic
tech gf180mcuB
timestamp 1698431365
<< properties >>
string GDS_END 3222036
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 3220816
<< end >>
