magic
tech gf180mcuA
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 453 1654 1094
<< pwell >>
rect -86 -86 1654 453
<< metal1 >>
rect 0 918 1568 1098
rect 49 710 95 918
rect 477 710 523 918
rect 757 664 803 872
rect 961 710 1007 918
rect 1185 664 1231 872
rect 1409 710 1455 918
rect 757 618 1231 664
rect 161 443 395 511
rect 161 354 306 443
rect 49 90 95 243
rect 1150 375 1231 618
rect 1150 335 1251 375
rect 757 289 1251 335
rect 533 90 579 243
rect 757 175 803 289
rect 981 90 1027 243
rect 1150 175 1251 289
rect 1429 90 1475 243
rect 0 -90 1568 90
<< obsm1 >>
rect 273 664 319 872
rect 273 618 487 664
rect 441 511 487 618
rect 441 443 949 511
rect 441 232 487 443
rect 262 186 487 232
<< labels >>
rlabel metal1 s 161 354 306 443 6 I
port 1 nsew default input
rlabel metal1 s 161 443 395 511 6 I
port 1 nsew default input
rlabel metal1 s 1150 175 1251 289 6 Z
port 2 nsew default output
rlabel metal1 s 757 175 803 289 6 Z
port 2 nsew default output
rlabel metal1 s 757 289 1251 335 6 Z
port 2 nsew default output
rlabel metal1 s 1150 335 1251 375 6 Z
port 2 nsew default output
rlabel metal1 s 1150 375 1231 618 6 Z
port 2 nsew default output
rlabel metal1 s 757 618 1231 664 6 Z
port 2 nsew default output
rlabel metal1 s 1185 664 1231 872 6 Z
port 2 nsew default output
rlabel metal1 s 757 664 803 872 6 Z
port 2 nsew default output
rlabel metal1 s 1409 710 1455 918 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 961 710 1007 918 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 477 710 523 918 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 710 95 918 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 918 1568 1098 6 VDD
port 3 nsew power bidirectional abutment
rlabel nwell s -86 453 1654 1094 6 VNW
port 4 nsew power bidirectional
rlabel pwell s -86 -86 1654 453 6 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 0 -90 1568 90 8 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1429 90 1475 243 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 981 90 1027 243 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 533 90 579 243 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 49 90 95 243 6 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1568 1008
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1395222
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1390928
<< end >>
