magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 453 5350 1094
<< pwell >>
rect -86 -86 5350 453
<< mvnmos >>
rect 124 156 244 274
rect 436 156 556 274
rect 604 156 724 274
rect 828 156 948 274
rect 996 156 1116 274
rect 1400 163 1520 321
rect 1712 156 1832 314
rect 2080 206 2200 324
rect 2304 206 2424 324
rect 2472 206 2592 324
rect 2640 206 2760 324
rect 2864 206 2984 324
rect 3088 206 3208 324
rect 3312 206 3432 324
rect 3540 206 3660 324
rect 3800 124 3920 324
rect 3968 124 4088 324
rect 4336 68 4456 332
rect 4560 68 4680 332
rect 4784 68 4904 332
rect 5008 68 5128 332
<< mvpmos >>
rect 173 652 273 852
rect 436 652 536 852
rect 584 652 684 852
rect 828 652 928 852
rect 976 652 1076 852
rect 1410 580 1510 856
rect 1614 580 1714 856
rect 2028 652 2128 852
rect 2232 652 2332 852
rect 2436 652 2536 852
rect 2640 652 2740 852
rect 2992 652 3092 852
rect 3196 652 3296 852
rect 3400 652 3500 852
rect 3604 652 3704 852
rect 3852 664 3952 940
rect 4056 664 4156 940
rect 4346 573 4446 939
rect 4570 573 4670 939
rect 4776 573 4876 939
rect 5000 573 5100 939
<< mvndiff >>
rect 1312 308 1400 321
rect 36 258 124 274
rect 36 212 49 258
rect 95 212 124 258
rect 36 156 124 212
rect 244 205 436 274
rect 244 159 317 205
rect 363 159 436 205
rect 244 156 436 159
rect 556 156 604 274
rect 724 258 828 274
rect 724 212 753 258
rect 799 212 828 258
rect 724 156 828 212
rect 948 156 996 274
rect 1116 156 1240 274
rect 1312 262 1325 308
rect 1371 262 1400 308
rect 1312 163 1400 262
rect 1520 314 1600 321
rect 1520 163 1712 314
rect 304 146 376 156
rect 1176 130 1240 156
rect 1176 118 1248 130
rect 1580 156 1712 163
rect 1832 296 1920 314
rect 1832 250 1861 296
rect 1907 250 1920 296
rect 1832 156 1920 250
rect 1992 265 2080 324
rect 1992 219 2005 265
rect 2051 219 2080 265
rect 1992 206 2080 219
rect 2200 271 2304 324
rect 2200 225 2229 271
rect 2275 225 2304 271
rect 2200 206 2304 225
rect 2424 206 2472 324
rect 2592 206 2640 324
rect 2760 265 2864 324
rect 2760 219 2789 265
rect 2835 219 2864 265
rect 2760 206 2864 219
rect 2984 311 3088 324
rect 2984 265 3013 311
rect 3059 265 3088 311
rect 2984 206 3088 265
rect 3208 311 3312 324
rect 3208 265 3237 311
rect 3283 265 3312 311
rect 3208 206 3312 265
rect 3432 311 3540 324
rect 3432 265 3465 311
rect 3511 265 3540 311
rect 3432 206 3540 265
rect 3660 265 3800 324
rect 3660 219 3689 265
rect 3735 219 3800 265
rect 3660 206 3800 219
rect 1176 72 1189 118
rect 1235 72 1248 118
rect 1176 59 1248 72
rect 1580 113 1652 156
rect 1580 67 1593 113
rect 1639 67 1652 113
rect 1580 54 1652 67
rect 3720 124 3800 206
rect 3920 124 3968 324
rect 4088 311 4176 324
rect 4088 171 4117 311
rect 4163 171 4176 311
rect 4088 124 4176 171
rect 4248 221 4336 332
rect 4248 81 4261 221
rect 4307 81 4336 221
rect 4248 68 4336 81
rect 4456 319 4560 332
rect 4456 179 4485 319
rect 4531 179 4560 319
rect 4456 68 4560 179
rect 4680 221 4784 332
rect 4680 81 4709 221
rect 4755 81 4784 221
rect 4680 68 4784 81
rect 4904 319 5008 332
rect 4904 179 4933 319
rect 4979 179 5008 319
rect 4904 68 5008 179
rect 5128 221 5216 332
rect 5128 81 5157 221
rect 5203 81 5216 221
rect 5128 68 5216 81
<< mvpdiff >>
rect 85 839 173 852
rect 85 699 98 839
rect 144 699 173 839
rect 85 652 173 699
rect 273 839 436 852
rect 273 699 302 839
rect 348 699 436 839
rect 273 652 436 699
rect 536 652 584 852
rect 684 839 828 852
rect 684 699 753 839
rect 799 699 828 839
rect 684 652 828 699
rect 928 652 976 852
rect 1076 839 1164 852
rect 1076 699 1105 839
rect 1151 699 1164 839
rect 1076 652 1164 699
rect 1322 639 1410 856
rect 1322 593 1335 639
rect 1381 593 1410 639
rect 1322 580 1410 593
rect 1510 834 1614 856
rect 1510 788 1539 834
rect 1585 788 1614 834
rect 1510 580 1614 788
rect 1714 639 1802 856
rect 3764 927 3852 940
rect 3764 881 3777 927
rect 3823 881 3852 927
rect 3764 852 3852 881
rect 1940 839 2028 852
rect 1940 699 1953 839
rect 1999 699 2028 839
rect 1940 652 2028 699
rect 2128 839 2232 852
rect 2128 699 2157 839
rect 2203 699 2232 839
rect 2128 652 2232 699
rect 2332 839 2436 852
rect 2332 699 2361 839
rect 2407 699 2436 839
rect 2332 652 2436 699
rect 2536 747 2640 852
rect 2536 701 2565 747
rect 2611 701 2640 747
rect 2536 652 2640 701
rect 2740 839 2828 852
rect 2740 699 2769 839
rect 2815 699 2828 839
rect 2740 652 2828 699
rect 2904 839 2992 852
rect 2904 699 2917 839
rect 2963 699 2992 839
rect 2904 652 2992 699
rect 3092 839 3196 852
rect 3092 699 3121 839
rect 3167 699 3196 839
rect 3092 652 3196 699
rect 3296 839 3400 852
rect 3296 699 3325 839
rect 3371 699 3400 839
rect 3296 652 3400 699
rect 3500 745 3604 852
rect 3500 699 3529 745
rect 3575 699 3604 745
rect 3500 652 3604 699
rect 3704 664 3852 852
rect 3952 729 4056 940
rect 3952 683 3981 729
rect 4027 683 4056 729
rect 3952 664 4056 683
rect 4156 939 4236 940
rect 4156 839 4346 939
rect 4156 699 4185 839
rect 4231 699 4346 839
rect 4156 664 4346 699
rect 3704 652 3784 664
rect 1714 593 1743 639
rect 1789 593 1802 639
rect 1714 580 1802 593
rect 4266 573 4346 664
rect 4446 839 4570 939
rect 4446 699 4485 839
rect 4531 699 4570 839
rect 4446 573 4570 699
rect 4670 839 4776 939
rect 4670 699 4699 839
rect 4745 699 4776 839
rect 4670 573 4776 699
rect 4876 839 5000 939
rect 4876 699 4905 839
rect 4951 699 5000 839
rect 4876 573 5000 699
rect 5100 839 5188 939
rect 5100 699 5129 839
rect 5175 699 5188 839
rect 5100 573 5188 699
<< mvndiffc >>
rect 49 212 95 258
rect 317 159 363 205
rect 753 212 799 258
rect 1325 262 1371 308
rect 1861 250 1907 296
rect 2005 219 2051 265
rect 2229 225 2275 271
rect 2789 219 2835 265
rect 3013 265 3059 311
rect 3237 265 3283 311
rect 3465 265 3511 311
rect 3689 219 3735 265
rect 1189 72 1235 118
rect 1593 67 1639 113
rect 4117 171 4163 311
rect 4261 81 4307 221
rect 4485 179 4531 319
rect 4709 81 4755 221
rect 4933 179 4979 319
rect 5157 81 5203 221
<< mvpdiffc >>
rect 98 699 144 839
rect 302 699 348 839
rect 753 699 799 839
rect 1105 699 1151 839
rect 1335 593 1381 639
rect 1539 788 1585 834
rect 3777 881 3823 927
rect 1953 699 1999 839
rect 2157 699 2203 839
rect 2361 699 2407 839
rect 2565 701 2611 747
rect 2769 699 2815 839
rect 2917 699 2963 839
rect 3121 699 3167 839
rect 3325 699 3371 839
rect 3529 699 3575 745
rect 3981 683 4027 729
rect 4185 699 4231 839
rect 1743 593 1789 639
rect 4485 699 4531 839
rect 4699 699 4745 839
rect 4905 699 4951 839
rect 5129 699 5175 839
<< polysilicon >>
rect 173 944 1076 984
rect 173 852 273 944
rect 436 852 536 896
rect 584 852 684 896
rect 828 852 928 896
rect 976 852 1076 944
rect 1614 944 3296 984
rect 1410 856 1510 900
rect 1614 856 1714 944
rect 173 559 273 652
rect 124 547 273 559
rect 436 547 536 652
rect 124 501 178 547
rect 224 501 244 547
rect 124 274 244 501
rect 436 501 449 547
rect 495 501 536 547
rect 436 318 536 501
rect 584 547 684 652
rect 584 501 597 547
rect 643 501 684 547
rect 584 488 684 501
rect 828 547 928 652
rect 976 608 1076 652
rect 2028 852 2128 896
rect 2232 852 2332 944
rect 2436 852 2536 896
rect 2640 852 2740 896
rect 2992 852 3092 896
rect 3196 852 3296 944
rect 3852 940 3952 984
rect 4056 940 4156 984
rect 3400 852 3500 896
rect 3604 852 3704 896
rect 4346 939 4446 983
rect 4570 939 4670 983
rect 4776 939 4876 983
rect 5000 939 5100 983
rect 828 501 841 547
rect 887 501 928 547
rect 828 318 928 501
rect 996 539 1116 552
rect 996 493 1029 539
rect 1075 493 1116 539
rect 436 274 556 318
rect 604 274 724 318
rect 828 274 948 318
rect 996 274 1116 493
rect 1410 547 1510 580
rect 1410 501 1423 547
rect 1469 501 1510 547
rect 1410 365 1510 501
rect 1614 547 1714 580
rect 1614 501 1627 547
rect 1673 501 1714 547
rect 1614 452 1714 501
rect 2028 560 2128 652
rect 2232 608 2332 652
rect 2436 608 2536 652
rect 2028 547 2424 560
rect 2028 501 2041 547
rect 2087 501 2424 547
rect 2028 488 2424 501
rect 1614 380 1832 452
rect 1400 321 1520 365
rect 1712 314 1832 380
rect 2304 403 2424 488
rect 2080 324 2200 368
rect 2304 357 2345 403
rect 2391 357 2424 403
rect 2304 324 2424 357
rect 2472 472 2536 608
rect 2472 460 2592 472
rect 2472 414 2485 460
rect 2531 414 2592 460
rect 2472 324 2592 414
rect 2640 368 2740 652
rect 2992 608 3092 652
rect 3196 608 3296 652
rect 2992 565 3032 608
rect 2864 552 3032 565
rect 2864 506 2897 552
rect 2943 506 3032 552
rect 2864 493 3032 506
rect 3088 547 3208 560
rect 3088 501 3121 547
rect 3167 501 3208 547
rect 2640 324 2760 368
rect 2864 324 2984 493
rect 3088 324 3208 501
rect 3256 424 3296 608
rect 3400 547 3500 652
rect 3604 608 3704 652
rect 3852 620 3952 664
rect 4056 620 4156 664
rect 3604 560 3660 608
rect 3852 560 3900 620
rect 4056 566 4128 620
rect 3400 501 3413 547
rect 3459 501 3500 547
rect 3400 488 3500 501
rect 3560 547 3660 560
rect 3560 501 3601 547
rect 3647 501 3660 547
rect 3256 384 3432 424
rect 3312 324 3432 384
rect 3560 368 3660 501
rect 3719 547 3900 560
rect 3719 501 3732 547
rect 3778 501 3900 547
rect 3719 500 3900 501
rect 3968 560 4128 566
rect 3968 514 4069 560
rect 4115 514 4128 560
rect 3968 501 4128 514
rect 3719 488 3840 500
rect 3540 324 3660 368
rect 3800 368 3840 488
rect 3800 324 3920 368
rect 3968 324 4088 501
rect 4346 464 4446 573
rect 4570 464 4670 573
rect 4776 464 4876 573
rect 5000 464 5100 573
rect 4346 456 5100 464
rect 4147 443 5100 456
rect 4147 397 4160 443
rect 4206 397 5100 443
rect 4147 392 5100 397
rect 4147 384 4218 392
rect 4336 332 4456 392
rect 4560 332 4680 392
rect 4784 332 4904 392
rect 5008 376 5100 392
rect 5008 332 5128 376
rect 124 64 244 156
rect 436 112 556 156
rect 604 64 724 156
rect 828 112 948 156
rect 996 112 1116 156
rect 1400 119 1520 163
rect 124 24 724 64
rect 1712 96 1832 156
rect 2080 96 2200 206
rect 2304 162 2424 206
rect 2472 162 2592 206
rect 1712 24 2200 96
rect 2640 64 2760 206
rect 2864 162 2984 206
rect 3088 162 3208 206
rect 3312 162 3432 206
rect 3540 162 3660 206
rect 3800 64 3920 124
rect 3968 80 4088 124
rect 2640 24 3920 64
rect 4336 24 4456 68
rect 4560 24 4680 68
rect 4784 24 4904 68
rect 5008 24 5128 68
<< polycontact >>
rect 178 501 224 547
rect 449 501 495 547
rect 597 501 643 547
rect 841 501 887 547
rect 1029 493 1075 539
rect 1423 501 1469 547
rect 1627 501 1673 547
rect 2041 501 2087 547
rect 2345 357 2391 403
rect 2485 414 2531 460
rect 2897 506 2943 552
rect 3121 501 3167 547
rect 3413 501 3459 547
rect 3601 501 3647 547
rect 3732 501 3778 547
rect 4069 514 4115 560
rect 4160 397 4206 443
<< metal1 >>
rect 0 927 5264 1098
rect 0 918 3777 927
rect 98 839 144 850
rect 98 639 144 699
rect 302 839 348 918
rect 302 688 348 699
rect 753 839 799 850
rect 753 642 799 699
rect 1105 839 1151 918
rect 1528 834 1596 918
rect 1528 788 1539 834
rect 1585 788 1596 834
rect 1953 839 1999 850
rect 1105 688 1151 699
rect 1197 699 1953 742
rect 1197 696 1999 699
rect 1197 642 1243 696
rect 1953 688 1999 696
rect 2157 839 2203 850
rect 98 593 643 639
rect 753 596 1243 642
rect 1743 639 1789 650
rect 1324 593 1335 639
rect 1381 593 1572 639
rect 597 547 643 593
rect 142 501 178 547
rect 224 501 235 547
rect 142 354 235 501
rect 366 501 449 547
rect 495 501 506 547
rect 366 354 506 501
rect 597 420 643 501
rect 702 501 841 547
rect 887 501 898 547
rect 702 466 898 501
rect 1029 539 1075 550
rect 1526 547 1572 593
rect 1743 547 1789 593
rect 2157 588 2203 699
rect 2361 839 2407 850
rect 2361 644 2407 699
rect 2565 747 2611 918
rect 2565 690 2611 701
rect 2769 839 2815 850
rect 2769 644 2815 699
rect 2917 839 2963 918
rect 3823 918 5264 927
rect 3777 870 3823 881
rect 2917 688 2963 699
rect 3121 839 3167 850
rect 3121 650 3167 699
rect 2361 598 2815 644
rect 3013 604 3167 650
rect 3325 849 3690 850
rect 3325 839 3736 849
rect 3371 824 3736 839
rect 4185 839 4231 918
rect 3849 824 4119 832
rect 3371 804 4119 824
rect 3680 786 4119 804
rect 3680 778 3875 786
rect 3325 623 3371 699
rect 2157 552 2274 588
rect 1029 420 1075 493
rect 597 374 1075 420
rect 1374 501 1423 547
rect 1469 501 1480 547
rect 1526 501 1627 547
rect 1673 501 1684 547
rect 1743 501 2041 547
rect 2087 501 2098 547
rect 2157 542 2897 552
rect 2229 506 2897 542
rect 2943 506 2954 552
rect 597 308 643 374
rect 1374 354 1480 501
rect 1638 308 1684 501
rect 49 262 643 308
rect 49 258 95 262
rect 753 258 799 269
rect 1314 262 1325 308
rect 1371 262 1684 308
rect 1861 296 1907 501
rect 49 201 95 212
rect 317 205 363 216
rect 1861 239 1907 250
rect 2005 265 2051 276
rect 799 216 1293 221
rect 799 212 1816 216
rect 753 193 1816 212
rect 2005 193 2051 219
rect 2229 271 2275 506
rect 3013 460 3059 604
rect 3237 577 3371 623
rect 3505 745 3575 756
rect 3505 699 3529 745
rect 3505 688 3575 699
rect 3981 729 4027 740
rect 2474 414 2485 460
rect 2531 414 3059 460
rect 2334 357 2345 403
rect 2391 368 2402 403
rect 2391 357 2967 368
rect 2334 322 2967 357
rect 2229 214 2275 225
rect 2789 265 2835 276
rect 753 175 2051 193
rect 1272 170 2051 175
rect 317 90 363 159
rect 1771 147 2051 170
rect 1189 118 1235 129
rect 0 72 1189 90
rect 1593 113 1639 124
rect 1235 72 1593 90
rect 0 67 1593 72
rect 2789 90 2835 219
rect 2921 208 2967 322
rect 3013 311 3059 414
rect 3013 254 3059 265
rect 3121 547 3167 558
rect 3121 208 3167 501
rect 3237 311 3283 577
rect 3413 547 3459 558
rect 3413 414 3459 501
rect 3237 254 3283 265
rect 3373 368 3459 414
rect 3373 208 3419 368
rect 3505 322 3551 688
rect 3981 650 4027 683
rect 3601 631 4027 650
rect 3601 604 4023 631
rect 3601 547 3647 604
rect 3601 490 3647 501
rect 3726 547 3778 558
rect 3726 501 3732 547
rect 3726 354 3778 501
rect 3977 443 4023 604
rect 4073 571 4119 786
rect 4185 688 4231 699
rect 4485 839 4531 850
rect 4069 560 4119 571
rect 4115 514 4119 560
rect 4069 503 4119 514
rect 3977 397 4160 443
rect 4206 397 4217 443
rect 3465 311 3551 322
rect 3511 265 3551 311
rect 4117 311 4163 397
rect 3465 254 3551 265
rect 3689 265 3735 276
rect 2921 162 3419 208
rect 3689 90 3735 219
rect 4485 324 4531 699
rect 4699 839 4745 918
rect 4699 688 4745 699
rect 4846 839 4979 850
rect 4846 699 4905 839
rect 4951 699 4979 839
rect 4846 324 4979 699
rect 5129 839 5175 918
rect 5129 688 5175 699
rect 4485 319 4979 324
rect 4117 160 4163 171
rect 4261 221 4307 232
rect 1639 81 4261 90
rect 4531 278 4933 319
rect 4846 242 4933 278
rect 4485 168 4531 179
rect 4709 221 4755 232
rect 4307 81 4709 90
rect 4933 168 4979 179
rect 5157 221 5203 232
rect 4755 81 5157 90
rect 5203 81 5264 90
rect 1639 67 5264 81
rect 0 -90 5264 67
<< labels >>
flabel metal1 s 1374 354 1480 547 0 FreeSans 200 0 0 0 CLK
port 5 nsew clock input
flabel metal1 s 702 466 898 547 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 4846 324 4979 850 0 FreeSans 200 0 0 0 Q
port 6 nsew default output
flabel metal1 s 3726 354 3778 558 0 FreeSans 200 0 0 0 RN
port 2 nsew default input
flabel metal1 s 142 354 235 547 0 FreeSans 200 0 0 0 SE
port 3 nsew default input
flabel metal1 s 366 354 506 547 0 FreeSans 200 0 0 0 SI
port 4 nsew default input
flabel metal1 s 0 918 5264 1098 0 FreeSans 200 0 0 0 VDD
port 7 nsew power bidirectional abutment
flabel metal1 s 3689 232 3735 276 0 FreeSans 200 0 0 0 VSS
port 10 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 8 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 9 nsew ground bidirectional
rlabel metal1 s 4485 324 4531 850 1 Q
port 6 nsew default output
rlabel metal1 s 4485 278 4979 324 1 Q
port 6 nsew default output
rlabel metal1 s 4846 242 4979 278 1 Q
port 6 nsew default output
rlabel metal1 s 4485 242 4531 278 1 Q
port 6 nsew default output
rlabel metal1 s 4933 168 4979 242 1 Q
port 6 nsew default output
rlabel metal1 s 4485 168 4531 242 1 Q
port 6 nsew default output
rlabel metal1 s 5129 870 5175 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4699 870 4745 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4185 870 4231 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3777 870 3823 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2917 870 2963 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2565 870 2611 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1528 870 1596 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1105 870 1151 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 302 870 348 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5129 788 5175 870 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4699 788 4745 870 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4185 788 4231 870 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2917 788 2963 870 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2565 788 2611 870 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1528 788 1596 870 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1105 788 1151 870 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 302 788 348 870 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5129 690 5175 788 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4699 690 4745 788 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4185 690 4231 788 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2917 690 2963 788 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2565 690 2611 788 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1105 690 1151 788 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 302 690 348 788 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5129 688 5175 690 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4699 688 4745 690 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4185 688 4231 690 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2917 688 2963 690 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1105 688 1151 690 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 302 688 348 690 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2789 232 2835 276 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 5157 216 5203 232 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 4709 216 4755 232 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 4261 216 4307 232 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 3689 216 3735 232 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 2789 216 2835 232 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 5157 129 5203 216 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 4709 129 4755 216 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 4261 129 4307 216 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 3689 129 3735 216 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 2789 129 2835 216 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 317 129 363 216 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 5157 124 5203 129 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 4709 124 4755 129 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 4261 124 4307 129 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 3689 124 3735 129 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 2789 124 2835 129 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 1189 124 1235 129 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 317 124 363 129 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 5157 90 5203 124 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 4709 90 4755 124 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 4261 90 4307 124 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 3689 90 3735 124 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 2789 90 2835 124 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 1593 90 1639 124 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 1189 90 1235 124 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 317 90 363 124 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 5264 90 1 VSS
port 10 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 5264 1008
string GDS_END 367660
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 355452
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
