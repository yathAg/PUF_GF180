magic
tech gf180mcuB
magscale 1 5
timestamp 1698431365
use 018SRAM_strap1_bndry_64x8m81  018SRAM_strap1_bndry_64x8m81_0
timestamp 1698431365
transform 1 0 0 0 -1 460
box -34 -34 334 484
use 018SRAM_strap1_bndry_64x8m81  018SRAM_strap1_bndry_64x8m81_1
timestamp 1698431365
transform 1 0 0 0 1 460
box -34 -34 334 484
<< properties >>
string GDS_END 1001350
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 1001236
<< end >>
