magic
tech gf180mcuA
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 453 5014 1094
<< pwell >>
rect -86 -86 5014 453
<< mvnmos >>
rect 124 156 244 272
rect 348 156 468 272
rect 516 156 636 272
rect 740 156 860 272
rect 908 156 1028 272
rect 1320 175 1440 333
rect 1632 175 1752 333
rect 2000 217 2120 333
rect 2224 217 2344 333
rect 2392 217 2512 333
rect 2692 217 2812 333
rect 2916 217 3036 333
rect 3140 217 3260 333
rect 3400 69 3520 333
rect 3624 69 3744 333
rect 3992 69 4112 333
rect 4216 69 4336 333
rect 4440 69 4560 333
rect 4664 69 4784 333
<< mvpmos >>
rect 200 652 300 852
rect 404 652 504 852
rect 552 652 652 852
rect 756 652 856 852
rect 918 652 1018 852
rect 1448 573 1548 849
rect 1652 573 1752 849
rect 2133 652 2233 852
rect 2340 652 2440 852
rect 2488 652 2588 852
rect 2692 652 2792 852
rect 2926 652 3026 852
rect 3140 652 3240 852
rect 3400 573 3500 939
rect 3618 573 3718 939
rect 4022 573 4122 939
rect 4226 573 4326 939
rect 4432 573 4532 939
rect 4657 573 4757 939
<< mvndiff >>
rect 1232 320 1320 333
rect 1232 274 1245 320
rect 1291 274 1320 320
rect 36 215 124 272
rect 36 169 49 215
rect 95 169 124 215
rect 36 156 124 169
rect 244 215 348 272
rect 244 169 273 215
rect 319 169 348 215
rect 244 156 348 169
rect 468 156 516 272
rect 636 215 740 272
rect 636 169 665 215
rect 711 169 740 215
rect 636 156 740 169
rect 860 156 908 272
rect 1028 156 1160 272
rect 1232 175 1320 274
rect 1440 175 1632 333
rect 1752 320 1840 333
rect 1752 274 1781 320
rect 1827 274 1840 320
rect 1752 175 1840 274
rect 1912 276 2000 333
rect 1912 230 1925 276
rect 1971 230 2000 276
rect 1912 217 2000 230
rect 2120 320 2224 333
rect 2120 274 2149 320
rect 2195 274 2224 320
rect 2120 217 2224 274
rect 2344 217 2392 333
rect 2512 217 2692 333
rect 2812 320 2916 333
rect 2812 274 2841 320
rect 2887 274 2916 320
rect 2812 217 2916 274
rect 3036 320 3140 333
rect 3036 274 3065 320
rect 3111 274 3140 320
rect 3036 217 3140 274
rect 3260 217 3400 333
rect 1088 114 1160 156
rect 1088 68 1101 114
rect 1147 68 1160 114
rect 1088 55 1160 68
rect 1500 114 1572 175
rect 1500 68 1513 114
rect 1559 68 1572 114
rect 1500 55 1572 68
rect 2572 127 2632 217
rect 2572 119 2643 127
rect 2571 114 2643 119
rect 2571 68 2584 114
rect 2630 68 2643 114
rect 3320 69 3400 217
rect 3520 268 3624 333
rect 3520 128 3549 268
rect 3595 128 3624 268
rect 3520 69 3624 128
rect 3744 309 3832 333
rect 3744 169 3773 309
rect 3819 169 3832 309
rect 3744 69 3832 169
rect 3904 309 3992 333
rect 3904 169 3917 309
rect 3963 169 3992 309
rect 3904 69 3992 169
rect 4112 320 4216 333
rect 4112 180 4141 320
rect 4187 180 4216 320
rect 4112 69 4216 180
rect 4336 222 4440 333
rect 4336 82 4365 222
rect 4411 82 4440 222
rect 4336 69 4440 82
rect 4560 320 4664 333
rect 4560 180 4589 320
rect 4635 180 4664 320
rect 4560 69 4664 180
rect 4784 222 4872 333
rect 4784 82 4813 222
rect 4859 82 4872 222
rect 4784 69 4872 82
rect 2571 55 2643 68
<< mvpdiff >>
rect 112 839 200 852
rect 112 699 125 839
rect 171 699 200 839
rect 112 652 200 699
rect 300 839 404 852
rect 300 699 329 839
rect 375 699 404 839
rect 300 652 404 699
rect 504 652 552 852
rect 652 839 756 852
rect 652 699 681 839
rect 727 699 756 839
rect 652 652 756 699
rect 856 652 918 852
rect 1018 838 1106 852
rect 3320 852 3400 939
rect 1018 792 1047 838
rect 1093 792 1106 838
rect 1018 652 1106 792
rect 1360 632 1448 849
rect 1360 586 1373 632
rect 1419 586 1448 632
rect 1360 573 1448 586
rect 1548 827 1652 849
rect 1548 781 1577 827
rect 1623 781 1652 827
rect 1548 573 1652 781
rect 1752 632 1840 849
rect 2045 746 2133 852
rect 2045 700 2058 746
rect 2104 700 2133 746
rect 2045 652 2133 700
rect 2233 839 2340 852
rect 2233 699 2265 839
rect 2311 699 2340 839
rect 2233 652 2340 699
rect 2440 652 2488 852
rect 2588 839 2692 852
rect 2588 699 2617 839
rect 2663 699 2692 839
rect 2588 652 2692 699
rect 2792 839 2926 852
rect 2792 699 2841 839
rect 2887 699 2926 839
rect 2792 652 2926 699
rect 3026 839 3140 852
rect 3026 699 3065 839
rect 3111 699 3140 839
rect 3026 652 3140 699
rect 3240 652 3400 852
rect 1752 586 1781 632
rect 1827 586 1840 632
rect 1752 573 1840 586
rect 3320 573 3400 652
rect 3500 861 3618 939
rect 3500 721 3529 861
rect 3575 721 3618 861
rect 3500 573 3618 721
rect 3718 839 3806 939
rect 3718 699 3747 839
rect 3793 699 3806 839
rect 3718 573 3806 699
rect 3934 926 4022 939
rect 3934 786 3947 926
rect 3993 786 4022 926
rect 3934 573 4022 786
rect 4122 839 4226 939
rect 4122 699 4151 839
rect 4197 699 4226 839
rect 4122 573 4226 699
rect 4326 926 4432 939
rect 4326 786 4355 926
rect 4401 786 4432 926
rect 4326 573 4432 786
rect 4532 839 4657 939
rect 4532 699 4561 839
rect 4607 699 4657 839
rect 4532 573 4657 699
rect 4757 926 4845 939
rect 4757 786 4786 926
rect 4832 786 4845 926
rect 4757 573 4845 786
<< mvndiffc >>
rect 1245 274 1291 320
rect 49 169 95 215
rect 273 169 319 215
rect 665 169 711 215
rect 1781 274 1827 320
rect 1925 230 1971 276
rect 2149 274 2195 320
rect 2841 274 2887 320
rect 3065 274 3111 320
rect 1101 68 1147 114
rect 1513 68 1559 114
rect 2584 68 2630 114
rect 3549 128 3595 268
rect 3773 169 3819 309
rect 3917 169 3963 309
rect 4141 180 4187 320
rect 4365 82 4411 222
rect 4589 180 4635 320
rect 4813 82 4859 222
<< mvpdiffc >>
rect 125 699 171 839
rect 329 699 375 839
rect 681 699 727 839
rect 1047 792 1093 838
rect 1373 586 1419 632
rect 1577 781 1623 827
rect 2058 700 2104 746
rect 2265 699 2311 839
rect 2617 699 2663 839
rect 2841 699 2887 839
rect 3065 699 3111 839
rect 1781 586 1827 632
rect 3529 721 3575 861
rect 3747 699 3793 839
rect 3947 786 3993 926
rect 4151 699 4197 839
rect 4355 786 4401 926
rect 4561 699 4607 839
rect 4786 786 4832 926
<< polysilicon >>
rect 200 944 856 984
rect 200 852 300 944
rect 404 852 504 896
rect 552 852 652 896
rect 756 852 856 944
rect 1652 944 3026 984
rect 918 852 1018 896
rect 1448 849 1548 893
rect 1652 849 1752 944
rect 2133 852 2233 896
rect 2340 852 2440 944
rect 2488 852 2588 896
rect 2692 852 2792 896
rect 2926 852 3026 944
rect 3400 939 3500 983
rect 3618 939 3718 983
rect 4022 939 4122 983
rect 4226 939 4326 983
rect 4432 939 4532 983
rect 4657 939 4757 983
rect 3140 852 3240 896
rect 200 476 300 652
rect 404 476 504 652
rect 24 463 300 476
rect 24 417 37 463
rect 83 419 300 463
rect 348 463 504 476
rect 83 417 244 419
rect 24 404 244 417
rect 124 272 244 404
rect 348 417 361 463
rect 407 443 504 463
rect 552 463 652 652
rect 756 608 856 652
rect 918 476 1018 652
rect 2133 608 2233 652
rect 2340 608 2440 652
rect 1448 476 1548 573
rect 1652 476 1752 573
rect 407 417 468 443
rect 348 272 468 417
rect 552 417 565 463
rect 611 436 652 463
rect 908 463 1018 476
rect 611 417 860 436
rect 552 364 860 417
rect 516 272 636 316
rect 740 272 860 364
rect 908 417 921 463
rect 967 417 1018 463
rect 908 316 1018 417
rect 1066 463 1548 476
rect 1066 417 1079 463
rect 1125 436 1548 463
rect 1632 463 1752 476
rect 1125 417 1440 436
rect 1066 404 1440 417
rect 1320 333 1440 404
rect 1632 417 1645 463
rect 1691 417 1752 463
rect 1632 333 1752 417
rect 2160 476 2233 608
rect 2160 463 2344 476
rect 2160 417 2173 463
rect 2219 417 2344 463
rect 2488 463 2588 652
rect 2488 461 2529 463
rect 2160 404 2344 417
rect 2000 333 2120 377
rect 2224 333 2344 404
rect 2392 417 2529 461
rect 2575 417 2588 463
rect 2392 393 2588 417
rect 2692 463 2792 652
rect 2692 417 2705 463
rect 2751 417 2792 463
rect 2926 465 3026 652
rect 3140 572 3240 652
rect 3140 526 3168 572
rect 3214 526 3240 572
rect 3140 513 3240 526
rect 2926 425 3260 465
rect 2392 333 2512 393
rect 2692 377 2792 417
rect 2692 333 2812 377
rect 2916 333 3036 377
rect 3140 333 3260 425
rect 3400 463 3500 573
rect 3400 417 3441 463
rect 3487 417 3500 463
rect 3400 377 3500 417
rect 3618 463 3718 573
rect 4022 476 4122 573
rect 3618 417 3631 463
rect 3677 417 3718 463
rect 3618 406 3718 417
rect 3624 377 3718 406
rect 3992 465 4122 476
rect 4226 465 4326 573
rect 4432 465 4532 573
rect 4657 465 4757 573
rect 3992 463 4757 465
rect 3992 417 4005 463
rect 4051 425 4757 463
rect 4051 417 4112 425
rect 3400 333 3520 377
rect 3624 333 3744 377
rect 3992 333 4112 417
rect 4216 333 4336 425
rect 4440 333 4560 425
rect 4664 377 4757 425
rect 4664 333 4784 377
rect 908 272 1028 316
rect 124 64 244 156
rect 348 112 468 156
rect 516 64 636 156
rect 740 112 860 156
rect 908 112 1028 156
rect 1320 131 1440 175
rect 124 24 636 64
rect 1632 96 1752 175
rect 2000 96 2120 217
rect 2224 184 2344 217
rect 2224 138 2285 184
rect 2331 138 2344 184
rect 2392 173 2512 217
rect 2224 125 2344 138
rect 2692 173 2812 217
rect 2916 184 3036 217
rect 2916 138 2957 184
rect 3003 138 3036 184
rect 3140 173 3260 217
rect 2916 125 3036 138
rect 1632 24 2120 96
rect 3400 25 3520 69
rect 3624 25 3744 69
rect 3992 25 4112 69
rect 4216 25 4336 69
rect 4440 25 4560 69
rect 4664 25 4784 69
<< polycontact >>
rect 37 417 83 463
rect 361 417 407 463
rect 565 417 611 463
rect 921 417 967 463
rect 1079 417 1125 463
rect 1645 417 1691 463
rect 2173 417 2219 463
rect 2529 417 2575 463
rect 2705 417 2751 463
rect 3168 526 3214 572
rect 3441 417 3487 463
rect 3631 417 3677 463
rect 4005 417 4051 463
rect 2285 138 2331 184
rect 2957 138 3003 184
<< metal1 >>
rect 0 926 4928 1098
rect 0 918 3947 926
rect 125 839 171 850
rect 125 642 171 699
rect 329 839 375 918
rect 329 688 375 699
rect 681 839 727 850
rect 1047 838 1093 918
rect 2265 839 2311 850
rect 1093 792 1577 827
rect 1047 781 1577 792
rect 1623 781 1634 827
rect 2058 746 2104 757
rect 727 700 2058 735
rect 727 699 2104 700
rect 681 689 2104 699
rect 681 688 727 689
rect 125 596 611 642
rect 30 463 83 542
rect 30 417 37 463
rect 30 354 83 417
rect 142 474 194 542
rect 142 463 407 474
rect 142 417 361 463
rect 142 406 407 417
rect 565 463 611 596
rect 1373 632 1691 643
rect 1419 586 1691 632
rect 1373 575 1691 586
rect 142 354 194 406
rect 565 307 611 417
rect 814 474 866 542
rect 814 463 967 474
rect 814 417 921 463
rect 814 406 967 417
rect 1038 463 1125 542
rect 1038 417 1079 463
rect 814 354 866 406
rect 1038 354 1125 417
rect 1645 463 1691 575
rect 1645 331 1691 417
rect 49 261 611 307
rect 1245 320 1691 331
rect 1291 274 1691 320
rect 1245 263 1691 274
rect 1781 632 1827 643
rect 1781 474 1827 586
rect 1781 463 2219 474
rect 1781 417 2173 463
rect 1781 406 2219 417
rect 1781 320 1827 406
rect 2265 360 2311 699
rect 2617 839 2663 918
rect 3529 861 3575 918
rect 2617 688 2663 699
rect 2841 839 2887 850
rect 2841 566 2887 699
rect 2529 520 2887 566
rect 2529 463 2575 520
rect 2529 406 2575 417
rect 2705 463 2751 474
rect 2705 360 2751 417
rect 2265 331 2751 360
rect 2149 320 2751 331
rect 1781 263 1827 274
rect 1925 276 1971 287
rect 49 215 95 261
rect 2195 314 2751 320
rect 2841 320 2887 520
rect 2195 274 2308 314
rect 2149 263 2308 274
rect 2841 263 2887 274
rect 3065 839 3111 850
rect 3529 710 3575 721
rect 3747 839 3793 850
rect 3065 664 3111 699
rect 3993 918 4355 926
rect 3947 775 3993 786
rect 4141 839 4197 850
rect 3065 618 3579 664
rect 3065 320 3111 618
rect 3065 263 3111 274
rect 3157 526 3168 572
rect 3214 526 3225 572
rect 665 217 711 226
rect 1925 217 1971 230
rect 3157 217 3225 526
rect 3441 463 3487 474
rect 3533 463 3579 618
rect 3747 474 3793 699
rect 4141 699 4151 839
rect 4401 918 4786 926
rect 4355 775 4401 786
rect 4561 839 4607 850
rect 4197 699 4561 729
rect 4832 918 4928 926
rect 4786 775 4832 786
rect 4141 683 4607 699
rect 3747 463 4051 474
rect 3533 417 3631 463
rect 3677 417 3688 463
rect 3747 417 4005 463
rect 3441 371 3487 417
rect 3747 406 4051 417
rect 4141 430 4187 683
rect 3747 371 3819 406
rect 3441 325 3819 371
rect 3773 309 3819 325
rect 4141 384 4562 430
rect 4141 320 4187 384
rect 665 215 1971 217
rect 49 158 95 169
rect 262 169 273 215
rect 319 169 330 215
rect 262 90 330 169
rect 711 171 1971 215
rect 2274 184 3225 217
rect 665 158 711 169
rect 2274 138 2285 184
rect 2331 171 2957 184
rect 2331 138 2342 171
rect 2946 138 2957 171
rect 3003 138 3225 184
rect 3549 268 3595 279
rect 3773 158 3819 169
rect 3917 309 3963 320
rect 4510 331 4562 384
rect 4510 320 4635 331
rect 4510 242 4589 320
rect 4141 169 4187 180
rect 4365 222 4411 233
rect 1101 114 1147 125
rect 0 68 1101 90
rect 1513 114 1559 125
rect 1147 68 1513 90
rect 2584 114 2630 125
rect 1559 68 2584 90
rect 3549 90 3595 128
rect 3917 90 3963 169
rect 2630 82 4365 90
rect 4589 169 4635 180
rect 4813 222 4859 233
rect 4411 82 4813 90
rect 4859 82 4928 90
rect 2630 68 4928 82
rect 0 -90 4928 68
<< labels >>
flabel metal1 s 1038 354 1125 542 0 FreeSans 200 0 0 0 CLK
port 4 nsew clock input
flabel metal1 s 814 474 866 542 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 4561 729 4607 850 0 FreeSans 200 0 0 0 Q
port 5 nsew default output
flabel metal1 s 30 354 83 542 0 FreeSans 200 0 0 0 SE
port 2 nsew default input
flabel metal1 s 142 474 194 542 0 FreeSans 200 0 0 0 SI
port 3 nsew default input
flabel metal1 s 0 918 4928 1098 0 FreeSans 200 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 3917 279 3963 320 0 FreeSans 200 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 7 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 8 nsew ground bidirectional
rlabel metal1 s 814 406 967 474 1 D
port 1 nsew default input
rlabel metal1 s 814 354 866 406 1 D
port 1 nsew default input
rlabel metal1 s 142 406 407 474 1 SI
port 3 nsew default input
rlabel metal1 s 142 354 194 406 1 SI
port 3 nsew default input
rlabel metal1 s 4141 729 4197 850 1 Q
port 5 nsew default output
rlabel metal1 s 4141 683 4607 729 1 Q
port 5 nsew default output
rlabel metal1 s 4141 430 4187 683 1 Q
port 5 nsew default output
rlabel metal1 s 4141 384 4562 430 1 Q
port 5 nsew default output
rlabel metal1 s 4510 331 4562 384 1 Q
port 5 nsew default output
rlabel metal1 s 4141 331 4187 384 1 Q
port 5 nsew default output
rlabel metal1 s 4510 242 4635 331 1 Q
port 5 nsew default output
rlabel metal1 s 4141 242 4187 331 1 Q
port 5 nsew default output
rlabel metal1 s 4589 169 4635 242 1 Q
port 5 nsew default output
rlabel metal1 s 4141 169 4187 242 1 Q
port 5 nsew default output
rlabel metal1 s 4786 827 4832 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4355 827 4401 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3947 827 3993 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3529 827 3575 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2617 827 2663 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1047 827 1093 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 329 827 375 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4786 781 4832 827 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4355 781 4401 827 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3947 781 3993 827 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3529 781 3575 827 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2617 781 2663 827 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1047 781 1634 827 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 329 781 375 827 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4786 775 4832 781 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4355 775 4401 781 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3947 775 3993 781 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3529 775 3575 781 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2617 775 2663 781 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 329 775 375 781 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3529 710 3575 775 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2617 710 2663 775 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 329 710 375 775 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2617 688 2663 710 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 329 688 375 710 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3917 233 3963 279 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3549 233 3595 279 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4813 215 4859 233 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4365 215 4411 233 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3917 215 3963 233 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3549 215 3595 233 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4813 125 4859 215 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4365 125 4411 215 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3917 125 3963 215 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3549 125 3595 215 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 262 125 330 215 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4813 90 4859 125 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4365 90 4411 125 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3917 90 3963 125 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3549 90 3595 125 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2584 90 2630 125 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1513 90 1559 125 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1101 90 1147 125 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 262 90 330 125 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 4928 90 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4928 1008
string GDS_END 333414
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 322692
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
