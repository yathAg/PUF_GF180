magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< polysilicon >>
rect 22205 59506 22518 59525
rect 22205 59371 22453 59506
rect 22434 59366 22453 59371
rect 22499 59366 22518 59506
rect 22434 59347 22518 59366
rect 22205 57848 22518 57983
rect 22205 57829 22453 57848
rect 22434 57725 22453 57829
rect 22205 57708 22453 57725
rect 22499 57708 22518 57848
rect 22205 57571 22518 57708
rect 22205 56082 22573 56183
rect 22205 56036 22454 56082
rect 22500 56036 22573 56082
rect 22205 56029 22573 56036
rect 22381 55925 22573 56029
rect 22205 55918 22573 55925
rect 22205 55872 22454 55918
rect 22500 55872 22573 55918
rect 22205 55771 22573 55872
rect 22205 54282 22573 54383
rect 22205 54236 22454 54282
rect 22500 54236 22573 54282
rect 22205 54229 22573 54236
rect 22381 54125 22573 54229
rect 22205 54118 22573 54125
rect 22205 54072 22454 54118
rect 22500 54072 22573 54118
rect 22205 53971 22573 54072
rect 22205 52482 22573 52583
rect 22205 52436 22454 52482
rect 22500 52436 22573 52482
rect 22205 52429 22573 52436
rect 22381 52325 22573 52429
rect 22205 52318 22573 52325
rect 22205 52272 22454 52318
rect 22500 52272 22573 52318
rect 22205 52171 22573 52272
rect 22205 50682 22573 50783
rect 22205 50636 22454 50682
rect 22500 50636 22573 50682
rect 22205 50629 22573 50636
rect 22381 50525 22573 50629
rect 22205 50518 22573 50525
rect 22205 50472 22454 50518
rect 22500 50472 22573 50518
rect 22205 50371 22573 50472
rect 22205 48882 22573 48983
rect 22205 48836 22454 48882
rect 22500 48836 22573 48882
rect 22205 48829 22573 48836
rect 22381 48725 22573 48829
rect 22205 48718 22573 48725
rect 22205 48672 22454 48718
rect 22500 48672 22573 48718
rect 22205 48571 22573 48672
rect 22205 47082 22573 47183
rect 22205 47036 22454 47082
rect 22500 47036 22573 47082
rect 22205 47029 22573 47036
rect 22381 46925 22573 47029
rect 22205 46918 22573 46925
rect 22205 46872 22454 46918
rect 22500 46872 22573 46918
rect 22205 46771 22573 46872
rect 22205 45282 22573 45383
rect 22205 45236 22454 45282
rect 22500 45236 22573 45282
rect 22205 45229 22573 45236
rect 22381 45125 22573 45229
rect 22205 45118 22573 45125
rect 22205 45072 22454 45118
rect 22500 45072 22573 45118
rect 22205 44971 22573 45072
rect 22205 43482 22573 43583
rect 22205 43436 22454 43482
rect 22500 43436 22573 43482
rect 22205 43429 22573 43436
rect 22381 43325 22573 43429
rect 22205 43318 22573 43325
rect 22205 43272 22454 43318
rect 22500 43272 22573 43318
rect 22205 43171 22573 43272
rect 22205 41682 22573 41783
rect 22205 41636 22454 41682
rect 22500 41636 22573 41682
rect 22205 41629 22573 41636
rect 22381 41525 22573 41629
rect 22205 41518 22573 41525
rect 22205 41472 22454 41518
rect 22500 41472 22573 41518
rect 22205 41371 22573 41472
rect 22205 39882 22573 39983
rect 22205 39836 22454 39882
rect 22500 39836 22573 39882
rect 22205 39829 22573 39836
rect 22381 39725 22573 39829
rect 22205 39718 22573 39725
rect 22205 39672 22454 39718
rect 22500 39672 22573 39718
rect 22205 39571 22573 39672
rect 22205 38082 22573 38183
rect 22205 38036 22454 38082
rect 22500 38036 22573 38082
rect 22205 38029 22573 38036
rect 22381 37925 22573 38029
rect 22205 37918 22573 37925
rect 22205 37872 22454 37918
rect 22500 37872 22573 37918
rect 22205 37771 22573 37872
rect 22205 36282 22573 36383
rect 22205 36236 22454 36282
rect 22500 36236 22573 36282
rect 22205 36229 22573 36236
rect 22381 36125 22573 36229
rect 22205 36118 22573 36125
rect 22205 36072 22454 36118
rect 22500 36072 22573 36118
rect 22205 35971 22573 36072
rect 22205 34482 22573 34583
rect 22205 34436 22454 34482
rect 22500 34436 22573 34482
rect 22205 34429 22573 34436
rect 22381 34325 22573 34429
rect 22205 34318 22573 34325
rect 22205 34272 22454 34318
rect 22500 34272 22573 34318
rect 22205 34171 22573 34272
rect 22205 32682 22573 32783
rect 22205 32636 22454 32682
rect 22500 32636 22573 32682
rect 22205 32629 22573 32636
rect 22381 32525 22573 32629
rect 22205 32518 22573 32525
rect 22205 32472 22454 32518
rect 22500 32472 22573 32518
rect 22205 32371 22573 32472
rect 22205 30882 22573 30983
rect 22205 30836 22454 30882
rect 22500 30836 22573 30882
rect 22205 30829 22573 30836
rect 22381 30725 22573 30829
rect 22205 30718 22573 30725
rect 22205 30672 22454 30718
rect 22500 30672 22573 30718
rect 22205 30571 22573 30672
rect 22205 29082 22573 29183
rect 22205 29036 22454 29082
rect 22500 29036 22573 29082
rect 22205 29029 22573 29036
rect 22381 28925 22573 29029
rect 22205 28918 22573 28925
rect 22205 28872 22454 28918
rect 22500 28872 22573 28918
rect 22205 28771 22573 28872
rect 22205 27282 22573 27383
rect 22205 27236 22454 27282
rect 22500 27236 22573 27282
rect 22205 27229 22573 27236
rect 22381 27125 22573 27229
rect 22205 27118 22573 27125
rect 22205 27072 22454 27118
rect 22500 27072 22573 27118
rect 22205 26971 22573 27072
rect 22205 25482 22573 25583
rect 22205 25436 22454 25482
rect 22500 25436 22573 25482
rect 22205 25429 22573 25436
rect 22381 25325 22573 25429
rect 22205 25318 22573 25325
rect 22205 25272 22454 25318
rect 22500 25272 22573 25318
rect 22205 25171 22573 25272
rect 22205 23682 22573 23783
rect 22205 23636 22454 23682
rect 22500 23636 22573 23682
rect 22205 23629 22573 23636
rect 22381 23525 22573 23629
rect 22205 23518 22573 23525
rect 22205 23472 22454 23518
rect 22500 23472 22573 23518
rect 22205 23371 22573 23472
rect 22205 21882 22573 21983
rect 22205 21836 22454 21882
rect 22500 21836 22573 21882
rect 22205 21829 22573 21836
rect 22381 21725 22573 21829
rect 22205 21718 22573 21725
rect 22205 21672 22454 21718
rect 22500 21672 22573 21718
rect 22205 21571 22573 21672
rect 22205 20082 22573 20183
rect 22205 20036 22454 20082
rect 22500 20036 22573 20082
rect 22205 20029 22573 20036
rect 22381 19925 22573 20029
rect 22205 19918 22573 19925
rect 22205 19872 22454 19918
rect 22500 19872 22573 19918
rect 22205 19771 22573 19872
rect 22205 18282 22573 18383
rect 22205 18236 22454 18282
rect 22500 18236 22573 18282
rect 22205 18229 22573 18236
rect 22381 18125 22573 18229
rect 22205 18118 22573 18125
rect 22205 18072 22454 18118
rect 22500 18072 22573 18118
rect 22205 17971 22573 18072
rect 22205 16482 22573 16583
rect 22205 16436 22454 16482
rect 22500 16436 22573 16482
rect 22205 16429 22573 16436
rect 22381 16325 22573 16429
rect 22205 16318 22573 16325
rect 22205 16272 22454 16318
rect 22500 16272 22573 16318
rect 22205 16171 22573 16272
rect 22205 14682 22573 14783
rect 22205 14636 22454 14682
rect 22500 14636 22573 14682
rect 22205 14629 22573 14636
rect 22381 14525 22573 14629
rect 22205 14518 22573 14525
rect 22205 14472 22454 14518
rect 22500 14472 22573 14518
rect 22205 14371 22573 14472
rect 22205 12882 22573 12983
rect 22205 12836 22454 12882
rect 22500 12836 22573 12882
rect 22205 12829 22573 12836
rect 22381 12725 22573 12829
rect 22205 12718 22573 12725
rect 22205 12672 22454 12718
rect 22500 12672 22573 12718
rect 22205 12571 22573 12672
rect 22205 11082 22573 11183
rect 22205 11036 22454 11082
rect 22500 11036 22573 11082
rect 22205 11029 22573 11036
rect 22381 10925 22573 11029
rect 22205 10918 22573 10925
rect 22205 10872 22454 10918
rect 22500 10872 22573 10918
rect 22205 10771 22573 10872
rect 22205 9282 22573 9383
rect 22205 9236 22454 9282
rect 22500 9236 22573 9282
rect 22205 9229 22573 9236
rect 22381 9125 22573 9229
rect 22205 9118 22573 9125
rect 22205 9072 22454 9118
rect 22500 9072 22573 9118
rect 22205 8971 22573 9072
rect 22205 7482 22573 7583
rect 22205 7436 22454 7482
rect 22500 7436 22573 7482
rect 22205 7429 22573 7436
rect 22381 7325 22573 7429
rect 22205 7318 22573 7325
rect 22205 7272 22454 7318
rect 22500 7272 22573 7318
rect 22205 7171 22573 7272
rect 22205 5682 22573 5783
rect 22205 5636 22454 5682
rect 22500 5636 22573 5682
rect 22205 5629 22573 5636
rect 22381 5525 22573 5629
rect 22205 5518 22573 5525
rect 22205 5472 22454 5518
rect 22500 5472 22573 5518
rect 22205 5371 22573 5472
rect 22205 3882 22573 3983
rect 22205 3836 22454 3882
rect 22500 3836 22573 3882
rect 22205 3829 22573 3836
rect 22381 3725 22573 3829
rect 22205 3718 22573 3725
rect 22205 3672 22454 3718
rect 22500 3672 22573 3718
rect 22205 3571 22573 3672
rect 22205 2082 22573 2183
rect 22205 2036 22454 2082
rect 22500 2036 22573 2082
rect 22205 2029 22573 2036
rect 22381 1925 22573 2029
rect 22205 1918 22573 1925
rect 22205 1872 22454 1918
rect 22500 1872 22573 1918
rect 22205 1771 22573 1872
rect 22381 522 22573 568
rect 22381 476 22454 522
rect 22500 476 22573 522
rect 22381 383 22573 476
rect 22205 358 22573 383
rect 22205 312 22454 358
rect 22500 312 22573 358
rect 22205 229 22573 312
<< polycontact >>
rect 22453 59366 22499 59506
rect 22453 57708 22499 57848
rect 22454 56036 22500 56082
rect 22454 55872 22500 55918
rect 22454 54236 22500 54282
rect 22454 54072 22500 54118
rect 22454 52436 22500 52482
rect 22454 52272 22500 52318
rect 22454 50636 22500 50682
rect 22454 50472 22500 50518
rect 22454 48836 22500 48882
rect 22454 48672 22500 48718
rect 22454 47036 22500 47082
rect 22454 46872 22500 46918
rect 22454 45236 22500 45282
rect 22454 45072 22500 45118
rect 22454 43436 22500 43482
rect 22454 43272 22500 43318
rect 22454 41636 22500 41682
rect 22454 41472 22500 41518
rect 22454 39836 22500 39882
rect 22454 39672 22500 39718
rect 22454 38036 22500 38082
rect 22454 37872 22500 37918
rect 22454 36236 22500 36282
rect 22454 36072 22500 36118
rect 22454 34436 22500 34482
rect 22454 34272 22500 34318
rect 22454 32636 22500 32682
rect 22454 32472 22500 32518
rect 22454 30836 22500 30882
rect 22454 30672 22500 30718
rect 22454 29036 22500 29082
rect 22454 28872 22500 28918
rect 22454 27236 22500 27282
rect 22454 27072 22500 27118
rect 22454 25436 22500 25482
rect 22454 25272 22500 25318
rect 22454 23636 22500 23682
rect 22454 23472 22500 23518
rect 22454 21836 22500 21882
rect 22454 21672 22500 21718
rect 22454 20036 22500 20082
rect 22454 19872 22500 19918
rect 22454 18236 22500 18282
rect 22454 18072 22500 18118
rect 22454 16436 22500 16482
rect 22454 16272 22500 16318
rect 22454 14636 22500 14682
rect 22454 14472 22500 14518
rect 22454 12836 22500 12882
rect 22454 12672 22500 12718
rect 22454 11036 22500 11082
rect 22454 10872 22500 10918
rect 22454 9236 22500 9282
rect 22454 9072 22500 9118
rect 22454 7436 22500 7482
rect 22454 7272 22500 7318
rect 22454 5636 22500 5682
rect 22454 5472 22500 5518
rect 22454 3836 22500 3882
rect 22454 3672 22500 3718
rect 22454 2036 22500 2082
rect 22454 1872 22500 1918
rect 22454 476 22500 522
rect 22454 312 22500 358
<< metal1 >>
rect 22438 59506 22514 59517
rect 22438 59505 22453 59506
rect 22499 59505 22514 59506
rect 22438 59245 22450 59505
rect 22502 59245 22514 59505
rect 22438 59233 22514 59245
rect 22413 57910 22537 57950
rect 22413 57858 22449 57910
rect 22501 57858 22537 57910
rect 22413 57848 22537 57858
rect 22413 57708 22453 57848
rect 22499 57708 22537 57848
rect 22413 57692 22537 57708
rect 22413 57640 22449 57692
rect 22501 57640 22537 57692
rect 22413 57600 22537 57640
rect 22413 56110 22537 56150
rect 22413 56058 22449 56110
rect 22501 56058 22537 56110
rect 22413 56036 22454 56058
rect 22500 56036 22537 56058
rect 22413 55918 22537 56036
rect 22413 55892 22454 55918
rect 22500 55892 22537 55918
rect 22413 55840 22449 55892
rect 22501 55840 22537 55892
rect 22413 55800 22537 55840
rect 22413 54310 22537 54350
rect 22413 54258 22449 54310
rect 22501 54258 22537 54310
rect 22413 54236 22454 54258
rect 22500 54236 22537 54258
rect 22413 54118 22537 54236
rect 22413 54092 22454 54118
rect 22500 54092 22537 54118
rect 22413 54040 22449 54092
rect 22501 54040 22537 54092
rect 22413 54000 22537 54040
rect 22413 52510 22537 52550
rect 22413 52458 22449 52510
rect 22501 52458 22537 52510
rect 22413 52436 22454 52458
rect 22500 52436 22537 52458
rect 22413 52318 22537 52436
rect 22413 52292 22454 52318
rect 22500 52292 22537 52318
rect 22413 52240 22449 52292
rect 22501 52240 22537 52292
rect 22413 52200 22537 52240
rect 22413 50710 22537 50750
rect 22413 50658 22449 50710
rect 22501 50658 22537 50710
rect 22413 50636 22454 50658
rect 22500 50636 22537 50658
rect 22413 50518 22537 50636
rect 22413 50492 22454 50518
rect 22500 50492 22537 50518
rect 22413 50440 22449 50492
rect 22501 50440 22537 50492
rect 22413 50400 22537 50440
rect 22413 48910 22537 48950
rect 22413 48858 22449 48910
rect 22501 48858 22537 48910
rect 22413 48836 22454 48858
rect 22500 48836 22537 48858
rect 22413 48718 22537 48836
rect 22413 48692 22454 48718
rect 22500 48692 22537 48718
rect 22413 48640 22449 48692
rect 22501 48640 22537 48692
rect 22413 48600 22537 48640
rect 22413 47110 22537 47150
rect 22413 47058 22449 47110
rect 22501 47058 22537 47110
rect 22413 47036 22454 47058
rect 22500 47036 22537 47058
rect 22413 46918 22537 47036
rect 22413 46892 22454 46918
rect 22500 46892 22537 46918
rect 22413 46840 22449 46892
rect 22501 46840 22537 46892
rect 22413 46800 22537 46840
rect 22413 45310 22537 45350
rect 22413 45258 22449 45310
rect 22501 45258 22537 45310
rect 22413 45236 22454 45258
rect 22500 45236 22537 45258
rect 22413 45118 22537 45236
rect 22413 45092 22454 45118
rect 22500 45092 22537 45118
rect 22413 45040 22449 45092
rect 22501 45040 22537 45092
rect 22413 45000 22537 45040
rect 22413 43510 22537 43550
rect 22413 43458 22449 43510
rect 22501 43458 22537 43510
rect 22413 43436 22454 43458
rect 22500 43436 22537 43458
rect 22413 43318 22537 43436
rect 22413 43292 22454 43318
rect 22500 43292 22537 43318
rect 22413 43240 22449 43292
rect 22501 43240 22537 43292
rect 22413 43200 22537 43240
rect 22413 41710 22537 41750
rect 22413 41658 22449 41710
rect 22501 41658 22537 41710
rect 22413 41636 22454 41658
rect 22500 41636 22537 41658
rect 22413 41518 22537 41636
rect 22413 41492 22454 41518
rect 22500 41492 22537 41518
rect 22413 41440 22449 41492
rect 22501 41440 22537 41492
rect 22413 41400 22537 41440
rect 22413 39910 22537 39950
rect 22413 39858 22449 39910
rect 22501 39858 22537 39910
rect 22413 39836 22454 39858
rect 22500 39836 22537 39858
rect 22413 39718 22537 39836
rect 22413 39692 22454 39718
rect 22500 39692 22537 39718
rect 22413 39640 22449 39692
rect 22501 39640 22537 39692
rect 22413 39600 22537 39640
rect 22413 38110 22537 38150
rect 22413 38058 22449 38110
rect 22501 38058 22537 38110
rect 22413 38036 22454 38058
rect 22500 38036 22537 38058
rect 22413 37918 22537 38036
rect 22413 37892 22454 37918
rect 22500 37892 22537 37918
rect 22413 37840 22449 37892
rect 22501 37840 22537 37892
rect 22413 37800 22537 37840
rect 22413 36310 22537 36350
rect 22413 36258 22449 36310
rect 22501 36258 22537 36310
rect 22413 36236 22454 36258
rect 22500 36236 22537 36258
rect 22413 36118 22537 36236
rect 22413 36092 22454 36118
rect 22500 36092 22537 36118
rect 22413 36040 22449 36092
rect 22501 36040 22537 36092
rect 22413 36000 22537 36040
rect 22413 34510 22537 34550
rect 22413 34458 22449 34510
rect 22501 34458 22537 34510
rect 22413 34436 22454 34458
rect 22500 34436 22537 34458
rect 22413 34318 22537 34436
rect 22413 34292 22454 34318
rect 22500 34292 22537 34318
rect 22413 34240 22449 34292
rect 22501 34240 22537 34292
rect 22413 34200 22537 34240
rect 22413 32710 22537 32750
rect 22413 32658 22449 32710
rect 22501 32658 22537 32710
rect 22413 32636 22454 32658
rect 22500 32636 22537 32658
rect 22413 32518 22537 32636
rect 22413 32492 22454 32518
rect 22500 32492 22537 32518
rect 22413 32440 22449 32492
rect 22501 32440 22537 32492
rect 22413 32400 22537 32440
rect 22413 30910 22537 30950
rect 22413 30858 22449 30910
rect 22501 30858 22537 30910
rect 22413 30836 22454 30858
rect 22500 30836 22537 30858
rect 22413 30718 22537 30836
rect 22413 30692 22454 30718
rect 22500 30692 22537 30718
rect 22413 30640 22449 30692
rect 22501 30640 22537 30692
rect 22413 30600 22537 30640
rect 22413 29110 22537 29150
rect 22413 29058 22449 29110
rect 22501 29058 22537 29110
rect 22413 29036 22454 29058
rect 22500 29036 22537 29058
rect 22413 28918 22537 29036
rect 22413 28892 22454 28918
rect 22500 28892 22537 28918
rect 22413 28840 22449 28892
rect 22501 28840 22537 28892
rect 22413 28800 22537 28840
rect 22413 27310 22537 27350
rect 22413 27258 22449 27310
rect 22501 27258 22537 27310
rect 22413 27236 22454 27258
rect 22500 27236 22537 27258
rect 22413 27118 22537 27236
rect 22413 27092 22454 27118
rect 22500 27092 22537 27118
rect 22413 27040 22449 27092
rect 22501 27040 22537 27092
rect 22413 27000 22537 27040
rect 22413 25514 22537 25554
rect 22413 25462 22449 25514
rect 22501 25462 22537 25514
rect 22413 25436 22454 25462
rect 22500 25436 22537 25462
rect 22413 25318 22537 25436
rect 22413 25296 22454 25318
rect 22500 25296 22537 25318
rect 22413 25244 22449 25296
rect 22501 25244 22537 25296
rect 22413 25204 22537 25244
rect 22413 23710 22537 23750
rect 22413 23658 22449 23710
rect 22501 23658 22537 23710
rect 22413 23636 22454 23658
rect 22500 23636 22537 23658
rect 22413 23518 22537 23636
rect 22413 23492 22454 23518
rect 22500 23492 22537 23518
rect 22413 23440 22449 23492
rect 22501 23440 22537 23492
rect 22413 23400 22537 23440
rect 22413 21914 22537 21954
rect 22413 21862 22449 21914
rect 22501 21862 22537 21914
rect 22413 21836 22454 21862
rect 22500 21836 22537 21862
rect 22413 21718 22537 21836
rect 22413 21696 22454 21718
rect 22500 21696 22537 21718
rect 22413 21644 22449 21696
rect 22501 21644 22537 21696
rect 22413 21604 22537 21644
rect 22413 20110 22537 20150
rect 22413 20058 22449 20110
rect 22501 20058 22537 20110
rect 22413 20036 22454 20058
rect 22500 20036 22537 20058
rect 22413 19918 22537 20036
rect 22413 19892 22454 19918
rect 22500 19892 22537 19918
rect 22413 19840 22449 19892
rect 22501 19840 22537 19892
rect 22413 19800 22537 19840
rect 22413 18314 22537 18354
rect 22413 18262 22449 18314
rect 22501 18262 22537 18314
rect 22413 18236 22454 18262
rect 22500 18236 22537 18262
rect 22413 18118 22537 18236
rect 22413 18096 22454 18118
rect 22500 18096 22537 18118
rect 22413 18044 22449 18096
rect 22501 18044 22537 18096
rect 22413 18004 22537 18044
rect 22413 16510 22537 16550
rect 22413 16458 22449 16510
rect 22501 16458 22537 16510
rect 22413 16436 22454 16458
rect 22500 16436 22537 16458
rect 22413 16318 22537 16436
rect 22413 16292 22454 16318
rect 22500 16292 22537 16318
rect 22413 16240 22449 16292
rect 22501 16240 22537 16292
rect 22413 16200 22537 16240
rect 22413 14714 22537 14754
rect 22413 14662 22449 14714
rect 22501 14662 22537 14714
rect 22413 14636 22454 14662
rect 22500 14636 22537 14662
rect 22413 14518 22537 14636
rect 22413 14496 22454 14518
rect 22500 14496 22537 14518
rect 22413 14444 22449 14496
rect 22501 14444 22537 14496
rect 22413 14404 22537 14444
rect 22413 12910 22537 12950
rect 22413 12858 22449 12910
rect 22501 12858 22537 12910
rect 22413 12836 22454 12858
rect 22500 12836 22537 12858
rect 22413 12718 22537 12836
rect 22413 12692 22454 12718
rect 22500 12692 22537 12718
rect 22413 12640 22449 12692
rect 22501 12640 22537 12692
rect 22413 12600 22537 12640
rect 22413 11114 22537 11154
rect 22413 11062 22449 11114
rect 22501 11062 22537 11114
rect 22413 11036 22454 11062
rect 22500 11036 22537 11062
rect 22413 10918 22537 11036
rect 22413 10896 22454 10918
rect 22500 10896 22537 10918
rect 22413 10844 22449 10896
rect 22501 10844 22537 10896
rect 22413 10804 22537 10844
rect 22413 9310 22537 9350
rect 22413 9258 22449 9310
rect 22501 9258 22537 9310
rect 22413 9236 22454 9258
rect 22500 9236 22537 9258
rect 22413 9118 22537 9236
rect 22413 9092 22454 9118
rect 22500 9092 22537 9118
rect 22413 9040 22449 9092
rect 22501 9040 22537 9092
rect 22413 9000 22537 9040
rect 22413 7514 22537 7554
rect 22413 7462 22449 7514
rect 22501 7462 22537 7514
rect 22413 7436 22454 7462
rect 22500 7436 22537 7462
rect 22413 7318 22537 7436
rect 22413 7296 22454 7318
rect 22500 7296 22537 7318
rect 22413 7244 22449 7296
rect 22501 7244 22537 7296
rect 22413 7204 22537 7244
rect 22413 5710 22537 5750
rect 22413 5658 22449 5710
rect 22501 5658 22537 5710
rect 22413 5636 22454 5658
rect 22500 5636 22537 5658
rect 22413 5518 22537 5636
rect 22413 5492 22454 5518
rect 22500 5492 22537 5518
rect 22413 5440 22449 5492
rect 22501 5440 22537 5492
rect 22413 5400 22537 5440
rect 22413 3914 22537 3954
rect 22413 3862 22449 3914
rect 22501 3862 22537 3914
rect 22413 3836 22454 3862
rect 22500 3836 22537 3862
rect 22413 3718 22537 3836
rect 22413 3696 22454 3718
rect 22500 3696 22537 3718
rect 22413 3644 22449 3696
rect 22501 3644 22537 3696
rect 22413 3604 22537 3644
rect 22413 2110 22537 2150
rect 22413 2058 22449 2110
rect 22501 2058 22537 2110
rect 22413 2036 22454 2058
rect 22500 2036 22537 2058
rect 22413 1918 22537 2036
rect 22413 1892 22454 1918
rect 22500 1892 22537 1918
rect 22413 1840 22449 1892
rect 22501 1840 22537 1892
rect 22413 1800 22537 1840
rect 22421 522 22533 559
rect 22421 476 22454 522
rect 22500 476 22533 522
rect 22421 455 22533 476
rect 22421 299 22449 455
rect 22501 299 22533 455
rect 22421 276 22533 299
<< via1 >>
rect 22450 59366 22453 59505
rect 22453 59366 22499 59505
rect 22499 59366 22502 59505
rect 22450 59245 22502 59366
rect 22449 57858 22501 57910
rect 22449 57640 22501 57692
rect 22449 56082 22501 56110
rect 22449 56058 22454 56082
rect 22454 56058 22500 56082
rect 22500 56058 22501 56082
rect 22449 55872 22454 55892
rect 22454 55872 22500 55892
rect 22500 55872 22501 55892
rect 22449 55840 22501 55872
rect 22449 54282 22501 54310
rect 22449 54258 22454 54282
rect 22454 54258 22500 54282
rect 22500 54258 22501 54282
rect 22449 54072 22454 54092
rect 22454 54072 22500 54092
rect 22500 54072 22501 54092
rect 22449 54040 22501 54072
rect 22449 52482 22501 52510
rect 22449 52458 22454 52482
rect 22454 52458 22500 52482
rect 22500 52458 22501 52482
rect 22449 52272 22454 52292
rect 22454 52272 22500 52292
rect 22500 52272 22501 52292
rect 22449 52240 22501 52272
rect 22449 50682 22501 50710
rect 22449 50658 22454 50682
rect 22454 50658 22500 50682
rect 22500 50658 22501 50682
rect 22449 50472 22454 50492
rect 22454 50472 22500 50492
rect 22500 50472 22501 50492
rect 22449 50440 22501 50472
rect 22449 48882 22501 48910
rect 22449 48858 22454 48882
rect 22454 48858 22500 48882
rect 22500 48858 22501 48882
rect 22449 48672 22454 48692
rect 22454 48672 22500 48692
rect 22500 48672 22501 48692
rect 22449 48640 22501 48672
rect 22449 47082 22501 47110
rect 22449 47058 22454 47082
rect 22454 47058 22500 47082
rect 22500 47058 22501 47082
rect 22449 46872 22454 46892
rect 22454 46872 22500 46892
rect 22500 46872 22501 46892
rect 22449 46840 22501 46872
rect 22449 45282 22501 45310
rect 22449 45258 22454 45282
rect 22454 45258 22500 45282
rect 22500 45258 22501 45282
rect 22449 45072 22454 45092
rect 22454 45072 22500 45092
rect 22500 45072 22501 45092
rect 22449 45040 22501 45072
rect 22449 43482 22501 43510
rect 22449 43458 22454 43482
rect 22454 43458 22500 43482
rect 22500 43458 22501 43482
rect 22449 43272 22454 43292
rect 22454 43272 22500 43292
rect 22500 43272 22501 43292
rect 22449 43240 22501 43272
rect 22449 41682 22501 41710
rect 22449 41658 22454 41682
rect 22454 41658 22500 41682
rect 22500 41658 22501 41682
rect 22449 41472 22454 41492
rect 22454 41472 22500 41492
rect 22500 41472 22501 41492
rect 22449 41440 22501 41472
rect 22449 39882 22501 39910
rect 22449 39858 22454 39882
rect 22454 39858 22500 39882
rect 22500 39858 22501 39882
rect 22449 39672 22454 39692
rect 22454 39672 22500 39692
rect 22500 39672 22501 39692
rect 22449 39640 22501 39672
rect 22449 38082 22501 38110
rect 22449 38058 22454 38082
rect 22454 38058 22500 38082
rect 22500 38058 22501 38082
rect 22449 37872 22454 37892
rect 22454 37872 22500 37892
rect 22500 37872 22501 37892
rect 22449 37840 22501 37872
rect 22449 36282 22501 36310
rect 22449 36258 22454 36282
rect 22454 36258 22500 36282
rect 22500 36258 22501 36282
rect 22449 36072 22454 36092
rect 22454 36072 22500 36092
rect 22500 36072 22501 36092
rect 22449 36040 22501 36072
rect 22449 34482 22501 34510
rect 22449 34458 22454 34482
rect 22454 34458 22500 34482
rect 22500 34458 22501 34482
rect 22449 34272 22454 34292
rect 22454 34272 22500 34292
rect 22500 34272 22501 34292
rect 22449 34240 22501 34272
rect 22449 32682 22501 32710
rect 22449 32658 22454 32682
rect 22454 32658 22500 32682
rect 22500 32658 22501 32682
rect 22449 32472 22454 32492
rect 22454 32472 22500 32492
rect 22500 32472 22501 32492
rect 22449 32440 22501 32472
rect 22449 30882 22501 30910
rect 22449 30858 22454 30882
rect 22454 30858 22500 30882
rect 22500 30858 22501 30882
rect 22449 30672 22454 30692
rect 22454 30672 22500 30692
rect 22500 30672 22501 30692
rect 22449 30640 22501 30672
rect 22449 29082 22501 29110
rect 22449 29058 22454 29082
rect 22454 29058 22500 29082
rect 22500 29058 22501 29082
rect 22449 28872 22454 28892
rect 22454 28872 22500 28892
rect 22500 28872 22501 28892
rect 22449 28840 22501 28872
rect 22449 27282 22501 27310
rect 22449 27258 22454 27282
rect 22454 27258 22500 27282
rect 22500 27258 22501 27282
rect 22449 27072 22454 27092
rect 22454 27072 22500 27092
rect 22500 27072 22501 27092
rect 22449 27040 22501 27072
rect 22449 25482 22501 25514
rect 22449 25462 22454 25482
rect 22454 25462 22500 25482
rect 22500 25462 22501 25482
rect 22449 25272 22454 25296
rect 22454 25272 22500 25296
rect 22500 25272 22501 25296
rect 22449 25244 22501 25272
rect 22449 23682 22501 23710
rect 22449 23658 22454 23682
rect 22454 23658 22500 23682
rect 22500 23658 22501 23682
rect 22449 23472 22454 23492
rect 22454 23472 22500 23492
rect 22500 23472 22501 23492
rect 22449 23440 22501 23472
rect 22449 21882 22501 21914
rect 22449 21862 22454 21882
rect 22454 21862 22500 21882
rect 22500 21862 22501 21882
rect 22449 21672 22454 21696
rect 22454 21672 22500 21696
rect 22500 21672 22501 21696
rect 22449 21644 22501 21672
rect 22449 20082 22501 20110
rect 22449 20058 22454 20082
rect 22454 20058 22500 20082
rect 22500 20058 22501 20082
rect 22449 19872 22454 19892
rect 22454 19872 22500 19892
rect 22500 19872 22501 19892
rect 22449 19840 22501 19872
rect 22449 18282 22501 18314
rect 22449 18262 22454 18282
rect 22454 18262 22500 18282
rect 22500 18262 22501 18282
rect 22449 18072 22454 18096
rect 22454 18072 22500 18096
rect 22500 18072 22501 18096
rect 22449 18044 22501 18072
rect 22449 16482 22501 16510
rect 22449 16458 22454 16482
rect 22454 16458 22500 16482
rect 22500 16458 22501 16482
rect 22449 16272 22454 16292
rect 22454 16272 22500 16292
rect 22500 16272 22501 16292
rect 22449 16240 22501 16272
rect 22449 14682 22501 14714
rect 22449 14662 22454 14682
rect 22454 14662 22500 14682
rect 22500 14662 22501 14682
rect 22449 14472 22454 14496
rect 22454 14472 22500 14496
rect 22500 14472 22501 14496
rect 22449 14444 22501 14472
rect 22449 12882 22501 12910
rect 22449 12858 22454 12882
rect 22454 12858 22500 12882
rect 22500 12858 22501 12882
rect 22449 12672 22454 12692
rect 22454 12672 22500 12692
rect 22500 12672 22501 12692
rect 22449 12640 22501 12672
rect 22449 11082 22501 11114
rect 22449 11062 22454 11082
rect 22454 11062 22500 11082
rect 22500 11062 22501 11082
rect 22449 10872 22454 10896
rect 22454 10872 22500 10896
rect 22500 10872 22501 10896
rect 22449 10844 22501 10872
rect 22449 9282 22501 9310
rect 22449 9258 22454 9282
rect 22454 9258 22500 9282
rect 22500 9258 22501 9282
rect 22449 9072 22454 9092
rect 22454 9072 22500 9092
rect 22500 9072 22501 9092
rect 22449 9040 22501 9072
rect 22449 7482 22501 7514
rect 22449 7462 22454 7482
rect 22454 7462 22500 7482
rect 22500 7462 22501 7482
rect 22449 7272 22454 7296
rect 22454 7272 22500 7296
rect 22500 7272 22501 7296
rect 22449 7244 22501 7272
rect 22449 5682 22501 5710
rect 22449 5658 22454 5682
rect 22454 5658 22500 5682
rect 22500 5658 22501 5682
rect 22449 5472 22454 5492
rect 22454 5472 22500 5492
rect 22500 5472 22501 5492
rect 22449 5440 22501 5472
rect 22449 3882 22501 3914
rect 22449 3862 22454 3882
rect 22454 3862 22500 3882
rect 22500 3862 22501 3882
rect 22449 3672 22454 3696
rect 22454 3672 22500 3696
rect 22500 3672 22501 3696
rect 22449 3644 22501 3672
rect 22449 2082 22501 2110
rect 22449 2058 22454 2082
rect 22454 2058 22500 2082
rect 22500 2058 22501 2082
rect 22449 1872 22454 1892
rect 22454 1872 22500 1892
rect 22500 1872 22501 1892
rect 22449 1840 22501 1872
rect 22449 358 22501 455
rect 22449 312 22454 358
rect 22454 312 22500 358
rect 22500 312 22501 358
rect 22449 299 22501 312
<< metal2 >>
rect 22412 59657 22537 59677
rect 22412 59497 22448 59657
rect 22504 59497 22537 59657
rect 22412 59245 22450 59497
rect 22502 59245 22537 59497
rect 22412 57910 22537 59245
rect 22412 57858 22449 57910
rect 22501 57858 22537 57910
rect 22412 57692 22537 57858
rect 22412 57640 22449 57692
rect 22501 57640 22537 57692
rect 22412 56110 22537 57640
rect 22412 56058 22449 56110
rect 22501 56058 22537 56110
rect 22412 55892 22537 56058
rect 22412 55840 22449 55892
rect 22501 55840 22537 55892
rect 22412 54310 22537 55840
rect 22412 54258 22449 54310
rect 22501 54258 22537 54310
rect 22412 54092 22537 54258
rect 22412 54040 22449 54092
rect 22501 54040 22537 54092
rect 22412 52510 22537 54040
rect 22412 52458 22449 52510
rect 22501 52458 22537 52510
rect 22412 52292 22537 52458
rect 22412 52240 22449 52292
rect 22501 52240 22537 52292
rect 22412 50710 22537 52240
rect 22412 50658 22449 50710
rect 22501 50658 22537 50710
rect 22412 50492 22537 50658
rect 22412 50440 22449 50492
rect 22501 50440 22537 50492
rect 22412 48910 22537 50440
rect 22412 48858 22449 48910
rect 22501 48858 22537 48910
rect 22412 48692 22537 48858
rect 22412 48640 22449 48692
rect 22501 48640 22537 48692
rect 22412 47110 22537 48640
rect 22412 47058 22449 47110
rect 22501 47058 22537 47110
rect 22412 46892 22537 47058
rect 22412 46840 22449 46892
rect 22501 46840 22537 46892
rect 22412 45310 22537 46840
rect 22412 45258 22449 45310
rect 22501 45258 22537 45310
rect 22412 45092 22537 45258
rect 22412 45040 22449 45092
rect 22501 45040 22537 45092
rect 22412 43510 22537 45040
rect 22412 43458 22449 43510
rect 22501 43458 22537 43510
rect 22412 43292 22537 43458
rect 22412 43240 22449 43292
rect 22501 43240 22537 43292
rect 22412 41710 22537 43240
rect 22412 41658 22449 41710
rect 22501 41658 22537 41710
rect 22412 41492 22537 41658
rect 22412 41440 22449 41492
rect 22501 41440 22537 41492
rect 22412 39910 22537 41440
rect 22412 39858 22449 39910
rect 22501 39858 22537 39910
rect 22412 39692 22537 39858
rect 22412 39640 22449 39692
rect 22501 39640 22537 39692
rect 22412 38110 22537 39640
rect 22412 38058 22449 38110
rect 22501 38058 22537 38110
rect 22412 37892 22537 38058
rect 22412 37840 22449 37892
rect 22501 37840 22537 37892
rect 22412 36310 22537 37840
rect 22412 36258 22449 36310
rect 22501 36258 22537 36310
rect 22412 36092 22537 36258
rect 22412 36040 22449 36092
rect 22501 36040 22537 36092
rect 22412 34510 22537 36040
rect 22412 34458 22449 34510
rect 22501 34458 22537 34510
rect 22412 34292 22537 34458
rect 22412 34240 22449 34292
rect 22501 34240 22537 34292
rect 22412 32710 22537 34240
rect 22412 32658 22449 32710
rect 22501 32658 22537 32710
rect 22412 32492 22537 32658
rect 22412 32440 22449 32492
rect 22501 32440 22537 32492
rect 22412 30910 22537 32440
rect 22412 30858 22449 30910
rect 22501 30858 22537 30910
rect 22412 30692 22537 30858
rect 22412 30640 22449 30692
rect 22501 30640 22537 30692
rect 22412 29110 22537 30640
rect 22412 29058 22449 29110
rect 22501 29058 22537 29110
rect 22412 28892 22537 29058
rect 22412 28840 22449 28892
rect 22501 28840 22537 28892
rect 22412 27310 22537 28840
rect 22412 27258 22449 27310
rect 22501 27258 22537 27310
rect 22412 27092 22537 27258
rect 22412 27040 22449 27092
rect 22501 27040 22537 27092
rect 22412 25514 22537 27040
rect 22412 25462 22449 25514
rect 22501 25462 22537 25514
rect 22412 25296 22537 25462
rect 22412 25244 22449 25296
rect 22501 25244 22537 25296
rect 22412 23710 22537 25244
rect 22412 23658 22449 23710
rect 22501 23658 22537 23710
rect 22412 23492 22537 23658
rect 22412 23440 22449 23492
rect 22501 23440 22537 23492
rect 22412 21914 22537 23440
rect 22412 21862 22449 21914
rect 22501 21862 22537 21914
rect 22412 21696 22537 21862
rect 22412 21644 22449 21696
rect 22501 21644 22537 21696
rect 22412 20110 22537 21644
rect 22412 20058 22449 20110
rect 22501 20058 22537 20110
rect 22412 19892 22537 20058
rect 22412 19840 22449 19892
rect 22501 19840 22537 19892
rect 22412 18314 22537 19840
rect 22412 18262 22449 18314
rect 22501 18262 22537 18314
rect 22412 18096 22537 18262
rect 22412 18044 22449 18096
rect 22501 18044 22537 18096
rect 22412 16510 22537 18044
rect 22412 16458 22449 16510
rect 22501 16458 22537 16510
rect 22412 16292 22537 16458
rect 22412 16240 22449 16292
rect 22501 16240 22537 16292
rect 22412 14714 22537 16240
rect 22412 14662 22449 14714
rect 22501 14662 22537 14714
rect 22412 14496 22537 14662
rect 22412 14444 22449 14496
rect 22501 14444 22537 14496
rect 22412 12910 22537 14444
rect 22412 12858 22449 12910
rect 22501 12858 22537 12910
rect 22412 12692 22537 12858
rect 22412 12640 22449 12692
rect 22501 12640 22537 12692
rect 22412 11114 22537 12640
rect 22412 11062 22449 11114
rect 22501 11062 22537 11114
rect 22412 10896 22537 11062
rect 22412 10844 22449 10896
rect 22501 10844 22537 10896
rect 22412 9310 22537 10844
rect 22412 9258 22449 9310
rect 22501 9258 22537 9310
rect 22412 9092 22537 9258
rect 22412 9040 22449 9092
rect 22501 9040 22537 9092
rect 22412 7514 22537 9040
rect 22412 7462 22449 7514
rect 22501 7462 22537 7514
rect 22412 7296 22537 7462
rect 22412 7244 22449 7296
rect 22501 7244 22537 7296
rect 22412 5710 22537 7244
rect 22412 5658 22449 5710
rect 22501 5658 22537 5710
rect 22412 5492 22537 5658
rect 22412 5440 22449 5492
rect 22501 5440 22537 5492
rect 22412 3914 22537 5440
rect 22412 3862 22449 3914
rect 22501 3862 22537 3914
rect 22412 3696 22537 3862
rect 22412 3644 22449 3696
rect 22501 3644 22537 3696
rect 22412 2110 22537 3644
rect 22412 2058 22449 2110
rect 22501 2058 22537 2110
rect 22412 1892 22537 2058
rect 22412 1840 22449 1892
rect 22501 1840 22537 1892
rect 22412 455 22537 1840
rect 22412 299 22449 455
rect 22501 299 22537 455
rect 22412 256 22537 299
rect 22412 96 22447 256
rect 22503 96 22537 256
rect 22412 76 22537 96
<< via2 >>
rect 22448 59505 22504 59657
rect 22448 59497 22450 59505
rect 22450 59497 22502 59505
rect 22502 59497 22504 59505
rect 22447 96 22503 256
<< metal3 >>
rect -636 59657 22538 59677
rect -636 59497 22448 59657
rect 22504 59497 22538 59657
rect -636 59477 22538 59497
rect -636 256 22537 277
rect -636 96 22447 256
rect 22503 96 22537 256
rect -636 77 22537 96
use 018SRAM_cell1_512x8m81  018SRAM_cell1_512x8m81_0
timestamp 1698431365
transform -1 0 22262 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_512x8m81  018SRAM_cell1_512x8m81_1
timestamp 1698431365
transform -1 0 22262 0 -1 59577
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_0
timestamp 1698431365
transform -1 0 13862 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_1
timestamp 1698431365
transform -1 0 12662 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_2
timestamp 1698431365
transform -1 0 13262 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_3
timestamp 1698431365
transform -1 0 12062 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_4
timestamp 1698431365
transform -1 0 16862 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_5
timestamp 1698431365
transform -1 0 17462 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_6
timestamp 1698431365
transform -1 0 18662 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_7
timestamp 1698431365
transform -1 0 18062 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_8
timestamp 1698431365
transform -1 0 19262 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_9
timestamp 1698431365
transform -1 0 19862 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_10
timestamp 1698431365
transform -1 0 20462 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_11
timestamp 1698431365
transform -1 0 21062 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_12
timestamp 1698431365
transform -1 0 15662 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_13
timestamp 1698431365
transform -1 0 15062 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_14
timestamp 1698431365
transform -1 0 14462 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_15
timestamp 1698431365
transform -1 0 662 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_16
timestamp 1698431365
transform -1 0 6062 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_17
timestamp 1698431365
transform -1 0 6662 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_18
timestamp 1698431365
transform -1 0 7862 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_19
timestamp 1698431365
transform -1 0 7262 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_20
timestamp 1698431365
transform -1 0 8462 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_21
timestamp 1698431365
transform -1 0 9062 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_22
timestamp 1698431365
transform -1 0 9662 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_23
timestamp 1698431365
transform -1 0 10262 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_24
timestamp 1698431365
transform -1 0 4862 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_25
timestamp 1698431365
transform -1 0 4262 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_26
timestamp 1698431365
transform -1 0 3662 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_27
timestamp 1698431365
transform -1 0 3062 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_28
timestamp 1698431365
transform -1 0 1862 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_29
timestamp 1698431365
transform -1 0 2462 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_30
timestamp 1698431365
transform -1 0 1262 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_31
timestamp 1698431365
transform -1 0 11462 0 1 177
box -68 -68 668 968
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_0
timestamp 1698431365
transform -1 0 16262 0 1 177
box -68 -68 668 968
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_1
timestamp 1698431365
transform 1 0 21062 0 1 177
box -68 -68 668 968
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_2
timestamp 1698431365
transform -1 0 10862 0 1 177
box -68 -68 668 968
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_3
timestamp 1698431365
transform -1 0 5462 0 1 177
box -68 -68 668 968
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_4
timestamp 1698431365
transform -1 0 62 0 1 177
box -68 -68 668 968
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_5
timestamp 1698431365
transform -1 0 62 0 -1 59577
box -68 -68 668 968
use array16_512_dummy_01_512x8m81  array16_512_dummy_01_512x8m81_0
timestamp 1698431365
transform 1 0 21594 0 1 1009
box 0 0 736 57736
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_0
timestamp 1698431365
transform 1 0 22477 0 -1 25377
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_1
timestamp 1698431365
transform 1 0 22477 0 -1 21777
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_2
timestamp 1698431365
transform 1 0 22477 0 -1 16377
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_3
timestamp 1698431365
transform 1 0 22477 0 -1 12777
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_4
timestamp 1698431365
transform 1 0 22477 0 -1 9177
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_5
timestamp 1698431365
transform 1 0 22477 0 -1 18177
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_6
timestamp 1698431365
transform 1 0 22477 0 -1 14577
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_7
timestamp 1698431365
transform 1 0 22477 0 -1 10977
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_8
timestamp 1698431365
transform 1 0 22477 0 -1 7377
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_9
timestamp 1698431365
transform 1 0 22477 0 -1 5577
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_10
timestamp 1698431365
transform 1 0 22477 0 -1 1977
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_11
timestamp 1698431365
transform 1 0 22477 0 -1 27177
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_12
timestamp 1698431365
transform 1 0 22477 0 -1 23577
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_13
timestamp 1698431365
transform 1 0 22477 0 -1 19977
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_14
timestamp 1698431365
transform 1 0 22477 0 -1 3777
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_15
timestamp 1698431365
transform 1 0 22477 0 -1 417
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_16
timestamp 1698431365
transform 1 0 22477 0 -1 28977
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_17
timestamp 1698431365
transform 1 0 22477 0 -1 32577
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_18
timestamp 1698431365
transform 1 0 22477 0 -1 34377
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_19
timestamp 1698431365
transform 1 0 22477 0 -1 36177
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_20
timestamp 1698431365
transform 1 0 22477 0 -1 37977
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_21
timestamp 1698431365
transform 1 0 22477 0 -1 39777
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_22
timestamp 1698431365
transform 1 0 22477 0 -1 41577
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_23
timestamp 1698431365
transform 1 0 22477 0 -1 43377
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_24
timestamp 1698431365
transform 1 0 22477 0 -1 45177
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_25
timestamp 1698431365
transform 1 0 22477 0 -1 46977
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_26
timestamp 1698431365
transform 1 0 22477 0 -1 48777
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_27
timestamp 1698431365
transform 1 0 22477 0 -1 50577
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_28
timestamp 1698431365
transform 1 0 22477 0 -1 52377
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_29
timestamp 1698431365
transform 1 0 22477 0 -1 54177
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_30
timestamp 1698431365
transform 1 0 22477 0 -1 55977
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_31
timestamp 1698431365
transform 1 0 22477 0 -1 30777
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_0
timestamp 1698431365
transform 1 0 22476 0 1 59436
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_1
timestamp 1698431365
transform 1 0 22476 0 1 57778
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_0
timestamp 1698431365
transform 1 0 22475 0 -1 7379
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_1
timestamp 1698431365
transform 1 0 22475 0 -1 21779
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_2
timestamp 1698431365
transform 1 0 22475 0 -1 28975
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_3
timestamp 1698431365
transform 1 0 22475 0 -1 14579
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_4
timestamp 1698431365
transform 1 0 22475 0 -1 3779
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_5
timestamp 1698431365
transform 1 0 22475 0 -1 18179
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_6
timestamp 1698431365
transform 1 0 22475 0 -1 25379
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_7
timestamp 1698431365
transform 1 0 22475 0 -1 10979
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_8
timestamp 1698431365
transform 1 0 22475 0 -1 1975
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_9
timestamp 1698431365
transform 1 0 22475 0 -1 5575
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_10
timestamp 1698431365
transform 1 0 22475 0 -1 9175
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_11
timestamp 1698431365
transform 1 0 22475 0 -1 12775
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_12
timestamp 1698431365
transform 1 0 22475 0 -1 16375
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_13
timestamp 1698431365
transform 1 0 22475 0 -1 19975
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_14
timestamp 1698431365
transform 1 0 22475 0 -1 23575
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_15
timestamp 1698431365
transform 1 0 22475 0 -1 27175
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_16
timestamp 1698431365
transform 1 0 22475 0 -1 32575
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_17
timestamp 1698431365
transform 1 0 22475 0 -1 34375
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_18
timestamp 1698431365
transform 1 0 22475 0 -1 36175
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_19
timestamp 1698431365
transform 1 0 22475 0 -1 37975
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_20
timestamp 1698431365
transform 1 0 22475 0 -1 39775
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_21
timestamp 1698431365
transform 1 0 22475 0 -1 41575
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_22
timestamp 1698431365
transform 1 0 22475 0 -1 43375
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_23
timestamp 1698431365
transform 1 0 22475 0 -1 45175
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_24
timestamp 1698431365
transform 1 0 22475 0 -1 46975
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_25
timestamp 1698431365
transform 1 0 22475 0 -1 48775
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_26
timestamp 1698431365
transform 1 0 22475 0 -1 50575
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_27
timestamp 1698431365
transform 1 0 22475 0 -1 52375
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_28
timestamp 1698431365
transform 1 0 22475 0 -1 54175
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_29
timestamp 1698431365
transform 1 0 22475 0 -1 55975
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_30
timestamp 1698431365
transform 1 0 22475 0 -1 57775
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_31
timestamp 1698431365
transform 1 0 22475 0 -1 30775
box 0 0 1 1
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_0
timestamp 1698431365
transform 1 0 22475 0 1 377
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_0
timestamp 1698431365
transform 1 0 22476 0 1 59375
box 0 0 1 1
use M3_M2431059130201_512x8m81  M3_M2431059130201_512x8m81_0
timestamp 1698431365
transform 1 0 22475 0 1 176
box 0 0 1 1
use M3_M2431059130201_512x8m81  M3_M2431059130201_512x8m81_1
timestamp 1698431365
transform 1 0 22476 0 1 59577
box 0 0 1 1
use new_dummyrow_unit_512x8m81  new_dummyrow_unit_512x8m81_0
timestamp 1698431365
transform 1 0 10800 0 -1 59754
box -6 109 10930 1145
use new_dummyrowunit01_512x8m81  new_dummyrowunit01_512x8m81_0
timestamp 1698431365
transform 1 0 0 0 -1 59754
box -6 109 10930 1145
<< properties >>
string GDS_END 2475994
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 2464766
<< end >>
