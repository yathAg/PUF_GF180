magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
use M1_NWELL$$46890028_128x8m81  M1_NWELL$$46890028_128x8m81_0
timestamp 1698431365
transform 1 0 8760 0 1 900
box 0 0 1 1
use M1_NWELL4310590548733_128x8m81  M1_NWELL4310590548733_128x8m81_0
timestamp 1698431365
transform 1 0 6202 0 1 900
box 0 0 1 1
use M1_PACTIVE$$204209196_128x8m81  M1_PACTIVE$$204209196_128x8m81_0
timestamp 1698431365
transform 1 0 4535 0 1 0
box 0 0 1 1
use M1_PACTIVE43105905487105_12_0  M1_PACTIVE43105905487105_12_0_0
timestamp 1698431365
transform 1 0 7811 0 1 900
box 0 0 1 1
use M1_POLY24310590548732_128x8m81  M1_POLY24310590548732_128x8m81_0
timestamp 1698431365
transform 1 0 9900 0 1 687
box 0 0 1 1
use M1_POLY24310590548732_128x8m81  M1_POLY24310590548732_128x8m81_1
timestamp 1698431365
transform 1 0 9463 0 1 256
box 0 0 1 1
use M1_POLY24310590548734_128x8m81  M1_POLY24310590548734_128x8m81_0
timestamp 1698431365
transform 1 0 14024 0 1 564
box 0 0 1 1
use M1_POLY24310590548734_128x8m81  M1_POLY24310590548734_128x8m81_1
timestamp 1698431365
transform 1 0 13039 0 1 759
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_0
timestamp 1698431365
transform 0 1 15130 -1 0 333
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_1
timestamp 1698431365
transform 1 0 6316 0 1 368
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_2
timestamp 1698431365
transform 1 0 8288 0 1 370
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_3
timestamp 1698431365
transform 1 0 18241 0 1 395
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_4
timestamp 1698431365
transform 1 0 6094 0 1 368
box 0 0 1 1
use M1_POLY243105905487104_128x8m81  M1_POLY243105905487104_128x8m81_0
timestamp 1698431365
transform 1 0 21219 0 1 516
box 0 0 1 1
use M1_POLY243105905487104_128x8m81  M1_POLY243105905487104_128x8m81_1
timestamp 1698431365
transform 1 0 3114 0 1 546
box 0 0 1 1
use M1_PSUB$$45111340_128x8m81  M1_PSUB$$45111340_128x8m81_0
timestamp 1698431365
transform -1 0 19779 0 1 0
box 0 0 1 1
use M1_PSUB$$49279020_128x8m81  M1_PSUB$$49279020_128x8m81_0
timestamp 1698431365
transform 1 0 11483 0 1 900
box 0 0 1 1
use M2_M1$$45004844_128x8m81  M2_M1$$45004844_128x8m81_0
timestamp 1698431365
transform 1 0 20179 0 1 900
box 0 0 1 1
use M2_M1$$46894124_128x8m81  M2_M1$$46894124_128x8m81_0
timestamp 1698431365
transform 1 0 6300 0 1 363
box 0 0 1 1
use M2_M1$$201262124_128x8m81  M2_M1$$201262124_128x8m81_0
timestamp 1698431365
transform 1 0 14667 0 1 438
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_0
timestamp 1698431365
transform 1 0 6300 0 1 363
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_1
timestamp 1698431365
transform 1 0 9397 0 1 662
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_0
timestamp 1698431365
transform 1 0 18218 0 1 385
box 0 0 1 1
use M2_M1$$204402732_128x8m81  M2_M1$$204402732_128x8m81_0
timestamp 1698431365
transform 1 0 22887 0 1 0
box 0 0 1 1
use M2_M1$$204402732_128x8m81  M2_M1$$204402732_128x8m81_1
timestamp 1698431365
transform 1 0 22887 0 1 900
box 0 0 1 1
use M2_M1$$204402732_128x8m81  M2_M1$$204402732_128x8m81_2
timestamp 1698431365
transform 1 0 1425 0 1 0
box 0 0 1 1
use M2_M1$$204402732_128x8m81  M2_M1$$204402732_128x8m81_3
timestamp 1698431365
transform 1 0 1425 0 1 900
box 0 0 1 1
use M2_M1$$204403756_128x8m81  M2_M1$$204403756_128x8m81_0
timestamp 1698431365
transform 1 0 7603 0 1 610
box 0 0 1 1
use M2_M1$$204403756_128x8m81  M2_M1$$204403756_128x8m81_1
timestamp 1698431365
transform 1 0 9965 0 1 900
box 0 0 1 1
use M2_M1$$204403756_128x8m81  M2_M1$$204403756_128x8m81_2
timestamp 1698431365
transform 1 0 21547 0 1 669
box 0 0 1 1
use M2_M1$$204403756_128x8m81  M2_M1$$204403756_128x8m81_3
timestamp 1698431365
transform 1 0 19850 0 1 0
box 0 0 1 1
use M2_M1$$204403756_128x8m81  M2_M1$$204403756_128x8m81_4
timestamp 1698431365
transform 1 0 8764 0 1 900
box 0 0 1 1
use M2_M1$$204403756_128x8m81  M2_M1$$204403756_128x8m81_5
timestamp 1698431365
transform 1 0 4467 0 1 0
box 0 0 1 1
use M2_M1$$204403756_128x8m81  M2_M1$$204403756_128x8m81_6
timestamp 1698431365
transform 1 0 7603 0 1 136
box 0 0 1 1
use M2_M1$$204403756_128x8m81  M2_M1$$204403756_128x8m81_7
timestamp 1698431365
transform 1 0 20785 0 1 676
box 0 0 1 1
use M2_M1$$204403756_128x8m81  M2_M1$$204403756_128x8m81_8
timestamp 1698431365
transform 1 0 2769 0 1 676
box 0 0 1 1
use M2_M1$$204403756_128x8m81  M2_M1$$204403756_128x8m81_9
timestamp 1698431365
transform 1 0 2769 0 1 228
box 0 0 1 1
use M2_M1$$204403756_128x8m81  M2_M1$$204403756_128x8m81_10
timestamp 1698431365
transform 1 0 3531 0 1 684
box 0 0 1 1
use M2_M1$$204403756_128x8m81  M2_M1$$204403756_128x8m81_11
timestamp 1698431365
transform 1 0 21547 0 1 206
box 0 0 1 1
use M2_M1$$204403756_R270_128x8m81  M2_M1$$204403756_R270_128x8m81_0
timestamp 1698431365
transform 0 -1 9616 1 0 354
box 0 0 1 1
use M2_M1$$204404780_128x8m81  M2_M1$$204404780_128x8m81_0
timestamp 1698431365
transform 1 0 13729 0 1 900
box 0 0 1 1
use M2_M1$$204404780_128x8m81  M2_M1$$204404780_128x8m81_1
timestamp 1698431365
transform 1 0 4223 0 1 900
box 0 0 1 1
use M2_M1$$204404780_128x8m81  M2_M1$$204404780_128x8m81_2
timestamp 1698431365
transform 1 0 6900 0 1 370
box 0 0 1 1
use M2_M1$$204405804_128x8m81  M2_M1$$204405804_128x8m81_0
timestamp 1698431365
transform 1 0 4069 0 1 438
box 0 0 1 1
use M2_M1$$204406828_128x8m81  M2_M1$$204406828_128x8m81_0
timestamp 1698431365
transform 1 0 18987 0 1 900
box 0 0 1 1
use M2_M1$$204406828_128x8m81  M2_M1$$204406828_128x8m81_1
timestamp 1698431365
transform 1 0 5369 0 1 900
box 0 0 1 1
use M2_M1$$204407852_128x8m81  M2_M1$$204407852_128x8m81_0
timestamp 1698431365
transform 1 0 5376 0 1 598
box 0 0 1 1
use M2_M1$$204407852_128x8m81  M2_M1$$204407852_128x8m81_1
timestamp 1698431365
transform 1 0 5376 0 1 138
box 0 0 1 1
use M2_M1$$204407852_128x8m81  M2_M1$$204407852_128x8m81_2
timestamp 1698431365
transform 1 0 18987 0 1 601
box 0 0 1 1
use M2_M1$$204407852_128x8m81  M2_M1$$204407852_128x8m81_3
timestamp 1698431365
transform 1 0 18987 0 1 138
box 0 0 1 1
use M2_M1$$204408876_128x8m81  M2_M1$$204408876_128x8m81_0
timestamp 1698431365
transform 1 0 14667 0 1 900
box 0 0 1 1
use M2_M1$$204408876_128x8m81  M2_M1$$204408876_128x8m81_1
timestamp 1698431365
transform 1 0 20133 0 1 438
box 0 0 1 1
use M2_M1$$204408876_128x8m81  M2_M1$$204408876_128x8m81_2
timestamp 1698431365
transform 1 0 8163 0 1 900
box 0 0 1 1
use M3_M2$$201251884_128x8m81  M3_M2$$201251884_128x8m81_0
timestamp 1698431365
transform 1 0 20102 0 1 0
box 0 0 1 1
use M3_M2$$201251884_128x8m81  M3_M2$$201251884_128x8m81_1
timestamp 1698431365
transform 1 0 13729 0 1 0
box 0 0 1 1
use M3_M2$$201251884_128x8m81  M3_M2$$201251884_128x8m81_2
timestamp 1698431365
transform 1 0 4223 0 1 0
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_0
timestamp 1698431365
transform 1 0 18218 0 1 385
box 0 0 1 1
use M3_M2$$204147756_128x8m81  M3_M2$$204147756_128x8m81_0
timestamp 1698431365
transform 1 0 14667 0 1 900
box 0 0 1 1
use M3_M2$$204147756_128x8m81  M3_M2$$204147756_128x8m81_1
timestamp 1698431365
transform 1 0 8163 0 1 0
box 0 0 1 1
use M3_M2$$204398636_128x8m81  M3_M2$$204398636_128x8m81_0
timestamp 1698431365
transform 1 0 9616 0 1 508
box 0 0 1 1
use M3_M2$$204398636_128x8m81  M3_M2$$204398636_128x8m81_1
timestamp 1698431365
transform 1 0 6300 0 1 508
box 0 0 1 1
use M3_M2$$204398636_128x8m81  M3_M2$$204398636_128x8m81_2
timestamp 1698431365
transform 1 0 9397 0 1 277
box 0 0 1 1
use M3_M2$$204399660_128x8m81  M3_M2$$204399660_128x8m81_0
timestamp 1698431365
transform 1 0 22887 0 1 900
box 0 0 1 1
use M3_M2$$204399660_128x8m81  M3_M2$$204399660_128x8m81_1
timestamp 1698431365
transform 1 0 1425 0 1 900
box 0 0 1 1
use M3_M2$$204400684_128x8m81  M3_M2$$204400684_128x8m81_0
timestamp 1698431365
transform 1 0 9965 0 1 0
box 0 0 1 1
use M3_M2$$204400684_128x8m81  M3_M2$$204400684_128x8m81_1
timestamp 1698431365
transform 1 0 7603 0 1 277
box 0 0 1 1
use M3_M2$$204400684_128x8m81  M3_M2$$204400684_128x8m81_2
timestamp 1698431365
transform 1 0 2769 0 1 467
box 0 0 1 1
use M3_M2$$204400684_128x8m81  M3_M2$$204400684_128x8m81_3
timestamp 1698431365
transform 1 0 3531 0 1 460
box 0 0 1 1
use M3_M2$$204400684_128x8m81  M3_M2$$204400684_128x8m81_4
timestamp 1698431365
transform 1 0 20785 0 1 460
box 0 0 1 1
use M3_M2$$204400684_128x8m81  M3_M2$$204400684_128x8m81_5
timestamp 1698431365
transform 1 0 8764 0 1 900
box 0 0 1 1
use M3_M2$$204400684_128x8m81  M3_M2$$204400684_128x8m81_6
timestamp 1698431365
transform 1 0 21547 0 1 460
box 0 0 1 1
use M3_M2$$204401708_128x8m81  M3_M2$$204401708_128x8m81_0
timestamp 1698431365
transform 1 0 18987 0 1 900
box 0 0 1 1
use M3_M2$$204401708_128x8m81  M3_M2$$204401708_128x8m81_1
timestamp 1698431365
transform 1 0 5369 0 1 900
box 0 0 1 1
use nmos_1p2$$49277996_R270_128x8m81  nmos_1p2$$49277996_R270_128x8m81_0
timestamp 1698431365
transform 0 -1 9763 1 0 759
box -31 0 -30 1
use nmos_5p043105905487107_128x8m81  nmos_5p043105905487107_128x8m81_0
timestamp 1698431365
transform 0 -1 9326 1 0 193
box 0 0 1 1
use nmos_5p043105905487108_128x8m81  nmos_5p043105905487108_128x8m81_0
timestamp 1698431365
transform 0 -1 4267 -1 0 848
box 0 0 1 1
use nmos_5p043105905487108_128x8m81  nmos_5p043105905487108_128x8m81_1
timestamp 1698431365
transform 0 1 20050 -1 0 848
box 0 0 1 1
use nmos_5p043105905487109_128x8m81  nmos_5p043105905487109_128x8m81_0
timestamp 1698431365
transform 0 -1 8152 1 0 193
box 0 0 1 1
use pmos_1p2$$49270828_R270_128x8m81  pmos_1p2$$49270828_R270_128x8m81_0
timestamp 1698431365
transform 0 -1 2932 1 0 311
box -31 0 -30 1
use pmos_1p2$$49271852_R270_128x8m81  pmos_1p2$$49271852_R270_128x8m81_0
timestamp 1698431365
transform 0 -1 7097 1 0 224
box -31 0 -30 1
use pmos_1p2$$49272876_R270_128x8m81  pmos_1p2$$49272876_R270_128x8m81_0
timestamp 1698431365
transform 0 1 18361 1 0 224
box -31 0 -30 1
use pmos_1p2$$49272876_R270_128x8m81  pmos_1p2$$49272876_R270_128x8m81_1
timestamp 1698431365
transform 0 -1 5956 1 0 224
box -31 0 -30 1
use pmos_5p043105905487103_128x8m81  pmos_5p043105905487103_128x8m81_0
timestamp 1698431365
transform 0 1 21385 1 0 280
box 0 0 1 1
use pmos_5p043105905487105_128x8m81  pmos_5p043105905487105_128x8m81_0
timestamp 1698431365
transform 0 1 14395 1 0 504
box 0 0 1 1
use pmos_5p043105905487105_128x8m81  pmos_5p043105905487105_128x8m81_1
timestamp 1698431365
transform 0 1 14395 1 0 728
box 0 0 1 1
use pmos_5p043105905487105_128x8m81  pmos_5p043105905487105_128x8m81_2
timestamp 1698431365
transform 0 1 14395 1 0 280
box 0 0 1 1
use pmos_5p043105905487110_128x8m81  pmos_5p043105905487110_128x8m81_0
timestamp 1698431365
transform 0 -1 8922 1 0 193
box 0 0 1 1
<< properties >>
string GDS_END 590122
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 572938
<< end >>
