magic
tech gf180mcuD
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 453 1318 1094
<< pwell >>
rect -86 -86 1318 453
<< metal1 >>
rect 0 918 1232 1098
rect 157 430 203 511
rect 30 354 203 430
rect 366 354 418 511
rect 590 443 667 542
rect 805 758 851 918
rect 273 90 319 172
rect 757 90 803 172
rect 1009 136 1090 872
rect 0 -90 1232 90
<< obsm1 >>
rect 58 769 759 815
rect 713 500 759 769
rect 713 454 950 500
rect 713 264 759 454
rect 49 218 759 264
rect 49 136 95 218
rect 497 136 543 218
<< labels >>
rlabel metal1 s 30 354 203 430 6 A1
port 1 nsew default input
rlabel metal1 s 157 430 203 511 6 A1
port 1 nsew default input
rlabel metal1 s 366 354 418 511 6 A2
port 2 nsew default input
rlabel metal1 s 590 443 667 542 6 A3
port 3 nsew default input
rlabel metal1 s 1009 136 1090 872 6 Z
port 4 nsew default output
rlabel metal1 s 805 758 851 918 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 918 1232 1098 6 VDD
port 5 nsew power bidirectional abutment
rlabel nwell s -86 453 1318 1094 6 VNW
port 6 nsew power bidirectional
rlabel pwell s -86 -86 1318 453 6 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 0 -90 1232 90 8 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 757 90 803 172 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 172 6 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1232 1008
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 278678
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 275220
<< end >>
