magic
tech gf180mcuB
magscale 1 10
timestamp 1698431365
<< metal1 >>
rect 3 3062 203 3074
rect 3 3010 15 3062
rect 67 3010 139 3062
rect 191 3010 203 3062
rect 3 2938 203 3010
rect 3 2886 15 2938
rect 67 2886 139 2938
rect 191 2886 203 2938
rect 3 2814 203 2886
rect 3 2762 15 2814
rect 67 2762 139 2814
rect 191 2762 203 2814
rect 3 2690 203 2762
rect 3 2638 15 2690
rect 67 2638 139 2690
rect 191 2638 203 2690
rect 3 2566 203 2638
rect 3 2514 15 2566
rect 67 2514 139 2566
rect 191 2514 203 2566
rect 3 2442 203 2514
rect 3 2390 15 2442
rect 67 2390 139 2442
rect 191 2390 203 2442
rect 3 2318 203 2390
rect 3 2266 15 2318
rect 67 2266 139 2318
rect 191 2266 203 2318
rect 3 2194 203 2266
rect 3 2142 15 2194
rect 67 2142 139 2194
rect 191 2142 203 2194
rect 3 2130 203 2142
rect 1020 3062 1220 3074
rect 1020 3010 1032 3062
rect 1084 3010 1156 3062
rect 1208 3010 1220 3062
rect 1020 2938 1220 3010
rect 1020 2886 1032 2938
rect 1084 2886 1156 2938
rect 1208 2886 1220 2938
rect 1020 2814 1220 2886
rect 1020 2762 1032 2814
rect 1084 2762 1156 2814
rect 1208 2762 1220 2814
rect 1020 2690 1220 2762
rect 1020 2638 1032 2690
rect 1084 2638 1156 2690
rect 1208 2638 1220 2690
rect 1020 2566 1220 2638
rect 1020 2514 1032 2566
rect 1084 2514 1156 2566
rect 1208 2514 1220 2566
rect 1020 2442 1220 2514
rect 1020 2390 1032 2442
rect 1084 2390 1156 2442
rect 1208 2390 1220 2442
rect 1020 2318 1220 2390
rect 1020 2266 1032 2318
rect 1084 2266 1156 2318
rect 1208 2266 1220 2318
rect 1020 2194 1220 2266
rect 1020 2142 1032 2194
rect 1084 2142 1156 2194
rect 1208 2142 1220 2194
rect 1020 2130 1220 2142
<< via1 >>
rect 15 3010 67 3062
rect 139 3010 191 3062
rect 15 2886 67 2938
rect 139 2886 191 2938
rect 15 2762 67 2814
rect 139 2762 191 2814
rect 15 2638 67 2690
rect 139 2638 191 2690
rect 15 2514 67 2566
rect 139 2514 191 2566
rect 15 2390 67 2442
rect 139 2390 191 2442
rect 15 2266 67 2318
rect 139 2266 191 2318
rect 15 2142 67 2194
rect 139 2142 191 2194
rect 1032 3010 1084 3062
rect 1156 3010 1208 3062
rect 1032 2886 1084 2938
rect 1156 2886 1208 2938
rect 1032 2762 1084 2814
rect 1156 2762 1208 2814
rect 1032 2638 1084 2690
rect 1156 2638 1208 2690
rect 1032 2514 1084 2566
rect 1156 2514 1208 2566
rect 1032 2390 1084 2442
rect 1156 2390 1208 2442
rect 1032 2266 1084 2318
rect 1156 2266 1208 2318
rect 1032 2142 1084 2194
rect 1156 2142 1208 2194
<< metal2 >>
rect 495 6267 719 7462
rect 495 6211 516 6267
rect 572 6211 640 6267
rect 696 6211 719 6267
rect 495 6143 719 6211
rect 495 6087 516 6143
rect 572 6087 640 6143
rect 696 6087 719 6143
rect 495 6019 719 6087
rect 495 5963 516 6019
rect 572 5963 640 6019
rect 696 5963 719 6019
rect -8 4667 216 5604
rect -8 4611 16 4667
rect 72 4611 140 4667
rect 196 4611 216 4667
rect -8 4543 216 4611
rect -8 4487 16 4543
rect 72 4487 140 4543
rect 196 4487 216 4543
rect -8 4419 216 4487
rect -8 4363 16 4419
rect 72 4363 140 4419
rect 196 4363 216 4419
rect -8 3062 216 4363
rect 495 4009 719 5963
rect 495 3953 516 4009
rect 572 3953 640 4009
rect 696 3953 719 4009
rect 495 3885 719 3953
rect 495 3829 516 3885
rect 572 3829 640 3885
rect 696 3829 719 3885
rect 495 3761 719 3829
rect 495 3705 516 3761
rect 572 3705 640 3761
rect 696 3705 719 3761
rect 495 3637 719 3705
rect 495 3581 516 3637
rect 572 3581 640 3637
rect 696 3581 719 3637
rect 495 3513 719 3581
rect 495 3457 516 3513
rect 572 3457 640 3513
rect 696 3457 719 3513
rect 495 3389 719 3457
rect 495 3333 516 3389
rect 572 3333 640 3389
rect 696 3333 719 3389
rect 495 3265 719 3333
rect 495 3209 516 3265
rect 572 3209 640 3265
rect 696 3209 719 3265
rect 495 3065 719 3209
rect 1011 4667 1235 5605
rect 1011 4611 1033 4667
rect 1089 4611 1157 4667
rect 1213 4611 1235 4667
rect 1011 4543 1235 4611
rect 1011 4487 1033 4543
rect 1089 4487 1157 4543
rect 1213 4487 1235 4543
rect 1011 4419 1235 4487
rect 1011 4363 1033 4419
rect 1089 4363 1157 4419
rect 1213 4363 1235 4419
rect -8 3010 15 3062
rect 67 3010 139 3062
rect 191 3010 216 3062
rect -8 2938 216 3010
rect -8 2886 15 2938
rect 67 2886 139 2938
rect 191 2886 216 2938
rect -8 2814 216 2886
rect -8 2762 15 2814
rect 67 2762 139 2814
rect 191 2762 216 2814
rect -8 2690 216 2762
rect -8 2638 15 2690
rect 67 2638 139 2690
rect 191 2638 216 2690
rect -8 2566 216 2638
rect -8 2514 15 2566
rect 67 2514 139 2566
rect 191 2514 216 2566
rect -8 2442 216 2514
rect -8 2390 15 2442
rect 67 2390 139 2442
rect 191 2390 216 2442
rect -8 2318 216 2390
rect -8 2266 15 2318
rect 67 2266 139 2318
rect 191 2266 216 2318
rect -8 2194 216 2266
rect -8 2142 15 2194
rect 67 2142 139 2194
rect 191 2142 216 2194
rect -8 2115 216 2142
rect 1011 3062 1235 4363
rect 1011 3010 1032 3062
rect 1084 3010 1156 3062
rect 1208 3010 1235 3062
rect 1011 2938 1235 3010
rect 1011 2886 1032 2938
rect 1084 2886 1156 2938
rect 1208 2886 1235 2938
rect 1011 2814 1235 2886
rect 1011 2762 1032 2814
rect 1084 2762 1156 2814
rect 1208 2762 1235 2814
rect 1011 2690 1235 2762
rect 1011 2638 1032 2690
rect 1084 2638 1156 2690
rect 1208 2638 1235 2690
rect 1011 2566 1235 2638
rect 1011 2514 1032 2566
rect 1084 2514 1156 2566
rect 1208 2514 1235 2566
rect 1011 2442 1235 2514
rect 1011 2390 1032 2442
rect 1084 2390 1156 2442
rect 1208 2390 1235 2442
rect 1011 2318 1235 2390
rect 1011 2266 1032 2318
rect 1084 2266 1156 2318
rect 1208 2266 1235 2318
rect 1011 2194 1235 2266
rect 1011 2142 1032 2194
rect 1084 2142 1156 2194
rect 1208 2142 1235 2194
rect 1011 2115 1235 2142
<< via2 >>
rect 516 6211 572 6267
rect 640 6211 696 6267
rect 516 6087 572 6143
rect 640 6087 696 6143
rect 516 5963 572 6019
rect 640 5963 696 6019
rect 16 4611 72 4667
rect 140 4611 196 4667
rect 16 4487 72 4543
rect 140 4487 196 4543
rect 16 4363 72 4419
rect 140 4363 196 4419
rect 516 3953 572 4009
rect 640 3953 696 4009
rect 516 3829 572 3885
rect 640 3829 696 3885
rect 516 3705 572 3761
rect 640 3705 696 3761
rect 516 3581 572 3637
rect 640 3581 696 3637
rect 516 3457 572 3513
rect 640 3457 696 3513
rect 516 3333 572 3389
rect 640 3333 696 3389
rect 516 3209 572 3265
rect 640 3209 696 3265
rect 1033 4611 1089 4667
rect 1157 4611 1213 4667
rect 1033 4487 1089 4543
rect 1157 4487 1213 4543
rect 1033 4363 1089 4419
rect 1157 4363 1213 4419
<< metal3 >>
rect 506 6267 706 6277
rect 506 6211 516 6267
rect 572 6211 640 6267
rect 696 6211 706 6267
rect 506 6143 706 6211
rect 506 6087 516 6143
rect 572 6087 640 6143
rect 696 6087 706 6143
rect 506 6019 706 6087
rect 506 5963 516 6019
rect 572 5963 640 6019
rect 696 5963 706 6019
rect 506 5953 706 5963
rect 6 4667 206 4677
rect 6 4611 16 4667
rect 72 4611 140 4667
rect 196 4611 206 4667
rect 6 4543 206 4611
rect 6 4487 16 4543
rect 72 4487 140 4543
rect 196 4487 206 4543
rect 6 4419 206 4487
rect 6 4363 16 4419
rect 72 4363 140 4419
rect 196 4363 206 4419
rect 6 4353 206 4363
rect 1023 4667 1223 4677
rect 1023 4611 1033 4667
rect 1089 4611 1157 4667
rect 1213 4611 1223 4667
rect 1023 4543 1223 4611
rect 1023 4487 1033 4543
rect 1089 4487 1157 4543
rect 1213 4487 1223 4543
rect 1023 4419 1223 4487
rect 1023 4363 1033 4419
rect 1089 4363 1157 4419
rect 1213 4363 1223 4419
rect 1023 4353 1223 4363
rect 506 4009 706 4019
rect 506 3953 516 4009
rect 572 3953 640 4009
rect 696 3953 706 4009
rect 506 3885 706 3953
rect 506 3829 516 3885
rect 572 3829 640 3885
rect 696 3829 706 3885
rect 506 3761 706 3829
rect 506 3705 516 3761
rect 572 3705 640 3761
rect 696 3705 706 3761
rect 506 3637 706 3705
rect 506 3581 516 3637
rect 572 3581 640 3637
rect 696 3581 706 3637
rect 506 3513 706 3581
rect 506 3457 516 3513
rect 572 3457 640 3513
rect 696 3457 706 3513
rect 506 3389 706 3457
rect 506 3333 516 3389
rect 572 3333 640 3389
rect 696 3333 706 3389
rect 506 3265 706 3333
rect 506 3209 516 3265
rect 572 3209 640 3265
rect 696 3209 706 3265
rect 506 3199 706 3209
use M2_M14310590878176_256x8m81  M2_M14310590878176_256x8m81_0
timestamp 1698431365
transform 1 0 1120 0 1 2602
box 0 0 1 1
use M2_M14310590878176_256x8m81  M2_M14310590878176_256x8m81_1
timestamp 1698431365
transform 1 0 103 0 1 2602
box 0 0 1 1
use M3_M24310590878171_256x8m81  M3_M24310590878171_256x8m81_0
timestamp 1698431365
transform 1 0 606 0 1 6115
box 0 0 1 1
use M3_M24310590878171_256x8m81  M3_M24310590878171_256x8m81_1
timestamp 1698431365
transform 1 0 1123 0 1 4515
box 0 0 1 1
use M3_M24310590878171_256x8m81  M3_M24310590878171_256x8m81_2
timestamp 1698431365
transform 1 0 106 0 1 4515
box 0 0 1 1
use M3_M24310590878196_256x8m81  M3_M24310590878196_256x8m81_0
timestamp 1698431365
transform 1 0 606 0 1 3609
box 0 0 1 1
<< properties >>
string GDS_END 1887046
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 1886568
string path 5.615 28.025 5.615 10.575 
<< end >>
