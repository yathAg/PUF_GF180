magic
tech gf180mcuD
magscale 1 10
timestamp 1698431365
<< psubdiff >>
rect 70 46083 85816 46102
rect 70 46037 89 46083
rect 135 46037 213 46083
rect 259 46037 337 46083
rect 383 46037 461 46083
rect 507 46037 585 46083
rect 631 46037 709 46083
rect 755 46037 833 46083
rect 879 46037 957 46083
rect 1003 46037 1081 46083
rect 1127 46037 1205 46083
rect 1251 46037 1329 46083
rect 1375 46037 1453 46083
rect 1499 46037 1577 46083
rect 1623 46037 1701 46083
rect 1747 46037 1825 46083
rect 1871 46037 1949 46083
rect 1995 46037 2073 46083
rect 2119 46037 2197 46083
rect 2243 46037 2321 46083
rect 2367 46037 2445 46083
rect 2491 46037 2569 46083
rect 2615 46037 2693 46083
rect 2739 46037 2817 46083
rect 2863 46037 2941 46083
rect 2987 46037 3065 46083
rect 3111 46037 3189 46083
rect 3235 46037 3313 46083
rect 3359 46037 3437 46083
rect 3483 46037 3561 46083
rect 3607 46037 3685 46083
rect 3731 46037 3809 46083
rect 3855 46037 3933 46083
rect 3979 46037 4057 46083
rect 4103 46037 4181 46083
rect 4227 46037 4305 46083
rect 4351 46037 4429 46083
rect 4475 46037 4553 46083
rect 4599 46037 4677 46083
rect 4723 46037 4801 46083
rect 4847 46037 4925 46083
rect 4971 46037 5049 46083
rect 5095 46037 5173 46083
rect 5219 46037 5297 46083
rect 5343 46037 5421 46083
rect 5467 46037 5545 46083
rect 5591 46037 5669 46083
rect 5715 46037 5793 46083
rect 5839 46037 5917 46083
rect 5963 46037 6041 46083
rect 6087 46037 6165 46083
rect 6211 46037 6289 46083
rect 6335 46037 6413 46083
rect 6459 46037 6537 46083
rect 6583 46037 6661 46083
rect 6707 46037 6785 46083
rect 6831 46037 6909 46083
rect 6955 46037 7033 46083
rect 7079 46037 7157 46083
rect 7203 46037 7281 46083
rect 7327 46037 7405 46083
rect 7451 46037 7529 46083
rect 7575 46037 7653 46083
rect 7699 46037 7777 46083
rect 7823 46037 7901 46083
rect 7947 46037 8025 46083
rect 8071 46037 8149 46083
rect 8195 46037 8273 46083
rect 8319 46037 8397 46083
rect 8443 46037 8521 46083
rect 8567 46037 8645 46083
rect 8691 46037 8769 46083
rect 8815 46037 8893 46083
rect 8939 46037 9017 46083
rect 9063 46037 9141 46083
rect 9187 46037 9265 46083
rect 9311 46037 9389 46083
rect 9435 46037 9513 46083
rect 9559 46037 9637 46083
rect 9683 46037 9761 46083
rect 9807 46037 9885 46083
rect 9931 46037 10009 46083
rect 10055 46037 10133 46083
rect 10179 46037 10257 46083
rect 10303 46037 10381 46083
rect 10427 46037 10505 46083
rect 10551 46037 10629 46083
rect 10675 46037 10753 46083
rect 10799 46037 10877 46083
rect 10923 46037 11001 46083
rect 11047 46037 11125 46083
rect 11171 46037 11249 46083
rect 11295 46037 11373 46083
rect 11419 46037 11497 46083
rect 11543 46037 11621 46083
rect 11667 46037 11745 46083
rect 11791 46037 11869 46083
rect 11915 46037 11993 46083
rect 12039 46037 12117 46083
rect 12163 46037 12241 46083
rect 12287 46037 12365 46083
rect 12411 46037 12489 46083
rect 12535 46037 12613 46083
rect 12659 46037 12737 46083
rect 12783 46037 12861 46083
rect 12907 46037 12985 46083
rect 13031 46037 13109 46083
rect 13155 46037 13233 46083
rect 13279 46037 13357 46083
rect 13403 46037 13481 46083
rect 13527 46037 13605 46083
rect 13651 46037 13729 46083
rect 13775 46037 13853 46083
rect 13899 46037 13977 46083
rect 14023 46037 14101 46083
rect 14147 46037 14225 46083
rect 14271 46037 14349 46083
rect 14395 46037 14473 46083
rect 14519 46037 14597 46083
rect 14643 46037 14721 46083
rect 14767 46037 14845 46083
rect 14891 46037 14969 46083
rect 15015 46037 15093 46083
rect 15139 46037 15217 46083
rect 15263 46037 15341 46083
rect 15387 46037 15465 46083
rect 15511 46037 15589 46083
rect 15635 46037 15713 46083
rect 15759 46037 15837 46083
rect 15883 46037 15961 46083
rect 16007 46037 16085 46083
rect 16131 46037 16209 46083
rect 16255 46037 16333 46083
rect 16379 46037 16457 46083
rect 16503 46037 16581 46083
rect 16627 46037 16705 46083
rect 16751 46037 16829 46083
rect 16875 46037 16953 46083
rect 16999 46037 17077 46083
rect 17123 46037 17201 46083
rect 17247 46037 17325 46083
rect 17371 46037 17449 46083
rect 17495 46037 17573 46083
rect 17619 46037 17697 46083
rect 17743 46037 17821 46083
rect 17867 46037 17945 46083
rect 17991 46037 18069 46083
rect 18115 46037 18193 46083
rect 18239 46037 18317 46083
rect 18363 46037 18441 46083
rect 18487 46037 18565 46083
rect 18611 46037 18689 46083
rect 18735 46037 18813 46083
rect 18859 46037 18937 46083
rect 18983 46037 19061 46083
rect 19107 46037 19185 46083
rect 19231 46037 19309 46083
rect 19355 46037 19433 46083
rect 19479 46037 19557 46083
rect 19603 46037 19681 46083
rect 19727 46037 19805 46083
rect 19851 46037 19929 46083
rect 19975 46037 20053 46083
rect 20099 46037 20177 46083
rect 20223 46037 20301 46083
rect 20347 46037 20425 46083
rect 20471 46037 20549 46083
rect 20595 46037 20673 46083
rect 20719 46037 20797 46083
rect 20843 46037 20921 46083
rect 20967 46037 21045 46083
rect 21091 46037 21169 46083
rect 21215 46037 21293 46083
rect 21339 46037 21417 46083
rect 21463 46037 21541 46083
rect 21587 46037 21665 46083
rect 21711 46037 21789 46083
rect 21835 46037 21913 46083
rect 21959 46037 22037 46083
rect 22083 46037 22161 46083
rect 22207 46037 22285 46083
rect 22331 46037 22409 46083
rect 22455 46037 22533 46083
rect 22579 46037 22657 46083
rect 22703 46037 22781 46083
rect 22827 46037 22905 46083
rect 22951 46037 23029 46083
rect 23075 46037 23153 46083
rect 23199 46037 23277 46083
rect 23323 46037 23401 46083
rect 23447 46037 23525 46083
rect 23571 46037 23649 46083
rect 23695 46037 23773 46083
rect 23819 46037 23897 46083
rect 23943 46037 24021 46083
rect 24067 46037 24145 46083
rect 24191 46037 24269 46083
rect 24315 46037 24393 46083
rect 24439 46037 24517 46083
rect 24563 46037 24641 46083
rect 24687 46037 24765 46083
rect 24811 46037 24889 46083
rect 24935 46037 25013 46083
rect 25059 46037 25137 46083
rect 25183 46037 25261 46083
rect 25307 46037 25385 46083
rect 25431 46037 25509 46083
rect 25555 46037 25633 46083
rect 25679 46037 25757 46083
rect 25803 46037 25881 46083
rect 25927 46037 26005 46083
rect 26051 46037 26129 46083
rect 26175 46037 26253 46083
rect 26299 46037 26377 46083
rect 26423 46037 26501 46083
rect 26547 46037 26625 46083
rect 26671 46037 26749 46083
rect 26795 46037 26873 46083
rect 26919 46037 26997 46083
rect 27043 46037 27121 46083
rect 27167 46037 27245 46083
rect 27291 46037 27369 46083
rect 27415 46037 27493 46083
rect 27539 46037 27617 46083
rect 27663 46037 27741 46083
rect 27787 46037 27865 46083
rect 27911 46037 27989 46083
rect 28035 46037 28113 46083
rect 28159 46037 28237 46083
rect 28283 46037 28361 46083
rect 28407 46037 28485 46083
rect 28531 46037 28609 46083
rect 28655 46037 28733 46083
rect 28779 46037 28857 46083
rect 28903 46037 28981 46083
rect 29027 46037 29105 46083
rect 29151 46037 29229 46083
rect 29275 46037 29353 46083
rect 29399 46037 29477 46083
rect 29523 46037 29601 46083
rect 29647 46037 29725 46083
rect 29771 46037 29849 46083
rect 29895 46037 29973 46083
rect 30019 46037 30097 46083
rect 30143 46037 30221 46083
rect 30267 46037 30345 46083
rect 30391 46037 30469 46083
rect 30515 46037 30593 46083
rect 30639 46037 30717 46083
rect 30763 46037 30841 46083
rect 30887 46037 30965 46083
rect 31011 46037 31089 46083
rect 31135 46037 31213 46083
rect 31259 46037 31337 46083
rect 31383 46037 31461 46083
rect 31507 46037 31585 46083
rect 31631 46037 31709 46083
rect 31755 46037 31833 46083
rect 31879 46037 31957 46083
rect 32003 46037 32081 46083
rect 32127 46037 32205 46083
rect 32251 46037 32329 46083
rect 32375 46037 32453 46083
rect 32499 46037 32577 46083
rect 32623 46037 32701 46083
rect 32747 46037 32825 46083
rect 32871 46037 32949 46083
rect 32995 46037 33073 46083
rect 33119 46037 33197 46083
rect 33243 46037 33321 46083
rect 33367 46037 33445 46083
rect 33491 46037 33569 46083
rect 33615 46037 33693 46083
rect 33739 46037 33817 46083
rect 33863 46037 33941 46083
rect 33987 46037 34065 46083
rect 34111 46037 34189 46083
rect 34235 46037 34313 46083
rect 34359 46037 34437 46083
rect 34483 46037 34561 46083
rect 34607 46037 34685 46083
rect 34731 46037 34809 46083
rect 34855 46037 34933 46083
rect 34979 46037 35057 46083
rect 35103 46037 35181 46083
rect 35227 46037 35305 46083
rect 35351 46037 35429 46083
rect 35475 46037 35553 46083
rect 35599 46037 35677 46083
rect 35723 46037 35801 46083
rect 35847 46037 35925 46083
rect 35971 46037 36049 46083
rect 36095 46037 36173 46083
rect 36219 46037 36297 46083
rect 36343 46037 36421 46083
rect 36467 46037 36545 46083
rect 36591 46037 36669 46083
rect 36715 46037 36793 46083
rect 36839 46037 36917 46083
rect 36963 46037 37041 46083
rect 37087 46037 37165 46083
rect 37211 46037 37289 46083
rect 37335 46037 37413 46083
rect 37459 46037 37537 46083
rect 37583 46037 37661 46083
rect 37707 46037 37785 46083
rect 37831 46037 37909 46083
rect 37955 46037 38033 46083
rect 38079 46037 38157 46083
rect 38203 46037 38281 46083
rect 38327 46037 38405 46083
rect 38451 46037 38529 46083
rect 38575 46037 38653 46083
rect 38699 46037 38777 46083
rect 38823 46037 38901 46083
rect 38947 46037 39025 46083
rect 39071 46037 39149 46083
rect 39195 46037 39273 46083
rect 39319 46037 39397 46083
rect 39443 46037 39521 46083
rect 39567 46037 39645 46083
rect 39691 46037 39769 46083
rect 39815 46037 39893 46083
rect 39939 46037 40017 46083
rect 40063 46037 40141 46083
rect 40187 46037 40265 46083
rect 40311 46037 40389 46083
rect 40435 46037 40513 46083
rect 40559 46037 40637 46083
rect 40683 46037 40761 46083
rect 40807 46037 40885 46083
rect 40931 46037 41009 46083
rect 41055 46037 41133 46083
rect 41179 46037 41257 46083
rect 41303 46037 41381 46083
rect 41427 46037 41505 46083
rect 41551 46037 41629 46083
rect 41675 46037 41753 46083
rect 41799 46037 41877 46083
rect 41923 46037 42001 46083
rect 42047 46037 42125 46083
rect 42171 46037 42249 46083
rect 42295 46037 42373 46083
rect 42419 46037 42497 46083
rect 42543 46037 42621 46083
rect 42667 46037 42745 46083
rect 42791 46037 42869 46083
rect 42915 46037 42993 46083
rect 43039 46037 43117 46083
rect 43163 46037 43241 46083
rect 43287 46037 43365 46083
rect 43411 46037 43489 46083
rect 43535 46037 43613 46083
rect 43659 46037 43737 46083
rect 43783 46037 43861 46083
rect 43907 46037 43985 46083
rect 44031 46037 44109 46083
rect 44155 46037 44233 46083
rect 44279 46037 44357 46083
rect 44403 46037 44481 46083
rect 44527 46037 44605 46083
rect 44651 46037 44729 46083
rect 44775 46037 44853 46083
rect 44899 46037 44977 46083
rect 45023 46037 45101 46083
rect 45147 46037 45225 46083
rect 45271 46037 45349 46083
rect 45395 46037 45473 46083
rect 45519 46037 45597 46083
rect 45643 46037 45721 46083
rect 45767 46037 45845 46083
rect 45891 46037 45969 46083
rect 46015 46037 46093 46083
rect 46139 46037 46217 46083
rect 46263 46037 46341 46083
rect 46387 46037 46465 46083
rect 46511 46037 46589 46083
rect 46635 46037 46713 46083
rect 46759 46037 46837 46083
rect 46883 46037 46961 46083
rect 47007 46037 47085 46083
rect 47131 46037 47209 46083
rect 47255 46037 47333 46083
rect 47379 46037 47457 46083
rect 47503 46037 47581 46083
rect 47627 46037 47705 46083
rect 47751 46037 47829 46083
rect 47875 46037 47953 46083
rect 47999 46037 48077 46083
rect 48123 46037 48201 46083
rect 48247 46037 48325 46083
rect 48371 46037 48449 46083
rect 48495 46037 48573 46083
rect 48619 46037 48697 46083
rect 48743 46037 48821 46083
rect 48867 46037 48945 46083
rect 48991 46037 49069 46083
rect 49115 46037 49193 46083
rect 49239 46037 49317 46083
rect 49363 46037 49441 46083
rect 49487 46037 49565 46083
rect 49611 46037 49689 46083
rect 49735 46037 49813 46083
rect 49859 46037 49937 46083
rect 49983 46037 50061 46083
rect 50107 46037 50185 46083
rect 50231 46037 50309 46083
rect 50355 46037 50433 46083
rect 50479 46037 50557 46083
rect 50603 46037 50681 46083
rect 50727 46037 50805 46083
rect 50851 46037 50929 46083
rect 50975 46037 51053 46083
rect 51099 46037 51177 46083
rect 51223 46037 51301 46083
rect 51347 46037 51425 46083
rect 51471 46037 51549 46083
rect 51595 46037 51673 46083
rect 51719 46037 51797 46083
rect 51843 46037 51921 46083
rect 51967 46037 52045 46083
rect 52091 46037 52169 46083
rect 52215 46037 52293 46083
rect 52339 46037 52417 46083
rect 52463 46037 52541 46083
rect 52587 46037 52665 46083
rect 52711 46037 52789 46083
rect 52835 46037 52913 46083
rect 52959 46037 53037 46083
rect 53083 46037 53161 46083
rect 53207 46037 53285 46083
rect 53331 46037 53409 46083
rect 53455 46037 53533 46083
rect 53579 46037 53657 46083
rect 53703 46037 53781 46083
rect 53827 46037 53905 46083
rect 53951 46037 54029 46083
rect 54075 46037 54153 46083
rect 54199 46037 54277 46083
rect 54323 46037 54401 46083
rect 54447 46037 54525 46083
rect 54571 46037 54649 46083
rect 54695 46037 54773 46083
rect 54819 46037 54897 46083
rect 54943 46037 55021 46083
rect 55067 46037 55145 46083
rect 55191 46037 55269 46083
rect 55315 46037 55393 46083
rect 55439 46037 55517 46083
rect 55563 46037 55641 46083
rect 55687 46037 55765 46083
rect 55811 46037 55889 46083
rect 55935 46037 56013 46083
rect 56059 46037 56137 46083
rect 56183 46037 56261 46083
rect 56307 46037 56385 46083
rect 56431 46037 56509 46083
rect 56555 46037 56633 46083
rect 56679 46037 56757 46083
rect 56803 46037 56881 46083
rect 56927 46037 57005 46083
rect 57051 46037 57129 46083
rect 57175 46037 57253 46083
rect 57299 46037 57377 46083
rect 57423 46037 57501 46083
rect 57547 46037 57625 46083
rect 57671 46037 57749 46083
rect 57795 46037 57873 46083
rect 57919 46037 57997 46083
rect 58043 46037 58121 46083
rect 58167 46037 58245 46083
rect 58291 46037 58369 46083
rect 58415 46037 58493 46083
rect 58539 46037 58617 46083
rect 58663 46037 58741 46083
rect 58787 46037 58865 46083
rect 58911 46037 58989 46083
rect 59035 46037 59113 46083
rect 59159 46037 59237 46083
rect 59283 46037 59361 46083
rect 59407 46037 59485 46083
rect 59531 46037 59609 46083
rect 59655 46037 59733 46083
rect 59779 46037 59857 46083
rect 59903 46037 59981 46083
rect 60027 46037 60105 46083
rect 60151 46037 60229 46083
rect 60275 46037 60353 46083
rect 60399 46037 60477 46083
rect 60523 46037 60601 46083
rect 60647 46037 60725 46083
rect 60771 46037 60849 46083
rect 60895 46037 60973 46083
rect 61019 46037 61097 46083
rect 61143 46037 61221 46083
rect 61267 46037 61345 46083
rect 61391 46037 61469 46083
rect 61515 46037 61593 46083
rect 61639 46037 61717 46083
rect 61763 46037 61841 46083
rect 61887 46037 61965 46083
rect 62011 46037 62089 46083
rect 62135 46037 62213 46083
rect 62259 46037 62337 46083
rect 62383 46037 62461 46083
rect 62507 46037 62585 46083
rect 62631 46037 62709 46083
rect 62755 46037 62833 46083
rect 62879 46037 62957 46083
rect 63003 46037 63081 46083
rect 63127 46037 63205 46083
rect 63251 46037 63329 46083
rect 63375 46037 63453 46083
rect 63499 46037 63577 46083
rect 63623 46037 63701 46083
rect 63747 46037 63825 46083
rect 63871 46037 63949 46083
rect 63995 46037 64073 46083
rect 64119 46037 64197 46083
rect 64243 46037 64321 46083
rect 64367 46037 64445 46083
rect 64491 46037 64569 46083
rect 64615 46037 64693 46083
rect 64739 46037 64817 46083
rect 64863 46037 64941 46083
rect 64987 46037 65065 46083
rect 65111 46037 65189 46083
rect 65235 46037 65313 46083
rect 65359 46037 65437 46083
rect 65483 46037 65561 46083
rect 65607 46037 65685 46083
rect 65731 46037 65809 46083
rect 65855 46037 65933 46083
rect 65979 46037 66057 46083
rect 66103 46037 66181 46083
rect 66227 46037 66305 46083
rect 66351 46037 66429 46083
rect 66475 46037 66553 46083
rect 66599 46037 66677 46083
rect 66723 46037 66801 46083
rect 66847 46037 66925 46083
rect 66971 46037 67049 46083
rect 67095 46037 67173 46083
rect 67219 46037 67297 46083
rect 67343 46037 67421 46083
rect 67467 46037 67545 46083
rect 67591 46037 67669 46083
rect 67715 46037 67793 46083
rect 67839 46037 67917 46083
rect 67963 46037 68041 46083
rect 68087 46037 68165 46083
rect 68211 46037 68289 46083
rect 68335 46037 68413 46083
rect 68459 46037 68537 46083
rect 68583 46037 68661 46083
rect 68707 46037 68785 46083
rect 68831 46037 68909 46083
rect 68955 46037 69033 46083
rect 69079 46037 69157 46083
rect 69203 46037 69281 46083
rect 69327 46037 69405 46083
rect 69451 46037 69529 46083
rect 69575 46037 69653 46083
rect 69699 46037 69777 46083
rect 69823 46037 69901 46083
rect 69947 46037 70025 46083
rect 70071 46037 70149 46083
rect 70195 46037 70273 46083
rect 70319 46037 70397 46083
rect 70443 46037 70521 46083
rect 70567 46037 70645 46083
rect 70691 46037 70769 46083
rect 70815 46037 70893 46083
rect 70939 46037 71017 46083
rect 71063 46037 71141 46083
rect 71187 46037 71265 46083
rect 71311 46037 71389 46083
rect 71435 46037 71513 46083
rect 71559 46037 71637 46083
rect 71683 46037 71761 46083
rect 71807 46037 71885 46083
rect 71931 46037 72009 46083
rect 72055 46037 72133 46083
rect 72179 46037 72257 46083
rect 72303 46037 72381 46083
rect 72427 46037 72505 46083
rect 72551 46037 72629 46083
rect 72675 46037 72753 46083
rect 72799 46037 72877 46083
rect 72923 46037 73001 46083
rect 73047 46037 73125 46083
rect 73171 46037 73249 46083
rect 73295 46037 73373 46083
rect 73419 46037 73497 46083
rect 73543 46037 73621 46083
rect 73667 46037 73745 46083
rect 73791 46037 73869 46083
rect 73915 46037 73993 46083
rect 74039 46037 74117 46083
rect 74163 46037 74241 46083
rect 74287 46037 74365 46083
rect 74411 46037 74489 46083
rect 74535 46037 74613 46083
rect 74659 46037 74737 46083
rect 74783 46037 74861 46083
rect 74907 46037 74985 46083
rect 75031 46037 75109 46083
rect 75155 46037 75233 46083
rect 75279 46037 75357 46083
rect 75403 46037 75481 46083
rect 75527 46037 75605 46083
rect 75651 46037 75729 46083
rect 75775 46037 75853 46083
rect 75899 46037 75977 46083
rect 76023 46037 76101 46083
rect 76147 46037 76225 46083
rect 76271 46037 76349 46083
rect 76395 46037 76473 46083
rect 76519 46037 76597 46083
rect 76643 46037 76721 46083
rect 76767 46037 76845 46083
rect 76891 46037 76969 46083
rect 77015 46037 77093 46083
rect 77139 46037 77217 46083
rect 77263 46037 77341 46083
rect 77387 46037 77465 46083
rect 77511 46037 77589 46083
rect 77635 46037 77713 46083
rect 77759 46037 77837 46083
rect 77883 46037 77961 46083
rect 78007 46037 78085 46083
rect 78131 46037 78209 46083
rect 78255 46037 78333 46083
rect 78379 46037 78457 46083
rect 78503 46037 78581 46083
rect 78627 46037 78705 46083
rect 78751 46037 78829 46083
rect 78875 46037 78953 46083
rect 78999 46037 79077 46083
rect 79123 46037 79201 46083
rect 79247 46037 79325 46083
rect 79371 46037 79449 46083
rect 79495 46037 79573 46083
rect 79619 46037 79697 46083
rect 79743 46037 79821 46083
rect 79867 46037 79945 46083
rect 79991 46037 80069 46083
rect 80115 46037 80193 46083
rect 80239 46037 80317 46083
rect 80363 46037 80441 46083
rect 80487 46037 80565 46083
rect 80611 46037 80689 46083
rect 80735 46037 80813 46083
rect 80859 46037 80937 46083
rect 80983 46037 81061 46083
rect 81107 46037 81185 46083
rect 81231 46037 81309 46083
rect 81355 46037 81433 46083
rect 81479 46037 81557 46083
rect 81603 46037 81681 46083
rect 81727 46037 81805 46083
rect 81851 46037 81929 46083
rect 81975 46037 82053 46083
rect 82099 46037 82177 46083
rect 82223 46037 82301 46083
rect 82347 46037 82425 46083
rect 82471 46037 82549 46083
rect 82595 46037 82673 46083
rect 82719 46037 82797 46083
rect 82843 46037 82921 46083
rect 82967 46037 83045 46083
rect 83091 46037 83169 46083
rect 83215 46037 83293 46083
rect 83339 46037 83417 46083
rect 83463 46037 83541 46083
rect 83587 46037 83665 46083
rect 83711 46037 83789 46083
rect 83835 46037 83913 46083
rect 83959 46037 84037 46083
rect 84083 46037 84161 46083
rect 84207 46037 84285 46083
rect 84331 46037 84409 46083
rect 84455 46037 84533 46083
rect 84579 46037 84657 46083
rect 84703 46037 84781 46083
rect 84827 46037 84905 46083
rect 84951 46037 85029 46083
rect 85075 46037 85153 46083
rect 85199 46037 85277 46083
rect 85323 46037 85401 46083
rect 85447 46037 85525 46083
rect 85571 46037 85649 46083
rect 85695 46037 85816 46083
rect 70 45959 85816 46037
rect 70 45913 89 45959
rect 135 45913 213 45959
rect 259 45913 337 45959
rect 383 45913 461 45959
rect 507 45913 585 45959
rect 631 45913 709 45959
rect 755 45913 833 45959
rect 879 45913 957 45959
rect 1003 45913 1081 45959
rect 1127 45913 1205 45959
rect 1251 45913 1329 45959
rect 1375 45913 1453 45959
rect 1499 45913 1577 45959
rect 1623 45913 1701 45959
rect 1747 45913 1825 45959
rect 1871 45913 1949 45959
rect 1995 45913 2073 45959
rect 2119 45913 2197 45959
rect 2243 45913 2321 45959
rect 2367 45913 2445 45959
rect 2491 45913 2569 45959
rect 2615 45913 2693 45959
rect 2739 45913 2817 45959
rect 2863 45913 2941 45959
rect 2987 45913 3065 45959
rect 3111 45913 3189 45959
rect 3235 45913 3313 45959
rect 3359 45913 3437 45959
rect 3483 45913 3561 45959
rect 3607 45913 3685 45959
rect 3731 45913 3809 45959
rect 3855 45913 3933 45959
rect 3979 45913 4057 45959
rect 4103 45913 4181 45959
rect 4227 45913 4305 45959
rect 4351 45913 4429 45959
rect 4475 45913 4553 45959
rect 4599 45913 4677 45959
rect 4723 45913 4801 45959
rect 4847 45913 4925 45959
rect 4971 45913 5049 45959
rect 5095 45913 5173 45959
rect 5219 45913 5297 45959
rect 5343 45913 5421 45959
rect 5467 45913 5545 45959
rect 5591 45913 5669 45959
rect 5715 45913 5793 45959
rect 5839 45913 5917 45959
rect 5963 45913 6041 45959
rect 6087 45913 6165 45959
rect 6211 45913 6289 45959
rect 6335 45913 6413 45959
rect 6459 45913 6537 45959
rect 6583 45913 6661 45959
rect 6707 45913 6785 45959
rect 6831 45913 6909 45959
rect 6955 45913 7033 45959
rect 7079 45913 7157 45959
rect 7203 45913 7281 45959
rect 7327 45913 7405 45959
rect 7451 45913 7529 45959
rect 7575 45913 7653 45959
rect 7699 45913 7777 45959
rect 7823 45913 7901 45959
rect 7947 45913 8025 45959
rect 8071 45913 8149 45959
rect 8195 45913 8273 45959
rect 8319 45913 8397 45959
rect 8443 45913 8521 45959
rect 8567 45913 8645 45959
rect 8691 45913 8769 45959
rect 8815 45913 8893 45959
rect 8939 45913 9017 45959
rect 9063 45913 9141 45959
rect 9187 45913 9265 45959
rect 9311 45913 9389 45959
rect 9435 45913 9513 45959
rect 9559 45913 9637 45959
rect 9683 45913 9761 45959
rect 9807 45913 9885 45959
rect 9931 45913 10009 45959
rect 10055 45913 10133 45959
rect 10179 45913 10257 45959
rect 10303 45913 10381 45959
rect 10427 45913 10505 45959
rect 10551 45913 10629 45959
rect 10675 45913 10753 45959
rect 10799 45913 10877 45959
rect 10923 45913 11001 45959
rect 11047 45913 11125 45959
rect 11171 45913 11249 45959
rect 11295 45913 11373 45959
rect 11419 45913 11497 45959
rect 11543 45913 11621 45959
rect 11667 45913 11745 45959
rect 11791 45913 11869 45959
rect 11915 45913 11993 45959
rect 12039 45913 12117 45959
rect 12163 45913 12241 45959
rect 12287 45913 12365 45959
rect 12411 45913 12489 45959
rect 12535 45913 12613 45959
rect 12659 45913 12737 45959
rect 12783 45913 12861 45959
rect 12907 45913 12985 45959
rect 13031 45913 13109 45959
rect 13155 45913 13233 45959
rect 13279 45913 13357 45959
rect 13403 45913 13481 45959
rect 13527 45913 13605 45959
rect 13651 45913 13729 45959
rect 13775 45913 13853 45959
rect 13899 45913 13977 45959
rect 14023 45913 14101 45959
rect 14147 45913 14225 45959
rect 14271 45913 14349 45959
rect 14395 45913 14473 45959
rect 14519 45913 14597 45959
rect 14643 45913 14721 45959
rect 14767 45913 14845 45959
rect 14891 45913 14969 45959
rect 15015 45913 15093 45959
rect 15139 45913 15217 45959
rect 15263 45913 15341 45959
rect 15387 45913 15465 45959
rect 15511 45913 15589 45959
rect 15635 45913 15713 45959
rect 15759 45913 15837 45959
rect 15883 45913 15961 45959
rect 16007 45913 16085 45959
rect 16131 45913 16209 45959
rect 16255 45913 16333 45959
rect 16379 45913 16457 45959
rect 16503 45913 16581 45959
rect 16627 45913 16705 45959
rect 16751 45913 16829 45959
rect 16875 45913 16953 45959
rect 16999 45913 17077 45959
rect 17123 45913 17201 45959
rect 17247 45913 17325 45959
rect 17371 45913 17449 45959
rect 17495 45913 17573 45959
rect 17619 45913 17697 45959
rect 17743 45913 17821 45959
rect 17867 45913 17945 45959
rect 17991 45913 18069 45959
rect 18115 45913 18193 45959
rect 18239 45913 18317 45959
rect 18363 45913 18441 45959
rect 18487 45913 18565 45959
rect 18611 45913 18689 45959
rect 18735 45913 18813 45959
rect 18859 45913 18937 45959
rect 18983 45913 19061 45959
rect 19107 45913 19185 45959
rect 19231 45913 19309 45959
rect 19355 45913 19433 45959
rect 19479 45913 19557 45959
rect 19603 45913 19681 45959
rect 19727 45913 19805 45959
rect 19851 45913 19929 45959
rect 19975 45913 20053 45959
rect 20099 45913 20177 45959
rect 20223 45913 20301 45959
rect 20347 45913 20425 45959
rect 20471 45913 20549 45959
rect 20595 45913 20673 45959
rect 20719 45913 20797 45959
rect 20843 45913 20921 45959
rect 20967 45913 21045 45959
rect 21091 45913 21169 45959
rect 21215 45913 21293 45959
rect 21339 45913 21417 45959
rect 21463 45913 21541 45959
rect 21587 45913 21665 45959
rect 21711 45913 21789 45959
rect 21835 45913 21913 45959
rect 21959 45913 22037 45959
rect 22083 45913 22161 45959
rect 22207 45913 22285 45959
rect 22331 45913 22409 45959
rect 22455 45913 22533 45959
rect 22579 45913 22657 45959
rect 22703 45913 22781 45959
rect 22827 45913 22905 45959
rect 22951 45913 23029 45959
rect 23075 45913 23153 45959
rect 23199 45913 23277 45959
rect 23323 45913 23401 45959
rect 23447 45913 23525 45959
rect 23571 45913 23649 45959
rect 23695 45913 23773 45959
rect 23819 45913 23897 45959
rect 23943 45913 24021 45959
rect 24067 45913 24145 45959
rect 24191 45913 24269 45959
rect 24315 45913 24393 45959
rect 24439 45913 24517 45959
rect 24563 45913 24641 45959
rect 24687 45913 24765 45959
rect 24811 45913 24889 45959
rect 24935 45913 25013 45959
rect 25059 45913 25137 45959
rect 25183 45913 25261 45959
rect 25307 45913 25385 45959
rect 25431 45913 25509 45959
rect 25555 45913 25633 45959
rect 25679 45913 25757 45959
rect 25803 45913 25881 45959
rect 25927 45913 26005 45959
rect 26051 45913 26129 45959
rect 26175 45913 26253 45959
rect 26299 45913 26377 45959
rect 26423 45913 26501 45959
rect 26547 45913 26625 45959
rect 26671 45913 26749 45959
rect 26795 45913 26873 45959
rect 26919 45913 26997 45959
rect 27043 45913 27121 45959
rect 27167 45913 27245 45959
rect 27291 45913 27369 45959
rect 27415 45913 27493 45959
rect 27539 45913 27617 45959
rect 27663 45913 27741 45959
rect 27787 45913 27865 45959
rect 27911 45913 27989 45959
rect 28035 45913 28113 45959
rect 28159 45913 28237 45959
rect 28283 45913 28361 45959
rect 28407 45913 28485 45959
rect 28531 45913 28609 45959
rect 28655 45913 28733 45959
rect 28779 45913 28857 45959
rect 28903 45913 28981 45959
rect 29027 45913 29105 45959
rect 29151 45913 29229 45959
rect 29275 45913 29353 45959
rect 29399 45913 29477 45959
rect 29523 45913 29601 45959
rect 29647 45913 29725 45959
rect 29771 45913 29849 45959
rect 29895 45913 29973 45959
rect 30019 45913 30097 45959
rect 30143 45913 30221 45959
rect 30267 45913 30345 45959
rect 30391 45913 30469 45959
rect 30515 45913 30593 45959
rect 30639 45913 30717 45959
rect 30763 45913 30841 45959
rect 30887 45913 30965 45959
rect 31011 45913 31089 45959
rect 31135 45913 31213 45959
rect 31259 45913 31337 45959
rect 31383 45913 31461 45959
rect 31507 45913 31585 45959
rect 31631 45913 31709 45959
rect 31755 45913 31833 45959
rect 31879 45913 31957 45959
rect 32003 45913 32081 45959
rect 32127 45913 32205 45959
rect 32251 45913 32329 45959
rect 32375 45913 32453 45959
rect 32499 45913 32577 45959
rect 32623 45913 32701 45959
rect 32747 45913 32825 45959
rect 32871 45913 32949 45959
rect 32995 45913 33073 45959
rect 33119 45913 33197 45959
rect 33243 45913 33321 45959
rect 33367 45913 33445 45959
rect 33491 45913 33569 45959
rect 33615 45913 33693 45959
rect 33739 45913 33817 45959
rect 33863 45913 33941 45959
rect 33987 45913 34065 45959
rect 34111 45913 34189 45959
rect 34235 45913 34313 45959
rect 34359 45913 34437 45959
rect 34483 45913 34561 45959
rect 34607 45913 34685 45959
rect 34731 45913 34809 45959
rect 34855 45913 34933 45959
rect 34979 45913 35057 45959
rect 35103 45913 35181 45959
rect 35227 45913 35305 45959
rect 35351 45913 35429 45959
rect 35475 45913 35553 45959
rect 35599 45913 35677 45959
rect 35723 45913 35801 45959
rect 35847 45913 35925 45959
rect 35971 45913 36049 45959
rect 36095 45913 36173 45959
rect 36219 45913 36297 45959
rect 36343 45913 36421 45959
rect 36467 45913 36545 45959
rect 36591 45913 36669 45959
rect 36715 45913 36793 45959
rect 36839 45913 36917 45959
rect 36963 45913 37041 45959
rect 37087 45913 37165 45959
rect 37211 45913 37289 45959
rect 37335 45913 37413 45959
rect 37459 45913 37537 45959
rect 37583 45913 37661 45959
rect 37707 45913 37785 45959
rect 37831 45913 37909 45959
rect 37955 45913 38033 45959
rect 38079 45913 38157 45959
rect 38203 45913 38281 45959
rect 38327 45913 38405 45959
rect 38451 45913 38529 45959
rect 38575 45913 38653 45959
rect 38699 45913 38777 45959
rect 38823 45913 38901 45959
rect 38947 45913 39025 45959
rect 39071 45913 39149 45959
rect 39195 45913 39273 45959
rect 39319 45913 39397 45959
rect 39443 45913 39521 45959
rect 39567 45913 39645 45959
rect 39691 45913 39769 45959
rect 39815 45913 39893 45959
rect 39939 45913 40017 45959
rect 40063 45913 40141 45959
rect 40187 45913 40265 45959
rect 40311 45913 40389 45959
rect 40435 45913 40513 45959
rect 40559 45913 40637 45959
rect 40683 45913 40761 45959
rect 40807 45913 40885 45959
rect 40931 45913 41009 45959
rect 41055 45913 41133 45959
rect 41179 45913 41257 45959
rect 41303 45913 41381 45959
rect 41427 45913 41505 45959
rect 41551 45913 41629 45959
rect 41675 45913 41753 45959
rect 41799 45913 41877 45959
rect 41923 45913 42001 45959
rect 42047 45913 42125 45959
rect 42171 45913 42249 45959
rect 42295 45913 42373 45959
rect 42419 45913 42497 45959
rect 42543 45913 42621 45959
rect 42667 45913 42745 45959
rect 42791 45913 42869 45959
rect 42915 45913 42993 45959
rect 43039 45913 43117 45959
rect 43163 45913 43241 45959
rect 43287 45913 43365 45959
rect 43411 45913 43489 45959
rect 43535 45913 43613 45959
rect 43659 45913 43737 45959
rect 43783 45913 43861 45959
rect 43907 45913 43985 45959
rect 44031 45913 44109 45959
rect 44155 45913 44233 45959
rect 44279 45913 44357 45959
rect 44403 45913 44481 45959
rect 44527 45913 44605 45959
rect 44651 45913 44729 45959
rect 44775 45913 44853 45959
rect 44899 45913 44977 45959
rect 45023 45913 45101 45959
rect 45147 45913 45225 45959
rect 45271 45913 45349 45959
rect 45395 45913 45473 45959
rect 45519 45913 45597 45959
rect 45643 45913 45721 45959
rect 45767 45913 45845 45959
rect 45891 45913 45969 45959
rect 46015 45913 46093 45959
rect 46139 45913 46217 45959
rect 46263 45913 46341 45959
rect 46387 45913 46465 45959
rect 46511 45913 46589 45959
rect 46635 45913 46713 45959
rect 46759 45913 46837 45959
rect 46883 45913 46961 45959
rect 47007 45913 47085 45959
rect 47131 45913 47209 45959
rect 47255 45913 47333 45959
rect 47379 45913 47457 45959
rect 47503 45913 47581 45959
rect 47627 45913 47705 45959
rect 47751 45913 47829 45959
rect 47875 45913 47953 45959
rect 47999 45913 48077 45959
rect 48123 45913 48201 45959
rect 48247 45913 48325 45959
rect 48371 45913 48449 45959
rect 48495 45913 48573 45959
rect 48619 45913 48697 45959
rect 48743 45913 48821 45959
rect 48867 45913 48945 45959
rect 48991 45913 49069 45959
rect 49115 45913 49193 45959
rect 49239 45913 49317 45959
rect 49363 45913 49441 45959
rect 49487 45913 49565 45959
rect 49611 45913 49689 45959
rect 49735 45913 49813 45959
rect 49859 45913 49937 45959
rect 49983 45913 50061 45959
rect 50107 45913 50185 45959
rect 50231 45913 50309 45959
rect 50355 45913 50433 45959
rect 50479 45913 50557 45959
rect 50603 45913 50681 45959
rect 50727 45913 50805 45959
rect 50851 45913 50929 45959
rect 50975 45913 51053 45959
rect 51099 45913 51177 45959
rect 51223 45913 51301 45959
rect 51347 45913 51425 45959
rect 51471 45913 51549 45959
rect 51595 45913 51673 45959
rect 51719 45913 51797 45959
rect 51843 45913 51921 45959
rect 51967 45913 52045 45959
rect 52091 45913 52169 45959
rect 52215 45913 52293 45959
rect 52339 45913 52417 45959
rect 52463 45913 52541 45959
rect 52587 45913 52665 45959
rect 52711 45913 52789 45959
rect 52835 45913 52913 45959
rect 52959 45913 53037 45959
rect 53083 45913 53161 45959
rect 53207 45913 53285 45959
rect 53331 45913 53409 45959
rect 53455 45913 53533 45959
rect 53579 45913 53657 45959
rect 53703 45913 53781 45959
rect 53827 45913 53905 45959
rect 53951 45913 54029 45959
rect 54075 45913 54153 45959
rect 54199 45913 54277 45959
rect 54323 45913 54401 45959
rect 54447 45913 54525 45959
rect 54571 45913 54649 45959
rect 54695 45913 54773 45959
rect 54819 45913 54897 45959
rect 54943 45913 55021 45959
rect 55067 45913 55145 45959
rect 55191 45913 55269 45959
rect 55315 45913 55393 45959
rect 55439 45913 55517 45959
rect 55563 45913 55641 45959
rect 55687 45913 55765 45959
rect 55811 45913 55889 45959
rect 55935 45913 56013 45959
rect 56059 45913 56137 45959
rect 56183 45913 56261 45959
rect 56307 45913 56385 45959
rect 56431 45913 56509 45959
rect 56555 45913 56633 45959
rect 56679 45913 56757 45959
rect 56803 45913 56881 45959
rect 56927 45913 57005 45959
rect 57051 45913 57129 45959
rect 57175 45913 57253 45959
rect 57299 45913 57377 45959
rect 57423 45913 57501 45959
rect 57547 45913 57625 45959
rect 57671 45913 57749 45959
rect 57795 45913 57873 45959
rect 57919 45913 57997 45959
rect 58043 45913 58121 45959
rect 58167 45913 58245 45959
rect 58291 45913 58369 45959
rect 58415 45913 58493 45959
rect 58539 45913 58617 45959
rect 58663 45913 58741 45959
rect 58787 45913 58865 45959
rect 58911 45913 58989 45959
rect 59035 45913 59113 45959
rect 59159 45913 59237 45959
rect 59283 45913 59361 45959
rect 59407 45913 59485 45959
rect 59531 45913 59609 45959
rect 59655 45913 59733 45959
rect 59779 45913 59857 45959
rect 59903 45913 59981 45959
rect 60027 45913 60105 45959
rect 60151 45913 60229 45959
rect 60275 45913 60353 45959
rect 60399 45913 60477 45959
rect 60523 45913 60601 45959
rect 60647 45913 60725 45959
rect 60771 45913 60849 45959
rect 60895 45913 60973 45959
rect 61019 45913 61097 45959
rect 61143 45913 61221 45959
rect 61267 45913 61345 45959
rect 61391 45913 61469 45959
rect 61515 45913 61593 45959
rect 61639 45913 61717 45959
rect 61763 45913 61841 45959
rect 61887 45913 61965 45959
rect 62011 45913 62089 45959
rect 62135 45913 62213 45959
rect 62259 45913 62337 45959
rect 62383 45913 62461 45959
rect 62507 45913 62585 45959
rect 62631 45913 62709 45959
rect 62755 45913 62833 45959
rect 62879 45913 62957 45959
rect 63003 45913 63081 45959
rect 63127 45913 63205 45959
rect 63251 45913 63329 45959
rect 63375 45913 63453 45959
rect 63499 45913 63577 45959
rect 63623 45913 63701 45959
rect 63747 45913 63825 45959
rect 63871 45913 63949 45959
rect 63995 45913 64073 45959
rect 64119 45913 64197 45959
rect 64243 45913 64321 45959
rect 64367 45913 64445 45959
rect 64491 45913 64569 45959
rect 64615 45913 64693 45959
rect 64739 45913 64817 45959
rect 64863 45913 64941 45959
rect 64987 45913 65065 45959
rect 65111 45913 65189 45959
rect 65235 45913 65313 45959
rect 65359 45913 65437 45959
rect 65483 45913 65561 45959
rect 65607 45913 65685 45959
rect 65731 45913 65809 45959
rect 65855 45913 65933 45959
rect 65979 45913 66057 45959
rect 66103 45913 66181 45959
rect 66227 45913 66305 45959
rect 66351 45913 66429 45959
rect 66475 45913 66553 45959
rect 66599 45913 66677 45959
rect 66723 45913 66801 45959
rect 66847 45913 66925 45959
rect 66971 45913 67049 45959
rect 67095 45913 67173 45959
rect 67219 45913 67297 45959
rect 67343 45913 67421 45959
rect 67467 45913 67545 45959
rect 67591 45913 67669 45959
rect 67715 45913 67793 45959
rect 67839 45913 67917 45959
rect 67963 45913 68041 45959
rect 68087 45913 68165 45959
rect 68211 45913 68289 45959
rect 68335 45913 68413 45959
rect 68459 45913 68537 45959
rect 68583 45913 68661 45959
rect 68707 45913 68785 45959
rect 68831 45913 68909 45959
rect 68955 45913 69033 45959
rect 69079 45913 69157 45959
rect 69203 45913 69281 45959
rect 69327 45913 69405 45959
rect 69451 45913 69529 45959
rect 69575 45913 69653 45959
rect 69699 45913 69777 45959
rect 69823 45913 69901 45959
rect 69947 45913 70025 45959
rect 70071 45913 70149 45959
rect 70195 45913 70273 45959
rect 70319 45913 70397 45959
rect 70443 45913 70521 45959
rect 70567 45913 70645 45959
rect 70691 45913 70769 45959
rect 70815 45913 70893 45959
rect 70939 45913 71017 45959
rect 71063 45913 71141 45959
rect 71187 45913 71265 45959
rect 71311 45913 71389 45959
rect 71435 45913 71513 45959
rect 71559 45913 71637 45959
rect 71683 45913 71761 45959
rect 71807 45913 71885 45959
rect 71931 45913 72009 45959
rect 72055 45913 72133 45959
rect 72179 45913 72257 45959
rect 72303 45913 72381 45959
rect 72427 45913 72505 45959
rect 72551 45913 72629 45959
rect 72675 45913 72753 45959
rect 72799 45913 72877 45959
rect 72923 45913 73001 45959
rect 73047 45913 73125 45959
rect 73171 45913 73249 45959
rect 73295 45913 73373 45959
rect 73419 45913 73497 45959
rect 73543 45913 73621 45959
rect 73667 45913 73745 45959
rect 73791 45913 73869 45959
rect 73915 45913 73993 45959
rect 74039 45913 74117 45959
rect 74163 45913 74241 45959
rect 74287 45913 74365 45959
rect 74411 45913 74489 45959
rect 74535 45913 74613 45959
rect 74659 45913 74737 45959
rect 74783 45913 74861 45959
rect 74907 45913 74985 45959
rect 75031 45913 75109 45959
rect 75155 45913 75233 45959
rect 75279 45913 75357 45959
rect 75403 45913 75481 45959
rect 75527 45913 75605 45959
rect 75651 45913 75729 45959
rect 75775 45913 75853 45959
rect 75899 45913 75977 45959
rect 76023 45913 76101 45959
rect 76147 45913 76225 45959
rect 76271 45913 76349 45959
rect 76395 45913 76473 45959
rect 76519 45913 76597 45959
rect 76643 45913 76721 45959
rect 76767 45913 76845 45959
rect 76891 45913 76969 45959
rect 77015 45913 77093 45959
rect 77139 45913 77217 45959
rect 77263 45913 77341 45959
rect 77387 45913 77465 45959
rect 77511 45913 77589 45959
rect 77635 45913 77713 45959
rect 77759 45913 77837 45959
rect 77883 45913 77961 45959
rect 78007 45913 78085 45959
rect 78131 45913 78209 45959
rect 78255 45913 78333 45959
rect 78379 45913 78457 45959
rect 78503 45913 78581 45959
rect 78627 45913 78705 45959
rect 78751 45913 78829 45959
rect 78875 45913 78953 45959
rect 78999 45913 79077 45959
rect 79123 45913 79201 45959
rect 79247 45913 79325 45959
rect 79371 45913 79449 45959
rect 79495 45913 79573 45959
rect 79619 45913 79697 45959
rect 79743 45913 79821 45959
rect 79867 45913 79945 45959
rect 79991 45913 80069 45959
rect 80115 45913 80193 45959
rect 80239 45913 80317 45959
rect 80363 45913 80441 45959
rect 80487 45913 80565 45959
rect 80611 45913 80689 45959
rect 80735 45913 80813 45959
rect 80859 45913 80937 45959
rect 80983 45913 81061 45959
rect 81107 45913 81185 45959
rect 81231 45913 81309 45959
rect 81355 45913 81433 45959
rect 81479 45913 81557 45959
rect 81603 45913 81681 45959
rect 81727 45913 81805 45959
rect 81851 45913 81929 45959
rect 81975 45913 82053 45959
rect 82099 45913 82177 45959
rect 82223 45913 82301 45959
rect 82347 45913 82425 45959
rect 82471 45913 82549 45959
rect 82595 45913 82673 45959
rect 82719 45913 82797 45959
rect 82843 45913 82921 45959
rect 82967 45913 83045 45959
rect 83091 45913 83169 45959
rect 83215 45913 83293 45959
rect 83339 45913 83417 45959
rect 83463 45913 83541 45959
rect 83587 45913 83665 45959
rect 83711 45913 83789 45959
rect 83835 45913 83913 45959
rect 83959 45913 84037 45959
rect 84083 45913 84161 45959
rect 84207 45913 84285 45959
rect 84331 45913 84409 45959
rect 84455 45913 84533 45959
rect 84579 45913 84657 45959
rect 84703 45913 84781 45959
rect 84827 45913 84905 45959
rect 84951 45913 85029 45959
rect 85075 45913 85153 45959
rect 85199 45913 85277 45959
rect 85323 45913 85401 45959
rect 85447 45913 85525 45959
rect 85571 45913 85649 45959
rect 85695 45913 85816 45959
rect 70 45835 85816 45913
rect 70 45789 89 45835
rect 135 45789 213 45835
rect 259 45789 337 45835
rect 383 45789 461 45835
rect 507 45789 585 45835
rect 631 45789 709 45835
rect 755 45789 833 45835
rect 879 45789 957 45835
rect 1003 45789 1081 45835
rect 1127 45789 1205 45835
rect 1251 45789 1329 45835
rect 1375 45789 1453 45835
rect 1499 45789 1577 45835
rect 1623 45789 1701 45835
rect 1747 45789 1825 45835
rect 1871 45789 1949 45835
rect 1995 45789 2073 45835
rect 2119 45789 2197 45835
rect 2243 45789 2321 45835
rect 2367 45789 2445 45835
rect 2491 45789 2569 45835
rect 2615 45789 2693 45835
rect 2739 45789 2817 45835
rect 2863 45789 2941 45835
rect 2987 45789 3065 45835
rect 3111 45789 3189 45835
rect 3235 45789 3313 45835
rect 3359 45789 3437 45835
rect 3483 45789 3561 45835
rect 3607 45789 3685 45835
rect 3731 45789 3809 45835
rect 3855 45789 3933 45835
rect 3979 45789 4057 45835
rect 4103 45789 4181 45835
rect 4227 45789 4305 45835
rect 4351 45789 4429 45835
rect 4475 45789 4553 45835
rect 4599 45789 4677 45835
rect 4723 45789 4801 45835
rect 4847 45789 4925 45835
rect 4971 45789 5049 45835
rect 5095 45789 5173 45835
rect 5219 45789 5297 45835
rect 5343 45789 5421 45835
rect 5467 45789 5545 45835
rect 5591 45789 5669 45835
rect 5715 45789 5793 45835
rect 5839 45789 5917 45835
rect 5963 45789 6041 45835
rect 6087 45789 6165 45835
rect 6211 45789 6289 45835
rect 6335 45789 6413 45835
rect 6459 45789 6537 45835
rect 6583 45789 6661 45835
rect 6707 45789 6785 45835
rect 6831 45789 6909 45835
rect 6955 45789 7033 45835
rect 7079 45789 7157 45835
rect 7203 45789 7281 45835
rect 7327 45789 7405 45835
rect 7451 45789 7529 45835
rect 7575 45789 7653 45835
rect 7699 45789 7777 45835
rect 7823 45789 7901 45835
rect 7947 45789 8025 45835
rect 8071 45789 8149 45835
rect 8195 45789 8273 45835
rect 8319 45789 8397 45835
rect 8443 45789 8521 45835
rect 8567 45789 8645 45835
rect 8691 45789 8769 45835
rect 8815 45789 8893 45835
rect 8939 45789 9017 45835
rect 9063 45789 9141 45835
rect 9187 45789 9265 45835
rect 9311 45789 9389 45835
rect 9435 45789 9513 45835
rect 9559 45789 9637 45835
rect 9683 45789 9761 45835
rect 9807 45789 9885 45835
rect 9931 45789 10009 45835
rect 10055 45789 10133 45835
rect 10179 45789 10257 45835
rect 10303 45789 10381 45835
rect 10427 45789 10505 45835
rect 10551 45789 10629 45835
rect 10675 45789 10753 45835
rect 10799 45789 10877 45835
rect 10923 45789 11001 45835
rect 11047 45789 11125 45835
rect 11171 45789 11249 45835
rect 11295 45789 11373 45835
rect 11419 45789 11497 45835
rect 11543 45789 11621 45835
rect 11667 45789 11745 45835
rect 11791 45789 11869 45835
rect 11915 45789 11993 45835
rect 12039 45789 12117 45835
rect 12163 45789 12241 45835
rect 12287 45789 12365 45835
rect 12411 45789 12489 45835
rect 12535 45789 12613 45835
rect 12659 45789 12737 45835
rect 12783 45789 12861 45835
rect 12907 45789 12985 45835
rect 13031 45789 13109 45835
rect 13155 45789 13233 45835
rect 13279 45789 13357 45835
rect 13403 45789 13481 45835
rect 13527 45789 13605 45835
rect 13651 45789 13729 45835
rect 13775 45789 13853 45835
rect 13899 45789 13977 45835
rect 14023 45789 14101 45835
rect 14147 45789 14225 45835
rect 14271 45789 14349 45835
rect 14395 45789 14473 45835
rect 14519 45789 14597 45835
rect 14643 45789 14721 45835
rect 14767 45789 14845 45835
rect 14891 45789 14969 45835
rect 15015 45789 15093 45835
rect 15139 45789 15217 45835
rect 15263 45789 15341 45835
rect 15387 45789 15465 45835
rect 15511 45789 15589 45835
rect 15635 45789 15713 45835
rect 15759 45789 15837 45835
rect 15883 45789 15961 45835
rect 16007 45789 16085 45835
rect 16131 45789 16209 45835
rect 16255 45789 16333 45835
rect 16379 45789 16457 45835
rect 16503 45789 16581 45835
rect 16627 45789 16705 45835
rect 16751 45789 16829 45835
rect 16875 45789 16953 45835
rect 16999 45789 17077 45835
rect 17123 45789 17201 45835
rect 17247 45789 17325 45835
rect 17371 45789 17449 45835
rect 17495 45789 17573 45835
rect 17619 45789 17697 45835
rect 17743 45789 17821 45835
rect 17867 45789 17945 45835
rect 17991 45789 18069 45835
rect 18115 45789 18193 45835
rect 18239 45789 18317 45835
rect 18363 45789 18441 45835
rect 18487 45789 18565 45835
rect 18611 45789 18689 45835
rect 18735 45789 18813 45835
rect 18859 45789 18937 45835
rect 18983 45789 19061 45835
rect 19107 45789 19185 45835
rect 19231 45789 19309 45835
rect 19355 45789 19433 45835
rect 19479 45789 19557 45835
rect 19603 45789 19681 45835
rect 19727 45789 19805 45835
rect 19851 45789 19929 45835
rect 19975 45789 20053 45835
rect 20099 45789 20177 45835
rect 20223 45789 20301 45835
rect 20347 45789 20425 45835
rect 20471 45789 20549 45835
rect 20595 45789 20673 45835
rect 20719 45789 20797 45835
rect 20843 45789 20921 45835
rect 20967 45789 21045 45835
rect 21091 45789 21169 45835
rect 21215 45789 21293 45835
rect 21339 45789 21417 45835
rect 21463 45789 21541 45835
rect 21587 45789 21665 45835
rect 21711 45789 21789 45835
rect 21835 45789 21913 45835
rect 21959 45789 22037 45835
rect 22083 45789 22161 45835
rect 22207 45789 22285 45835
rect 22331 45789 22409 45835
rect 22455 45789 22533 45835
rect 22579 45789 22657 45835
rect 22703 45789 22781 45835
rect 22827 45789 22905 45835
rect 22951 45789 23029 45835
rect 23075 45789 23153 45835
rect 23199 45789 23277 45835
rect 23323 45789 23401 45835
rect 23447 45789 23525 45835
rect 23571 45789 23649 45835
rect 23695 45789 23773 45835
rect 23819 45789 23897 45835
rect 23943 45789 24021 45835
rect 24067 45789 24145 45835
rect 24191 45789 24269 45835
rect 24315 45789 24393 45835
rect 24439 45789 24517 45835
rect 24563 45789 24641 45835
rect 24687 45789 24765 45835
rect 24811 45789 24889 45835
rect 24935 45789 25013 45835
rect 25059 45789 25137 45835
rect 25183 45789 25261 45835
rect 25307 45789 25385 45835
rect 25431 45789 25509 45835
rect 25555 45789 25633 45835
rect 25679 45789 25757 45835
rect 25803 45789 25881 45835
rect 25927 45789 26005 45835
rect 26051 45789 26129 45835
rect 26175 45789 26253 45835
rect 26299 45789 26377 45835
rect 26423 45789 26501 45835
rect 26547 45789 26625 45835
rect 26671 45789 26749 45835
rect 26795 45789 26873 45835
rect 26919 45789 26997 45835
rect 27043 45789 27121 45835
rect 27167 45789 27245 45835
rect 27291 45789 27369 45835
rect 27415 45789 27493 45835
rect 27539 45789 27617 45835
rect 27663 45789 27741 45835
rect 27787 45789 27865 45835
rect 27911 45789 27989 45835
rect 28035 45789 28113 45835
rect 28159 45789 28237 45835
rect 28283 45789 28361 45835
rect 28407 45789 28485 45835
rect 28531 45789 28609 45835
rect 28655 45789 28733 45835
rect 28779 45789 28857 45835
rect 28903 45789 28981 45835
rect 29027 45789 29105 45835
rect 29151 45789 29229 45835
rect 29275 45789 29353 45835
rect 29399 45789 29477 45835
rect 29523 45789 29601 45835
rect 29647 45789 29725 45835
rect 29771 45789 29849 45835
rect 29895 45789 29973 45835
rect 30019 45789 30097 45835
rect 30143 45789 30221 45835
rect 30267 45789 30345 45835
rect 30391 45789 30469 45835
rect 30515 45789 30593 45835
rect 30639 45789 30717 45835
rect 30763 45789 30841 45835
rect 30887 45789 30965 45835
rect 31011 45789 31089 45835
rect 31135 45789 31213 45835
rect 31259 45789 31337 45835
rect 31383 45789 31461 45835
rect 31507 45789 31585 45835
rect 31631 45789 31709 45835
rect 31755 45789 31833 45835
rect 31879 45789 31957 45835
rect 32003 45789 32081 45835
rect 32127 45789 32205 45835
rect 32251 45789 32329 45835
rect 32375 45789 32453 45835
rect 32499 45789 32577 45835
rect 32623 45789 32701 45835
rect 32747 45789 32825 45835
rect 32871 45789 32949 45835
rect 32995 45789 33073 45835
rect 33119 45789 33197 45835
rect 33243 45789 33321 45835
rect 33367 45789 33445 45835
rect 33491 45789 33569 45835
rect 33615 45789 33693 45835
rect 33739 45789 33817 45835
rect 33863 45789 33941 45835
rect 33987 45789 34065 45835
rect 34111 45789 34189 45835
rect 34235 45789 34313 45835
rect 34359 45789 34437 45835
rect 34483 45789 34561 45835
rect 34607 45789 34685 45835
rect 34731 45789 34809 45835
rect 34855 45789 34933 45835
rect 34979 45789 35057 45835
rect 35103 45789 35181 45835
rect 35227 45789 35305 45835
rect 35351 45789 35429 45835
rect 35475 45789 35553 45835
rect 35599 45789 35677 45835
rect 35723 45789 35801 45835
rect 35847 45789 35925 45835
rect 35971 45789 36049 45835
rect 36095 45789 36173 45835
rect 36219 45789 36297 45835
rect 36343 45789 36421 45835
rect 36467 45789 36545 45835
rect 36591 45789 36669 45835
rect 36715 45789 36793 45835
rect 36839 45789 36917 45835
rect 36963 45789 37041 45835
rect 37087 45789 37165 45835
rect 37211 45789 37289 45835
rect 37335 45789 37413 45835
rect 37459 45789 37537 45835
rect 37583 45789 37661 45835
rect 37707 45789 37785 45835
rect 37831 45789 37909 45835
rect 37955 45789 38033 45835
rect 38079 45789 38157 45835
rect 38203 45789 38281 45835
rect 38327 45789 38405 45835
rect 38451 45789 38529 45835
rect 38575 45789 38653 45835
rect 38699 45789 38777 45835
rect 38823 45789 38901 45835
rect 38947 45789 39025 45835
rect 39071 45789 39149 45835
rect 39195 45789 39273 45835
rect 39319 45789 39397 45835
rect 39443 45789 39521 45835
rect 39567 45789 39645 45835
rect 39691 45789 39769 45835
rect 39815 45789 39893 45835
rect 39939 45789 40017 45835
rect 40063 45789 40141 45835
rect 40187 45789 40265 45835
rect 40311 45789 40389 45835
rect 40435 45789 40513 45835
rect 40559 45789 40637 45835
rect 40683 45789 40761 45835
rect 40807 45789 40885 45835
rect 40931 45789 41009 45835
rect 41055 45789 41133 45835
rect 41179 45789 41257 45835
rect 41303 45789 41381 45835
rect 41427 45789 41505 45835
rect 41551 45789 41629 45835
rect 41675 45789 41753 45835
rect 41799 45789 41877 45835
rect 41923 45789 42001 45835
rect 42047 45789 42125 45835
rect 42171 45789 42249 45835
rect 42295 45789 42373 45835
rect 42419 45789 42497 45835
rect 42543 45789 42621 45835
rect 42667 45789 42745 45835
rect 42791 45789 42869 45835
rect 42915 45789 42993 45835
rect 43039 45789 43117 45835
rect 43163 45789 43241 45835
rect 43287 45789 43365 45835
rect 43411 45789 43489 45835
rect 43535 45789 43613 45835
rect 43659 45789 43737 45835
rect 43783 45789 43861 45835
rect 43907 45789 43985 45835
rect 44031 45789 44109 45835
rect 44155 45789 44233 45835
rect 44279 45789 44357 45835
rect 44403 45789 44481 45835
rect 44527 45789 44605 45835
rect 44651 45789 44729 45835
rect 44775 45789 44853 45835
rect 44899 45789 44977 45835
rect 45023 45789 45101 45835
rect 45147 45789 45225 45835
rect 45271 45789 45349 45835
rect 45395 45789 45473 45835
rect 45519 45789 45597 45835
rect 45643 45789 45721 45835
rect 45767 45789 45845 45835
rect 45891 45789 45969 45835
rect 46015 45789 46093 45835
rect 46139 45789 46217 45835
rect 46263 45789 46341 45835
rect 46387 45789 46465 45835
rect 46511 45789 46589 45835
rect 46635 45789 46713 45835
rect 46759 45789 46837 45835
rect 46883 45789 46961 45835
rect 47007 45789 47085 45835
rect 47131 45789 47209 45835
rect 47255 45789 47333 45835
rect 47379 45789 47457 45835
rect 47503 45789 47581 45835
rect 47627 45789 47705 45835
rect 47751 45789 47829 45835
rect 47875 45789 47953 45835
rect 47999 45789 48077 45835
rect 48123 45789 48201 45835
rect 48247 45789 48325 45835
rect 48371 45789 48449 45835
rect 48495 45789 48573 45835
rect 48619 45789 48697 45835
rect 48743 45789 48821 45835
rect 48867 45789 48945 45835
rect 48991 45789 49069 45835
rect 49115 45789 49193 45835
rect 49239 45789 49317 45835
rect 49363 45789 49441 45835
rect 49487 45789 49565 45835
rect 49611 45789 49689 45835
rect 49735 45789 49813 45835
rect 49859 45789 49937 45835
rect 49983 45789 50061 45835
rect 50107 45789 50185 45835
rect 50231 45789 50309 45835
rect 50355 45789 50433 45835
rect 50479 45789 50557 45835
rect 50603 45789 50681 45835
rect 50727 45789 50805 45835
rect 50851 45789 50929 45835
rect 50975 45789 51053 45835
rect 51099 45789 51177 45835
rect 51223 45789 51301 45835
rect 51347 45789 51425 45835
rect 51471 45789 51549 45835
rect 51595 45789 51673 45835
rect 51719 45789 51797 45835
rect 51843 45789 51921 45835
rect 51967 45789 52045 45835
rect 52091 45789 52169 45835
rect 52215 45789 52293 45835
rect 52339 45789 52417 45835
rect 52463 45789 52541 45835
rect 52587 45789 52665 45835
rect 52711 45789 52789 45835
rect 52835 45789 52913 45835
rect 52959 45789 53037 45835
rect 53083 45789 53161 45835
rect 53207 45789 53285 45835
rect 53331 45789 53409 45835
rect 53455 45789 53533 45835
rect 53579 45789 53657 45835
rect 53703 45789 53781 45835
rect 53827 45789 53905 45835
rect 53951 45789 54029 45835
rect 54075 45789 54153 45835
rect 54199 45789 54277 45835
rect 54323 45789 54401 45835
rect 54447 45789 54525 45835
rect 54571 45789 54649 45835
rect 54695 45789 54773 45835
rect 54819 45789 54897 45835
rect 54943 45789 55021 45835
rect 55067 45789 55145 45835
rect 55191 45789 55269 45835
rect 55315 45789 55393 45835
rect 55439 45789 55517 45835
rect 55563 45789 55641 45835
rect 55687 45789 55765 45835
rect 55811 45789 55889 45835
rect 55935 45789 56013 45835
rect 56059 45789 56137 45835
rect 56183 45789 56261 45835
rect 56307 45789 56385 45835
rect 56431 45789 56509 45835
rect 56555 45789 56633 45835
rect 56679 45789 56757 45835
rect 56803 45789 56881 45835
rect 56927 45789 57005 45835
rect 57051 45789 57129 45835
rect 57175 45789 57253 45835
rect 57299 45789 57377 45835
rect 57423 45789 57501 45835
rect 57547 45789 57625 45835
rect 57671 45789 57749 45835
rect 57795 45789 57873 45835
rect 57919 45789 57997 45835
rect 58043 45789 58121 45835
rect 58167 45789 58245 45835
rect 58291 45789 58369 45835
rect 58415 45789 58493 45835
rect 58539 45789 58617 45835
rect 58663 45789 58741 45835
rect 58787 45789 58865 45835
rect 58911 45789 58989 45835
rect 59035 45789 59113 45835
rect 59159 45789 59237 45835
rect 59283 45789 59361 45835
rect 59407 45789 59485 45835
rect 59531 45789 59609 45835
rect 59655 45789 59733 45835
rect 59779 45789 59857 45835
rect 59903 45789 59981 45835
rect 60027 45789 60105 45835
rect 60151 45789 60229 45835
rect 60275 45789 60353 45835
rect 60399 45789 60477 45835
rect 60523 45789 60601 45835
rect 60647 45789 60725 45835
rect 60771 45789 60849 45835
rect 60895 45789 60973 45835
rect 61019 45789 61097 45835
rect 61143 45789 61221 45835
rect 61267 45789 61345 45835
rect 61391 45789 61469 45835
rect 61515 45789 61593 45835
rect 61639 45789 61717 45835
rect 61763 45789 61841 45835
rect 61887 45789 61965 45835
rect 62011 45789 62089 45835
rect 62135 45789 62213 45835
rect 62259 45789 62337 45835
rect 62383 45789 62461 45835
rect 62507 45789 62585 45835
rect 62631 45789 62709 45835
rect 62755 45789 62833 45835
rect 62879 45789 62957 45835
rect 63003 45789 63081 45835
rect 63127 45789 63205 45835
rect 63251 45789 63329 45835
rect 63375 45789 63453 45835
rect 63499 45789 63577 45835
rect 63623 45789 63701 45835
rect 63747 45789 63825 45835
rect 63871 45789 63949 45835
rect 63995 45789 64073 45835
rect 64119 45789 64197 45835
rect 64243 45789 64321 45835
rect 64367 45789 64445 45835
rect 64491 45789 64569 45835
rect 64615 45789 64693 45835
rect 64739 45789 64817 45835
rect 64863 45789 64941 45835
rect 64987 45789 65065 45835
rect 65111 45789 65189 45835
rect 65235 45789 65313 45835
rect 65359 45789 65437 45835
rect 65483 45789 65561 45835
rect 65607 45789 65685 45835
rect 65731 45789 65809 45835
rect 65855 45789 65933 45835
rect 65979 45789 66057 45835
rect 66103 45789 66181 45835
rect 66227 45789 66305 45835
rect 66351 45789 66429 45835
rect 66475 45789 66553 45835
rect 66599 45789 66677 45835
rect 66723 45789 66801 45835
rect 66847 45789 66925 45835
rect 66971 45789 67049 45835
rect 67095 45789 67173 45835
rect 67219 45789 67297 45835
rect 67343 45789 67421 45835
rect 67467 45789 67545 45835
rect 67591 45789 67669 45835
rect 67715 45789 67793 45835
rect 67839 45789 67917 45835
rect 67963 45789 68041 45835
rect 68087 45789 68165 45835
rect 68211 45789 68289 45835
rect 68335 45789 68413 45835
rect 68459 45789 68537 45835
rect 68583 45789 68661 45835
rect 68707 45789 68785 45835
rect 68831 45789 68909 45835
rect 68955 45789 69033 45835
rect 69079 45789 69157 45835
rect 69203 45789 69281 45835
rect 69327 45789 69405 45835
rect 69451 45789 69529 45835
rect 69575 45789 69653 45835
rect 69699 45789 69777 45835
rect 69823 45789 69901 45835
rect 69947 45789 70025 45835
rect 70071 45789 70149 45835
rect 70195 45789 70273 45835
rect 70319 45789 70397 45835
rect 70443 45789 70521 45835
rect 70567 45789 70645 45835
rect 70691 45789 70769 45835
rect 70815 45789 70893 45835
rect 70939 45789 71017 45835
rect 71063 45789 71141 45835
rect 71187 45789 71265 45835
rect 71311 45789 71389 45835
rect 71435 45789 71513 45835
rect 71559 45789 71637 45835
rect 71683 45789 71761 45835
rect 71807 45789 71885 45835
rect 71931 45789 72009 45835
rect 72055 45789 72133 45835
rect 72179 45789 72257 45835
rect 72303 45789 72381 45835
rect 72427 45789 72505 45835
rect 72551 45789 72629 45835
rect 72675 45789 72753 45835
rect 72799 45789 72877 45835
rect 72923 45789 73001 45835
rect 73047 45789 73125 45835
rect 73171 45789 73249 45835
rect 73295 45789 73373 45835
rect 73419 45789 73497 45835
rect 73543 45789 73621 45835
rect 73667 45789 73745 45835
rect 73791 45789 73869 45835
rect 73915 45789 73993 45835
rect 74039 45789 74117 45835
rect 74163 45789 74241 45835
rect 74287 45789 74365 45835
rect 74411 45789 74489 45835
rect 74535 45789 74613 45835
rect 74659 45789 74737 45835
rect 74783 45789 74861 45835
rect 74907 45789 74985 45835
rect 75031 45789 75109 45835
rect 75155 45789 75233 45835
rect 75279 45789 75357 45835
rect 75403 45789 75481 45835
rect 75527 45789 75605 45835
rect 75651 45789 75729 45835
rect 75775 45789 75853 45835
rect 75899 45789 75977 45835
rect 76023 45789 76101 45835
rect 76147 45789 76225 45835
rect 76271 45789 76349 45835
rect 76395 45789 76473 45835
rect 76519 45789 76597 45835
rect 76643 45789 76721 45835
rect 76767 45789 76845 45835
rect 76891 45789 76969 45835
rect 77015 45789 77093 45835
rect 77139 45789 77217 45835
rect 77263 45789 77341 45835
rect 77387 45789 77465 45835
rect 77511 45789 77589 45835
rect 77635 45789 77713 45835
rect 77759 45789 77837 45835
rect 77883 45789 77961 45835
rect 78007 45789 78085 45835
rect 78131 45789 78209 45835
rect 78255 45789 78333 45835
rect 78379 45789 78457 45835
rect 78503 45789 78581 45835
rect 78627 45789 78705 45835
rect 78751 45789 78829 45835
rect 78875 45789 78953 45835
rect 78999 45789 79077 45835
rect 79123 45789 79201 45835
rect 79247 45789 79325 45835
rect 79371 45789 79449 45835
rect 79495 45789 79573 45835
rect 79619 45789 79697 45835
rect 79743 45789 79821 45835
rect 79867 45789 79945 45835
rect 79991 45789 80069 45835
rect 80115 45789 80193 45835
rect 80239 45789 80317 45835
rect 80363 45789 80441 45835
rect 80487 45789 80565 45835
rect 80611 45789 80689 45835
rect 80735 45789 80813 45835
rect 80859 45789 80937 45835
rect 80983 45789 81061 45835
rect 81107 45789 81185 45835
rect 81231 45789 81309 45835
rect 81355 45789 81433 45835
rect 81479 45789 81557 45835
rect 81603 45789 81681 45835
rect 81727 45789 81805 45835
rect 81851 45789 81929 45835
rect 81975 45789 82053 45835
rect 82099 45789 82177 45835
rect 82223 45789 82301 45835
rect 82347 45789 82425 45835
rect 82471 45789 82549 45835
rect 82595 45789 82673 45835
rect 82719 45789 82797 45835
rect 82843 45789 82921 45835
rect 82967 45789 83045 45835
rect 83091 45789 83169 45835
rect 83215 45789 83293 45835
rect 83339 45789 83417 45835
rect 83463 45789 83541 45835
rect 83587 45789 83665 45835
rect 83711 45789 83789 45835
rect 83835 45789 83913 45835
rect 83959 45789 84037 45835
rect 84083 45789 84161 45835
rect 84207 45789 84285 45835
rect 84331 45789 84409 45835
rect 84455 45789 84533 45835
rect 84579 45789 84657 45835
rect 84703 45789 84781 45835
rect 84827 45789 84905 45835
rect 84951 45789 85029 45835
rect 85075 45789 85153 45835
rect 85199 45789 85277 45835
rect 85323 45789 85401 45835
rect 85447 45789 85525 45835
rect 85571 45789 85649 45835
rect 85695 45789 85816 45835
rect 70 45711 85816 45789
rect 70 45665 89 45711
rect 135 45665 213 45711
rect 259 45665 337 45711
rect 383 45665 461 45711
rect 507 45665 585 45711
rect 631 45665 709 45711
rect 755 45665 833 45711
rect 879 45665 957 45711
rect 1003 45665 1081 45711
rect 1127 45665 1205 45711
rect 1251 45665 1329 45711
rect 1375 45665 1453 45711
rect 1499 45665 1577 45711
rect 1623 45665 1701 45711
rect 1747 45665 1825 45711
rect 1871 45665 1949 45711
rect 1995 45665 2073 45711
rect 2119 45665 2197 45711
rect 2243 45665 2321 45711
rect 2367 45665 2445 45711
rect 2491 45665 2569 45711
rect 2615 45665 2693 45711
rect 2739 45665 2817 45711
rect 2863 45665 2941 45711
rect 2987 45665 3065 45711
rect 3111 45665 3189 45711
rect 3235 45665 3313 45711
rect 3359 45665 3437 45711
rect 3483 45665 3561 45711
rect 3607 45665 3685 45711
rect 3731 45665 3809 45711
rect 3855 45665 3933 45711
rect 3979 45665 4057 45711
rect 4103 45665 4181 45711
rect 4227 45665 4305 45711
rect 4351 45665 4429 45711
rect 4475 45665 4553 45711
rect 4599 45665 4677 45711
rect 4723 45665 4801 45711
rect 4847 45665 4925 45711
rect 4971 45665 5049 45711
rect 5095 45665 5173 45711
rect 5219 45665 5297 45711
rect 5343 45665 5421 45711
rect 5467 45665 5545 45711
rect 5591 45665 5669 45711
rect 5715 45665 5793 45711
rect 5839 45665 5917 45711
rect 5963 45665 6041 45711
rect 6087 45665 6165 45711
rect 6211 45665 6289 45711
rect 6335 45665 6413 45711
rect 6459 45665 6537 45711
rect 6583 45665 6661 45711
rect 6707 45665 6785 45711
rect 6831 45665 6909 45711
rect 6955 45665 7033 45711
rect 7079 45665 7157 45711
rect 7203 45665 7281 45711
rect 7327 45665 7405 45711
rect 7451 45665 7529 45711
rect 7575 45665 7653 45711
rect 7699 45665 7777 45711
rect 7823 45665 7901 45711
rect 7947 45665 8025 45711
rect 8071 45665 8149 45711
rect 8195 45665 8273 45711
rect 8319 45665 8397 45711
rect 8443 45665 8521 45711
rect 8567 45665 8645 45711
rect 8691 45665 8769 45711
rect 8815 45665 8893 45711
rect 8939 45665 9017 45711
rect 9063 45665 9141 45711
rect 9187 45665 9265 45711
rect 9311 45665 9389 45711
rect 9435 45665 9513 45711
rect 9559 45665 9637 45711
rect 9683 45665 9761 45711
rect 9807 45665 9885 45711
rect 9931 45665 10009 45711
rect 10055 45665 10133 45711
rect 10179 45665 10257 45711
rect 10303 45665 10381 45711
rect 10427 45665 10505 45711
rect 10551 45665 10629 45711
rect 10675 45665 10753 45711
rect 10799 45665 10877 45711
rect 10923 45665 11001 45711
rect 11047 45665 11125 45711
rect 11171 45665 11249 45711
rect 11295 45665 11373 45711
rect 11419 45665 11497 45711
rect 11543 45665 11621 45711
rect 11667 45665 11745 45711
rect 11791 45665 11869 45711
rect 11915 45665 11993 45711
rect 12039 45665 12117 45711
rect 12163 45665 12241 45711
rect 12287 45665 12365 45711
rect 12411 45665 12489 45711
rect 12535 45665 12613 45711
rect 12659 45665 12737 45711
rect 12783 45665 12861 45711
rect 12907 45665 12985 45711
rect 13031 45665 13109 45711
rect 13155 45665 13233 45711
rect 13279 45665 13357 45711
rect 13403 45665 13481 45711
rect 13527 45665 13605 45711
rect 13651 45665 13729 45711
rect 13775 45665 13853 45711
rect 13899 45665 13977 45711
rect 14023 45665 14101 45711
rect 14147 45665 14225 45711
rect 14271 45665 14349 45711
rect 14395 45665 14473 45711
rect 14519 45665 14597 45711
rect 14643 45665 14721 45711
rect 14767 45665 14845 45711
rect 14891 45665 14969 45711
rect 15015 45665 15093 45711
rect 15139 45665 15217 45711
rect 15263 45665 15341 45711
rect 15387 45665 15465 45711
rect 15511 45665 15589 45711
rect 15635 45665 15713 45711
rect 15759 45665 15837 45711
rect 15883 45665 15961 45711
rect 16007 45665 16085 45711
rect 16131 45665 16209 45711
rect 16255 45665 16333 45711
rect 16379 45665 16457 45711
rect 16503 45665 16581 45711
rect 16627 45665 16705 45711
rect 16751 45665 16829 45711
rect 16875 45665 16953 45711
rect 16999 45665 17077 45711
rect 17123 45665 17201 45711
rect 17247 45665 17325 45711
rect 17371 45665 17449 45711
rect 17495 45665 17573 45711
rect 17619 45665 17697 45711
rect 17743 45665 17821 45711
rect 17867 45665 17945 45711
rect 17991 45665 18069 45711
rect 18115 45665 18193 45711
rect 18239 45665 18317 45711
rect 18363 45665 18441 45711
rect 18487 45665 18565 45711
rect 18611 45665 18689 45711
rect 18735 45665 18813 45711
rect 18859 45665 18937 45711
rect 18983 45665 19061 45711
rect 19107 45665 19185 45711
rect 19231 45665 19309 45711
rect 19355 45665 19433 45711
rect 19479 45665 19557 45711
rect 19603 45665 19681 45711
rect 19727 45665 19805 45711
rect 19851 45665 19929 45711
rect 19975 45665 20053 45711
rect 20099 45665 20177 45711
rect 20223 45665 20301 45711
rect 20347 45665 20425 45711
rect 20471 45665 20549 45711
rect 20595 45665 20673 45711
rect 20719 45665 20797 45711
rect 20843 45665 20921 45711
rect 20967 45665 21045 45711
rect 21091 45665 21169 45711
rect 21215 45665 21293 45711
rect 21339 45665 21417 45711
rect 21463 45665 21541 45711
rect 21587 45665 21665 45711
rect 21711 45665 21789 45711
rect 21835 45665 21913 45711
rect 21959 45665 22037 45711
rect 22083 45665 22161 45711
rect 22207 45665 22285 45711
rect 22331 45665 22409 45711
rect 22455 45665 22533 45711
rect 22579 45665 22657 45711
rect 22703 45665 22781 45711
rect 22827 45665 22905 45711
rect 22951 45665 23029 45711
rect 23075 45665 23153 45711
rect 23199 45665 23277 45711
rect 23323 45665 23401 45711
rect 23447 45665 23525 45711
rect 23571 45665 23649 45711
rect 23695 45665 23773 45711
rect 23819 45665 23897 45711
rect 23943 45665 24021 45711
rect 24067 45665 24145 45711
rect 24191 45665 24269 45711
rect 24315 45665 24393 45711
rect 24439 45665 24517 45711
rect 24563 45665 24641 45711
rect 24687 45665 24765 45711
rect 24811 45665 24889 45711
rect 24935 45665 25013 45711
rect 25059 45665 25137 45711
rect 25183 45665 25261 45711
rect 25307 45665 25385 45711
rect 25431 45665 25509 45711
rect 25555 45665 25633 45711
rect 25679 45665 25757 45711
rect 25803 45665 25881 45711
rect 25927 45665 26005 45711
rect 26051 45665 26129 45711
rect 26175 45665 26253 45711
rect 26299 45665 26377 45711
rect 26423 45665 26501 45711
rect 26547 45665 26625 45711
rect 26671 45665 26749 45711
rect 26795 45665 26873 45711
rect 26919 45665 26997 45711
rect 27043 45665 27121 45711
rect 27167 45665 27245 45711
rect 27291 45665 27369 45711
rect 27415 45665 27493 45711
rect 27539 45665 27617 45711
rect 27663 45665 27741 45711
rect 27787 45665 27865 45711
rect 27911 45665 27989 45711
rect 28035 45665 28113 45711
rect 28159 45665 28237 45711
rect 28283 45665 28361 45711
rect 28407 45665 28485 45711
rect 28531 45665 28609 45711
rect 28655 45665 28733 45711
rect 28779 45665 28857 45711
rect 28903 45665 28981 45711
rect 29027 45665 29105 45711
rect 29151 45665 29229 45711
rect 29275 45665 29353 45711
rect 29399 45665 29477 45711
rect 29523 45665 29601 45711
rect 29647 45665 29725 45711
rect 29771 45665 29849 45711
rect 29895 45665 29973 45711
rect 30019 45665 30097 45711
rect 30143 45665 30221 45711
rect 30267 45665 30345 45711
rect 30391 45665 30469 45711
rect 30515 45665 30593 45711
rect 30639 45665 30717 45711
rect 30763 45665 30841 45711
rect 30887 45665 30965 45711
rect 31011 45665 31089 45711
rect 31135 45665 31213 45711
rect 31259 45665 31337 45711
rect 31383 45665 31461 45711
rect 31507 45665 31585 45711
rect 31631 45665 31709 45711
rect 31755 45665 31833 45711
rect 31879 45665 31957 45711
rect 32003 45665 32081 45711
rect 32127 45665 32205 45711
rect 32251 45665 32329 45711
rect 32375 45665 32453 45711
rect 32499 45665 32577 45711
rect 32623 45665 32701 45711
rect 32747 45665 32825 45711
rect 32871 45665 32949 45711
rect 32995 45665 33073 45711
rect 33119 45665 33197 45711
rect 33243 45665 33321 45711
rect 33367 45665 33445 45711
rect 33491 45665 33569 45711
rect 33615 45665 33693 45711
rect 33739 45665 33817 45711
rect 33863 45665 33941 45711
rect 33987 45665 34065 45711
rect 34111 45665 34189 45711
rect 34235 45665 34313 45711
rect 34359 45665 34437 45711
rect 34483 45665 34561 45711
rect 34607 45665 34685 45711
rect 34731 45665 34809 45711
rect 34855 45665 34933 45711
rect 34979 45665 35057 45711
rect 35103 45665 35181 45711
rect 35227 45665 35305 45711
rect 35351 45665 35429 45711
rect 35475 45665 35553 45711
rect 35599 45665 35677 45711
rect 35723 45665 35801 45711
rect 35847 45665 35925 45711
rect 35971 45665 36049 45711
rect 36095 45665 36173 45711
rect 36219 45665 36297 45711
rect 36343 45665 36421 45711
rect 36467 45665 36545 45711
rect 36591 45665 36669 45711
rect 36715 45665 36793 45711
rect 36839 45665 36917 45711
rect 36963 45665 37041 45711
rect 37087 45665 37165 45711
rect 37211 45665 37289 45711
rect 37335 45665 37413 45711
rect 37459 45665 37537 45711
rect 37583 45665 37661 45711
rect 37707 45665 37785 45711
rect 37831 45665 37909 45711
rect 37955 45665 38033 45711
rect 38079 45665 38157 45711
rect 38203 45665 38281 45711
rect 38327 45665 38405 45711
rect 38451 45665 38529 45711
rect 38575 45665 38653 45711
rect 38699 45665 38777 45711
rect 38823 45665 38901 45711
rect 38947 45665 39025 45711
rect 39071 45665 39149 45711
rect 39195 45665 39273 45711
rect 39319 45665 39397 45711
rect 39443 45665 39521 45711
rect 39567 45665 39645 45711
rect 39691 45665 39769 45711
rect 39815 45665 39893 45711
rect 39939 45665 40017 45711
rect 40063 45665 40141 45711
rect 40187 45665 40265 45711
rect 40311 45665 40389 45711
rect 40435 45665 40513 45711
rect 40559 45665 40637 45711
rect 40683 45665 40761 45711
rect 40807 45665 40885 45711
rect 40931 45665 41009 45711
rect 41055 45665 41133 45711
rect 41179 45665 41257 45711
rect 41303 45665 41381 45711
rect 41427 45665 41505 45711
rect 41551 45665 41629 45711
rect 41675 45665 41753 45711
rect 41799 45665 41877 45711
rect 41923 45665 42001 45711
rect 42047 45665 42125 45711
rect 42171 45665 42249 45711
rect 42295 45665 42373 45711
rect 42419 45665 42497 45711
rect 42543 45665 42621 45711
rect 42667 45665 42745 45711
rect 42791 45665 42869 45711
rect 42915 45665 42993 45711
rect 43039 45665 43117 45711
rect 43163 45665 43241 45711
rect 43287 45665 43365 45711
rect 43411 45665 43489 45711
rect 43535 45665 43613 45711
rect 43659 45665 43737 45711
rect 43783 45665 43861 45711
rect 43907 45665 43985 45711
rect 44031 45665 44109 45711
rect 44155 45665 44233 45711
rect 44279 45665 44357 45711
rect 44403 45665 44481 45711
rect 44527 45665 44605 45711
rect 44651 45665 44729 45711
rect 44775 45665 44853 45711
rect 44899 45665 44977 45711
rect 45023 45665 45101 45711
rect 45147 45665 45225 45711
rect 45271 45665 45349 45711
rect 45395 45665 45473 45711
rect 45519 45665 45597 45711
rect 45643 45665 45721 45711
rect 45767 45665 45845 45711
rect 45891 45665 45969 45711
rect 46015 45665 46093 45711
rect 46139 45665 46217 45711
rect 46263 45665 46341 45711
rect 46387 45665 46465 45711
rect 46511 45665 46589 45711
rect 46635 45665 46713 45711
rect 46759 45665 46837 45711
rect 46883 45665 46961 45711
rect 47007 45665 47085 45711
rect 47131 45665 47209 45711
rect 47255 45665 47333 45711
rect 47379 45665 47457 45711
rect 47503 45665 47581 45711
rect 47627 45665 47705 45711
rect 47751 45665 47829 45711
rect 47875 45665 47953 45711
rect 47999 45665 48077 45711
rect 48123 45665 48201 45711
rect 48247 45665 48325 45711
rect 48371 45665 48449 45711
rect 48495 45665 48573 45711
rect 48619 45665 48697 45711
rect 48743 45665 48821 45711
rect 48867 45665 48945 45711
rect 48991 45665 49069 45711
rect 49115 45665 49193 45711
rect 49239 45665 49317 45711
rect 49363 45665 49441 45711
rect 49487 45665 49565 45711
rect 49611 45665 49689 45711
rect 49735 45665 49813 45711
rect 49859 45665 49937 45711
rect 49983 45665 50061 45711
rect 50107 45665 50185 45711
rect 50231 45665 50309 45711
rect 50355 45665 50433 45711
rect 50479 45665 50557 45711
rect 50603 45665 50681 45711
rect 50727 45665 50805 45711
rect 50851 45665 50929 45711
rect 50975 45665 51053 45711
rect 51099 45665 51177 45711
rect 51223 45665 51301 45711
rect 51347 45665 51425 45711
rect 51471 45665 51549 45711
rect 51595 45665 51673 45711
rect 51719 45665 51797 45711
rect 51843 45665 51921 45711
rect 51967 45665 52045 45711
rect 52091 45665 52169 45711
rect 52215 45665 52293 45711
rect 52339 45665 52417 45711
rect 52463 45665 52541 45711
rect 52587 45665 52665 45711
rect 52711 45665 52789 45711
rect 52835 45665 52913 45711
rect 52959 45665 53037 45711
rect 53083 45665 53161 45711
rect 53207 45665 53285 45711
rect 53331 45665 53409 45711
rect 53455 45665 53533 45711
rect 53579 45665 53657 45711
rect 53703 45665 53781 45711
rect 53827 45665 53905 45711
rect 53951 45665 54029 45711
rect 54075 45665 54153 45711
rect 54199 45665 54277 45711
rect 54323 45665 54401 45711
rect 54447 45665 54525 45711
rect 54571 45665 54649 45711
rect 54695 45665 54773 45711
rect 54819 45665 54897 45711
rect 54943 45665 55021 45711
rect 55067 45665 55145 45711
rect 55191 45665 55269 45711
rect 55315 45665 55393 45711
rect 55439 45665 55517 45711
rect 55563 45665 55641 45711
rect 55687 45665 55765 45711
rect 55811 45665 55889 45711
rect 55935 45665 56013 45711
rect 56059 45665 56137 45711
rect 56183 45665 56261 45711
rect 56307 45665 56385 45711
rect 56431 45665 56509 45711
rect 56555 45665 56633 45711
rect 56679 45665 56757 45711
rect 56803 45665 56881 45711
rect 56927 45665 57005 45711
rect 57051 45665 57129 45711
rect 57175 45665 57253 45711
rect 57299 45665 57377 45711
rect 57423 45665 57501 45711
rect 57547 45665 57625 45711
rect 57671 45665 57749 45711
rect 57795 45665 57873 45711
rect 57919 45665 57997 45711
rect 58043 45665 58121 45711
rect 58167 45665 58245 45711
rect 58291 45665 58369 45711
rect 58415 45665 58493 45711
rect 58539 45665 58617 45711
rect 58663 45665 58741 45711
rect 58787 45665 58865 45711
rect 58911 45665 58989 45711
rect 59035 45665 59113 45711
rect 59159 45665 59237 45711
rect 59283 45665 59361 45711
rect 59407 45665 59485 45711
rect 59531 45665 59609 45711
rect 59655 45665 59733 45711
rect 59779 45665 59857 45711
rect 59903 45665 59981 45711
rect 60027 45665 60105 45711
rect 60151 45665 60229 45711
rect 60275 45665 60353 45711
rect 60399 45665 60477 45711
rect 60523 45665 60601 45711
rect 60647 45665 60725 45711
rect 60771 45665 60849 45711
rect 60895 45665 60973 45711
rect 61019 45665 61097 45711
rect 61143 45665 61221 45711
rect 61267 45665 61345 45711
rect 61391 45665 61469 45711
rect 61515 45665 61593 45711
rect 61639 45665 61717 45711
rect 61763 45665 61841 45711
rect 61887 45665 61965 45711
rect 62011 45665 62089 45711
rect 62135 45665 62213 45711
rect 62259 45665 62337 45711
rect 62383 45665 62461 45711
rect 62507 45665 62585 45711
rect 62631 45665 62709 45711
rect 62755 45665 62833 45711
rect 62879 45665 62957 45711
rect 63003 45665 63081 45711
rect 63127 45665 63205 45711
rect 63251 45665 63329 45711
rect 63375 45665 63453 45711
rect 63499 45665 63577 45711
rect 63623 45665 63701 45711
rect 63747 45665 63825 45711
rect 63871 45665 63949 45711
rect 63995 45665 64073 45711
rect 64119 45665 64197 45711
rect 64243 45665 64321 45711
rect 64367 45665 64445 45711
rect 64491 45665 64569 45711
rect 64615 45665 64693 45711
rect 64739 45665 64817 45711
rect 64863 45665 64941 45711
rect 64987 45665 65065 45711
rect 65111 45665 65189 45711
rect 65235 45665 65313 45711
rect 65359 45665 65437 45711
rect 65483 45665 65561 45711
rect 65607 45665 65685 45711
rect 65731 45665 65809 45711
rect 65855 45665 65933 45711
rect 65979 45665 66057 45711
rect 66103 45665 66181 45711
rect 66227 45665 66305 45711
rect 66351 45665 66429 45711
rect 66475 45665 66553 45711
rect 66599 45665 66677 45711
rect 66723 45665 66801 45711
rect 66847 45665 66925 45711
rect 66971 45665 67049 45711
rect 67095 45665 67173 45711
rect 67219 45665 67297 45711
rect 67343 45665 67421 45711
rect 67467 45665 67545 45711
rect 67591 45665 67669 45711
rect 67715 45665 67793 45711
rect 67839 45665 67917 45711
rect 67963 45665 68041 45711
rect 68087 45665 68165 45711
rect 68211 45665 68289 45711
rect 68335 45665 68413 45711
rect 68459 45665 68537 45711
rect 68583 45665 68661 45711
rect 68707 45665 68785 45711
rect 68831 45665 68909 45711
rect 68955 45665 69033 45711
rect 69079 45665 69157 45711
rect 69203 45665 69281 45711
rect 69327 45665 69405 45711
rect 69451 45665 69529 45711
rect 69575 45665 69653 45711
rect 69699 45665 69777 45711
rect 69823 45665 69901 45711
rect 69947 45665 70025 45711
rect 70071 45665 70149 45711
rect 70195 45665 70273 45711
rect 70319 45665 70397 45711
rect 70443 45665 70521 45711
rect 70567 45665 70645 45711
rect 70691 45665 70769 45711
rect 70815 45665 70893 45711
rect 70939 45665 71017 45711
rect 71063 45665 71141 45711
rect 71187 45665 71265 45711
rect 71311 45665 71389 45711
rect 71435 45665 71513 45711
rect 71559 45665 71637 45711
rect 71683 45665 71761 45711
rect 71807 45665 71885 45711
rect 71931 45665 72009 45711
rect 72055 45665 72133 45711
rect 72179 45665 72257 45711
rect 72303 45665 72381 45711
rect 72427 45665 72505 45711
rect 72551 45665 72629 45711
rect 72675 45665 72753 45711
rect 72799 45665 72877 45711
rect 72923 45665 73001 45711
rect 73047 45665 73125 45711
rect 73171 45665 73249 45711
rect 73295 45665 73373 45711
rect 73419 45665 73497 45711
rect 73543 45665 73621 45711
rect 73667 45665 73745 45711
rect 73791 45665 73869 45711
rect 73915 45665 73993 45711
rect 74039 45665 74117 45711
rect 74163 45665 74241 45711
rect 74287 45665 74365 45711
rect 74411 45665 74489 45711
rect 74535 45665 74613 45711
rect 74659 45665 74737 45711
rect 74783 45665 74861 45711
rect 74907 45665 74985 45711
rect 75031 45665 75109 45711
rect 75155 45665 75233 45711
rect 75279 45665 75357 45711
rect 75403 45665 75481 45711
rect 75527 45665 75605 45711
rect 75651 45665 75729 45711
rect 75775 45665 75853 45711
rect 75899 45665 75977 45711
rect 76023 45665 76101 45711
rect 76147 45665 76225 45711
rect 76271 45665 76349 45711
rect 76395 45665 76473 45711
rect 76519 45665 76597 45711
rect 76643 45665 76721 45711
rect 76767 45665 76845 45711
rect 76891 45665 76969 45711
rect 77015 45665 77093 45711
rect 77139 45665 77217 45711
rect 77263 45665 77341 45711
rect 77387 45665 77465 45711
rect 77511 45665 77589 45711
rect 77635 45665 77713 45711
rect 77759 45665 77837 45711
rect 77883 45665 77961 45711
rect 78007 45665 78085 45711
rect 78131 45665 78209 45711
rect 78255 45665 78333 45711
rect 78379 45665 78457 45711
rect 78503 45665 78581 45711
rect 78627 45665 78705 45711
rect 78751 45665 78829 45711
rect 78875 45665 78953 45711
rect 78999 45665 79077 45711
rect 79123 45665 79201 45711
rect 79247 45665 79325 45711
rect 79371 45665 79449 45711
rect 79495 45665 79573 45711
rect 79619 45665 79697 45711
rect 79743 45665 79821 45711
rect 79867 45665 79945 45711
rect 79991 45665 80069 45711
rect 80115 45665 80193 45711
rect 80239 45665 80317 45711
rect 80363 45665 80441 45711
rect 80487 45665 80565 45711
rect 80611 45665 80689 45711
rect 80735 45665 80813 45711
rect 80859 45665 80937 45711
rect 80983 45665 81061 45711
rect 81107 45665 81185 45711
rect 81231 45665 81309 45711
rect 81355 45665 81433 45711
rect 81479 45665 81557 45711
rect 81603 45665 81681 45711
rect 81727 45665 81805 45711
rect 81851 45665 81929 45711
rect 81975 45665 82053 45711
rect 82099 45665 82177 45711
rect 82223 45665 82301 45711
rect 82347 45665 82425 45711
rect 82471 45665 82549 45711
rect 82595 45665 82673 45711
rect 82719 45665 82797 45711
rect 82843 45665 82921 45711
rect 82967 45665 83045 45711
rect 83091 45665 83169 45711
rect 83215 45665 83293 45711
rect 83339 45665 83417 45711
rect 83463 45665 83541 45711
rect 83587 45665 83665 45711
rect 83711 45665 83789 45711
rect 83835 45665 83913 45711
rect 83959 45665 84037 45711
rect 84083 45665 84161 45711
rect 84207 45665 84285 45711
rect 84331 45665 84409 45711
rect 84455 45665 84533 45711
rect 84579 45665 84657 45711
rect 84703 45665 84781 45711
rect 84827 45665 84905 45711
rect 84951 45665 85029 45711
rect 85075 45665 85153 45711
rect 85199 45665 85277 45711
rect 85323 45665 85401 45711
rect 85447 45665 85525 45711
rect 85571 45665 85649 45711
rect 85695 45665 85816 45711
rect 70 45646 85816 45665
rect 70 45563 454 45646
rect 70 1117 89 45563
rect 435 1117 454 45563
rect 70 1034 454 1117
rect 85432 45563 85816 45646
rect 85432 1117 85451 45563
rect 85797 1117 85816 45563
rect 85432 1034 85816 1117
rect 70 1015 85816 1034
rect 70 969 89 1015
rect 135 969 213 1015
rect 259 969 337 1015
rect 383 969 461 1015
rect 507 969 585 1015
rect 631 969 709 1015
rect 755 969 833 1015
rect 879 969 957 1015
rect 1003 969 1081 1015
rect 1127 969 1205 1015
rect 1251 969 1329 1015
rect 1375 969 1453 1015
rect 1499 969 1577 1015
rect 1623 969 1701 1015
rect 1747 969 1825 1015
rect 1871 969 1949 1015
rect 1995 969 2073 1015
rect 2119 969 2197 1015
rect 2243 969 2321 1015
rect 2367 969 2445 1015
rect 2491 969 2569 1015
rect 2615 969 2693 1015
rect 2739 969 2817 1015
rect 2863 969 2941 1015
rect 2987 969 3065 1015
rect 3111 969 3189 1015
rect 3235 969 3313 1015
rect 3359 969 3437 1015
rect 3483 969 3561 1015
rect 3607 969 3685 1015
rect 3731 969 3809 1015
rect 3855 969 3933 1015
rect 3979 969 4057 1015
rect 4103 969 4181 1015
rect 4227 969 4305 1015
rect 4351 969 4429 1015
rect 4475 969 4553 1015
rect 4599 969 4677 1015
rect 4723 969 4801 1015
rect 4847 969 4925 1015
rect 4971 969 5049 1015
rect 5095 969 5173 1015
rect 5219 969 5297 1015
rect 5343 969 5421 1015
rect 5467 969 5545 1015
rect 5591 969 5669 1015
rect 5715 969 5793 1015
rect 5839 969 5917 1015
rect 5963 969 6041 1015
rect 6087 969 6165 1015
rect 6211 969 6289 1015
rect 6335 969 6413 1015
rect 6459 969 6537 1015
rect 6583 969 6661 1015
rect 6707 969 6785 1015
rect 6831 969 6909 1015
rect 6955 969 7033 1015
rect 7079 969 7157 1015
rect 7203 969 7281 1015
rect 7327 969 7405 1015
rect 7451 969 7529 1015
rect 7575 969 7653 1015
rect 7699 969 7777 1015
rect 7823 969 7901 1015
rect 7947 969 8025 1015
rect 8071 969 8149 1015
rect 8195 969 8273 1015
rect 8319 969 8397 1015
rect 8443 969 8521 1015
rect 8567 969 8645 1015
rect 8691 969 8769 1015
rect 8815 969 8893 1015
rect 8939 969 9017 1015
rect 9063 969 9141 1015
rect 9187 969 9265 1015
rect 9311 969 9389 1015
rect 9435 969 9513 1015
rect 9559 969 9637 1015
rect 9683 969 9761 1015
rect 9807 969 9885 1015
rect 9931 969 10009 1015
rect 10055 969 10133 1015
rect 10179 969 10257 1015
rect 10303 969 10381 1015
rect 10427 969 10505 1015
rect 10551 969 10629 1015
rect 10675 969 10753 1015
rect 10799 969 10877 1015
rect 10923 969 11001 1015
rect 11047 969 11125 1015
rect 11171 969 11249 1015
rect 11295 969 11373 1015
rect 11419 969 11497 1015
rect 11543 969 11621 1015
rect 11667 969 11745 1015
rect 11791 969 11869 1015
rect 11915 969 11993 1015
rect 12039 969 12117 1015
rect 12163 969 12241 1015
rect 12287 969 12365 1015
rect 12411 969 12489 1015
rect 12535 969 12613 1015
rect 12659 969 12737 1015
rect 12783 969 12861 1015
rect 12907 969 12985 1015
rect 13031 969 13109 1015
rect 13155 969 13233 1015
rect 13279 969 13357 1015
rect 13403 969 13481 1015
rect 13527 969 13605 1015
rect 13651 969 13729 1015
rect 13775 969 13853 1015
rect 13899 969 13977 1015
rect 14023 969 14101 1015
rect 14147 969 14225 1015
rect 14271 969 14349 1015
rect 14395 969 14473 1015
rect 14519 969 14597 1015
rect 14643 969 14721 1015
rect 14767 969 14845 1015
rect 14891 969 14969 1015
rect 15015 969 15093 1015
rect 15139 969 15217 1015
rect 15263 969 15341 1015
rect 15387 969 15465 1015
rect 15511 969 15589 1015
rect 15635 969 15713 1015
rect 15759 969 15837 1015
rect 15883 969 15961 1015
rect 16007 969 16085 1015
rect 16131 969 16209 1015
rect 16255 969 16333 1015
rect 16379 969 16457 1015
rect 16503 969 16581 1015
rect 16627 969 16705 1015
rect 16751 969 16829 1015
rect 16875 969 16953 1015
rect 16999 969 17077 1015
rect 17123 969 17201 1015
rect 17247 969 17325 1015
rect 17371 969 17449 1015
rect 17495 969 17573 1015
rect 17619 969 17697 1015
rect 17743 969 17821 1015
rect 17867 969 17945 1015
rect 17991 969 18069 1015
rect 18115 969 18193 1015
rect 18239 969 18317 1015
rect 18363 969 18441 1015
rect 18487 969 18565 1015
rect 18611 969 18689 1015
rect 18735 969 18813 1015
rect 18859 969 18937 1015
rect 18983 969 19061 1015
rect 19107 969 19185 1015
rect 19231 969 19309 1015
rect 19355 969 19433 1015
rect 19479 969 19557 1015
rect 19603 969 19681 1015
rect 19727 969 19805 1015
rect 19851 969 19929 1015
rect 19975 969 20053 1015
rect 20099 969 20177 1015
rect 20223 969 20301 1015
rect 20347 969 20425 1015
rect 20471 969 20549 1015
rect 20595 969 20673 1015
rect 20719 969 20797 1015
rect 20843 969 20921 1015
rect 20967 969 21045 1015
rect 21091 969 21169 1015
rect 21215 969 21293 1015
rect 21339 969 21417 1015
rect 21463 969 21541 1015
rect 21587 969 21665 1015
rect 21711 969 21789 1015
rect 21835 969 21913 1015
rect 21959 969 22037 1015
rect 22083 969 22161 1015
rect 22207 969 22285 1015
rect 22331 969 22409 1015
rect 22455 969 22533 1015
rect 22579 969 22657 1015
rect 22703 969 22781 1015
rect 22827 969 22905 1015
rect 22951 969 23029 1015
rect 23075 969 23153 1015
rect 23199 969 23277 1015
rect 23323 969 23401 1015
rect 23447 969 23525 1015
rect 23571 969 23649 1015
rect 23695 969 23773 1015
rect 23819 969 23897 1015
rect 23943 969 24021 1015
rect 24067 969 24145 1015
rect 24191 969 24269 1015
rect 24315 969 24393 1015
rect 24439 969 24517 1015
rect 24563 969 24641 1015
rect 24687 969 24765 1015
rect 24811 969 24889 1015
rect 24935 969 25013 1015
rect 25059 969 25137 1015
rect 25183 969 25261 1015
rect 25307 969 25385 1015
rect 25431 969 25509 1015
rect 25555 969 25633 1015
rect 25679 969 25757 1015
rect 25803 969 25881 1015
rect 25927 969 26005 1015
rect 26051 969 26129 1015
rect 26175 969 26253 1015
rect 26299 969 26377 1015
rect 26423 969 26501 1015
rect 26547 969 26625 1015
rect 26671 969 26749 1015
rect 26795 969 26873 1015
rect 26919 969 26997 1015
rect 27043 969 27121 1015
rect 27167 969 27245 1015
rect 27291 969 27369 1015
rect 27415 969 27493 1015
rect 27539 969 27617 1015
rect 27663 969 27741 1015
rect 27787 969 27865 1015
rect 27911 969 27989 1015
rect 28035 969 28113 1015
rect 28159 969 28237 1015
rect 28283 969 28361 1015
rect 28407 969 28485 1015
rect 28531 969 28609 1015
rect 28655 969 28733 1015
rect 28779 969 28857 1015
rect 28903 969 28981 1015
rect 29027 969 29105 1015
rect 29151 969 29229 1015
rect 29275 969 29353 1015
rect 29399 969 29477 1015
rect 29523 969 29601 1015
rect 29647 969 29725 1015
rect 29771 969 29849 1015
rect 29895 969 29973 1015
rect 30019 969 30097 1015
rect 30143 969 30221 1015
rect 30267 969 30345 1015
rect 30391 969 30469 1015
rect 30515 969 30593 1015
rect 30639 969 30717 1015
rect 30763 969 30841 1015
rect 30887 969 30965 1015
rect 31011 969 31089 1015
rect 31135 969 31213 1015
rect 31259 969 31337 1015
rect 31383 969 31461 1015
rect 31507 969 31585 1015
rect 31631 969 31709 1015
rect 31755 969 31833 1015
rect 31879 969 31957 1015
rect 32003 969 32081 1015
rect 32127 969 32205 1015
rect 32251 969 32329 1015
rect 32375 969 32453 1015
rect 32499 969 32577 1015
rect 32623 969 32701 1015
rect 32747 969 32825 1015
rect 32871 969 32949 1015
rect 32995 969 33073 1015
rect 33119 969 33197 1015
rect 33243 969 33321 1015
rect 33367 969 33445 1015
rect 33491 969 33569 1015
rect 33615 969 33693 1015
rect 33739 969 33817 1015
rect 33863 969 33941 1015
rect 33987 969 34065 1015
rect 34111 969 34189 1015
rect 34235 969 34313 1015
rect 34359 969 34437 1015
rect 34483 969 34561 1015
rect 34607 969 34685 1015
rect 34731 969 34809 1015
rect 34855 969 34933 1015
rect 34979 969 35057 1015
rect 35103 969 35181 1015
rect 35227 969 35305 1015
rect 35351 969 35429 1015
rect 35475 969 35553 1015
rect 35599 969 35677 1015
rect 35723 969 35801 1015
rect 35847 969 35925 1015
rect 35971 969 36049 1015
rect 36095 969 36173 1015
rect 36219 969 36297 1015
rect 36343 969 36421 1015
rect 36467 969 36545 1015
rect 36591 969 36669 1015
rect 36715 969 36793 1015
rect 36839 969 36917 1015
rect 36963 969 37041 1015
rect 37087 969 37165 1015
rect 37211 969 37289 1015
rect 37335 969 37413 1015
rect 37459 969 37537 1015
rect 37583 969 37661 1015
rect 37707 969 37785 1015
rect 37831 969 37909 1015
rect 37955 969 38033 1015
rect 38079 969 38157 1015
rect 38203 969 38281 1015
rect 38327 969 38405 1015
rect 38451 969 38529 1015
rect 38575 969 38653 1015
rect 38699 969 38777 1015
rect 38823 969 38901 1015
rect 38947 969 39025 1015
rect 39071 969 39149 1015
rect 39195 969 39273 1015
rect 39319 969 39397 1015
rect 39443 969 39521 1015
rect 39567 969 39645 1015
rect 39691 969 39769 1015
rect 39815 969 39893 1015
rect 39939 969 40017 1015
rect 40063 969 40141 1015
rect 40187 969 40265 1015
rect 40311 969 40389 1015
rect 40435 969 40513 1015
rect 40559 969 40637 1015
rect 40683 969 40761 1015
rect 40807 969 40885 1015
rect 40931 969 41009 1015
rect 41055 969 41133 1015
rect 41179 969 41257 1015
rect 41303 969 41381 1015
rect 41427 969 41505 1015
rect 41551 969 41629 1015
rect 41675 969 41753 1015
rect 41799 969 41877 1015
rect 41923 969 42001 1015
rect 42047 969 42125 1015
rect 42171 969 42249 1015
rect 42295 969 42373 1015
rect 42419 969 42497 1015
rect 42543 969 42621 1015
rect 42667 969 42745 1015
rect 42791 969 42869 1015
rect 42915 969 42993 1015
rect 43039 969 43117 1015
rect 43163 969 43241 1015
rect 43287 969 43365 1015
rect 43411 969 43489 1015
rect 43535 969 43613 1015
rect 43659 969 43737 1015
rect 43783 969 43861 1015
rect 43907 969 43985 1015
rect 44031 969 44109 1015
rect 44155 969 44233 1015
rect 44279 969 44357 1015
rect 44403 969 44481 1015
rect 44527 969 44605 1015
rect 44651 969 44729 1015
rect 44775 969 44853 1015
rect 44899 969 44977 1015
rect 45023 969 45101 1015
rect 45147 969 45225 1015
rect 45271 969 45349 1015
rect 45395 969 45473 1015
rect 45519 969 45597 1015
rect 45643 969 45721 1015
rect 45767 969 45845 1015
rect 45891 969 45969 1015
rect 46015 969 46093 1015
rect 46139 969 46217 1015
rect 46263 969 46341 1015
rect 46387 969 46465 1015
rect 46511 969 46589 1015
rect 46635 969 46713 1015
rect 46759 969 46837 1015
rect 46883 969 46961 1015
rect 47007 969 47085 1015
rect 47131 969 47209 1015
rect 47255 969 47333 1015
rect 47379 969 47457 1015
rect 47503 969 47581 1015
rect 47627 969 47705 1015
rect 47751 969 47829 1015
rect 47875 969 47953 1015
rect 47999 969 48077 1015
rect 48123 969 48201 1015
rect 48247 969 48325 1015
rect 48371 969 48449 1015
rect 48495 969 48573 1015
rect 48619 969 48697 1015
rect 48743 969 48821 1015
rect 48867 969 48945 1015
rect 48991 969 49069 1015
rect 49115 969 49193 1015
rect 49239 969 49317 1015
rect 49363 969 49441 1015
rect 49487 969 49565 1015
rect 49611 969 49689 1015
rect 49735 969 49813 1015
rect 49859 969 49937 1015
rect 49983 969 50061 1015
rect 50107 969 50185 1015
rect 50231 969 50309 1015
rect 50355 969 50433 1015
rect 50479 969 50557 1015
rect 50603 969 50681 1015
rect 50727 969 50805 1015
rect 50851 969 50929 1015
rect 50975 969 51053 1015
rect 51099 969 51177 1015
rect 51223 969 51301 1015
rect 51347 969 51425 1015
rect 51471 969 51549 1015
rect 51595 969 51673 1015
rect 51719 969 51797 1015
rect 51843 969 51921 1015
rect 51967 969 52045 1015
rect 52091 969 52169 1015
rect 52215 969 52293 1015
rect 52339 969 52417 1015
rect 52463 969 52541 1015
rect 52587 969 52665 1015
rect 52711 969 52789 1015
rect 52835 969 52913 1015
rect 52959 969 53037 1015
rect 53083 969 53161 1015
rect 53207 969 53285 1015
rect 53331 969 53409 1015
rect 53455 969 53533 1015
rect 53579 969 53657 1015
rect 53703 969 53781 1015
rect 53827 969 53905 1015
rect 53951 969 54029 1015
rect 54075 969 54153 1015
rect 54199 969 54277 1015
rect 54323 969 54401 1015
rect 54447 969 54525 1015
rect 54571 969 54649 1015
rect 54695 969 54773 1015
rect 54819 969 54897 1015
rect 54943 969 55021 1015
rect 55067 969 55145 1015
rect 55191 969 55269 1015
rect 55315 969 55393 1015
rect 55439 969 55517 1015
rect 55563 969 55641 1015
rect 55687 969 55765 1015
rect 55811 969 55889 1015
rect 55935 969 56013 1015
rect 56059 969 56137 1015
rect 56183 969 56261 1015
rect 56307 969 56385 1015
rect 56431 969 56509 1015
rect 56555 969 56633 1015
rect 56679 969 56757 1015
rect 56803 969 56881 1015
rect 56927 969 57005 1015
rect 57051 969 57129 1015
rect 57175 969 57253 1015
rect 57299 969 57377 1015
rect 57423 969 57501 1015
rect 57547 969 57625 1015
rect 57671 969 57749 1015
rect 57795 969 57873 1015
rect 57919 969 57997 1015
rect 58043 969 58121 1015
rect 58167 969 58245 1015
rect 58291 969 58369 1015
rect 58415 969 58493 1015
rect 58539 969 58617 1015
rect 58663 969 58741 1015
rect 58787 969 58865 1015
rect 58911 969 58989 1015
rect 59035 969 59113 1015
rect 59159 969 59237 1015
rect 59283 969 59361 1015
rect 59407 969 59485 1015
rect 59531 969 59609 1015
rect 59655 969 59733 1015
rect 59779 969 59857 1015
rect 59903 969 59981 1015
rect 60027 969 60105 1015
rect 60151 969 60229 1015
rect 60275 969 60353 1015
rect 60399 969 60477 1015
rect 60523 969 60601 1015
rect 60647 969 60725 1015
rect 60771 969 60849 1015
rect 60895 969 60973 1015
rect 61019 969 61097 1015
rect 61143 969 61221 1015
rect 61267 969 61345 1015
rect 61391 969 61469 1015
rect 61515 969 61593 1015
rect 61639 969 61717 1015
rect 61763 969 61841 1015
rect 61887 969 61965 1015
rect 62011 969 62089 1015
rect 62135 969 62213 1015
rect 62259 969 62337 1015
rect 62383 969 62461 1015
rect 62507 969 62585 1015
rect 62631 969 62709 1015
rect 62755 969 62833 1015
rect 62879 969 62957 1015
rect 63003 969 63081 1015
rect 63127 969 63205 1015
rect 63251 969 63329 1015
rect 63375 969 63453 1015
rect 63499 969 63577 1015
rect 63623 969 63701 1015
rect 63747 969 63825 1015
rect 63871 969 63949 1015
rect 63995 969 64073 1015
rect 64119 969 64197 1015
rect 64243 969 64321 1015
rect 64367 969 64445 1015
rect 64491 969 64569 1015
rect 64615 969 64693 1015
rect 64739 969 64817 1015
rect 64863 969 64941 1015
rect 64987 969 65065 1015
rect 65111 969 65189 1015
rect 65235 969 65313 1015
rect 65359 969 65437 1015
rect 65483 969 65561 1015
rect 65607 969 65685 1015
rect 65731 969 65809 1015
rect 65855 969 65933 1015
rect 65979 969 66057 1015
rect 66103 969 66181 1015
rect 66227 969 66305 1015
rect 66351 969 66429 1015
rect 66475 969 66553 1015
rect 66599 969 66677 1015
rect 66723 969 66801 1015
rect 66847 969 66925 1015
rect 66971 969 67049 1015
rect 67095 969 67173 1015
rect 67219 969 67297 1015
rect 67343 969 67421 1015
rect 67467 969 67545 1015
rect 67591 969 67669 1015
rect 67715 969 67793 1015
rect 67839 969 67917 1015
rect 67963 969 68041 1015
rect 68087 969 68165 1015
rect 68211 969 68289 1015
rect 68335 969 68413 1015
rect 68459 969 68537 1015
rect 68583 969 68661 1015
rect 68707 969 68785 1015
rect 68831 969 68909 1015
rect 68955 969 69033 1015
rect 69079 969 69157 1015
rect 69203 969 69281 1015
rect 69327 969 69405 1015
rect 69451 969 69529 1015
rect 69575 969 69653 1015
rect 69699 969 69777 1015
rect 69823 969 69901 1015
rect 69947 969 70025 1015
rect 70071 969 70149 1015
rect 70195 969 70273 1015
rect 70319 969 70397 1015
rect 70443 969 70521 1015
rect 70567 969 70645 1015
rect 70691 969 70769 1015
rect 70815 969 70893 1015
rect 70939 969 71017 1015
rect 71063 969 71141 1015
rect 71187 969 71265 1015
rect 71311 969 71389 1015
rect 71435 969 71513 1015
rect 71559 969 71637 1015
rect 71683 969 71761 1015
rect 71807 969 71885 1015
rect 71931 969 72009 1015
rect 72055 969 72133 1015
rect 72179 969 72257 1015
rect 72303 969 72381 1015
rect 72427 969 72505 1015
rect 72551 969 72629 1015
rect 72675 969 72753 1015
rect 72799 969 72877 1015
rect 72923 969 73001 1015
rect 73047 969 73125 1015
rect 73171 969 73249 1015
rect 73295 969 73373 1015
rect 73419 969 73497 1015
rect 73543 969 73621 1015
rect 73667 969 73745 1015
rect 73791 969 73869 1015
rect 73915 969 73993 1015
rect 74039 969 74117 1015
rect 74163 969 74241 1015
rect 74287 969 74365 1015
rect 74411 969 74489 1015
rect 74535 969 74613 1015
rect 74659 969 74737 1015
rect 74783 969 74861 1015
rect 74907 969 74985 1015
rect 75031 969 75109 1015
rect 75155 969 75233 1015
rect 75279 969 75357 1015
rect 75403 969 75481 1015
rect 75527 969 75605 1015
rect 75651 969 75729 1015
rect 75775 969 75853 1015
rect 75899 969 75977 1015
rect 76023 969 76101 1015
rect 76147 969 76225 1015
rect 76271 969 76349 1015
rect 76395 969 76473 1015
rect 76519 969 76597 1015
rect 76643 969 76721 1015
rect 76767 969 76845 1015
rect 76891 969 76969 1015
rect 77015 969 77093 1015
rect 77139 969 77217 1015
rect 77263 969 77341 1015
rect 77387 969 77465 1015
rect 77511 969 77589 1015
rect 77635 969 77713 1015
rect 77759 969 77837 1015
rect 77883 969 77961 1015
rect 78007 969 78085 1015
rect 78131 969 78209 1015
rect 78255 969 78333 1015
rect 78379 969 78457 1015
rect 78503 969 78581 1015
rect 78627 969 78705 1015
rect 78751 969 78829 1015
rect 78875 969 78953 1015
rect 78999 969 79077 1015
rect 79123 969 79201 1015
rect 79247 969 79325 1015
rect 79371 969 79449 1015
rect 79495 969 79573 1015
rect 79619 969 79697 1015
rect 79743 969 79821 1015
rect 79867 969 79945 1015
rect 79991 969 80069 1015
rect 80115 969 80193 1015
rect 80239 969 80317 1015
rect 80363 969 80441 1015
rect 80487 969 80565 1015
rect 80611 969 80689 1015
rect 80735 969 80813 1015
rect 80859 969 80937 1015
rect 80983 969 81061 1015
rect 81107 969 81185 1015
rect 81231 969 81309 1015
rect 81355 969 81433 1015
rect 81479 969 81557 1015
rect 81603 969 81681 1015
rect 81727 969 81805 1015
rect 81851 969 81929 1015
rect 81975 969 82053 1015
rect 82099 969 82177 1015
rect 82223 969 82301 1015
rect 82347 969 82425 1015
rect 82471 969 82549 1015
rect 82595 969 82673 1015
rect 82719 969 82797 1015
rect 82843 969 82921 1015
rect 82967 969 83045 1015
rect 83091 969 83169 1015
rect 83215 969 83293 1015
rect 83339 969 83417 1015
rect 83463 969 83541 1015
rect 83587 969 83665 1015
rect 83711 969 83789 1015
rect 83835 969 83913 1015
rect 83959 969 84037 1015
rect 84083 969 84161 1015
rect 84207 969 84285 1015
rect 84331 969 84409 1015
rect 84455 969 84533 1015
rect 84579 969 84657 1015
rect 84703 969 84781 1015
rect 84827 969 84905 1015
rect 84951 969 85029 1015
rect 85075 969 85153 1015
rect 85199 969 85277 1015
rect 85323 969 85401 1015
rect 85447 969 85525 1015
rect 85571 969 85649 1015
rect 85695 969 85816 1015
rect 70 891 85816 969
rect 70 845 89 891
rect 135 845 213 891
rect 259 845 337 891
rect 383 845 461 891
rect 507 845 585 891
rect 631 845 709 891
rect 755 845 833 891
rect 879 845 957 891
rect 1003 845 1081 891
rect 1127 845 1205 891
rect 1251 845 1329 891
rect 1375 845 1453 891
rect 1499 845 1577 891
rect 1623 845 1701 891
rect 1747 845 1825 891
rect 1871 845 1949 891
rect 1995 845 2073 891
rect 2119 845 2197 891
rect 2243 845 2321 891
rect 2367 845 2445 891
rect 2491 845 2569 891
rect 2615 845 2693 891
rect 2739 845 2817 891
rect 2863 845 2941 891
rect 2987 845 3065 891
rect 3111 845 3189 891
rect 3235 845 3313 891
rect 3359 845 3437 891
rect 3483 845 3561 891
rect 3607 845 3685 891
rect 3731 845 3809 891
rect 3855 845 3933 891
rect 3979 845 4057 891
rect 4103 845 4181 891
rect 4227 845 4305 891
rect 4351 845 4429 891
rect 4475 845 4553 891
rect 4599 845 4677 891
rect 4723 845 4801 891
rect 4847 845 4925 891
rect 4971 845 5049 891
rect 5095 845 5173 891
rect 5219 845 5297 891
rect 5343 845 5421 891
rect 5467 845 5545 891
rect 5591 845 5669 891
rect 5715 845 5793 891
rect 5839 845 5917 891
rect 5963 845 6041 891
rect 6087 845 6165 891
rect 6211 845 6289 891
rect 6335 845 6413 891
rect 6459 845 6537 891
rect 6583 845 6661 891
rect 6707 845 6785 891
rect 6831 845 6909 891
rect 6955 845 7033 891
rect 7079 845 7157 891
rect 7203 845 7281 891
rect 7327 845 7405 891
rect 7451 845 7529 891
rect 7575 845 7653 891
rect 7699 845 7777 891
rect 7823 845 7901 891
rect 7947 845 8025 891
rect 8071 845 8149 891
rect 8195 845 8273 891
rect 8319 845 8397 891
rect 8443 845 8521 891
rect 8567 845 8645 891
rect 8691 845 8769 891
rect 8815 845 8893 891
rect 8939 845 9017 891
rect 9063 845 9141 891
rect 9187 845 9265 891
rect 9311 845 9389 891
rect 9435 845 9513 891
rect 9559 845 9637 891
rect 9683 845 9761 891
rect 9807 845 9885 891
rect 9931 845 10009 891
rect 10055 845 10133 891
rect 10179 845 10257 891
rect 10303 845 10381 891
rect 10427 845 10505 891
rect 10551 845 10629 891
rect 10675 845 10753 891
rect 10799 845 10877 891
rect 10923 845 11001 891
rect 11047 845 11125 891
rect 11171 845 11249 891
rect 11295 845 11373 891
rect 11419 845 11497 891
rect 11543 845 11621 891
rect 11667 845 11745 891
rect 11791 845 11869 891
rect 11915 845 11993 891
rect 12039 845 12117 891
rect 12163 845 12241 891
rect 12287 845 12365 891
rect 12411 845 12489 891
rect 12535 845 12613 891
rect 12659 845 12737 891
rect 12783 845 12861 891
rect 12907 845 12985 891
rect 13031 845 13109 891
rect 13155 845 13233 891
rect 13279 845 13357 891
rect 13403 845 13481 891
rect 13527 845 13605 891
rect 13651 845 13729 891
rect 13775 845 13853 891
rect 13899 845 13977 891
rect 14023 845 14101 891
rect 14147 845 14225 891
rect 14271 845 14349 891
rect 14395 845 14473 891
rect 14519 845 14597 891
rect 14643 845 14721 891
rect 14767 845 14845 891
rect 14891 845 14969 891
rect 15015 845 15093 891
rect 15139 845 15217 891
rect 15263 845 15341 891
rect 15387 845 15465 891
rect 15511 845 15589 891
rect 15635 845 15713 891
rect 15759 845 15837 891
rect 15883 845 15961 891
rect 16007 845 16085 891
rect 16131 845 16209 891
rect 16255 845 16333 891
rect 16379 845 16457 891
rect 16503 845 16581 891
rect 16627 845 16705 891
rect 16751 845 16829 891
rect 16875 845 16953 891
rect 16999 845 17077 891
rect 17123 845 17201 891
rect 17247 845 17325 891
rect 17371 845 17449 891
rect 17495 845 17573 891
rect 17619 845 17697 891
rect 17743 845 17821 891
rect 17867 845 17945 891
rect 17991 845 18069 891
rect 18115 845 18193 891
rect 18239 845 18317 891
rect 18363 845 18441 891
rect 18487 845 18565 891
rect 18611 845 18689 891
rect 18735 845 18813 891
rect 18859 845 18937 891
rect 18983 845 19061 891
rect 19107 845 19185 891
rect 19231 845 19309 891
rect 19355 845 19433 891
rect 19479 845 19557 891
rect 19603 845 19681 891
rect 19727 845 19805 891
rect 19851 845 19929 891
rect 19975 845 20053 891
rect 20099 845 20177 891
rect 20223 845 20301 891
rect 20347 845 20425 891
rect 20471 845 20549 891
rect 20595 845 20673 891
rect 20719 845 20797 891
rect 20843 845 20921 891
rect 20967 845 21045 891
rect 21091 845 21169 891
rect 21215 845 21293 891
rect 21339 845 21417 891
rect 21463 845 21541 891
rect 21587 845 21665 891
rect 21711 845 21789 891
rect 21835 845 21913 891
rect 21959 845 22037 891
rect 22083 845 22161 891
rect 22207 845 22285 891
rect 22331 845 22409 891
rect 22455 845 22533 891
rect 22579 845 22657 891
rect 22703 845 22781 891
rect 22827 845 22905 891
rect 22951 845 23029 891
rect 23075 845 23153 891
rect 23199 845 23277 891
rect 23323 845 23401 891
rect 23447 845 23525 891
rect 23571 845 23649 891
rect 23695 845 23773 891
rect 23819 845 23897 891
rect 23943 845 24021 891
rect 24067 845 24145 891
rect 24191 845 24269 891
rect 24315 845 24393 891
rect 24439 845 24517 891
rect 24563 845 24641 891
rect 24687 845 24765 891
rect 24811 845 24889 891
rect 24935 845 25013 891
rect 25059 845 25137 891
rect 25183 845 25261 891
rect 25307 845 25385 891
rect 25431 845 25509 891
rect 25555 845 25633 891
rect 25679 845 25757 891
rect 25803 845 25881 891
rect 25927 845 26005 891
rect 26051 845 26129 891
rect 26175 845 26253 891
rect 26299 845 26377 891
rect 26423 845 26501 891
rect 26547 845 26625 891
rect 26671 845 26749 891
rect 26795 845 26873 891
rect 26919 845 26997 891
rect 27043 845 27121 891
rect 27167 845 27245 891
rect 27291 845 27369 891
rect 27415 845 27493 891
rect 27539 845 27617 891
rect 27663 845 27741 891
rect 27787 845 27865 891
rect 27911 845 27989 891
rect 28035 845 28113 891
rect 28159 845 28237 891
rect 28283 845 28361 891
rect 28407 845 28485 891
rect 28531 845 28609 891
rect 28655 845 28733 891
rect 28779 845 28857 891
rect 28903 845 28981 891
rect 29027 845 29105 891
rect 29151 845 29229 891
rect 29275 845 29353 891
rect 29399 845 29477 891
rect 29523 845 29601 891
rect 29647 845 29725 891
rect 29771 845 29849 891
rect 29895 845 29973 891
rect 30019 845 30097 891
rect 30143 845 30221 891
rect 30267 845 30345 891
rect 30391 845 30469 891
rect 30515 845 30593 891
rect 30639 845 30717 891
rect 30763 845 30841 891
rect 30887 845 30965 891
rect 31011 845 31089 891
rect 31135 845 31213 891
rect 31259 845 31337 891
rect 31383 845 31461 891
rect 31507 845 31585 891
rect 31631 845 31709 891
rect 31755 845 31833 891
rect 31879 845 31957 891
rect 32003 845 32081 891
rect 32127 845 32205 891
rect 32251 845 32329 891
rect 32375 845 32453 891
rect 32499 845 32577 891
rect 32623 845 32701 891
rect 32747 845 32825 891
rect 32871 845 32949 891
rect 32995 845 33073 891
rect 33119 845 33197 891
rect 33243 845 33321 891
rect 33367 845 33445 891
rect 33491 845 33569 891
rect 33615 845 33693 891
rect 33739 845 33817 891
rect 33863 845 33941 891
rect 33987 845 34065 891
rect 34111 845 34189 891
rect 34235 845 34313 891
rect 34359 845 34437 891
rect 34483 845 34561 891
rect 34607 845 34685 891
rect 34731 845 34809 891
rect 34855 845 34933 891
rect 34979 845 35057 891
rect 35103 845 35181 891
rect 35227 845 35305 891
rect 35351 845 35429 891
rect 35475 845 35553 891
rect 35599 845 35677 891
rect 35723 845 35801 891
rect 35847 845 35925 891
rect 35971 845 36049 891
rect 36095 845 36173 891
rect 36219 845 36297 891
rect 36343 845 36421 891
rect 36467 845 36545 891
rect 36591 845 36669 891
rect 36715 845 36793 891
rect 36839 845 36917 891
rect 36963 845 37041 891
rect 37087 845 37165 891
rect 37211 845 37289 891
rect 37335 845 37413 891
rect 37459 845 37537 891
rect 37583 845 37661 891
rect 37707 845 37785 891
rect 37831 845 37909 891
rect 37955 845 38033 891
rect 38079 845 38157 891
rect 38203 845 38281 891
rect 38327 845 38405 891
rect 38451 845 38529 891
rect 38575 845 38653 891
rect 38699 845 38777 891
rect 38823 845 38901 891
rect 38947 845 39025 891
rect 39071 845 39149 891
rect 39195 845 39273 891
rect 39319 845 39397 891
rect 39443 845 39521 891
rect 39567 845 39645 891
rect 39691 845 39769 891
rect 39815 845 39893 891
rect 39939 845 40017 891
rect 40063 845 40141 891
rect 40187 845 40265 891
rect 40311 845 40389 891
rect 40435 845 40513 891
rect 40559 845 40637 891
rect 40683 845 40761 891
rect 40807 845 40885 891
rect 40931 845 41009 891
rect 41055 845 41133 891
rect 41179 845 41257 891
rect 41303 845 41381 891
rect 41427 845 41505 891
rect 41551 845 41629 891
rect 41675 845 41753 891
rect 41799 845 41877 891
rect 41923 845 42001 891
rect 42047 845 42125 891
rect 42171 845 42249 891
rect 42295 845 42373 891
rect 42419 845 42497 891
rect 42543 845 42621 891
rect 42667 845 42745 891
rect 42791 845 42869 891
rect 42915 845 42993 891
rect 43039 845 43117 891
rect 43163 845 43241 891
rect 43287 845 43365 891
rect 43411 845 43489 891
rect 43535 845 43613 891
rect 43659 845 43737 891
rect 43783 845 43861 891
rect 43907 845 43985 891
rect 44031 845 44109 891
rect 44155 845 44233 891
rect 44279 845 44357 891
rect 44403 845 44481 891
rect 44527 845 44605 891
rect 44651 845 44729 891
rect 44775 845 44853 891
rect 44899 845 44977 891
rect 45023 845 45101 891
rect 45147 845 45225 891
rect 45271 845 45349 891
rect 45395 845 45473 891
rect 45519 845 45597 891
rect 45643 845 45721 891
rect 45767 845 45845 891
rect 45891 845 45969 891
rect 46015 845 46093 891
rect 46139 845 46217 891
rect 46263 845 46341 891
rect 46387 845 46465 891
rect 46511 845 46589 891
rect 46635 845 46713 891
rect 46759 845 46837 891
rect 46883 845 46961 891
rect 47007 845 47085 891
rect 47131 845 47209 891
rect 47255 845 47333 891
rect 47379 845 47457 891
rect 47503 845 47581 891
rect 47627 845 47705 891
rect 47751 845 47829 891
rect 47875 845 47953 891
rect 47999 845 48077 891
rect 48123 845 48201 891
rect 48247 845 48325 891
rect 48371 845 48449 891
rect 48495 845 48573 891
rect 48619 845 48697 891
rect 48743 845 48821 891
rect 48867 845 48945 891
rect 48991 845 49069 891
rect 49115 845 49193 891
rect 49239 845 49317 891
rect 49363 845 49441 891
rect 49487 845 49565 891
rect 49611 845 49689 891
rect 49735 845 49813 891
rect 49859 845 49937 891
rect 49983 845 50061 891
rect 50107 845 50185 891
rect 50231 845 50309 891
rect 50355 845 50433 891
rect 50479 845 50557 891
rect 50603 845 50681 891
rect 50727 845 50805 891
rect 50851 845 50929 891
rect 50975 845 51053 891
rect 51099 845 51177 891
rect 51223 845 51301 891
rect 51347 845 51425 891
rect 51471 845 51549 891
rect 51595 845 51673 891
rect 51719 845 51797 891
rect 51843 845 51921 891
rect 51967 845 52045 891
rect 52091 845 52169 891
rect 52215 845 52293 891
rect 52339 845 52417 891
rect 52463 845 52541 891
rect 52587 845 52665 891
rect 52711 845 52789 891
rect 52835 845 52913 891
rect 52959 845 53037 891
rect 53083 845 53161 891
rect 53207 845 53285 891
rect 53331 845 53409 891
rect 53455 845 53533 891
rect 53579 845 53657 891
rect 53703 845 53781 891
rect 53827 845 53905 891
rect 53951 845 54029 891
rect 54075 845 54153 891
rect 54199 845 54277 891
rect 54323 845 54401 891
rect 54447 845 54525 891
rect 54571 845 54649 891
rect 54695 845 54773 891
rect 54819 845 54897 891
rect 54943 845 55021 891
rect 55067 845 55145 891
rect 55191 845 55269 891
rect 55315 845 55393 891
rect 55439 845 55517 891
rect 55563 845 55641 891
rect 55687 845 55765 891
rect 55811 845 55889 891
rect 55935 845 56013 891
rect 56059 845 56137 891
rect 56183 845 56261 891
rect 56307 845 56385 891
rect 56431 845 56509 891
rect 56555 845 56633 891
rect 56679 845 56757 891
rect 56803 845 56881 891
rect 56927 845 57005 891
rect 57051 845 57129 891
rect 57175 845 57253 891
rect 57299 845 57377 891
rect 57423 845 57501 891
rect 57547 845 57625 891
rect 57671 845 57749 891
rect 57795 845 57873 891
rect 57919 845 57997 891
rect 58043 845 58121 891
rect 58167 845 58245 891
rect 58291 845 58369 891
rect 58415 845 58493 891
rect 58539 845 58617 891
rect 58663 845 58741 891
rect 58787 845 58865 891
rect 58911 845 58989 891
rect 59035 845 59113 891
rect 59159 845 59237 891
rect 59283 845 59361 891
rect 59407 845 59485 891
rect 59531 845 59609 891
rect 59655 845 59733 891
rect 59779 845 59857 891
rect 59903 845 59981 891
rect 60027 845 60105 891
rect 60151 845 60229 891
rect 60275 845 60353 891
rect 60399 845 60477 891
rect 60523 845 60601 891
rect 60647 845 60725 891
rect 60771 845 60849 891
rect 60895 845 60973 891
rect 61019 845 61097 891
rect 61143 845 61221 891
rect 61267 845 61345 891
rect 61391 845 61469 891
rect 61515 845 61593 891
rect 61639 845 61717 891
rect 61763 845 61841 891
rect 61887 845 61965 891
rect 62011 845 62089 891
rect 62135 845 62213 891
rect 62259 845 62337 891
rect 62383 845 62461 891
rect 62507 845 62585 891
rect 62631 845 62709 891
rect 62755 845 62833 891
rect 62879 845 62957 891
rect 63003 845 63081 891
rect 63127 845 63205 891
rect 63251 845 63329 891
rect 63375 845 63453 891
rect 63499 845 63577 891
rect 63623 845 63701 891
rect 63747 845 63825 891
rect 63871 845 63949 891
rect 63995 845 64073 891
rect 64119 845 64197 891
rect 64243 845 64321 891
rect 64367 845 64445 891
rect 64491 845 64569 891
rect 64615 845 64693 891
rect 64739 845 64817 891
rect 64863 845 64941 891
rect 64987 845 65065 891
rect 65111 845 65189 891
rect 65235 845 65313 891
rect 65359 845 65437 891
rect 65483 845 65561 891
rect 65607 845 65685 891
rect 65731 845 65809 891
rect 65855 845 65933 891
rect 65979 845 66057 891
rect 66103 845 66181 891
rect 66227 845 66305 891
rect 66351 845 66429 891
rect 66475 845 66553 891
rect 66599 845 66677 891
rect 66723 845 66801 891
rect 66847 845 66925 891
rect 66971 845 67049 891
rect 67095 845 67173 891
rect 67219 845 67297 891
rect 67343 845 67421 891
rect 67467 845 67545 891
rect 67591 845 67669 891
rect 67715 845 67793 891
rect 67839 845 67917 891
rect 67963 845 68041 891
rect 68087 845 68165 891
rect 68211 845 68289 891
rect 68335 845 68413 891
rect 68459 845 68537 891
rect 68583 845 68661 891
rect 68707 845 68785 891
rect 68831 845 68909 891
rect 68955 845 69033 891
rect 69079 845 69157 891
rect 69203 845 69281 891
rect 69327 845 69405 891
rect 69451 845 69529 891
rect 69575 845 69653 891
rect 69699 845 69777 891
rect 69823 845 69901 891
rect 69947 845 70025 891
rect 70071 845 70149 891
rect 70195 845 70273 891
rect 70319 845 70397 891
rect 70443 845 70521 891
rect 70567 845 70645 891
rect 70691 845 70769 891
rect 70815 845 70893 891
rect 70939 845 71017 891
rect 71063 845 71141 891
rect 71187 845 71265 891
rect 71311 845 71389 891
rect 71435 845 71513 891
rect 71559 845 71637 891
rect 71683 845 71761 891
rect 71807 845 71885 891
rect 71931 845 72009 891
rect 72055 845 72133 891
rect 72179 845 72257 891
rect 72303 845 72381 891
rect 72427 845 72505 891
rect 72551 845 72629 891
rect 72675 845 72753 891
rect 72799 845 72877 891
rect 72923 845 73001 891
rect 73047 845 73125 891
rect 73171 845 73249 891
rect 73295 845 73373 891
rect 73419 845 73497 891
rect 73543 845 73621 891
rect 73667 845 73745 891
rect 73791 845 73869 891
rect 73915 845 73993 891
rect 74039 845 74117 891
rect 74163 845 74241 891
rect 74287 845 74365 891
rect 74411 845 74489 891
rect 74535 845 74613 891
rect 74659 845 74737 891
rect 74783 845 74861 891
rect 74907 845 74985 891
rect 75031 845 75109 891
rect 75155 845 75233 891
rect 75279 845 75357 891
rect 75403 845 75481 891
rect 75527 845 75605 891
rect 75651 845 75729 891
rect 75775 845 75853 891
rect 75899 845 75977 891
rect 76023 845 76101 891
rect 76147 845 76225 891
rect 76271 845 76349 891
rect 76395 845 76473 891
rect 76519 845 76597 891
rect 76643 845 76721 891
rect 76767 845 76845 891
rect 76891 845 76969 891
rect 77015 845 77093 891
rect 77139 845 77217 891
rect 77263 845 77341 891
rect 77387 845 77465 891
rect 77511 845 77589 891
rect 77635 845 77713 891
rect 77759 845 77837 891
rect 77883 845 77961 891
rect 78007 845 78085 891
rect 78131 845 78209 891
rect 78255 845 78333 891
rect 78379 845 78457 891
rect 78503 845 78581 891
rect 78627 845 78705 891
rect 78751 845 78829 891
rect 78875 845 78953 891
rect 78999 845 79077 891
rect 79123 845 79201 891
rect 79247 845 79325 891
rect 79371 845 79449 891
rect 79495 845 79573 891
rect 79619 845 79697 891
rect 79743 845 79821 891
rect 79867 845 79945 891
rect 79991 845 80069 891
rect 80115 845 80193 891
rect 80239 845 80317 891
rect 80363 845 80441 891
rect 80487 845 80565 891
rect 80611 845 80689 891
rect 80735 845 80813 891
rect 80859 845 80937 891
rect 80983 845 81061 891
rect 81107 845 81185 891
rect 81231 845 81309 891
rect 81355 845 81433 891
rect 81479 845 81557 891
rect 81603 845 81681 891
rect 81727 845 81805 891
rect 81851 845 81929 891
rect 81975 845 82053 891
rect 82099 845 82177 891
rect 82223 845 82301 891
rect 82347 845 82425 891
rect 82471 845 82549 891
rect 82595 845 82673 891
rect 82719 845 82797 891
rect 82843 845 82921 891
rect 82967 845 83045 891
rect 83091 845 83169 891
rect 83215 845 83293 891
rect 83339 845 83417 891
rect 83463 845 83541 891
rect 83587 845 83665 891
rect 83711 845 83789 891
rect 83835 845 83913 891
rect 83959 845 84037 891
rect 84083 845 84161 891
rect 84207 845 84285 891
rect 84331 845 84409 891
rect 84455 845 84533 891
rect 84579 845 84657 891
rect 84703 845 84781 891
rect 84827 845 84905 891
rect 84951 845 85029 891
rect 85075 845 85153 891
rect 85199 845 85277 891
rect 85323 845 85401 891
rect 85447 845 85525 891
rect 85571 845 85649 891
rect 85695 845 85816 891
rect 70 767 85816 845
rect 70 721 89 767
rect 135 721 213 767
rect 259 721 337 767
rect 383 721 461 767
rect 507 721 585 767
rect 631 721 709 767
rect 755 721 833 767
rect 879 721 957 767
rect 1003 721 1081 767
rect 1127 721 1205 767
rect 1251 721 1329 767
rect 1375 721 1453 767
rect 1499 721 1577 767
rect 1623 721 1701 767
rect 1747 721 1825 767
rect 1871 721 1949 767
rect 1995 721 2073 767
rect 2119 721 2197 767
rect 2243 721 2321 767
rect 2367 721 2445 767
rect 2491 721 2569 767
rect 2615 721 2693 767
rect 2739 721 2817 767
rect 2863 721 2941 767
rect 2987 721 3065 767
rect 3111 721 3189 767
rect 3235 721 3313 767
rect 3359 721 3437 767
rect 3483 721 3561 767
rect 3607 721 3685 767
rect 3731 721 3809 767
rect 3855 721 3933 767
rect 3979 721 4057 767
rect 4103 721 4181 767
rect 4227 721 4305 767
rect 4351 721 4429 767
rect 4475 721 4553 767
rect 4599 721 4677 767
rect 4723 721 4801 767
rect 4847 721 4925 767
rect 4971 721 5049 767
rect 5095 721 5173 767
rect 5219 721 5297 767
rect 5343 721 5421 767
rect 5467 721 5545 767
rect 5591 721 5669 767
rect 5715 721 5793 767
rect 5839 721 5917 767
rect 5963 721 6041 767
rect 6087 721 6165 767
rect 6211 721 6289 767
rect 6335 721 6413 767
rect 6459 721 6537 767
rect 6583 721 6661 767
rect 6707 721 6785 767
rect 6831 721 6909 767
rect 6955 721 7033 767
rect 7079 721 7157 767
rect 7203 721 7281 767
rect 7327 721 7405 767
rect 7451 721 7529 767
rect 7575 721 7653 767
rect 7699 721 7777 767
rect 7823 721 7901 767
rect 7947 721 8025 767
rect 8071 721 8149 767
rect 8195 721 8273 767
rect 8319 721 8397 767
rect 8443 721 8521 767
rect 8567 721 8645 767
rect 8691 721 8769 767
rect 8815 721 8893 767
rect 8939 721 9017 767
rect 9063 721 9141 767
rect 9187 721 9265 767
rect 9311 721 9389 767
rect 9435 721 9513 767
rect 9559 721 9637 767
rect 9683 721 9761 767
rect 9807 721 9885 767
rect 9931 721 10009 767
rect 10055 721 10133 767
rect 10179 721 10257 767
rect 10303 721 10381 767
rect 10427 721 10505 767
rect 10551 721 10629 767
rect 10675 721 10753 767
rect 10799 721 10877 767
rect 10923 721 11001 767
rect 11047 721 11125 767
rect 11171 721 11249 767
rect 11295 721 11373 767
rect 11419 721 11497 767
rect 11543 721 11621 767
rect 11667 721 11745 767
rect 11791 721 11869 767
rect 11915 721 11993 767
rect 12039 721 12117 767
rect 12163 721 12241 767
rect 12287 721 12365 767
rect 12411 721 12489 767
rect 12535 721 12613 767
rect 12659 721 12737 767
rect 12783 721 12861 767
rect 12907 721 12985 767
rect 13031 721 13109 767
rect 13155 721 13233 767
rect 13279 721 13357 767
rect 13403 721 13481 767
rect 13527 721 13605 767
rect 13651 721 13729 767
rect 13775 721 13853 767
rect 13899 721 13977 767
rect 14023 721 14101 767
rect 14147 721 14225 767
rect 14271 721 14349 767
rect 14395 721 14473 767
rect 14519 721 14597 767
rect 14643 721 14721 767
rect 14767 721 14845 767
rect 14891 721 14969 767
rect 15015 721 15093 767
rect 15139 721 15217 767
rect 15263 721 15341 767
rect 15387 721 15465 767
rect 15511 721 15589 767
rect 15635 721 15713 767
rect 15759 721 15837 767
rect 15883 721 15961 767
rect 16007 721 16085 767
rect 16131 721 16209 767
rect 16255 721 16333 767
rect 16379 721 16457 767
rect 16503 721 16581 767
rect 16627 721 16705 767
rect 16751 721 16829 767
rect 16875 721 16953 767
rect 16999 721 17077 767
rect 17123 721 17201 767
rect 17247 721 17325 767
rect 17371 721 17449 767
rect 17495 721 17573 767
rect 17619 721 17697 767
rect 17743 721 17821 767
rect 17867 721 17945 767
rect 17991 721 18069 767
rect 18115 721 18193 767
rect 18239 721 18317 767
rect 18363 721 18441 767
rect 18487 721 18565 767
rect 18611 721 18689 767
rect 18735 721 18813 767
rect 18859 721 18937 767
rect 18983 721 19061 767
rect 19107 721 19185 767
rect 19231 721 19309 767
rect 19355 721 19433 767
rect 19479 721 19557 767
rect 19603 721 19681 767
rect 19727 721 19805 767
rect 19851 721 19929 767
rect 19975 721 20053 767
rect 20099 721 20177 767
rect 20223 721 20301 767
rect 20347 721 20425 767
rect 20471 721 20549 767
rect 20595 721 20673 767
rect 20719 721 20797 767
rect 20843 721 20921 767
rect 20967 721 21045 767
rect 21091 721 21169 767
rect 21215 721 21293 767
rect 21339 721 21417 767
rect 21463 721 21541 767
rect 21587 721 21665 767
rect 21711 721 21789 767
rect 21835 721 21913 767
rect 21959 721 22037 767
rect 22083 721 22161 767
rect 22207 721 22285 767
rect 22331 721 22409 767
rect 22455 721 22533 767
rect 22579 721 22657 767
rect 22703 721 22781 767
rect 22827 721 22905 767
rect 22951 721 23029 767
rect 23075 721 23153 767
rect 23199 721 23277 767
rect 23323 721 23401 767
rect 23447 721 23525 767
rect 23571 721 23649 767
rect 23695 721 23773 767
rect 23819 721 23897 767
rect 23943 721 24021 767
rect 24067 721 24145 767
rect 24191 721 24269 767
rect 24315 721 24393 767
rect 24439 721 24517 767
rect 24563 721 24641 767
rect 24687 721 24765 767
rect 24811 721 24889 767
rect 24935 721 25013 767
rect 25059 721 25137 767
rect 25183 721 25261 767
rect 25307 721 25385 767
rect 25431 721 25509 767
rect 25555 721 25633 767
rect 25679 721 25757 767
rect 25803 721 25881 767
rect 25927 721 26005 767
rect 26051 721 26129 767
rect 26175 721 26253 767
rect 26299 721 26377 767
rect 26423 721 26501 767
rect 26547 721 26625 767
rect 26671 721 26749 767
rect 26795 721 26873 767
rect 26919 721 26997 767
rect 27043 721 27121 767
rect 27167 721 27245 767
rect 27291 721 27369 767
rect 27415 721 27493 767
rect 27539 721 27617 767
rect 27663 721 27741 767
rect 27787 721 27865 767
rect 27911 721 27989 767
rect 28035 721 28113 767
rect 28159 721 28237 767
rect 28283 721 28361 767
rect 28407 721 28485 767
rect 28531 721 28609 767
rect 28655 721 28733 767
rect 28779 721 28857 767
rect 28903 721 28981 767
rect 29027 721 29105 767
rect 29151 721 29229 767
rect 29275 721 29353 767
rect 29399 721 29477 767
rect 29523 721 29601 767
rect 29647 721 29725 767
rect 29771 721 29849 767
rect 29895 721 29973 767
rect 30019 721 30097 767
rect 30143 721 30221 767
rect 30267 721 30345 767
rect 30391 721 30469 767
rect 30515 721 30593 767
rect 30639 721 30717 767
rect 30763 721 30841 767
rect 30887 721 30965 767
rect 31011 721 31089 767
rect 31135 721 31213 767
rect 31259 721 31337 767
rect 31383 721 31461 767
rect 31507 721 31585 767
rect 31631 721 31709 767
rect 31755 721 31833 767
rect 31879 721 31957 767
rect 32003 721 32081 767
rect 32127 721 32205 767
rect 32251 721 32329 767
rect 32375 721 32453 767
rect 32499 721 32577 767
rect 32623 721 32701 767
rect 32747 721 32825 767
rect 32871 721 32949 767
rect 32995 721 33073 767
rect 33119 721 33197 767
rect 33243 721 33321 767
rect 33367 721 33445 767
rect 33491 721 33569 767
rect 33615 721 33693 767
rect 33739 721 33817 767
rect 33863 721 33941 767
rect 33987 721 34065 767
rect 34111 721 34189 767
rect 34235 721 34313 767
rect 34359 721 34437 767
rect 34483 721 34561 767
rect 34607 721 34685 767
rect 34731 721 34809 767
rect 34855 721 34933 767
rect 34979 721 35057 767
rect 35103 721 35181 767
rect 35227 721 35305 767
rect 35351 721 35429 767
rect 35475 721 35553 767
rect 35599 721 35677 767
rect 35723 721 35801 767
rect 35847 721 35925 767
rect 35971 721 36049 767
rect 36095 721 36173 767
rect 36219 721 36297 767
rect 36343 721 36421 767
rect 36467 721 36545 767
rect 36591 721 36669 767
rect 36715 721 36793 767
rect 36839 721 36917 767
rect 36963 721 37041 767
rect 37087 721 37165 767
rect 37211 721 37289 767
rect 37335 721 37413 767
rect 37459 721 37537 767
rect 37583 721 37661 767
rect 37707 721 37785 767
rect 37831 721 37909 767
rect 37955 721 38033 767
rect 38079 721 38157 767
rect 38203 721 38281 767
rect 38327 721 38405 767
rect 38451 721 38529 767
rect 38575 721 38653 767
rect 38699 721 38777 767
rect 38823 721 38901 767
rect 38947 721 39025 767
rect 39071 721 39149 767
rect 39195 721 39273 767
rect 39319 721 39397 767
rect 39443 721 39521 767
rect 39567 721 39645 767
rect 39691 721 39769 767
rect 39815 721 39893 767
rect 39939 721 40017 767
rect 40063 721 40141 767
rect 40187 721 40265 767
rect 40311 721 40389 767
rect 40435 721 40513 767
rect 40559 721 40637 767
rect 40683 721 40761 767
rect 40807 721 40885 767
rect 40931 721 41009 767
rect 41055 721 41133 767
rect 41179 721 41257 767
rect 41303 721 41381 767
rect 41427 721 41505 767
rect 41551 721 41629 767
rect 41675 721 41753 767
rect 41799 721 41877 767
rect 41923 721 42001 767
rect 42047 721 42125 767
rect 42171 721 42249 767
rect 42295 721 42373 767
rect 42419 721 42497 767
rect 42543 721 42621 767
rect 42667 721 42745 767
rect 42791 721 42869 767
rect 42915 721 42993 767
rect 43039 721 43117 767
rect 43163 721 43241 767
rect 43287 721 43365 767
rect 43411 721 43489 767
rect 43535 721 43613 767
rect 43659 721 43737 767
rect 43783 721 43861 767
rect 43907 721 43985 767
rect 44031 721 44109 767
rect 44155 721 44233 767
rect 44279 721 44357 767
rect 44403 721 44481 767
rect 44527 721 44605 767
rect 44651 721 44729 767
rect 44775 721 44853 767
rect 44899 721 44977 767
rect 45023 721 45101 767
rect 45147 721 45225 767
rect 45271 721 45349 767
rect 45395 721 45473 767
rect 45519 721 45597 767
rect 45643 721 45721 767
rect 45767 721 45845 767
rect 45891 721 45969 767
rect 46015 721 46093 767
rect 46139 721 46217 767
rect 46263 721 46341 767
rect 46387 721 46465 767
rect 46511 721 46589 767
rect 46635 721 46713 767
rect 46759 721 46837 767
rect 46883 721 46961 767
rect 47007 721 47085 767
rect 47131 721 47209 767
rect 47255 721 47333 767
rect 47379 721 47457 767
rect 47503 721 47581 767
rect 47627 721 47705 767
rect 47751 721 47829 767
rect 47875 721 47953 767
rect 47999 721 48077 767
rect 48123 721 48201 767
rect 48247 721 48325 767
rect 48371 721 48449 767
rect 48495 721 48573 767
rect 48619 721 48697 767
rect 48743 721 48821 767
rect 48867 721 48945 767
rect 48991 721 49069 767
rect 49115 721 49193 767
rect 49239 721 49317 767
rect 49363 721 49441 767
rect 49487 721 49565 767
rect 49611 721 49689 767
rect 49735 721 49813 767
rect 49859 721 49937 767
rect 49983 721 50061 767
rect 50107 721 50185 767
rect 50231 721 50309 767
rect 50355 721 50433 767
rect 50479 721 50557 767
rect 50603 721 50681 767
rect 50727 721 50805 767
rect 50851 721 50929 767
rect 50975 721 51053 767
rect 51099 721 51177 767
rect 51223 721 51301 767
rect 51347 721 51425 767
rect 51471 721 51549 767
rect 51595 721 51673 767
rect 51719 721 51797 767
rect 51843 721 51921 767
rect 51967 721 52045 767
rect 52091 721 52169 767
rect 52215 721 52293 767
rect 52339 721 52417 767
rect 52463 721 52541 767
rect 52587 721 52665 767
rect 52711 721 52789 767
rect 52835 721 52913 767
rect 52959 721 53037 767
rect 53083 721 53161 767
rect 53207 721 53285 767
rect 53331 721 53409 767
rect 53455 721 53533 767
rect 53579 721 53657 767
rect 53703 721 53781 767
rect 53827 721 53905 767
rect 53951 721 54029 767
rect 54075 721 54153 767
rect 54199 721 54277 767
rect 54323 721 54401 767
rect 54447 721 54525 767
rect 54571 721 54649 767
rect 54695 721 54773 767
rect 54819 721 54897 767
rect 54943 721 55021 767
rect 55067 721 55145 767
rect 55191 721 55269 767
rect 55315 721 55393 767
rect 55439 721 55517 767
rect 55563 721 55641 767
rect 55687 721 55765 767
rect 55811 721 55889 767
rect 55935 721 56013 767
rect 56059 721 56137 767
rect 56183 721 56261 767
rect 56307 721 56385 767
rect 56431 721 56509 767
rect 56555 721 56633 767
rect 56679 721 56757 767
rect 56803 721 56881 767
rect 56927 721 57005 767
rect 57051 721 57129 767
rect 57175 721 57253 767
rect 57299 721 57377 767
rect 57423 721 57501 767
rect 57547 721 57625 767
rect 57671 721 57749 767
rect 57795 721 57873 767
rect 57919 721 57997 767
rect 58043 721 58121 767
rect 58167 721 58245 767
rect 58291 721 58369 767
rect 58415 721 58493 767
rect 58539 721 58617 767
rect 58663 721 58741 767
rect 58787 721 58865 767
rect 58911 721 58989 767
rect 59035 721 59113 767
rect 59159 721 59237 767
rect 59283 721 59361 767
rect 59407 721 59485 767
rect 59531 721 59609 767
rect 59655 721 59733 767
rect 59779 721 59857 767
rect 59903 721 59981 767
rect 60027 721 60105 767
rect 60151 721 60229 767
rect 60275 721 60353 767
rect 60399 721 60477 767
rect 60523 721 60601 767
rect 60647 721 60725 767
rect 60771 721 60849 767
rect 60895 721 60973 767
rect 61019 721 61097 767
rect 61143 721 61221 767
rect 61267 721 61345 767
rect 61391 721 61469 767
rect 61515 721 61593 767
rect 61639 721 61717 767
rect 61763 721 61841 767
rect 61887 721 61965 767
rect 62011 721 62089 767
rect 62135 721 62213 767
rect 62259 721 62337 767
rect 62383 721 62461 767
rect 62507 721 62585 767
rect 62631 721 62709 767
rect 62755 721 62833 767
rect 62879 721 62957 767
rect 63003 721 63081 767
rect 63127 721 63205 767
rect 63251 721 63329 767
rect 63375 721 63453 767
rect 63499 721 63577 767
rect 63623 721 63701 767
rect 63747 721 63825 767
rect 63871 721 63949 767
rect 63995 721 64073 767
rect 64119 721 64197 767
rect 64243 721 64321 767
rect 64367 721 64445 767
rect 64491 721 64569 767
rect 64615 721 64693 767
rect 64739 721 64817 767
rect 64863 721 64941 767
rect 64987 721 65065 767
rect 65111 721 65189 767
rect 65235 721 65313 767
rect 65359 721 65437 767
rect 65483 721 65561 767
rect 65607 721 65685 767
rect 65731 721 65809 767
rect 65855 721 65933 767
rect 65979 721 66057 767
rect 66103 721 66181 767
rect 66227 721 66305 767
rect 66351 721 66429 767
rect 66475 721 66553 767
rect 66599 721 66677 767
rect 66723 721 66801 767
rect 66847 721 66925 767
rect 66971 721 67049 767
rect 67095 721 67173 767
rect 67219 721 67297 767
rect 67343 721 67421 767
rect 67467 721 67545 767
rect 67591 721 67669 767
rect 67715 721 67793 767
rect 67839 721 67917 767
rect 67963 721 68041 767
rect 68087 721 68165 767
rect 68211 721 68289 767
rect 68335 721 68413 767
rect 68459 721 68537 767
rect 68583 721 68661 767
rect 68707 721 68785 767
rect 68831 721 68909 767
rect 68955 721 69033 767
rect 69079 721 69157 767
rect 69203 721 69281 767
rect 69327 721 69405 767
rect 69451 721 69529 767
rect 69575 721 69653 767
rect 69699 721 69777 767
rect 69823 721 69901 767
rect 69947 721 70025 767
rect 70071 721 70149 767
rect 70195 721 70273 767
rect 70319 721 70397 767
rect 70443 721 70521 767
rect 70567 721 70645 767
rect 70691 721 70769 767
rect 70815 721 70893 767
rect 70939 721 71017 767
rect 71063 721 71141 767
rect 71187 721 71265 767
rect 71311 721 71389 767
rect 71435 721 71513 767
rect 71559 721 71637 767
rect 71683 721 71761 767
rect 71807 721 71885 767
rect 71931 721 72009 767
rect 72055 721 72133 767
rect 72179 721 72257 767
rect 72303 721 72381 767
rect 72427 721 72505 767
rect 72551 721 72629 767
rect 72675 721 72753 767
rect 72799 721 72877 767
rect 72923 721 73001 767
rect 73047 721 73125 767
rect 73171 721 73249 767
rect 73295 721 73373 767
rect 73419 721 73497 767
rect 73543 721 73621 767
rect 73667 721 73745 767
rect 73791 721 73869 767
rect 73915 721 73993 767
rect 74039 721 74117 767
rect 74163 721 74241 767
rect 74287 721 74365 767
rect 74411 721 74489 767
rect 74535 721 74613 767
rect 74659 721 74737 767
rect 74783 721 74861 767
rect 74907 721 74985 767
rect 75031 721 75109 767
rect 75155 721 75233 767
rect 75279 721 75357 767
rect 75403 721 75481 767
rect 75527 721 75605 767
rect 75651 721 75729 767
rect 75775 721 75853 767
rect 75899 721 75977 767
rect 76023 721 76101 767
rect 76147 721 76225 767
rect 76271 721 76349 767
rect 76395 721 76473 767
rect 76519 721 76597 767
rect 76643 721 76721 767
rect 76767 721 76845 767
rect 76891 721 76969 767
rect 77015 721 77093 767
rect 77139 721 77217 767
rect 77263 721 77341 767
rect 77387 721 77465 767
rect 77511 721 77589 767
rect 77635 721 77713 767
rect 77759 721 77837 767
rect 77883 721 77961 767
rect 78007 721 78085 767
rect 78131 721 78209 767
rect 78255 721 78333 767
rect 78379 721 78457 767
rect 78503 721 78581 767
rect 78627 721 78705 767
rect 78751 721 78829 767
rect 78875 721 78953 767
rect 78999 721 79077 767
rect 79123 721 79201 767
rect 79247 721 79325 767
rect 79371 721 79449 767
rect 79495 721 79573 767
rect 79619 721 79697 767
rect 79743 721 79821 767
rect 79867 721 79945 767
rect 79991 721 80069 767
rect 80115 721 80193 767
rect 80239 721 80317 767
rect 80363 721 80441 767
rect 80487 721 80565 767
rect 80611 721 80689 767
rect 80735 721 80813 767
rect 80859 721 80937 767
rect 80983 721 81061 767
rect 81107 721 81185 767
rect 81231 721 81309 767
rect 81355 721 81433 767
rect 81479 721 81557 767
rect 81603 721 81681 767
rect 81727 721 81805 767
rect 81851 721 81929 767
rect 81975 721 82053 767
rect 82099 721 82177 767
rect 82223 721 82301 767
rect 82347 721 82425 767
rect 82471 721 82549 767
rect 82595 721 82673 767
rect 82719 721 82797 767
rect 82843 721 82921 767
rect 82967 721 83045 767
rect 83091 721 83169 767
rect 83215 721 83293 767
rect 83339 721 83417 767
rect 83463 721 83541 767
rect 83587 721 83665 767
rect 83711 721 83789 767
rect 83835 721 83913 767
rect 83959 721 84037 767
rect 84083 721 84161 767
rect 84207 721 84285 767
rect 84331 721 84409 767
rect 84455 721 84533 767
rect 84579 721 84657 767
rect 84703 721 84781 767
rect 84827 721 84905 767
rect 84951 721 85029 767
rect 85075 721 85153 767
rect 85199 721 85277 767
rect 85323 721 85401 767
rect 85447 721 85525 767
rect 85571 721 85649 767
rect 85695 721 85816 767
rect 70 643 85816 721
rect 70 597 89 643
rect 135 597 213 643
rect 259 597 337 643
rect 383 597 461 643
rect 507 597 585 643
rect 631 597 709 643
rect 755 597 833 643
rect 879 597 957 643
rect 1003 597 1081 643
rect 1127 597 1205 643
rect 1251 597 1329 643
rect 1375 597 1453 643
rect 1499 597 1577 643
rect 1623 597 1701 643
rect 1747 597 1825 643
rect 1871 597 1949 643
rect 1995 597 2073 643
rect 2119 597 2197 643
rect 2243 597 2321 643
rect 2367 597 2445 643
rect 2491 597 2569 643
rect 2615 597 2693 643
rect 2739 597 2817 643
rect 2863 597 2941 643
rect 2987 597 3065 643
rect 3111 597 3189 643
rect 3235 597 3313 643
rect 3359 597 3437 643
rect 3483 597 3561 643
rect 3607 597 3685 643
rect 3731 597 3809 643
rect 3855 597 3933 643
rect 3979 597 4057 643
rect 4103 597 4181 643
rect 4227 597 4305 643
rect 4351 597 4429 643
rect 4475 597 4553 643
rect 4599 597 4677 643
rect 4723 597 4801 643
rect 4847 597 4925 643
rect 4971 597 5049 643
rect 5095 597 5173 643
rect 5219 597 5297 643
rect 5343 597 5421 643
rect 5467 597 5545 643
rect 5591 597 5669 643
rect 5715 597 5793 643
rect 5839 597 5917 643
rect 5963 597 6041 643
rect 6087 597 6165 643
rect 6211 597 6289 643
rect 6335 597 6413 643
rect 6459 597 6537 643
rect 6583 597 6661 643
rect 6707 597 6785 643
rect 6831 597 6909 643
rect 6955 597 7033 643
rect 7079 597 7157 643
rect 7203 597 7281 643
rect 7327 597 7405 643
rect 7451 597 7529 643
rect 7575 597 7653 643
rect 7699 597 7777 643
rect 7823 597 7901 643
rect 7947 597 8025 643
rect 8071 597 8149 643
rect 8195 597 8273 643
rect 8319 597 8397 643
rect 8443 597 8521 643
rect 8567 597 8645 643
rect 8691 597 8769 643
rect 8815 597 8893 643
rect 8939 597 9017 643
rect 9063 597 9141 643
rect 9187 597 9265 643
rect 9311 597 9389 643
rect 9435 597 9513 643
rect 9559 597 9637 643
rect 9683 597 9761 643
rect 9807 597 9885 643
rect 9931 597 10009 643
rect 10055 597 10133 643
rect 10179 597 10257 643
rect 10303 597 10381 643
rect 10427 597 10505 643
rect 10551 597 10629 643
rect 10675 597 10753 643
rect 10799 597 10877 643
rect 10923 597 11001 643
rect 11047 597 11125 643
rect 11171 597 11249 643
rect 11295 597 11373 643
rect 11419 597 11497 643
rect 11543 597 11621 643
rect 11667 597 11745 643
rect 11791 597 11869 643
rect 11915 597 11993 643
rect 12039 597 12117 643
rect 12163 597 12241 643
rect 12287 597 12365 643
rect 12411 597 12489 643
rect 12535 597 12613 643
rect 12659 597 12737 643
rect 12783 597 12861 643
rect 12907 597 12985 643
rect 13031 597 13109 643
rect 13155 597 13233 643
rect 13279 597 13357 643
rect 13403 597 13481 643
rect 13527 597 13605 643
rect 13651 597 13729 643
rect 13775 597 13853 643
rect 13899 597 13977 643
rect 14023 597 14101 643
rect 14147 597 14225 643
rect 14271 597 14349 643
rect 14395 597 14473 643
rect 14519 597 14597 643
rect 14643 597 14721 643
rect 14767 597 14845 643
rect 14891 597 14969 643
rect 15015 597 15093 643
rect 15139 597 15217 643
rect 15263 597 15341 643
rect 15387 597 15465 643
rect 15511 597 15589 643
rect 15635 597 15713 643
rect 15759 597 15837 643
rect 15883 597 15961 643
rect 16007 597 16085 643
rect 16131 597 16209 643
rect 16255 597 16333 643
rect 16379 597 16457 643
rect 16503 597 16581 643
rect 16627 597 16705 643
rect 16751 597 16829 643
rect 16875 597 16953 643
rect 16999 597 17077 643
rect 17123 597 17201 643
rect 17247 597 17325 643
rect 17371 597 17449 643
rect 17495 597 17573 643
rect 17619 597 17697 643
rect 17743 597 17821 643
rect 17867 597 17945 643
rect 17991 597 18069 643
rect 18115 597 18193 643
rect 18239 597 18317 643
rect 18363 597 18441 643
rect 18487 597 18565 643
rect 18611 597 18689 643
rect 18735 597 18813 643
rect 18859 597 18937 643
rect 18983 597 19061 643
rect 19107 597 19185 643
rect 19231 597 19309 643
rect 19355 597 19433 643
rect 19479 597 19557 643
rect 19603 597 19681 643
rect 19727 597 19805 643
rect 19851 597 19929 643
rect 19975 597 20053 643
rect 20099 597 20177 643
rect 20223 597 20301 643
rect 20347 597 20425 643
rect 20471 597 20549 643
rect 20595 597 20673 643
rect 20719 597 20797 643
rect 20843 597 20921 643
rect 20967 597 21045 643
rect 21091 597 21169 643
rect 21215 597 21293 643
rect 21339 597 21417 643
rect 21463 597 21541 643
rect 21587 597 21665 643
rect 21711 597 21789 643
rect 21835 597 21913 643
rect 21959 597 22037 643
rect 22083 597 22161 643
rect 22207 597 22285 643
rect 22331 597 22409 643
rect 22455 597 22533 643
rect 22579 597 22657 643
rect 22703 597 22781 643
rect 22827 597 22905 643
rect 22951 597 23029 643
rect 23075 597 23153 643
rect 23199 597 23277 643
rect 23323 597 23401 643
rect 23447 597 23525 643
rect 23571 597 23649 643
rect 23695 597 23773 643
rect 23819 597 23897 643
rect 23943 597 24021 643
rect 24067 597 24145 643
rect 24191 597 24269 643
rect 24315 597 24393 643
rect 24439 597 24517 643
rect 24563 597 24641 643
rect 24687 597 24765 643
rect 24811 597 24889 643
rect 24935 597 25013 643
rect 25059 597 25137 643
rect 25183 597 25261 643
rect 25307 597 25385 643
rect 25431 597 25509 643
rect 25555 597 25633 643
rect 25679 597 25757 643
rect 25803 597 25881 643
rect 25927 597 26005 643
rect 26051 597 26129 643
rect 26175 597 26253 643
rect 26299 597 26377 643
rect 26423 597 26501 643
rect 26547 597 26625 643
rect 26671 597 26749 643
rect 26795 597 26873 643
rect 26919 597 26997 643
rect 27043 597 27121 643
rect 27167 597 27245 643
rect 27291 597 27369 643
rect 27415 597 27493 643
rect 27539 597 27617 643
rect 27663 597 27741 643
rect 27787 597 27865 643
rect 27911 597 27989 643
rect 28035 597 28113 643
rect 28159 597 28237 643
rect 28283 597 28361 643
rect 28407 597 28485 643
rect 28531 597 28609 643
rect 28655 597 28733 643
rect 28779 597 28857 643
rect 28903 597 28981 643
rect 29027 597 29105 643
rect 29151 597 29229 643
rect 29275 597 29353 643
rect 29399 597 29477 643
rect 29523 597 29601 643
rect 29647 597 29725 643
rect 29771 597 29849 643
rect 29895 597 29973 643
rect 30019 597 30097 643
rect 30143 597 30221 643
rect 30267 597 30345 643
rect 30391 597 30469 643
rect 30515 597 30593 643
rect 30639 597 30717 643
rect 30763 597 30841 643
rect 30887 597 30965 643
rect 31011 597 31089 643
rect 31135 597 31213 643
rect 31259 597 31337 643
rect 31383 597 31461 643
rect 31507 597 31585 643
rect 31631 597 31709 643
rect 31755 597 31833 643
rect 31879 597 31957 643
rect 32003 597 32081 643
rect 32127 597 32205 643
rect 32251 597 32329 643
rect 32375 597 32453 643
rect 32499 597 32577 643
rect 32623 597 32701 643
rect 32747 597 32825 643
rect 32871 597 32949 643
rect 32995 597 33073 643
rect 33119 597 33197 643
rect 33243 597 33321 643
rect 33367 597 33445 643
rect 33491 597 33569 643
rect 33615 597 33693 643
rect 33739 597 33817 643
rect 33863 597 33941 643
rect 33987 597 34065 643
rect 34111 597 34189 643
rect 34235 597 34313 643
rect 34359 597 34437 643
rect 34483 597 34561 643
rect 34607 597 34685 643
rect 34731 597 34809 643
rect 34855 597 34933 643
rect 34979 597 35057 643
rect 35103 597 35181 643
rect 35227 597 35305 643
rect 35351 597 35429 643
rect 35475 597 35553 643
rect 35599 597 35677 643
rect 35723 597 35801 643
rect 35847 597 35925 643
rect 35971 597 36049 643
rect 36095 597 36173 643
rect 36219 597 36297 643
rect 36343 597 36421 643
rect 36467 597 36545 643
rect 36591 597 36669 643
rect 36715 597 36793 643
rect 36839 597 36917 643
rect 36963 597 37041 643
rect 37087 597 37165 643
rect 37211 597 37289 643
rect 37335 597 37413 643
rect 37459 597 37537 643
rect 37583 597 37661 643
rect 37707 597 37785 643
rect 37831 597 37909 643
rect 37955 597 38033 643
rect 38079 597 38157 643
rect 38203 597 38281 643
rect 38327 597 38405 643
rect 38451 597 38529 643
rect 38575 597 38653 643
rect 38699 597 38777 643
rect 38823 597 38901 643
rect 38947 597 39025 643
rect 39071 597 39149 643
rect 39195 597 39273 643
rect 39319 597 39397 643
rect 39443 597 39521 643
rect 39567 597 39645 643
rect 39691 597 39769 643
rect 39815 597 39893 643
rect 39939 597 40017 643
rect 40063 597 40141 643
rect 40187 597 40265 643
rect 40311 597 40389 643
rect 40435 597 40513 643
rect 40559 597 40637 643
rect 40683 597 40761 643
rect 40807 597 40885 643
rect 40931 597 41009 643
rect 41055 597 41133 643
rect 41179 597 41257 643
rect 41303 597 41381 643
rect 41427 597 41505 643
rect 41551 597 41629 643
rect 41675 597 41753 643
rect 41799 597 41877 643
rect 41923 597 42001 643
rect 42047 597 42125 643
rect 42171 597 42249 643
rect 42295 597 42373 643
rect 42419 597 42497 643
rect 42543 597 42621 643
rect 42667 597 42745 643
rect 42791 597 42869 643
rect 42915 597 42993 643
rect 43039 597 43117 643
rect 43163 597 43241 643
rect 43287 597 43365 643
rect 43411 597 43489 643
rect 43535 597 43613 643
rect 43659 597 43737 643
rect 43783 597 43861 643
rect 43907 597 43985 643
rect 44031 597 44109 643
rect 44155 597 44233 643
rect 44279 597 44357 643
rect 44403 597 44481 643
rect 44527 597 44605 643
rect 44651 597 44729 643
rect 44775 597 44853 643
rect 44899 597 44977 643
rect 45023 597 45101 643
rect 45147 597 45225 643
rect 45271 597 45349 643
rect 45395 597 45473 643
rect 45519 597 45597 643
rect 45643 597 45721 643
rect 45767 597 45845 643
rect 45891 597 45969 643
rect 46015 597 46093 643
rect 46139 597 46217 643
rect 46263 597 46341 643
rect 46387 597 46465 643
rect 46511 597 46589 643
rect 46635 597 46713 643
rect 46759 597 46837 643
rect 46883 597 46961 643
rect 47007 597 47085 643
rect 47131 597 47209 643
rect 47255 597 47333 643
rect 47379 597 47457 643
rect 47503 597 47581 643
rect 47627 597 47705 643
rect 47751 597 47829 643
rect 47875 597 47953 643
rect 47999 597 48077 643
rect 48123 597 48201 643
rect 48247 597 48325 643
rect 48371 597 48449 643
rect 48495 597 48573 643
rect 48619 597 48697 643
rect 48743 597 48821 643
rect 48867 597 48945 643
rect 48991 597 49069 643
rect 49115 597 49193 643
rect 49239 597 49317 643
rect 49363 597 49441 643
rect 49487 597 49565 643
rect 49611 597 49689 643
rect 49735 597 49813 643
rect 49859 597 49937 643
rect 49983 597 50061 643
rect 50107 597 50185 643
rect 50231 597 50309 643
rect 50355 597 50433 643
rect 50479 597 50557 643
rect 50603 597 50681 643
rect 50727 597 50805 643
rect 50851 597 50929 643
rect 50975 597 51053 643
rect 51099 597 51177 643
rect 51223 597 51301 643
rect 51347 597 51425 643
rect 51471 597 51549 643
rect 51595 597 51673 643
rect 51719 597 51797 643
rect 51843 597 51921 643
rect 51967 597 52045 643
rect 52091 597 52169 643
rect 52215 597 52293 643
rect 52339 597 52417 643
rect 52463 597 52541 643
rect 52587 597 52665 643
rect 52711 597 52789 643
rect 52835 597 52913 643
rect 52959 597 53037 643
rect 53083 597 53161 643
rect 53207 597 53285 643
rect 53331 597 53409 643
rect 53455 597 53533 643
rect 53579 597 53657 643
rect 53703 597 53781 643
rect 53827 597 53905 643
rect 53951 597 54029 643
rect 54075 597 54153 643
rect 54199 597 54277 643
rect 54323 597 54401 643
rect 54447 597 54525 643
rect 54571 597 54649 643
rect 54695 597 54773 643
rect 54819 597 54897 643
rect 54943 597 55021 643
rect 55067 597 55145 643
rect 55191 597 55269 643
rect 55315 597 55393 643
rect 55439 597 55517 643
rect 55563 597 55641 643
rect 55687 597 55765 643
rect 55811 597 55889 643
rect 55935 597 56013 643
rect 56059 597 56137 643
rect 56183 597 56261 643
rect 56307 597 56385 643
rect 56431 597 56509 643
rect 56555 597 56633 643
rect 56679 597 56757 643
rect 56803 597 56881 643
rect 56927 597 57005 643
rect 57051 597 57129 643
rect 57175 597 57253 643
rect 57299 597 57377 643
rect 57423 597 57501 643
rect 57547 597 57625 643
rect 57671 597 57749 643
rect 57795 597 57873 643
rect 57919 597 57997 643
rect 58043 597 58121 643
rect 58167 597 58245 643
rect 58291 597 58369 643
rect 58415 597 58493 643
rect 58539 597 58617 643
rect 58663 597 58741 643
rect 58787 597 58865 643
rect 58911 597 58989 643
rect 59035 597 59113 643
rect 59159 597 59237 643
rect 59283 597 59361 643
rect 59407 597 59485 643
rect 59531 597 59609 643
rect 59655 597 59733 643
rect 59779 597 59857 643
rect 59903 597 59981 643
rect 60027 597 60105 643
rect 60151 597 60229 643
rect 60275 597 60353 643
rect 60399 597 60477 643
rect 60523 597 60601 643
rect 60647 597 60725 643
rect 60771 597 60849 643
rect 60895 597 60973 643
rect 61019 597 61097 643
rect 61143 597 61221 643
rect 61267 597 61345 643
rect 61391 597 61469 643
rect 61515 597 61593 643
rect 61639 597 61717 643
rect 61763 597 61841 643
rect 61887 597 61965 643
rect 62011 597 62089 643
rect 62135 597 62213 643
rect 62259 597 62337 643
rect 62383 597 62461 643
rect 62507 597 62585 643
rect 62631 597 62709 643
rect 62755 597 62833 643
rect 62879 597 62957 643
rect 63003 597 63081 643
rect 63127 597 63205 643
rect 63251 597 63329 643
rect 63375 597 63453 643
rect 63499 597 63577 643
rect 63623 597 63701 643
rect 63747 597 63825 643
rect 63871 597 63949 643
rect 63995 597 64073 643
rect 64119 597 64197 643
rect 64243 597 64321 643
rect 64367 597 64445 643
rect 64491 597 64569 643
rect 64615 597 64693 643
rect 64739 597 64817 643
rect 64863 597 64941 643
rect 64987 597 65065 643
rect 65111 597 65189 643
rect 65235 597 65313 643
rect 65359 597 65437 643
rect 65483 597 65561 643
rect 65607 597 65685 643
rect 65731 597 65809 643
rect 65855 597 65933 643
rect 65979 597 66057 643
rect 66103 597 66181 643
rect 66227 597 66305 643
rect 66351 597 66429 643
rect 66475 597 66553 643
rect 66599 597 66677 643
rect 66723 597 66801 643
rect 66847 597 66925 643
rect 66971 597 67049 643
rect 67095 597 67173 643
rect 67219 597 67297 643
rect 67343 597 67421 643
rect 67467 597 67545 643
rect 67591 597 67669 643
rect 67715 597 67793 643
rect 67839 597 67917 643
rect 67963 597 68041 643
rect 68087 597 68165 643
rect 68211 597 68289 643
rect 68335 597 68413 643
rect 68459 597 68537 643
rect 68583 597 68661 643
rect 68707 597 68785 643
rect 68831 597 68909 643
rect 68955 597 69033 643
rect 69079 597 69157 643
rect 69203 597 69281 643
rect 69327 597 69405 643
rect 69451 597 69529 643
rect 69575 597 69653 643
rect 69699 597 69777 643
rect 69823 597 69901 643
rect 69947 597 70025 643
rect 70071 597 70149 643
rect 70195 597 70273 643
rect 70319 597 70397 643
rect 70443 597 70521 643
rect 70567 597 70645 643
rect 70691 597 70769 643
rect 70815 597 70893 643
rect 70939 597 71017 643
rect 71063 597 71141 643
rect 71187 597 71265 643
rect 71311 597 71389 643
rect 71435 597 71513 643
rect 71559 597 71637 643
rect 71683 597 71761 643
rect 71807 597 71885 643
rect 71931 597 72009 643
rect 72055 597 72133 643
rect 72179 597 72257 643
rect 72303 597 72381 643
rect 72427 597 72505 643
rect 72551 597 72629 643
rect 72675 597 72753 643
rect 72799 597 72877 643
rect 72923 597 73001 643
rect 73047 597 73125 643
rect 73171 597 73249 643
rect 73295 597 73373 643
rect 73419 597 73497 643
rect 73543 597 73621 643
rect 73667 597 73745 643
rect 73791 597 73869 643
rect 73915 597 73993 643
rect 74039 597 74117 643
rect 74163 597 74241 643
rect 74287 597 74365 643
rect 74411 597 74489 643
rect 74535 597 74613 643
rect 74659 597 74737 643
rect 74783 597 74861 643
rect 74907 597 74985 643
rect 75031 597 75109 643
rect 75155 597 75233 643
rect 75279 597 75357 643
rect 75403 597 75481 643
rect 75527 597 75605 643
rect 75651 597 75729 643
rect 75775 597 75853 643
rect 75899 597 75977 643
rect 76023 597 76101 643
rect 76147 597 76225 643
rect 76271 597 76349 643
rect 76395 597 76473 643
rect 76519 597 76597 643
rect 76643 597 76721 643
rect 76767 597 76845 643
rect 76891 597 76969 643
rect 77015 597 77093 643
rect 77139 597 77217 643
rect 77263 597 77341 643
rect 77387 597 77465 643
rect 77511 597 77589 643
rect 77635 597 77713 643
rect 77759 597 77837 643
rect 77883 597 77961 643
rect 78007 597 78085 643
rect 78131 597 78209 643
rect 78255 597 78333 643
rect 78379 597 78457 643
rect 78503 597 78581 643
rect 78627 597 78705 643
rect 78751 597 78829 643
rect 78875 597 78953 643
rect 78999 597 79077 643
rect 79123 597 79201 643
rect 79247 597 79325 643
rect 79371 597 79449 643
rect 79495 597 79573 643
rect 79619 597 79697 643
rect 79743 597 79821 643
rect 79867 597 79945 643
rect 79991 597 80069 643
rect 80115 597 80193 643
rect 80239 597 80317 643
rect 80363 597 80441 643
rect 80487 597 80565 643
rect 80611 597 80689 643
rect 80735 597 80813 643
rect 80859 597 80937 643
rect 80983 597 81061 643
rect 81107 597 81185 643
rect 81231 597 81309 643
rect 81355 597 81433 643
rect 81479 597 81557 643
rect 81603 597 81681 643
rect 81727 597 81805 643
rect 81851 597 81929 643
rect 81975 597 82053 643
rect 82099 597 82177 643
rect 82223 597 82301 643
rect 82347 597 82425 643
rect 82471 597 82549 643
rect 82595 597 82673 643
rect 82719 597 82797 643
rect 82843 597 82921 643
rect 82967 597 83045 643
rect 83091 597 83169 643
rect 83215 597 83293 643
rect 83339 597 83417 643
rect 83463 597 83541 643
rect 83587 597 83665 643
rect 83711 597 83789 643
rect 83835 597 83913 643
rect 83959 597 84037 643
rect 84083 597 84161 643
rect 84207 597 84285 643
rect 84331 597 84409 643
rect 84455 597 84533 643
rect 84579 597 84657 643
rect 84703 597 84781 643
rect 84827 597 84905 643
rect 84951 597 85029 643
rect 85075 597 85153 643
rect 85199 597 85277 643
rect 85323 597 85401 643
rect 85447 597 85525 643
rect 85571 597 85649 643
rect 85695 597 85816 643
rect 70 578 85816 597
<< psubdiffcont >>
rect 89 46037 135 46083
rect 213 46037 259 46083
rect 337 46037 383 46083
rect 461 46037 507 46083
rect 585 46037 631 46083
rect 709 46037 755 46083
rect 833 46037 879 46083
rect 957 46037 1003 46083
rect 1081 46037 1127 46083
rect 1205 46037 1251 46083
rect 1329 46037 1375 46083
rect 1453 46037 1499 46083
rect 1577 46037 1623 46083
rect 1701 46037 1747 46083
rect 1825 46037 1871 46083
rect 1949 46037 1995 46083
rect 2073 46037 2119 46083
rect 2197 46037 2243 46083
rect 2321 46037 2367 46083
rect 2445 46037 2491 46083
rect 2569 46037 2615 46083
rect 2693 46037 2739 46083
rect 2817 46037 2863 46083
rect 2941 46037 2987 46083
rect 3065 46037 3111 46083
rect 3189 46037 3235 46083
rect 3313 46037 3359 46083
rect 3437 46037 3483 46083
rect 3561 46037 3607 46083
rect 3685 46037 3731 46083
rect 3809 46037 3855 46083
rect 3933 46037 3979 46083
rect 4057 46037 4103 46083
rect 4181 46037 4227 46083
rect 4305 46037 4351 46083
rect 4429 46037 4475 46083
rect 4553 46037 4599 46083
rect 4677 46037 4723 46083
rect 4801 46037 4847 46083
rect 4925 46037 4971 46083
rect 5049 46037 5095 46083
rect 5173 46037 5219 46083
rect 5297 46037 5343 46083
rect 5421 46037 5467 46083
rect 5545 46037 5591 46083
rect 5669 46037 5715 46083
rect 5793 46037 5839 46083
rect 5917 46037 5963 46083
rect 6041 46037 6087 46083
rect 6165 46037 6211 46083
rect 6289 46037 6335 46083
rect 6413 46037 6459 46083
rect 6537 46037 6583 46083
rect 6661 46037 6707 46083
rect 6785 46037 6831 46083
rect 6909 46037 6955 46083
rect 7033 46037 7079 46083
rect 7157 46037 7203 46083
rect 7281 46037 7327 46083
rect 7405 46037 7451 46083
rect 7529 46037 7575 46083
rect 7653 46037 7699 46083
rect 7777 46037 7823 46083
rect 7901 46037 7947 46083
rect 8025 46037 8071 46083
rect 8149 46037 8195 46083
rect 8273 46037 8319 46083
rect 8397 46037 8443 46083
rect 8521 46037 8567 46083
rect 8645 46037 8691 46083
rect 8769 46037 8815 46083
rect 8893 46037 8939 46083
rect 9017 46037 9063 46083
rect 9141 46037 9187 46083
rect 9265 46037 9311 46083
rect 9389 46037 9435 46083
rect 9513 46037 9559 46083
rect 9637 46037 9683 46083
rect 9761 46037 9807 46083
rect 9885 46037 9931 46083
rect 10009 46037 10055 46083
rect 10133 46037 10179 46083
rect 10257 46037 10303 46083
rect 10381 46037 10427 46083
rect 10505 46037 10551 46083
rect 10629 46037 10675 46083
rect 10753 46037 10799 46083
rect 10877 46037 10923 46083
rect 11001 46037 11047 46083
rect 11125 46037 11171 46083
rect 11249 46037 11295 46083
rect 11373 46037 11419 46083
rect 11497 46037 11543 46083
rect 11621 46037 11667 46083
rect 11745 46037 11791 46083
rect 11869 46037 11915 46083
rect 11993 46037 12039 46083
rect 12117 46037 12163 46083
rect 12241 46037 12287 46083
rect 12365 46037 12411 46083
rect 12489 46037 12535 46083
rect 12613 46037 12659 46083
rect 12737 46037 12783 46083
rect 12861 46037 12907 46083
rect 12985 46037 13031 46083
rect 13109 46037 13155 46083
rect 13233 46037 13279 46083
rect 13357 46037 13403 46083
rect 13481 46037 13527 46083
rect 13605 46037 13651 46083
rect 13729 46037 13775 46083
rect 13853 46037 13899 46083
rect 13977 46037 14023 46083
rect 14101 46037 14147 46083
rect 14225 46037 14271 46083
rect 14349 46037 14395 46083
rect 14473 46037 14519 46083
rect 14597 46037 14643 46083
rect 14721 46037 14767 46083
rect 14845 46037 14891 46083
rect 14969 46037 15015 46083
rect 15093 46037 15139 46083
rect 15217 46037 15263 46083
rect 15341 46037 15387 46083
rect 15465 46037 15511 46083
rect 15589 46037 15635 46083
rect 15713 46037 15759 46083
rect 15837 46037 15883 46083
rect 15961 46037 16007 46083
rect 16085 46037 16131 46083
rect 16209 46037 16255 46083
rect 16333 46037 16379 46083
rect 16457 46037 16503 46083
rect 16581 46037 16627 46083
rect 16705 46037 16751 46083
rect 16829 46037 16875 46083
rect 16953 46037 16999 46083
rect 17077 46037 17123 46083
rect 17201 46037 17247 46083
rect 17325 46037 17371 46083
rect 17449 46037 17495 46083
rect 17573 46037 17619 46083
rect 17697 46037 17743 46083
rect 17821 46037 17867 46083
rect 17945 46037 17991 46083
rect 18069 46037 18115 46083
rect 18193 46037 18239 46083
rect 18317 46037 18363 46083
rect 18441 46037 18487 46083
rect 18565 46037 18611 46083
rect 18689 46037 18735 46083
rect 18813 46037 18859 46083
rect 18937 46037 18983 46083
rect 19061 46037 19107 46083
rect 19185 46037 19231 46083
rect 19309 46037 19355 46083
rect 19433 46037 19479 46083
rect 19557 46037 19603 46083
rect 19681 46037 19727 46083
rect 19805 46037 19851 46083
rect 19929 46037 19975 46083
rect 20053 46037 20099 46083
rect 20177 46037 20223 46083
rect 20301 46037 20347 46083
rect 20425 46037 20471 46083
rect 20549 46037 20595 46083
rect 20673 46037 20719 46083
rect 20797 46037 20843 46083
rect 20921 46037 20967 46083
rect 21045 46037 21091 46083
rect 21169 46037 21215 46083
rect 21293 46037 21339 46083
rect 21417 46037 21463 46083
rect 21541 46037 21587 46083
rect 21665 46037 21711 46083
rect 21789 46037 21835 46083
rect 21913 46037 21959 46083
rect 22037 46037 22083 46083
rect 22161 46037 22207 46083
rect 22285 46037 22331 46083
rect 22409 46037 22455 46083
rect 22533 46037 22579 46083
rect 22657 46037 22703 46083
rect 22781 46037 22827 46083
rect 22905 46037 22951 46083
rect 23029 46037 23075 46083
rect 23153 46037 23199 46083
rect 23277 46037 23323 46083
rect 23401 46037 23447 46083
rect 23525 46037 23571 46083
rect 23649 46037 23695 46083
rect 23773 46037 23819 46083
rect 23897 46037 23943 46083
rect 24021 46037 24067 46083
rect 24145 46037 24191 46083
rect 24269 46037 24315 46083
rect 24393 46037 24439 46083
rect 24517 46037 24563 46083
rect 24641 46037 24687 46083
rect 24765 46037 24811 46083
rect 24889 46037 24935 46083
rect 25013 46037 25059 46083
rect 25137 46037 25183 46083
rect 25261 46037 25307 46083
rect 25385 46037 25431 46083
rect 25509 46037 25555 46083
rect 25633 46037 25679 46083
rect 25757 46037 25803 46083
rect 25881 46037 25927 46083
rect 26005 46037 26051 46083
rect 26129 46037 26175 46083
rect 26253 46037 26299 46083
rect 26377 46037 26423 46083
rect 26501 46037 26547 46083
rect 26625 46037 26671 46083
rect 26749 46037 26795 46083
rect 26873 46037 26919 46083
rect 26997 46037 27043 46083
rect 27121 46037 27167 46083
rect 27245 46037 27291 46083
rect 27369 46037 27415 46083
rect 27493 46037 27539 46083
rect 27617 46037 27663 46083
rect 27741 46037 27787 46083
rect 27865 46037 27911 46083
rect 27989 46037 28035 46083
rect 28113 46037 28159 46083
rect 28237 46037 28283 46083
rect 28361 46037 28407 46083
rect 28485 46037 28531 46083
rect 28609 46037 28655 46083
rect 28733 46037 28779 46083
rect 28857 46037 28903 46083
rect 28981 46037 29027 46083
rect 29105 46037 29151 46083
rect 29229 46037 29275 46083
rect 29353 46037 29399 46083
rect 29477 46037 29523 46083
rect 29601 46037 29647 46083
rect 29725 46037 29771 46083
rect 29849 46037 29895 46083
rect 29973 46037 30019 46083
rect 30097 46037 30143 46083
rect 30221 46037 30267 46083
rect 30345 46037 30391 46083
rect 30469 46037 30515 46083
rect 30593 46037 30639 46083
rect 30717 46037 30763 46083
rect 30841 46037 30887 46083
rect 30965 46037 31011 46083
rect 31089 46037 31135 46083
rect 31213 46037 31259 46083
rect 31337 46037 31383 46083
rect 31461 46037 31507 46083
rect 31585 46037 31631 46083
rect 31709 46037 31755 46083
rect 31833 46037 31879 46083
rect 31957 46037 32003 46083
rect 32081 46037 32127 46083
rect 32205 46037 32251 46083
rect 32329 46037 32375 46083
rect 32453 46037 32499 46083
rect 32577 46037 32623 46083
rect 32701 46037 32747 46083
rect 32825 46037 32871 46083
rect 32949 46037 32995 46083
rect 33073 46037 33119 46083
rect 33197 46037 33243 46083
rect 33321 46037 33367 46083
rect 33445 46037 33491 46083
rect 33569 46037 33615 46083
rect 33693 46037 33739 46083
rect 33817 46037 33863 46083
rect 33941 46037 33987 46083
rect 34065 46037 34111 46083
rect 34189 46037 34235 46083
rect 34313 46037 34359 46083
rect 34437 46037 34483 46083
rect 34561 46037 34607 46083
rect 34685 46037 34731 46083
rect 34809 46037 34855 46083
rect 34933 46037 34979 46083
rect 35057 46037 35103 46083
rect 35181 46037 35227 46083
rect 35305 46037 35351 46083
rect 35429 46037 35475 46083
rect 35553 46037 35599 46083
rect 35677 46037 35723 46083
rect 35801 46037 35847 46083
rect 35925 46037 35971 46083
rect 36049 46037 36095 46083
rect 36173 46037 36219 46083
rect 36297 46037 36343 46083
rect 36421 46037 36467 46083
rect 36545 46037 36591 46083
rect 36669 46037 36715 46083
rect 36793 46037 36839 46083
rect 36917 46037 36963 46083
rect 37041 46037 37087 46083
rect 37165 46037 37211 46083
rect 37289 46037 37335 46083
rect 37413 46037 37459 46083
rect 37537 46037 37583 46083
rect 37661 46037 37707 46083
rect 37785 46037 37831 46083
rect 37909 46037 37955 46083
rect 38033 46037 38079 46083
rect 38157 46037 38203 46083
rect 38281 46037 38327 46083
rect 38405 46037 38451 46083
rect 38529 46037 38575 46083
rect 38653 46037 38699 46083
rect 38777 46037 38823 46083
rect 38901 46037 38947 46083
rect 39025 46037 39071 46083
rect 39149 46037 39195 46083
rect 39273 46037 39319 46083
rect 39397 46037 39443 46083
rect 39521 46037 39567 46083
rect 39645 46037 39691 46083
rect 39769 46037 39815 46083
rect 39893 46037 39939 46083
rect 40017 46037 40063 46083
rect 40141 46037 40187 46083
rect 40265 46037 40311 46083
rect 40389 46037 40435 46083
rect 40513 46037 40559 46083
rect 40637 46037 40683 46083
rect 40761 46037 40807 46083
rect 40885 46037 40931 46083
rect 41009 46037 41055 46083
rect 41133 46037 41179 46083
rect 41257 46037 41303 46083
rect 41381 46037 41427 46083
rect 41505 46037 41551 46083
rect 41629 46037 41675 46083
rect 41753 46037 41799 46083
rect 41877 46037 41923 46083
rect 42001 46037 42047 46083
rect 42125 46037 42171 46083
rect 42249 46037 42295 46083
rect 42373 46037 42419 46083
rect 42497 46037 42543 46083
rect 42621 46037 42667 46083
rect 42745 46037 42791 46083
rect 42869 46037 42915 46083
rect 42993 46037 43039 46083
rect 43117 46037 43163 46083
rect 43241 46037 43287 46083
rect 43365 46037 43411 46083
rect 43489 46037 43535 46083
rect 43613 46037 43659 46083
rect 43737 46037 43783 46083
rect 43861 46037 43907 46083
rect 43985 46037 44031 46083
rect 44109 46037 44155 46083
rect 44233 46037 44279 46083
rect 44357 46037 44403 46083
rect 44481 46037 44527 46083
rect 44605 46037 44651 46083
rect 44729 46037 44775 46083
rect 44853 46037 44899 46083
rect 44977 46037 45023 46083
rect 45101 46037 45147 46083
rect 45225 46037 45271 46083
rect 45349 46037 45395 46083
rect 45473 46037 45519 46083
rect 45597 46037 45643 46083
rect 45721 46037 45767 46083
rect 45845 46037 45891 46083
rect 45969 46037 46015 46083
rect 46093 46037 46139 46083
rect 46217 46037 46263 46083
rect 46341 46037 46387 46083
rect 46465 46037 46511 46083
rect 46589 46037 46635 46083
rect 46713 46037 46759 46083
rect 46837 46037 46883 46083
rect 46961 46037 47007 46083
rect 47085 46037 47131 46083
rect 47209 46037 47255 46083
rect 47333 46037 47379 46083
rect 47457 46037 47503 46083
rect 47581 46037 47627 46083
rect 47705 46037 47751 46083
rect 47829 46037 47875 46083
rect 47953 46037 47999 46083
rect 48077 46037 48123 46083
rect 48201 46037 48247 46083
rect 48325 46037 48371 46083
rect 48449 46037 48495 46083
rect 48573 46037 48619 46083
rect 48697 46037 48743 46083
rect 48821 46037 48867 46083
rect 48945 46037 48991 46083
rect 49069 46037 49115 46083
rect 49193 46037 49239 46083
rect 49317 46037 49363 46083
rect 49441 46037 49487 46083
rect 49565 46037 49611 46083
rect 49689 46037 49735 46083
rect 49813 46037 49859 46083
rect 49937 46037 49983 46083
rect 50061 46037 50107 46083
rect 50185 46037 50231 46083
rect 50309 46037 50355 46083
rect 50433 46037 50479 46083
rect 50557 46037 50603 46083
rect 50681 46037 50727 46083
rect 50805 46037 50851 46083
rect 50929 46037 50975 46083
rect 51053 46037 51099 46083
rect 51177 46037 51223 46083
rect 51301 46037 51347 46083
rect 51425 46037 51471 46083
rect 51549 46037 51595 46083
rect 51673 46037 51719 46083
rect 51797 46037 51843 46083
rect 51921 46037 51967 46083
rect 52045 46037 52091 46083
rect 52169 46037 52215 46083
rect 52293 46037 52339 46083
rect 52417 46037 52463 46083
rect 52541 46037 52587 46083
rect 52665 46037 52711 46083
rect 52789 46037 52835 46083
rect 52913 46037 52959 46083
rect 53037 46037 53083 46083
rect 53161 46037 53207 46083
rect 53285 46037 53331 46083
rect 53409 46037 53455 46083
rect 53533 46037 53579 46083
rect 53657 46037 53703 46083
rect 53781 46037 53827 46083
rect 53905 46037 53951 46083
rect 54029 46037 54075 46083
rect 54153 46037 54199 46083
rect 54277 46037 54323 46083
rect 54401 46037 54447 46083
rect 54525 46037 54571 46083
rect 54649 46037 54695 46083
rect 54773 46037 54819 46083
rect 54897 46037 54943 46083
rect 55021 46037 55067 46083
rect 55145 46037 55191 46083
rect 55269 46037 55315 46083
rect 55393 46037 55439 46083
rect 55517 46037 55563 46083
rect 55641 46037 55687 46083
rect 55765 46037 55811 46083
rect 55889 46037 55935 46083
rect 56013 46037 56059 46083
rect 56137 46037 56183 46083
rect 56261 46037 56307 46083
rect 56385 46037 56431 46083
rect 56509 46037 56555 46083
rect 56633 46037 56679 46083
rect 56757 46037 56803 46083
rect 56881 46037 56927 46083
rect 57005 46037 57051 46083
rect 57129 46037 57175 46083
rect 57253 46037 57299 46083
rect 57377 46037 57423 46083
rect 57501 46037 57547 46083
rect 57625 46037 57671 46083
rect 57749 46037 57795 46083
rect 57873 46037 57919 46083
rect 57997 46037 58043 46083
rect 58121 46037 58167 46083
rect 58245 46037 58291 46083
rect 58369 46037 58415 46083
rect 58493 46037 58539 46083
rect 58617 46037 58663 46083
rect 58741 46037 58787 46083
rect 58865 46037 58911 46083
rect 58989 46037 59035 46083
rect 59113 46037 59159 46083
rect 59237 46037 59283 46083
rect 59361 46037 59407 46083
rect 59485 46037 59531 46083
rect 59609 46037 59655 46083
rect 59733 46037 59779 46083
rect 59857 46037 59903 46083
rect 59981 46037 60027 46083
rect 60105 46037 60151 46083
rect 60229 46037 60275 46083
rect 60353 46037 60399 46083
rect 60477 46037 60523 46083
rect 60601 46037 60647 46083
rect 60725 46037 60771 46083
rect 60849 46037 60895 46083
rect 60973 46037 61019 46083
rect 61097 46037 61143 46083
rect 61221 46037 61267 46083
rect 61345 46037 61391 46083
rect 61469 46037 61515 46083
rect 61593 46037 61639 46083
rect 61717 46037 61763 46083
rect 61841 46037 61887 46083
rect 61965 46037 62011 46083
rect 62089 46037 62135 46083
rect 62213 46037 62259 46083
rect 62337 46037 62383 46083
rect 62461 46037 62507 46083
rect 62585 46037 62631 46083
rect 62709 46037 62755 46083
rect 62833 46037 62879 46083
rect 62957 46037 63003 46083
rect 63081 46037 63127 46083
rect 63205 46037 63251 46083
rect 63329 46037 63375 46083
rect 63453 46037 63499 46083
rect 63577 46037 63623 46083
rect 63701 46037 63747 46083
rect 63825 46037 63871 46083
rect 63949 46037 63995 46083
rect 64073 46037 64119 46083
rect 64197 46037 64243 46083
rect 64321 46037 64367 46083
rect 64445 46037 64491 46083
rect 64569 46037 64615 46083
rect 64693 46037 64739 46083
rect 64817 46037 64863 46083
rect 64941 46037 64987 46083
rect 65065 46037 65111 46083
rect 65189 46037 65235 46083
rect 65313 46037 65359 46083
rect 65437 46037 65483 46083
rect 65561 46037 65607 46083
rect 65685 46037 65731 46083
rect 65809 46037 65855 46083
rect 65933 46037 65979 46083
rect 66057 46037 66103 46083
rect 66181 46037 66227 46083
rect 66305 46037 66351 46083
rect 66429 46037 66475 46083
rect 66553 46037 66599 46083
rect 66677 46037 66723 46083
rect 66801 46037 66847 46083
rect 66925 46037 66971 46083
rect 67049 46037 67095 46083
rect 67173 46037 67219 46083
rect 67297 46037 67343 46083
rect 67421 46037 67467 46083
rect 67545 46037 67591 46083
rect 67669 46037 67715 46083
rect 67793 46037 67839 46083
rect 67917 46037 67963 46083
rect 68041 46037 68087 46083
rect 68165 46037 68211 46083
rect 68289 46037 68335 46083
rect 68413 46037 68459 46083
rect 68537 46037 68583 46083
rect 68661 46037 68707 46083
rect 68785 46037 68831 46083
rect 68909 46037 68955 46083
rect 69033 46037 69079 46083
rect 69157 46037 69203 46083
rect 69281 46037 69327 46083
rect 69405 46037 69451 46083
rect 69529 46037 69575 46083
rect 69653 46037 69699 46083
rect 69777 46037 69823 46083
rect 69901 46037 69947 46083
rect 70025 46037 70071 46083
rect 70149 46037 70195 46083
rect 70273 46037 70319 46083
rect 70397 46037 70443 46083
rect 70521 46037 70567 46083
rect 70645 46037 70691 46083
rect 70769 46037 70815 46083
rect 70893 46037 70939 46083
rect 71017 46037 71063 46083
rect 71141 46037 71187 46083
rect 71265 46037 71311 46083
rect 71389 46037 71435 46083
rect 71513 46037 71559 46083
rect 71637 46037 71683 46083
rect 71761 46037 71807 46083
rect 71885 46037 71931 46083
rect 72009 46037 72055 46083
rect 72133 46037 72179 46083
rect 72257 46037 72303 46083
rect 72381 46037 72427 46083
rect 72505 46037 72551 46083
rect 72629 46037 72675 46083
rect 72753 46037 72799 46083
rect 72877 46037 72923 46083
rect 73001 46037 73047 46083
rect 73125 46037 73171 46083
rect 73249 46037 73295 46083
rect 73373 46037 73419 46083
rect 73497 46037 73543 46083
rect 73621 46037 73667 46083
rect 73745 46037 73791 46083
rect 73869 46037 73915 46083
rect 73993 46037 74039 46083
rect 74117 46037 74163 46083
rect 74241 46037 74287 46083
rect 74365 46037 74411 46083
rect 74489 46037 74535 46083
rect 74613 46037 74659 46083
rect 74737 46037 74783 46083
rect 74861 46037 74907 46083
rect 74985 46037 75031 46083
rect 75109 46037 75155 46083
rect 75233 46037 75279 46083
rect 75357 46037 75403 46083
rect 75481 46037 75527 46083
rect 75605 46037 75651 46083
rect 75729 46037 75775 46083
rect 75853 46037 75899 46083
rect 75977 46037 76023 46083
rect 76101 46037 76147 46083
rect 76225 46037 76271 46083
rect 76349 46037 76395 46083
rect 76473 46037 76519 46083
rect 76597 46037 76643 46083
rect 76721 46037 76767 46083
rect 76845 46037 76891 46083
rect 76969 46037 77015 46083
rect 77093 46037 77139 46083
rect 77217 46037 77263 46083
rect 77341 46037 77387 46083
rect 77465 46037 77511 46083
rect 77589 46037 77635 46083
rect 77713 46037 77759 46083
rect 77837 46037 77883 46083
rect 77961 46037 78007 46083
rect 78085 46037 78131 46083
rect 78209 46037 78255 46083
rect 78333 46037 78379 46083
rect 78457 46037 78503 46083
rect 78581 46037 78627 46083
rect 78705 46037 78751 46083
rect 78829 46037 78875 46083
rect 78953 46037 78999 46083
rect 79077 46037 79123 46083
rect 79201 46037 79247 46083
rect 79325 46037 79371 46083
rect 79449 46037 79495 46083
rect 79573 46037 79619 46083
rect 79697 46037 79743 46083
rect 79821 46037 79867 46083
rect 79945 46037 79991 46083
rect 80069 46037 80115 46083
rect 80193 46037 80239 46083
rect 80317 46037 80363 46083
rect 80441 46037 80487 46083
rect 80565 46037 80611 46083
rect 80689 46037 80735 46083
rect 80813 46037 80859 46083
rect 80937 46037 80983 46083
rect 81061 46037 81107 46083
rect 81185 46037 81231 46083
rect 81309 46037 81355 46083
rect 81433 46037 81479 46083
rect 81557 46037 81603 46083
rect 81681 46037 81727 46083
rect 81805 46037 81851 46083
rect 81929 46037 81975 46083
rect 82053 46037 82099 46083
rect 82177 46037 82223 46083
rect 82301 46037 82347 46083
rect 82425 46037 82471 46083
rect 82549 46037 82595 46083
rect 82673 46037 82719 46083
rect 82797 46037 82843 46083
rect 82921 46037 82967 46083
rect 83045 46037 83091 46083
rect 83169 46037 83215 46083
rect 83293 46037 83339 46083
rect 83417 46037 83463 46083
rect 83541 46037 83587 46083
rect 83665 46037 83711 46083
rect 83789 46037 83835 46083
rect 83913 46037 83959 46083
rect 84037 46037 84083 46083
rect 84161 46037 84207 46083
rect 84285 46037 84331 46083
rect 84409 46037 84455 46083
rect 84533 46037 84579 46083
rect 84657 46037 84703 46083
rect 84781 46037 84827 46083
rect 84905 46037 84951 46083
rect 85029 46037 85075 46083
rect 85153 46037 85199 46083
rect 85277 46037 85323 46083
rect 85401 46037 85447 46083
rect 85525 46037 85571 46083
rect 85649 46037 85695 46083
rect 89 45913 135 45959
rect 213 45913 259 45959
rect 337 45913 383 45959
rect 461 45913 507 45959
rect 585 45913 631 45959
rect 709 45913 755 45959
rect 833 45913 879 45959
rect 957 45913 1003 45959
rect 1081 45913 1127 45959
rect 1205 45913 1251 45959
rect 1329 45913 1375 45959
rect 1453 45913 1499 45959
rect 1577 45913 1623 45959
rect 1701 45913 1747 45959
rect 1825 45913 1871 45959
rect 1949 45913 1995 45959
rect 2073 45913 2119 45959
rect 2197 45913 2243 45959
rect 2321 45913 2367 45959
rect 2445 45913 2491 45959
rect 2569 45913 2615 45959
rect 2693 45913 2739 45959
rect 2817 45913 2863 45959
rect 2941 45913 2987 45959
rect 3065 45913 3111 45959
rect 3189 45913 3235 45959
rect 3313 45913 3359 45959
rect 3437 45913 3483 45959
rect 3561 45913 3607 45959
rect 3685 45913 3731 45959
rect 3809 45913 3855 45959
rect 3933 45913 3979 45959
rect 4057 45913 4103 45959
rect 4181 45913 4227 45959
rect 4305 45913 4351 45959
rect 4429 45913 4475 45959
rect 4553 45913 4599 45959
rect 4677 45913 4723 45959
rect 4801 45913 4847 45959
rect 4925 45913 4971 45959
rect 5049 45913 5095 45959
rect 5173 45913 5219 45959
rect 5297 45913 5343 45959
rect 5421 45913 5467 45959
rect 5545 45913 5591 45959
rect 5669 45913 5715 45959
rect 5793 45913 5839 45959
rect 5917 45913 5963 45959
rect 6041 45913 6087 45959
rect 6165 45913 6211 45959
rect 6289 45913 6335 45959
rect 6413 45913 6459 45959
rect 6537 45913 6583 45959
rect 6661 45913 6707 45959
rect 6785 45913 6831 45959
rect 6909 45913 6955 45959
rect 7033 45913 7079 45959
rect 7157 45913 7203 45959
rect 7281 45913 7327 45959
rect 7405 45913 7451 45959
rect 7529 45913 7575 45959
rect 7653 45913 7699 45959
rect 7777 45913 7823 45959
rect 7901 45913 7947 45959
rect 8025 45913 8071 45959
rect 8149 45913 8195 45959
rect 8273 45913 8319 45959
rect 8397 45913 8443 45959
rect 8521 45913 8567 45959
rect 8645 45913 8691 45959
rect 8769 45913 8815 45959
rect 8893 45913 8939 45959
rect 9017 45913 9063 45959
rect 9141 45913 9187 45959
rect 9265 45913 9311 45959
rect 9389 45913 9435 45959
rect 9513 45913 9559 45959
rect 9637 45913 9683 45959
rect 9761 45913 9807 45959
rect 9885 45913 9931 45959
rect 10009 45913 10055 45959
rect 10133 45913 10179 45959
rect 10257 45913 10303 45959
rect 10381 45913 10427 45959
rect 10505 45913 10551 45959
rect 10629 45913 10675 45959
rect 10753 45913 10799 45959
rect 10877 45913 10923 45959
rect 11001 45913 11047 45959
rect 11125 45913 11171 45959
rect 11249 45913 11295 45959
rect 11373 45913 11419 45959
rect 11497 45913 11543 45959
rect 11621 45913 11667 45959
rect 11745 45913 11791 45959
rect 11869 45913 11915 45959
rect 11993 45913 12039 45959
rect 12117 45913 12163 45959
rect 12241 45913 12287 45959
rect 12365 45913 12411 45959
rect 12489 45913 12535 45959
rect 12613 45913 12659 45959
rect 12737 45913 12783 45959
rect 12861 45913 12907 45959
rect 12985 45913 13031 45959
rect 13109 45913 13155 45959
rect 13233 45913 13279 45959
rect 13357 45913 13403 45959
rect 13481 45913 13527 45959
rect 13605 45913 13651 45959
rect 13729 45913 13775 45959
rect 13853 45913 13899 45959
rect 13977 45913 14023 45959
rect 14101 45913 14147 45959
rect 14225 45913 14271 45959
rect 14349 45913 14395 45959
rect 14473 45913 14519 45959
rect 14597 45913 14643 45959
rect 14721 45913 14767 45959
rect 14845 45913 14891 45959
rect 14969 45913 15015 45959
rect 15093 45913 15139 45959
rect 15217 45913 15263 45959
rect 15341 45913 15387 45959
rect 15465 45913 15511 45959
rect 15589 45913 15635 45959
rect 15713 45913 15759 45959
rect 15837 45913 15883 45959
rect 15961 45913 16007 45959
rect 16085 45913 16131 45959
rect 16209 45913 16255 45959
rect 16333 45913 16379 45959
rect 16457 45913 16503 45959
rect 16581 45913 16627 45959
rect 16705 45913 16751 45959
rect 16829 45913 16875 45959
rect 16953 45913 16999 45959
rect 17077 45913 17123 45959
rect 17201 45913 17247 45959
rect 17325 45913 17371 45959
rect 17449 45913 17495 45959
rect 17573 45913 17619 45959
rect 17697 45913 17743 45959
rect 17821 45913 17867 45959
rect 17945 45913 17991 45959
rect 18069 45913 18115 45959
rect 18193 45913 18239 45959
rect 18317 45913 18363 45959
rect 18441 45913 18487 45959
rect 18565 45913 18611 45959
rect 18689 45913 18735 45959
rect 18813 45913 18859 45959
rect 18937 45913 18983 45959
rect 19061 45913 19107 45959
rect 19185 45913 19231 45959
rect 19309 45913 19355 45959
rect 19433 45913 19479 45959
rect 19557 45913 19603 45959
rect 19681 45913 19727 45959
rect 19805 45913 19851 45959
rect 19929 45913 19975 45959
rect 20053 45913 20099 45959
rect 20177 45913 20223 45959
rect 20301 45913 20347 45959
rect 20425 45913 20471 45959
rect 20549 45913 20595 45959
rect 20673 45913 20719 45959
rect 20797 45913 20843 45959
rect 20921 45913 20967 45959
rect 21045 45913 21091 45959
rect 21169 45913 21215 45959
rect 21293 45913 21339 45959
rect 21417 45913 21463 45959
rect 21541 45913 21587 45959
rect 21665 45913 21711 45959
rect 21789 45913 21835 45959
rect 21913 45913 21959 45959
rect 22037 45913 22083 45959
rect 22161 45913 22207 45959
rect 22285 45913 22331 45959
rect 22409 45913 22455 45959
rect 22533 45913 22579 45959
rect 22657 45913 22703 45959
rect 22781 45913 22827 45959
rect 22905 45913 22951 45959
rect 23029 45913 23075 45959
rect 23153 45913 23199 45959
rect 23277 45913 23323 45959
rect 23401 45913 23447 45959
rect 23525 45913 23571 45959
rect 23649 45913 23695 45959
rect 23773 45913 23819 45959
rect 23897 45913 23943 45959
rect 24021 45913 24067 45959
rect 24145 45913 24191 45959
rect 24269 45913 24315 45959
rect 24393 45913 24439 45959
rect 24517 45913 24563 45959
rect 24641 45913 24687 45959
rect 24765 45913 24811 45959
rect 24889 45913 24935 45959
rect 25013 45913 25059 45959
rect 25137 45913 25183 45959
rect 25261 45913 25307 45959
rect 25385 45913 25431 45959
rect 25509 45913 25555 45959
rect 25633 45913 25679 45959
rect 25757 45913 25803 45959
rect 25881 45913 25927 45959
rect 26005 45913 26051 45959
rect 26129 45913 26175 45959
rect 26253 45913 26299 45959
rect 26377 45913 26423 45959
rect 26501 45913 26547 45959
rect 26625 45913 26671 45959
rect 26749 45913 26795 45959
rect 26873 45913 26919 45959
rect 26997 45913 27043 45959
rect 27121 45913 27167 45959
rect 27245 45913 27291 45959
rect 27369 45913 27415 45959
rect 27493 45913 27539 45959
rect 27617 45913 27663 45959
rect 27741 45913 27787 45959
rect 27865 45913 27911 45959
rect 27989 45913 28035 45959
rect 28113 45913 28159 45959
rect 28237 45913 28283 45959
rect 28361 45913 28407 45959
rect 28485 45913 28531 45959
rect 28609 45913 28655 45959
rect 28733 45913 28779 45959
rect 28857 45913 28903 45959
rect 28981 45913 29027 45959
rect 29105 45913 29151 45959
rect 29229 45913 29275 45959
rect 29353 45913 29399 45959
rect 29477 45913 29523 45959
rect 29601 45913 29647 45959
rect 29725 45913 29771 45959
rect 29849 45913 29895 45959
rect 29973 45913 30019 45959
rect 30097 45913 30143 45959
rect 30221 45913 30267 45959
rect 30345 45913 30391 45959
rect 30469 45913 30515 45959
rect 30593 45913 30639 45959
rect 30717 45913 30763 45959
rect 30841 45913 30887 45959
rect 30965 45913 31011 45959
rect 31089 45913 31135 45959
rect 31213 45913 31259 45959
rect 31337 45913 31383 45959
rect 31461 45913 31507 45959
rect 31585 45913 31631 45959
rect 31709 45913 31755 45959
rect 31833 45913 31879 45959
rect 31957 45913 32003 45959
rect 32081 45913 32127 45959
rect 32205 45913 32251 45959
rect 32329 45913 32375 45959
rect 32453 45913 32499 45959
rect 32577 45913 32623 45959
rect 32701 45913 32747 45959
rect 32825 45913 32871 45959
rect 32949 45913 32995 45959
rect 33073 45913 33119 45959
rect 33197 45913 33243 45959
rect 33321 45913 33367 45959
rect 33445 45913 33491 45959
rect 33569 45913 33615 45959
rect 33693 45913 33739 45959
rect 33817 45913 33863 45959
rect 33941 45913 33987 45959
rect 34065 45913 34111 45959
rect 34189 45913 34235 45959
rect 34313 45913 34359 45959
rect 34437 45913 34483 45959
rect 34561 45913 34607 45959
rect 34685 45913 34731 45959
rect 34809 45913 34855 45959
rect 34933 45913 34979 45959
rect 35057 45913 35103 45959
rect 35181 45913 35227 45959
rect 35305 45913 35351 45959
rect 35429 45913 35475 45959
rect 35553 45913 35599 45959
rect 35677 45913 35723 45959
rect 35801 45913 35847 45959
rect 35925 45913 35971 45959
rect 36049 45913 36095 45959
rect 36173 45913 36219 45959
rect 36297 45913 36343 45959
rect 36421 45913 36467 45959
rect 36545 45913 36591 45959
rect 36669 45913 36715 45959
rect 36793 45913 36839 45959
rect 36917 45913 36963 45959
rect 37041 45913 37087 45959
rect 37165 45913 37211 45959
rect 37289 45913 37335 45959
rect 37413 45913 37459 45959
rect 37537 45913 37583 45959
rect 37661 45913 37707 45959
rect 37785 45913 37831 45959
rect 37909 45913 37955 45959
rect 38033 45913 38079 45959
rect 38157 45913 38203 45959
rect 38281 45913 38327 45959
rect 38405 45913 38451 45959
rect 38529 45913 38575 45959
rect 38653 45913 38699 45959
rect 38777 45913 38823 45959
rect 38901 45913 38947 45959
rect 39025 45913 39071 45959
rect 39149 45913 39195 45959
rect 39273 45913 39319 45959
rect 39397 45913 39443 45959
rect 39521 45913 39567 45959
rect 39645 45913 39691 45959
rect 39769 45913 39815 45959
rect 39893 45913 39939 45959
rect 40017 45913 40063 45959
rect 40141 45913 40187 45959
rect 40265 45913 40311 45959
rect 40389 45913 40435 45959
rect 40513 45913 40559 45959
rect 40637 45913 40683 45959
rect 40761 45913 40807 45959
rect 40885 45913 40931 45959
rect 41009 45913 41055 45959
rect 41133 45913 41179 45959
rect 41257 45913 41303 45959
rect 41381 45913 41427 45959
rect 41505 45913 41551 45959
rect 41629 45913 41675 45959
rect 41753 45913 41799 45959
rect 41877 45913 41923 45959
rect 42001 45913 42047 45959
rect 42125 45913 42171 45959
rect 42249 45913 42295 45959
rect 42373 45913 42419 45959
rect 42497 45913 42543 45959
rect 42621 45913 42667 45959
rect 42745 45913 42791 45959
rect 42869 45913 42915 45959
rect 42993 45913 43039 45959
rect 43117 45913 43163 45959
rect 43241 45913 43287 45959
rect 43365 45913 43411 45959
rect 43489 45913 43535 45959
rect 43613 45913 43659 45959
rect 43737 45913 43783 45959
rect 43861 45913 43907 45959
rect 43985 45913 44031 45959
rect 44109 45913 44155 45959
rect 44233 45913 44279 45959
rect 44357 45913 44403 45959
rect 44481 45913 44527 45959
rect 44605 45913 44651 45959
rect 44729 45913 44775 45959
rect 44853 45913 44899 45959
rect 44977 45913 45023 45959
rect 45101 45913 45147 45959
rect 45225 45913 45271 45959
rect 45349 45913 45395 45959
rect 45473 45913 45519 45959
rect 45597 45913 45643 45959
rect 45721 45913 45767 45959
rect 45845 45913 45891 45959
rect 45969 45913 46015 45959
rect 46093 45913 46139 45959
rect 46217 45913 46263 45959
rect 46341 45913 46387 45959
rect 46465 45913 46511 45959
rect 46589 45913 46635 45959
rect 46713 45913 46759 45959
rect 46837 45913 46883 45959
rect 46961 45913 47007 45959
rect 47085 45913 47131 45959
rect 47209 45913 47255 45959
rect 47333 45913 47379 45959
rect 47457 45913 47503 45959
rect 47581 45913 47627 45959
rect 47705 45913 47751 45959
rect 47829 45913 47875 45959
rect 47953 45913 47999 45959
rect 48077 45913 48123 45959
rect 48201 45913 48247 45959
rect 48325 45913 48371 45959
rect 48449 45913 48495 45959
rect 48573 45913 48619 45959
rect 48697 45913 48743 45959
rect 48821 45913 48867 45959
rect 48945 45913 48991 45959
rect 49069 45913 49115 45959
rect 49193 45913 49239 45959
rect 49317 45913 49363 45959
rect 49441 45913 49487 45959
rect 49565 45913 49611 45959
rect 49689 45913 49735 45959
rect 49813 45913 49859 45959
rect 49937 45913 49983 45959
rect 50061 45913 50107 45959
rect 50185 45913 50231 45959
rect 50309 45913 50355 45959
rect 50433 45913 50479 45959
rect 50557 45913 50603 45959
rect 50681 45913 50727 45959
rect 50805 45913 50851 45959
rect 50929 45913 50975 45959
rect 51053 45913 51099 45959
rect 51177 45913 51223 45959
rect 51301 45913 51347 45959
rect 51425 45913 51471 45959
rect 51549 45913 51595 45959
rect 51673 45913 51719 45959
rect 51797 45913 51843 45959
rect 51921 45913 51967 45959
rect 52045 45913 52091 45959
rect 52169 45913 52215 45959
rect 52293 45913 52339 45959
rect 52417 45913 52463 45959
rect 52541 45913 52587 45959
rect 52665 45913 52711 45959
rect 52789 45913 52835 45959
rect 52913 45913 52959 45959
rect 53037 45913 53083 45959
rect 53161 45913 53207 45959
rect 53285 45913 53331 45959
rect 53409 45913 53455 45959
rect 53533 45913 53579 45959
rect 53657 45913 53703 45959
rect 53781 45913 53827 45959
rect 53905 45913 53951 45959
rect 54029 45913 54075 45959
rect 54153 45913 54199 45959
rect 54277 45913 54323 45959
rect 54401 45913 54447 45959
rect 54525 45913 54571 45959
rect 54649 45913 54695 45959
rect 54773 45913 54819 45959
rect 54897 45913 54943 45959
rect 55021 45913 55067 45959
rect 55145 45913 55191 45959
rect 55269 45913 55315 45959
rect 55393 45913 55439 45959
rect 55517 45913 55563 45959
rect 55641 45913 55687 45959
rect 55765 45913 55811 45959
rect 55889 45913 55935 45959
rect 56013 45913 56059 45959
rect 56137 45913 56183 45959
rect 56261 45913 56307 45959
rect 56385 45913 56431 45959
rect 56509 45913 56555 45959
rect 56633 45913 56679 45959
rect 56757 45913 56803 45959
rect 56881 45913 56927 45959
rect 57005 45913 57051 45959
rect 57129 45913 57175 45959
rect 57253 45913 57299 45959
rect 57377 45913 57423 45959
rect 57501 45913 57547 45959
rect 57625 45913 57671 45959
rect 57749 45913 57795 45959
rect 57873 45913 57919 45959
rect 57997 45913 58043 45959
rect 58121 45913 58167 45959
rect 58245 45913 58291 45959
rect 58369 45913 58415 45959
rect 58493 45913 58539 45959
rect 58617 45913 58663 45959
rect 58741 45913 58787 45959
rect 58865 45913 58911 45959
rect 58989 45913 59035 45959
rect 59113 45913 59159 45959
rect 59237 45913 59283 45959
rect 59361 45913 59407 45959
rect 59485 45913 59531 45959
rect 59609 45913 59655 45959
rect 59733 45913 59779 45959
rect 59857 45913 59903 45959
rect 59981 45913 60027 45959
rect 60105 45913 60151 45959
rect 60229 45913 60275 45959
rect 60353 45913 60399 45959
rect 60477 45913 60523 45959
rect 60601 45913 60647 45959
rect 60725 45913 60771 45959
rect 60849 45913 60895 45959
rect 60973 45913 61019 45959
rect 61097 45913 61143 45959
rect 61221 45913 61267 45959
rect 61345 45913 61391 45959
rect 61469 45913 61515 45959
rect 61593 45913 61639 45959
rect 61717 45913 61763 45959
rect 61841 45913 61887 45959
rect 61965 45913 62011 45959
rect 62089 45913 62135 45959
rect 62213 45913 62259 45959
rect 62337 45913 62383 45959
rect 62461 45913 62507 45959
rect 62585 45913 62631 45959
rect 62709 45913 62755 45959
rect 62833 45913 62879 45959
rect 62957 45913 63003 45959
rect 63081 45913 63127 45959
rect 63205 45913 63251 45959
rect 63329 45913 63375 45959
rect 63453 45913 63499 45959
rect 63577 45913 63623 45959
rect 63701 45913 63747 45959
rect 63825 45913 63871 45959
rect 63949 45913 63995 45959
rect 64073 45913 64119 45959
rect 64197 45913 64243 45959
rect 64321 45913 64367 45959
rect 64445 45913 64491 45959
rect 64569 45913 64615 45959
rect 64693 45913 64739 45959
rect 64817 45913 64863 45959
rect 64941 45913 64987 45959
rect 65065 45913 65111 45959
rect 65189 45913 65235 45959
rect 65313 45913 65359 45959
rect 65437 45913 65483 45959
rect 65561 45913 65607 45959
rect 65685 45913 65731 45959
rect 65809 45913 65855 45959
rect 65933 45913 65979 45959
rect 66057 45913 66103 45959
rect 66181 45913 66227 45959
rect 66305 45913 66351 45959
rect 66429 45913 66475 45959
rect 66553 45913 66599 45959
rect 66677 45913 66723 45959
rect 66801 45913 66847 45959
rect 66925 45913 66971 45959
rect 67049 45913 67095 45959
rect 67173 45913 67219 45959
rect 67297 45913 67343 45959
rect 67421 45913 67467 45959
rect 67545 45913 67591 45959
rect 67669 45913 67715 45959
rect 67793 45913 67839 45959
rect 67917 45913 67963 45959
rect 68041 45913 68087 45959
rect 68165 45913 68211 45959
rect 68289 45913 68335 45959
rect 68413 45913 68459 45959
rect 68537 45913 68583 45959
rect 68661 45913 68707 45959
rect 68785 45913 68831 45959
rect 68909 45913 68955 45959
rect 69033 45913 69079 45959
rect 69157 45913 69203 45959
rect 69281 45913 69327 45959
rect 69405 45913 69451 45959
rect 69529 45913 69575 45959
rect 69653 45913 69699 45959
rect 69777 45913 69823 45959
rect 69901 45913 69947 45959
rect 70025 45913 70071 45959
rect 70149 45913 70195 45959
rect 70273 45913 70319 45959
rect 70397 45913 70443 45959
rect 70521 45913 70567 45959
rect 70645 45913 70691 45959
rect 70769 45913 70815 45959
rect 70893 45913 70939 45959
rect 71017 45913 71063 45959
rect 71141 45913 71187 45959
rect 71265 45913 71311 45959
rect 71389 45913 71435 45959
rect 71513 45913 71559 45959
rect 71637 45913 71683 45959
rect 71761 45913 71807 45959
rect 71885 45913 71931 45959
rect 72009 45913 72055 45959
rect 72133 45913 72179 45959
rect 72257 45913 72303 45959
rect 72381 45913 72427 45959
rect 72505 45913 72551 45959
rect 72629 45913 72675 45959
rect 72753 45913 72799 45959
rect 72877 45913 72923 45959
rect 73001 45913 73047 45959
rect 73125 45913 73171 45959
rect 73249 45913 73295 45959
rect 73373 45913 73419 45959
rect 73497 45913 73543 45959
rect 73621 45913 73667 45959
rect 73745 45913 73791 45959
rect 73869 45913 73915 45959
rect 73993 45913 74039 45959
rect 74117 45913 74163 45959
rect 74241 45913 74287 45959
rect 74365 45913 74411 45959
rect 74489 45913 74535 45959
rect 74613 45913 74659 45959
rect 74737 45913 74783 45959
rect 74861 45913 74907 45959
rect 74985 45913 75031 45959
rect 75109 45913 75155 45959
rect 75233 45913 75279 45959
rect 75357 45913 75403 45959
rect 75481 45913 75527 45959
rect 75605 45913 75651 45959
rect 75729 45913 75775 45959
rect 75853 45913 75899 45959
rect 75977 45913 76023 45959
rect 76101 45913 76147 45959
rect 76225 45913 76271 45959
rect 76349 45913 76395 45959
rect 76473 45913 76519 45959
rect 76597 45913 76643 45959
rect 76721 45913 76767 45959
rect 76845 45913 76891 45959
rect 76969 45913 77015 45959
rect 77093 45913 77139 45959
rect 77217 45913 77263 45959
rect 77341 45913 77387 45959
rect 77465 45913 77511 45959
rect 77589 45913 77635 45959
rect 77713 45913 77759 45959
rect 77837 45913 77883 45959
rect 77961 45913 78007 45959
rect 78085 45913 78131 45959
rect 78209 45913 78255 45959
rect 78333 45913 78379 45959
rect 78457 45913 78503 45959
rect 78581 45913 78627 45959
rect 78705 45913 78751 45959
rect 78829 45913 78875 45959
rect 78953 45913 78999 45959
rect 79077 45913 79123 45959
rect 79201 45913 79247 45959
rect 79325 45913 79371 45959
rect 79449 45913 79495 45959
rect 79573 45913 79619 45959
rect 79697 45913 79743 45959
rect 79821 45913 79867 45959
rect 79945 45913 79991 45959
rect 80069 45913 80115 45959
rect 80193 45913 80239 45959
rect 80317 45913 80363 45959
rect 80441 45913 80487 45959
rect 80565 45913 80611 45959
rect 80689 45913 80735 45959
rect 80813 45913 80859 45959
rect 80937 45913 80983 45959
rect 81061 45913 81107 45959
rect 81185 45913 81231 45959
rect 81309 45913 81355 45959
rect 81433 45913 81479 45959
rect 81557 45913 81603 45959
rect 81681 45913 81727 45959
rect 81805 45913 81851 45959
rect 81929 45913 81975 45959
rect 82053 45913 82099 45959
rect 82177 45913 82223 45959
rect 82301 45913 82347 45959
rect 82425 45913 82471 45959
rect 82549 45913 82595 45959
rect 82673 45913 82719 45959
rect 82797 45913 82843 45959
rect 82921 45913 82967 45959
rect 83045 45913 83091 45959
rect 83169 45913 83215 45959
rect 83293 45913 83339 45959
rect 83417 45913 83463 45959
rect 83541 45913 83587 45959
rect 83665 45913 83711 45959
rect 83789 45913 83835 45959
rect 83913 45913 83959 45959
rect 84037 45913 84083 45959
rect 84161 45913 84207 45959
rect 84285 45913 84331 45959
rect 84409 45913 84455 45959
rect 84533 45913 84579 45959
rect 84657 45913 84703 45959
rect 84781 45913 84827 45959
rect 84905 45913 84951 45959
rect 85029 45913 85075 45959
rect 85153 45913 85199 45959
rect 85277 45913 85323 45959
rect 85401 45913 85447 45959
rect 85525 45913 85571 45959
rect 85649 45913 85695 45959
rect 89 45789 135 45835
rect 213 45789 259 45835
rect 337 45789 383 45835
rect 461 45789 507 45835
rect 585 45789 631 45835
rect 709 45789 755 45835
rect 833 45789 879 45835
rect 957 45789 1003 45835
rect 1081 45789 1127 45835
rect 1205 45789 1251 45835
rect 1329 45789 1375 45835
rect 1453 45789 1499 45835
rect 1577 45789 1623 45835
rect 1701 45789 1747 45835
rect 1825 45789 1871 45835
rect 1949 45789 1995 45835
rect 2073 45789 2119 45835
rect 2197 45789 2243 45835
rect 2321 45789 2367 45835
rect 2445 45789 2491 45835
rect 2569 45789 2615 45835
rect 2693 45789 2739 45835
rect 2817 45789 2863 45835
rect 2941 45789 2987 45835
rect 3065 45789 3111 45835
rect 3189 45789 3235 45835
rect 3313 45789 3359 45835
rect 3437 45789 3483 45835
rect 3561 45789 3607 45835
rect 3685 45789 3731 45835
rect 3809 45789 3855 45835
rect 3933 45789 3979 45835
rect 4057 45789 4103 45835
rect 4181 45789 4227 45835
rect 4305 45789 4351 45835
rect 4429 45789 4475 45835
rect 4553 45789 4599 45835
rect 4677 45789 4723 45835
rect 4801 45789 4847 45835
rect 4925 45789 4971 45835
rect 5049 45789 5095 45835
rect 5173 45789 5219 45835
rect 5297 45789 5343 45835
rect 5421 45789 5467 45835
rect 5545 45789 5591 45835
rect 5669 45789 5715 45835
rect 5793 45789 5839 45835
rect 5917 45789 5963 45835
rect 6041 45789 6087 45835
rect 6165 45789 6211 45835
rect 6289 45789 6335 45835
rect 6413 45789 6459 45835
rect 6537 45789 6583 45835
rect 6661 45789 6707 45835
rect 6785 45789 6831 45835
rect 6909 45789 6955 45835
rect 7033 45789 7079 45835
rect 7157 45789 7203 45835
rect 7281 45789 7327 45835
rect 7405 45789 7451 45835
rect 7529 45789 7575 45835
rect 7653 45789 7699 45835
rect 7777 45789 7823 45835
rect 7901 45789 7947 45835
rect 8025 45789 8071 45835
rect 8149 45789 8195 45835
rect 8273 45789 8319 45835
rect 8397 45789 8443 45835
rect 8521 45789 8567 45835
rect 8645 45789 8691 45835
rect 8769 45789 8815 45835
rect 8893 45789 8939 45835
rect 9017 45789 9063 45835
rect 9141 45789 9187 45835
rect 9265 45789 9311 45835
rect 9389 45789 9435 45835
rect 9513 45789 9559 45835
rect 9637 45789 9683 45835
rect 9761 45789 9807 45835
rect 9885 45789 9931 45835
rect 10009 45789 10055 45835
rect 10133 45789 10179 45835
rect 10257 45789 10303 45835
rect 10381 45789 10427 45835
rect 10505 45789 10551 45835
rect 10629 45789 10675 45835
rect 10753 45789 10799 45835
rect 10877 45789 10923 45835
rect 11001 45789 11047 45835
rect 11125 45789 11171 45835
rect 11249 45789 11295 45835
rect 11373 45789 11419 45835
rect 11497 45789 11543 45835
rect 11621 45789 11667 45835
rect 11745 45789 11791 45835
rect 11869 45789 11915 45835
rect 11993 45789 12039 45835
rect 12117 45789 12163 45835
rect 12241 45789 12287 45835
rect 12365 45789 12411 45835
rect 12489 45789 12535 45835
rect 12613 45789 12659 45835
rect 12737 45789 12783 45835
rect 12861 45789 12907 45835
rect 12985 45789 13031 45835
rect 13109 45789 13155 45835
rect 13233 45789 13279 45835
rect 13357 45789 13403 45835
rect 13481 45789 13527 45835
rect 13605 45789 13651 45835
rect 13729 45789 13775 45835
rect 13853 45789 13899 45835
rect 13977 45789 14023 45835
rect 14101 45789 14147 45835
rect 14225 45789 14271 45835
rect 14349 45789 14395 45835
rect 14473 45789 14519 45835
rect 14597 45789 14643 45835
rect 14721 45789 14767 45835
rect 14845 45789 14891 45835
rect 14969 45789 15015 45835
rect 15093 45789 15139 45835
rect 15217 45789 15263 45835
rect 15341 45789 15387 45835
rect 15465 45789 15511 45835
rect 15589 45789 15635 45835
rect 15713 45789 15759 45835
rect 15837 45789 15883 45835
rect 15961 45789 16007 45835
rect 16085 45789 16131 45835
rect 16209 45789 16255 45835
rect 16333 45789 16379 45835
rect 16457 45789 16503 45835
rect 16581 45789 16627 45835
rect 16705 45789 16751 45835
rect 16829 45789 16875 45835
rect 16953 45789 16999 45835
rect 17077 45789 17123 45835
rect 17201 45789 17247 45835
rect 17325 45789 17371 45835
rect 17449 45789 17495 45835
rect 17573 45789 17619 45835
rect 17697 45789 17743 45835
rect 17821 45789 17867 45835
rect 17945 45789 17991 45835
rect 18069 45789 18115 45835
rect 18193 45789 18239 45835
rect 18317 45789 18363 45835
rect 18441 45789 18487 45835
rect 18565 45789 18611 45835
rect 18689 45789 18735 45835
rect 18813 45789 18859 45835
rect 18937 45789 18983 45835
rect 19061 45789 19107 45835
rect 19185 45789 19231 45835
rect 19309 45789 19355 45835
rect 19433 45789 19479 45835
rect 19557 45789 19603 45835
rect 19681 45789 19727 45835
rect 19805 45789 19851 45835
rect 19929 45789 19975 45835
rect 20053 45789 20099 45835
rect 20177 45789 20223 45835
rect 20301 45789 20347 45835
rect 20425 45789 20471 45835
rect 20549 45789 20595 45835
rect 20673 45789 20719 45835
rect 20797 45789 20843 45835
rect 20921 45789 20967 45835
rect 21045 45789 21091 45835
rect 21169 45789 21215 45835
rect 21293 45789 21339 45835
rect 21417 45789 21463 45835
rect 21541 45789 21587 45835
rect 21665 45789 21711 45835
rect 21789 45789 21835 45835
rect 21913 45789 21959 45835
rect 22037 45789 22083 45835
rect 22161 45789 22207 45835
rect 22285 45789 22331 45835
rect 22409 45789 22455 45835
rect 22533 45789 22579 45835
rect 22657 45789 22703 45835
rect 22781 45789 22827 45835
rect 22905 45789 22951 45835
rect 23029 45789 23075 45835
rect 23153 45789 23199 45835
rect 23277 45789 23323 45835
rect 23401 45789 23447 45835
rect 23525 45789 23571 45835
rect 23649 45789 23695 45835
rect 23773 45789 23819 45835
rect 23897 45789 23943 45835
rect 24021 45789 24067 45835
rect 24145 45789 24191 45835
rect 24269 45789 24315 45835
rect 24393 45789 24439 45835
rect 24517 45789 24563 45835
rect 24641 45789 24687 45835
rect 24765 45789 24811 45835
rect 24889 45789 24935 45835
rect 25013 45789 25059 45835
rect 25137 45789 25183 45835
rect 25261 45789 25307 45835
rect 25385 45789 25431 45835
rect 25509 45789 25555 45835
rect 25633 45789 25679 45835
rect 25757 45789 25803 45835
rect 25881 45789 25927 45835
rect 26005 45789 26051 45835
rect 26129 45789 26175 45835
rect 26253 45789 26299 45835
rect 26377 45789 26423 45835
rect 26501 45789 26547 45835
rect 26625 45789 26671 45835
rect 26749 45789 26795 45835
rect 26873 45789 26919 45835
rect 26997 45789 27043 45835
rect 27121 45789 27167 45835
rect 27245 45789 27291 45835
rect 27369 45789 27415 45835
rect 27493 45789 27539 45835
rect 27617 45789 27663 45835
rect 27741 45789 27787 45835
rect 27865 45789 27911 45835
rect 27989 45789 28035 45835
rect 28113 45789 28159 45835
rect 28237 45789 28283 45835
rect 28361 45789 28407 45835
rect 28485 45789 28531 45835
rect 28609 45789 28655 45835
rect 28733 45789 28779 45835
rect 28857 45789 28903 45835
rect 28981 45789 29027 45835
rect 29105 45789 29151 45835
rect 29229 45789 29275 45835
rect 29353 45789 29399 45835
rect 29477 45789 29523 45835
rect 29601 45789 29647 45835
rect 29725 45789 29771 45835
rect 29849 45789 29895 45835
rect 29973 45789 30019 45835
rect 30097 45789 30143 45835
rect 30221 45789 30267 45835
rect 30345 45789 30391 45835
rect 30469 45789 30515 45835
rect 30593 45789 30639 45835
rect 30717 45789 30763 45835
rect 30841 45789 30887 45835
rect 30965 45789 31011 45835
rect 31089 45789 31135 45835
rect 31213 45789 31259 45835
rect 31337 45789 31383 45835
rect 31461 45789 31507 45835
rect 31585 45789 31631 45835
rect 31709 45789 31755 45835
rect 31833 45789 31879 45835
rect 31957 45789 32003 45835
rect 32081 45789 32127 45835
rect 32205 45789 32251 45835
rect 32329 45789 32375 45835
rect 32453 45789 32499 45835
rect 32577 45789 32623 45835
rect 32701 45789 32747 45835
rect 32825 45789 32871 45835
rect 32949 45789 32995 45835
rect 33073 45789 33119 45835
rect 33197 45789 33243 45835
rect 33321 45789 33367 45835
rect 33445 45789 33491 45835
rect 33569 45789 33615 45835
rect 33693 45789 33739 45835
rect 33817 45789 33863 45835
rect 33941 45789 33987 45835
rect 34065 45789 34111 45835
rect 34189 45789 34235 45835
rect 34313 45789 34359 45835
rect 34437 45789 34483 45835
rect 34561 45789 34607 45835
rect 34685 45789 34731 45835
rect 34809 45789 34855 45835
rect 34933 45789 34979 45835
rect 35057 45789 35103 45835
rect 35181 45789 35227 45835
rect 35305 45789 35351 45835
rect 35429 45789 35475 45835
rect 35553 45789 35599 45835
rect 35677 45789 35723 45835
rect 35801 45789 35847 45835
rect 35925 45789 35971 45835
rect 36049 45789 36095 45835
rect 36173 45789 36219 45835
rect 36297 45789 36343 45835
rect 36421 45789 36467 45835
rect 36545 45789 36591 45835
rect 36669 45789 36715 45835
rect 36793 45789 36839 45835
rect 36917 45789 36963 45835
rect 37041 45789 37087 45835
rect 37165 45789 37211 45835
rect 37289 45789 37335 45835
rect 37413 45789 37459 45835
rect 37537 45789 37583 45835
rect 37661 45789 37707 45835
rect 37785 45789 37831 45835
rect 37909 45789 37955 45835
rect 38033 45789 38079 45835
rect 38157 45789 38203 45835
rect 38281 45789 38327 45835
rect 38405 45789 38451 45835
rect 38529 45789 38575 45835
rect 38653 45789 38699 45835
rect 38777 45789 38823 45835
rect 38901 45789 38947 45835
rect 39025 45789 39071 45835
rect 39149 45789 39195 45835
rect 39273 45789 39319 45835
rect 39397 45789 39443 45835
rect 39521 45789 39567 45835
rect 39645 45789 39691 45835
rect 39769 45789 39815 45835
rect 39893 45789 39939 45835
rect 40017 45789 40063 45835
rect 40141 45789 40187 45835
rect 40265 45789 40311 45835
rect 40389 45789 40435 45835
rect 40513 45789 40559 45835
rect 40637 45789 40683 45835
rect 40761 45789 40807 45835
rect 40885 45789 40931 45835
rect 41009 45789 41055 45835
rect 41133 45789 41179 45835
rect 41257 45789 41303 45835
rect 41381 45789 41427 45835
rect 41505 45789 41551 45835
rect 41629 45789 41675 45835
rect 41753 45789 41799 45835
rect 41877 45789 41923 45835
rect 42001 45789 42047 45835
rect 42125 45789 42171 45835
rect 42249 45789 42295 45835
rect 42373 45789 42419 45835
rect 42497 45789 42543 45835
rect 42621 45789 42667 45835
rect 42745 45789 42791 45835
rect 42869 45789 42915 45835
rect 42993 45789 43039 45835
rect 43117 45789 43163 45835
rect 43241 45789 43287 45835
rect 43365 45789 43411 45835
rect 43489 45789 43535 45835
rect 43613 45789 43659 45835
rect 43737 45789 43783 45835
rect 43861 45789 43907 45835
rect 43985 45789 44031 45835
rect 44109 45789 44155 45835
rect 44233 45789 44279 45835
rect 44357 45789 44403 45835
rect 44481 45789 44527 45835
rect 44605 45789 44651 45835
rect 44729 45789 44775 45835
rect 44853 45789 44899 45835
rect 44977 45789 45023 45835
rect 45101 45789 45147 45835
rect 45225 45789 45271 45835
rect 45349 45789 45395 45835
rect 45473 45789 45519 45835
rect 45597 45789 45643 45835
rect 45721 45789 45767 45835
rect 45845 45789 45891 45835
rect 45969 45789 46015 45835
rect 46093 45789 46139 45835
rect 46217 45789 46263 45835
rect 46341 45789 46387 45835
rect 46465 45789 46511 45835
rect 46589 45789 46635 45835
rect 46713 45789 46759 45835
rect 46837 45789 46883 45835
rect 46961 45789 47007 45835
rect 47085 45789 47131 45835
rect 47209 45789 47255 45835
rect 47333 45789 47379 45835
rect 47457 45789 47503 45835
rect 47581 45789 47627 45835
rect 47705 45789 47751 45835
rect 47829 45789 47875 45835
rect 47953 45789 47999 45835
rect 48077 45789 48123 45835
rect 48201 45789 48247 45835
rect 48325 45789 48371 45835
rect 48449 45789 48495 45835
rect 48573 45789 48619 45835
rect 48697 45789 48743 45835
rect 48821 45789 48867 45835
rect 48945 45789 48991 45835
rect 49069 45789 49115 45835
rect 49193 45789 49239 45835
rect 49317 45789 49363 45835
rect 49441 45789 49487 45835
rect 49565 45789 49611 45835
rect 49689 45789 49735 45835
rect 49813 45789 49859 45835
rect 49937 45789 49983 45835
rect 50061 45789 50107 45835
rect 50185 45789 50231 45835
rect 50309 45789 50355 45835
rect 50433 45789 50479 45835
rect 50557 45789 50603 45835
rect 50681 45789 50727 45835
rect 50805 45789 50851 45835
rect 50929 45789 50975 45835
rect 51053 45789 51099 45835
rect 51177 45789 51223 45835
rect 51301 45789 51347 45835
rect 51425 45789 51471 45835
rect 51549 45789 51595 45835
rect 51673 45789 51719 45835
rect 51797 45789 51843 45835
rect 51921 45789 51967 45835
rect 52045 45789 52091 45835
rect 52169 45789 52215 45835
rect 52293 45789 52339 45835
rect 52417 45789 52463 45835
rect 52541 45789 52587 45835
rect 52665 45789 52711 45835
rect 52789 45789 52835 45835
rect 52913 45789 52959 45835
rect 53037 45789 53083 45835
rect 53161 45789 53207 45835
rect 53285 45789 53331 45835
rect 53409 45789 53455 45835
rect 53533 45789 53579 45835
rect 53657 45789 53703 45835
rect 53781 45789 53827 45835
rect 53905 45789 53951 45835
rect 54029 45789 54075 45835
rect 54153 45789 54199 45835
rect 54277 45789 54323 45835
rect 54401 45789 54447 45835
rect 54525 45789 54571 45835
rect 54649 45789 54695 45835
rect 54773 45789 54819 45835
rect 54897 45789 54943 45835
rect 55021 45789 55067 45835
rect 55145 45789 55191 45835
rect 55269 45789 55315 45835
rect 55393 45789 55439 45835
rect 55517 45789 55563 45835
rect 55641 45789 55687 45835
rect 55765 45789 55811 45835
rect 55889 45789 55935 45835
rect 56013 45789 56059 45835
rect 56137 45789 56183 45835
rect 56261 45789 56307 45835
rect 56385 45789 56431 45835
rect 56509 45789 56555 45835
rect 56633 45789 56679 45835
rect 56757 45789 56803 45835
rect 56881 45789 56927 45835
rect 57005 45789 57051 45835
rect 57129 45789 57175 45835
rect 57253 45789 57299 45835
rect 57377 45789 57423 45835
rect 57501 45789 57547 45835
rect 57625 45789 57671 45835
rect 57749 45789 57795 45835
rect 57873 45789 57919 45835
rect 57997 45789 58043 45835
rect 58121 45789 58167 45835
rect 58245 45789 58291 45835
rect 58369 45789 58415 45835
rect 58493 45789 58539 45835
rect 58617 45789 58663 45835
rect 58741 45789 58787 45835
rect 58865 45789 58911 45835
rect 58989 45789 59035 45835
rect 59113 45789 59159 45835
rect 59237 45789 59283 45835
rect 59361 45789 59407 45835
rect 59485 45789 59531 45835
rect 59609 45789 59655 45835
rect 59733 45789 59779 45835
rect 59857 45789 59903 45835
rect 59981 45789 60027 45835
rect 60105 45789 60151 45835
rect 60229 45789 60275 45835
rect 60353 45789 60399 45835
rect 60477 45789 60523 45835
rect 60601 45789 60647 45835
rect 60725 45789 60771 45835
rect 60849 45789 60895 45835
rect 60973 45789 61019 45835
rect 61097 45789 61143 45835
rect 61221 45789 61267 45835
rect 61345 45789 61391 45835
rect 61469 45789 61515 45835
rect 61593 45789 61639 45835
rect 61717 45789 61763 45835
rect 61841 45789 61887 45835
rect 61965 45789 62011 45835
rect 62089 45789 62135 45835
rect 62213 45789 62259 45835
rect 62337 45789 62383 45835
rect 62461 45789 62507 45835
rect 62585 45789 62631 45835
rect 62709 45789 62755 45835
rect 62833 45789 62879 45835
rect 62957 45789 63003 45835
rect 63081 45789 63127 45835
rect 63205 45789 63251 45835
rect 63329 45789 63375 45835
rect 63453 45789 63499 45835
rect 63577 45789 63623 45835
rect 63701 45789 63747 45835
rect 63825 45789 63871 45835
rect 63949 45789 63995 45835
rect 64073 45789 64119 45835
rect 64197 45789 64243 45835
rect 64321 45789 64367 45835
rect 64445 45789 64491 45835
rect 64569 45789 64615 45835
rect 64693 45789 64739 45835
rect 64817 45789 64863 45835
rect 64941 45789 64987 45835
rect 65065 45789 65111 45835
rect 65189 45789 65235 45835
rect 65313 45789 65359 45835
rect 65437 45789 65483 45835
rect 65561 45789 65607 45835
rect 65685 45789 65731 45835
rect 65809 45789 65855 45835
rect 65933 45789 65979 45835
rect 66057 45789 66103 45835
rect 66181 45789 66227 45835
rect 66305 45789 66351 45835
rect 66429 45789 66475 45835
rect 66553 45789 66599 45835
rect 66677 45789 66723 45835
rect 66801 45789 66847 45835
rect 66925 45789 66971 45835
rect 67049 45789 67095 45835
rect 67173 45789 67219 45835
rect 67297 45789 67343 45835
rect 67421 45789 67467 45835
rect 67545 45789 67591 45835
rect 67669 45789 67715 45835
rect 67793 45789 67839 45835
rect 67917 45789 67963 45835
rect 68041 45789 68087 45835
rect 68165 45789 68211 45835
rect 68289 45789 68335 45835
rect 68413 45789 68459 45835
rect 68537 45789 68583 45835
rect 68661 45789 68707 45835
rect 68785 45789 68831 45835
rect 68909 45789 68955 45835
rect 69033 45789 69079 45835
rect 69157 45789 69203 45835
rect 69281 45789 69327 45835
rect 69405 45789 69451 45835
rect 69529 45789 69575 45835
rect 69653 45789 69699 45835
rect 69777 45789 69823 45835
rect 69901 45789 69947 45835
rect 70025 45789 70071 45835
rect 70149 45789 70195 45835
rect 70273 45789 70319 45835
rect 70397 45789 70443 45835
rect 70521 45789 70567 45835
rect 70645 45789 70691 45835
rect 70769 45789 70815 45835
rect 70893 45789 70939 45835
rect 71017 45789 71063 45835
rect 71141 45789 71187 45835
rect 71265 45789 71311 45835
rect 71389 45789 71435 45835
rect 71513 45789 71559 45835
rect 71637 45789 71683 45835
rect 71761 45789 71807 45835
rect 71885 45789 71931 45835
rect 72009 45789 72055 45835
rect 72133 45789 72179 45835
rect 72257 45789 72303 45835
rect 72381 45789 72427 45835
rect 72505 45789 72551 45835
rect 72629 45789 72675 45835
rect 72753 45789 72799 45835
rect 72877 45789 72923 45835
rect 73001 45789 73047 45835
rect 73125 45789 73171 45835
rect 73249 45789 73295 45835
rect 73373 45789 73419 45835
rect 73497 45789 73543 45835
rect 73621 45789 73667 45835
rect 73745 45789 73791 45835
rect 73869 45789 73915 45835
rect 73993 45789 74039 45835
rect 74117 45789 74163 45835
rect 74241 45789 74287 45835
rect 74365 45789 74411 45835
rect 74489 45789 74535 45835
rect 74613 45789 74659 45835
rect 74737 45789 74783 45835
rect 74861 45789 74907 45835
rect 74985 45789 75031 45835
rect 75109 45789 75155 45835
rect 75233 45789 75279 45835
rect 75357 45789 75403 45835
rect 75481 45789 75527 45835
rect 75605 45789 75651 45835
rect 75729 45789 75775 45835
rect 75853 45789 75899 45835
rect 75977 45789 76023 45835
rect 76101 45789 76147 45835
rect 76225 45789 76271 45835
rect 76349 45789 76395 45835
rect 76473 45789 76519 45835
rect 76597 45789 76643 45835
rect 76721 45789 76767 45835
rect 76845 45789 76891 45835
rect 76969 45789 77015 45835
rect 77093 45789 77139 45835
rect 77217 45789 77263 45835
rect 77341 45789 77387 45835
rect 77465 45789 77511 45835
rect 77589 45789 77635 45835
rect 77713 45789 77759 45835
rect 77837 45789 77883 45835
rect 77961 45789 78007 45835
rect 78085 45789 78131 45835
rect 78209 45789 78255 45835
rect 78333 45789 78379 45835
rect 78457 45789 78503 45835
rect 78581 45789 78627 45835
rect 78705 45789 78751 45835
rect 78829 45789 78875 45835
rect 78953 45789 78999 45835
rect 79077 45789 79123 45835
rect 79201 45789 79247 45835
rect 79325 45789 79371 45835
rect 79449 45789 79495 45835
rect 79573 45789 79619 45835
rect 79697 45789 79743 45835
rect 79821 45789 79867 45835
rect 79945 45789 79991 45835
rect 80069 45789 80115 45835
rect 80193 45789 80239 45835
rect 80317 45789 80363 45835
rect 80441 45789 80487 45835
rect 80565 45789 80611 45835
rect 80689 45789 80735 45835
rect 80813 45789 80859 45835
rect 80937 45789 80983 45835
rect 81061 45789 81107 45835
rect 81185 45789 81231 45835
rect 81309 45789 81355 45835
rect 81433 45789 81479 45835
rect 81557 45789 81603 45835
rect 81681 45789 81727 45835
rect 81805 45789 81851 45835
rect 81929 45789 81975 45835
rect 82053 45789 82099 45835
rect 82177 45789 82223 45835
rect 82301 45789 82347 45835
rect 82425 45789 82471 45835
rect 82549 45789 82595 45835
rect 82673 45789 82719 45835
rect 82797 45789 82843 45835
rect 82921 45789 82967 45835
rect 83045 45789 83091 45835
rect 83169 45789 83215 45835
rect 83293 45789 83339 45835
rect 83417 45789 83463 45835
rect 83541 45789 83587 45835
rect 83665 45789 83711 45835
rect 83789 45789 83835 45835
rect 83913 45789 83959 45835
rect 84037 45789 84083 45835
rect 84161 45789 84207 45835
rect 84285 45789 84331 45835
rect 84409 45789 84455 45835
rect 84533 45789 84579 45835
rect 84657 45789 84703 45835
rect 84781 45789 84827 45835
rect 84905 45789 84951 45835
rect 85029 45789 85075 45835
rect 85153 45789 85199 45835
rect 85277 45789 85323 45835
rect 85401 45789 85447 45835
rect 85525 45789 85571 45835
rect 85649 45789 85695 45835
rect 89 45665 135 45711
rect 213 45665 259 45711
rect 337 45665 383 45711
rect 461 45665 507 45711
rect 585 45665 631 45711
rect 709 45665 755 45711
rect 833 45665 879 45711
rect 957 45665 1003 45711
rect 1081 45665 1127 45711
rect 1205 45665 1251 45711
rect 1329 45665 1375 45711
rect 1453 45665 1499 45711
rect 1577 45665 1623 45711
rect 1701 45665 1747 45711
rect 1825 45665 1871 45711
rect 1949 45665 1995 45711
rect 2073 45665 2119 45711
rect 2197 45665 2243 45711
rect 2321 45665 2367 45711
rect 2445 45665 2491 45711
rect 2569 45665 2615 45711
rect 2693 45665 2739 45711
rect 2817 45665 2863 45711
rect 2941 45665 2987 45711
rect 3065 45665 3111 45711
rect 3189 45665 3235 45711
rect 3313 45665 3359 45711
rect 3437 45665 3483 45711
rect 3561 45665 3607 45711
rect 3685 45665 3731 45711
rect 3809 45665 3855 45711
rect 3933 45665 3979 45711
rect 4057 45665 4103 45711
rect 4181 45665 4227 45711
rect 4305 45665 4351 45711
rect 4429 45665 4475 45711
rect 4553 45665 4599 45711
rect 4677 45665 4723 45711
rect 4801 45665 4847 45711
rect 4925 45665 4971 45711
rect 5049 45665 5095 45711
rect 5173 45665 5219 45711
rect 5297 45665 5343 45711
rect 5421 45665 5467 45711
rect 5545 45665 5591 45711
rect 5669 45665 5715 45711
rect 5793 45665 5839 45711
rect 5917 45665 5963 45711
rect 6041 45665 6087 45711
rect 6165 45665 6211 45711
rect 6289 45665 6335 45711
rect 6413 45665 6459 45711
rect 6537 45665 6583 45711
rect 6661 45665 6707 45711
rect 6785 45665 6831 45711
rect 6909 45665 6955 45711
rect 7033 45665 7079 45711
rect 7157 45665 7203 45711
rect 7281 45665 7327 45711
rect 7405 45665 7451 45711
rect 7529 45665 7575 45711
rect 7653 45665 7699 45711
rect 7777 45665 7823 45711
rect 7901 45665 7947 45711
rect 8025 45665 8071 45711
rect 8149 45665 8195 45711
rect 8273 45665 8319 45711
rect 8397 45665 8443 45711
rect 8521 45665 8567 45711
rect 8645 45665 8691 45711
rect 8769 45665 8815 45711
rect 8893 45665 8939 45711
rect 9017 45665 9063 45711
rect 9141 45665 9187 45711
rect 9265 45665 9311 45711
rect 9389 45665 9435 45711
rect 9513 45665 9559 45711
rect 9637 45665 9683 45711
rect 9761 45665 9807 45711
rect 9885 45665 9931 45711
rect 10009 45665 10055 45711
rect 10133 45665 10179 45711
rect 10257 45665 10303 45711
rect 10381 45665 10427 45711
rect 10505 45665 10551 45711
rect 10629 45665 10675 45711
rect 10753 45665 10799 45711
rect 10877 45665 10923 45711
rect 11001 45665 11047 45711
rect 11125 45665 11171 45711
rect 11249 45665 11295 45711
rect 11373 45665 11419 45711
rect 11497 45665 11543 45711
rect 11621 45665 11667 45711
rect 11745 45665 11791 45711
rect 11869 45665 11915 45711
rect 11993 45665 12039 45711
rect 12117 45665 12163 45711
rect 12241 45665 12287 45711
rect 12365 45665 12411 45711
rect 12489 45665 12535 45711
rect 12613 45665 12659 45711
rect 12737 45665 12783 45711
rect 12861 45665 12907 45711
rect 12985 45665 13031 45711
rect 13109 45665 13155 45711
rect 13233 45665 13279 45711
rect 13357 45665 13403 45711
rect 13481 45665 13527 45711
rect 13605 45665 13651 45711
rect 13729 45665 13775 45711
rect 13853 45665 13899 45711
rect 13977 45665 14023 45711
rect 14101 45665 14147 45711
rect 14225 45665 14271 45711
rect 14349 45665 14395 45711
rect 14473 45665 14519 45711
rect 14597 45665 14643 45711
rect 14721 45665 14767 45711
rect 14845 45665 14891 45711
rect 14969 45665 15015 45711
rect 15093 45665 15139 45711
rect 15217 45665 15263 45711
rect 15341 45665 15387 45711
rect 15465 45665 15511 45711
rect 15589 45665 15635 45711
rect 15713 45665 15759 45711
rect 15837 45665 15883 45711
rect 15961 45665 16007 45711
rect 16085 45665 16131 45711
rect 16209 45665 16255 45711
rect 16333 45665 16379 45711
rect 16457 45665 16503 45711
rect 16581 45665 16627 45711
rect 16705 45665 16751 45711
rect 16829 45665 16875 45711
rect 16953 45665 16999 45711
rect 17077 45665 17123 45711
rect 17201 45665 17247 45711
rect 17325 45665 17371 45711
rect 17449 45665 17495 45711
rect 17573 45665 17619 45711
rect 17697 45665 17743 45711
rect 17821 45665 17867 45711
rect 17945 45665 17991 45711
rect 18069 45665 18115 45711
rect 18193 45665 18239 45711
rect 18317 45665 18363 45711
rect 18441 45665 18487 45711
rect 18565 45665 18611 45711
rect 18689 45665 18735 45711
rect 18813 45665 18859 45711
rect 18937 45665 18983 45711
rect 19061 45665 19107 45711
rect 19185 45665 19231 45711
rect 19309 45665 19355 45711
rect 19433 45665 19479 45711
rect 19557 45665 19603 45711
rect 19681 45665 19727 45711
rect 19805 45665 19851 45711
rect 19929 45665 19975 45711
rect 20053 45665 20099 45711
rect 20177 45665 20223 45711
rect 20301 45665 20347 45711
rect 20425 45665 20471 45711
rect 20549 45665 20595 45711
rect 20673 45665 20719 45711
rect 20797 45665 20843 45711
rect 20921 45665 20967 45711
rect 21045 45665 21091 45711
rect 21169 45665 21215 45711
rect 21293 45665 21339 45711
rect 21417 45665 21463 45711
rect 21541 45665 21587 45711
rect 21665 45665 21711 45711
rect 21789 45665 21835 45711
rect 21913 45665 21959 45711
rect 22037 45665 22083 45711
rect 22161 45665 22207 45711
rect 22285 45665 22331 45711
rect 22409 45665 22455 45711
rect 22533 45665 22579 45711
rect 22657 45665 22703 45711
rect 22781 45665 22827 45711
rect 22905 45665 22951 45711
rect 23029 45665 23075 45711
rect 23153 45665 23199 45711
rect 23277 45665 23323 45711
rect 23401 45665 23447 45711
rect 23525 45665 23571 45711
rect 23649 45665 23695 45711
rect 23773 45665 23819 45711
rect 23897 45665 23943 45711
rect 24021 45665 24067 45711
rect 24145 45665 24191 45711
rect 24269 45665 24315 45711
rect 24393 45665 24439 45711
rect 24517 45665 24563 45711
rect 24641 45665 24687 45711
rect 24765 45665 24811 45711
rect 24889 45665 24935 45711
rect 25013 45665 25059 45711
rect 25137 45665 25183 45711
rect 25261 45665 25307 45711
rect 25385 45665 25431 45711
rect 25509 45665 25555 45711
rect 25633 45665 25679 45711
rect 25757 45665 25803 45711
rect 25881 45665 25927 45711
rect 26005 45665 26051 45711
rect 26129 45665 26175 45711
rect 26253 45665 26299 45711
rect 26377 45665 26423 45711
rect 26501 45665 26547 45711
rect 26625 45665 26671 45711
rect 26749 45665 26795 45711
rect 26873 45665 26919 45711
rect 26997 45665 27043 45711
rect 27121 45665 27167 45711
rect 27245 45665 27291 45711
rect 27369 45665 27415 45711
rect 27493 45665 27539 45711
rect 27617 45665 27663 45711
rect 27741 45665 27787 45711
rect 27865 45665 27911 45711
rect 27989 45665 28035 45711
rect 28113 45665 28159 45711
rect 28237 45665 28283 45711
rect 28361 45665 28407 45711
rect 28485 45665 28531 45711
rect 28609 45665 28655 45711
rect 28733 45665 28779 45711
rect 28857 45665 28903 45711
rect 28981 45665 29027 45711
rect 29105 45665 29151 45711
rect 29229 45665 29275 45711
rect 29353 45665 29399 45711
rect 29477 45665 29523 45711
rect 29601 45665 29647 45711
rect 29725 45665 29771 45711
rect 29849 45665 29895 45711
rect 29973 45665 30019 45711
rect 30097 45665 30143 45711
rect 30221 45665 30267 45711
rect 30345 45665 30391 45711
rect 30469 45665 30515 45711
rect 30593 45665 30639 45711
rect 30717 45665 30763 45711
rect 30841 45665 30887 45711
rect 30965 45665 31011 45711
rect 31089 45665 31135 45711
rect 31213 45665 31259 45711
rect 31337 45665 31383 45711
rect 31461 45665 31507 45711
rect 31585 45665 31631 45711
rect 31709 45665 31755 45711
rect 31833 45665 31879 45711
rect 31957 45665 32003 45711
rect 32081 45665 32127 45711
rect 32205 45665 32251 45711
rect 32329 45665 32375 45711
rect 32453 45665 32499 45711
rect 32577 45665 32623 45711
rect 32701 45665 32747 45711
rect 32825 45665 32871 45711
rect 32949 45665 32995 45711
rect 33073 45665 33119 45711
rect 33197 45665 33243 45711
rect 33321 45665 33367 45711
rect 33445 45665 33491 45711
rect 33569 45665 33615 45711
rect 33693 45665 33739 45711
rect 33817 45665 33863 45711
rect 33941 45665 33987 45711
rect 34065 45665 34111 45711
rect 34189 45665 34235 45711
rect 34313 45665 34359 45711
rect 34437 45665 34483 45711
rect 34561 45665 34607 45711
rect 34685 45665 34731 45711
rect 34809 45665 34855 45711
rect 34933 45665 34979 45711
rect 35057 45665 35103 45711
rect 35181 45665 35227 45711
rect 35305 45665 35351 45711
rect 35429 45665 35475 45711
rect 35553 45665 35599 45711
rect 35677 45665 35723 45711
rect 35801 45665 35847 45711
rect 35925 45665 35971 45711
rect 36049 45665 36095 45711
rect 36173 45665 36219 45711
rect 36297 45665 36343 45711
rect 36421 45665 36467 45711
rect 36545 45665 36591 45711
rect 36669 45665 36715 45711
rect 36793 45665 36839 45711
rect 36917 45665 36963 45711
rect 37041 45665 37087 45711
rect 37165 45665 37211 45711
rect 37289 45665 37335 45711
rect 37413 45665 37459 45711
rect 37537 45665 37583 45711
rect 37661 45665 37707 45711
rect 37785 45665 37831 45711
rect 37909 45665 37955 45711
rect 38033 45665 38079 45711
rect 38157 45665 38203 45711
rect 38281 45665 38327 45711
rect 38405 45665 38451 45711
rect 38529 45665 38575 45711
rect 38653 45665 38699 45711
rect 38777 45665 38823 45711
rect 38901 45665 38947 45711
rect 39025 45665 39071 45711
rect 39149 45665 39195 45711
rect 39273 45665 39319 45711
rect 39397 45665 39443 45711
rect 39521 45665 39567 45711
rect 39645 45665 39691 45711
rect 39769 45665 39815 45711
rect 39893 45665 39939 45711
rect 40017 45665 40063 45711
rect 40141 45665 40187 45711
rect 40265 45665 40311 45711
rect 40389 45665 40435 45711
rect 40513 45665 40559 45711
rect 40637 45665 40683 45711
rect 40761 45665 40807 45711
rect 40885 45665 40931 45711
rect 41009 45665 41055 45711
rect 41133 45665 41179 45711
rect 41257 45665 41303 45711
rect 41381 45665 41427 45711
rect 41505 45665 41551 45711
rect 41629 45665 41675 45711
rect 41753 45665 41799 45711
rect 41877 45665 41923 45711
rect 42001 45665 42047 45711
rect 42125 45665 42171 45711
rect 42249 45665 42295 45711
rect 42373 45665 42419 45711
rect 42497 45665 42543 45711
rect 42621 45665 42667 45711
rect 42745 45665 42791 45711
rect 42869 45665 42915 45711
rect 42993 45665 43039 45711
rect 43117 45665 43163 45711
rect 43241 45665 43287 45711
rect 43365 45665 43411 45711
rect 43489 45665 43535 45711
rect 43613 45665 43659 45711
rect 43737 45665 43783 45711
rect 43861 45665 43907 45711
rect 43985 45665 44031 45711
rect 44109 45665 44155 45711
rect 44233 45665 44279 45711
rect 44357 45665 44403 45711
rect 44481 45665 44527 45711
rect 44605 45665 44651 45711
rect 44729 45665 44775 45711
rect 44853 45665 44899 45711
rect 44977 45665 45023 45711
rect 45101 45665 45147 45711
rect 45225 45665 45271 45711
rect 45349 45665 45395 45711
rect 45473 45665 45519 45711
rect 45597 45665 45643 45711
rect 45721 45665 45767 45711
rect 45845 45665 45891 45711
rect 45969 45665 46015 45711
rect 46093 45665 46139 45711
rect 46217 45665 46263 45711
rect 46341 45665 46387 45711
rect 46465 45665 46511 45711
rect 46589 45665 46635 45711
rect 46713 45665 46759 45711
rect 46837 45665 46883 45711
rect 46961 45665 47007 45711
rect 47085 45665 47131 45711
rect 47209 45665 47255 45711
rect 47333 45665 47379 45711
rect 47457 45665 47503 45711
rect 47581 45665 47627 45711
rect 47705 45665 47751 45711
rect 47829 45665 47875 45711
rect 47953 45665 47999 45711
rect 48077 45665 48123 45711
rect 48201 45665 48247 45711
rect 48325 45665 48371 45711
rect 48449 45665 48495 45711
rect 48573 45665 48619 45711
rect 48697 45665 48743 45711
rect 48821 45665 48867 45711
rect 48945 45665 48991 45711
rect 49069 45665 49115 45711
rect 49193 45665 49239 45711
rect 49317 45665 49363 45711
rect 49441 45665 49487 45711
rect 49565 45665 49611 45711
rect 49689 45665 49735 45711
rect 49813 45665 49859 45711
rect 49937 45665 49983 45711
rect 50061 45665 50107 45711
rect 50185 45665 50231 45711
rect 50309 45665 50355 45711
rect 50433 45665 50479 45711
rect 50557 45665 50603 45711
rect 50681 45665 50727 45711
rect 50805 45665 50851 45711
rect 50929 45665 50975 45711
rect 51053 45665 51099 45711
rect 51177 45665 51223 45711
rect 51301 45665 51347 45711
rect 51425 45665 51471 45711
rect 51549 45665 51595 45711
rect 51673 45665 51719 45711
rect 51797 45665 51843 45711
rect 51921 45665 51967 45711
rect 52045 45665 52091 45711
rect 52169 45665 52215 45711
rect 52293 45665 52339 45711
rect 52417 45665 52463 45711
rect 52541 45665 52587 45711
rect 52665 45665 52711 45711
rect 52789 45665 52835 45711
rect 52913 45665 52959 45711
rect 53037 45665 53083 45711
rect 53161 45665 53207 45711
rect 53285 45665 53331 45711
rect 53409 45665 53455 45711
rect 53533 45665 53579 45711
rect 53657 45665 53703 45711
rect 53781 45665 53827 45711
rect 53905 45665 53951 45711
rect 54029 45665 54075 45711
rect 54153 45665 54199 45711
rect 54277 45665 54323 45711
rect 54401 45665 54447 45711
rect 54525 45665 54571 45711
rect 54649 45665 54695 45711
rect 54773 45665 54819 45711
rect 54897 45665 54943 45711
rect 55021 45665 55067 45711
rect 55145 45665 55191 45711
rect 55269 45665 55315 45711
rect 55393 45665 55439 45711
rect 55517 45665 55563 45711
rect 55641 45665 55687 45711
rect 55765 45665 55811 45711
rect 55889 45665 55935 45711
rect 56013 45665 56059 45711
rect 56137 45665 56183 45711
rect 56261 45665 56307 45711
rect 56385 45665 56431 45711
rect 56509 45665 56555 45711
rect 56633 45665 56679 45711
rect 56757 45665 56803 45711
rect 56881 45665 56927 45711
rect 57005 45665 57051 45711
rect 57129 45665 57175 45711
rect 57253 45665 57299 45711
rect 57377 45665 57423 45711
rect 57501 45665 57547 45711
rect 57625 45665 57671 45711
rect 57749 45665 57795 45711
rect 57873 45665 57919 45711
rect 57997 45665 58043 45711
rect 58121 45665 58167 45711
rect 58245 45665 58291 45711
rect 58369 45665 58415 45711
rect 58493 45665 58539 45711
rect 58617 45665 58663 45711
rect 58741 45665 58787 45711
rect 58865 45665 58911 45711
rect 58989 45665 59035 45711
rect 59113 45665 59159 45711
rect 59237 45665 59283 45711
rect 59361 45665 59407 45711
rect 59485 45665 59531 45711
rect 59609 45665 59655 45711
rect 59733 45665 59779 45711
rect 59857 45665 59903 45711
rect 59981 45665 60027 45711
rect 60105 45665 60151 45711
rect 60229 45665 60275 45711
rect 60353 45665 60399 45711
rect 60477 45665 60523 45711
rect 60601 45665 60647 45711
rect 60725 45665 60771 45711
rect 60849 45665 60895 45711
rect 60973 45665 61019 45711
rect 61097 45665 61143 45711
rect 61221 45665 61267 45711
rect 61345 45665 61391 45711
rect 61469 45665 61515 45711
rect 61593 45665 61639 45711
rect 61717 45665 61763 45711
rect 61841 45665 61887 45711
rect 61965 45665 62011 45711
rect 62089 45665 62135 45711
rect 62213 45665 62259 45711
rect 62337 45665 62383 45711
rect 62461 45665 62507 45711
rect 62585 45665 62631 45711
rect 62709 45665 62755 45711
rect 62833 45665 62879 45711
rect 62957 45665 63003 45711
rect 63081 45665 63127 45711
rect 63205 45665 63251 45711
rect 63329 45665 63375 45711
rect 63453 45665 63499 45711
rect 63577 45665 63623 45711
rect 63701 45665 63747 45711
rect 63825 45665 63871 45711
rect 63949 45665 63995 45711
rect 64073 45665 64119 45711
rect 64197 45665 64243 45711
rect 64321 45665 64367 45711
rect 64445 45665 64491 45711
rect 64569 45665 64615 45711
rect 64693 45665 64739 45711
rect 64817 45665 64863 45711
rect 64941 45665 64987 45711
rect 65065 45665 65111 45711
rect 65189 45665 65235 45711
rect 65313 45665 65359 45711
rect 65437 45665 65483 45711
rect 65561 45665 65607 45711
rect 65685 45665 65731 45711
rect 65809 45665 65855 45711
rect 65933 45665 65979 45711
rect 66057 45665 66103 45711
rect 66181 45665 66227 45711
rect 66305 45665 66351 45711
rect 66429 45665 66475 45711
rect 66553 45665 66599 45711
rect 66677 45665 66723 45711
rect 66801 45665 66847 45711
rect 66925 45665 66971 45711
rect 67049 45665 67095 45711
rect 67173 45665 67219 45711
rect 67297 45665 67343 45711
rect 67421 45665 67467 45711
rect 67545 45665 67591 45711
rect 67669 45665 67715 45711
rect 67793 45665 67839 45711
rect 67917 45665 67963 45711
rect 68041 45665 68087 45711
rect 68165 45665 68211 45711
rect 68289 45665 68335 45711
rect 68413 45665 68459 45711
rect 68537 45665 68583 45711
rect 68661 45665 68707 45711
rect 68785 45665 68831 45711
rect 68909 45665 68955 45711
rect 69033 45665 69079 45711
rect 69157 45665 69203 45711
rect 69281 45665 69327 45711
rect 69405 45665 69451 45711
rect 69529 45665 69575 45711
rect 69653 45665 69699 45711
rect 69777 45665 69823 45711
rect 69901 45665 69947 45711
rect 70025 45665 70071 45711
rect 70149 45665 70195 45711
rect 70273 45665 70319 45711
rect 70397 45665 70443 45711
rect 70521 45665 70567 45711
rect 70645 45665 70691 45711
rect 70769 45665 70815 45711
rect 70893 45665 70939 45711
rect 71017 45665 71063 45711
rect 71141 45665 71187 45711
rect 71265 45665 71311 45711
rect 71389 45665 71435 45711
rect 71513 45665 71559 45711
rect 71637 45665 71683 45711
rect 71761 45665 71807 45711
rect 71885 45665 71931 45711
rect 72009 45665 72055 45711
rect 72133 45665 72179 45711
rect 72257 45665 72303 45711
rect 72381 45665 72427 45711
rect 72505 45665 72551 45711
rect 72629 45665 72675 45711
rect 72753 45665 72799 45711
rect 72877 45665 72923 45711
rect 73001 45665 73047 45711
rect 73125 45665 73171 45711
rect 73249 45665 73295 45711
rect 73373 45665 73419 45711
rect 73497 45665 73543 45711
rect 73621 45665 73667 45711
rect 73745 45665 73791 45711
rect 73869 45665 73915 45711
rect 73993 45665 74039 45711
rect 74117 45665 74163 45711
rect 74241 45665 74287 45711
rect 74365 45665 74411 45711
rect 74489 45665 74535 45711
rect 74613 45665 74659 45711
rect 74737 45665 74783 45711
rect 74861 45665 74907 45711
rect 74985 45665 75031 45711
rect 75109 45665 75155 45711
rect 75233 45665 75279 45711
rect 75357 45665 75403 45711
rect 75481 45665 75527 45711
rect 75605 45665 75651 45711
rect 75729 45665 75775 45711
rect 75853 45665 75899 45711
rect 75977 45665 76023 45711
rect 76101 45665 76147 45711
rect 76225 45665 76271 45711
rect 76349 45665 76395 45711
rect 76473 45665 76519 45711
rect 76597 45665 76643 45711
rect 76721 45665 76767 45711
rect 76845 45665 76891 45711
rect 76969 45665 77015 45711
rect 77093 45665 77139 45711
rect 77217 45665 77263 45711
rect 77341 45665 77387 45711
rect 77465 45665 77511 45711
rect 77589 45665 77635 45711
rect 77713 45665 77759 45711
rect 77837 45665 77883 45711
rect 77961 45665 78007 45711
rect 78085 45665 78131 45711
rect 78209 45665 78255 45711
rect 78333 45665 78379 45711
rect 78457 45665 78503 45711
rect 78581 45665 78627 45711
rect 78705 45665 78751 45711
rect 78829 45665 78875 45711
rect 78953 45665 78999 45711
rect 79077 45665 79123 45711
rect 79201 45665 79247 45711
rect 79325 45665 79371 45711
rect 79449 45665 79495 45711
rect 79573 45665 79619 45711
rect 79697 45665 79743 45711
rect 79821 45665 79867 45711
rect 79945 45665 79991 45711
rect 80069 45665 80115 45711
rect 80193 45665 80239 45711
rect 80317 45665 80363 45711
rect 80441 45665 80487 45711
rect 80565 45665 80611 45711
rect 80689 45665 80735 45711
rect 80813 45665 80859 45711
rect 80937 45665 80983 45711
rect 81061 45665 81107 45711
rect 81185 45665 81231 45711
rect 81309 45665 81355 45711
rect 81433 45665 81479 45711
rect 81557 45665 81603 45711
rect 81681 45665 81727 45711
rect 81805 45665 81851 45711
rect 81929 45665 81975 45711
rect 82053 45665 82099 45711
rect 82177 45665 82223 45711
rect 82301 45665 82347 45711
rect 82425 45665 82471 45711
rect 82549 45665 82595 45711
rect 82673 45665 82719 45711
rect 82797 45665 82843 45711
rect 82921 45665 82967 45711
rect 83045 45665 83091 45711
rect 83169 45665 83215 45711
rect 83293 45665 83339 45711
rect 83417 45665 83463 45711
rect 83541 45665 83587 45711
rect 83665 45665 83711 45711
rect 83789 45665 83835 45711
rect 83913 45665 83959 45711
rect 84037 45665 84083 45711
rect 84161 45665 84207 45711
rect 84285 45665 84331 45711
rect 84409 45665 84455 45711
rect 84533 45665 84579 45711
rect 84657 45665 84703 45711
rect 84781 45665 84827 45711
rect 84905 45665 84951 45711
rect 85029 45665 85075 45711
rect 85153 45665 85199 45711
rect 85277 45665 85323 45711
rect 85401 45665 85447 45711
rect 85525 45665 85571 45711
rect 85649 45665 85695 45711
rect 89 1117 435 45563
rect 85451 1117 85797 45563
rect 89 969 135 1015
rect 213 969 259 1015
rect 337 969 383 1015
rect 461 969 507 1015
rect 585 969 631 1015
rect 709 969 755 1015
rect 833 969 879 1015
rect 957 969 1003 1015
rect 1081 969 1127 1015
rect 1205 969 1251 1015
rect 1329 969 1375 1015
rect 1453 969 1499 1015
rect 1577 969 1623 1015
rect 1701 969 1747 1015
rect 1825 969 1871 1015
rect 1949 969 1995 1015
rect 2073 969 2119 1015
rect 2197 969 2243 1015
rect 2321 969 2367 1015
rect 2445 969 2491 1015
rect 2569 969 2615 1015
rect 2693 969 2739 1015
rect 2817 969 2863 1015
rect 2941 969 2987 1015
rect 3065 969 3111 1015
rect 3189 969 3235 1015
rect 3313 969 3359 1015
rect 3437 969 3483 1015
rect 3561 969 3607 1015
rect 3685 969 3731 1015
rect 3809 969 3855 1015
rect 3933 969 3979 1015
rect 4057 969 4103 1015
rect 4181 969 4227 1015
rect 4305 969 4351 1015
rect 4429 969 4475 1015
rect 4553 969 4599 1015
rect 4677 969 4723 1015
rect 4801 969 4847 1015
rect 4925 969 4971 1015
rect 5049 969 5095 1015
rect 5173 969 5219 1015
rect 5297 969 5343 1015
rect 5421 969 5467 1015
rect 5545 969 5591 1015
rect 5669 969 5715 1015
rect 5793 969 5839 1015
rect 5917 969 5963 1015
rect 6041 969 6087 1015
rect 6165 969 6211 1015
rect 6289 969 6335 1015
rect 6413 969 6459 1015
rect 6537 969 6583 1015
rect 6661 969 6707 1015
rect 6785 969 6831 1015
rect 6909 969 6955 1015
rect 7033 969 7079 1015
rect 7157 969 7203 1015
rect 7281 969 7327 1015
rect 7405 969 7451 1015
rect 7529 969 7575 1015
rect 7653 969 7699 1015
rect 7777 969 7823 1015
rect 7901 969 7947 1015
rect 8025 969 8071 1015
rect 8149 969 8195 1015
rect 8273 969 8319 1015
rect 8397 969 8443 1015
rect 8521 969 8567 1015
rect 8645 969 8691 1015
rect 8769 969 8815 1015
rect 8893 969 8939 1015
rect 9017 969 9063 1015
rect 9141 969 9187 1015
rect 9265 969 9311 1015
rect 9389 969 9435 1015
rect 9513 969 9559 1015
rect 9637 969 9683 1015
rect 9761 969 9807 1015
rect 9885 969 9931 1015
rect 10009 969 10055 1015
rect 10133 969 10179 1015
rect 10257 969 10303 1015
rect 10381 969 10427 1015
rect 10505 969 10551 1015
rect 10629 969 10675 1015
rect 10753 969 10799 1015
rect 10877 969 10923 1015
rect 11001 969 11047 1015
rect 11125 969 11171 1015
rect 11249 969 11295 1015
rect 11373 969 11419 1015
rect 11497 969 11543 1015
rect 11621 969 11667 1015
rect 11745 969 11791 1015
rect 11869 969 11915 1015
rect 11993 969 12039 1015
rect 12117 969 12163 1015
rect 12241 969 12287 1015
rect 12365 969 12411 1015
rect 12489 969 12535 1015
rect 12613 969 12659 1015
rect 12737 969 12783 1015
rect 12861 969 12907 1015
rect 12985 969 13031 1015
rect 13109 969 13155 1015
rect 13233 969 13279 1015
rect 13357 969 13403 1015
rect 13481 969 13527 1015
rect 13605 969 13651 1015
rect 13729 969 13775 1015
rect 13853 969 13899 1015
rect 13977 969 14023 1015
rect 14101 969 14147 1015
rect 14225 969 14271 1015
rect 14349 969 14395 1015
rect 14473 969 14519 1015
rect 14597 969 14643 1015
rect 14721 969 14767 1015
rect 14845 969 14891 1015
rect 14969 969 15015 1015
rect 15093 969 15139 1015
rect 15217 969 15263 1015
rect 15341 969 15387 1015
rect 15465 969 15511 1015
rect 15589 969 15635 1015
rect 15713 969 15759 1015
rect 15837 969 15883 1015
rect 15961 969 16007 1015
rect 16085 969 16131 1015
rect 16209 969 16255 1015
rect 16333 969 16379 1015
rect 16457 969 16503 1015
rect 16581 969 16627 1015
rect 16705 969 16751 1015
rect 16829 969 16875 1015
rect 16953 969 16999 1015
rect 17077 969 17123 1015
rect 17201 969 17247 1015
rect 17325 969 17371 1015
rect 17449 969 17495 1015
rect 17573 969 17619 1015
rect 17697 969 17743 1015
rect 17821 969 17867 1015
rect 17945 969 17991 1015
rect 18069 969 18115 1015
rect 18193 969 18239 1015
rect 18317 969 18363 1015
rect 18441 969 18487 1015
rect 18565 969 18611 1015
rect 18689 969 18735 1015
rect 18813 969 18859 1015
rect 18937 969 18983 1015
rect 19061 969 19107 1015
rect 19185 969 19231 1015
rect 19309 969 19355 1015
rect 19433 969 19479 1015
rect 19557 969 19603 1015
rect 19681 969 19727 1015
rect 19805 969 19851 1015
rect 19929 969 19975 1015
rect 20053 969 20099 1015
rect 20177 969 20223 1015
rect 20301 969 20347 1015
rect 20425 969 20471 1015
rect 20549 969 20595 1015
rect 20673 969 20719 1015
rect 20797 969 20843 1015
rect 20921 969 20967 1015
rect 21045 969 21091 1015
rect 21169 969 21215 1015
rect 21293 969 21339 1015
rect 21417 969 21463 1015
rect 21541 969 21587 1015
rect 21665 969 21711 1015
rect 21789 969 21835 1015
rect 21913 969 21959 1015
rect 22037 969 22083 1015
rect 22161 969 22207 1015
rect 22285 969 22331 1015
rect 22409 969 22455 1015
rect 22533 969 22579 1015
rect 22657 969 22703 1015
rect 22781 969 22827 1015
rect 22905 969 22951 1015
rect 23029 969 23075 1015
rect 23153 969 23199 1015
rect 23277 969 23323 1015
rect 23401 969 23447 1015
rect 23525 969 23571 1015
rect 23649 969 23695 1015
rect 23773 969 23819 1015
rect 23897 969 23943 1015
rect 24021 969 24067 1015
rect 24145 969 24191 1015
rect 24269 969 24315 1015
rect 24393 969 24439 1015
rect 24517 969 24563 1015
rect 24641 969 24687 1015
rect 24765 969 24811 1015
rect 24889 969 24935 1015
rect 25013 969 25059 1015
rect 25137 969 25183 1015
rect 25261 969 25307 1015
rect 25385 969 25431 1015
rect 25509 969 25555 1015
rect 25633 969 25679 1015
rect 25757 969 25803 1015
rect 25881 969 25927 1015
rect 26005 969 26051 1015
rect 26129 969 26175 1015
rect 26253 969 26299 1015
rect 26377 969 26423 1015
rect 26501 969 26547 1015
rect 26625 969 26671 1015
rect 26749 969 26795 1015
rect 26873 969 26919 1015
rect 26997 969 27043 1015
rect 27121 969 27167 1015
rect 27245 969 27291 1015
rect 27369 969 27415 1015
rect 27493 969 27539 1015
rect 27617 969 27663 1015
rect 27741 969 27787 1015
rect 27865 969 27911 1015
rect 27989 969 28035 1015
rect 28113 969 28159 1015
rect 28237 969 28283 1015
rect 28361 969 28407 1015
rect 28485 969 28531 1015
rect 28609 969 28655 1015
rect 28733 969 28779 1015
rect 28857 969 28903 1015
rect 28981 969 29027 1015
rect 29105 969 29151 1015
rect 29229 969 29275 1015
rect 29353 969 29399 1015
rect 29477 969 29523 1015
rect 29601 969 29647 1015
rect 29725 969 29771 1015
rect 29849 969 29895 1015
rect 29973 969 30019 1015
rect 30097 969 30143 1015
rect 30221 969 30267 1015
rect 30345 969 30391 1015
rect 30469 969 30515 1015
rect 30593 969 30639 1015
rect 30717 969 30763 1015
rect 30841 969 30887 1015
rect 30965 969 31011 1015
rect 31089 969 31135 1015
rect 31213 969 31259 1015
rect 31337 969 31383 1015
rect 31461 969 31507 1015
rect 31585 969 31631 1015
rect 31709 969 31755 1015
rect 31833 969 31879 1015
rect 31957 969 32003 1015
rect 32081 969 32127 1015
rect 32205 969 32251 1015
rect 32329 969 32375 1015
rect 32453 969 32499 1015
rect 32577 969 32623 1015
rect 32701 969 32747 1015
rect 32825 969 32871 1015
rect 32949 969 32995 1015
rect 33073 969 33119 1015
rect 33197 969 33243 1015
rect 33321 969 33367 1015
rect 33445 969 33491 1015
rect 33569 969 33615 1015
rect 33693 969 33739 1015
rect 33817 969 33863 1015
rect 33941 969 33987 1015
rect 34065 969 34111 1015
rect 34189 969 34235 1015
rect 34313 969 34359 1015
rect 34437 969 34483 1015
rect 34561 969 34607 1015
rect 34685 969 34731 1015
rect 34809 969 34855 1015
rect 34933 969 34979 1015
rect 35057 969 35103 1015
rect 35181 969 35227 1015
rect 35305 969 35351 1015
rect 35429 969 35475 1015
rect 35553 969 35599 1015
rect 35677 969 35723 1015
rect 35801 969 35847 1015
rect 35925 969 35971 1015
rect 36049 969 36095 1015
rect 36173 969 36219 1015
rect 36297 969 36343 1015
rect 36421 969 36467 1015
rect 36545 969 36591 1015
rect 36669 969 36715 1015
rect 36793 969 36839 1015
rect 36917 969 36963 1015
rect 37041 969 37087 1015
rect 37165 969 37211 1015
rect 37289 969 37335 1015
rect 37413 969 37459 1015
rect 37537 969 37583 1015
rect 37661 969 37707 1015
rect 37785 969 37831 1015
rect 37909 969 37955 1015
rect 38033 969 38079 1015
rect 38157 969 38203 1015
rect 38281 969 38327 1015
rect 38405 969 38451 1015
rect 38529 969 38575 1015
rect 38653 969 38699 1015
rect 38777 969 38823 1015
rect 38901 969 38947 1015
rect 39025 969 39071 1015
rect 39149 969 39195 1015
rect 39273 969 39319 1015
rect 39397 969 39443 1015
rect 39521 969 39567 1015
rect 39645 969 39691 1015
rect 39769 969 39815 1015
rect 39893 969 39939 1015
rect 40017 969 40063 1015
rect 40141 969 40187 1015
rect 40265 969 40311 1015
rect 40389 969 40435 1015
rect 40513 969 40559 1015
rect 40637 969 40683 1015
rect 40761 969 40807 1015
rect 40885 969 40931 1015
rect 41009 969 41055 1015
rect 41133 969 41179 1015
rect 41257 969 41303 1015
rect 41381 969 41427 1015
rect 41505 969 41551 1015
rect 41629 969 41675 1015
rect 41753 969 41799 1015
rect 41877 969 41923 1015
rect 42001 969 42047 1015
rect 42125 969 42171 1015
rect 42249 969 42295 1015
rect 42373 969 42419 1015
rect 42497 969 42543 1015
rect 42621 969 42667 1015
rect 42745 969 42791 1015
rect 42869 969 42915 1015
rect 42993 969 43039 1015
rect 43117 969 43163 1015
rect 43241 969 43287 1015
rect 43365 969 43411 1015
rect 43489 969 43535 1015
rect 43613 969 43659 1015
rect 43737 969 43783 1015
rect 43861 969 43907 1015
rect 43985 969 44031 1015
rect 44109 969 44155 1015
rect 44233 969 44279 1015
rect 44357 969 44403 1015
rect 44481 969 44527 1015
rect 44605 969 44651 1015
rect 44729 969 44775 1015
rect 44853 969 44899 1015
rect 44977 969 45023 1015
rect 45101 969 45147 1015
rect 45225 969 45271 1015
rect 45349 969 45395 1015
rect 45473 969 45519 1015
rect 45597 969 45643 1015
rect 45721 969 45767 1015
rect 45845 969 45891 1015
rect 45969 969 46015 1015
rect 46093 969 46139 1015
rect 46217 969 46263 1015
rect 46341 969 46387 1015
rect 46465 969 46511 1015
rect 46589 969 46635 1015
rect 46713 969 46759 1015
rect 46837 969 46883 1015
rect 46961 969 47007 1015
rect 47085 969 47131 1015
rect 47209 969 47255 1015
rect 47333 969 47379 1015
rect 47457 969 47503 1015
rect 47581 969 47627 1015
rect 47705 969 47751 1015
rect 47829 969 47875 1015
rect 47953 969 47999 1015
rect 48077 969 48123 1015
rect 48201 969 48247 1015
rect 48325 969 48371 1015
rect 48449 969 48495 1015
rect 48573 969 48619 1015
rect 48697 969 48743 1015
rect 48821 969 48867 1015
rect 48945 969 48991 1015
rect 49069 969 49115 1015
rect 49193 969 49239 1015
rect 49317 969 49363 1015
rect 49441 969 49487 1015
rect 49565 969 49611 1015
rect 49689 969 49735 1015
rect 49813 969 49859 1015
rect 49937 969 49983 1015
rect 50061 969 50107 1015
rect 50185 969 50231 1015
rect 50309 969 50355 1015
rect 50433 969 50479 1015
rect 50557 969 50603 1015
rect 50681 969 50727 1015
rect 50805 969 50851 1015
rect 50929 969 50975 1015
rect 51053 969 51099 1015
rect 51177 969 51223 1015
rect 51301 969 51347 1015
rect 51425 969 51471 1015
rect 51549 969 51595 1015
rect 51673 969 51719 1015
rect 51797 969 51843 1015
rect 51921 969 51967 1015
rect 52045 969 52091 1015
rect 52169 969 52215 1015
rect 52293 969 52339 1015
rect 52417 969 52463 1015
rect 52541 969 52587 1015
rect 52665 969 52711 1015
rect 52789 969 52835 1015
rect 52913 969 52959 1015
rect 53037 969 53083 1015
rect 53161 969 53207 1015
rect 53285 969 53331 1015
rect 53409 969 53455 1015
rect 53533 969 53579 1015
rect 53657 969 53703 1015
rect 53781 969 53827 1015
rect 53905 969 53951 1015
rect 54029 969 54075 1015
rect 54153 969 54199 1015
rect 54277 969 54323 1015
rect 54401 969 54447 1015
rect 54525 969 54571 1015
rect 54649 969 54695 1015
rect 54773 969 54819 1015
rect 54897 969 54943 1015
rect 55021 969 55067 1015
rect 55145 969 55191 1015
rect 55269 969 55315 1015
rect 55393 969 55439 1015
rect 55517 969 55563 1015
rect 55641 969 55687 1015
rect 55765 969 55811 1015
rect 55889 969 55935 1015
rect 56013 969 56059 1015
rect 56137 969 56183 1015
rect 56261 969 56307 1015
rect 56385 969 56431 1015
rect 56509 969 56555 1015
rect 56633 969 56679 1015
rect 56757 969 56803 1015
rect 56881 969 56927 1015
rect 57005 969 57051 1015
rect 57129 969 57175 1015
rect 57253 969 57299 1015
rect 57377 969 57423 1015
rect 57501 969 57547 1015
rect 57625 969 57671 1015
rect 57749 969 57795 1015
rect 57873 969 57919 1015
rect 57997 969 58043 1015
rect 58121 969 58167 1015
rect 58245 969 58291 1015
rect 58369 969 58415 1015
rect 58493 969 58539 1015
rect 58617 969 58663 1015
rect 58741 969 58787 1015
rect 58865 969 58911 1015
rect 58989 969 59035 1015
rect 59113 969 59159 1015
rect 59237 969 59283 1015
rect 59361 969 59407 1015
rect 59485 969 59531 1015
rect 59609 969 59655 1015
rect 59733 969 59779 1015
rect 59857 969 59903 1015
rect 59981 969 60027 1015
rect 60105 969 60151 1015
rect 60229 969 60275 1015
rect 60353 969 60399 1015
rect 60477 969 60523 1015
rect 60601 969 60647 1015
rect 60725 969 60771 1015
rect 60849 969 60895 1015
rect 60973 969 61019 1015
rect 61097 969 61143 1015
rect 61221 969 61267 1015
rect 61345 969 61391 1015
rect 61469 969 61515 1015
rect 61593 969 61639 1015
rect 61717 969 61763 1015
rect 61841 969 61887 1015
rect 61965 969 62011 1015
rect 62089 969 62135 1015
rect 62213 969 62259 1015
rect 62337 969 62383 1015
rect 62461 969 62507 1015
rect 62585 969 62631 1015
rect 62709 969 62755 1015
rect 62833 969 62879 1015
rect 62957 969 63003 1015
rect 63081 969 63127 1015
rect 63205 969 63251 1015
rect 63329 969 63375 1015
rect 63453 969 63499 1015
rect 63577 969 63623 1015
rect 63701 969 63747 1015
rect 63825 969 63871 1015
rect 63949 969 63995 1015
rect 64073 969 64119 1015
rect 64197 969 64243 1015
rect 64321 969 64367 1015
rect 64445 969 64491 1015
rect 64569 969 64615 1015
rect 64693 969 64739 1015
rect 64817 969 64863 1015
rect 64941 969 64987 1015
rect 65065 969 65111 1015
rect 65189 969 65235 1015
rect 65313 969 65359 1015
rect 65437 969 65483 1015
rect 65561 969 65607 1015
rect 65685 969 65731 1015
rect 65809 969 65855 1015
rect 65933 969 65979 1015
rect 66057 969 66103 1015
rect 66181 969 66227 1015
rect 66305 969 66351 1015
rect 66429 969 66475 1015
rect 66553 969 66599 1015
rect 66677 969 66723 1015
rect 66801 969 66847 1015
rect 66925 969 66971 1015
rect 67049 969 67095 1015
rect 67173 969 67219 1015
rect 67297 969 67343 1015
rect 67421 969 67467 1015
rect 67545 969 67591 1015
rect 67669 969 67715 1015
rect 67793 969 67839 1015
rect 67917 969 67963 1015
rect 68041 969 68087 1015
rect 68165 969 68211 1015
rect 68289 969 68335 1015
rect 68413 969 68459 1015
rect 68537 969 68583 1015
rect 68661 969 68707 1015
rect 68785 969 68831 1015
rect 68909 969 68955 1015
rect 69033 969 69079 1015
rect 69157 969 69203 1015
rect 69281 969 69327 1015
rect 69405 969 69451 1015
rect 69529 969 69575 1015
rect 69653 969 69699 1015
rect 69777 969 69823 1015
rect 69901 969 69947 1015
rect 70025 969 70071 1015
rect 70149 969 70195 1015
rect 70273 969 70319 1015
rect 70397 969 70443 1015
rect 70521 969 70567 1015
rect 70645 969 70691 1015
rect 70769 969 70815 1015
rect 70893 969 70939 1015
rect 71017 969 71063 1015
rect 71141 969 71187 1015
rect 71265 969 71311 1015
rect 71389 969 71435 1015
rect 71513 969 71559 1015
rect 71637 969 71683 1015
rect 71761 969 71807 1015
rect 71885 969 71931 1015
rect 72009 969 72055 1015
rect 72133 969 72179 1015
rect 72257 969 72303 1015
rect 72381 969 72427 1015
rect 72505 969 72551 1015
rect 72629 969 72675 1015
rect 72753 969 72799 1015
rect 72877 969 72923 1015
rect 73001 969 73047 1015
rect 73125 969 73171 1015
rect 73249 969 73295 1015
rect 73373 969 73419 1015
rect 73497 969 73543 1015
rect 73621 969 73667 1015
rect 73745 969 73791 1015
rect 73869 969 73915 1015
rect 73993 969 74039 1015
rect 74117 969 74163 1015
rect 74241 969 74287 1015
rect 74365 969 74411 1015
rect 74489 969 74535 1015
rect 74613 969 74659 1015
rect 74737 969 74783 1015
rect 74861 969 74907 1015
rect 74985 969 75031 1015
rect 75109 969 75155 1015
rect 75233 969 75279 1015
rect 75357 969 75403 1015
rect 75481 969 75527 1015
rect 75605 969 75651 1015
rect 75729 969 75775 1015
rect 75853 969 75899 1015
rect 75977 969 76023 1015
rect 76101 969 76147 1015
rect 76225 969 76271 1015
rect 76349 969 76395 1015
rect 76473 969 76519 1015
rect 76597 969 76643 1015
rect 76721 969 76767 1015
rect 76845 969 76891 1015
rect 76969 969 77015 1015
rect 77093 969 77139 1015
rect 77217 969 77263 1015
rect 77341 969 77387 1015
rect 77465 969 77511 1015
rect 77589 969 77635 1015
rect 77713 969 77759 1015
rect 77837 969 77883 1015
rect 77961 969 78007 1015
rect 78085 969 78131 1015
rect 78209 969 78255 1015
rect 78333 969 78379 1015
rect 78457 969 78503 1015
rect 78581 969 78627 1015
rect 78705 969 78751 1015
rect 78829 969 78875 1015
rect 78953 969 78999 1015
rect 79077 969 79123 1015
rect 79201 969 79247 1015
rect 79325 969 79371 1015
rect 79449 969 79495 1015
rect 79573 969 79619 1015
rect 79697 969 79743 1015
rect 79821 969 79867 1015
rect 79945 969 79991 1015
rect 80069 969 80115 1015
rect 80193 969 80239 1015
rect 80317 969 80363 1015
rect 80441 969 80487 1015
rect 80565 969 80611 1015
rect 80689 969 80735 1015
rect 80813 969 80859 1015
rect 80937 969 80983 1015
rect 81061 969 81107 1015
rect 81185 969 81231 1015
rect 81309 969 81355 1015
rect 81433 969 81479 1015
rect 81557 969 81603 1015
rect 81681 969 81727 1015
rect 81805 969 81851 1015
rect 81929 969 81975 1015
rect 82053 969 82099 1015
rect 82177 969 82223 1015
rect 82301 969 82347 1015
rect 82425 969 82471 1015
rect 82549 969 82595 1015
rect 82673 969 82719 1015
rect 82797 969 82843 1015
rect 82921 969 82967 1015
rect 83045 969 83091 1015
rect 83169 969 83215 1015
rect 83293 969 83339 1015
rect 83417 969 83463 1015
rect 83541 969 83587 1015
rect 83665 969 83711 1015
rect 83789 969 83835 1015
rect 83913 969 83959 1015
rect 84037 969 84083 1015
rect 84161 969 84207 1015
rect 84285 969 84331 1015
rect 84409 969 84455 1015
rect 84533 969 84579 1015
rect 84657 969 84703 1015
rect 84781 969 84827 1015
rect 84905 969 84951 1015
rect 85029 969 85075 1015
rect 85153 969 85199 1015
rect 85277 969 85323 1015
rect 85401 969 85447 1015
rect 85525 969 85571 1015
rect 85649 969 85695 1015
rect 89 845 135 891
rect 213 845 259 891
rect 337 845 383 891
rect 461 845 507 891
rect 585 845 631 891
rect 709 845 755 891
rect 833 845 879 891
rect 957 845 1003 891
rect 1081 845 1127 891
rect 1205 845 1251 891
rect 1329 845 1375 891
rect 1453 845 1499 891
rect 1577 845 1623 891
rect 1701 845 1747 891
rect 1825 845 1871 891
rect 1949 845 1995 891
rect 2073 845 2119 891
rect 2197 845 2243 891
rect 2321 845 2367 891
rect 2445 845 2491 891
rect 2569 845 2615 891
rect 2693 845 2739 891
rect 2817 845 2863 891
rect 2941 845 2987 891
rect 3065 845 3111 891
rect 3189 845 3235 891
rect 3313 845 3359 891
rect 3437 845 3483 891
rect 3561 845 3607 891
rect 3685 845 3731 891
rect 3809 845 3855 891
rect 3933 845 3979 891
rect 4057 845 4103 891
rect 4181 845 4227 891
rect 4305 845 4351 891
rect 4429 845 4475 891
rect 4553 845 4599 891
rect 4677 845 4723 891
rect 4801 845 4847 891
rect 4925 845 4971 891
rect 5049 845 5095 891
rect 5173 845 5219 891
rect 5297 845 5343 891
rect 5421 845 5467 891
rect 5545 845 5591 891
rect 5669 845 5715 891
rect 5793 845 5839 891
rect 5917 845 5963 891
rect 6041 845 6087 891
rect 6165 845 6211 891
rect 6289 845 6335 891
rect 6413 845 6459 891
rect 6537 845 6583 891
rect 6661 845 6707 891
rect 6785 845 6831 891
rect 6909 845 6955 891
rect 7033 845 7079 891
rect 7157 845 7203 891
rect 7281 845 7327 891
rect 7405 845 7451 891
rect 7529 845 7575 891
rect 7653 845 7699 891
rect 7777 845 7823 891
rect 7901 845 7947 891
rect 8025 845 8071 891
rect 8149 845 8195 891
rect 8273 845 8319 891
rect 8397 845 8443 891
rect 8521 845 8567 891
rect 8645 845 8691 891
rect 8769 845 8815 891
rect 8893 845 8939 891
rect 9017 845 9063 891
rect 9141 845 9187 891
rect 9265 845 9311 891
rect 9389 845 9435 891
rect 9513 845 9559 891
rect 9637 845 9683 891
rect 9761 845 9807 891
rect 9885 845 9931 891
rect 10009 845 10055 891
rect 10133 845 10179 891
rect 10257 845 10303 891
rect 10381 845 10427 891
rect 10505 845 10551 891
rect 10629 845 10675 891
rect 10753 845 10799 891
rect 10877 845 10923 891
rect 11001 845 11047 891
rect 11125 845 11171 891
rect 11249 845 11295 891
rect 11373 845 11419 891
rect 11497 845 11543 891
rect 11621 845 11667 891
rect 11745 845 11791 891
rect 11869 845 11915 891
rect 11993 845 12039 891
rect 12117 845 12163 891
rect 12241 845 12287 891
rect 12365 845 12411 891
rect 12489 845 12535 891
rect 12613 845 12659 891
rect 12737 845 12783 891
rect 12861 845 12907 891
rect 12985 845 13031 891
rect 13109 845 13155 891
rect 13233 845 13279 891
rect 13357 845 13403 891
rect 13481 845 13527 891
rect 13605 845 13651 891
rect 13729 845 13775 891
rect 13853 845 13899 891
rect 13977 845 14023 891
rect 14101 845 14147 891
rect 14225 845 14271 891
rect 14349 845 14395 891
rect 14473 845 14519 891
rect 14597 845 14643 891
rect 14721 845 14767 891
rect 14845 845 14891 891
rect 14969 845 15015 891
rect 15093 845 15139 891
rect 15217 845 15263 891
rect 15341 845 15387 891
rect 15465 845 15511 891
rect 15589 845 15635 891
rect 15713 845 15759 891
rect 15837 845 15883 891
rect 15961 845 16007 891
rect 16085 845 16131 891
rect 16209 845 16255 891
rect 16333 845 16379 891
rect 16457 845 16503 891
rect 16581 845 16627 891
rect 16705 845 16751 891
rect 16829 845 16875 891
rect 16953 845 16999 891
rect 17077 845 17123 891
rect 17201 845 17247 891
rect 17325 845 17371 891
rect 17449 845 17495 891
rect 17573 845 17619 891
rect 17697 845 17743 891
rect 17821 845 17867 891
rect 17945 845 17991 891
rect 18069 845 18115 891
rect 18193 845 18239 891
rect 18317 845 18363 891
rect 18441 845 18487 891
rect 18565 845 18611 891
rect 18689 845 18735 891
rect 18813 845 18859 891
rect 18937 845 18983 891
rect 19061 845 19107 891
rect 19185 845 19231 891
rect 19309 845 19355 891
rect 19433 845 19479 891
rect 19557 845 19603 891
rect 19681 845 19727 891
rect 19805 845 19851 891
rect 19929 845 19975 891
rect 20053 845 20099 891
rect 20177 845 20223 891
rect 20301 845 20347 891
rect 20425 845 20471 891
rect 20549 845 20595 891
rect 20673 845 20719 891
rect 20797 845 20843 891
rect 20921 845 20967 891
rect 21045 845 21091 891
rect 21169 845 21215 891
rect 21293 845 21339 891
rect 21417 845 21463 891
rect 21541 845 21587 891
rect 21665 845 21711 891
rect 21789 845 21835 891
rect 21913 845 21959 891
rect 22037 845 22083 891
rect 22161 845 22207 891
rect 22285 845 22331 891
rect 22409 845 22455 891
rect 22533 845 22579 891
rect 22657 845 22703 891
rect 22781 845 22827 891
rect 22905 845 22951 891
rect 23029 845 23075 891
rect 23153 845 23199 891
rect 23277 845 23323 891
rect 23401 845 23447 891
rect 23525 845 23571 891
rect 23649 845 23695 891
rect 23773 845 23819 891
rect 23897 845 23943 891
rect 24021 845 24067 891
rect 24145 845 24191 891
rect 24269 845 24315 891
rect 24393 845 24439 891
rect 24517 845 24563 891
rect 24641 845 24687 891
rect 24765 845 24811 891
rect 24889 845 24935 891
rect 25013 845 25059 891
rect 25137 845 25183 891
rect 25261 845 25307 891
rect 25385 845 25431 891
rect 25509 845 25555 891
rect 25633 845 25679 891
rect 25757 845 25803 891
rect 25881 845 25927 891
rect 26005 845 26051 891
rect 26129 845 26175 891
rect 26253 845 26299 891
rect 26377 845 26423 891
rect 26501 845 26547 891
rect 26625 845 26671 891
rect 26749 845 26795 891
rect 26873 845 26919 891
rect 26997 845 27043 891
rect 27121 845 27167 891
rect 27245 845 27291 891
rect 27369 845 27415 891
rect 27493 845 27539 891
rect 27617 845 27663 891
rect 27741 845 27787 891
rect 27865 845 27911 891
rect 27989 845 28035 891
rect 28113 845 28159 891
rect 28237 845 28283 891
rect 28361 845 28407 891
rect 28485 845 28531 891
rect 28609 845 28655 891
rect 28733 845 28779 891
rect 28857 845 28903 891
rect 28981 845 29027 891
rect 29105 845 29151 891
rect 29229 845 29275 891
rect 29353 845 29399 891
rect 29477 845 29523 891
rect 29601 845 29647 891
rect 29725 845 29771 891
rect 29849 845 29895 891
rect 29973 845 30019 891
rect 30097 845 30143 891
rect 30221 845 30267 891
rect 30345 845 30391 891
rect 30469 845 30515 891
rect 30593 845 30639 891
rect 30717 845 30763 891
rect 30841 845 30887 891
rect 30965 845 31011 891
rect 31089 845 31135 891
rect 31213 845 31259 891
rect 31337 845 31383 891
rect 31461 845 31507 891
rect 31585 845 31631 891
rect 31709 845 31755 891
rect 31833 845 31879 891
rect 31957 845 32003 891
rect 32081 845 32127 891
rect 32205 845 32251 891
rect 32329 845 32375 891
rect 32453 845 32499 891
rect 32577 845 32623 891
rect 32701 845 32747 891
rect 32825 845 32871 891
rect 32949 845 32995 891
rect 33073 845 33119 891
rect 33197 845 33243 891
rect 33321 845 33367 891
rect 33445 845 33491 891
rect 33569 845 33615 891
rect 33693 845 33739 891
rect 33817 845 33863 891
rect 33941 845 33987 891
rect 34065 845 34111 891
rect 34189 845 34235 891
rect 34313 845 34359 891
rect 34437 845 34483 891
rect 34561 845 34607 891
rect 34685 845 34731 891
rect 34809 845 34855 891
rect 34933 845 34979 891
rect 35057 845 35103 891
rect 35181 845 35227 891
rect 35305 845 35351 891
rect 35429 845 35475 891
rect 35553 845 35599 891
rect 35677 845 35723 891
rect 35801 845 35847 891
rect 35925 845 35971 891
rect 36049 845 36095 891
rect 36173 845 36219 891
rect 36297 845 36343 891
rect 36421 845 36467 891
rect 36545 845 36591 891
rect 36669 845 36715 891
rect 36793 845 36839 891
rect 36917 845 36963 891
rect 37041 845 37087 891
rect 37165 845 37211 891
rect 37289 845 37335 891
rect 37413 845 37459 891
rect 37537 845 37583 891
rect 37661 845 37707 891
rect 37785 845 37831 891
rect 37909 845 37955 891
rect 38033 845 38079 891
rect 38157 845 38203 891
rect 38281 845 38327 891
rect 38405 845 38451 891
rect 38529 845 38575 891
rect 38653 845 38699 891
rect 38777 845 38823 891
rect 38901 845 38947 891
rect 39025 845 39071 891
rect 39149 845 39195 891
rect 39273 845 39319 891
rect 39397 845 39443 891
rect 39521 845 39567 891
rect 39645 845 39691 891
rect 39769 845 39815 891
rect 39893 845 39939 891
rect 40017 845 40063 891
rect 40141 845 40187 891
rect 40265 845 40311 891
rect 40389 845 40435 891
rect 40513 845 40559 891
rect 40637 845 40683 891
rect 40761 845 40807 891
rect 40885 845 40931 891
rect 41009 845 41055 891
rect 41133 845 41179 891
rect 41257 845 41303 891
rect 41381 845 41427 891
rect 41505 845 41551 891
rect 41629 845 41675 891
rect 41753 845 41799 891
rect 41877 845 41923 891
rect 42001 845 42047 891
rect 42125 845 42171 891
rect 42249 845 42295 891
rect 42373 845 42419 891
rect 42497 845 42543 891
rect 42621 845 42667 891
rect 42745 845 42791 891
rect 42869 845 42915 891
rect 42993 845 43039 891
rect 43117 845 43163 891
rect 43241 845 43287 891
rect 43365 845 43411 891
rect 43489 845 43535 891
rect 43613 845 43659 891
rect 43737 845 43783 891
rect 43861 845 43907 891
rect 43985 845 44031 891
rect 44109 845 44155 891
rect 44233 845 44279 891
rect 44357 845 44403 891
rect 44481 845 44527 891
rect 44605 845 44651 891
rect 44729 845 44775 891
rect 44853 845 44899 891
rect 44977 845 45023 891
rect 45101 845 45147 891
rect 45225 845 45271 891
rect 45349 845 45395 891
rect 45473 845 45519 891
rect 45597 845 45643 891
rect 45721 845 45767 891
rect 45845 845 45891 891
rect 45969 845 46015 891
rect 46093 845 46139 891
rect 46217 845 46263 891
rect 46341 845 46387 891
rect 46465 845 46511 891
rect 46589 845 46635 891
rect 46713 845 46759 891
rect 46837 845 46883 891
rect 46961 845 47007 891
rect 47085 845 47131 891
rect 47209 845 47255 891
rect 47333 845 47379 891
rect 47457 845 47503 891
rect 47581 845 47627 891
rect 47705 845 47751 891
rect 47829 845 47875 891
rect 47953 845 47999 891
rect 48077 845 48123 891
rect 48201 845 48247 891
rect 48325 845 48371 891
rect 48449 845 48495 891
rect 48573 845 48619 891
rect 48697 845 48743 891
rect 48821 845 48867 891
rect 48945 845 48991 891
rect 49069 845 49115 891
rect 49193 845 49239 891
rect 49317 845 49363 891
rect 49441 845 49487 891
rect 49565 845 49611 891
rect 49689 845 49735 891
rect 49813 845 49859 891
rect 49937 845 49983 891
rect 50061 845 50107 891
rect 50185 845 50231 891
rect 50309 845 50355 891
rect 50433 845 50479 891
rect 50557 845 50603 891
rect 50681 845 50727 891
rect 50805 845 50851 891
rect 50929 845 50975 891
rect 51053 845 51099 891
rect 51177 845 51223 891
rect 51301 845 51347 891
rect 51425 845 51471 891
rect 51549 845 51595 891
rect 51673 845 51719 891
rect 51797 845 51843 891
rect 51921 845 51967 891
rect 52045 845 52091 891
rect 52169 845 52215 891
rect 52293 845 52339 891
rect 52417 845 52463 891
rect 52541 845 52587 891
rect 52665 845 52711 891
rect 52789 845 52835 891
rect 52913 845 52959 891
rect 53037 845 53083 891
rect 53161 845 53207 891
rect 53285 845 53331 891
rect 53409 845 53455 891
rect 53533 845 53579 891
rect 53657 845 53703 891
rect 53781 845 53827 891
rect 53905 845 53951 891
rect 54029 845 54075 891
rect 54153 845 54199 891
rect 54277 845 54323 891
rect 54401 845 54447 891
rect 54525 845 54571 891
rect 54649 845 54695 891
rect 54773 845 54819 891
rect 54897 845 54943 891
rect 55021 845 55067 891
rect 55145 845 55191 891
rect 55269 845 55315 891
rect 55393 845 55439 891
rect 55517 845 55563 891
rect 55641 845 55687 891
rect 55765 845 55811 891
rect 55889 845 55935 891
rect 56013 845 56059 891
rect 56137 845 56183 891
rect 56261 845 56307 891
rect 56385 845 56431 891
rect 56509 845 56555 891
rect 56633 845 56679 891
rect 56757 845 56803 891
rect 56881 845 56927 891
rect 57005 845 57051 891
rect 57129 845 57175 891
rect 57253 845 57299 891
rect 57377 845 57423 891
rect 57501 845 57547 891
rect 57625 845 57671 891
rect 57749 845 57795 891
rect 57873 845 57919 891
rect 57997 845 58043 891
rect 58121 845 58167 891
rect 58245 845 58291 891
rect 58369 845 58415 891
rect 58493 845 58539 891
rect 58617 845 58663 891
rect 58741 845 58787 891
rect 58865 845 58911 891
rect 58989 845 59035 891
rect 59113 845 59159 891
rect 59237 845 59283 891
rect 59361 845 59407 891
rect 59485 845 59531 891
rect 59609 845 59655 891
rect 59733 845 59779 891
rect 59857 845 59903 891
rect 59981 845 60027 891
rect 60105 845 60151 891
rect 60229 845 60275 891
rect 60353 845 60399 891
rect 60477 845 60523 891
rect 60601 845 60647 891
rect 60725 845 60771 891
rect 60849 845 60895 891
rect 60973 845 61019 891
rect 61097 845 61143 891
rect 61221 845 61267 891
rect 61345 845 61391 891
rect 61469 845 61515 891
rect 61593 845 61639 891
rect 61717 845 61763 891
rect 61841 845 61887 891
rect 61965 845 62011 891
rect 62089 845 62135 891
rect 62213 845 62259 891
rect 62337 845 62383 891
rect 62461 845 62507 891
rect 62585 845 62631 891
rect 62709 845 62755 891
rect 62833 845 62879 891
rect 62957 845 63003 891
rect 63081 845 63127 891
rect 63205 845 63251 891
rect 63329 845 63375 891
rect 63453 845 63499 891
rect 63577 845 63623 891
rect 63701 845 63747 891
rect 63825 845 63871 891
rect 63949 845 63995 891
rect 64073 845 64119 891
rect 64197 845 64243 891
rect 64321 845 64367 891
rect 64445 845 64491 891
rect 64569 845 64615 891
rect 64693 845 64739 891
rect 64817 845 64863 891
rect 64941 845 64987 891
rect 65065 845 65111 891
rect 65189 845 65235 891
rect 65313 845 65359 891
rect 65437 845 65483 891
rect 65561 845 65607 891
rect 65685 845 65731 891
rect 65809 845 65855 891
rect 65933 845 65979 891
rect 66057 845 66103 891
rect 66181 845 66227 891
rect 66305 845 66351 891
rect 66429 845 66475 891
rect 66553 845 66599 891
rect 66677 845 66723 891
rect 66801 845 66847 891
rect 66925 845 66971 891
rect 67049 845 67095 891
rect 67173 845 67219 891
rect 67297 845 67343 891
rect 67421 845 67467 891
rect 67545 845 67591 891
rect 67669 845 67715 891
rect 67793 845 67839 891
rect 67917 845 67963 891
rect 68041 845 68087 891
rect 68165 845 68211 891
rect 68289 845 68335 891
rect 68413 845 68459 891
rect 68537 845 68583 891
rect 68661 845 68707 891
rect 68785 845 68831 891
rect 68909 845 68955 891
rect 69033 845 69079 891
rect 69157 845 69203 891
rect 69281 845 69327 891
rect 69405 845 69451 891
rect 69529 845 69575 891
rect 69653 845 69699 891
rect 69777 845 69823 891
rect 69901 845 69947 891
rect 70025 845 70071 891
rect 70149 845 70195 891
rect 70273 845 70319 891
rect 70397 845 70443 891
rect 70521 845 70567 891
rect 70645 845 70691 891
rect 70769 845 70815 891
rect 70893 845 70939 891
rect 71017 845 71063 891
rect 71141 845 71187 891
rect 71265 845 71311 891
rect 71389 845 71435 891
rect 71513 845 71559 891
rect 71637 845 71683 891
rect 71761 845 71807 891
rect 71885 845 71931 891
rect 72009 845 72055 891
rect 72133 845 72179 891
rect 72257 845 72303 891
rect 72381 845 72427 891
rect 72505 845 72551 891
rect 72629 845 72675 891
rect 72753 845 72799 891
rect 72877 845 72923 891
rect 73001 845 73047 891
rect 73125 845 73171 891
rect 73249 845 73295 891
rect 73373 845 73419 891
rect 73497 845 73543 891
rect 73621 845 73667 891
rect 73745 845 73791 891
rect 73869 845 73915 891
rect 73993 845 74039 891
rect 74117 845 74163 891
rect 74241 845 74287 891
rect 74365 845 74411 891
rect 74489 845 74535 891
rect 74613 845 74659 891
rect 74737 845 74783 891
rect 74861 845 74907 891
rect 74985 845 75031 891
rect 75109 845 75155 891
rect 75233 845 75279 891
rect 75357 845 75403 891
rect 75481 845 75527 891
rect 75605 845 75651 891
rect 75729 845 75775 891
rect 75853 845 75899 891
rect 75977 845 76023 891
rect 76101 845 76147 891
rect 76225 845 76271 891
rect 76349 845 76395 891
rect 76473 845 76519 891
rect 76597 845 76643 891
rect 76721 845 76767 891
rect 76845 845 76891 891
rect 76969 845 77015 891
rect 77093 845 77139 891
rect 77217 845 77263 891
rect 77341 845 77387 891
rect 77465 845 77511 891
rect 77589 845 77635 891
rect 77713 845 77759 891
rect 77837 845 77883 891
rect 77961 845 78007 891
rect 78085 845 78131 891
rect 78209 845 78255 891
rect 78333 845 78379 891
rect 78457 845 78503 891
rect 78581 845 78627 891
rect 78705 845 78751 891
rect 78829 845 78875 891
rect 78953 845 78999 891
rect 79077 845 79123 891
rect 79201 845 79247 891
rect 79325 845 79371 891
rect 79449 845 79495 891
rect 79573 845 79619 891
rect 79697 845 79743 891
rect 79821 845 79867 891
rect 79945 845 79991 891
rect 80069 845 80115 891
rect 80193 845 80239 891
rect 80317 845 80363 891
rect 80441 845 80487 891
rect 80565 845 80611 891
rect 80689 845 80735 891
rect 80813 845 80859 891
rect 80937 845 80983 891
rect 81061 845 81107 891
rect 81185 845 81231 891
rect 81309 845 81355 891
rect 81433 845 81479 891
rect 81557 845 81603 891
rect 81681 845 81727 891
rect 81805 845 81851 891
rect 81929 845 81975 891
rect 82053 845 82099 891
rect 82177 845 82223 891
rect 82301 845 82347 891
rect 82425 845 82471 891
rect 82549 845 82595 891
rect 82673 845 82719 891
rect 82797 845 82843 891
rect 82921 845 82967 891
rect 83045 845 83091 891
rect 83169 845 83215 891
rect 83293 845 83339 891
rect 83417 845 83463 891
rect 83541 845 83587 891
rect 83665 845 83711 891
rect 83789 845 83835 891
rect 83913 845 83959 891
rect 84037 845 84083 891
rect 84161 845 84207 891
rect 84285 845 84331 891
rect 84409 845 84455 891
rect 84533 845 84579 891
rect 84657 845 84703 891
rect 84781 845 84827 891
rect 84905 845 84951 891
rect 85029 845 85075 891
rect 85153 845 85199 891
rect 85277 845 85323 891
rect 85401 845 85447 891
rect 85525 845 85571 891
rect 85649 845 85695 891
rect 89 721 135 767
rect 213 721 259 767
rect 337 721 383 767
rect 461 721 507 767
rect 585 721 631 767
rect 709 721 755 767
rect 833 721 879 767
rect 957 721 1003 767
rect 1081 721 1127 767
rect 1205 721 1251 767
rect 1329 721 1375 767
rect 1453 721 1499 767
rect 1577 721 1623 767
rect 1701 721 1747 767
rect 1825 721 1871 767
rect 1949 721 1995 767
rect 2073 721 2119 767
rect 2197 721 2243 767
rect 2321 721 2367 767
rect 2445 721 2491 767
rect 2569 721 2615 767
rect 2693 721 2739 767
rect 2817 721 2863 767
rect 2941 721 2987 767
rect 3065 721 3111 767
rect 3189 721 3235 767
rect 3313 721 3359 767
rect 3437 721 3483 767
rect 3561 721 3607 767
rect 3685 721 3731 767
rect 3809 721 3855 767
rect 3933 721 3979 767
rect 4057 721 4103 767
rect 4181 721 4227 767
rect 4305 721 4351 767
rect 4429 721 4475 767
rect 4553 721 4599 767
rect 4677 721 4723 767
rect 4801 721 4847 767
rect 4925 721 4971 767
rect 5049 721 5095 767
rect 5173 721 5219 767
rect 5297 721 5343 767
rect 5421 721 5467 767
rect 5545 721 5591 767
rect 5669 721 5715 767
rect 5793 721 5839 767
rect 5917 721 5963 767
rect 6041 721 6087 767
rect 6165 721 6211 767
rect 6289 721 6335 767
rect 6413 721 6459 767
rect 6537 721 6583 767
rect 6661 721 6707 767
rect 6785 721 6831 767
rect 6909 721 6955 767
rect 7033 721 7079 767
rect 7157 721 7203 767
rect 7281 721 7327 767
rect 7405 721 7451 767
rect 7529 721 7575 767
rect 7653 721 7699 767
rect 7777 721 7823 767
rect 7901 721 7947 767
rect 8025 721 8071 767
rect 8149 721 8195 767
rect 8273 721 8319 767
rect 8397 721 8443 767
rect 8521 721 8567 767
rect 8645 721 8691 767
rect 8769 721 8815 767
rect 8893 721 8939 767
rect 9017 721 9063 767
rect 9141 721 9187 767
rect 9265 721 9311 767
rect 9389 721 9435 767
rect 9513 721 9559 767
rect 9637 721 9683 767
rect 9761 721 9807 767
rect 9885 721 9931 767
rect 10009 721 10055 767
rect 10133 721 10179 767
rect 10257 721 10303 767
rect 10381 721 10427 767
rect 10505 721 10551 767
rect 10629 721 10675 767
rect 10753 721 10799 767
rect 10877 721 10923 767
rect 11001 721 11047 767
rect 11125 721 11171 767
rect 11249 721 11295 767
rect 11373 721 11419 767
rect 11497 721 11543 767
rect 11621 721 11667 767
rect 11745 721 11791 767
rect 11869 721 11915 767
rect 11993 721 12039 767
rect 12117 721 12163 767
rect 12241 721 12287 767
rect 12365 721 12411 767
rect 12489 721 12535 767
rect 12613 721 12659 767
rect 12737 721 12783 767
rect 12861 721 12907 767
rect 12985 721 13031 767
rect 13109 721 13155 767
rect 13233 721 13279 767
rect 13357 721 13403 767
rect 13481 721 13527 767
rect 13605 721 13651 767
rect 13729 721 13775 767
rect 13853 721 13899 767
rect 13977 721 14023 767
rect 14101 721 14147 767
rect 14225 721 14271 767
rect 14349 721 14395 767
rect 14473 721 14519 767
rect 14597 721 14643 767
rect 14721 721 14767 767
rect 14845 721 14891 767
rect 14969 721 15015 767
rect 15093 721 15139 767
rect 15217 721 15263 767
rect 15341 721 15387 767
rect 15465 721 15511 767
rect 15589 721 15635 767
rect 15713 721 15759 767
rect 15837 721 15883 767
rect 15961 721 16007 767
rect 16085 721 16131 767
rect 16209 721 16255 767
rect 16333 721 16379 767
rect 16457 721 16503 767
rect 16581 721 16627 767
rect 16705 721 16751 767
rect 16829 721 16875 767
rect 16953 721 16999 767
rect 17077 721 17123 767
rect 17201 721 17247 767
rect 17325 721 17371 767
rect 17449 721 17495 767
rect 17573 721 17619 767
rect 17697 721 17743 767
rect 17821 721 17867 767
rect 17945 721 17991 767
rect 18069 721 18115 767
rect 18193 721 18239 767
rect 18317 721 18363 767
rect 18441 721 18487 767
rect 18565 721 18611 767
rect 18689 721 18735 767
rect 18813 721 18859 767
rect 18937 721 18983 767
rect 19061 721 19107 767
rect 19185 721 19231 767
rect 19309 721 19355 767
rect 19433 721 19479 767
rect 19557 721 19603 767
rect 19681 721 19727 767
rect 19805 721 19851 767
rect 19929 721 19975 767
rect 20053 721 20099 767
rect 20177 721 20223 767
rect 20301 721 20347 767
rect 20425 721 20471 767
rect 20549 721 20595 767
rect 20673 721 20719 767
rect 20797 721 20843 767
rect 20921 721 20967 767
rect 21045 721 21091 767
rect 21169 721 21215 767
rect 21293 721 21339 767
rect 21417 721 21463 767
rect 21541 721 21587 767
rect 21665 721 21711 767
rect 21789 721 21835 767
rect 21913 721 21959 767
rect 22037 721 22083 767
rect 22161 721 22207 767
rect 22285 721 22331 767
rect 22409 721 22455 767
rect 22533 721 22579 767
rect 22657 721 22703 767
rect 22781 721 22827 767
rect 22905 721 22951 767
rect 23029 721 23075 767
rect 23153 721 23199 767
rect 23277 721 23323 767
rect 23401 721 23447 767
rect 23525 721 23571 767
rect 23649 721 23695 767
rect 23773 721 23819 767
rect 23897 721 23943 767
rect 24021 721 24067 767
rect 24145 721 24191 767
rect 24269 721 24315 767
rect 24393 721 24439 767
rect 24517 721 24563 767
rect 24641 721 24687 767
rect 24765 721 24811 767
rect 24889 721 24935 767
rect 25013 721 25059 767
rect 25137 721 25183 767
rect 25261 721 25307 767
rect 25385 721 25431 767
rect 25509 721 25555 767
rect 25633 721 25679 767
rect 25757 721 25803 767
rect 25881 721 25927 767
rect 26005 721 26051 767
rect 26129 721 26175 767
rect 26253 721 26299 767
rect 26377 721 26423 767
rect 26501 721 26547 767
rect 26625 721 26671 767
rect 26749 721 26795 767
rect 26873 721 26919 767
rect 26997 721 27043 767
rect 27121 721 27167 767
rect 27245 721 27291 767
rect 27369 721 27415 767
rect 27493 721 27539 767
rect 27617 721 27663 767
rect 27741 721 27787 767
rect 27865 721 27911 767
rect 27989 721 28035 767
rect 28113 721 28159 767
rect 28237 721 28283 767
rect 28361 721 28407 767
rect 28485 721 28531 767
rect 28609 721 28655 767
rect 28733 721 28779 767
rect 28857 721 28903 767
rect 28981 721 29027 767
rect 29105 721 29151 767
rect 29229 721 29275 767
rect 29353 721 29399 767
rect 29477 721 29523 767
rect 29601 721 29647 767
rect 29725 721 29771 767
rect 29849 721 29895 767
rect 29973 721 30019 767
rect 30097 721 30143 767
rect 30221 721 30267 767
rect 30345 721 30391 767
rect 30469 721 30515 767
rect 30593 721 30639 767
rect 30717 721 30763 767
rect 30841 721 30887 767
rect 30965 721 31011 767
rect 31089 721 31135 767
rect 31213 721 31259 767
rect 31337 721 31383 767
rect 31461 721 31507 767
rect 31585 721 31631 767
rect 31709 721 31755 767
rect 31833 721 31879 767
rect 31957 721 32003 767
rect 32081 721 32127 767
rect 32205 721 32251 767
rect 32329 721 32375 767
rect 32453 721 32499 767
rect 32577 721 32623 767
rect 32701 721 32747 767
rect 32825 721 32871 767
rect 32949 721 32995 767
rect 33073 721 33119 767
rect 33197 721 33243 767
rect 33321 721 33367 767
rect 33445 721 33491 767
rect 33569 721 33615 767
rect 33693 721 33739 767
rect 33817 721 33863 767
rect 33941 721 33987 767
rect 34065 721 34111 767
rect 34189 721 34235 767
rect 34313 721 34359 767
rect 34437 721 34483 767
rect 34561 721 34607 767
rect 34685 721 34731 767
rect 34809 721 34855 767
rect 34933 721 34979 767
rect 35057 721 35103 767
rect 35181 721 35227 767
rect 35305 721 35351 767
rect 35429 721 35475 767
rect 35553 721 35599 767
rect 35677 721 35723 767
rect 35801 721 35847 767
rect 35925 721 35971 767
rect 36049 721 36095 767
rect 36173 721 36219 767
rect 36297 721 36343 767
rect 36421 721 36467 767
rect 36545 721 36591 767
rect 36669 721 36715 767
rect 36793 721 36839 767
rect 36917 721 36963 767
rect 37041 721 37087 767
rect 37165 721 37211 767
rect 37289 721 37335 767
rect 37413 721 37459 767
rect 37537 721 37583 767
rect 37661 721 37707 767
rect 37785 721 37831 767
rect 37909 721 37955 767
rect 38033 721 38079 767
rect 38157 721 38203 767
rect 38281 721 38327 767
rect 38405 721 38451 767
rect 38529 721 38575 767
rect 38653 721 38699 767
rect 38777 721 38823 767
rect 38901 721 38947 767
rect 39025 721 39071 767
rect 39149 721 39195 767
rect 39273 721 39319 767
rect 39397 721 39443 767
rect 39521 721 39567 767
rect 39645 721 39691 767
rect 39769 721 39815 767
rect 39893 721 39939 767
rect 40017 721 40063 767
rect 40141 721 40187 767
rect 40265 721 40311 767
rect 40389 721 40435 767
rect 40513 721 40559 767
rect 40637 721 40683 767
rect 40761 721 40807 767
rect 40885 721 40931 767
rect 41009 721 41055 767
rect 41133 721 41179 767
rect 41257 721 41303 767
rect 41381 721 41427 767
rect 41505 721 41551 767
rect 41629 721 41675 767
rect 41753 721 41799 767
rect 41877 721 41923 767
rect 42001 721 42047 767
rect 42125 721 42171 767
rect 42249 721 42295 767
rect 42373 721 42419 767
rect 42497 721 42543 767
rect 42621 721 42667 767
rect 42745 721 42791 767
rect 42869 721 42915 767
rect 42993 721 43039 767
rect 43117 721 43163 767
rect 43241 721 43287 767
rect 43365 721 43411 767
rect 43489 721 43535 767
rect 43613 721 43659 767
rect 43737 721 43783 767
rect 43861 721 43907 767
rect 43985 721 44031 767
rect 44109 721 44155 767
rect 44233 721 44279 767
rect 44357 721 44403 767
rect 44481 721 44527 767
rect 44605 721 44651 767
rect 44729 721 44775 767
rect 44853 721 44899 767
rect 44977 721 45023 767
rect 45101 721 45147 767
rect 45225 721 45271 767
rect 45349 721 45395 767
rect 45473 721 45519 767
rect 45597 721 45643 767
rect 45721 721 45767 767
rect 45845 721 45891 767
rect 45969 721 46015 767
rect 46093 721 46139 767
rect 46217 721 46263 767
rect 46341 721 46387 767
rect 46465 721 46511 767
rect 46589 721 46635 767
rect 46713 721 46759 767
rect 46837 721 46883 767
rect 46961 721 47007 767
rect 47085 721 47131 767
rect 47209 721 47255 767
rect 47333 721 47379 767
rect 47457 721 47503 767
rect 47581 721 47627 767
rect 47705 721 47751 767
rect 47829 721 47875 767
rect 47953 721 47999 767
rect 48077 721 48123 767
rect 48201 721 48247 767
rect 48325 721 48371 767
rect 48449 721 48495 767
rect 48573 721 48619 767
rect 48697 721 48743 767
rect 48821 721 48867 767
rect 48945 721 48991 767
rect 49069 721 49115 767
rect 49193 721 49239 767
rect 49317 721 49363 767
rect 49441 721 49487 767
rect 49565 721 49611 767
rect 49689 721 49735 767
rect 49813 721 49859 767
rect 49937 721 49983 767
rect 50061 721 50107 767
rect 50185 721 50231 767
rect 50309 721 50355 767
rect 50433 721 50479 767
rect 50557 721 50603 767
rect 50681 721 50727 767
rect 50805 721 50851 767
rect 50929 721 50975 767
rect 51053 721 51099 767
rect 51177 721 51223 767
rect 51301 721 51347 767
rect 51425 721 51471 767
rect 51549 721 51595 767
rect 51673 721 51719 767
rect 51797 721 51843 767
rect 51921 721 51967 767
rect 52045 721 52091 767
rect 52169 721 52215 767
rect 52293 721 52339 767
rect 52417 721 52463 767
rect 52541 721 52587 767
rect 52665 721 52711 767
rect 52789 721 52835 767
rect 52913 721 52959 767
rect 53037 721 53083 767
rect 53161 721 53207 767
rect 53285 721 53331 767
rect 53409 721 53455 767
rect 53533 721 53579 767
rect 53657 721 53703 767
rect 53781 721 53827 767
rect 53905 721 53951 767
rect 54029 721 54075 767
rect 54153 721 54199 767
rect 54277 721 54323 767
rect 54401 721 54447 767
rect 54525 721 54571 767
rect 54649 721 54695 767
rect 54773 721 54819 767
rect 54897 721 54943 767
rect 55021 721 55067 767
rect 55145 721 55191 767
rect 55269 721 55315 767
rect 55393 721 55439 767
rect 55517 721 55563 767
rect 55641 721 55687 767
rect 55765 721 55811 767
rect 55889 721 55935 767
rect 56013 721 56059 767
rect 56137 721 56183 767
rect 56261 721 56307 767
rect 56385 721 56431 767
rect 56509 721 56555 767
rect 56633 721 56679 767
rect 56757 721 56803 767
rect 56881 721 56927 767
rect 57005 721 57051 767
rect 57129 721 57175 767
rect 57253 721 57299 767
rect 57377 721 57423 767
rect 57501 721 57547 767
rect 57625 721 57671 767
rect 57749 721 57795 767
rect 57873 721 57919 767
rect 57997 721 58043 767
rect 58121 721 58167 767
rect 58245 721 58291 767
rect 58369 721 58415 767
rect 58493 721 58539 767
rect 58617 721 58663 767
rect 58741 721 58787 767
rect 58865 721 58911 767
rect 58989 721 59035 767
rect 59113 721 59159 767
rect 59237 721 59283 767
rect 59361 721 59407 767
rect 59485 721 59531 767
rect 59609 721 59655 767
rect 59733 721 59779 767
rect 59857 721 59903 767
rect 59981 721 60027 767
rect 60105 721 60151 767
rect 60229 721 60275 767
rect 60353 721 60399 767
rect 60477 721 60523 767
rect 60601 721 60647 767
rect 60725 721 60771 767
rect 60849 721 60895 767
rect 60973 721 61019 767
rect 61097 721 61143 767
rect 61221 721 61267 767
rect 61345 721 61391 767
rect 61469 721 61515 767
rect 61593 721 61639 767
rect 61717 721 61763 767
rect 61841 721 61887 767
rect 61965 721 62011 767
rect 62089 721 62135 767
rect 62213 721 62259 767
rect 62337 721 62383 767
rect 62461 721 62507 767
rect 62585 721 62631 767
rect 62709 721 62755 767
rect 62833 721 62879 767
rect 62957 721 63003 767
rect 63081 721 63127 767
rect 63205 721 63251 767
rect 63329 721 63375 767
rect 63453 721 63499 767
rect 63577 721 63623 767
rect 63701 721 63747 767
rect 63825 721 63871 767
rect 63949 721 63995 767
rect 64073 721 64119 767
rect 64197 721 64243 767
rect 64321 721 64367 767
rect 64445 721 64491 767
rect 64569 721 64615 767
rect 64693 721 64739 767
rect 64817 721 64863 767
rect 64941 721 64987 767
rect 65065 721 65111 767
rect 65189 721 65235 767
rect 65313 721 65359 767
rect 65437 721 65483 767
rect 65561 721 65607 767
rect 65685 721 65731 767
rect 65809 721 65855 767
rect 65933 721 65979 767
rect 66057 721 66103 767
rect 66181 721 66227 767
rect 66305 721 66351 767
rect 66429 721 66475 767
rect 66553 721 66599 767
rect 66677 721 66723 767
rect 66801 721 66847 767
rect 66925 721 66971 767
rect 67049 721 67095 767
rect 67173 721 67219 767
rect 67297 721 67343 767
rect 67421 721 67467 767
rect 67545 721 67591 767
rect 67669 721 67715 767
rect 67793 721 67839 767
rect 67917 721 67963 767
rect 68041 721 68087 767
rect 68165 721 68211 767
rect 68289 721 68335 767
rect 68413 721 68459 767
rect 68537 721 68583 767
rect 68661 721 68707 767
rect 68785 721 68831 767
rect 68909 721 68955 767
rect 69033 721 69079 767
rect 69157 721 69203 767
rect 69281 721 69327 767
rect 69405 721 69451 767
rect 69529 721 69575 767
rect 69653 721 69699 767
rect 69777 721 69823 767
rect 69901 721 69947 767
rect 70025 721 70071 767
rect 70149 721 70195 767
rect 70273 721 70319 767
rect 70397 721 70443 767
rect 70521 721 70567 767
rect 70645 721 70691 767
rect 70769 721 70815 767
rect 70893 721 70939 767
rect 71017 721 71063 767
rect 71141 721 71187 767
rect 71265 721 71311 767
rect 71389 721 71435 767
rect 71513 721 71559 767
rect 71637 721 71683 767
rect 71761 721 71807 767
rect 71885 721 71931 767
rect 72009 721 72055 767
rect 72133 721 72179 767
rect 72257 721 72303 767
rect 72381 721 72427 767
rect 72505 721 72551 767
rect 72629 721 72675 767
rect 72753 721 72799 767
rect 72877 721 72923 767
rect 73001 721 73047 767
rect 73125 721 73171 767
rect 73249 721 73295 767
rect 73373 721 73419 767
rect 73497 721 73543 767
rect 73621 721 73667 767
rect 73745 721 73791 767
rect 73869 721 73915 767
rect 73993 721 74039 767
rect 74117 721 74163 767
rect 74241 721 74287 767
rect 74365 721 74411 767
rect 74489 721 74535 767
rect 74613 721 74659 767
rect 74737 721 74783 767
rect 74861 721 74907 767
rect 74985 721 75031 767
rect 75109 721 75155 767
rect 75233 721 75279 767
rect 75357 721 75403 767
rect 75481 721 75527 767
rect 75605 721 75651 767
rect 75729 721 75775 767
rect 75853 721 75899 767
rect 75977 721 76023 767
rect 76101 721 76147 767
rect 76225 721 76271 767
rect 76349 721 76395 767
rect 76473 721 76519 767
rect 76597 721 76643 767
rect 76721 721 76767 767
rect 76845 721 76891 767
rect 76969 721 77015 767
rect 77093 721 77139 767
rect 77217 721 77263 767
rect 77341 721 77387 767
rect 77465 721 77511 767
rect 77589 721 77635 767
rect 77713 721 77759 767
rect 77837 721 77883 767
rect 77961 721 78007 767
rect 78085 721 78131 767
rect 78209 721 78255 767
rect 78333 721 78379 767
rect 78457 721 78503 767
rect 78581 721 78627 767
rect 78705 721 78751 767
rect 78829 721 78875 767
rect 78953 721 78999 767
rect 79077 721 79123 767
rect 79201 721 79247 767
rect 79325 721 79371 767
rect 79449 721 79495 767
rect 79573 721 79619 767
rect 79697 721 79743 767
rect 79821 721 79867 767
rect 79945 721 79991 767
rect 80069 721 80115 767
rect 80193 721 80239 767
rect 80317 721 80363 767
rect 80441 721 80487 767
rect 80565 721 80611 767
rect 80689 721 80735 767
rect 80813 721 80859 767
rect 80937 721 80983 767
rect 81061 721 81107 767
rect 81185 721 81231 767
rect 81309 721 81355 767
rect 81433 721 81479 767
rect 81557 721 81603 767
rect 81681 721 81727 767
rect 81805 721 81851 767
rect 81929 721 81975 767
rect 82053 721 82099 767
rect 82177 721 82223 767
rect 82301 721 82347 767
rect 82425 721 82471 767
rect 82549 721 82595 767
rect 82673 721 82719 767
rect 82797 721 82843 767
rect 82921 721 82967 767
rect 83045 721 83091 767
rect 83169 721 83215 767
rect 83293 721 83339 767
rect 83417 721 83463 767
rect 83541 721 83587 767
rect 83665 721 83711 767
rect 83789 721 83835 767
rect 83913 721 83959 767
rect 84037 721 84083 767
rect 84161 721 84207 767
rect 84285 721 84331 767
rect 84409 721 84455 767
rect 84533 721 84579 767
rect 84657 721 84703 767
rect 84781 721 84827 767
rect 84905 721 84951 767
rect 85029 721 85075 767
rect 85153 721 85199 767
rect 85277 721 85323 767
rect 85401 721 85447 767
rect 85525 721 85571 767
rect 85649 721 85695 767
rect 89 597 135 643
rect 213 597 259 643
rect 337 597 383 643
rect 461 597 507 643
rect 585 597 631 643
rect 709 597 755 643
rect 833 597 879 643
rect 957 597 1003 643
rect 1081 597 1127 643
rect 1205 597 1251 643
rect 1329 597 1375 643
rect 1453 597 1499 643
rect 1577 597 1623 643
rect 1701 597 1747 643
rect 1825 597 1871 643
rect 1949 597 1995 643
rect 2073 597 2119 643
rect 2197 597 2243 643
rect 2321 597 2367 643
rect 2445 597 2491 643
rect 2569 597 2615 643
rect 2693 597 2739 643
rect 2817 597 2863 643
rect 2941 597 2987 643
rect 3065 597 3111 643
rect 3189 597 3235 643
rect 3313 597 3359 643
rect 3437 597 3483 643
rect 3561 597 3607 643
rect 3685 597 3731 643
rect 3809 597 3855 643
rect 3933 597 3979 643
rect 4057 597 4103 643
rect 4181 597 4227 643
rect 4305 597 4351 643
rect 4429 597 4475 643
rect 4553 597 4599 643
rect 4677 597 4723 643
rect 4801 597 4847 643
rect 4925 597 4971 643
rect 5049 597 5095 643
rect 5173 597 5219 643
rect 5297 597 5343 643
rect 5421 597 5467 643
rect 5545 597 5591 643
rect 5669 597 5715 643
rect 5793 597 5839 643
rect 5917 597 5963 643
rect 6041 597 6087 643
rect 6165 597 6211 643
rect 6289 597 6335 643
rect 6413 597 6459 643
rect 6537 597 6583 643
rect 6661 597 6707 643
rect 6785 597 6831 643
rect 6909 597 6955 643
rect 7033 597 7079 643
rect 7157 597 7203 643
rect 7281 597 7327 643
rect 7405 597 7451 643
rect 7529 597 7575 643
rect 7653 597 7699 643
rect 7777 597 7823 643
rect 7901 597 7947 643
rect 8025 597 8071 643
rect 8149 597 8195 643
rect 8273 597 8319 643
rect 8397 597 8443 643
rect 8521 597 8567 643
rect 8645 597 8691 643
rect 8769 597 8815 643
rect 8893 597 8939 643
rect 9017 597 9063 643
rect 9141 597 9187 643
rect 9265 597 9311 643
rect 9389 597 9435 643
rect 9513 597 9559 643
rect 9637 597 9683 643
rect 9761 597 9807 643
rect 9885 597 9931 643
rect 10009 597 10055 643
rect 10133 597 10179 643
rect 10257 597 10303 643
rect 10381 597 10427 643
rect 10505 597 10551 643
rect 10629 597 10675 643
rect 10753 597 10799 643
rect 10877 597 10923 643
rect 11001 597 11047 643
rect 11125 597 11171 643
rect 11249 597 11295 643
rect 11373 597 11419 643
rect 11497 597 11543 643
rect 11621 597 11667 643
rect 11745 597 11791 643
rect 11869 597 11915 643
rect 11993 597 12039 643
rect 12117 597 12163 643
rect 12241 597 12287 643
rect 12365 597 12411 643
rect 12489 597 12535 643
rect 12613 597 12659 643
rect 12737 597 12783 643
rect 12861 597 12907 643
rect 12985 597 13031 643
rect 13109 597 13155 643
rect 13233 597 13279 643
rect 13357 597 13403 643
rect 13481 597 13527 643
rect 13605 597 13651 643
rect 13729 597 13775 643
rect 13853 597 13899 643
rect 13977 597 14023 643
rect 14101 597 14147 643
rect 14225 597 14271 643
rect 14349 597 14395 643
rect 14473 597 14519 643
rect 14597 597 14643 643
rect 14721 597 14767 643
rect 14845 597 14891 643
rect 14969 597 15015 643
rect 15093 597 15139 643
rect 15217 597 15263 643
rect 15341 597 15387 643
rect 15465 597 15511 643
rect 15589 597 15635 643
rect 15713 597 15759 643
rect 15837 597 15883 643
rect 15961 597 16007 643
rect 16085 597 16131 643
rect 16209 597 16255 643
rect 16333 597 16379 643
rect 16457 597 16503 643
rect 16581 597 16627 643
rect 16705 597 16751 643
rect 16829 597 16875 643
rect 16953 597 16999 643
rect 17077 597 17123 643
rect 17201 597 17247 643
rect 17325 597 17371 643
rect 17449 597 17495 643
rect 17573 597 17619 643
rect 17697 597 17743 643
rect 17821 597 17867 643
rect 17945 597 17991 643
rect 18069 597 18115 643
rect 18193 597 18239 643
rect 18317 597 18363 643
rect 18441 597 18487 643
rect 18565 597 18611 643
rect 18689 597 18735 643
rect 18813 597 18859 643
rect 18937 597 18983 643
rect 19061 597 19107 643
rect 19185 597 19231 643
rect 19309 597 19355 643
rect 19433 597 19479 643
rect 19557 597 19603 643
rect 19681 597 19727 643
rect 19805 597 19851 643
rect 19929 597 19975 643
rect 20053 597 20099 643
rect 20177 597 20223 643
rect 20301 597 20347 643
rect 20425 597 20471 643
rect 20549 597 20595 643
rect 20673 597 20719 643
rect 20797 597 20843 643
rect 20921 597 20967 643
rect 21045 597 21091 643
rect 21169 597 21215 643
rect 21293 597 21339 643
rect 21417 597 21463 643
rect 21541 597 21587 643
rect 21665 597 21711 643
rect 21789 597 21835 643
rect 21913 597 21959 643
rect 22037 597 22083 643
rect 22161 597 22207 643
rect 22285 597 22331 643
rect 22409 597 22455 643
rect 22533 597 22579 643
rect 22657 597 22703 643
rect 22781 597 22827 643
rect 22905 597 22951 643
rect 23029 597 23075 643
rect 23153 597 23199 643
rect 23277 597 23323 643
rect 23401 597 23447 643
rect 23525 597 23571 643
rect 23649 597 23695 643
rect 23773 597 23819 643
rect 23897 597 23943 643
rect 24021 597 24067 643
rect 24145 597 24191 643
rect 24269 597 24315 643
rect 24393 597 24439 643
rect 24517 597 24563 643
rect 24641 597 24687 643
rect 24765 597 24811 643
rect 24889 597 24935 643
rect 25013 597 25059 643
rect 25137 597 25183 643
rect 25261 597 25307 643
rect 25385 597 25431 643
rect 25509 597 25555 643
rect 25633 597 25679 643
rect 25757 597 25803 643
rect 25881 597 25927 643
rect 26005 597 26051 643
rect 26129 597 26175 643
rect 26253 597 26299 643
rect 26377 597 26423 643
rect 26501 597 26547 643
rect 26625 597 26671 643
rect 26749 597 26795 643
rect 26873 597 26919 643
rect 26997 597 27043 643
rect 27121 597 27167 643
rect 27245 597 27291 643
rect 27369 597 27415 643
rect 27493 597 27539 643
rect 27617 597 27663 643
rect 27741 597 27787 643
rect 27865 597 27911 643
rect 27989 597 28035 643
rect 28113 597 28159 643
rect 28237 597 28283 643
rect 28361 597 28407 643
rect 28485 597 28531 643
rect 28609 597 28655 643
rect 28733 597 28779 643
rect 28857 597 28903 643
rect 28981 597 29027 643
rect 29105 597 29151 643
rect 29229 597 29275 643
rect 29353 597 29399 643
rect 29477 597 29523 643
rect 29601 597 29647 643
rect 29725 597 29771 643
rect 29849 597 29895 643
rect 29973 597 30019 643
rect 30097 597 30143 643
rect 30221 597 30267 643
rect 30345 597 30391 643
rect 30469 597 30515 643
rect 30593 597 30639 643
rect 30717 597 30763 643
rect 30841 597 30887 643
rect 30965 597 31011 643
rect 31089 597 31135 643
rect 31213 597 31259 643
rect 31337 597 31383 643
rect 31461 597 31507 643
rect 31585 597 31631 643
rect 31709 597 31755 643
rect 31833 597 31879 643
rect 31957 597 32003 643
rect 32081 597 32127 643
rect 32205 597 32251 643
rect 32329 597 32375 643
rect 32453 597 32499 643
rect 32577 597 32623 643
rect 32701 597 32747 643
rect 32825 597 32871 643
rect 32949 597 32995 643
rect 33073 597 33119 643
rect 33197 597 33243 643
rect 33321 597 33367 643
rect 33445 597 33491 643
rect 33569 597 33615 643
rect 33693 597 33739 643
rect 33817 597 33863 643
rect 33941 597 33987 643
rect 34065 597 34111 643
rect 34189 597 34235 643
rect 34313 597 34359 643
rect 34437 597 34483 643
rect 34561 597 34607 643
rect 34685 597 34731 643
rect 34809 597 34855 643
rect 34933 597 34979 643
rect 35057 597 35103 643
rect 35181 597 35227 643
rect 35305 597 35351 643
rect 35429 597 35475 643
rect 35553 597 35599 643
rect 35677 597 35723 643
rect 35801 597 35847 643
rect 35925 597 35971 643
rect 36049 597 36095 643
rect 36173 597 36219 643
rect 36297 597 36343 643
rect 36421 597 36467 643
rect 36545 597 36591 643
rect 36669 597 36715 643
rect 36793 597 36839 643
rect 36917 597 36963 643
rect 37041 597 37087 643
rect 37165 597 37211 643
rect 37289 597 37335 643
rect 37413 597 37459 643
rect 37537 597 37583 643
rect 37661 597 37707 643
rect 37785 597 37831 643
rect 37909 597 37955 643
rect 38033 597 38079 643
rect 38157 597 38203 643
rect 38281 597 38327 643
rect 38405 597 38451 643
rect 38529 597 38575 643
rect 38653 597 38699 643
rect 38777 597 38823 643
rect 38901 597 38947 643
rect 39025 597 39071 643
rect 39149 597 39195 643
rect 39273 597 39319 643
rect 39397 597 39443 643
rect 39521 597 39567 643
rect 39645 597 39691 643
rect 39769 597 39815 643
rect 39893 597 39939 643
rect 40017 597 40063 643
rect 40141 597 40187 643
rect 40265 597 40311 643
rect 40389 597 40435 643
rect 40513 597 40559 643
rect 40637 597 40683 643
rect 40761 597 40807 643
rect 40885 597 40931 643
rect 41009 597 41055 643
rect 41133 597 41179 643
rect 41257 597 41303 643
rect 41381 597 41427 643
rect 41505 597 41551 643
rect 41629 597 41675 643
rect 41753 597 41799 643
rect 41877 597 41923 643
rect 42001 597 42047 643
rect 42125 597 42171 643
rect 42249 597 42295 643
rect 42373 597 42419 643
rect 42497 597 42543 643
rect 42621 597 42667 643
rect 42745 597 42791 643
rect 42869 597 42915 643
rect 42993 597 43039 643
rect 43117 597 43163 643
rect 43241 597 43287 643
rect 43365 597 43411 643
rect 43489 597 43535 643
rect 43613 597 43659 643
rect 43737 597 43783 643
rect 43861 597 43907 643
rect 43985 597 44031 643
rect 44109 597 44155 643
rect 44233 597 44279 643
rect 44357 597 44403 643
rect 44481 597 44527 643
rect 44605 597 44651 643
rect 44729 597 44775 643
rect 44853 597 44899 643
rect 44977 597 45023 643
rect 45101 597 45147 643
rect 45225 597 45271 643
rect 45349 597 45395 643
rect 45473 597 45519 643
rect 45597 597 45643 643
rect 45721 597 45767 643
rect 45845 597 45891 643
rect 45969 597 46015 643
rect 46093 597 46139 643
rect 46217 597 46263 643
rect 46341 597 46387 643
rect 46465 597 46511 643
rect 46589 597 46635 643
rect 46713 597 46759 643
rect 46837 597 46883 643
rect 46961 597 47007 643
rect 47085 597 47131 643
rect 47209 597 47255 643
rect 47333 597 47379 643
rect 47457 597 47503 643
rect 47581 597 47627 643
rect 47705 597 47751 643
rect 47829 597 47875 643
rect 47953 597 47999 643
rect 48077 597 48123 643
rect 48201 597 48247 643
rect 48325 597 48371 643
rect 48449 597 48495 643
rect 48573 597 48619 643
rect 48697 597 48743 643
rect 48821 597 48867 643
rect 48945 597 48991 643
rect 49069 597 49115 643
rect 49193 597 49239 643
rect 49317 597 49363 643
rect 49441 597 49487 643
rect 49565 597 49611 643
rect 49689 597 49735 643
rect 49813 597 49859 643
rect 49937 597 49983 643
rect 50061 597 50107 643
rect 50185 597 50231 643
rect 50309 597 50355 643
rect 50433 597 50479 643
rect 50557 597 50603 643
rect 50681 597 50727 643
rect 50805 597 50851 643
rect 50929 597 50975 643
rect 51053 597 51099 643
rect 51177 597 51223 643
rect 51301 597 51347 643
rect 51425 597 51471 643
rect 51549 597 51595 643
rect 51673 597 51719 643
rect 51797 597 51843 643
rect 51921 597 51967 643
rect 52045 597 52091 643
rect 52169 597 52215 643
rect 52293 597 52339 643
rect 52417 597 52463 643
rect 52541 597 52587 643
rect 52665 597 52711 643
rect 52789 597 52835 643
rect 52913 597 52959 643
rect 53037 597 53083 643
rect 53161 597 53207 643
rect 53285 597 53331 643
rect 53409 597 53455 643
rect 53533 597 53579 643
rect 53657 597 53703 643
rect 53781 597 53827 643
rect 53905 597 53951 643
rect 54029 597 54075 643
rect 54153 597 54199 643
rect 54277 597 54323 643
rect 54401 597 54447 643
rect 54525 597 54571 643
rect 54649 597 54695 643
rect 54773 597 54819 643
rect 54897 597 54943 643
rect 55021 597 55067 643
rect 55145 597 55191 643
rect 55269 597 55315 643
rect 55393 597 55439 643
rect 55517 597 55563 643
rect 55641 597 55687 643
rect 55765 597 55811 643
rect 55889 597 55935 643
rect 56013 597 56059 643
rect 56137 597 56183 643
rect 56261 597 56307 643
rect 56385 597 56431 643
rect 56509 597 56555 643
rect 56633 597 56679 643
rect 56757 597 56803 643
rect 56881 597 56927 643
rect 57005 597 57051 643
rect 57129 597 57175 643
rect 57253 597 57299 643
rect 57377 597 57423 643
rect 57501 597 57547 643
rect 57625 597 57671 643
rect 57749 597 57795 643
rect 57873 597 57919 643
rect 57997 597 58043 643
rect 58121 597 58167 643
rect 58245 597 58291 643
rect 58369 597 58415 643
rect 58493 597 58539 643
rect 58617 597 58663 643
rect 58741 597 58787 643
rect 58865 597 58911 643
rect 58989 597 59035 643
rect 59113 597 59159 643
rect 59237 597 59283 643
rect 59361 597 59407 643
rect 59485 597 59531 643
rect 59609 597 59655 643
rect 59733 597 59779 643
rect 59857 597 59903 643
rect 59981 597 60027 643
rect 60105 597 60151 643
rect 60229 597 60275 643
rect 60353 597 60399 643
rect 60477 597 60523 643
rect 60601 597 60647 643
rect 60725 597 60771 643
rect 60849 597 60895 643
rect 60973 597 61019 643
rect 61097 597 61143 643
rect 61221 597 61267 643
rect 61345 597 61391 643
rect 61469 597 61515 643
rect 61593 597 61639 643
rect 61717 597 61763 643
rect 61841 597 61887 643
rect 61965 597 62011 643
rect 62089 597 62135 643
rect 62213 597 62259 643
rect 62337 597 62383 643
rect 62461 597 62507 643
rect 62585 597 62631 643
rect 62709 597 62755 643
rect 62833 597 62879 643
rect 62957 597 63003 643
rect 63081 597 63127 643
rect 63205 597 63251 643
rect 63329 597 63375 643
rect 63453 597 63499 643
rect 63577 597 63623 643
rect 63701 597 63747 643
rect 63825 597 63871 643
rect 63949 597 63995 643
rect 64073 597 64119 643
rect 64197 597 64243 643
rect 64321 597 64367 643
rect 64445 597 64491 643
rect 64569 597 64615 643
rect 64693 597 64739 643
rect 64817 597 64863 643
rect 64941 597 64987 643
rect 65065 597 65111 643
rect 65189 597 65235 643
rect 65313 597 65359 643
rect 65437 597 65483 643
rect 65561 597 65607 643
rect 65685 597 65731 643
rect 65809 597 65855 643
rect 65933 597 65979 643
rect 66057 597 66103 643
rect 66181 597 66227 643
rect 66305 597 66351 643
rect 66429 597 66475 643
rect 66553 597 66599 643
rect 66677 597 66723 643
rect 66801 597 66847 643
rect 66925 597 66971 643
rect 67049 597 67095 643
rect 67173 597 67219 643
rect 67297 597 67343 643
rect 67421 597 67467 643
rect 67545 597 67591 643
rect 67669 597 67715 643
rect 67793 597 67839 643
rect 67917 597 67963 643
rect 68041 597 68087 643
rect 68165 597 68211 643
rect 68289 597 68335 643
rect 68413 597 68459 643
rect 68537 597 68583 643
rect 68661 597 68707 643
rect 68785 597 68831 643
rect 68909 597 68955 643
rect 69033 597 69079 643
rect 69157 597 69203 643
rect 69281 597 69327 643
rect 69405 597 69451 643
rect 69529 597 69575 643
rect 69653 597 69699 643
rect 69777 597 69823 643
rect 69901 597 69947 643
rect 70025 597 70071 643
rect 70149 597 70195 643
rect 70273 597 70319 643
rect 70397 597 70443 643
rect 70521 597 70567 643
rect 70645 597 70691 643
rect 70769 597 70815 643
rect 70893 597 70939 643
rect 71017 597 71063 643
rect 71141 597 71187 643
rect 71265 597 71311 643
rect 71389 597 71435 643
rect 71513 597 71559 643
rect 71637 597 71683 643
rect 71761 597 71807 643
rect 71885 597 71931 643
rect 72009 597 72055 643
rect 72133 597 72179 643
rect 72257 597 72303 643
rect 72381 597 72427 643
rect 72505 597 72551 643
rect 72629 597 72675 643
rect 72753 597 72799 643
rect 72877 597 72923 643
rect 73001 597 73047 643
rect 73125 597 73171 643
rect 73249 597 73295 643
rect 73373 597 73419 643
rect 73497 597 73543 643
rect 73621 597 73667 643
rect 73745 597 73791 643
rect 73869 597 73915 643
rect 73993 597 74039 643
rect 74117 597 74163 643
rect 74241 597 74287 643
rect 74365 597 74411 643
rect 74489 597 74535 643
rect 74613 597 74659 643
rect 74737 597 74783 643
rect 74861 597 74907 643
rect 74985 597 75031 643
rect 75109 597 75155 643
rect 75233 597 75279 643
rect 75357 597 75403 643
rect 75481 597 75527 643
rect 75605 597 75651 643
rect 75729 597 75775 643
rect 75853 597 75899 643
rect 75977 597 76023 643
rect 76101 597 76147 643
rect 76225 597 76271 643
rect 76349 597 76395 643
rect 76473 597 76519 643
rect 76597 597 76643 643
rect 76721 597 76767 643
rect 76845 597 76891 643
rect 76969 597 77015 643
rect 77093 597 77139 643
rect 77217 597 77263 643
rect 77341 597 77387 643
rect 77465 597 77511 643
rect 77589 597 77635 643
rect 77713 597 77759 643
rect 77837 597 77883 643
rect 77961 597 78007 643
rect 78085 597 78131 643
rect 78209 597 78255 643
rect 78333 597 78379 643
rect 78457 597 78503 643
rect 78581 597 78627 643
rect 78705 597 78751 643
rect 78829 597 78875 643
rect 78953 597 78999 643
rect 79077 597 79123 643
rect 79201 597 79247 643
rect 79325 597 79371 643
rect 79449 597 79495 643
rect 79573 597 79619 643
rect 79697 597 79743 643
rect 79821 597 79867 643
rect 79945 597 79991 643
rect 80069 597 80115 643
rect 80193 597 80239 643
rect 80317 597 80363 643
rect 80441 597 80487 643
rect 80565 597 80611 643
rect 80689 597 80735 643
rect 80813 597 80859 643
rect 80937 597 80983 643
rect 81061 597 81107 643
rect 81185 597 81231 643
rect 81309 597 81355 643
rect 81433 597 81479 643
rect 81557 597 81603 643
rect 81681 597 81727 643
rect 81805 597 81851 643
rect 81929 597 81975 643
rect 82053 597 82099 643
rect 82177 597 82223 643
rect 82301 597 82347 643
rect 82425 597 82471 643
rect 82549 597 82595 643
rect 82673 597 82719 643
rect 82797 597 82843 643
rect 82921 597 82967 643
rect 83045 597 83091 643
rect 83169 597 83215 643
rect 83293 597 83339 643
rect 83417 597 83463 643
rect 83541 597 83587 643
rect 83665 597 83711 643
rect 83789 597 83835 643
rect 83913 597 83959 643
rect 84037 597 84083 643
rect 84161 597 84207 643
rect 84285 597 84331 643
rect 84409 597 84455 643
rect 84533 597 84579 643
rect 84657 597 84703 643
rect 84781 597 84827 643
rect 84905 597 84951 643
rect 85029 597 85075 643
rect 85153 597 85199 643
rect 85277 597 85323 643
rect 85401 597 85447 643
rect 85525 597 85571 643
rect 85649 597 85695 643
<< metal1 >>
rect 0 46094 1000 46294
rect 0 46083 85706 46094
rect 0 46037 89 46083
rect 135 46037 213 46083
rect 259 46037 337 46083
rect 383 46037 461 46083
rect 507 46037 585 46083
rect 631 46037 709 46083
rect 755 46037 833 46083
rect 879 46037 957 46083
rect 1003 46037 1081 46083
rect 1127 46037 1205 46083
rect 1251 46037 1329 46083
rect 1375 46037 1453 46083
rect 1499 46037 1577 46083
rect 1623 46037 1701 46083
rect 1747 46037 1825 46083
rect 1871 46037 1949 46083
rect 1995 46037 2073 46083
rect 2119 46037 2197 46083
rect 2243 46037 2321 46083
rect 2367 46037 2445 46083
rect 2491 46037 2569 46083
rect 2615 46037 2693 46083
rect 2739 46037 2817 46083
rect 2863 46037 2941 46083
rect 2987 46037 3065 46083
rect 3111 46037 3189 46083
rect 3235 46037 3313 46083
rect 3359 46037 3437 46083
rect 3483 46037 3561 46083
rect 3607 46037 3685 46083
rect 3731 46037 3809 46083
rect 3855 46037 3933 46083
rect 3979 46037 4057 46083
rect 4103 46037 4181 46083
rect 4227 46037 4305 46083
rect 4351 46037 4429 46083
rect 4475 46037 4553 46083
rect 4599 46037 4677 46083
rect 4723 46037 4801 46083
rect 4847 46037 4925 46083
rect 4971 46037 5049 46083
rect 5095 46037 5173 46083
rect 5219 46037 5297 46083
rect 5343 46037 5421 46083
rect 5467 46037 5545 46083
rect 5591 46037 5669 46083
rect 5715 46037 5793 46083
rect 5839 46037 5917 46083
rect 5963 46037 6041 46083
rect 6087 46037 6165 46083
rect 6211 46037 6289 46083
rect 6335 46037 6413 46083
rect 6459 46037 6537 46083
rect 6583 46037 6661 46083
rect 6707 46037 6785 46083
rect 6831 46037 6909 46083
rect 6955 46037 7033 46083
rect 7079 46037 7157 46083
rect 7203 46037 7281 46083
rect 7327 46037 7405 46083
rect 7451 46037 7529 46083
rect 7575 46037 7653 46083
rect 7699 46037 7777 46083
rect 7823 46037 7901 46083
rect 7947 46037 8025 46083
rect 8071 46037 8149 46083
rect 8195 46037 8273 46083
rect 8319 46037 8397 46083
rect 8443 46037 8521 46083
rect 8567 46037 8645 46083
rect 8691 46037 8769 46083
rect 8815 46037 8893 46083
rect 8939 46037 9017 46083
rect 9063 46037 9141 46083
rect 9187 46037 9265 46083
rect 9311 46037 9389 46083
rect 9435 46037 9513 46083
rect 9559 46037 9637 46083
rect 9683 46037 9761 46083
rect 9807 46037 9885 46083
rect 9931 46037 10009 46083
rect 10055 46037 10133 46083
rect 10179 46037 10257 46083
rect 10303 46037 10381 46083
rect 10427 46037 10505 46083
rect 10551 46037 10629 46083
rect 10675 46037 10753 46083
rect 10799 46037 10877 46083
rect 10923 46037 11001 46083
rect 11047 46037 11125 46083
rect 11171 46037 11249 46083
rect 11295 46037 11373 46083
rect 11419 46037 11497 46083
rect 11543 46037 11621 46083
rect 11667 46037 11745 46083
rect 11791 46037 11869 46083
rect 11915 46037 11993 46083
rect 12039 46037 12117 46083
rect 12163 46037 12241 46083
rect 12287 46037 12365 46083
rect 12411 46037 12489 46083
rect 12535 46037 12613 46083
rect 12659 46037 12737 46083
rect 12783 46037 12861 46083
rect 12907 46037 12985 46083
rect 13031 46037 13109 46083
rect 13155 46037 13233 46083
rect 13279 46037 13357 46083
rect 13403 46037 13481 46083
rect 13527 46037 13605 46083
rect 13651 46037 13729 46083
rect 13775 46037 13853 46083
rect 13899 46037 13977 46083
rect 14023 46037 14101 46083
rect 14147 46037 14225 46083
rect 14271 46037 14349 46083
rect 14395 46037 14473 46083
rect 14519 46037 14597 46083
rect 14643 46037 14721 46083
rect 14767 46037 14845 46083
rect 14891 46037 14969 46083
rect 15015 46037 15093 46083
rect 15139 46037 15217 46083
rect 15263 46037 15341 46083
rect 15387 46037 15465 46083
rect 15511 46037 15589 46083
rect 15635 46037 15713 46083
rect 15759 46037 15837 46083
rect 15883 46037 15961 46083
rect 16007 46037 16085 46083
rect 16131 46037 16209 46083
rect 16255 46037 16333 46083
rect 16379 46037 16457 46083
rect 16503 46037 16581 46083
rect 16627 46037 16705 46083
rect 16751 46037 16829 46083
rect 16875 46037 16953 46083
rect 16999 46037 17077 46083
rect 17123 46037 17201 46083
rect 17247 46037 17325 46083
rect 17371 46037 17449 46083
rect 17495 46037 17573 46083
rect 17619 46037 17697 46083
rect 17743 46037 17821 46083
rect 17867 46037 17945 46083
rect 17991 46037 18069 46083
rect 18115 46037 18193 46083
rect 18239 46037 18317 46083
rect 18363 46037 18441 46083
rect 18487 46037 18565 46083
rect 18611 46037 18689 46083
rect 18735 46037 18813 46083
rect 18859 46037 18937 46083
rect 18983 46037 19061 46083
rect 19107 46037 19185 46083
rect 19231 46037 19309 46083
rect 19355 46037 19433 46083
rect 19479 46037 19557 46083
rect 19603 46037 19681 46083
rect 19727 46037 19805 46083
rect 19851 46037 19929 46083
rect 19975 46037 20053 46083
rect 20099 46037 20177 46083
rect 20223 46037 20301 46083
rect 20347 46037 20425 46083
rect 20471 46037 20549 46083
rect 20595 46037 20673 46083
rect 20719 46037 20797 46083
rect 20843 46037 20921 46083
rect 20967 46037 21045 46083
rect 21091 46037 21169 46083
rect 21215 46037 21293 46083
rect 21339 46037 21417 46083
rect 21463 46037 21541 46083
rect 21587 46037 21665 46083
rect 21711 46037 21789 46083
rect 21835 46037 21913 46083
rect 21959 46037 22037 46083
rect 22083 46037 22161 46083
rect 22207 46037 22285 46083
rect 22331 46037 22409 46083
rect 22455 46037 22533 46083
rect 22579 46037 22657 46083
rect 22703 46037 22781 46083
rect 22827 46037 22905 46083
rect 22951 46037 23029 46083
rect 23075 46037 23153 46083
rect 23199 46037 23277 46083
rect 23323 46037 23401 46083
rect 23447 46037 23525 46083
rect 23571 46037 23649 46083
rect 23695 46037 23773 46083
rect 23819 46037 23897 46083
rect 23943 46037 24021 46083
rect 24067 46037 24145 46083
rect 24191 46037 24269 46083
rect 24315 46037 24393 46083
rect 24439 46037 24517 46083
rect 24563 46037 24641 46083
rect 24687 46037 24765 46083
rect 24811 46037 24889 46083
rect 24935 46037 25013 46083
rect 25059 46037 25137 46083
rect 25183 46037 25261 46083
rect 25307 46037 25385 46083
rect 25431 46037 25509 46083
rect 25555 46037 25633 46083
rect 25679 46037 25757 46083
rect 25803 46037 25881 46083
rect 25927 46037 26005 46083
rect 26051 46037 26129 46083
rect 26175 46037 26253 46083
rect 26299 46037 26377 46083
rect 26423 46037 26501 46083
rect 26547 46037 26625 46083
rect 26671 46037 26749 46083
rect 26795 46037 26873 46083
rect 26919 46037 26997 46083
rect 27043 46037 27121 46083
rect 27167 46037 27245 46083
rect 27291 46037 27369 46083
rect 27415 46037 27493 46083
rect 27539 46037 27617 46083
rect 27663 46037 27741 46083
rect 27787 46037 27865 46083
rect 27911 46037 27989 46083
rect 28035 46037 28113 46083
rect 28159 46037 28237 46083
rect 28283 46037 28361 46083
rect 28407 46037 28485 46083
rect 28531 46037 28609 46083
rect 28655 46037 28733 46083
rect 28779 46037 28857 46083
rect 28903 46037 28981 46083
rect 29027 46037 29105 46083
rect 29151 46037 29229 46083
rect 29275 46037 29353 46083
rect 29399 46037 29477 46083
rect 29523 46037 29601 46083
rect 29647 46037 29725 46083
rect 29771 46037 29849 46083
rect 29895 46037 29973 46083
rect 30019 46037 30097 46083
rect 30143 46037 30221 46083
rect 30267 46037 30345 46083
rect 30391 46037 30469 46083
rect 30515 46037 30593 46083
rect 30639 46037 30717 46083
rect 30763 46037 30841 46083
rect 30887 46037 30965 46083
rect 31011 46037 31089 46083
rect 31135 46037 31213 46083
rect 31259 46037 31337 46083
rect 31383 46037 31461 46083
rect 31507 46037 31585 46083
rect 31631 46037 31709 46083
rect 31755 46037 31833 46083
rect 31879 46037 31957 46083
rect 32003 46037 32081 46083
rect 32127 46037 32205 46083
rect 32251 46037 32329 46083
rect 32375 46037 32453 46083
rect 32499 46037 32577 46083
rect 32623 46037 32701 46083
rect 32747 46037 32825 46083
rect 32871 46037 32949 46083
rect 32995 46037 33073 46083
rect 33119 46037 33197 46083
rect 33243 46037 33321 46083
rect 33367 46037 33445 46083
rect 33491 46037 33569 46083
rect 33615 46037 33693 46083
rect 33739 46037 33817 46083
rect 33863 46037 33941 46083
rect 33987 46037 34065 46083
rect 34111 46037 34189 46083
rect 34235 46037 34313 46083
rect 34359 46037 34437 46083
rect 34483 46037 34561 46083
rect 34607 46037 34685 46083
rect 34731 46037 34809 46083
rect 34855 46037 34933 46083
rect 34979 46037 35057 46083
rect 35103 46037 35181 46083
rect 35227 46037 35305 46083
rect 35351 46037 35429 46083
rect 35475 46037 35553 46083
rect 35599 46037 35677 46083
rect 35723 46037 35801 46083
rect 35847 46037 35925 46083
rect 35971 46037 36049 46083
rect 36095 46037 36173 46083
rect 36219 46037 36297 46083
rect 36343 46037 36421 46083
rect 36467 46037 36545 46083
rect 36591 46037 36669 46083
rect 36715 46037 36793 46083
rect 36839 46037 36917 46083
rect 36963 46037 37041 46083
rect 37087 46037 37165 46083
rect 37211 46037 37289 46083
rect 37335 46037 37413 46083
rect 37459 46037 37537 46083
rect 37583 46037 37661 46083
rect 37707 46037 37785 46083
rect 37831 46037 37909 46083
rect 37955 46037 38033 46083
rect 38079 46037 38157 46083
rect 38203 46037 38281 46083
rect 38327 46037 38405 46083
rect 38451 46037 38529 46083
rect 38575 46037 38653 46083
rect 38699 46037 38777 46083
rect 38823 46037 38901 46083
rect 38947 46037 39025 46083
rect 39071 46037 39149 46083
rect 39195 46037 39273 46083
rect 39319 46037 39397 46083
rect 39443 46037 39521 46083
rect 39567 46037 39645 46083
rect 39691 46037 39769 46083
rect 39815 46037 39893 46083
rect 39939 46037 40017 46083
rect 40063 46037 40141 46083
rect 40187 46037 40265 46083
rect 40311 46037 40389 46083
rect 40435 46037 40513 46083
rect 40559 46037 40637 46083
rect 40683 46037 40761 46083
rect 40807 46037 40885 46083
rect 40931 46037 41009 46083
rect 41055 46037 41133 46083
rect 41179 46037 41257 46083
rect 41303 46037 41381 46083
rect 41427 46037 41505 46083
rect 41551 46037 41629 46083
rect 41675 46037 41753 46083
rect 41799 46037 41877 46083
rect 41923 46037 42001 46083
rect 42047 46037 42125 46083
rect 42171 46037 42249 46083
rect 42295 46037 42373 46083
rect 42419 46037 42497 46083
rect 42543 46037 42621 46083
rect 42667 46037 42745 46083
rect 42791 46037 42869 46083
rect 42915 46037 42993 46083
rect 43039 46037 43117 46083
rect 43163 46037 43241 46083
rect 43287 46037 43365 46083
rect 43411 46037 43489 46083
rect 43535 46037 43613 46083
rect 43659 46037 43737 46083
rect 43783 46037 43861 46083
rect 43907 46037 43985 46083
rect 44031 46037 44109 46083
rect 44155 46037 44233 46083
rect 44279 46037 44357 46083
rect 44403 46037 44481 46083
rect 44527 46037 44605 46083
rect 44651 46037 44729 46083
rect 44775 46037 44853 46083
rect 44899 46037 44977 46083
rect 45023 46037 45101 46083
rect 45147 46037 45225 46083
rect 45271 46037 45349 46083
rect 45395 46037 45473 46083
rect 45519 46037 45597 46083
rect 45643 46037 45721 46083
rect 45767 46037 45845 46083
rect 45891 46037 45969 46083
rect 46015 46037 46093 46083
rect 46139 46037 46217 46083
rect 46263 46037 46341 46083
rect 46387 46037 46465 46083
rect 46511 46037 46589 46083
rect 46635 46037 46713 46083
rect 46759 46037 46837 46083
rect 46883 46037 46961 46083
rect 47007 46037 47085 46083
rect 47131 46037 47209 46083
rect 47255 46037 47333 46083
rect 47379 46037 47457 46083
rect 47503 46037 47581 46083
rect 47627 46037 47705 46083
rect 47751 46037 47829 46083
rect 47875 46037 47953 46083
rect 47999 46037 48077 46083
rect 48123 46037 48201 46083
rect 48247 46037 48325 46083
rect 48371 46037 48449 46083
rect 48495 46037 48573 46083
rect 48619 46037 48697 46083
rect 48743 46037 48821 46083
rect 48867 46037 48945 46083
rect 48991 46037 49069 46083
rect 49115 46037 49193 46083
rect 49239 46037 49317 46083
rect 49363 46037 49441 46083
rect 49487 46037 49565 46083
rect 49611 46037 49689 46083
rect 49735 46037 49813 46083
rect 49859 46037 49937 46083
rect 49983 46037 50061 46083
rect 50107 46037 50185 46083
rect 50231 46037 50309 46083
rect 50355 46037 50433 46083
rect 50479 46037 50557 46083
rect 50603 46037 50681 46083
rect 50727 46037 50805 46083
rect 50851 46037 50929 46083
rect 50975 46037 51053 46083
rect 51099 46037 51177 46083
rect 51223 46037 51301 46083
rect 51347 46037 51425 46083
rect 51471 46037 51549 46083
rect 51595 46037 51673 46083
rect 51719 46037 51797 46083
rect 51843 46037 51921 46083
rect 51967 46037 52045 46083
rect 52091 46037 52169 46083
rect 52215 46037 52293 46083
rect 52339 46037 52417 46083
rect 52463 46037 52541 46083
rect 52587 46037 52665 46083
rect 52711 46037 52789 46083
rect 52835 46037 52913 46083
rect 52959 46037 53037 46083
rect 53083 46037 53161 46083
rect 53207 46037 53285 46083
rect 53331 46037 53409 46083
rect 53455 46037 53533 46083
rect 53579 46037 53657 46083
rect 53703 46037 53781 46083
rect 53827 46037 53905 46083
rect 53951 46037 54029 46083
rect 54075 46037 54153 46083
rect 54199 46037 54277 46083
rect 54323 46037 54401 46083
rect 54447 46037 54525 46083
rect 54571 46037 54649 46083
rect 54695 46037 54773 46083
rect 54819 46037 54897 46083
rect 54943 46037 55021 46083
rect 55067 46037 55145 46083
rect 55191 46037 55269 46083
rect 55315 46037 55393 46083
rect 55439 46037 55517 46083
rect 55563 46037 55641 46083
rect 55687 46037 55765 46083
rect 55811 46037 55889 46083
rect 55935 46037 56013 46083
rect 56059 46037 56137 46083
rect 56183 46037 56261 46083
rect 56307 46037 56385 46083
rect 56431 46037 56509 46083
rect 56555 46037 56633 46083
rect 56679 46037 56757 46083
rect 56803 46037 56881 46083
rect 56927 46037 57005 46083
rect 57051 46037 57129 46083
rect 57175 46037 57253 46083
rect 57299 46037 57377 46083
rect 57423 46037 57501 46083
rect 57547 46037 57625 46083
rect 57671 46037 57749 46083
rect 57795 46037 57873 46083
rect 57919 46037 57997 46083
rect 58043 46037 58121 46083
rect 58167 46037 58245 46083
rect 58291 46037 58369 46083
rect 58415 46037 58493 46083
rect 58539 46037 58617 46083
rect 58663 46037 58741 46083
rect 58787 46037 58865 46083
rect 58911 46037 58989 46083
rect 59035 46037 59113 46083
rect 59159 46037 59237 46083
rect 59283 46037 59361 46083
rect 59407 46037 59485 46083
rect 59531 46037 59609 46083
rect 59655 46037 59733 46083
rect 59779 46037 59857 46083
rect 59903 46037 59981 46083
rect 60027 46037 60105 46083
rect 60151 46037 60229 46083
rect 60275 46037 60353 46083
rect 60399 46037 60477 46083
rect 60523 46037 60601 46083
rect 60647 46037 60725 46083
rect 60771 46037 60849 46083
rect 60895 46037 60973 46083
rect 61019 46037 61097 46083
rect 61143 46037 61221 46083
rect 61267 46037 61345 46083
rect 61391 46037 61469 46083
rect 61515 46037 61593 46083
rect 61639 46037 61717 46083
rect 61763 46037 61841 46083
rect 61887 46037 61965 46083
rect 62011 46037 62089 46083
rect 62135 46037 62213 46083
rect 62259 46037 62337 46083
rect 62383 46037 62461 46083
rect 62507 46037 62585 46083
rect 62631 46037 62709 46083
rect 62755 46037 62833 46083
rect 62879 46037 62957 46083
rect 63003 46037 63081 46083
rect 63127 46037 63205 46083
rect 63251 46037 63329 46083
rect 63375 46037 63453 46083
rect 63499 46037 63577 46083
rect 63623 46037 63701 46083
rect 63747 46037 63825 46083
rect 63871 46037 63949 46083
rect 63995 46037 64073 46083
rect 64119 46037 64197 46083
rect 64243 46037 64321 46083
rect 64367 46037 64445 46083
rect 64491 46037 64569 46083
rect 64615 46037 64693 46083
rect 64739 46037 64817 46083
rect 64863 46037 64941 46083
rect 64987 46037 65065 46083
rect 65111 46037 65189 46083
rect 65235 46037 65313 46083
rect 65359 46037 65437 46083
rect 65483 46037 65561 46083
rect 65607 46037 65685 46083
rect 65731 46037 65809 46083
rect 65855 46037 65933 46083
rect 65979 46037 66057 46083
rect 66103 46037 66181 46083
rect 66227 46037 66305 46083
rect 66351 46037 66429 46083
rect 66475 46037 66553 46083
rect 66599 46037 66677 46083
rect 66723 46037 66801 46083
rect 66847 46037 66925 46083
rect 66971 46037 67049 46083
rect 67095 46037 67173 46083
rect 67219 46037 67297 46083
rect 67343 46037 67421 46083
rect 67467 46037 67545 46083
rect 67591 46037 67669 46083
rect 67715 46037 67793 46083
rect 67839 46037 67917 46083
rect 67963 46037 68041 46083
rect 68087 46037 68165 46083
rect 68211 46037 68289 46083
rect 68335 46037 68413 46083
rect 68459 46037 68537 46083
rect 68583 46037 68661 46083
rect 68707 46037 68785 46083
rect 68831 46037 68909 46083
rect 68955 46037 69033 46083
rect 69079 46037 69157 46083
rect 69203 46037 69281 46083
rect 69327 46037 69405 46083
rect 69451 46037 69529 46083
rect 69575 46037 69653 46083
rect 69699 46037 69777 46083
rect 69823 46037 69901 46083
rect 69947 46037 70025 46083
rect 70071 46037 70149 46083
rect 70195 46037 70273 46083
rect 70319 46037 70397 46083
rect 70443 46037 70521 46083
rect 70567 46037 70645 46083
rect 70691 46037 70769 46083
rect 70815 46037 70893 46083
rect 70939 46037 71017 46083
rect 71063 46037 71141 46083
rect 71187 46037 71265 46083
rect 71311 46037 71389 46083
rect 71435 46037 71513 46083
rect 71559 46037 71637 46083
rect 71683 46037 71761 46083
rect 71807 46037 71885 46083
rect 71931 46037 72009 46083
rect 72055 46037 72133 46083
rect 72179 46037 72257 46083
rect 72303 46037 72381 46083
rect 72427 46037 72505 46083
rect 72551 46037 72629 46083
rect 72675 46037 72753 46083
rect 72799 46037 72877 46083
rect 72923 46037 73001 46083
rect 73047 46037 73125 46083
rect 73171 46037 73249 46083
rect 73295 46037 73373 46083
rect 73419 46037 73497 46083
rect 73543 46037 73621 46083
rect 73667 46037 73745 46083
rect 73791 46037 73869 46083
rect 73915 46037 73993 46083
rect 74039 46037 74117 46083
rect 74163 46037 74241 46083
rect 74287 46037 74365 46083
rect 74411 46037 74489 46083
rect 74535 46037 74613 46083
rect 74659 46037 74737 46083
rect 74783 46037 74861 46083
rect 74907 46037 74985 46083
rect 75031 46037 75109 46083
rect 75155 46037 75233 46083
rect 75279 46037 75357 46083
rect 75403 46037 75481 46083
rect 75527 46037 75605 46083
rect 75651 46037 75729 46083
rect 75775 46037 75853 46083
rect 75899 46037 75977 46083
rect 76023 46037 76101 46083
rect 76147 46037 76225 46083
rect 76271 46037 76349 46083
rect 76395 46037 76473 46083
rect 76519 46037 76597 46083
rect 76643 46037 76721 46083
rect 76767 46037 76845 46083
rect 76891 46037 76969 46083
rect 77015 46037 77093 46083
rect 77139 46037 77217 46083
rect 77263 46037 77341 46083
rect 77387 46037 77465 46083
rect 77511 46037 77589 46083
rect 77635 46037 77713 46083
rect 77759 46037 77837 46083
rect 77883 46037 77961 46083
rect 78007 46037 78085 46083
rect 78131 46037 78209 46083
rect 78255 46037 78333 46083
rect 78379 46037 78457 46083
rect 78503 46037 78581 46083
rect 78627 46037 78705 46083
rect 78751 46037 78829 46083
rect 78875 46037 78953 46083
rect 78999 46037 79077 46083
rect 79123 46037 79201 46083
rect 79247 46037 79325 46083
rect 79371 46037 79449 46083
rect 79495 46037 79573 46083
rect 79619 46037 79697 46083
rect 79743 46037 79821 46083
rect 79867 46037 79945 46083
rect 79991 46037 80069 46083
rect 80115 46037 80193 46083
rect 80239 46037 80317 46083
rect 80363 46037 80441 46083
rect 80487 46037 80565 46083
rect 80611 46037 80689 46083
rect 80735 46037 80813 46083
rect 80859 46037 80937 46083
rect 80983 46037 81061 46083
rect 81107 46037 81185 46083
rect 81231 46037 81309 46083
rect 81355 46037 81433 46083
rect 81479 46037 81557 46083
rect 81603 46037 81681 46083
rect 81727 46037 81805 46083
rect 81851 46037 81929 46083
rect 81975 46037 82053 46083
rect 82099 46037 82177 46083
rect 82223 46037 82301 46083
rect 82347 46037 82425 46083
rect 82471 46037 82549 46083
rect 82595 46037 82673 46083
rect 82719 46037 82797 46083
rect 82843 46037 82921 46083
rect 82967 46037 83045 46083
rect 83091 46037 83169 46083
rect 83215 46037 83293 46083
rect 83339 46037 83417 46083
rect 83463 46037 83541 46083
rect 83587 46037 83665 46083
rect 83711 46037 83789 46083
rect 83835 46037 83913 46083
rect 83959 46037 84037 46083
rect 84083 46037 84161 46083
rect 84207 46037 84285 46083
rect 84331 46037 84409 46083
rect 84455 46037 84533 46083
rect 84579 46037 84657 46083
rect 84703 46037 84781 46083
rect 84827 46037 84905 46083
rect 84951 46037 85029 46083
rect 85075 46037 85153 46083
rect 85199 46037 85277 46083
rect 85323 46037 85401 46083
rect 85447 46037 85525 46083
rect 85571 46037 85649 46083
rect 85695 46037 85706 46083
rect 0 45959 85706 46037
rect 0 45913 89 45959
rect 135 45913 213 45959
rect 259 45913 337 45959
rect 383 45913 461 45959
rect 507 45913 585 45959
rect 631 45913 709 45959
rect 755 45913 833 45959
rect 879 45913 957 45959
rect 1003 45913 1081 45959
rect 1127 45913 1205 45959
rect 1251 45913 1329 45959
rect 1375 45913 1453 45959
rect 1499 45913 1577 45959
rect 1623 45913 1701 45959
rect 1747 45913 1825 45959
rect 1871 45913 1949 45959
rect 1995 45913 2073 45959
rect 2119 45913 2197 45959
rect 2243 45913 2321 45959
rect 2367 45913 2445 45959
rect 2491 45913 2569 45959
rect 2615 45913 2693 45959
rect 2739 45913 2817 45959
rect 2863 45913 2941 45959
rect 2987 45913 3065 45959
rect 3111 45913 3189 45959
rect 3235 45913 3313 45959
rect 3359 45913 3437 45959
rect 3483 45913 3561 45959
rect 3607 45913 3685 45959
rect 3731 45913 3809 45959
rect 3855 45913 3933 45959
rect 3979 45913 4057 45959
rect 4103 45913 4181 45959
rect 4227 45913 4305 45959
rect 4351 45913 4429 45959
rect 4475 45913 4553 45959
rect 4599 45913 4677 45959
rect 4723 45913 4801 45959
rect 4847 45913 4925 45959
rect 4971 45913 5049 45959
rect 5095 45913 5173 45959
rect 5219 45913 5297 45959
rect 5343 45913 5421 45959
rect 5467 45913 5545 45959
rect 5591 45913 5669 45959
rect 5715 45913 5793 45959
rect 5839 45913 5917 45959
rect 5963 45913 6041 45959
rect 6087 45913 6165 45959
rect 6211 45913 6289 45959
rect 6335 45913 6413 45959
rect 6459 45913 6537 45959
rect 6583 45913 6661 45959
rect 6707 45913 6785 45959
rect 6831 45913 6909 45959
rect 6955 45913 7033 45959
rect 7079 45913 7157 45959
rect 7203 45913 7281 45959
rect 7327 45913 7405 45959
rect 7451 45913 7529 45959
rect 7575 45913 7653 45959
rect 7699 45913 7777 45959
rect 7823 45913 7901 45959
rect 7947 45913 8025 45959
rect 8071 45913 8149 45959
rect 8195 45913 8273 45959
rect 8319 45913 8397 45959
rect 8443 45913 8521 45959
rect 8567 45913 8645 45959
rect 8691 45913 8769 45959
rect 8815 45913 8893 45959
rect 8939 45913 9017 45959
rect 9063 45913 9141 45959
rect 9187 45913 9265 45959
rect 9311 45913 9389 45959
rect 9435 45913 9513 45959
rect 9559 45913 9637 45959
rect 9683 45913 9761 45959
rect 9807 45913 9885 45959
rect 9931 45913 10009 45959
rect 10055 45913 10133 45959
rect 10179 45913 10257 45959
rect 10303 45913 10381 45959
rect 10427 45913 10505 45959
rect 10551 45913 10629 45959
rect 10675 45913 10753 45959
rect 10799 45913 10877 45959
rect 10923 45913 11001 45959
rect 11047 45913 11125 45959
rect 11171 45913 11249 45959
rect 11295 45913 11373 45959
rect 11419 45913 11497 45959
rect 11543 45913 11621 45959
rect 11667 45913 11745 45959
rect 11791 45913 11869 45959
rect 11915 45913 11993 45959
rect 12039 45913 12117 45959
rect 12163 45913 12241 45959
rect 12287 45913 12365 45959
rect 12411 45913 12489 45959
rect 12535 45913 12613 45959
rect 12659 45913 12737 45959
rect 12783 45913 12861 45959
rect 12907 45913 12985 45959
rect 13031 45913 13109 45959
rect 13155 45913 13233 45959
rect 13279 45913 13357 45959
rect 13403 45913 13481 45959
rect 13527 45913 13605 45959
rect 13651 45913 13729 45959
rect 13775 45913 13853 45959
rect 13899 45913 13977 45959
rect 14023 45913 14101 45959
rect 14147 45913 14225 45959
rect 14271 45913 14349 45959
rect 14395 45913 14473 45959
rect 14519 45913 14597 45959
rect 14643 45913 14721 45959
rect 14767 45913 14845 45959
rect 14891 45913 14969 45959
rect 15015 45913 15093 45959
rect 15139 45913 15217 45959
rect 15263 45913 15341 45959
rect 15387 45913 15465 45959
rect 15511 45913 15589 45959
rect 15635 45913 15713 45959
rect 15759 45913 15837 45959
rect 15883 45913 15961 45959
rect 16007 45913 16085 45959
rect 16131 45913 16209 45959
rect 16255 45913 16333 45959
rect 16379 45913 16457 45959
rect 16503 45913 16581 45959
rect 16627 45913 16705 45959
rect 16751 45913 16829 45959
rect 16875 45913 16953 45959
rect 16999 45913 17077 45959
rect 17123 45913 17201 45959
rect 17247 45913 17325 45959
rect 17371 45913 17449 45959
rect 17495 45913 17573 45959
rect 17619 45913 17697 45959
rect 17743 45913 17821 45959
rect 17867 45913 17945 45959
rect 17991 45913 18069 45959
rect 18115 45913 18193 45959
rect 18239 45913 18317 45959
rect 18363 45913 18441 45959
rect 18487 45913 18565 45959
rect 18611 45913 18689 45959
rect 18735 45913 18813 45959
rect 18859 45913 18937 45959
rect 18983 45913 19061 45959
rect 19107 45913 19185 45959
rect 19231 45913 19309 45959
rect 19355 45913 19433 45959
rect 19479 45913 19557 45959
rect 19603 45913 19681 45959
rect 19727 45913 19805 45959
rect 19851 45913 19929 45959
rect 19975 45913 20053 45959
rect 20099 45913 20177 45959
rect 20223 45913 20301 45959
rect 20347 45913 20425 45959
rect 20471 45913 20549 45959
rect 20595 45913 20673 45959
rect 20719 45913 20797 45959
rect 20843 45913 20921 45959
rect 20967 45913 21045 45959
rect 21091 45913 21169 45959
rect 21215 45913 21293 45959
rect 21339 45913 21417 45959
rect 21463 45913 21541 45959
rect 21587 45913 21665 45959
rect 21711 45913 21789 45959
rect 21835 45913 21913 45959
rect 21959 45913 22037 45959
rect 22083 45913 22161 45959
rect 22207 45913 22285 45959
rect 22331 45913 22409 45959
rect 22455 45913 22533 45959
rect 22579 45913 22657 45959
rect 22703 45913 22781 45959
rect 22827 45913 22905 45959
rect 22951 45913 23029 45959
rect 23075 45913 23153 45959
rect 23199 45913 23277 45959
rect 23323 45913 23401 45959
rect 23447 45913 23525 45959
rect 23571 45913 23649 45959
rect 23695 45913 23773 45959
rect 23819 45913 23897 45959
rect 23943 45913 24021 45959
rect 24067 45913 24145 45959
rect 24191 45913 24269 45959
rect 24315 45913 24393 45959
rect 24439 45913 24517 45959
rect 24563 45913 24641 45959
rect 24687 45913 24765 45959
rect 24811 45913 24889 45959
rect 24935 45913 25013 45959
rect 25059 45913 25137 45959
rect 25183 45913 25261 45959
rect 25307 45913 25385 45959
rect 25431 45913 25509 45959
rect 25555 45913 25633 45959
rect 25679 45913 25757 45959
rect 25803 45913 25881 45959
rect 25927 45913 26005 45959
rect 26051 45913 26129 45959
rect 26175 45913 26253 45959
rect 26299 45913 26377 45959
rect 26423 45913 26501 45959
rect 26547 45913 26625 45959
rect 26671 45913 26749 45959
rect 26795 45913 26873 45959
rect 26919 45913 26997 45959
rect 27043 45913 27121 45959
rect 27167 45913 27245 45959
rect 27291 45913 27369 45959
rect 27415 45913 27493 45959
rect 27539 45913 27617 45959
rect 27663 45913 27741 45959
rect 27787 45913 27865 45959
rect 27911 45913 27989 45959
rect 28035 45913 28113 45959
rect 28159 45913 28237 45959
rect 28283 45913 28361 45959
rect 28407 45913 28485 45959
rect 28531 45913 28609 45959
rect 28655 45913 28733 45959
rect 28779 45913 28857 45959
rect 28903 45913 28981 45959
rect 29027 45913 29105 45959
rect 29151 45913 29229 45959
rect 29275 45913 29353 45959
rect 29399 45913 29477 45959
rect 29523 45913 29601 45959
rect 29647 45913 29725 45959
rect 29771 45913 29849 45959
rect 29895 45913 29973 45959
rect 30019 45913 30097 45959
rect 30143 45913 30221 45959
rect 30267 45913 30345 45959
rect 30391 45913 30469 45959
rect 30515 45913 30593 45959
rect 30639 45913 30717 45959
rect 30763 45913 30841 45959
rect 30887 45913 30965 45959
rect 31011 45913 31089 45959
rect 31135 45913 31213 45959
rect 31259 45913 31337 45959
rect 31383 45913 31461 45959
rect 31507 45913 31585 45959
rect 31631 45913 31709 45959
rect 31755 45913 31833 45959
rect 31879 45913 31957 45959
rect 32003 45913 32081 45959
rect 32127 45913 32205 45959
rect 32251 45913 32329 45959
rect 32375 45913 32453 45959
rect 32499 45913 32577 45959
rect 32623 45913 32701 45959
rect 32747 45913 32825 45959
rect 32871 45913 32949 45959
rect 32995 45913 33073 45959
rect 33119 45913 33197 45959
rect 33243 45913 33321 45959
rect 33367 45913 33445 45959
rect 33491 45913 33569 45959
rect 33615 45913 33693 45959
rect 33739 45913 33817 45959
rect 33863 45913 33941 45959
rect 33987 45913 34065 45959
rect 34111 45913 34189 45959
rect 34235 45913 34313 45959
rect 34359 45913 34437 45959
rect 34483 45913 34561 45959
rect 34607 45913 34685 45959
rect 34731 45913 34809 45959
rect 34855 45913 34933 45959
rect 34979 45913 35057 45959
rect 35103 45913 35181 45959
rect 35227 45913 35305 45959
rect 35351 45913 35429 45959
rect 35475 45913 35553 45959
rect 35599 45913 35677 45959
rect 35723 45913 35801 45959
rect 35847 45913 35925 45959
rect 35971 45913 36049 45959
rect 36095 45913 36173 45959
rect 36219 45913 36297 45959
rect 36343 45913 36421 45959
rect 36467 45913 36545 45959
rect 36591 45913 36669 45959
rect 36715 45913 36793 45959
rect 36839 45913 36917 45959
rect 36963 45913 37041 45959
rect 37087 45913 37165 45959
rect 37211 45913 37289 45959
rect 37335 45913 37413 45959
rect 37459 45913 37537 45959
rect 37583 45913 37661 45959
rect 37707 45913 37785 45959
rect 37831 45913 37909 45959
rect 37955 45913 38033 45959
rect 38079 45913 38157 45959
rect 38203 45913 38281 45959
rect 38327 45913 38405 45959
rect 38451 45913 38529 45959
rect 38575 45913 38653 45959
rect 38699 45913 38777 45959
rect 38823 45913 38901 45959
rect 38947 45913 39025 45959
rect 39071 45913 39149 45959
rect 39195 45913 39273 45959
rect 39319 45913 39397 45959
rect 39443 45913 39521 45959
rect 39567 45913 39645 45959
rect 39691 45913 39769 45959
rect 39815 45913 39893 45959
rect 39939 45913 40017 45959
rect 40063 45913 40141 45959
rect 40187 45913 40265 45959
rect 40311 45913 40389 45959
rect 40435 45913 40513 45959
rect 40559 45913 40637 45959
rect 40683 45913 40761 45959
rect 40807 45913 40885 45959
rect 40931 45913 41009 45959
rect 41055 45913 41133 45959
rect 41179 45913 41257 45959
rect 41303 45913 41381 45959
rect 41427 45913 41505 45959
rect 41551 45913 41629 45959
rect 41675 45913 41753 45959
rect 41799 45913 41877 45959
rect 41923 45913 42001 45959
rect 42047 45913 42125 45959
rect 42171 45913 42249 45959
rect 42295 45913 42373 45959
rect 42419 45913 42497 45959
rect 42543 45913 42621 45959
rect 42667 45913 42745 45959
rect 42791 45913 42869 45959
rect 42915 45913 42993 45959
rect 43039 45913 43117 45959
rect 43163 45913 43241 45959
rect 43287 45913 43365 45959
rect 43411 45913 43489 45959
rect 43535 45913 43613 45959
rect 43659 45913 43737 45959
rect 43783 45913 43861 45959
rect 43907 45913 43985 45959
rect 44031 45913 44109 45959
rect 44155 45913 44233 45959
rect 44279 45913 44357 45959
rect 44403 45913 44481 45959
rect 44527 45913 44605 45959
rect 44651 45913 44729 45959
rect 44775 45913 44853 45959
rect 44899 45913 44977 45959
rect 45023 45913 45101 45959
rect 45147 45913 45225 45959
rect 45271 45913 45349 45959
rect 45395 45913 45473 45959
rect 45519 45913 45597 45959
rect 45643 45913 45721 45959
rect 45767 45913 45845 45959
rect 45891 45913 45969 45959
rect 46015 45913 46093 45959
rect 46139 45913 46217 45959
rect 46263 45913 46341 45959
rect 46387 45913 46465 45959
rect 46511 45913 46589 45959
rect 46635 45913 46713 45959
rect 46759 45913 46837 45959
rect 46883 45913 46961 45959
rect 47007 45913 47085 45959
rect 47131 45913 47209 45959
rect 47255 45913 47333 45959
rect 47379 45913 47457 45959
rect 47503 45913 47581 45959
rect 47627 45913 47705 45959
rect 47751 45913 47829 45959
rect 47875 45913 47953 45959
rect 47999 45913 48077 45959
rect 48123 45913 48201 45959
rect 48247 45913 48325 45959
rect 48371 45913 48449 45959
rect 48495 45913 48573 45959
rect 48619 45913 48697 45959
rect 48743 45913 48821 45959
rect 48867 45913 48945 45959
rect 48991 45913 49069 45959
rect 49115 45913 49193 45959
rect 49239 45913 49317 45959
rect 49363 45913 49441 45959
rect 49487 45913 49565 45959
rect 49611 45913 49689 45959
rect 49735 45913 49813 45959
rect 49859 45913 49937 45959
rect 49983 45913 50061 45959
rect 50107 45913 50185 45959
rect 50231 45913 50309 45959
rect 50355 45913 50433 45959
rect 50479 45913 50557 45959
rect 50603 45913 50681 45959
rect 50727 45913 50805 45959
rect 50851 45913 50929 45959
rect 50975 45913 51053 45959
rect 51099 45913 51177 45959
rect 51223 45913 51301 45959
rect 51347 45913 51425 45959
rect 51471 45913 51549 45959
rect 51595 45913 51673 45959
rect 51719 45913 51797 45959
rect 51843 45913 51921 45959
rect 51967 45913 52045 45959
rect 52091 45913 52169 45959
rect 52215 45913 52293 45959
rect 52339 45913 52417 45959
rect 52463 45913 52541 45959
rect 52587 45913 52665 45959
rect 52711 45913 52789 45959
rect 52835 45913 52913 45959
rect 52959 45913 53037 45959
rect 53083 45913 53161 45959
rect 53207 45913 53285 45959
rect 53331 45913 53409 45959
rect 53455 45913 53533 45959
rect 53579 45913 53657 45959
rect 53703 45913 53781 45959
rect 53827 45913 53905 45959
rect 53951 45913 54029 45959
rect 54075 45913 54153 45959
rect 54199 45913 54277 45959
rect 54323 45913 54401 45959
rect 54447 45913 54525 45959
rect 54571 45913 54649 45959
rect 54695 45913 54773 45959
rect 54819 45913 54897 45959
rect 54943 45913 55021 45959
rect 55067 45913 55145 45959
rect 55191 45913 55269 45959
rect 55315 45913 55393 45959
rect 55439 45913 55517 45959
rect 55563 45913 55641 45959
rect 55687 45913 55765 45959
rect 55811 45913 55889 45959
rect 55935 45913 56013 45959
rect 56059 45913 56137 45959
rect 56183 45913 56261 45959
rect 56307 45913 56385 45959
rect 56431 45913 56509 45959
rect 56555 45913 56633 45959
rect 56679 45913 56757 45959
rect 56803 45913 56881 45959
rect 56927 45913 57005 45959
rect 57051 45913 57129 45959
rect 57175 45913 57253 45959
rect 57299 45913 57377 45959
rect 57423 45913 57501 45959
rect 57547 45913 57625 45959
rect 57671 45913 57749 45959
rect 57795 45913 57873 45959
rect 57919 45913 57997 45959
rect 58043 45913 58121 45959
rect 58167 45913 58245 45959
rect 58291 45913 58369 45959
rect 58415 45913 58493 45959
rect 58539 45913 58617 45959
rect 58663 45913 58741 45959
rect 58787 45913 58865 45959
rect 58911 45913 58989 45959
rect 59035 45913 59113 45959
rect 59159 45913 59237 45959
rect 59283 45913 59361 45959
rect 59407 45913 59485 45959
rect 59531 45913 59609 45959
rect 59655 45913 59733 45959
rect 59779 45913 59857 45959
rect 59903 45913 59981 45959
rect 60027 45913 60105 45959
rect 60151 45913 60229 45959
rect 60275 45913 60353 45959
rect 60399 45913 60477 45959
rect 60523 45913 60601 45959
rect 60647 45913 60725 45959
rect 60771 45913 60849 45959
rect 60895 45913 60973 45959
rect 61019 45913 61097 45959
rect 61143 45913 61221 45959
rect 61267 45913 61345 45959
rect 61391 45913 61469 45959
rect 61515 45913 61593 45959
rect 61639 45913 61717 45959
rect 61763 45913 61841 45959
rect 61887 45913 61965 45959
rect 62011 45913 62089 45959
rect 62135 45913 62213 45959
rect 62259 45913 62337 45959
rect 62383 45913 62461 45959
rect 62507 45913 62585 45959
rect 62631 45913 62709 45959
rect 62755 45913 62833 45959
rect 62879 45913 62957 45959
rect 63003 45913 63081 45959
rect 63127 45913 63205 45959
rect 63251 45913 63329 45959
rect 63375 45913 63453 45959
rect 63499 45913 63577 45959
rect 63623 45913 63701 45959
rect 63747 45913 63825 45959
rect 63871 45913 63949 45959
rect 63995 45913 64073 45959
rect 64119 45913 64197 45959
rect 64243 45913 64321 45959
rect 64367 45913 64445 45959
rect 64491 45913 64569 45959
rect 64615 45913 64693 45959
rect 64739 45913 64817 45959
rect 64863 45913 64941 45959
rect 64987 45913 65065 45959
rect 65111 45913 65189 45959
rect 65235 45913 65313 45959
rect 65359 45913 65437 45959
rect 65483 45913 65561 45959
rect 65607 45913 65685 45959
rect 65731 45913 65809 45959
rect 65855 45913 65933 45959
rect 65979 45913 66057 45959
rect 66103 45913 66181 45959
rect 66227 45913 66305 45959
rect 66351 45913 66429 45959
rect 66475 45913 66553 45959
rect 66599 45913 66677 45959
rect 66723 45913 66801 45959
rect 66847 45913 66925 45959
rect 66971 45913 67049 45959
rect 67095 45913 67173 45959
rect 67219 45913 67297 45959
rect 67343 45913 67421 45959
rect 67467 45913 67545 45959
rect 67591 45913 67669 45959
rect 67715 45913 67793 45959
rect 67839 45913 67917 45959
rect 67963 45913 68041 45959
rect 68087 45913 68165 45959
rect 68211 45913 68289 45959
rect 68335 45913 68413 45959
rect 68459 45913 68537 45959
rect 68583 45913 68661 45959
rect 68707 45913 68785 45959
rect 68831 45913 68909 45959
rect 68955 45913 69033 45959
rect 69079 45913 69157 45959
rect 69203 45913 69281 45959
rect 69327 45913 69405 45959
rect 69451 45913 69529 45959
rect 69575 45913 69653 45959
rect 69699 45913 69777 45959
rect 69823 45913 69901 45959
rect 69947 45913 70025 45959
rect 70071 45913 70149 45959
rect 70195 45913 70273 45959
rect 70319 45913 70397 45959
rect 70443 45913 70521 45959
rect 70567 45913 70645 45959
rect 70691 45913 70769 45959
rect 70815 45913 70893 45959
rect 70939 45913 71017 45959
rect 71063 45913 71141 45959
rect 71187 45913 71265 45959
rect 71311 45913 71389 45959
rect 71435 45913 71513 45959
rect 71559 45913 71637 45959
rect 71683 45913 71761 45959
rect 71807 45913 71885 45959
rect 71931 45913 72009 45959
rect 72055 45913 72133 45959
rect 72179 45913 72257 45959
rect 72303 45913 72381 45959
rect 72427 45913 72505 45959
rect 72551 45913 72629 45959
rect 72675 45913 72753 45959
rect 72799 45913 72877 45959
rect 72923 45913 73001 45959
rect 73047 45913 73125 45959
rect 73171 45913 73249 45959
rect 73295 45913 73373 45959
rect 73419 45913 73497 45959
rect 73543 45913 73621 45959
rect 73667 45913 73745 45959
rect 73791 45913 73869 45959
rect 73915 45913 73993 45959
rect 74039 45913 74117 45959
rect 74163 45913 74241 45959
rect 74287 45913 74365 45959
rect 74411 45913 74489 45959
rect 74535 45913 74613 45959
rect 74659 45913 74737 45959
rect 74783 45913 74861 45959
rect 74907 45913 74985 45959
rect 75031 45913 75109 45959
rect 75155 45913 75233 45959
rect 75279 45913 75357 45959
rect 75403 45913 75481 45959
rect 75527 45913 75605 45959
rect 75651 45913 75729 45959
rect 75775 45913 75853 45959
rect 75899 45913 75977 45959
rect 76023 45913 76101 45959
rect 76147 45913 76225 45959
rect 76271 45913 76349 45959
rect 76395 45913 76473 45959
rect 76519 45913 76597 45959
rect 76643 45913 76721 45959
rect 76767 45913 76845 45959
rect 76891 45913 76969 45959
rect 77015 45913 77093 45959
rect 77139 45913 77217 45959
rect 77263 45913 77341 45959
rect 77387 45913 77465 45959
rect 77511 45913 77589 45959
rect 77635 45913 77713 45959
rect 77759 45913 77837 45959
rect 77883 45913 77961 45959
rect 78007 45913 78085 45959
rect 78131 45913 78209 45959
rect 78255 45913 78333 45959
rect 78379 45913 78457 45959
rect 78503 45913 78581 45959
rect 78627 45913 78705 45959
rect 78751 45913 78829 45959
rect 78875 45913 78953 45959
rect 78999 45913 79077 45959
rect 79123 45913 79201 45959
rect 79247 45913 79325 45959
rect 79371 45913 79449 45959
rect 79495 45913 79573 45959
rect 79619 45913 79697 45959
rect 79743 45913 79821 45959
rect 79867 45913 79945 45959
rect 79991 45913 80069 45959
rect 80115 45913 80193 45959
rect 80239 45913 80317 45959
rect 80363 45913 80441 45959
rect 80487 45913 80565 45959
rect 80611 45913 80689 45959
rect 80735 45913 80813 45959
rect 80859 45913 80937 45959
rect 80983 45913 81061 45959
rect 81107 45913 81185 45959
rect 81231 45913 81309 45959
rect 81355 45913 81433 45959
rect 81479 45913 81557 45959
rect 81603 45913 81681 45959
rect 81727 45913 81805 45959
rect 81851 45913 81929 45959
rect 81975 45913 82053 45959
rect 82099 45913 82177 45959
rect 82223 45913 82301 45959
rect 82347 45913 82425 45959
rect 82471 45913 82549 45959
rect 82595 45913 82673 45959
rect 82719 45913 82797 45959
rect 82843 45913 82921 45959
rect 82967 45913 83045 45959
rect 83091 45913 83169 45959
rect 83215 45913 83293 45959
rect 83339 45913 83417 45959
rect 83463 45913 83541 45959
rect 83587 45913 83665 45959
rect 83711 45913 83789 45959
rect 83835 45913 83913 45959
rect 83959 45913 84037 45959
rect 84083 45913 84161 45959
rect 84207 45913 84285 45959
rect 84331 45913 84409 45959
rect 84455 45913 84533 45959
rect 84579 45913 84657 45959
rect 84703 45913 84781 45959
rect 84827 45913 84905 45959
rect 84951 45913 85029 45959
rect 85075 45913 85153 45959
rect 85199 45913 85277 45959
rect 85323 45913 85401 45959
rect 85447 45913 85525 45959
rect 85571 45913 85649 45959
rect 85695 45913 85706 45959
rect 0 45835 85706 45913
rect 0 45789 89 45835
rect 135 45789 213 45835
rect 259 45789 337 45835
rect 383 45789 461 45835
rect 507 45789 585 45835
rect 631 45789 709 45835
rect 755 45789 833 45835
rect 879 45789 957 45835
rect 1003 45789 1081 45835
rect 1127 45789 1205 45835
rect 1251 45789 1329 45835
rect 1375 45789 1453 45835
rect 1499 45789 1577 45835
rect 1623 45789 1701 45835
rect 1747 45789 1825 45835
rect 1871 45789 1949 45835
rect 1995 45789 2073 45835
rect 2119 45789 2197 45835
rect 2243 45789 2321 45835
rect 2367 45789 2445 45835
rect 2491 45789 2569 45835
rect 2615 45789 2693 45835
rect 2739 45789 2817 45835
rect 2863 45789 2941 45835
rect 2987 45789 3065 45835
rect 3111 45789 3189 45835
rect 3235 45789 3313 45835
rect 3359 45789 3437 45835
rect 3483 45789 3561 45835
rect 3607 45789 3685 45835
rect 3731 45789 3809 45835
rect 3855 45789 3933 45835
rect 3979 45789 4057 45835
rect 4103 45789 4181 45835
rect 4227 45789 4305 45835
rect 4351 45789 4429 45835
rect 4475 45789 4553 45835
rect 4599 45789 4677 45835
rect 4723 45789 4801 45835
rect 4847 45789 4925 45835
rect 4971 45789 5049 45835
rect 5095 45789 5173 45835
rect 5219 45789 5297 45835
rect 5343 45789 5421 45835
rect 5467 45789 5545 45835
rect 5591 45789 5669 45835
rect 5715 45789 5793 45835
rect 5839 45789 5917 45835
rect 5963 45789 6041 45835
rect 6087 45789 6165 45835
rect 6211 45789 6289 45835
rect 6335 45789 6413 45835
rect 6459 45789 6537 45835
rect 6583 45789 6661 45835
rect 6707 45789 6785 45835
rect 6831 45789 6909 45835
rect 6955 45789 7033 45835
rect 7079 45789 7157 45835
rect 7203 45789 7281 45835
rect 7327 45789 7405 45835
rect 7451 45789 7529 45835
rect 7575 45789 7653 45835
rect 7699 45789 7777 45835
rect 7823 45789 7901 45835
rect 7947 45789 8025 45835
rect 8071 45789 8149 45835
rect 8195 45789 8273 45835
rect 8319 45789 8397 45835
rect 8443 45789 8521 45835
rect 8567 45789 8645 45835
rect 8691 45789 8769 45835
rect 8815 45789 8893 45835
rect 8939 45789 9017 45835
rect 9063 45789 9141 45835
rect 9187 45789 9265 45835
rect 9311 45789 9389 45835
rect 9435 45789 9513 45835
rect 9559 45789 9637 45835
rect 9683 45789 9761 45835
rect 9807 45789 9885 45835
rect 9931 45789 10009 45835
rect 10055 45789 10133 45835
rect 10179 45789 10257 45835
rect 10303 45789 10381 45835
rect 10427 45789 10505 45835
rect 10551 45789 10629 45835
rect 10675 45789 10753 45835
rect 10799 45789 10877 45835
rect 10923 45789 11001 45835
rect 11047 45789 11125 45835
rect 11171 45789 11249 45835
rect 11295 45789 11373 45835
rect 11419 45789 11497 45835
rect 11543 45789 11621 45835
rect 11667 45789 11745 45835
rect 11791 45789 11869 45835
rect 11915 45789 11993 45835
rect 12039 45789 12117 45835
rect 12163 45789 12241 45835
rect 12287 45789 12365 45835
rect 12411 45789 12489 45835
rect 12535 45789 12613 45835
rect 12659 45789 12737 45835
rect 12783 45789 12861 45835
rect 12907 45789 12985 45835
rect 13031 45789 13109 45835
rect 13155 45789 13233 45835
rect 13279 45789 13357 45835
rect 13403 45789 13481 45835
rect 13527 45789 13605 45835
rect 13651 45789 13729 45835
rect 13775 45789 13853 45835
rect 13899 45789 13977 45835
rect 14023 45789 14101 45835
rect 14147 45789 14225 45835
rect 14271 45789 14349 45835
rect 14395 45789 14473 45835
rect 14519 45789 14597 45835
rect 14643 45789 14721 45835
rect 14767 45789 14845 45835
rect 14891 45789 14969 45835
rect 15015 45789 15093 45835
rect 15139 45789 15217 45835
rect 15263 45789 15341 45835
rect 15387 45789 15465 45835
rect 15511 45789 15589 45835
rect 15635 45789 15713 45835
rect 15759 45789 15837 45835
rect 15883 45789 15961 45835
rect 16007 45789 16085 45835
rect 16131 45789 16209 45835
rect 16255 45789 16333 45835
rect 16379 45789 16457 45835
rect 16503 45789 16581 45835
rect 16627 45789 16705 45835
rect 16751 45789 16829 45835
rect 16875 45789 16953 45835
rect 16999 45789 17077 45835
rect 17123 45789 17201 45835
rect 17247 45789 17325 45835
rect 17371 45789 17449 45835
rect 17495 45789 17573 45835
rect 17619 45789 17697 45835
rect 17743 45789 17821 45835
rect 17867 45789 17945 45835
rect 17991 45789 18069 45835
rect 18115 45789 18193 45835
rect 18239 45789 18317 45835
rect 18363 45789 18441 45835
rect 18487 45789 18565 45835
rect 18611 45789 18689 45835
rect 18735 45789 18813 45835
rect 18859 45789 18937 45835
rect 18983 45789 19061 45835
rect 19107 45789 19185 45835
rect 19231 45789 19309 45835
rect 19355 45789 19433 45835
rect 19479 45789 19557 45835
rect 19603 45789 19681 45835
rect 19727 45789 19805 45835
rect 19851 45789 19929 45835
rect 19975 45789 20053 45835
rect 20099 45789 20177 45835
rect 20223 45789 20301 45835
rect 20347 45789 20425 45835
rect 20471 45789 20549 45835
rect 20595 45789 20673 45835
rect 20719 45789 20797 45835
rect 20843 45789 20921 45835
rect 20967 45789 21045 45835
rect 21091 45789 21169 45835
rect 21215 45789 21293 45835
rect 21339 45789 21417 45835
rect 21463 45789 21541 45835
rect 21587 45789 21665 45835
rect 21711 45789 21789 45835
rect 21835 45789 21913 45835
rect 21959 45789 22037 45835
rect 22083 45789 22161 45835
rect 22207 45789 22285 45835
rect 22331 45789 22409 45835
rect 22455 45789 22533 45835
rect 22579 45789 22657 45835
rect 22703 45789 22781 45835
rect 22827 45789 22905 45835
rect 22951 45789 23029 45835
rect 23075 45789 23153 45835
rect 23199 45789 23277 45835
rect 23323 45789 23401 45835
rect 23447 45789 23525 45835
rect 23571 45789 23649 45835
rect 23695 45789 23773 45835
rect 23819 45789 23897 45835
rect 23943 45789 24021 45835
rect 24067 45789 24145 45835
rect 24191 45789 24269 45835
rect 24315 45789 24393 45835
rect 24439 45789 24517 45835
rect 24563 45789 24641 45835
rect 24687 45789 24765 45835
rect 24811 45789 24889 45835
rect 24935 45789 25013 45835
rect 25059 45789 25137 45835
rect 25183 45789 25261 45835
rect 25307 45789 25385 45835
rect 25431 45789 25509 45835
rect 25555 45789 25633 45835
rect 25679 45789 25757 45835
rect 25803 45789 25881 45835
rect 25927 45789 26005 45835
rect 26051 45789 26129 45835
rect 26175 45789 26253 45835
rect 26299 45789 26377 45835
rect 26423 45789 26501 45835
rect 26547 45789 26625 45835
rect 26671 45789 26749 45835
rect 26795 45789 26873 45835
rect 26919 45789 26997 45835
rect 27043 45789 27121 45835
rect 27167 45789 27245 45835
rect 27291 45789 27369 45835
rect 27415 45789 27493 45835
rect 27539 45789 27617 45835
rect 27663 45789 27741 45835
rect 27787 45789 27865 45835
rect 27911 45789 27989 45835
rect 28035 45789 28113 45835
rect 28159 45789 28237 45835
rect 28283 45789 28361 45835
rect 28407 45789 28485 45835
rect 28531 45789 28609 45835
rect 28655 45789 28733 45835
rect 28779 45789 28857 45835
rect 28903 45789 28981 45835
rect 29027 45789 29105 45835
rect 29151 45789 29229 45835
rect 29275 45789 29353 45835
rect 29399 45789 29477 45835
rect 29523 45789 29601 45835
rect 29647 45789 29725 45835
rect 29771 45789 29849 45835
rect 29895 45789 29973 45835
rect 30019 45789 30097 45835
rect 30143 45789 30221 45835
rect 30267 45789 30345 45835
rect 30391 45789 30469 45835
rect 30515 45789 30593 45835
rect 30639 45789 30717 45835
rect 30763 45789 30841 45835
rect 30887 45789 30965 45835
rect 31011 45789 31089 45835
rect 31135 45789 31213 45835
rect 31259 45789 31337 45835
rect 31383 45789 31461 45835
rect 31507 45789 31585 45835
rect 31631 45789 31709 45835
rect 31755 45789 31833 45835
rect 31879 45789 31957 45835
rect 32003 45789 32081 45835
rect 32127 45789 32205 45835
rect 32251 45789 32329 45835
rect 32375 45789 32453 45835
rect 32499 45789 32577 45835
rect 32623 45789 32701 45835
rect 32747 45789 32825 45835
rect 32871 45789 32949 45835
rect 32995 45789 33073 45835
rect 33119 45789 33197 45835
rect 33243 45789 33321 45835
rect 33367 45789 33445 45835
rect 33491 45789 33569 45835
rect 33615 45789 33693 45835
rect 33739 45789 33817 45835
rect 33863 45789 33941 45835
rect 33987 45789 34065 45835
rect 34111 45789 34189 45835
rect 34235 45789 34313 45835
rect 34359 45789 34437 45835
rect 34483 45789 34561 45835
rect 34607 45789 34685 45835
rect 34731 45789 34809 45835
rect 34855 45789 34933 45835
rect 34979 45789 35057 45835
rect 35103 45789 35181 45835
rect 35227 45789 35305 45835
rect 35351 45789 35429 45835
rect 35475 45789 35553 45835
rect 35599 45789 35677 45835
rect 35723 45789 35801 45835
rect 35847 45789 35925 45835
rect 35971 45789 36049 45835
rect 36095 45789 36173 45835
rect 36219 45789 36297 45835
rect 36343 45789 36421 45835
rect 36467 45789 36545 45835
rect 36591 45789 36669 45835
rect 36715 45789 36793 45835
rect 36839 45789 36917 45835
rect 36963 45789 37041 45835
rect 37087 45789 37165 45835
rect 37211 45789 37289 45835
rect 37335 45789 37413 45835
rect 37459 45789 37537 45835
rect 37583 45789 37661 45835
rect 37707 45789 37785 45835
rect 37831 45789 37909 45835
rect 37955 45789 38033 45835
rect 38079 45789 38157 45835
rect 38203 45789 38281 45835
rect 38327 45789 38405 45835
rect 38451 45789 38529 45835
rect 38575 45789 38653 45835
rect 38699 45789 38777 45835
rect 38823 45789 38901 45835
rect 38947 45789 39025 45835
rect 39071 45789 39149 45835
rect 39195 45789 39273 45835
rect 39319 45789 39397 45835
rect 39443 45789 39521 45835
rect 39567 45789 39645 45835
rect 39691 45789 39769 45835
rect 39815 45789 39893 45835
rect 39939 45789 40017 45835
rect 40063 45789 40141 45835
rect 40187 45789 40265 45835
rect 40311 45789 40389 45835
rect 40435 45789 40513 45835
rect 40559 45789 40637 45835
rect 40683 45789 40761 45835
rect 40807 45789 40885 45835
rect 40931 45789 41009 45835
rect 41055 45789 41133 45835
rect 41179 45789 41257 45835
rect 41303 45789 41381 45835
rect 41427 45789 41505 45835
rect 41551 45789 41629 45835
rect 41675 45789 41753 45835
rect 41799 45789 41877 45835
rect 41923 45789 42001 45835
rect 42047 45789 42125 45835
rect 42171 45789 42249 45835
rect 42295 45789 42373 45835
rect 42419 45789 42497 45835
rect 42543 45789 42621 45835
rect 42667 45789 42745 45835
rect 42791 45789 42869 45835
rect 42915 45789 42993 45835
rect 43039 45789 43117 45835
rect 43163 45789 43241 45835
rect 43287 45789 43365 45835
rect 43411 45789 43489 45835
rect 43535 45789 43613 45835
rect 43659 45789 43737 45835
rect 43783 45789 43861 45835
rect 43907 45789 43985 45835
rect 44031 45789 44109 45835
rect 44155 45789 44233 45835
rect 44279 45789 44357 45835
rect 44403 45789 44481 45835
rect 44527 45789 44605 45835
rect 44651 45789 44729 45835
rect 44775 45789 44853 45835
rect 44899 45789 44977 45835
rect 45023 45789 45101 45835
rect 45147 45789 45225 45835
rect 45271 45789 45349 45835
rect 45395 45789 45473 45835
rect 45519 45789 45597 45835
rect 45643 45789 45721 45835
rect 45767 45789 45845 45835
rect 45891 45789 45969 45835
rect 46015 45789 46093 45835
rect 46139 45789 46217 45835
rect 46263 45789 46341 45835
rect 46387 45789 46465 45835
rect 46511 45789 46589 45835
rect 46635 45789 46713 45835
rect 46759 45789 46837 45835
rect 46883 45789 46961 45835
rect 47007 45789 47085 45835
rect 47131 45789 47209 45835
rect 47255 45789 47333 45835
rect 47379 45789 47457 45835
rect 47503 45789 47581 45835
rect 47627 45789 47705 45835
rect 47751 45789 47829 45835
rect 47875 45789 47953 45835
rect 47999 45789 48077 45835
rect 48123 45789 48201 45835
rect 48247 45789 48325 45835
rect 48371 45789 48449 45835
rect 48495 45789 48573 45835
rect 48619 45789 48697 45835
rect 48743 45789 48821 45835
rect 48867 45789 48945 45835
rect 48991 45789 49069 45835
rect 49115 45789 49193 45835
rect 49239 45789 49317 45835
rect 49363 45789 49441 45835
rect 49487 45789 49565 45835
rect 49611 45789 49689 45835
rect 49735 45789 49813 45835
rect 49859 45789 49937 45835
rect 49983 45789 50061 45835
rect 50107 45789 50185 45835
rect 50231 45789 50309 45835
rect 50355 45789 50433 45835
rect 50479 45789 50557 45835
rect 50603 45789 50681 45835
rect 50727 45789 50805 45835
rect 50851 45789 50929 45835
rect 50975 45789 51053 45835
rect 51099 45789 51177 45835
rect 51223 45789 51301 45835
rect 51347 45789 51425 45835
rect 51471 45789 51549 45835
rect 51595 45789 51673 45835
rect 51719 45789 51797 45835
rect 51843 45789 51921 45835
rect 51967 45789 52045 45835
rect 52091 45789 52169 45835
rect 52215 45789 52293 45835
rect 52339 45789 52417 45835
rect 52463 45789 52541 45835
rect 52587 45789 52665 45835
rect 52711 45789 52789 45835
rect 52835 45789 52913 45835
rect 52959 45789 53037 45835
rect 53083 45789 53161 45835
rect 53207 45789 53285 45835
rect 53331 45789 53409 45835
rect 53455 45789 53533 45835
rect 53579 45789 53657 45835
rect 53703 45789 53781 45835
rect 53827 45789 53905 45835
rect 53951 45789 54029 45835
rect 54075 45789 54153 45835
rect 54199 45789 54277 45835
rect 54323 45789 54401 45835
rect 54447 45789 54525 45835
rect 54571 45789 54649 45835
rect 54695 45789 54773 45835
rect 54819 45789 54897 45835
rect 54943 45789 55021 45835
rect 55067 45789 55145 45835
rect 55191 45789 55269 45835
rect 55315 45789 55393 45835
rect 55439 45789 55517 45835
rect 55563 45789 55641 45835
rect 55687 45789 55765 45835
rect 55811 45789 55889 45835
rect 55935 45789 56013 45835
rect 56059 45789 56137 45835
rect 56183 45789 56261 45835
rect 56307 45789 56385 45835
rect 56431 45789 56509 45835
rect 56555 45789 56633 45835
rect 56679 45789 56757 45835
rect 56803 45789 56881 45835
rect 56927 45789 57005 45835
rect 57051 45789 57129 45835
rect 57175 45789 57253 45835
rect 57299 45789 57377 45835
rect 57423 45789 57501 45835
rect 57547 45789 57625 45835
rect 57671 45789 57749 45835
rect 57795 45789 57873 45835
rect 57919 45789 57997 45835
rect 58043 45789 58121 45835
rect 58167 45789 58245 45835
rect 58291 45789 58369 45835
rect 58415 45789 58493 45835
rect 58539 45789 58617 45835
rect 58663 45789 58741 45835
rect 58787 45789 58865 45835
rect 58911 45789 58989 45835
rect 59035 45789 59113 45835
rect 59159 45789 59237 45835
rect 59283 45789 59361 45835
rect 59407 45789 59485 45835
rect 59531 45789 59609 45835
rect 59655 45789 59733 45835
rect 59779 45789 59857 45835
rect 59903 45789 59981 45835
rect 60027 45789 60105 45835
rect 60151 45789 60229 45835
rect 60275 45789 60353 45835
rect 60399 45789 60477 45835
rect 60523 45789 60601 45835
rect 60647 45789 60725 45835
rect 60771 45789 60849 45835
rect 60895 45789 60973 45835
rect 61019 45789 61097 45835
rect 61143 45789 61221 45835
rect 61267 45789 61345 45835
rect 61391 45789 61469 45835
rect 61515 45789 61593 45835
rect 61639 45789 61717 45835
rect 61763 45789 61841 45835
rect 61887 45789 61965 45835
rect 62011 45789 62089 45835
rect 62135 45789 62213 45835
rect 62259 45789 62337 45835
rect 62383 45789 62461 45835
rect 62507 45789 62585 45835
rect 62631 45789 62709 45835
rect 62755 45789 62833 45835
rect 62879 45789 62957 45835
rect 63003 45789 63081 45835
rect 63127 45789 63205 45835
rect 63251 45789 63329 45835
rect 63375 45789 63453 45835
rect 63499 45789 63577 45835
rect 63623 45789 63701 45835
rect 63747 45789 63825 45835
rect 63871 45789 63949 45835
rect 63995 45789 64073 45835
rect 64119 45789 64197 45835
rect 64243 45789 64321 45835
rect 64367 45789 64445 45835
rect 64491 45789 64569 45835
rect 64615 45789 64693 45835
rect 64739 45789 64817 45835
rect 64863 45789 64941 45835
rect 64987 45789 65065 45835
rect 65111 45789 65189 45835
rect 65235 45789 65313 45835
rect 65359 45789 65437 45835
rect 65483 45789 65561 45835
rect 65607 45789 65685 45835
rect 65731 45789 65809 45835
rect 65855 45789 65933 45835
rect 65979 45789 66057 45835
rect 66103 45789 66181 45835
rect 66227 45789 66305 45835
rect 66351 45789 66429 45835
rect 66475 45789 66553 45835
rect 66599 45789 66677 45835
rect 66723 45789 66801 45835
rect 66847 45789 66925 45835
rect 66971 45789 67049 45835
rect 67095 45789 67173 45835
rect 67219 45789 67297 45835
rect 67343 45789 67421 45835
rect 67467 45789 67545 45835
rect 67591 45789 67669 45835
rect 67715 45789 67793 45835
rect 67839 45789 67917 45835
rect 67963 45789 68041 45835
rect 68087 45789 68165 45835
rect 68211 45789 68289 45835
rect 68335 45789 68413 45835
rect 68459 45789 68537 45835
rect 68583 45789 68661 45835
rect 68707 45789 68785 45835
rect 68831 45789 68909 45835
rect 68955 45789 69033 45835
rect 69079 45789 69157 45835
rect 69203 45789 69281 45835
rect 69327 45789 69405 45835
rect 69451 45789 69529 45835
rect 69575 45789 69653 45835
rect 69699 45789 69777 45835
rect 69823 45789 69901 45835
rect 69947 45789 70025 45835
rect 70071 45789 70149 45835
rect 70195 45789 70273 45835
rect 70319 45789 70397 45835
rect 70443 45789 70521 45835
rect 70567 45789 70645 45835
rect 70691 45789 70769 45835
rect 70815 45789 70893 45835
rect 70939 45789 71017 45835
rect 71063 45789 71141 45835
rect 71187 45789 71265 45835
rect 71311 45789 71389 45835
rect 71435 45789 71513 45835
rect 71559 45789 71637 45835
rect 71683 45789 71761 45835
rect 71807 45789 71885 45835
rect 71931 45789 72009 45835
rect 72055 45789 72133 45835
rect 72179 45789 72257 45835
rect 72303 45789 72381 45835
rect 72427 45789 72505 45835
rect 72551 45789 72629 45835
rect 72675 45789 72753 45835
rect 72799 45789 72877 45835
rect 72923 45789 73001 45835
rect 73047 45789 73125 45835
rect 73171 45789 73249 45835
rect 73295 45789 73373 45835
rect 73419 45789 73497 45835
rect 73543 45789 73621 45835
rect 73667 45789 73745 45835
rect 73791 45789 73869 45835
rect 73915 45789 73993 45835
rect 74039 45789 74117 45835
rect 74163 45789 74241 45835
rect 74287 45789 74365 45835
rect 74411 45789 74489 45835
rect 74535 45789 74613 45835
rect 74659 45789 74737 45835
rect 74783 45789 74861 45835
rect 74907 45789 74985 45835
rect 75031 45789 75109 45835
rect 75155 45789 75233 45835
rect 75279 45789 75357 45835
rect 75403 45789 75481 45835
rect 75527 45789 75605 45835
rect 75651 45789 75729 45835
rect 75775 45789 75853 45835
rect 75899 45789 75977 45835
rect 76023 45789 76101 45835
rect 76147 45789 76225 45835
rect 76271 45789 76349 45835
rect 76395 45789 76473 45835
rect 76519 45789 76597 45835
rect 76643 45789 76721 45835
rect 76767 45789 76845 45835
rect 76891 45789 76969 45835
rect 77015 45789 77093 45835
rect 77139 45789 77217 45835
rect 77263 45789 77341 45835
rect 77387 45789 77465 45835
rect 77511 45789 77589 45835
rect 77635 45789 77713 45835
rect 77759 45789 77837 45835
rect 77883 45789 77961 45835
rect 78007 45789 78085 45835
rect 78131 45789 78209 45835
rect 78255 45789 78333 45835
rect 78379 45789 78457 45835
rect 78503 45789 78581 45835
rect 78627 45789 78705 45835
rect 78751 45789 78829 45835
rect 78875 45789 78953 45835
rect 78999 45789 79077 45835
rect 79123 45789 79201 45835
rect 79247 45789 79325 45835
rect 79371 45789 79449 45835
rect 79495 45789 79573 45835
rect 79619 45789 79697 45835
rect 79743 45789 79821 45835
rect 79867 45789 79945 45835
rect 79991 45789 80069 45835
rect 80115 45789 80193 45835
rect 80239 45789 80317 45835
rect 80363 45789 80441 45835
rect 80487 45789 80565 45835
rect 80611 45789 80689 45835
rect 80735 45789 80813 45835
rect 80859 45789 80937 45835
rect 80983 45789 81061 45835
rect 81107 45789 81185 45835
rect 81231 45789 81309 45835
rect 81355 45789 81433 45835
rect 81479 45789 81557 45835
rect 81603 45789 81681 45835
rect 81727 45789 81805 45835
rect 81851 45789 81929 45835
rect 81975 45789 82053 45835
rect 82099 45789 82177 45835
rect 82223 45789 82301 45835
rect 82347 45789 82425 45835
rect 82471 45789 82549 45835
rect 82595 45789 82673 45835
rect 82719 45789 82797 45835
rect 82843 45789 82921 45835
rect 82967 45789 83045 45835
rect 83091 45789 83169 45835
rect 83215 45789 83293 45835
rect 83339 45789 83417 45835
rect 83463 45789 83541 45835
rect 83587 45789 83665 45835
rect 83711 45789 83789 45835
rect 83835 45789 83913 45835
rect 83959 45789 84037 45835
rect 84083 45789 84161 45835
rect 84207 45789 84285 45835
rect 84331 45789 84409 45835
rect 84455 45789 84533 45835
rect 84579 45789 84657 45835
rect 84703 45789 84781 45835
rect 84827 45789 84905 45835
rect 84951 45789 85029 45835
rect 85075 45789 85153 45835
rect 85199 45789 85277 45835
rect 85323 45789 85401 45835
rect 85447 45789 85525 45835
rect 85571 45789 85649 45835
rect 85695 45789 85706 45835
rect 0 45711 85706 45789
rect 0 45665 89 45711
rect 135 45665 213 45711
rect 259 45665 337 45711
rect 383 45665 461 45711
rect 507 45665 585 45711
rect 631 45665 709 45711
rect 755 45665 833 45711
rect 879 45665 957 45711
rect 1003 45665 1081 45711
rect 1127 45665 1205 45711
rect 1251 45665 1329 45711
rect 1375 45665 1453 45711
rect 1499 45665 1577 45711
rect 1623 45665 1701 45711
rect 1747 45665 1825 45711
rect 1871 45665 1949 45711
rect 1995 45665 2073 45711
rect 2119 45665 2197 45711
rect 2243 45665 2321 45711
rect 2367 45665 2445 45711
rect 2491 45665 2569 45711
rect 2615 45665 2693 45711
rect 2739 45665 2817 45711
rect 2863 45665 2941 45711
rect 2987 45665 3065 45711
rect 3111 45665 3189 45711
rect 3235 45665 3313 45711
rect 3359 45665 3437 45711
rect 3483 45665 3561 45711
rect 3607 45665 3685 45711
rect 3731 45665 3809 45711
rect 3855 45665 3933 45711
rect 3979 45665 4057 45711
rect 4103 45665 4181 45711
rect 4227 45665 4305 45711
rect 4351 45665 4429 45711
rect 4475 45665 4553 45711
rect 4599 45665 4677 45711
rect 4723 45665 4801 45711
rect 4847 45665 4925 45711
rect 4971 45665 5049 45711
rect 5095 45665 5173 45711
rect 5219 45665 5297 45711
rect 5343 45665 5421 45711
rect 5467 45665 5545 45711
rect 5591 45665 5669 45711
rect 5715 45665 5793 45711
rect 5839 45665 5917 45711
rect 5963 45665 6041 45711
rect 6087 45665 6165 45711
rect 6211 45665 6289 45711
rect 6335 45665 6413 45711
rect 6459 45665 6537 45711
rect 6583 45665 6661 45711
rect 6707 45665 6785 45711
rect 6831 45665 6909 45711
rect 6955 45665 7033 45711
rect 7079 45665 7157 45711
rect 7203 45665 7281 45711
rect 7327 45665 7405 45711
rect 7451 45665 7529 45711
rect 7575 45665 7653 45711
rect 7699 45665 7777 45711
rect 7823 45665 7901 45711
rect 7947 45665 8025 45711
rect 8071 45665 8149 45711
rect 8195 45665 8273 45711
rect 8319 45665 8397 45711
rect 8443 45665 8521 45711
rect 8567 45665 8645 45711
rect 8691 45665 8769 45711
rect 8815 45665 8893 45711
rect 8939 45665 9017 45711
rect 9063 45665 9141 45711
rect 9187 45665 9265 45711
rect 9311 45665 9389 45711
rect 9435 45665 9513 45711
rect 9559 45665 9637 45711
rect 9683 45665 9761 45711
rect 9807 45665 9885 45711
rect 9931 45665 10009 45711
rect 10055 45665 10133 45711
rect 10179 45665 10257 45711
rect 10303 45665 10381 45711
rect 10427 45665 10505 45711
rect 10551 45665 10629 45711
rect 10675 45665 10753 45711
rect 10799 45665 10877 45711
rect 10923 45665 11001 45711
rect 11047 45665 11125 45711
rect 11171 45665 11249 45711
rect 11295 45665 11373 45711
rect 11419 45665 11497 45711
rect 11543 45665 11621 45711
rect 11667 45665 11745 45711
rect 11791 45665 11869 45711
rect 11915 45665 11993 45711
rect 12039 45665 12117 45711
rect 12163 45665 12241 45711
rect 12287 45665 12365 45711
rect 12411 45665 12489 45711
rect 12535 45665 12613 45711
rect 12659 45665 12737 45711
rect 12783 45665 12861 45711
rect 12907 45665 12985 45711
rect 13031 45665 13109 45711
rect 13155 45665 13233 45711
rect 13279 45665 13357 45711
rect 13403 45665 13481 45711
rect 13527 45665 13605 45711
rect 13651 45665 13729 45711
rect 13775 45665 13853 45711
rect 13899 45665 13977 45711
rect 14023 45665 14101 45711
rect 14147 45665 14225 45711
rect 14271 45665 14349 45711
rect 14395 45665 14473 45711
rect 14519 45665 14597 45711
rect 14643 45665 14721 45711
rect 14767 45665 14845 45711
rect 14891 45665 14969 45711
rect 15015 45665 15093 45711
rect 15139 45665 15217 45711
rect 15263 45665 15341 45711
rect 15387 45665 15465 45711
rect 15511 45665 15589 45711
rect 15635 45665 15713 45711
rect 15759 45665 15837 45711
rect 15883 45665 15961 45711
rect 16007 45665 16085 45711
rect 16131 45665 16209 45711
rect 16255 45665 16333 45711
rect 16379 45665 16457 45711
rect 16503 45665 16581 45711
rect 16627 45665 16705 45711
rect 16751 45665 16829 45711
rect 16875 45665 16953 45711
rect 16999 45665 17077 45711
rect 17123 45665 17201 45711
rect 17247 45665 17325 45711
rect 17371 45665 17449 45711
rect 17495 45665 17573 45711
rect 17619 45665 17697 45711
rect 17743 45665 17821 45711
rect 17867 45665 17945 45711
rect 17991 45665 18069 45711
rect 18115 45665 18193 45711
rect 18239 45665 18317 45711
rect 18363 45665 18441 45711
rect 18487 45665 18565 45711
rect 18611 45665 18689 45711
rect 18735 45665 18813 45711
rect 18859 45665 18937 45711
rect 18983 45665 19061 45711
rect 19107 45665 19185 45711
rect 19231 45665 19309 45711
rect 19355 45665 19433 45711
rect 19479 45665 19557 45711
rect 19603 45665 19681 45711
rect 19727 45665 19805 45711
rect 19851 45665 19929 45711
rect 19975 45665 20053 45711
rect 20099 45665 20177 45711
rect 20223 45665 20301 45711
rect 20347 45665 20425 45711
rect 20471 45665 20549 45711
rect 20595 45665 20673 45711
rect 20719 45665 20797 45711
rect 20843 45665 20921 45711
rect 20967 45665 21045 45711
rect 21091 45665 21169 45711
rect 21215 45665 21293 45711
rect 21339 45665 21417 45711
rect 21463 45665 21541 45711
rect 21587 45665 21665 45711
rect 21711 45665 21789 45711
rect 21835 45665 21913 45711
rect 21959 45665 22037 45711
rect 22083 45665 22161 45711
rect 22207 45665 22285 45711
rect 22331 45665 22409 45711
rect 22455 45665 22533 45711
rect 22579 45665 22657 45711
rect 22703 45665 22781 45711
rect 22827 45665 22905 45711
rect 22951 45665 23029 45711
rect 23075 45665 23153 45711
rect 23199 45665 23277 45711
rect 23323 45665 23401 45711
rect 23447 45665 23525 45711
rect 23571 45665 23649 45711
rect 23695 45665 23773 45711
rect 23819 45665 23897 45711
rect 23943 45665 24021 45711
rect 24067 45665 24145 45711
rect 24191 45665 24269 45711
rect 24315 45665 24393 45711
rect 24439 45665 24517 45711
rect 24563 45665 24641 45711
rect 24687 45665 24765 45711
rect 24811 45665 24889 45711
rect 24935 45665 25013 45711
rect 25059 45665 25137 45711
rect 25183 45665 25261 45711
rect 25307 45665 25385 45711
rect 25431 45665 25509 45711
rect 25555 45665 25633 45711
rect 25679 45665 25757 45711
rect 25803 45665 25881 45711
rect 25927 45665 26005 45711
rect 26051 45665 26129 45711
rect 26175 45665 26253 45711
rect 26299 45665 26377 45711
rect 26423 45665 26501 45711
rect 26547 45665 26625 45711
rect 26671 45665 26749 45711
rect 26795 45665 26873 45711
rect 26919 45665 26997 45711
rect 27043 45665 27121 45711
rect 27167 45665 27245 45711
rect 27291 45665 27369 45711
rect 27415 45665 27493 45711
rect 27539 45665 27617 45711
rect 27663 45665 27741 45711
rect 27787 45665 27865 45711
rect 27911 45665 27989 45711
rect 28035 45665 28113 45711
rect 28159 45665 28237 45711
rect 28283 45665 28361 45711
rect 28407 45665 28485 45711
rect 28531 45665 28609 45711
rect 28655 45665 28733 45711
rect 28779 45665 28857 45711
rect 28903 45665 28981 45711
rect 29027 45665 29105 45711
rect 29151 45665 29229 45711
rect 29275 45665 29353 45711
rect 29399 45665 29477 45711
rect 29523 45665 29601 45711
rect 29647 45665 29725 45711
rect 29771 45665 29849 45711
rect 29895 45665 29973 45711
rect 30019 45665 30097 45711
rect 30143 45665 30221 45711
rect 30267 45665 30345 45711
rect 30391 45665 30469 45711
rect 30515 45665 30593 45711
rect 30639 45665 30717 45711
rect 30763 45665 30841 45711
rect 30887 45665 30965 45711
rect 31011 45665 31089 45711
rect 31135 45665 31213 45711
rect 31259 45665 31337 45711
rect 31383 45665 31461 45711
rect 31507 45665 31585 45711
rect 31631 45665 31709 45711
rect 31755 45665 31833 45711
rect 31879 45665 31957 45711
rect 32003 45665 32081 45711
rect 32127 45665 32205 45711
rect 32251 45665 32329 45711
rect 32375 45665 32453 45711
rect 32499 45665 32577 45711
rect 32623 45665 32701 45711
rect 32747 45665 32825 45711
rect 32871 45665 32949 45711
rect 32995 45665 33073 45711
rect 33119 45665 33197 45711
rect 33243 45665 33321 45711
rect 33367 45665 33445 45711
rect 33491 45665 33569 45711
rect 33615 45665 33693 45711
rect 33739 45665 33817 45711
rect 33863 45665 33941 45711
rect 33987 45665 34065 45711
rect 34111 45665 34189 45711
rect 34235 45665 34313 45711
rect 34359 45665 34437 45711
rect 34483 45665 34561 45711
rect 34607 45665 34685 45711
rect 34731 45665 34809 45711
rect 34855 45665 34933 45711
rect 34979 45665 35057 45711
rect 35103 45665 35181 45711
rect 35227 45665 35305 45711
rect 35351 45665 35429 45711
rect 35475 45665 35553 45711
rect 35599 45665 35677 45711
rect 35723 45665 35801 45711
rect 35847 45665 35925 45711
rect 35971 45665 36049 45711
rect 36095 45665 36173 45711
rect 36219 45665 36297 45711
rect 36343 45665 36421 45711
rect 36467 45665 36545 45711
rect 36591 45665 36669 45711
rect 36715 45665 36793 45711
rect 36839 45665 36917 45711
rect 36963 45665 37041 45711
rect 37087 45665 37165 45711
rect 37211 45665 37289 45711
rect 37335 45665 37413 45711
rect 37459 45665 37537 45711
rect 37583 45665 37661 45711
rect 37707 45665 37785 45711
rect 37831 45665 37909 45711
rect 37955 45665 38033 45711
rect 38079 45665 38157 45711
rect 38203 45665 38281 45711
rect 38327 45665 38405 45711
rect 38451 45665 38529 45711
rect 38575 45665 38653 45711
rect 38699 45665 38777 45711
rect 38823 45665 38901 45711
rect 38947 45665 39025 45711
rect 39071 45665 39149 45711
rect 39195 45665 39273 45711
rect 39319 45665 39397 45711
rect 39443 45665 39521 45711
rect 39567 45665 39645 45711
rect 39691 45665 39769 45711
rect 39815 45665 39893 45711
rect 39939 45665 40017 45711
rect 40063 45665 40141 45711
rect 40187 45665 40265 45711
rect 40311 45665 40389 45711
rect 40435 45665 40513 45711
rect 40559 45665 40637 45711
rect 40683 45665 40761 45711
rect 40807 45665 40885 45711
rect 40931 45665 41009 45711
rect 41055 45665 41133 45711
rect 41179 45665 41257 45711
rect 41303 45665 41381 45711
rect 41427 45665 41505 45711
rect 41551 45665 41629 45711
rect 41675 45665 41753 45711
rect 41799 45665 41877 45711
rect 41923 45665 42001 45711
rect 42047 45665 42125 45711
rect 42171 45665 42249 45711
rect 42295 45665 42373 45711
rect 42419 45665 42497 45711
rect 42543 45665 42621 45711
rect 42667 45665 42745 45711
rect 42791 45665 42869 45711
rect 42915 45665 42993 45711
rect 43039 45665 43117 45711
rect 43163 45665 43241 45711
rect 43287 45665 43365 45711
rect 43411 45665 43489 45711
rect 43535 45665 43613 45711
rect 43659 45665 43737 45711
rect 43783 45665 43861 45711
rect 43907 45665 43985 45711
rect 44031 45665 44109 45711
rect 44155 45665 44233 45711
rect 44279 45665 44357 45711
rect 44403 45665 44481 45711
rect 44527 45665 44605 45711
rect 44651 45665 44729 45711
rect 44775 45665 44853 45711
rect 44899 45665 44977 45711
rect 45023 45665 45101 45711
rect 45147 45665 45225 45711
rect 45271 45665 45349 45711
rect 45395 45665 45473 45711
rect 45519 45665 45597 45711
rect 45643 45665 45721 45711
rect 45767 45665 45845 45711
rect 45891 45665 45969 45711
rect 46015 45665 46093 45711
rect 46139 45665 46217 45711
rect 46263 45665 46341 45711
rect 46387 45665 46465 45711
rect 46511 45665 46589 45711
rect 46635 45665 46713 45711
rect 46759 45665 46837 45711
rect 46883 45665 46961 45711
rect 47007 45665 47085 45711
rect 47131 45665 47209 45711
rect 47255 45665 47333 45711
rect 47379 45665 47457 45711
rect 47503 45665 47581 45711
rect 47627 45665 47705 45711
rect 47751 45665 47829 45711
rect 47875 45665 47953 45711
rect 47999 45665 48077 45711
rect 48123 45665 48201 45711
rect 48247 45665 48325 45711
rect 48371 45665 48449 45711
rect 48495 45665 48573 45711
rect 48619 45665 48697 45711
rect 48743 45665 48821 45711
rect 48867 45665 48945 45711
rect 48991 45665 49069 45711
rect 49115 45665 49193 45711
rect 49239 45665 49317 45711
rect 49363 45665 49441 45711
rect 49487 45665 49565 45711
rect 49611 45665 49689 45711
rect 49735 45665 49813 45711
rect 49859 45665 49937 45711
rect 49983 45665 50061 45711
rect 50107 45665 50185 45711
rect 50231 45665 50309 45711
rect 50355 45665 50433 45711
rect 50479 45665 50557 45711
rect 50603 45665 50681 45711
rect 50727 45665 50805 45711
rect 50851 45665 50929 45711
rect 50975 45665 51053 45711
rect 51099 45665 51177 45711
rect 51223 45665 51301 45711
rect 51347 45665 51425 45711
rect 51471 45665 51549 45711
rect 51595 45665 51673 45711
rect 51719 45665 51797 45711
rect 51843 45665 51921 45711
rect 51967 45665 52045 45711
rect 52091 45665 52169 45711
rect 52215 45665 52293 45711
rect 52339 45665 52417 45711
rect 52463 45665 52541 45711
rect 52587 45665 52665 45711
rect 52711 45665 52789 45711
rect 52835 45665 52913 45711
rect 52959 45665 53037 45711
rect 53083 45665 53161 45711
rect 53207 45665 53285 45711
rect 53331 45665 53409 45711
rect 53455 45665 53533 45711
rect 53579 45665 53657 45711
rect 53703 45665 53781 45711
rect 53827 45665 53905 45711
rect 53951 45665 54029 45711
rect 54075 45665 54153 45711
rect 54199 45665 54277 45711
rect 54323 45665 54401 45711
rect 54447 45665 54525 45711
rect 54571 45665 54649 45711
rect 54695 45665 54773 45711
rect 54819 45665 54897 45711
rect 54943 45665 55021 45711
rect 55067 45665 55145 45711
rect 55191 45665 55269 45711
rect 55315 45665 55393 45711
rect 55439 45665 55517 45711
rect 55563 45665 55641 45711
rect 55687 45665 55765 45711
rect 55811 45665 55889 45711
rect 55935 45665 56013 45711
rect 56059 45665 56137 45711
rect 56183 45665 56261 45711
rect 56307 45665 56385 45711
rect 56431 45665 56509 45711
rect 56555 45665 56633 45711
rect 56679 45665 56757 45711
rect 56803 45665 56881 45711
rect 56927 45665 57005 45711
rect 57051 45665 57129 45711
rect 57175 45665 57253 45711
rect 57299 45665 57377 45711
rect 57423 45665 57501 45711
rect 57547 45665 57625 45711
rect 57671 45665 57749 45711
rect 57795 45665 57873 45711
rect 57919 45665 57997 45711
rect 58043 45665 58121 45711
rect 58167 45665 58245 45711
rect 58291 45665 58369 45711
rect 58415 45665 58493 45711
rect 58539 45665 58617 45711
rect 58663 45665 58741 45711
rect 58787 45665 58865 45711
rect 58911 45665 58989 45711
rect 59035 45665 59113 45711
rect 59159 45665 59237 45711
rect 59283 45665 59361 45711
rect 59407 45665 59485 45711
rect 59531 45665 59609 45711
rect 59655 45665 59733 45711
rect 59779 45665 59857 45711
rect 59903 45665 59981 45711
rect 60027 45665 60105 45711
rect 60151 45665 60229 45711
rect 60275 45665 60353 45711
rect 60399 45665 60477 45711
rect 60523 45665 60601 45711
rect 60647 45665 60725 45711
rect 60771 45665 60849 45711
rect 60895 45665 60973 45711
rect 61019 45665 61097 45711
rect 61143 45665 61221 45711
rect 61267 45665 61345 45711
rect 61391 45665 61469 45711
rect 61515 45665 61593 45711
rect 61639 45665 61717 45711
rect 61763 45665 61841 45711
rect 61887 45665 61965 45711
rect 62011 45665 62089 45711
rect 62135 45665 62213 45711
rect 62259 45665 62337 45711
rect 62383 45665 62461 45711
rect 62507 45665 62585 45711
rect 62631 45665 62709 45711
rect 62755 45665 62833 45711
rect 62879 45665 62957 45711
rect 63003 45665 63081 45711
rect 63127 45665 63205 45711
rect 63251 45665 63329 45711
rect 63375 45665 63453 45711
rect 63499 45665 63577 45711
rect 63623 45665 63701 45711
rect 63747 45665 63825 45711
rect 63871 45665 63949 45711
rect 63995 45665 64073 45711
rect 64119 45665 64197 45711
rect 64243 45665 64321 45711
rect 64367 45665 64445 45711
rect 64491 45665 64569 45711
rect 64615 45665 64693 45711
rect 64739 45665 64817 45711
rect 64863 45665 64941 45711
rect 64987 45665 65065 45711
rect 65111 45665 65189 45711
rect 65235 45665 65313 45711
rect 65359 45665 65437 45711
rect 65483 45665 65561 45711
rect 65607 45665 65685 45711
rect 65731 45665 65809 45711
rect 65855 45665 65933 45711
rect 65979 45665 66057 45711
rect 66103 45665 66181 45711
rect 66227 45665 66305 45711
rect 66351 45665 66429 45711
rect 66475 45665 66553 45711
rect 66599 45665 66677 45711
rect 66723 45665 66801 45711
rect 66847 45665 66925 45711
rect 66971 45665 67049 45711
rect 67095 45665 67173 45711
rect 67219 45665 67297 45711
rect 67343 45665 67421 45711
rect 67467 45665 67545 45711
rect 67591 45665 67669 45711
rect 67715 45665 67793 45711
rect 67839 45665 67917 45711
rect 67963 45665 68041 45711
rect 68087 45665 68165 45711
rect 68211 45665 68289 45711
rect 68335 45665 68413 45711
rect 68459 45665 68537 45711
rect 68583 45665 68661 45711
rect 68707 45665 68785 45711
rect 68831 45665 68909 45711
rect 68955 45665 69033 45711
rect 69079 45665 69157 45711
rect 69203 45665 69281 45711
rect 69327 45665 69405 45711
rect 69451 45665 69529 45711
rect 69575 45665 69653 45711
rect 69699 45665 69777 45711
rect 69823 45665 69901 45711
rect 69947 45665 70025 45711
rect 70071 45665 70149 45711
rect 70195 45665 70273 45711
rect 70319 45665 70397 45711
rect 70443 45665 70521 45711
rect 70567 45665 70645 45711
rect 70691 45665 70769 45711
rect 70815 45665 70893 45711
rect 70939 45665 71017 45711
rect 71063 45665 71141 45711
rect 71187 45665 71265 45711
rect 71311 45665 71389 45711
rect 71435 45665 71513 45711
rect 71559 45665 71637 45711
rect 71683 45665 71761 45711
rect 71807 45665 71885 45711
rect 71931 45665 72009 45711
rect 72055 45665 72133 45711
rect 72179 45665 72257 45711
rect 72303 45665 72381 45711
rect 72427 45665 72505 45711
rect 72551 45665 72629 45711
rect 72675 45665 72753 45711
rect 72799 45665 72877 45711
rect 72923 45665 73001 45711
rect 73047 45665 73125 45711
rect 73171 45665 73249 45711
rect 73295 45665 73373 45711
rect 73419 45665 73497 45711
rect 73543 45665 73621 45711
rect 73667 45665 73745 45711
rect 73791 45665 73869 45711
rect 73915 45665 73993 45711
rect 74039 45665 74117 45711
rect 74163 45665 74241 45711
rect 74287 45665 74365 45711
rect 74411 45665 74489 45711
rect 74535 45665 74613 45711
rect 74659 45665 74737 45711
rect 74783 45665 74861 45711
rect 74907 45665 74985 45711
rect 75031 45665 75109 45711
rect 75155 45665 75233 45711
rect 75279 45665 75357 45711
rect 75403 45665 75481 45711
rect 75527 45665 75605 45711
rect 75651 45665 75729 45711
rect 75775 45665 75853 45711
rect 75899 45665 75977 45711
rect 76023 45665 76101 45711
rect 76147 45665 76225 45711
rect 76271 45665 76349 45711
rect 76395 45665 76473 45711
rect 76519 45665 76597 45711
rect 76643 45665 76721 45711
rect 76767 45665 76845 45711
rect 76891 45665 76969 45711
rect 77015 45665 77093 45711
rect 77139 45665 77217 45711
rect 77263 45665 77341 45711
rect 77387 45665 77465 45711
rect 77511 45665 77589 45711
rect 77635 45665 77713 45711
rect 77759 45665 77837 45711
rect 77883 45665 77961 45711
rect 78007 45665 78085 45711
rect 78131 45665 78209 45711
rect 78255 45665 78333 45711
rect 78379 45665 78457 45711
rect 78503 45665 78581 45711
rect 78627 45665 78705 45711
rect 78751 45665 78829 45711
rect 78875 45665 78953 45711
rect 78999 45665 79077 45711
rect 79123 45665 79201 45711
rect 79247 45665 79325 45711
rect 79371 45665 79449 45711
rect 79495 45665 79573 45711
rect 79619 45665 79697 45711
rect 79743 45665 79821 45711
rect 79867 45665 79945 45711
rect 79991 45665 80069 45711
rect 80115 45665 80193 45711
rect 80239 45665 80317 45711
rect 80363 45665 80441 45711
rect 80487 45665 80565 45711
rect 80611 45665 80689 45711
rect 80735 45665 80813 45711
rect 80859 45665 80937 45711
rect 80983 45665 81061 45711
rect 81107 45665 81185 45711
rect 81231 45665 81309 45711
rect 81355 45665 81433 45711
rect 81479 45665 81557 45711
rect 81603 45665 81681 45711
rect 81727 45665 81805 45711
rect 81851 45665 81929 45711
rect 81975 45665 82053 45711
rect 82099 45665 82177 45711
rect 82223 45665 82301 45711
rect 82347 45665 82425 45711
rect 82471 45665 82549 45711
rect 82595 45665 82673 45711
rect 82719 45665 82797 45711
rect 82843 45665 82921 45711
rect 82967 45665 83045 45711
rect 83091 45665 83169 45711
rect 83215 45665 83293 45711
rect 83339 45665 83417 45711
rect 83463 45665 83541 45711
rect 83587 45665 83665 45711
rect 83711 45665 83789 45711
rect 83835 45665 83913 45711
rect 83959 45665 84037 45711
rect 84083 45665 84161 45711
rect 84207 45665 84285 45711
rect 84331 45665 84409 45711
rect 84455 45665 84533 45711
rect 84579 45665 84657 45711
rect 84703 45665 84781 45711
rect 84827 45665 84905 45711
rect 84951 45665 85029 45711
rect 85075 45665 85153 45711
rect 85199 45665 85277 45711
rect 85323 45665 85401 45711
rect 85447 45665 85525 45711
rect 85571 45665 85649 45711
rect 85695 45665 85706 45711
rect 0 45654 85706 45665
rect 0 45563 1000 45654
rect 0 1117 89 45563
rect 435 1117 1000 45563
rect 0 1026 1000 1117
rect 85440 45563 85808 45574
rect 85440 1117 85451 45563
rect 85797 1117 85808 45563
rect 85440 1106 85808 1117
rect 0 1015 85706 1026
rect 0 969 89 1015
rect 135 969 213 1015
rect 259 969 337 1015
rect 383 969 461 1015
rect 507 969 585 1015
rect 631 969 709 1015
rect 755 969 833 1015
rect 879 969 957 1015
rect 1003 969 1081 1015
rect 1127 969 1205 1015
rect 1251 969 1329 1015
rect 1375 969 1453 1015
rect 1499 969 1577 1015
rect 1623 969 1701 1015
rect 1747 969 1825 1015
rect 1871 969 1949 1015
rect 1995 969 2073 1015
rect 2119 969 2197 1015
rect 2243 969 2321 1015
rect 2367 969 2445 1015
rect 2491 969 2569 1015
rect 2615 969 2693 1015
rect 2739 969 2817 1015
rect 2863 969 2941 1015
rect 2987 969 3065 1015
rect 3111 969 3189 1015
rect 3235 969 3313 1015
rect 3359 969 3437 1015
rect 3483 969 3561 1015
rect 3607 969 3685 1015
rect 3731 969 3809 1015
rect 3855 969 3933 1015
rect 3979 969 4057 1015
rect 4103 969 4181 1015
rect 4227 969 4305 1015
rect 4351 969 4429 1015
rect 4475 969 4553 1015
rect 4599 969 4677 1015
rect 4723 969 4801 1015
rect 4847 969 4925 1015
rect 4971 969 5049 1015
rect 5095 969 5173 1015
rect 5219 969 5297 1015
rect 5343 969 5421 1015
rect 5467 969 5545 1015
rect 5591 969 5669 1015
rect 5715 969 5793 1015
rect 5839 969 5917 1015
rect 5963 969 6041 1015
rect 6087 969 6165 1015
rect 6211 969 6289 1015
rect 6335 969 6413 1015
rect 6459 969 6537 1015
rect 6583 969 6661 1015
rect 6707 969 6785 1015
rect 6831 969 6909 1015
rect 6955 969 7033 1015
rect 7079 969 7157 1015
rect 7203 969 7281 1015
rect 7327 969 7405 1015
rect 7451 969 7529 1015
rect 7575 969 7653 1015
rect 7699 969 7777 1015
rect 7823 969 7901 1015
rect 7947 969 8025 1015
rect 8071 969 8149 1015
rect 8195 969 8273 1015
rect 8319 969 8397 1015
rect 8443 969 8521 1015
rect 8567 969 8645 1015
rect 8691 969 8769 1015
rect 8815 969 8893 1015
rect 8939 969 9017 1015
rect 9063 969 9141 1015
rect 9187 969 9265 1015
rect 9311 969 9389 1015
rect 9435 969 9513 1015
rect 9559 969 9637 1015
rect 9683 969 9761 1015
rect 9807 969 9885 1015
rect 9931 969 10009 1015
rect 10055 969 10133 1015
rect 10179 969 10257 1015
rect 10303 969 10381 1015
rect 10427 969 10505 1015
rect 10551 969 10629 1015
rect 10675 969 10753 1015
rect 10799 969 10877 1015
rect 10923 969 11001 1015
rect 11047 969 11125 1015
rect 11171 969 11249 1015
rect 11295 969 11373 1015
rect 11419 969 11497 1015
rect 11543 969 11621 1015
rect 11667 969 11745 1015
rect 11791 969 11869 1015
rect 11915 969 11993 1015
rect 12039 969 12117 1015
rect 12163 969 12241 1015
rect 12287 969 12365 1015
rect 12411 969 12489 1015
rect 12535 969 12613 1015
rect 12659 969 12737 1015
rect 12783 969 12861 1015
rect 12907 969 12985 1015
rect 13031 969 13109 1015
rect 13155 969 13233 1015
rect 13279 969 13357 1015
rect 13403 969 13481 1015
rect 13527 969 13605 1015
rect 13651 969 13729 1015
rect 13775 969 13853 1015
rect 13899 969 13977 1015
rect 14023 969 14101 1015
rect 14147 969 14225 1015
rect 14271 969 14349 1015
rect 14395 969 14473 1015
rect 14519 969 14597 1015
rect 14643 969 14721 1015
rect 14767 969 14845 1015
rect 14891 969 14969 1015
rect 15015 969 15093 1015
rect 15139 969 15217 1015
rect 15263 969 15341 1015
rect 15387 969 15465 1015
rect 15511 969 15589 1015
rect 15635 969 15713 1015
rect 15759 969 15837 1015
rect 15883 969 15961 1015
rect 16007 969 16085 1015
rect 16131 969 16209 1015
rect 16255 969 16333 1015
rect 16379 969 16457 1015
rect 16503 969 16581 1015
rect 16627 969 16705 1015
rect 16751 969 16829 1015
rect 16875 969 16953 1015
rect 16999 969 17077 1015
rect 17123 969 17201 1015
rect 17247 969 17325 1015
rect 17371 969 17449 1015
rect 17495 969 17573 1015
rect 17619 969 17697 1015
rect 17743 969 17821 1015
rect 17867 969 17945 1015
rect 17991 969 18069 1015
rect 18115 969 18193 1015
rect 18239 969 18317 1015
rect 18363 969 18441 1015
rect 18487 969 18565 1015
rect 18611 969 18689 1015
rect 18735 969 18813 1015
rect 18859 969 18937 1015
rect 18983 969 19061 1015
rect 19107 969 19185 1015
rect 19231 969 19309 1015
rect 19355 969 19433 1015
rect 19479 969 19557 1015
rect 19603 969 19681 1015
rect 19727 969 19805 1015
rect 19851 969 19929 1015
rect 19975 969 20053 1015
rect 20099 969 20177 1015
rect 20223 969 20301 1015
rect 20347 969 20425 1015
rect 20471 969 20549 1015
rect 20595 969 20673 1015
rect 20719 969 20797 1015
rect 20843 969 20921 1015
rect 20967 969 21045 1015
rect 21091 969 21169 1015
rect 21215 969 21293 1015
rect 21339 969 21417 1015
rect 21463 969 21541 1015
rect 21587 969 21665 1015
rect 21711 969 21789 1015
rect 21835 969 21913 1015
rect 21959 969 22037 1015
rect 22083 969 22161 1015
rect 22207 969 22285 1015
rect 22331 969 22409 1015
rect 22455 969 22533 1015
rect 22579 969 22657 1015
rect 22703 969 22781 1015
rect 22827 969 22905 1015
rect 22951 969 23029 1015
rect 23075 969 23153 1015
rect 23199 969 23277 1015
rect 23323 969 23401 1015
rect 23447 969 23525 1015
rect 23571 969 23649 1015
rect 23695 969 23773 1015
rect 23819 969 23897 1015
rect 23943 969 24021 1015
rect 24067 969 24145 1015
rect 24191 969 24269 1015
rect 24315 969 24393 1015
rect 24439 969 24517 1015
rect 24563 969 24641 1015
rect 24687 969 24765 1015
rect 24811 969 24889 1015
rect 24935 969 25013 1015
rect 25059 969 25137 1015
rect 25183 969 25261 1015
rect 25307 969 25385 1015
rect 25431 969 25509 1015
rect 25555 969 25633 1015
rect 25679 969 25757 1015
rect 25803 969 25881 1015
rect 25927 969 26005 1015
rect 26051 969 26129 1015
rect 26175 969 26253 1015
rect 26299 969 26377 1015
rect 26423 969 26501 1015
rect 26547 969 26625 1015
rect 26671 969 26749 1015
rect 26795 969 26873 1015
rect 26919 969 26997 1015
rect 27043 969 27121 1015
rect 27167 969 27245 1015
rect 27291 969 27369 1015
rect 27415 969 27493 1015
rect 27539 969 27617 1015
rect 27663 969 27741 1015
rect 27787 969 27865 1015
rect 27911 969 27989 1015
rect 28035 969 28113 1015
rect 28159 969 28237 1015
rect 28283 969 28361 1015
rect 28407 969 28485 1015
rect 28531 969 28609 1015
rect 28655 969 28733 1015
rect 28779 969 28857 1015
rect 28903 969 28981 1015
rect 29027 969 29105 1015
rect 29151 969 29229 1015
rect 29275 969 29353 1015
rect 29399 969 29477 1015
rect 29523 969 29601 1015
rect 29647 969 29725 1015
rect 29771 969 29849 1015
rect 29895 969 29973 1015
rect 30019 969 30097 1015
rect 30143 969 30221 1015
rect 30267 969 30345 1015
rect 30391 969 30469 1015
rect 30515 969 30593 1015
rect 30639 969 30717 1015
rect 30763 969 30841 1015
rect 30887 969 30965 1015
rect 31011 969 31089 1015
rect 31135 969 31213 1015
rect 31259 969 31337 1015
rect 31383 969 31461 1015
rect 31507 969 31585 1015
rect 31631 969 31709 1015
rect 31755 969 31833 1015
rect 31879 969 31957 1015
rect 32003 969 32081 1015
rect 32127 969 32205 1015
rect 32251 969 32329 1015
rect 32375 969 32453 1015
rect 32499 969 32577 1015
rect 32623 969 32701 1015
rect 32747 969 32825 1015
rect 32871 969 32949 1015
rect 32995 969 33073 1015
rect 33119 969 33197 1015
rect 33243 969 33321 1015
rect 33367 969 33445 1015
rect 33491 969 33569 1015
rect 33615 969 33693 1015
rect 33739 969 33817 1015
rect 33863 969 33941 1015
rect 33987 969 34065 1015
rect 34111 969 34189 1015
rect 34235 969 34313 1015
rect 34359 969 34437 1015
rect 34483 969 34561 1015
rect 34607 969 34685 1015
rect 34731 969 34809 1015
rect 34855 969 34933 1015
rect 34979 969 35057 1015
rect 35103 969 35181 1015
rect 35227 969 35305 1015
rect 35351 969 35429 1015
rect 35475 969 35553 1015
rect 35599 969 35677 1015
rect 35723 969 35801 1015
rect 35847 969 35925 1015
rect 35971 969 36049 1015
rect 36095 969 36173 1015
rect 36219 969 36297 1015
rect 36343 969 36421 1015
rect 36467 969 36545 1015
rect 36591 969 36669 1015
rect 36715 969 36793 1015
rect 36839 969 36917 1015
rect 36963 969 37041 1015
rect 37087 969 37165 1015
rect 37211 969 37289 1015
rect 37335 969 37413 1015
rect 37459 969 37537 1015
rect 37583 969 37661 1015
rect 37707 969 37785 1015
rect 37831 969 37909 1015
rect 37955 969 38033 1015
rect 38079 969 38157 1015
rect 38203 969 38281 1015
rect 38327 969 38405 1015
rect 38451 969 38529 1015
rect 38575 969 38653 1015
rect 38699 969 38777 1015
rect 38823 969 38901 1015
rect 38947 969 39025 1015
rect 39071 969 39149 1015
rect 39195 969 39273 1015
rect 39319 969 39397 1015
rect 39443 969 39521 1015
rect 39567 969 39645 1015
rect 39691 969 39769 1015
rect 39815 969 39893 1015
rect 39939 969 40017 1015
rect 40063 969 40141 1015
rect 40187 969 40265 1015
rect 40311 969 40389 1015
rect 40435 969 40513 1015
rect 40559 969 40637 1015
rect 40683 969 40761 1015
rect 40807 969 40885 1015
rect 40931 969 41009 1015
rect 41055 969 41133 1015
rect 41179 969 41257 1015
rect 41303 969 41381 1015
rect 41427 969 41505 1015
rect 41551 969 41629 1015
rect 41675 969 41753 1015
rect 41799 969 41877 1015
rect 41923 969 42001 1015
rect 42047 969 42125 1015
rect 42171 969 42249 1015
rect 42295 969 42373 1015
rect 42419 969 42497 1015
rect 42543 969 42621 1015
rect 42667 969 42745 1015
rect 42791 969 42869 1015
rect 42915 969 42993 1015
rect 43039 969 43117 1015
rect 43163 969 43241 1015
rect 43287 969 43365 1015
rect 43411 969 43489 1015
rect 43535 969 43613 1015
rect 43659 969 43737 1015
rect 43783 969 43861 1015
rect 43907 969 43985 1015
rect 44031 969 44109 1015
rect 44155 969 44233 1015
rect 44279 969 44357 1015
rect 44403 969 44481 1015
rect 44527 969 44605 1015
rect 44651 969 44729 1015
rect 44775 969 44853 1015
rect 44899 969 44977 1015
rect 45023 969 45101 1015
rect 45147 969 45225 1015
rect 45271 969 45349 1015
rect 45395 969 45473 1015
rect 45519 969 45597 1015
rect 45643 969 45721 1015
rect 45767 969 45845 1015
rect 45891 969 45969 1015
rect 46015 969 46093 1015
rect 46139 969 46217 1015
rect 46263 969 46341 1015
rect 46387 969 46465 1015
rect 46511 969 46589 1015
rect 46635 969 46713 1015
rect 46759 969 46837 1015
rect 46883 969 46961 1015
rect 47007 969 47085 1015
rect 47131 969 47209 1015
rect 47255 969 47333 1015
rect 47379 969 47457 1015
rect 47503 969 47581 1015
rect 47627 969 47705 1015
rect 47751 969 47829 1015
rect 47875 969 47953 1015
rect 47999 969 48077 1015
rect 48123 969 48201 1015
rect 48247 969 48325 1015
rect 48371 969 48449 1015
rect 48495 969 48573 1015
rect 48619 969 48697 1015
rect 48743 969 48821 1015
rect 48867 969 48945 1015
rect 48991 969 49069 1015
rect 49115 969 49193 1015
rect 49239 969 49317 1015
rect 49363 969 49441 1015
rect 49487 969 49565 1015
rect 49611 969 49689 1015
rect 49735 969 49813 1015
rect 49859 969 49937 1015
rect 49983 969 50061 1015
rect 50107 969 50185 1015
rect 50231 969 50309 1015
rect 50355 969 50433 1015
rect 50479 969 50557 1015
rect 50603 969 50681 1015
rect 50727 969 50805 1015
rect 50851 969 50929 1015
rect 50975 969 51053 1015
rect 51099 969 51177 1015
rect 51223 969 51301 1015
rect 51347 969 51425 1015
rect 51471 969 51549 1015
rect 51595 969 51673 1015
rect 51719 969 51797 1015
rect 51843 969 51921 1015
rect 51967 969 52045 1015
rect 52091 969 52169 1015
rect 52215 969 52293 1015
rect 52339 969 52417 1015
rect 52463 969 52541 1015
rect 52587 969 52665 1015
rect 52711 969 52789 1015
rect 52835 969 52913 1015
rect 52959 969 53037 1015
rect 53083 969 53161 1015
rect 53207 969 53285 1015
rect 53331 969 53409 1015
rect 53455 969 53533 1015
rect 53579 969 53657 1015
rect 53703 969 53781 1015
rect 53827 969 53905 1015
rect 53951 969 54029 1015
rect 54075 969 54153 1015
rect 54199 969 54277 1015
rect 54323 969 54401 1015
rect 54447 969 54525 1015
rect 54571 969 54649 1015
rect 54695 969 54773 1015
rect 54819 969 54897 1015
rect 54943 969 55021 1015
rect 55067 969 55145 1015
rect 55191 969 55269 1015
rect 55315 969 55393 1015
rect 55439 969 55517 1015
rect 55563 969 55641 1015
rect 55687 969 55765 1015
rect 55811 969 55889 1015
rect 55935 969 56013 1015
rect 56059 969 56137 1015
rect 56183 969 56261 1015
rect 56307 969 56385 1015
rect 56431 969 56509 1015
rect 56555 969 56633 1015
rect 56679 969 56757 1015
rect 56803 969 56881 1015
rect 56927 969 57005 1015
rect 57051 969 57129 1015
rect 57175 969 57253 1015
rect 57299 969 57377 1015
rect 57423 969 57501 1015
rect 57547 969 57625 1015
rect 57671 969 57749 1015
rect 57795 969 57873 1015
rect 57919 969 57997 1015
rect 58043 969 58121 1015
rect 58167 969 58245 1015
rect 58291 969 58369 1015
rect 58415 969 58493 1015
rect 58539 969 58617 1015
rect 58663 969 58741 1015
rect 58787 969 58865 1015
rect 58911 969 58989 1015
rect 59035 969 59113 1015
rect 59159 969 59237 1015
rect 59283 969 59361 1015
rect 59407 969 59485 1015
rect 59531 969 59609 1015
rect 59655 969 59733 1015
rect 59779 969 59857 1015
rect 59903 969 59981 1015
rect 60027 969 60105 1015
rect 60151 969 60229 1015
rect 60275 969 60353 1015
rect 60399 969 60477 1015
rect 60523 969 60601 1015
rect 60647 969 60725 1015
rect 60771 969 60849 1015
rect 60895 969 60973 1015
rect 61019 969 61097 1015
rect 61143 969 61221 1015
rect 61267 969 61345 1015
rect 61391 969 61469 1015
rect 61515 969 61593 1015
rect 61639 969 61717 1015
rect 61763 969 61841 1015
rect 61887 969 61965 1015
rect 62011 969 62089 1015
rect 62135 969 62213 1015
rect 62259 969 62337 1015
rect 62383 969 62461 1015
rect 62507 969 62585 1015
rect 62631 969 62709 1015
rect 62755 969 62833 1015
rect 62879 969 62957 1015
rect 63003 969 63081 1015
rect 63127 969 63205 1015
rect 63251 969 63329 1015
rect 63375 969 63453 1015
rect 63499 969 63577 1015
rect 63623 969 63701 1015
rect 63747 969 63825 1015
rect 63871 969 63949 1015
rect 63995 969 64073 1015
rect 64119 969 64197 1015
rect 64243 969 64321 1015
rect 64367 969 64445 1015
rect 64491 969 64569 1015
rect 64615 969 64693 1015
rect 64739 969 64817 1015
rect 64863 969 64941 1015
rect 64987 969 65065 1015
rect 65111 969 65189 1015
rect 65235 969 65313 1015
rect 65359 969 65437 1015
rect 65483 969 65561 1015
rect 65607 969 65685 1015
rect 65731 969 65809 1015
rect 65855 969 65933 1015
rect 65979 969 66057 1015
rect 66103 969 66181 1015
rect 66227 969 66305 1015
rect 66351 969 66429 1015
rect 66475 969 66553 1015
rect 66599 969 66677 1015
rect 66723 969 66801 1015
rect 66847 969 66925 1015
rect 66971 969 67049 1015
rect 67095 969 67173 1015
rect 67219 969 67297 1015
rect 67343 969 67421 1015
rect 67467 969 67545 1015
rect 67591 969 67669 1015
rect 67715 969 67793 1015
rect 67839 969 67917 1015
rect 67963 969 68041 1015
rect 68087 969 68165 1015
rect 68211 969 68289 1015
rect 68335 969 68413 1015
rect 68459 969 68537 1015
rect 68583 969 68661 1015
rect 68707 969 68785 1015
rect 68831 969 68909 1015
rect 68955 969 69033 1015
rect 69079 969 69157 1015
rect 69203 969 69281 1015
rect 69327 969 69405 1015
rect 69451 969 69529 1015
rect 69575 969 69653 1015
rect 69699 969 69777 1015
rect 69823 969 69901 1015
rect 69947 969 70025 1015
rect 70071 969 70149 1015
rect 70195 969 70273 1015
rect 70319 969 70397 1015
rect 70443 969 70521 1015
rect 70567 969 70645 1015
rect 70691 969 70769 1015
rect 70815 969 70893 1015
rect 70939 969 71017 1015
rect 71063 969 71141 1015
rect 71187 969 71265 1015
rect 71311 969 71389 1015
rect 71435 969 71513 1015
rect 71559 969 71637 1015
rect 71683 969 71761 1015
rect 71807 969 71885 1015
rect 71931 969 72009 1015
rect 72055 969 72133 1015
rect 72179 969 72257 1015
rect 72303 969 72381 1015
rect 72427 969 72505 1015
rect 72551 969 72629 1015
rect 72675 969 72753 1015
rect 72799 969 72877 1015
rect 72923 969 73001 1015
rect 73047 969 73125 1015
rect 73171 969 73249 1015
rect 73295 969 73373 1015
rect 73419 969 73497 1015
rect 73543 969 73621 1015
rect 73667 969 73745 1015
rect 73791 969 73869 1015
rect 73915 969 73993 1015
rect 74039 969 74117 1015
rect 74163 969 74241 1015
rect 74287 969 74365 1015
rect 74411 969 74489 1015
rect 74535 969 74613 1015
rect 74659 969 74737 1015
rect 74783 969 74861 1015
rect 74907 969 74985 1015
rect 75031 969 75109 1015
rect 75155 969 75233 1015
rect 75279 969 75357 1015
rect 75403 969 75481 1015
rect 75527 969 75605 1015
rect 75651 969 75729 1015
rect 75775 969 75853 1015
rect 75899 969 75977 1015
rect 76023 969 76101 1015
rect 76147 969 76225 1015
rect 76271 969 76349 1015
rect 76395 969 76473 1015
rect 76519 969 76597 1015
rect 76643 969 76721 1015
rect 76767 969 76845 1015
rect 76891 969 76969 1015
rect 77015 969 77093 1015
rect 77139 969 77217 1015
rect 77263 969 77341 1015
rect 77387 969 77465 1015
rect 77511 969 77589 1015
rect 77635 969 77713 1015
rect 77759 969 77837 1015
rect 77883 969 77961 1015
rect 78007 969 78085 1015
rect 78131 969 78209 1015
rect 78255 969 78333 1015
rect 78379 969 78457 1015
rect 78503 969 78581 1015
rect 78627 969 78705 1015
rect 78751 969 78829 1015
rect 78875 969 78953 1015
rect 78999 969 79077 1015
rect 79123 969 79201 1015
rect 79247 969 79325 1015
rect 79371 969 79449 1015
rect 79495 969 79573 1015
rect 79619 969 79697 1015
rect 79743 969 79821 1015
rect 79867 969 79945 1015
rect 79991 969 80069 1015
rect 80115 969 80193 1015
rect 80239 969 80317 1015
rect 80363 969 80441 1015
rect 80487 969 80565 1015
rect 80611 969 80689 1015
rect 80735 969 80813 1015
rect 80859 969 80937 1015
rect 80983 969 81061 1015
rect 81107 969 81185 1015
rect 81231 969 81309 1015
rect 81355 969 81433 1015
rect 81479 969 81557 1015
rect 81603 969 81681 1015
rect 81727 969 81805 1015
rect 81851 969 81929 1015
rect 81975 969 82053 1015
rect 82099 969 82177 1015
rect 82223 969 82301 1015
rect 82347 969 82425 1015
rect 82471 969 82549 1015
rect 82595 969 82673 1015
rect 82719 969 82797 1015
rect 82843 969 82921 1015
rect 82967 969 83045 1015
rect 83091 969 83169 1015
rect 83215 969 83293 1015
rect 83339 969 83417 1015
rect 83463 969 83541 1015
rect 83587 969 83665 1015
rect 83711 969 83789 1015
rect 83835 969 83913 1015
rect 83959 969 84037 1015
rect 84083 969 84161 1015
rect 84207 969 84285 1015
rect 84331 969 84409 1015
rect 84455 969 84533 1015
rect 84579 969 84657 1015
rect 84703 969 84781 1015
rect 84827 969 84905 1015
rect 84951 969 85029 1015
rect 85075 969 85153 1015
rect 85199 969 85277 1015
rect 85323 969 85401 1015
rect 85447 969 85525 1015
rect 85571 969 85649 1015
rect 85695 969 85706 1015
rect 0 891 85706 969
rect 0 845 89 891
rect 135 845 213 891
rect 259 845 337 891
rect 383 845 461 891
rect 507 845 585 891
rect 631 845 709 891
rect 755 845 833 891
rect 879 845 957 891
rect 1003 845 1081 891
rect 1127 845 1205 891
rect 1251 845 1329 891
rect 1375 845 1453 891
rect 1499 845 1577 891
rect 1623 845 1701 891
rect 1747 845 1825 891
rect 1871 845 1949 891
rect 1995 845 2073 891
rect 2119 845 2197 891
rect 2243 845 2321 891
rect 2367 845 2445 891
rect 2491 845 2569 891
rect 2615 845 2693 891
rect 2739 845 2817 891
rect 2863 845 2941 891
rect 2987 845 3065 891
rect 3111 845 3189 891
rect 3235 845 3313 891
rect 3359 845 3437 891
rect 3483 845 3561 891
rect 3607 845 3685 891
rect 3731 845 3809 891
rect 3855 845 3933 891
rect 3979 845 4057 891
rect 4103 845 4181 891
rect 4227 845 4305 891
rect 4351 845 4429 891
rect 4475 845 4553 891
rect 4599 845 4677 891
rect 4723 845 4801 891
rect 4847 845 4925 891
rect 4971 845 5049 891
rect 5095 845 5173 891
rect 5219 845 5297 891
rect 5343 845 5421 891
rect 5467 845 5545 891
rect 5591 845 5669 891
rect 5715 845 5793 891
rect 5839 845 5917 891
rect 5963 845 6041 891
rect 6087 845 6165 891
rect 6211 845 6289 891
rect 6335 845 6413 891
rect 6459 845 6537 891
rect 6583 845 6661 891
rect 6707 845 6785 891
rect 6831 845 6909 891
rect 6955 845 7033 891
rect 7079 845 7157 891
rect 7203 845 7281 891
rect 7327 845 7405 891
rect 7451 845 7529 891
rect 7575 845 7653 891
rect 7699 845 7777 891
rect 7823 845 7901 891
rect 7947 845 8025 891
rect 8071 845 8149 891
rect 8195 845 8273 891
rect 8319 845 8397 891
rect 8443 845 8521 891
rect 8567 845 8645 891
rect 8691 845 8769 891
rect 8815 845 8893 891
rect 8939 845 9017 891
rect 9063 845 9141 891
rect 9187 845 9265 891
rect 9311 845 9389 891
rect 9435 845 9513 891
rect 9559 845 9637 891
rect 9683 845 9761 891
rect 9807 845 9885 891
rect 9931 845 10009 891
rect 10055 845 10133 891
rect 10179 845 10257 891
rect 10303 845 10381 891
rect 10427 845 10505 891
rect 10551 845 10629 891
rect 10675 845 10753 891
rect 10799 845 10877 891
rect 10923 845 11001 891
rect 11047 845 11125 891
rect 11171 845 11249 891
rect 11295 845 11373 891
rect 11419 845 11497 891
rect 11543 845 11621 891
rect 11667 845 11745 891
rect 11791 845 11869 891
rect 11915 845 11993 891
rect 12039 845 12117 891
rect 12163 845 12241 891
rect 12287 845 12365 891
rect 12411 845 12489 891
rect 12535 845 12613 891
rect 12659 845 12737 891
rect 12783 845 12861 891
rect 12907 845 12985 891
rect 13031 845 13109 891
rect 13155 845 13233 891
rect 13279 845 13357 891
rect 13403 845 13481 891
rect 13527 845 13605 891
rect 13651 845 13729 891
rect 13775 845 13853 891
rect 13899 845 13977 891
rect 14023 845 14101 891
rect 14147 845 14225 891
rect 14271 845 14349 891
rect 14395 845 14473 891
rect 14519 845 14597 891
rect 14643 845 14721 891
rect 14767 845 14845 891
rect 14891 845 14969 891
rect 15015 845 15093 891
rect 15139 845 15217 891
rect 15263 845 15341 891
rect 15387 845 15465 891
rect 15511 845 15589 891
rect 15635 845 15713 891
rect 15759 845 15837 891
rect 15883 845 15961 891
rect 16007 845 16085 891
rect 16131 845 16209 891
rect 16255 845 16333 891
rect 16379 845 16457 891
rect 16503 845 16581 891
rect 16627 845 16705 891
rect 16751 845 16829 891
rect 16875 845 16953 891
rect 16999 845 17077 891
rect 17123 845 17201 891
rect 17247 845 17325 891
rect 17371 845 17449 891
rect 17495 845 17573 891
rect 17619 845 17697 891
rect 17743 845 17821 891
rect 17867 845 17945 891
rect 17991 845 18069 891
rect 18115 845 18193 891
rect 18239 845 18317 891
rect 18363 845 18441 891
rect 18487 845 18565 891
rect 18611 845 18689 891
rect 18735 845 18813 891
rect 18859 845 18937 891
rect 18983 845 19061 891
rect 19107 845 19185 891
rect 19231 845 19309 891
rect 19355 845 19433 891
rect 19479 845 19557 891
rect 19603 845 19681 891
rect 19727 845 19805 891
rect 19851 845 19929 891
rect 19975 845 20053 891
rect 20099 845 20177 891
rect 20223 845 20301 891
rect 20347 845 20425 891
rect 20471 845 20549 891
rect 20595 845 20673 891
rect 20719 845 20797 891
rect 20843 845 20921 891
rect 20967 845 21045 891
rect 21091 845 21169 891
rect 21215 845 21293 891
rect 21339 845 21417 891
rect 21463 845 21541 891
rect 21587 845 21665 891
rect 21711 845 21789 891
rect 21835 845 21913 891
rect 21959 845 22037 891
rect 22083 845 22161 891
rect 22207 845 22285 891
rect 22331 845 22409 891
rect 22455 845 22533 891
rect 22579 845 22657 891
rect 22703 845 22781 891
rect 22827 845 22905 891
rect 22951 845 23029 891
rect 23075 845 23153 891
rect 23199 845 23277 891
rect 23323 845 23401 891
rect 23447 845 23525 891
rect 23571 845 23649 891
rect 23695 845 23773 891
rect 23819 845 23897 891
rect 23943 845 24021 891
rect 24067 845 24145 891
rect 24191 845 24269 891
rect 24315 845 24393 891
rect 24439 845 24517 891
rect 24563 845 24641 891
rect 24687 845 24765 891
rect 24811 845 24889 891
rect 24935 845 25013 891
rect 25059 845 25137 891
rect 25183 845 25261 891
rect 25307 845 25385 891
rect 25431 845 25509 891
rect 25555 845 25633 891
rect 25679 845 25757 891
rect 25803 845 25881 891
rect 25927 845 26005 891
rect 26051 845 26129 891
rect 26175 845 26253 891
rect 26299 845 26377 891
rect 26423 845 26501 891
rect 26547 845 26625 891
rect 26671 845 26749 891
rect 26795 845 26873 891
rect 26919 845 26997 891
rect 27043 845 27121 891
rect 27167 845 27245 891
rect 27291 845 27369 891
rect 27415 845 27493 891
rect 27539 845 27617 891
rect 27663 845 27741 891
rect 27787 845 27865 891
rect 27911 845 27989 891
rect 28035 845 28113 891
rect 28159 845 28237 891
rect 28283 845 28361 891
rect 28407 845 28485 891
rect 28531 845 28609 891
rect 28655 845 28733 891
rect 28779 845 28857 891
rect 28903 845 28981 891
rect 29027 845 29105 891
rect 29151 845 29229 891
rect 29275 845 29353 891
rect 29399 845 29477 891
rect 29523 845 29601 891
rect 29647 845 29725 891
rect 29771 845 29849 891
rect 29895 845 29973 891
rect 30019 845 30097 891
rect 30143 845 30221 891
rect 30267 845 30345 891
rect 30391 845 30469 891
rect 30515 845 30593 891
rect 30639 845 30717 891
rect 30763 845 30841 891
rect 30887 845 30965 891
rect 31011 845 31089 891
rect 31135 845 31213 891
rect 31259 845 31337 891
rect 31383 845 31461 891
rect 31507 845 31585 891
rect 31631 845 31709 891
rect 31755 845 31833 891
rect 31879 845 31957 891
rect 32003 845 32081 891
rect 32127 845 32205 891
rect 32251 845 32329 891
rect 32375 845 32453 891
rect 32499 845 32577 891
rect 32623 845 32701 891
rect 32747 845 32825 891
rect 32871 845 32949 891
rect 32995 845 33073 891
rect 33119 845 33197 891
rect 33243 845 33321 891
rect 33367 845 33445 891
rect 33491 845 33569 891
rect 33615 845 33693 891
rect 33739 845 33817 891
rect 33863 845 33941 891
rect 33987 845 34065 891
rect 34111 845 34189 891
rect 34235 845 34313 891
rect 34359 845 34437 891
rect 34483 845 34561 891
rect 34607 845 34685 891
rect 34731 845 34809 891
rect 34855 845 34933 891
rect 34979 845 35057 891
rect 35103 845 35181 891
rect 35227 845 35305 891
rect 35351 845 35429 891
rect 35475 845 35553 891
rect 35599 845 35677 891
rect 35723 845 35801 891
rect 35847 845 35925 891
rect 35971 845 36049 891
rect 36095 845 36173 891
rect 36219 845 36297 891
rect 36343 845 36421 891
rect 36467 845 36545 891
rect 36591 845 36669 891
rect 36715 845 36793 891
rect 36839 845 36917 891
rect 36963 845 37041 891
rect 37087 845 37165 891
rect 37211 845 37289 891
rect 37335 845 37413 891
rect 37459 845 37537 891
rect 37583 845 37661 891
rect 37707 845 37785 891
rect 37831 845 37909 891
rect 37955 845 38033 891
rect 38079 845 38157 891
rect 38203 845 38281 891
rect 38327 845 38405 891
rect 38451 845 38529 891
rect 38575 845 38653 891
rect 38699 845 38777 891
rect 38823 845 38901 891
rect 38947 845 39025 891
rect 39071 845 39149 891
rect 39195 845 39273 891
rect 39319 845 39397 891
rect 39443 845 39521 891
rect 39567 845 39645 891
rect 39691 845 39769 891
rect 39815 845 39893 891
rect 39939 845 40017 891
rect 40063 845 40141 891
rect 40187 845 40265 891
rect 40311 845 40389 891
rect 40435 845 40513 891
rect 40559 845 40637 891
rect 40683 845 40761 891
rect 40807 845 40885 891
rect 40931 845 41009 891
rect 41055 845 41133 891
rect 41179 845 41257 891
rect 41303 845 41381 891
rect 41427 845 41505 891
rect 41551 845 41629 891
rect 41675 845 41753 891
rect 41799 845 41877 891
rect 41923 845 42001 891
rect 42047 845 42125 891
rect 42171 845 42249 891
rect 42295 845 42373 891
rect 42419 845 42497 891
rect 42543 845 42621 891
rect 42667 845 42745 891
rect 42791 845 42869 891
rect 42915 845 42993 891
rect 43039 845 43117 891
rect 43163 845 43241 891
rect 43287 845 43365 891
rect 43411 845 43489 891
rect 43535 845 43613 891
rect 43659 845 43737 891
rect 43783 845 43861 891
rect 43907 845 43985 891
rect 44031 845 44109 891
rect 44155 845 44233 891
rect 44279 845 44357 891
rect 44403 845 44481 891
rect 44527 845 44605 891
rect 44651 845 44729 891
rect 44775 845 44853 891
rect 44899 845 44977 891
rect 45023 845 45101 891
rect 45147 845 45225 891
rect 45271 845 45349 891
rect 45395 845 45473 891
rect 45519 845 45597 891
rect 45643 845 45721 891
rect 45767 845 45845 891
rect 45891 845 45969 891
rect 46015 845 46093 891
rect 46139 845 46217 891
rect 46263 845 46341 891
rect 46387 845 46465 891
rect 46511 845 46589 891
rect 46635 845 46713 891
rect 46759 845 46837 891
rect 46883 845 46961 891
rect 47007 845 47085 891
rect 47131 845 47209 891
rect 47255 845 47333 891
rect 47379 845 47457 891
rect 47503 845 47581 891
rect 47627 845 47705 891
rect 47751 845 47829 891
rect 47875 845 47953 891
rect 47999 845 48077 891
rect 48123 845 48201 891
rect 48247 845 48325 891
rect 48371 845 48449 891
rect 48495 845 48573 891
rect 48619 845 48697 891
rect 48743 845 48821 891
rect 48867 845 48945 891
rect 48991 845 49069 891
rect 49115 845 49193 891
rect 49239 845 49317 891
rect 49363 845 49441 891
rect 49487 845 49565 891
rect 49611 845 49689 891
rect 49735 845 49813 891
rect 49859 845 49937 891
rect 49983 845 50061 891
rect 50107 845 50185 891
rect 50231 845 50309 891
rect 50355 845 50433 891
rect 50479 845 50557 891
rect 50603 845 50681 891
rect 50727 845 50805 891
rect 50851 845 50929 891
rect 50975 845 51053 891
rect 51099 845 51177 891
rect 51223 845 51301 891
rect 51347 845 51425 891
rect 51471 845 51549 891
rect 51595 845 51673 891
rect 51719 845 51797 891
rect 51843 845 51921 891
rect 51967 845 52045 891
rect 52091 845 52169 891
rect 52215 845 52293 891
rect 52339 845 52417 891
rect 52463 845 52541 891
rect 52587 845 52665 891
rect 52711 845 52789 891
rect 52835 845 52913 891
rect 52959 845 53037 891
rect 53083 845 53161 891
rect 53207 845 53285 891
rect 53331 845 53409 891
rect 53455 845 53533 891
rect 53579 845 53657 891
rect 53703 845 53781 891
rect 53827 845 53905 891
rect 53951 845 54029 891
rect 54075 845 54153 891
rect 54199 845 54277 891
rect 54323 845 54401 891
rect 54447 845 54525 891
rect 54571 845 54649 891
rect 54695 845 54773 891
rect 54819 845 54897 891
rect 54943 845 55021 891
rect 55067 845 55145 891
rect 55191 845 55269 891
rect 55315 845 55393 891
rect 55439 845 55517 891
rect 55563 845 55641 891
rect 55687 845 55765 891
rect 55811 845 55889 891
rect 55935 845 56013 891
rect 56059 845 56137 891
rect 56183 845 56261 891
rect 56307 845 56385 891
rect 56431 845 56509 891
rect 56555 845 56633 891
rect 56679 845 56757 891
rect 56803 845 56881 891
rect 56927 845 57005 891
rect 57051 845 57129 891
rect 57175 845 57253 891
rect 57299 845 57377 891
rect 57423 845 57501 891
rect 57547 845 57625 891
rect 57671 845 57749 891
rect 57795 845 57873 891
rect 57919 845 57997 891
rect 58043 845 58121 891
rect 58167 845 58245 891
rect 58291 845 58369 891
rect 58415 845 58493 891
rect 58539 845 58617 891
rect 58663 845 58741 891
rect 58787 845 58865 891
rect 58911 845 58989 891
rect 59035 845 59113 891
rect 59159 845 59237 891
rect 59283 845 59361 891
rect 59407 845 59485 891
rect 59531 845 59609 891
rect 59655 845 59733 891
rect 59779 845 59857 891
rect 59903 845 59981 891
rect 60027 845 60105 891
rect 60151 845 60229 891
rect 60275 845 60353 891
rect 60399 845 60477 891
rect 60523 845 60601 891
rect 60647 845 60725 891
rect 60771 845 60849 891
rect 60895 845 60973 891
rect 61019 845 61097 891
rect 61143 845 61221 891
rect 61267 845 61345 891
rect 61391 845 61469 891
rect 61515 845 61593 891
rect 61639 845 61717 891
rect 61763 845 61841 891
rect 61887 845 61965 891
rect 62011 845 62089 891
rect 62135 845 62213 891
rect 62259 845 62337 891
rect 62383 845 62461 891
rect 62507 845 62585 891
rect 62631 845 62709 891
rect 62755 845 62833 891
rect 62879 845 62957 891
rect 63003 845 63081 891
rect 63127 845 63205 891
rect 63251 845 63329 891
rect 63375 845 63453 891
rect 63499 845 63577 891
rect 63623 845 63701 891
rect 63747 845 63825 891
rect 63871 845 63949 891
rect 63995 845 64073 891
rect 64119 845 64197 891
rect 64243 845 64321 891
rect 64367 845 64445 891
rect 64491 845 64569 891
rect 64615 845 64693 891
rect 64739 845 64817 891
rect 64863 845 64941 891
rect 64987 845 65065 891
rect 65111 845 65189 891
rect 65235 845 65313 891
rect 65359 845 65437 891
rect 65483 845 65561 891
rect 65607 845 65685 891
rect 65731 845 65809 891
rect 65855 845 65933 891
rect 65979 845 66057 891
rect 66103 845 66181 891
rect 66227 845 66305 891
rect 66351 845 66429 891
rect 66475 845 66553 891
rect 66599 845 66677 891
rect 66723 845 66801 891
rect 66847 845 66925 891
rect 66971 845 67049 891
rect 67095 845 67173 891
rect 67219 845 67297 891
rect 67343 845 67421 891
rect 67467 845 67545 891
rect 67591 845 67669 891
rect 67715 845 67793 891
rect 67839 845 67917 891
rect 67963 845 68041 891
rect 68087 845 68165 891
rect 68211 845 68289 891
rect 68335 845 68413 891
rect 68459 845 68537 891
rect 68583 845 68661 891
rect 68707 845 68785 891
rect 68831 845 68909 891
rect 68955 845 69033 891
rect 69079 845 69157 891
rect 69203 845 69281 891
rect 69327 845 69405 891
rect 69451 845 69529 891
rect 69575 845 69653 891
rect 69699 845 69777 891
rect 69823 845 69901 891
rect 69947 845 70025 891
rect 70071 845 70149 891
rect 70195 845 70273 891
rect 70319 845 70397 891
rect 70443 845 70521 891
rect 70567 845 70645 891
rect 70691 845 70769 891
rect 70815 845 70893 891
rect 70939 845 71017 891
rect 71063 845 71141 891
rect 71187 845 71265 891
rect 71311 845 71389 891
rect 71435 845 71513 891
rect 71559 845 71637 891
rect 71683 845 71761 891
rect 71807 845 71885 891
rect 71931 845 72009 891
rect 72055 845 72133 891
rect 72179 845 72257 891
rect 72303 845 72381 891
rect 72427 845 72505 891
rect 72551 845 72629 891
rect 72675 845 72753 891
rect 72799 845 72877 891
rect 72923 845 73001 891
rect 73047 845 73125 891
rect 73171 845 73249 891
rect 73295 845 73373 891
rect 73419 845 73497 891
rect 73543 845 73621 891
rect 73667 845 73745 891
rect 73791 845 73869 891
rect 73915 845 73993 891
rect 74039 845 74117 891
rect 74163 845 74241 891
rect 74287 845 74365 891
rect 74411 845 74489 891
rect 74535 845 74613 891
rect 74659 845 74737 891
rect 74783 845 74861 891
rect 74907 845 74985 891
rect 75031 845 75109 891
rect 75155 845 75233 891
rect 75279 845 75357 891
rect 75403 845 75481 891
rect 75527 845 75605 891
rect 75651 845 75729 891
rect 75775 845 75853 891
rect 75899 845 75977 891
rect 76023 845 76101 891
rect 76147 845 76225 891
rect 76271 845 76349 891
rect 76395 845 76473 891
rect 76519 845 76597 891
rect 76643 845 76721 891
rect 76767 845 76845 891
rect 76891 845 76969 891
rect 77015 845 77093 891
rect 77139 845 77217 891
rect 77263 845 77341 891
rect 77387 845 77465 891
rect 77511 845 77589 891
rect 77635 845 77713 891
rect 77759 845 77837 891
rect 77883 845 77961 891
rect 78007 845 78085 891
rect 78131 845 78209 891
rect 78255 845 78333 891
rect 78379 845 78457 891
rect 78503 845 78581 891
rect 78627 845 78705 891
rect 78751 845 78829 891
rect 78875 845 78953 891
rect 78999 845 79077 891
rect 79123 845 79201 891
rect 79247 845 79325 891
rect 79371 845 79449 891
rect 79495 845 79573 891
rect 79619 845 79697 891
rect 79743 845 79821 891
rect 79867 845 79945 891
rect 79991 845 80069 891
rect 80115 845 80193 891
rect 80239 845 80317 891
rect 80363 845 80441 891
rect 80487 845 80565 891
rect 80611 845 80689 891
rect 80735 845 80813 891
rect 80859 845 80937 891
rect 80983 845 81061 891
rect 81107 845 81185 891
rect 81231 845 81309 891
rect 81355 845 81433 891
rect 81479 845 81557 891
rect 81603 845 81681 891
rect 81727 845 81805 891
rect 81851 845 81929 891
rect 81975 845 82053 891
rect 82099 845 82177 891
rect 82223 845 82301 891
rect 82347 845 82425 891
rect 82471 845 82549 891
rect 82595 845 82673 891
rect 82719 845 82797 891
rect 82843 845 82921 891
rect 82967 845 83045 891
rect 83091 845 83169 891
rect 83215 845 83293 891
rect 83339 845 83417 891
rect 83463 845 83541 891
rect 83587 845 83665 891
rect 83711 845 83789 891
rect 83835 845 83913 891
rect 83959 845 84037 891
rect 84083 845 84161 891
rect 84207 845 84285 891
rect 84331 845 84409 891
rect 84455 845 84533 891
rect 84579 845 84657 891
rect 84703 845 84781 891
rect 84827 845 84905 891
rect 84951 845 85029 891
rect 85075 845 85153 891
rect 85199 845 85277 891
rect 85323 845 85401 891
rect 85447 845 85525 891
rect 85571 845 85649 891
rect 85695 845 85706 891
rect 0 767 85706 845
rect 0 721 89 767
rect 135 721 213 767
rect 259 721 337 767
rect 383 721 461 767
rect 507 721 585 767
rect 631 721 709 767
rect 755 721 833 767
rect 879 721 957 767
rect 1003 721 1081 767
rect 1127 721 1205 767
rect 1251 721 1329 767
rect 1375 721 1453 767
rect 1499 721 1577 767
rect 1623 721 1701 767
rect 1747 721 1825 767
rect 1871 721 1949 767
rect 1995 721 2073 767
rect 2119 721 2197 767
rect 2243 721 2321 767
rect 2367 721 2445 767
rect 2491 721 2569 767
rect 2615 721 2693 767
rect 2739 721 2817 767
rect 2863 721 2941 767
rect 2987 721 3065 767
rect 3111 721 3189 767
rect 3235 721 3313 767
rect 3359 721 3437 767
rect 3483 721 3561 767
rect 3607 721 3685 767
rect 3731 721 3809 767
rect 3855 721 3933 767
rect 3979 721 4057 767
rect 4103 721 4181 767
rect 4227 721 4305 767
rect 4351 721 4429 767
rect 4475 721 4553 767
rect 4599 721 4677 767
rect 4723 721 4801 767
rect 4847 721 4925 767
rect 4971 721 5049 767
rect 5095 721 5173 767
rect 5219 721 5297 767
rect 5343 721 5421 767
rect 5467 721 5545 767
rect 5591 721 5669 767
rect 5715 721 5793 767
rect 5839 721 5917 767
rect 5963 721 6041 767
rect 6087 721 6165 767
rect 6211 721 6289 767
rect 6335 721 6413 767
rect 6459 721 6537 767
rect 6583 721 6661 767
rect 6707 721 6785 767
rect 6831 721 6909 767
rect 6955 721 7033 767
rect 7079 721 7157 767
rect 7203 721 7281 767
rect 7327 721 7405 767
rect 7451 721 7529 767
rect 7575 721 7653 767
rect 7699 721 7777 767
rect 7823 721 7901 767
rect 7947 721 8025 767
rect 8071 721 8149 767
rect 8195 721 8273 767
rect 8319 721 8397 767
rect 8443 721 8521 767
rect 8567 721 8645 767
rect 8691 721 8769 767
rect 8815 721 8893 767
rect 8939 721 9017 767
rect 9063 721 9141 767
rect 9187 721 9265 767
rect 9311 721 9389 767
rect 9435 721 9513 767
rect 9559 721 9637 767
rect 9683 721 9761 767
rect 9807 721 9885 767
rect 9931 721 10009 767
rect 10055 721 10133 767
rect 10179 721 10257 767
rect 10303 721 10381 767
rect 10427 721 10505 767
rect 10551 721 10629 767
rect 10675 721 10753 767
rect 10799 721 10877 767
rect 10923 721 11001 767
rect 11047 721 11125 767
rect 11171 721 11249 767
rect 11295 721 11373 767
rect 11419 721 11497 767
rect 11543 721 11621 767
rect 11667 721 11745 767
rect 11791 721 11869 767
rect 11915 721 11993 767
rect 12039 721 12117 767
rect 12163 721 12241 767
rect 12287 721 12365 767
rect 12411 721 12489 767
rect 12535 721 12613 767
rect 12659 721 12737 767
rect 12783 721 12861 767
rect 12907 721 12985 767
rect 13031 721 13109 767
rect 13155 721 13233 767
rect 13279 721 13357 767
rect 13403 721 13481 767
rect 13527 721 13605 767
rect 13651 721 13729 767
rect 13775 721 13853 767
rect 13899 721 13977 767
rect 14023 721 14101 767
rect 14147 721 14225 767
rect 14271 721 14349 767
rect 14395 721 14473 767
rect 14519 721 14597 767
rect 14643 721 14721 767
rect 14767 721 14845 767
rect 14891 721 14969 767
rect 15015 721 15093 767
rect 15139 721 15217 767
rect 15263 721 15341 767
rect 15387 721 15465 767
rect 15511 721 15589 767
rect 15635 721 15713 767
rect 15759 721 15837 767
rect 15883 721 15961 767
rect 16007 721 16085 767
rect 16131 721 16209 767
rect 16255 721 16333 767
rect 16379 721 16457 767
rect 16503 721 16581 767
rect 16627 721 16705 767
rect 16751 721 16829 767
rect 16875 721 16953 767
rect 16999 721 17077 767
rect 17123 721 17201 767
rect 17247 721 17325 767
rect 17371 721 17449 767
rect 17495 721 17573 767
rect 17619 721 17697 767
rect 17743 721 17821 767
rect 17867 721 17945 767
rect 17991 721 18069 767
rect 18115 721 18193 767
rect 18239 721 18317 767
rect 18363 721 18441 767
rect 18487 721 18565 767
rect 18611 721 18689 767
rect 18735 721 18813 767
rect 18859 721 18937 767
rect 18983 721 19061 767
rect 19107 721 19185 767
rect 19231 721 19309 767
rect 19355 721 19433 767
rect 19479 721 19557 767
rect 19603 721 19681 767
rect 19727 721 19805 767
rect 19851 721 19929 767
rect 19975 721 20053 767
rect 20099 721 20177 767
rect 20223 721 20301 767
rect 20347 721 20425 767
rect 20471 721 20549 767
rect 20595 721 20673 767
rect 20719 721 20797 767
rect 20843 721 20921 767
rect 20967 721 21045 767
rect 21091 721 21169 767
rect 21215 721 21293 767
rect 21339 721 21417 767
rect 21463 721 21541 767
rect 21587 721 21665 767
rect 21711 721 21789 767
rect 21835 721 21913 767
rect 21959 721 22037 767
rect 22083 721 22161 767
rect 22207 721 22285 767
rect 22331 721 22409 767
rect 22455 721 22533 767
rect 22579 721 22657 767
rect 22703 721 22781 767
rect 22827 721 22905 767
rect 22951 721 23029 767
rect 23075 721 23153 767
rect 23199 721 23277 767
rect 23323 721 23401 767
rect 23447 721 23525 767
rect 23571 721 23649 767
rect 23695 721 23773 767
rect 23819 721 23897 767
rect 23943 721 24021 767
rect 24067 721 24145 767
rect 24191 721 24269 767
rect 24315 721 24393 767
rect 24439 721 24517 767
rect 24563 721 24641 767
rect 24687 721 24765 767
rect 24811 721 24889 767
rect 24935 721 25013 767
rect 25059 721 25137 767
rect 25183 721 25261 767
rect 25307 721 25385 767
rect 25431 721 25509 767
rect 25555 721 25633 767
rect 25679 721 25757 767
rect 25803 721 25881 767
rect 25927 721 26005 767
rect 26051 721 26129 767
rect 26175 721 26253 767
rect 26299 721 26377 767
rect 26423 721 26501 767
rect 26547 721 26625 767
rect 26671 721 26749 767
rect 26795 721 26873 767
rect 26919 721 26997 767
rect 27043 721 27121 767
rect 27167 721 27245 767
rect 27291 721 27369 767
rect 27415 721 27493 767
rect 27539 721 27617 767
rect 27663 721 27741 767
rect 27787 721 27865 767
rect 27911 721 27989 767
rect 28035 721 28113 767
rect 28159 721 28237 767
rect 28283 721 28361 767
rect 28407 721 28485 767
rect 28531 721 28609 767
rect 28655 721 28733 767
rect 28779 721 28857 767
rect 28903 721 28981 767
rect 29027 721 29105 767
rect 29151 721 29229 767
rect 29275 721 29353 767
rect 29399 721 29477 767
rect 29523 721 29601 767
rect 29647 721 29725 767
rect 29771 721 29849 767
rect 29895 721 29973 767
rect 30019 721 30097 767
rect 30143 721 30221 767
rect 30267 721 30345 767
rect 30391 721 30469 767
rect 30515 721 30593 767
rect 30639 721 30717 767
rect 30763 721 30841 767
rect 30887 721 30965 767
rect 31011 721 31089 767
rect 31135 721 31213 767
rect 31259 721 31337 767
rect 31383 721 31461 767
rect 31507 721 31585 767
rect 31631 721 31709 767
rect 31755 721 31833 767
rect 31879 721 31957 767
rect 32003 721 32081 767
rect 32127 721 32205 767
rect 32251 721 32329 767
rect 32375 721 32453 767
rect 32499 721 32577 767
rect 32623 721 32701 767
rect 32747 721 32825 767
rect 32871 721 32949 767
rect 32995 721 33073 767
rect 33119 721 33197 767
rect 33243 721 33321 767
rect 33367 721 33445 767
rect 33491 721 33569 767
rect 33615 721 33693 767
rect 33739 721 33817 767
rect 33863 721 33941 767
rect 33987 721 34065 767
rect 34111 721 34189 767
rect 34235 721 34313 767
rect 34359 721 34437 767
rect 34483 721 34561 767
rect 34607 721 34685 767
rect 34731 721 34809 767
rect 34855 721 34933 767
rect 34979 721 35057 767
rect 35103 721 35181 767
rect 35227 721 35305 767
rect 35351 721 35429 767
rect 35475 721 35553 767
rect 35599 721 35677 767
rect 35723 721 35801 767
rect 35847 721 35925 767
rect 35971 721 36049 767
rect 36095 721 36173 767
rect 36219 721 36297 767
rect 36343 721 36421 767
rect 36467 721 36545 767
rect 36591 721 36669 767
rect 36715 721 36793 767
rect 36839 721 36917 767
rect 36963 721 37041 767
rect 37087 721 37165 767
rect 37211 721 37289 767
rect 37335 721 37413 767
rect 37459 721 37537 767
rect 37583 721 37661 767
rect 37707 721 37785 767
rect 37831 721 37909 767
rect 37955 721 38033 767
rect 38079 721 38157 767
rect 38203 721 38281 767
rect 38327 721 38405 767
rect 38451 721 38529 767
rect 38575 721 38653 767
rect 38699 721 38777 767
rect 38823 721 38901 767
rect 38947 721 39025 767
rect 39071 721 39149 767
rect 39195 721 39273 767
rect 39319 721 39397 767
rect 39443 721 39521 767
rect 39567 721 39645 767
rect 39691 721 39769 767
rect 39815 721 39893 767
rect 39939 721 40017 767
rect 40063 721 40141 767
rect 40187 721 40265 767
rect 40311 721 40389 767
rect 40435 721 40513 767
rect 40559 721 40637 767
rect 40683 721 40761 767
rect 40807 721 40885 767
rect 40931 721 41009 767
rect 41055 721 41133 767
rect 41179 721 41257 767
rect 41303 721 41381 767
rect 41427 721 41505 767
rect 41551 721 41629 767
rect 41675 721 41753 767
rect 41799 721 41877 767
rect 41923 721 42001 767
rect 42047 721 42125 767
rect 42171 721 42249 767
rect 42295 721 42373 767
rect 42419 721 42497 767
rect 42543 721 42621 767
rect 42667 721 42745 767
rect 42791 721 42869 767
rect 42915 721 42993 767
rect 43039 721 43117 767
rect 43163 721 43241 767
rect 43287 721 43365 767
rect 43411 721 43489 767
rect 43535 721 43613 767
rect 43659 721 43737 767
rect 43783 721 43861 767
rect 43907 721 43985 767
rect 44031 721 44109 767
rect 44155 721 44233 767
rect 44279 721 44357 767
rect 44403 721 44481 767
rect 44527 721 44605 767
rect 44651 721 44729 767
rect 44775 721 44853 767
rect 44899 721 44977 767
rect 45023 721 45101 767
rect 45147 721 45225 767
rect 45271 721 45349 767
rect 45395 721 45473 767
rect 45519 721 45597 767
rect 45643 721 45721 767
rect 45767 721 45845 767
rect 45891 721 45969 767
rect 46015 721 46093 767
rect 46139 721 46217 767
rect 46263 721 46341 767
rect 46387 721 46465 767
rect 46511 721 46589 767
rect 46635 721 46713 767
rect 46759 721 46837 767
rect 46883 721 46961 767
rect 47007 721 47085 767
rect 47131 721 47209 767
rect 47255 721 47333 767
rect 47379 721 47457 767
rect 47503 721 47581 767
rect 47627 721 47705 767
rect 47751 721 47829 767
rect 47875 721 47953 767
rect 47999 721 48077 767
rect 48123 721 48201 767
rect 48247 721 48325 767
rect 48371 721 48449 767
rect 48495 721 48573 767
rect 48619 721 48697 767
rect 48743 721 48821 767
rect 48867 721 48945 767
rect 48991 721 49069 767
rect 49115 721 49193 767
rect 49239 721 49317 767
rect 49363 721 49441 767
rect 49487 721 49565 767
rect 49611 721 49689 767
rect 49735 721 49813 767
rect 49859 721 49937 767
rect 49983 721 50061 767
rect 50107 721 50185 767
rect 50231 721 50309 767
rect 50355 721 50433 767
rect 50479 721 50557 767
rect 50603 721 50681 767
rect 50727 721 50805 767
rect 50851 721 50929 767
rect 50975 721 51053 767
rect 51099 721 51177 767
rect 51223 721 51301 767
rect 51347 721 51425 767
rect 51471 721 51549 767
rect 51595 721 51673 767
rect 51719 721 51797 767
rect 51843 721 51921 767
rect 51967 721 52045 767
rect 52091 721 52169 767
rect 52215 721 52293 767
rect 52339 721 52417 767
rect 52463 721 52541 767
rect 52587 721 52665 767
rect 52711 721 52789 767
rect 52835 721 52913 767
rect 52959 721 53037 767
rect 53083 721 53161 767
rect 53207 721 53285 767
rect 53331 721 53409 767
rect 53455 721 53533 767
rect 53579 721 53657 767
rect 53703 721 53781 767
rect 53827 721 53905 767
rect 53951 721 54029 767
rect 54075 721 54153 767
rect 54199 721 54277 767
rect 54323 721 54401 767
rect 54447 721 54525 767
rect 54571 721 54649 767
rect 54695 721 54773 767
rect 54819 721 54897 767
rect 54943 721 55021 767
rect 55067 721 55145 767
rect 55191 721 55269 767
rect 55315 721 55393 767
rect 55439 721 55517 767
rect 55563 721 55641 767
rect 55687 721 55765 767
rect 55811 721 55889 767
rect 55935 721 56013 767
rect 56059 721 56137 767
rect 56183 721 56261 767
rect 56307 721 56385 767
rect 56431 721 56509 767
rect 56555 721 56633 767
rect 56679 721 56757 767
rect 56803 721 56881 767
rect 56927 721 57005 767
rect 57051 721 57129 767
rect 57175 721 57253 767
rect 57299 721 57377 767
rect 57423 721 57501 767
rect 57547 721 57625 767
rect 57671 721 57749 767
rect 57795 721 57873 767
rect 57919 721 57997 767
rect 58043 721 58121 767
rect 58167 721 58245 767
rect 58291 721 58369 767
rect 58415 721 58493 767
rect 58539 721 58617 767
rect 58663 721 58741 767
rect 58787 721 58865 767
rect 58911 721 58989 767
rect 59035 721 59113 767
rect 59159 721 59237 767
rect 59283 721 59361 767
rect 59407 721 59485 767
rect 59531 721 59609 767
rect 59655 721 59733 767
rect 59779 721 59857 767
rect 59903 721 59981 767
rect 60027 721 60105 767
rect 60151 721 60229 767
rect 60275 721 60353 767
rect 60399 721 60477 767
rect 60523 721 60601 767
rect 60647 721 60725 767
rect 60771 721 60849 767
rect 60895 721 60973 767
rect 61019 721 61097 767
rect 61143 721 61221 767
rect 61267 721 61345 767
rect 61391 721 61469 767
rect 61515 721 61593 767
rect 61639 721 61717 767
rect 61763 721 61841 767
rect 61887 721 61965 767
rect 62011 721 62089 767
rect 62135 721 62213 767
rect 62259 721 62337 767
rect 62383 721 62461 767
rect 62507 721 62585 767
rect 62631 721 62709 767
rect 62755 721 62833 767
rect 62879 721 62957 767
rect 63003 721 63081 767
rect 63127 721 63205 767
rect 63251 721 63329 767
rect 63375 721 63453 767
rect 63499 721 63577 767
rect 63623 721 63701 767
rect 63747 721 63825 767
rect 63871 721 63949 767
rect 63995 721 64073 767
rect 64119 721 64197 767
rect 64243 721 64321 767
rect 64367 721 64445 767
rect 64491 721 64569 767
rect 64615 721 64693 767
rect 64739 721 64817 767
rect 64863 721 64941 767
rect 64987 721 65065 767
rect 65111 721 65189 767
rect 65235 721 65313 767
rect 65359 721 65437 767
rect 65483 721 65561 767
rect 65607 721 65685 767
rect 65731 721 65809 767
rect 65855 721 65933 767
rect 65979 721 66057 767
rect 66103 721 66181 767
rect 66227 721 66305 767
rect 66351 721 66429 767
rect 66475 721 66553 767
rect 66599 721 66677 767
rect 66723 721 66801 767
rect 66847 721 66925 767
rect 66971 721 67049 767
rect 67095 721 67173 767
rect 67219 721 67297 767
rect 67343 721 67421 767
rect 67467 721 67545 767
rect 67591 721 67669 767
rect 67715 721 67793 767
rect 67839 721 67917 767
rect 67963 721 68041 767
rect 68087 721 68165 767
rect 68211 721 68289 767
rect 68335 721 68413 767
rect 68459 721 68537 767
rect 68583 721 68661 767
rect 68707 721 68785 767
rect 68831 721 68909 767
rect 68955 721 69033 767
rect 69079 721 69157 767
rect 69203 721 69281 767
rect 69327 721 69405 767
rect 69451 721 69529 767
rect 69575 721 69653 767
rect 69699 721 69777 767
rect 69823 721 69901 767
rect 69947 721 70025 767
rect 70071 721 70149 767
rect 70195 721 70273 767
rect 70319 721 70397 767
rect 70443 721 70521 767
rect 70567 721 70645 767
rect 70691 721 70769 767
rect 70815 721 70893 767
rect 70939 721 71017 767
rect 71063 721 71141 767
rect 71187 721 71265 767
rect 71311 721 71389 767
rect 71435 721 71513 767
rect 71559 721 71637 767
rect 71683 721 71761 767
rect 71807 721 71885 767
rect 71931 721 72009 767
rect 72055 721 72133 767
rect 72179 721 72257 767
rect 72303 721 72381 767
rect 72427 721 72505 767
rect 72551 721 72629 767
rect 72675 721 72753 767
rect 72799 721 72877 767
rect 72923 721 73001 767
rect 73047 721 73125 767
rect 73171 721 73249 767
rect 73295 721 73373 767
rect 73419 721 73497 767
rect 73543 721 73621 767
rect 73667 721 73745 767
rect 73791 721 73869 767
rect 73915 721 73993 767
rect 74039 721 74117 767
rect 74163 721 74241 767
rect 74287 721 74365 767
rect 74411 721 74489 767
rect 74535 721 74613 767
rect 74659 721 74737 767
rect 74783 721 74861 767
rect 74907 721 74985 767
rect 75031 721 75109 767
rect 75155 721 75233 767
rect 75279 721 75357 767
rect 75403 721 75481 767
rect 75527 721 75605 767
rect 75651 721 75729 767
rect 75775 721 75853 767
rect 75899 721 75977 767
rect 76023 721 76101 767
rect 76147 721 76225 767
rect 76271 721 76349 767
rect 76395 721 76473 767
rect 76519 721 76597 767
rect 76643 721 76721 767
rect 76767 721 76845 767
rect 76891 721 76969 767
rect 77015 721 77093 767
rect 77139 721 77217 767
rect 77263 721 77341 767
rect 77387 721 77465 767
rect 77511 721 77589 767
rect 77635 721 77713 767
rect 77759 721 77837 767
rect 77883 721 77961 767
rect 78007 721 78085 767
rect 78131 721 78209 767
rect 78255 721 78333 767
rect 78379 721 78457 767
rect 78503 721 78581 767
rect 78627 721 78705 767
rect 78751 721 78829 767
rect 78875 721 78953 767
rect 78999 721 79077 767
rect 79123 721 79201 767
rect 79247 721 79325 767
rect 79371 721 79449 767
rect 79495 721 79573 767
rect 79619 721 79697 767
rect 79743 721 79821 767
rect 79867 721 79945 767
rect 79991 721 80069 767
rect 80115 721 80193 767
rect 80239 721 80317 767
rect 80363 721 80441 767
rect 80487 721 80565 767
rect 80611 721 80689 767
rect 80735 721 80813 767
rect 80859 721 80937 767
rect 80983 721 81061 767
rect 81107 721 81185 767
rect 81231 721 81309 767
rect 81355 721 81433 767
rect 81479 721 81557 767
rect 81603 721 81681 767
rect 81727 721 81805 767
rect 81851 721 81929 767
rect 81975 721 82053 767
rect 82099 721 82177 767
rect 82223 721 82301 767
rect 82347 721 82425 767
rect 82471 721 82549 767
rect 82595 721 82673 767
rect 82719 721 82797 767
rect 82843 721 82921 767
rect 82967 721 83045 767
rect 83091 721 83169 767
rect 83215 721 83293 767
rect 83339 721 83417 767
rect 83463 721 83541 767
rect 83587 721 83665 767
rect 83711 721 83789 767
rect 83835 721 83913 767
rect 83959 721 84037 767
rect 84083 721 84161 767
rect 84207 721 84285 767
rect 84331 721 84409 767
rect 84455 721 84533 767
rect 84579 721 84657 767
rect 84703 721 84781 767
rect 84827 721 84905 767
rect 84951 721 85029 767
rect 85075 721 85153 767
rect 85199 721 85277 767
rect 85323 721 85401 767
rect 85447 721 85525 767
rect 85571 721 85649 767
rect 85695 721 85706 767
rect 0 643 85706 721
rect 0 597 89 643
rect 135 597 213 643
rect 259 597 337 643
rect 383 597 461 643
rect 507 597 585 643
rect 631 597 709 643
rect 755 597 833 643
rect 879 597 957 643
rect 1003 597 1081 643
rect 1127 597 1205 643
rect 1251 597 1329 643
rect 1375 597 1453 643
rect 1499 597 1577 643
rect 1623 597 1701 643
rect 1747 597 1825 643
rect 1871 597 1949 643
rect 1995 597 2073 643
rect 2119 597 2197 643
rect 2243 597 2321 643
rect 2367 597 2445 643
rect 2491 597 2569 643
rect 2615 597 2693 643
rect 2739 597 2817 643
rect 2863 597 2941 643
rect 2987 597 3065 643
rect 3111 597 3189 643
rect 3235 597 3313 643
rect 3359 597 3437 643
rect 3483 597 3561 643
rect 3607 597 3685 643
rect 3731 597 3809 643
rect 3855 597 3933 643
rect 3979 597 4057 643
rect 4103 597 4181 643
rect 4227 597 4305 643
rect 4351 597 4429 643
rect 4475 597 4553 643
rect 4599 597 4677 643
rect 4723 597 4801 643
rect 4847 597 4925 643
rect 4971 597 5049 643
rect 5095 597 5173 643
rect 5219 597 5297 643
rect 5343 597 5421 643
rect 5467 597 5545 643
rect 5591 597 5669 643
rect 5715 597 5793 643
rect 5839 597 5917 643
rect 5963 597 6041 643
rect 6087 597 6165 643
rect 6211 597 6289 643
rect 6335 597 6413 643
rect 6459 597 6537 643
rect 6583 597 6661 643
rect 6707 597 6785 643
rect 6831 597 6909 643
rect 6955 597 7033 643
rect 7079 597 7157 643
rect 7203 597 7281 643
rect 7327 597 7405 643
rect 7451 597 7529 643
rect 7575 597 7653 643
rect 7699 597 7777 643
rect 7823 597 7901 643
rect 7947 597 8025 643
rect 8071 597 8149 643
rect 8195 597 8273 643
rect 8319 597 8397 643
rect 8443 597 8521 643
rect 8567 597 8645 643
rect 8691 597 8769 643
rect 8815 597 8893 643
rect 8939 597 9017 643
rect 9063 597 9141 643
rect 9187 597 9265 643
rect 9311 597 9389 643
rect 9435 597 9513 643
rect 9559 597 9637 643
rect 9683 597 9761 643
rect 9807 597 9885 643
rect 9931 597 10009 643
rect 10055 597 10133 643
rect 10179 597 10257 643
rect 10303 597 10381 643
rect 10427 597 10505 643
rect 10551 597 10629 643
rect 10675 597 10753 643
rect 10799 597 10877 643
rect 10923 597 11001 643
rect 11047 597 11125 643
rect 11171 597 11249 643
rect 11295 597 11373 643
rect 11419 597 11497 643
rect 11543 597 11621 643
rect 11667 597 11745 643
rect 11791 597 11869 643
rect 11915 597 11993 643
rect 12039 597 12117 643
rect 12163 597 12241 643
rect 12287 597 12365 643
rect 12411 597 12489 643
rect 12535 597 12613 643
rect 12659 597 12737 643
rect 12783 597 12861 643
rect 12907 597 12985 643
rect 13031 597 13109 643
rect 13155 597 13233 643
rect 13279 597 13357 643
rect 13403 597 13481 643
rect 13527 597 13605 643
rect 13651 597 13729 643
rect 13775 597 13853 643
rect 13899 597 13977 643
rect 14023 597 14101 643
rect 14147 597 14225 643
rect 14271 597 14349 643
rect 14395 597 14473 643
rect 14519 597 14597 643
rect 14643 597 14721 643
rect 14767 597 14845 643
rect 14891 597 14969 643
rect 15015 597 15093 643
rect 15139 597 15217 643
rect 15263 597 15341 643
rect 15387 597 15465 643
rect 15511 597 15589 643
rect 15635 597 15713 643
rect 15759 597 15837 643
rect 15883 597 15961 643
rect 16007 597 16085 643
rect 16131 597 16209 643
rect 16255 597 16333 643
rect 16379 597 16457 643
rect 16503 597 16581 643
rect 16627 597 16705 643
rect 16751 597 16829 643
rect 16875 597 16953 643
rect 16999 597 17077 643
rect 17123 597 17201 643
rect 17247 597 17325 643
rect 17371 597 17449 643
rect 17495 597 17573 643
rect 17619 597 17697 643
rect 17743 597 17821 643
rect 17867 597 17945 643
rect 17991 597 18069 643
rect 18115 597 18193 643
rect 18239 597 18317 643
rect 18363 597 18441 643
rect 18487 597 18565 643
rect 18611 597 18689 643
rect 18735 597 18813 643
rect 18859 597 18937 643
rect 18983 597 19061 643
rect 19107 597 19185 643
rect 19231 597 19309 643
rect 19355 597 19433 643
rect 19479 597 19557 643
rect 19603 597 19681 643
rect 19727 597 19805 643
rect 19851 597 19929 643
rect 19975 597 20053 643
rect 20099 597 20177 643
rect 20223 597 20301 643
rect 20347 597 20425 643
rect 20471 597 20549 643
rect 20595 597 20673 643
rect 20719 597 20797 643
rect 20843 597 20921 643
rect 20967 597 21045 643
rect 21091 597 21169 643
rect 21215 597 21293 643
rect 21339 597 21417 643
rect 21463 597 21541 643
rect 21587 597 21665 643
rect 21711 597 21789 643
rect 21835 597 21913 643
rect 21959 597 22037 643
rect 22083 597 22161 643
rect 22207 597 22285 643
rect 22331 597 22409 643
rect 22455 597 22533 643
rect 22579 597 22657 643
rect 22703 597 22781 643
rect 22827 597 22905 643
rect 22951 597 23029 643
rect 23075 597 23153 643
rect 23199 597 23277 643
rect 23323 597 23401 643
rect 23447 597 23525 643
rect 23571 597 23649 643
rect 23695 597 23773 643
rect 23819 597 23897 643
rect 23943 597 24021 643
rect 24067 597 24145 643
rect 24191 597 24269 643
rect 24315 597 24393 643
rect 24439 597 24517 643
rect 24563 597 24641 643
rect 24687 597 24765 643
rect 24811 597 24889 643
rect 24935 597 25013 643
rect 25059 597 25137 643
rect 25183 597 25261 643
rect 25307 597 25385 643
rect 25431 597 25509 643
rect 25555 597 25633 643
rect 25679 597 25757 643
rect 25803 597 25881 643
rect 25927 597 26005 643
rect 26051 597 26129 643
rect 26175 597 26253 643
rect 26299 597 26377 643
rect 26423 597 26501 643
rect 26547 597 26625 643
rect 26671 597 26749 643
rect 26795 597 26873 643
rect 26919 597 26997 643
rect 27043 597 27121 643
rect 27167 597 27245 643
rect 27291 597 27369 643
rect 27415 597 27493 643
rect 27539 597 27617 643
rect 27663 597 27741 643
rect 27787 597 27865 643
rect 27911 597 27989 643
rect 28035 597 28113 643
rect 28159 597 28237 643
rect 28283 597 28361 643
rect 28407 597 28485 643
rect 28531 597 28609 643
rect 28655 597 28733 643
rect 28779 597 28857 643
rect 28903 597 28981 643
rect 29027 597 29105 643
rect 29151 597 29229 643
rect 29275 597 29353 643
rect 29399 597 29477 643
rect 29523 597 29601 643
rect 29647 597 29725 643
rect 29771 597 29849 643
rect 29895 597 29973 643
rect 30019 597 30097 643
rect 30143 597 30221 643
rect 30267 597 30345 643
rect 30391 597 30469 643
rect 30515 597 30593 643
rect 30639 597 30717 643
rect 30763 597 30841 643
rect 30887 597 30965 643
rect 31011 597 31089 643
rect 31135 597 31213 643
rect 31259 597 31337 643
rect 31383 597 31461 643
rect 31507 597 31585 643
rect 31631 597 31709 643
rect 31755 597 31833 643
rect 31879 597 31957 643
rect 32003 597 32081 643
rect 32127 597 32205 643
rect 32251 597 32329 643
rect 32375 597 32453 643
rect 32499 597 32577 643
rect 32623 597 32701 643
rect 32747 597 32825 643
rect 32871 597 32949 643
rect 32995 597 33073 643
rect 33119 597 33197 643
rect 33243 597 33321 643
rect 33367 597 33445 643
rect 33491 597 33569 643
rect 33615 597 33693 643
rect 33739 597 33817 643
rect 33863 597 33941 643
rect 33987 597 34065 643
rect 34111 597 34189 643
rect 34235 597 34313 643
rect 34359 597 34437 643
rect 34483 597 34561 643
rect 34607 597 34685 643
rect 34731 597 34809 643
rect 34855 597 34933 643
rect 34979 597 35057 643
rect 35103 597 35181 643
rect 35227 597 35305 643
rect 35351 597 35429 643
rect 35475 597 35553 643
rect 35599 597 35677 643
rect 35723 597 35801 643
rect 35847 597 35925 643
rect 35971 597 36049 643
rect 36095 597 36173 643
rect 36219 597 36297 643
rect 36343 597 36421 643
rect 36467 597 36545 643
rect 36591 597 36669 643
rect 36715 597 36793 643
rect 36839 597 36917 643
rect 36963 597 37041 643
rect 37087 597 37165 643
rect 37211 597 37289 643
rect 37335 597 37413 643
rect 37459 597 37537 643
rect 37583 597 37661 643
rect 37707 597 37785 643
rect 37831 597 37909 643
rect 37955 597 38033 643
rect 38079 597 38157 643
rect 38203 597 38281 643
rect 38327 597 38405 643
rect 38451 597 38529 643
rect 38575 597 38653 643
rect 38699 597 38777 643
rect 38823 597 38901 643
rect 38947 597 39025 643
rect 39071 597 39149 643
rect 39195 597 39273 643
rect 39319 597 39397 643
rect 39443 597 39521 643
rect 39567 597 39645 643
rect 39691 597 39769 643
rect 39815 597 39893 643
rect 39939 597 40017 643
rect 40063 597 40141 643
rect 40187 597 40265 643
rect 40311 597 40389 643
rect 40435 597 40513 643
rect 40559 597 40637 643
rect 40683 597 40761 643
rect 40807 597 40885 643
rect 40931 597 41009 643
rect 41055 597 41133 643
rect 41179 597 41257 643
rect 41303 597 41381 643
rect 41427 597 41505 643
rect 41551 597 41629 643
rect 41675 597 41753 643
rect 41799 597 41877 643
rect 41923 597 42001 643
rect 42047 597 42125 643
rect 42171 597 42249 643
rect 42295 597 42373 643
rect 42419 597 42497 643
rect 42543 597 42621 643
rect 42667 597 42745 643
rect 42791 597 42869 643
rect 42915 597 42993 643
rect 43039 597 43117 643
rect 43163 597 43241 643
rect 43287 597 43365 643
rect 43411 597 43489 643
rect 43535 597 43613 643
rect 43659 597 43737 643
rect 43783 597 43861 643
rect 43907 597 43985 643
rect 44031 597 44109 643
rect 44155 597 44233 643
rect 44279 597 44357 643
rect 44403 597 44481 643
rect 44527 597 44605 643
rect 44651 597 44729 643
rect 44775 597 44853 643
rect 44899 597 44977 643
rect 45023 597 45101 643
rect 45147 597 45225 643
rect 45271 597 45349 643
rect 45395 597 45473 643
rect 45519 597 45597 643
rect 45643 597 45721 643
rect 45767 597 45845 643
rect 45891 597 45969 643
rect 46015 597 46093 643
rect 46139 597 46217 643
rect 46263 597 46341 643
rect 46387 597 46465 643
rect 46511 597 46589 643
rect 46635 597 46713 643
rect 46759 597 46837 643
rect 46883 597 46961 643
rect 47007 597 47085 643
rect 47131 597 47209 643
rect 47255 597 47333 643
rect 47379 597 47457 643
rect 47503 597 47581 643
rect 47627 597 47705 643
rect 47751 597 47829 643
rect 47875 597 47953 643
rect 47999 597 48077 643
rect 48123 597 48201 643
rect 48247 597 48325 643
rect 48371 597 48449 643
rect 48495 597 48573 643
rect 48619 597 48697 643
rect 48743 597 48821 643
rect 48867 597 48945 643
rect 48991 597 49069 643
rect 49115 597 49193 643
rect 49239 597 49317 643
rect 49363 597 49441 643
rect 49487 597 49565 643
rect 49611 597 49689 643
rect 49735 597 49813 643
rect 49859 597 49937 643
rect 49983 597 50061 643
rect 50107 597 50185 643
rect 50231 597 50309 643
rect 50355 597 50433 643
rect 50479 597 50557 643
rect 50603 597 50681 643
rect 50727 597 50805 643
rect 50851 597 50929 643
rect 50975 597 51053 643
rect 51099 597 51177 643
rect 51223 597 51301 643
rect 51347 597 51425 643
rect 51471 597 51549 643
rect 51595 597 51673 643
rect 51719 597 51797 643
rect 51843 597 51921 643
rect 51967 597 52045 643
rect 52091 597 52169 643
rect 52215 597 52293 643
rect 52339 597 52417 643
rect 52463 597 52541 643
rect 52587 597 52665 643
rect 52711 597 52789 643
rect 52835 597 52913 643
rect 52959 597 53037 643
rect 53083 597 53161 643
rect 53207 597 53285 643
rect 53331 597 53409 643
rect 53455 597 53533 643
rect 53579 597 53657 643
rect 53703 597 53781 643
rect 53827 597 53905 643
rect 53951 597 54029 643
rect 54075 597 54153 643
rect 54199 597 54277 643
rect 54323 597 54401 643
rect 54447 597 54525 643
rect 54571 597 54649 643
rect 54695 597 54773 643
rect 54819 597 54897 643
rect 54943 597 55021 643
rect 55067 597 55145 643
rect 55191 597 55269 643
rect 55315 597 55393 643
rect 55439 597 55517 643
rect 55563 597 55641 643
rect 55687 597 55765 643
rect 55811 597 55889 643
rect 55935 597 56013 643
rect 56059 597 56137 643
rect 56183 597 56261 643
rect 56307 597 56385 643
rect 56431 597 56509 643
rect 56555 597 56633 643
rect 56679 597 56757 643
rect 56803 597 56881 643
rect 56927 597 57005 643
rect 57051 597 57129 643
rect 57175 597 57253 643
rect 57299 597 57377 643
rect 57423 597 57501 643
rect 57547 597 57625 643
rect 57671 597 57749 643
rect 57795 597 57873 643
rect 57919 597 57997 643
rect 58043 597 58121 643
rect 58167 597 58245 643
rect 58291 597 58369 643
rect 58415 597 58493 643
rect 58539 597 58617 643
rect 58663 597 58741 643
rect 58787 597 58865 643
rect 58911 597 58989 643
rect 59035 597 59113 643
rect 59159 597 59237 643
rect 59283 597 59361 643
rect 59407 597 59485 643
rect 59531 597 59609 643
rect 59655 597 59733 643
rect 59779 597 59857 643
rect 59903 597 59981 643
rect 60027 597 60105 643
rect 60151 597 60229 643
rect 60275 597 60353 643
rect 60399 597 60477 643
rect 60523 597 60601 643
rect 60647 597 60725 643
rect 60771 597 60849 643
rect 60895 597 60973 643
rect 61019 597 61097 643
rect 61143 597 61221 643
rect 61267 597 61345 643
rect 61391 597 61469 643
rect 61515 597 61593 643
rect 61639 597 61717 643
rect 61763 597 61841 643
rect 61887 597 61965 643
rect 62011 597 62089 643
rect 62135 597 62213 643
rect 62259 597 62337 643
rect 62383 597 62461 643
rect 62507 597 62585 643
rect 62631 597 62709 643
rect 62755 597 62833 643
rect 62879 597 62957 643
rect 63003 597 63081 643
rect 63127 597 63205 643
rect 63251 597 63329 643
rect 63375 597 63453 643
rect 63499 597 63577 643
rect 63623 597 63701 643
rect 63747 597 63825 643
rect 63871 597 63949 643
rect 63995 597 64073 643
rect 64119 597 64197 643
rect 64243 597 64321 643
rect 64367 597 64445 643
rect 64491 597 64569 643
rect 64615 597 64693 643
rect 64739 597 64817 643
rect 64863 597 64941 643
rect 64987 597 65065 643
rect 65111 597 65189 643
rect 65235 597 65313 643
rect 65359 597 65437 643
rect 65483 597 65561 643
rect 65607 597 65685 643
rect 65731 597 65809 643
rect 65855 597 65933 643
rect 65979 597 66057 643
rect 66103 597 66181 643
rect 66227 597 66305 643
rect 66351 597 66429 643
rect 66475 597 66553 643
rect 66599 597 66677 643
rect 66723 597 66801 643
rect 66847 597 66925 643
rect 66971 597 67049 643
rect 67095 597 67173 643
rect 67219 597 67297 643
rect 67343 597 67421 643
rect 67467 597 67545 643
rect 67591 597 67669 643
rect 67715 597 67793 643
rect 67839 597 67917 643
rect 67963 597 68041 643
rect 68087 597 68165 643
rect 68211 597 68289 643
rect 68335 597 68413 643
rect 68459 597 68537 643
rect 68583 597 68661 643
rect 68707 597 68785 643
rect 68831 597 68909 643
rect 68955 597 69033 643
rect 69079 597 69157 643
rect 69203 597 69281 643
rect 69327 597 69405 643
rect 69451 597 69529 643
rect 69575 597 69653 643
rect 69699 597 69777 643
rect 69823 597 69901 643
rect 69947 597 70025 643
rect 70071 597 70149 643
rect 70195 597 70273 643
rect 70319 597 70397 643
rect 70443 597 70521 643
rect 70567 597 70645 643
rect 70691 597 70769 643
rect 70815 597 70893 643
rect 70939 597 71017 643
rect 71063 597 71141 643
rect 71187 597 71265 643
rect 71311 597 71389 643
rect 71435 597 71513 643
rect 71559 597 71637 643
rect 71683 597 71761 643
rect 71807 597 71885 643
rect 71931 597 72009 643
rect 72055 597 72133 643
rect 72179 597 72257 643
rect 72303 597 72381 643
rect 72427 597 72505 643
rect 72551 597 72629 643
rect 72675 597 72753 643
rect 72799 597 72877 643
rect 72923 597 73001 643
rect 73047 597 73125 643
rect 73171 597 73249 643
rect 73295 597 73373 643
rect 73419 597 73497 643
rect 73543 597 73621 643
rect 73667 597 73745 643
rect 73791 597 73869 643
rect 73915 597 73993 643
rect 74039 597 74117 643
rect 74163 597 74241 643
rect 74287 597 74365 643
rect 74411 597 74489 643
rect 74535 597 74613 643
rect 74659 597 74737 643
rect 74783 597 74861 643
rect 74907 597 74985 643
rect 75031 597 75109 643
rect 75155 597 75233 643
rect 75279 597 75357 643
rect 75403 597 75481 643
rect 75527 597 75605 643
rect 75651 597 75729 643
rect 75775 597 75853 643
rect 75899 597 75977 643
rect 76023 597 76101 643
rect 76147 597 76225 643
rect 76271 597 76349 643
rect 76395 597 76473 643
rect 76519 597 76597 643
rect 76643 597 76721 643
rect 76767 597 76845 643
rect 76891 597 76969 643
rect 77015 597 77093 643
rect 77139 597 77217 643
rect 77263 597 77341 643
rect 77387 597 77465 643
rect 77511 597 77589 643
rect 77635 597 77713 643
rect 77759 597 77837 643
rect 77883 597 77961 643
rect 78007 597 78085 643
rect 78131 597 78209 643
rect 78255 597 78333 643
rect 78379 597 78457 643
rect 78503 597 78581 643
rect 78627 597 78705 643
rect 78751 597 78829 643
rect 78875 597 78953 643
rect 78999 597 79077 643
rect 79123 597 79201 643
rect 79247 597 79325 643
rect 79371 597 79449 643
rect 79495 597 79573 643
rect 79619 597 79697 643
rect 79743 597 79821 643
rect 79867 597 79945 643
rect 79991 597 80069 643
rect 80115 597 80193 643
rect 80239 597 80317 643
rect 80363 597 80441 643
rect 80487 597 80565 643
rect 80611 597 80689 643
rect 80735 597 80813 643
rect 80859 597 80937 643
rect 80983 597 81061 643
rect 81107 597 81185 643
rect 81231 597 81309 643
rect 81355 597 81433 643
rect 81479 597 81557 643
rect 81603 597 81681 643
rect 81727 597 81805 643
rect 81851 597 81929 643
rect 81975 597 82053 643
rect 82099 597 82177 643
rect 82223 597 82301 643
rect 82347 597 82425 643
rect 82471 597 82549 643
rect 82595 597 82673 643
rect 82719 597 82797 643
rect 82843 597 82921 643
rect 82967 597 83045 643
rect 83091 597 83169 643
rect 83215 597 83293 643
rect 83339 597 83417 643
rect 83463 597 83541 643
rect 83587 597 83665 643
rect 83711 597 83789 643
rect 83835 597 83913 643
rect 83959 597 84037 643
rect 84083 597 84161 643
rect 84207 597 84285 643
rect 84331 597 84409 643
rect 84455 597 84533 643
rect 84579 597 84657 643
rect 84703 597 84781 643
rect 84827 597 84905 643
rect 84951 597 85029 643
rect 85075 597 85153 643
rect 85199 597 85277 643
rect 85323 597 85401 643
rect 85447 597 85525 643
rect 85571 597 85649 643
rect 85695 597 85706 643
rect 0 586 85706 597
rect 0 403 1000 586
<< metal2 >>
rect 424 403 1424 45776
<< metal3 >>
rect 424 0 1424 2232
use M1_PSUB43105899832108_64x8m81  M1_PSUB43105899832108_64x8m81_0
timestamp 1698431365
transform -1 0 85672 0 1 45688
box 0 0 1 1
use M1_PSUB43105899832108_64x8m81  M1_PSUB43105899832108_64x8m81_1
timestamp 1698431365
transform -1 0 85672 0 1 620
box 0 0 1 1
use M1_PSUB43105899832109_64x8m81  M1_PSUB43105899832109_64x8m81_0
timestamp 1698431365
transform 1 0 85474 0 1 1140
box 0 0 1 1
use M1_PSUB43105899832109_64x8m81  M1_PSUB43105899832109_64x8m81_1
timestamp 1698431365
transform 1 0 112 0 1 1140
box 0 0 1 1
<< labels >>
flabel metal3 s 924 178 924 178 0 FreeSans 448 0 0 0 VDD
port 1 nsew
<< properties >>
string GDS_END 2255372
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 2254716
string path 4.620 11.160 4.620 0.000 
<< end >>
