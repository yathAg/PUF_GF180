magic
tech gf180mcuA
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 352 3670 870
<< pwell >>
rect -86 -86 3670 352
<< mvnmos >>
rect 124 93 244 165
rect 348 93 468 165
rect 572 93 692 165
rect 796 93 916 165
rect 980 93 1100 165
rect 1366 93 1486 165
rect 1590 93 1710 165
rect 1859 68 1979 232
rect 2083 68 2203 232
rect 2267 68 2387 232
rect 2643 68 2763 232
rect 2867 68 2987 232
rect 3091 68 3211 232
rect 3315 68 3435 232
<< mvpmos >>
rect 144 532 244 604
rect 348 532 448 604
rect 592 527 692 604
rect 796 527 896 604
rect 1000 527 1100 604
rect 1467 527 1567 604
rect 1631 527 1731 604
rect 1879 472 1979 716
rect 2083 472 2183 716
rect 2287 472 2387 716
rect 2663 472 2763 716
rect 2877 472 2977 716
rect 3101 472 3201 716
rect 3315 472 3415 716
<< mvndiff >>
rect 1770 165 1859 232
rect 36 152 124 165
rect 36 106 49 152
rect 95 106 124 152
rect 36 93 124 106
rect 244 152 348 165
rect 244 106 273 152
rect 319 106 348 152
rect 244 93 348 106
rect 468 152 572 165
rect 468 106 497 152
rect 543 106 572 152
rect 468 93 572 106
rect 692 152 796 165
rect 692 106 721 152
rect 767 106 796 152
rect 692 93 796 106
rect 916 93 980 165
rect 1100 152 1188 165
rect 1100 106 1129 152
rect 1175 106 1188 152
rect 1100 93 1188 106
rect 1278 152 1366 165
rect 1278 106 1291 152
rect 1337 106 1366 152
rect 1278 93 1366 106
rect 1486 152 1590 165
rect 1486 106 1515 152
rect 1561 106 1590 152
rect 1486 93 1590 106
rect 1710 152 1859 165
rect 1710 106 1783 152
rect 1829 106 1859 152
rect 1710 93 1859 106
rect 1770 68 1859 93
rect 1979 152 2083 232
rect 1979 106 2008 152
rect 2054 106 2083 152
rect 1979 68 2083 106
rect 2203 68 2267 232
rect 2387 128 2475 232
rect 2387 82 2416 128
rect 2462 82 2475 128
rect 2387 68 2475 82
rect 2555 191 2643 232
rect 2555 145 2568 191
rect 2614 145 2643 191
rect 2555 68 2643 145
rect 2763 157 2867 232
rect 2763 111 2792 157
rect 2838 111 2867 157
rect 2763 68 2867 111
rect 2987 191 3091 232
rect 2987 145 3016 191
rect 3062 145 3091 191
rect 2987 68 3091 145
rect 3211 157 3315 232
rect 3211 111 3240 157
rect 3286 111 3315 157
rect 3211 68 3315 111
rect 3435 191 3523 232
rect 3435 145 3464 191
rect 3510 145 3523 191
rect 3435 68 3523 145
<< mvpdiff >>
rect 1791 703 1879 716
rect 1791 604 1804 703
rect 56 591 144 604
rect 56 545 69 591
rect 115 545 144 591
rect 56 532 144 545
rect 244 532 348 604
rect 448 591 592 604
rect 448 545 477 591
rect 523 545 592 591
rect 448 532 592 545
rect 512 527 592 532
rect 692 591 796 604
rect 692 545 721 591
rect 767 545 796 591
rect 692 527 796 545
rect 896 586 1000 604
rect 896 540 925 586
rect 971 540 1000 586
rect 896 527 1000 540
rect 1100 591 1235 604
rect 1100 545 1176 591
rect 1222 545 1235 591
rect 1100 527 1235 545
rect 1379 586 1467 604
rect 1379 540 1392 586
rect 1438 540 1467 586
rect 1379 527 1467 540
rect 1567 527 1631 604
rect 1731 563 1804 604
rect 1850 563 1879 703
rect 1731 527 1879 563
rect 1791 472 1879 527
rect 1979 678 2083 716
rect 1979 632 2008 678
rect 2054 632 2083 678
rect 1979 472 2083 632
rect 2183 586 2287 716
rect 2183 540 2212 586
rect 2258 540 2287 586
rect 2183 472 2287 540
rect 2387 678 2475 716
rect 2387 632 2416 678
rect 2462 632 2475 678
rect 2387 472 2475 632
rect 2575 665 2663 716
rect 2575 525 2588 665
rect 2634 525 2663 665
rect 2575 472 2663 525
rect 2763 665 2877 716
rect 2763 619 2792 665
rect 2838 619 2877 665
rect 2763 472 2877 619
rect 2977 665 3101 716
rect 2977 525 3006 665
rect 3052 525 3101 665
rect 2977 472 3101 525
rect 3201 665 3315 716
rect 3201 619 3230 665
rect 3276 619 3315 665
rect 3201 472 3315 619
rect 3415 665 3503 716
rect 3415 525 3444 665
rect 3490 525 3503 665
rect 3415 472 3503 525
<< mvndiffc >>
rect 49 106 95 152
rect 273 106 319 152
rect 497 106 543 152
rect 721 106 767 152
rect 1129 106 1175 152
rect 1291 106 1337 152
rect 1515 106 1561 152
rect 1783 106 1829 152
rect 2008 106 2054 152
rect 2416 82 2462 128
rect 2568 145 2614 191
rect 2792 111 2838 157
rect 3016 145 3062 191
rect 3240 111 3286 157
rect 3464 145 3510 191
<< mvpdiffc >>
rect 69 545 115 591
rect 477 545 523 591
rect 721 545 767 591
rect 925 540 971 586
rect 1176 545 1222 591
rect 1392 540 1438 586
rect 1804 563 1850 703
rect 2008 632 2054 678
rect 2212 540 2258 586
rect 2416 632 2462 678
rect 2588 525 2634 665
rect 2792 619 2838 665
rect 3006 525 3052 665
rect 3230 619 3276 665
rect 3444 525 3490 665
<< polysilicon >>
rect 1879 716 1979 760
rect 2083 716 2183 760
rect 2287 716 2387 760
rect 2663 716 2763 760
rect 2877 716 2977 760
rect 3101 716 3201 760
rect 3315 716 3415 760
rect 144 604 244 648
rect 348 604 448 648
rect 592 604 692 648
rect 796 604 896 648
rect 1000 604 1100 648
rect 1467 604 1567 648
rect 1631 604 1731 648
rect 144 378 244 532
rect 144 332 175 378
rect 221 332 244 378
rect 144 209 244 332
rect 124 165 244 209
rect 348 303 448 532
rect 592 418 692 527
rect 348 257 387 303
rect 433 257 448 303
rect 348 209 448 257
rect 572 403 692 418
rect 572 357 587 403
rect 633 357 692 403
rect 348 165 468 209
rect 572 165 692 357
rect 796 304 896 527
rect 1000 467 1100 527
rect 796 258 809 304
rect 855 258 896 304
rect 796 209 896 258
rect 980 412 1100 467
rect 980 366 995 412
rect 1041 366 1100 412
rect 796 165 916 209
rect 980 165 1100 366
rect 1467 322 1567 527
rect 1366 307 1567 322
rect 1366 261 1393 307
rect 1439 282 1567 307
rect 1631 483 1731 527
rect 1631 412 1710 483
rect 1631 366 1651 412
rect 1697 366 1710 412
rect 1439 261 1486 282
rect 1366 165 1486 261
rect 1631 232 1710 366
rect 1879 312 1979 472
rect 1879 288 1892 312
rect 1859 266 1892 288
rect 1938 266 1979 312
rect 1859 232 1979 266
rect 2083 312 2183 472
rect 2083 266 2110 312
rect 2156 288 2183 312
rect 2287 423 2387 472
rect 2287 377 2300 423
rect 2346 377 2387 423
rect 2287 288 2387 377
rect 2663 412 2763 472
rect 2877 412 2977 472
rect 3101 412 3201 472
rect 3315 412 3415 472
rect 2663 399 3415 412
rect 2663 353 2683 399
rect 3387 353 3415 399
rect 2663 340 3415 353
rect 2663 288 2763 340
rect 2156 266 2203 288
rect 2083 232 2203 266
rect 2267 232 2387 288
rect 2643 232 2763 288
rect 2867 232 2987 340
rect 3091 232 3211 340
rect 3315 288 3415 340
rect 3315 232 3435 288
rect 1590 165 1710 232
rect 124 49 244 93
rect 348 49 468 93
rect 572 49 692 93
rect 796 49 916 93
rect 980 49 1100 93
rect 1366 49 1486 93
rect 1590 49 1710 93
rect 1859 24 1979 68
rect 2083 24 2203 68
rect 2267 24 2387 68
rect 2643 24 2763 68
rect 2867 24 2987 68
rect 3091 24 3211 68
rect 3315 24 3435 68
<< polycontact >>
rect 175 332 221 378
rect 387 257 433 303
rect 587 357 633 403
rect 809 258 855 304
rect 995 366 1041 412
rect 1393 261 1439 307
rect 1651 366 1697 412
rect 1892 266 1938 312
rect 2110 266 2156 312
rect 2300 377 2346 423
rect 2683 353 3387 399
<< metal1 >>
rect 0 724 3584 844
rect 69 591 115 603
rect 466 591 534 724
rect 1793 703 1861 724
rect 466 545 477 591
rect 523 545 534 591
rect 710 632 1233 678
rect 710 591 778 632
rect 710 545 721 591
rect 767 545 778 591
rect 1165 591 1233 632
rect 69 245 115 545
rect 914 540 925 586
rect 971 540 982 586
rect 1165 545 1176 591
rect 1222 545 1233 591
rect 1279 632 1678 678
rect 914 511 982 540
rect 914 499 1134 511
rect 1279 499 1325 632
rect 175 453 778 499
rect 914 465 1325 499
rect 1088 453 1325 465
rect 175 378 221 453
rect 690 419 778 453
rect 690 412 1052 419
rect 175 313 221 332
rect 284 403 644 407
rect 284 357 587 403
rect 633 357 644 403
rect 690 366 995 412
rect 1041 366 1052 412
rect 690 364 1052 366
rect 284 353 644 357
rect 284 245 330 353
rect 1279 307 1325 453
rect 1381 540 1392 586
rect 1438 540 1449 586
rect 1381 419 1449 540
rect 1623 511 1678 632
rect 1793 563 1804 703
rect 1850 563 1861 703
rect 1979 632 2008 678
rect 2054 632 2416 678
rect 2462 632 2475 678
rect 2588 665 2634 676
rect 1793 557 1861 563
rect 2183 540 2212 586
rect 2258 540 2475 586
rect 1623 465 2147 511
rect 2101 436 2147 465
rect 2101 423 2352 436
rect 1381 360 1572 419
rect 1635 412 2055 419
rect 1635 366 1651 412
rect 1697 366 2055 412
rect 1635 360 2055 366
rect 2101 377 2300 423
rect 2346 377 2352 423
rect 2101 364 2352 377
rect 2429 399 2475 540
rect 2792 665 2838 724
rect 2792 603 2838 619
rect 3006 665 3052 676
rect 2634 525 3006 536
rect 3230 665 3276 724
rect 3230 603 3276 619
rect 3444 665 3555 676
rect 3052 525 3444 536
rect 3490 525 3555 665
rect 2588 472 3555 525
rect 376 304 884 307
rect 376 303 809 304
rect 376 257 387 303
rect 433 258 809 303
rect 855 258 884 304
rect 433 257 884 258
rect 376 248 884 257
rect 1023 261 1393 307
rect 1439 261 1455 307
rect 1023 260 1455 261
rect 1504 261 1572 360
rect 2004 313 2055 360
rect 2429 353 2683 399
rect 3387 353 3412 399
rect 2004 312 2230 313
rect 1881 266 1892 312
rect 1938 266 1949 312
rect 1881 261 1949 266
rect 69 198 330 245
rect 262 152 330 198
rect 1023 152 1069 260
rect 1504 215 1949 261
rect 2004 266 2110 312
rect 2156 266 2230 312
rect 2429 297 2475 353
rect 3464 307 3555 472
rect 2004 251 2230 266
rect 2313 251 2475 297
rect 2568 252 3555 307
rect 1504 152 1572 215
rect 38 106 49 152
rect 95 106 106 152
rect 262 106 273 152
rect 319 106 330 152
rect 486 106 497 152
rect 543 106 554 152
rect 710 106 721 152
rect 767 106 1069 152
rect 1118 106 1129 152
rect 1175 106 1291 152
rect 1337 106 1348 152
rect 1504 106 1515 152
rect 1561 106 1572 152
rect 1783 152 1829 168
rect 2313 152 2359 251
rect 1979 106 2008 152
rect 2054 106 2359 152
rect 2568 191 2614 252
rect 3016 191 3062 252
rect 2568 131 2614 145
rect 2792 157 2838 181
rect 38 60 106 106
rect 486 60 554 106
rect 1118 60 1348 106
rect 1783 60 1829 106
rect 2405 82 2416 128
rect 2462 82 2473 128
rect 2405 60 2473 82
rect 3464 191 3555 252
rect 3016 131 3062 145
rect 3240 157 3286 181
rect 2792 60 2838 111
rect 3510 145 3555 191
rect 3464 120 3555 145
rect 3240 60 3286 111
rect 0 -60 3584 60
<< labels >>
flabel metal1 s 1635 360 2055 419 0 FreeSans 400 0 0 0 A3
port 3 nsew default input
flabel metal1 s 0 724 3584 844 0 FreeSans 400 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 3240 168 3286 181 0 FreeSans 400 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel metal1 s 3444 536 3555 676 0 FreeSans 400 0 0 0 ZN
port 4 nsew default output
flabel metal1 s 376 248 884 307 0 FreeSans 400 0 0 0 A1
port 1 nsew default input
flabel metal1 s 175 453 778 499 0 FreeSans 400 0 0 0 A2
port 2 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 6 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 690 419 778 453 1 A2
port 2 nsew default input
rlabel metal1 s 175 419 221 453 1 A2
port 2 nsew default input
rlabel metal1 s 690 364 1052 419 1 A2
port 2 nsew default input
rlabel metal1 s 175 364 221 419 1 A2
port 2 nsew default input
rlabel metal1 s 175 313 221 364 1 A2
port 2 nsew default input
rlabel metal1 s 2004 313 2055 360 1 A3
port 3 nsew default input
rlabel metal1 s 2004 251 2230 313 1 A3
port 3 nsew default input
rlabel metal1 s 3006 536 3052 676 1 ZN
port 4 nsew default output
rlabel metal1 s 2588 536 2634 676 1 ZN
port 4 nsew default output
rlabel metal1 s 2588 472 3555 536 1 ZN
port 4 nsew default output
rlabel metal1 s 3464 307 3555 472 1 ZN
port 4 nsew default output
rlabel metal1 s 2568 252 3555 307 1 ZN
port 4 nsew default output
rlabel metal1 s 3464 131 3555 252 1 ZN
port 4 nsew default output
rlabel metal1 s 3016 131 3062 252 1 ZN
port 4 nsew default output
rlabel metal1 s 2568 131 2614 252 1 ZN
port 4 nsew default output
rlabel metal1 s 3464 120 3555 131 1 ZN
port 4 nsew default output
rlabel metal1 s 3230 603 3276 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2792 603 2838 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1793 603 1861 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 466 603 534 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1793 557 1861 603 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 466 557 534 603 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 466 545 534 557 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2792 168 2838 181 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3240 152 3286 168 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2792 152 2838 168 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1783 152 1829 168 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3240 128 3286 152 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2792 128 2838 152 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1783 128 1829 152 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1118 128 1348 152 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 486 128 554 152 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 38 128 106 152 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3240 60 3286 128 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2792 60 2838 128 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2405 60 2473 128 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1783 60 1829 128 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1118 60 1348 128 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 486 60 554 128 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 38 60 106 128 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3584 60 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3584 784
string GDS_END 356348
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 348300
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
