magic
tech gf180mcuA
magscale 1 10
timestamp 1698431365
<< nwell >>
rect 1980 15510 4160 15514
rect 461 14569 4160 15510
rect 6583 15258 9560 15532
rect 13849 15258 15116 15548
rect 23608 15510 25788 15514
rect 6583 14608 11141 15258
rect 13849 15181 15441 15258
rect 13850 14608 15441 15181
rect 6583 14607 9382 14608
rect 461 -209 2610 14569
rect 6583 14558 8962 14607
rect 16520 14576 21087 15503
rect 23608 14569 27308 15510
rect 25159 -209 27308 14569
<< mvnmos >>
rect 4324 14872 6346 14992
rect 11385 14872 11913 14992
rect 12286 14873 13604 14993
rect 15755 14872 16283 14992
rect 21324 14872 23346 14992
<< mvpmos >>
rect 597 14456 1696 15244
rect 6719 15096 9245 15216
rect 6719 14872 9245 14992
rect 9686 14872 11004 14992
rect 13986 14872 15304 14992
rect 16656 14872 17974 14992
rect 18424 15096 20950 15216
rect 18424 14872 20950 14992
rect 597 13556 1696 14344
rect 597 12656 1696 13444
rect 597 11756 1696 12544
rect 597 10856 1696 11644
rect 597 9956 1696 10744
rect 597 9056 1696 9844
rect 597 8156 1696 8944
rect 597 7256 1696 8044
rect 597 6356 1696 7144
rect 597 5456 1696 6244
rect 597 4556 1696 5344
rect 597 3656 1696 4444
rect 597 2756 1696 3544
rect 597 1856 1696 2644
rect 597 956 1696 1744
rect 597 56 1696 844
rect 26073 14456 27172 15244
rect 26073 13556 27172 14344
rect 26073 12656 27172 13444
rect 26073 11756 27172 12544
rect 26073 10856 27172 11644
rect 26073 9956 27172 10744
rect 26073 9056 27172 9844
rect 26073 8156 27172 8944
rect 26073 7256 27172 8044
rect 26073 6356 27172 7144
rect 26073 5456 27172 6244
rect 26073 4556 27172 5344
rect 26073 3656 27172 4444
rect 26073 2756 27172 3544
rect 26073 1856 27172 2644
rect 26073 956 27172 1744
rect 26073 56 27172 844
<< mvndiff >>
rect 4324 15067 6346 15080
rect 4324 15021 4337 15067
rect 5097 15021 5154 15067
rect 5200 15021 5257 15067
rect 5303 15021 5360 15067
rect 5406 15021 5463 15067
rect 5509 15021 5566 15067
rect 5612 15021 5669 15067
rect 5715 15021 5772 15067
rect 5818 15021 5875 15067
rect 5921 15021 5978 15067
rect 6024 15021 6081 15067
rect 6127 15021 6184 15067
rect 6230 15021 6287 15067
rect 6333 15021 6346 15067
rect 4324 14992 6346 15021
rect 11385 15067 11913 15080
rect 11385 15021 11398 15067
rect 11444 15021 11512 15067
rect 11558 15021 11626 15067
rect 11672 15021 11740 15067
rect 11786 15021 11854 15067
rect 11900 15021 11913 15067
rect 12286 15068 13604 15081
rect 11385 14992 11913 15021
rect 12286 15022 12299 15068
rect 12345 15022 12402 15068
rect 12448 15022 12505 15068
rect 12551 15022 12609 15068
rect 12655 15022 12713 15068
rect 12759 15022 12817 15068
rect 12863 15022 12921 15068
rect 12967 15022 13025 15068
rect 13071 15022 13129 15068
rect 13175 15022 13233 15068
rect 13279 15022 13337 15068
rect 13383 15022 13441 15068
rect 13487 15022 13545 15068
rect 13591 15022 13604 15068
rect 12286 14993 13604 15022
rect 4324 14843 6346 14872
rect 4324 14797 4337 14843
rect 5097 14797 5154 14843
rect 5200 14797 5257 14843
rect 5303 14797 5360 14843
rect 5406 14797 5463 14843
rect 5509 14797 5566 14843
rect 5612 14797 5669 14843
rect 5715 14797 5772 14843
rect 5818 14797 5875 14843
rect 5921 14797 5978 14843
rect 6024 14797 6081 14843
rect 6127 14797 6184 14843
rect 6230 14797 6287 14843
rect 6333 14797 6346 14843
rect 4324 14784 6346 14797
rect 11385 14843 11913 14872
rect 11385 14797 11398 14843
rect 11444 14797 11512 14843
rect 11558 14797 11626 14843
rect 11672 14797 11740 14843
rect 11786 14797 11854 14843
rect 11900 14797 11913 14843
rect 11385 14784 11913 14797
rect 12286 14844 13604 14873
rect 15755 15067 16283 15080
rect 15755 15021 15768 15067
rect 15814 15021 15882 15067
rect 15928 15021 15996 15067
rect 16042 15021 16110 15067
rect 16156 15021 16224 15067
rect 16270 15021 16283 15067
rect 15755 14992 16283 15021
rect 21324 15067 23346 15080
rect 21324 15021 21337 15067
rect 22097 15021 22154 15067
rect 22200 15021 22257 15067
rect 22303 15021 22360 15067
rect 22406 15021 22463 15067
rect 22509 15021 22566 15067
rect 22612 15021 22669 15067
rect 22715 15021 22772 15067
rect 22818 15021 22875 15067
rect 22921 15021 22978 15067
rect 23024 15021 23081 15067
rect 23127 15021 23184 15067
rect 23230 15021 23287 15067
rect 23333 15021 23346 15067
rect 21324 14992 23346 15021
rect 12286 14798 12299 14844
rect 12345 14798 12402 14844
rect 12448 14798 12505 14844
rect 12551 14798 12609 14844
rect 12655 14798 12713 14844
rect 12759 14798 12817 14844
rect 12863 14798 12921 14844
rect 12967 14798 13025 14844
rect 13071 14798 13129 14844
rect 13175 14798 13233 14844
rect 13279 14798 13337 14844
rect 13383 14798 13441 14844
rect 13487 14798 13545 14844
rect 13591 14798 13604 14844
rect 12286 14785 13604 14798
rect 15755 14843 16283 14872
rect 15755 14797 15768 14843
rect 15814 14797 15882 14843
rect 15928 14797 15996 14843
rect 16042 14797 16110 14843
rect 16156 14797 16224 14843
rect 16270 14797 16283 14843
rect 15755 14784 16283 14797
rect 21324 14843 23346 14872
rect 21324 14797 21337 14843
rect 22097 14797 22154 14843
rect 22200 14797 22257 14843
rect 22303 14797 22360 14843
rect 22406 14797 22463 14843
rect 22509 14797 22566 14843
rect 22612 14797 22669 14843
rect 22715 14797 22772 14843
rect 22818 14797 22875 14843
rect 22921 14797 22978 14843
rect 23024 14797 23081 14843
rect 23127 14797 23184 14843
rect 23230 14797 23287 14843
rect 23333 14797 23346 14843
rect 21324 14784 23346 14797
<< mvpdiff >>
rect 597 15323 1696 15369
rect 597 15277 640 15323
rect 686 15277 801 15323
rect 847 15277 961 15323
rect 1007 15277 1121 15323
rect 1167 15277 1282 15323
rect 1328 15277 1444 15323
rect 1490 15277 1607 15323
rect 1653 15277 1696 15323
rect 597 15244 1696 15277
rect 6719 15291 9245 15304
rect 6719 15245 6732 15291
rect 8614 15245 8671 15291
rect 8717 15245 8774 15291
rect 8820 15245 8877 15291
rect 8923 15245 8980 15291
rect 9026 15245 9083 15291
rect 9129 15245 9186 15291
rect 9232 15245 9245 15291
rect 6719 15216 9245 15245
rect 6719 15067 9245 15096
rect 6719 15021 6732 15067
rect 8614 15021 8671 15067
rect 8717 15021 8774 15067
rect 8820 15021 8877 15067
rect 8923 15021 8980 15067
rect 9026 15021 9083 15067
rect 9129 15021 9186 15067
rect 9232 15021 9245 15067
rect 6719 14992 9245 15021
rect 9686 15067 11004 15080
rect 9686 15021 9699 15067
rect 9745 15021 9802 15067
rect 9848 15021 9905 15067
rect 9951 15021 10009 15067
rect 10055 15021 10113 15067
rect 10159 15021 10217 15067
rect 10263 15021 10321 15067
rect 10367 15021 10425 15067
rect 10471 15021 10529 15067
rect 10575 15021 10633 15067
rect 10679 15021 10737 15067
rect 10783 15021 10841 15067
rect 10887 15021 10945 15067
rect 10991 15021 11004 15067
rect 9686 14992 11004 15021
rect 13986 15067 15304 15080
rect 13986 15021 13999 15067
rect 14045 15021 14102 15067
rect 14148 15021 14205 15067
rect 14251 15021 14309 15067
rect 14355 15021 14413 15067
rect 14459 15021 14517 15067
rect 14563 15021 14621 15067
rect 14667 15021 14725 15067
rect 14771 15021 14829 15067
rect 14875 15021 14933 15067
rect 14979 15021 15037 15067
rect 15083 15021 15141 15067
rect 15187 15021 15245 15067
rect 15291 15021 15304 15067
rect 13986 14992 15304 15021
rect 18424 15291 20950 15304
rect 18424 15245 18437 15291
rect 20319 15245 20376 15291
rect 20422 15245 20479 15291
rect 20525 15245 20582 15291
rect 20628 15245 20685 15291
rect 20731 15245 20788 15291
rect 20834 15245 20891 15291
rect 20937 15245 20950 15291
rect 18424 15216 20950 15245
rect 6719 14843 9245 14872
rect 6719 14797 6732 14843
rect 8614 14797 8671 14843
rect 8717 14797 8774 14843
rect 8820 14797 8877 14843
rect 8923 14797 8980 14843
rect 9026 14797 9083 14843
rect 9129 14797 9186 14843
rect 9232 14797 9245 14843
rect 6719 14784 9245 14797
rect 9686 14843 11004 14872
rect 9686 14797 9699 14843
rect 9745 14797 9802 14843
rect 9848 14797 9905 14843
rect 9951 14797 10009 14843
rect 10055 14797 10113 14843
rect 10159 14797 10217 14843
rect 10263 14797 10321 14843
rect 10367 14797 10425 14843
rect 10471 14797 10529 14843
rect 10575 14797 10633 14843
rect 10679 14797 10737 14843
rect 10783 14797 10841 14843
rect 10887 14797 10945 14843
rect 10991 14797 11004 14843
rect 9686 14784 11004 14797
rect 16656 15067 17974 15080
rect 16656 15021 16669 15067
rect 16715 15021 16772 15067
rect 16818 15021 16875 15067
rect 16921 15021 16979 15067
rect 17025 15021 17083 15067
rect 17129 15021 17187 15067
rect 17233 15021 17291 15067
rect 17337 15021 17395 15067
rect 17441 15021 17499 15067
rect 17545 15021 17603 15067
rect 17649 15021 17707 15067
rect 17753 15021 17811 15067
rect 17857 15021 17915 15067
rect 17961 15021 17974 15067
rect 16656 14992 17974 15021
rect 18424 15067 20950 15096
rect 18424 15021 18437 15067
rect 20319 15021 20376 15067
rect 20422 15021 20479 15067
rect 20525 15021 20582 15067
rect 20628 15021 20685 15067
rect 20731 15021 20788 15067
rect 20834 15021 20891 15067
rect 20937 15021 20950 15067
rect 18424 14992 20950 15021
rect 26073 15323 27172 15369
rect 26073 15277 26116 15323
rect 26162 15277 26279 15323
rect 26325 15277 26441 15323
rect 26487 15277 26602 15323
rect 26648 15277 26762 15323
rect 26808 15277 26922 15323
rect 26968 15277 27083 15323
rect 27129 15277 27172 15323
rect 26073 15244 27172 15277
rect 13986 14843 15304 14872
rect 13986 14797 13999 14843
rect 14045 14797 14102 14843
rect 14148 14797 14205 14843
rect 14251 14797 14309 14843
rect 14355 14797 14413 14843
rect 14459 14797 14517 14843
rect 14563 14797 14621 14843
rect 14667 14797 14725 14843
rect 14771 14797 14829 14843
rect 14875 14797 14933 14843
rect 14979 14797 15037 14843
rect 15083 14797 15141 14843
rect 15187 14797 15245 14843
rect 15291 14797 15304 14843
rect 13986 14784 15304 14797
rect 16656 14843 17974 14872
rect 16656 14797 16669 14843
rect 16715 14797 16772 14843
rect 16818 14797 16875 14843
rect 16921 14797 16979 14843
rect 17025 14797 17083 14843
rect 17129 14797 17187 14843
rect 17233 14797 17291 14843
rect 17337 14797 17395 14843
rect 17441 14797 17499 14843
rect 17545 14797 17603 14843
rect 17649 14797 17707 14843
rect 17753 14797 17811 14843
rect 17857 14797 17915 14843
rect 17961 14797 17974 14843
rect 16656 14784 17974 14797
rect 18424 14843 20950 14872
rect 18424 14797 18437 14843
rect 20319 14797 20376 14843
rect 20422 14797 20479 14843
rect 20525 14797 20582 14843
rect 20628 14797 20685 14843
rect 20731 14797 20788 14843
rect 20834 14797 20891 14843
rect 20937 14797 20950 14843
rect 18424 14784 20950 14797
rect 597 14423 1696 14456
rect 597 14377 640 14423
rect 686 14377 801 14423
rect 847 14377 961 14423
rect 1007 14377 1121 14423
rect 1167 14377 1282 14423
rect 1328 14377 1444 14423
rect 1490 14377 1607 14423
rect 1653 14377 1696 14423
rect 597 14344 1696 14377
rect 597 13523 1696 13556
rect 597 13477 640 13523
rect 686 13477 801 13523
rect 847 13477 961 13523
rect 1007 13477 1121 13523
rect 1167 13477 1282 13523
rect 1328 13477 1444 13523
rect 1490 13477 1607 13523
rect 1653 13477 1696 13523
rect 597 13444 1696 13477
rect 597 12623 1696 12656
rect 597 12577 640 12623
rect 686 12577 801 12623
rect 847 12577 961 12623
rect 1007 12577 1121 12623
rect 1167 12577 1282 12623
rect 1328 12577 1444 12623
rect 1490 12577 1607 12623
rect 1653 12577 1696 12623
rect 597 12544 1696 12577
rect 597 11723 1696 11756
rect 597 11677 640 11723
rect 686 11677 801 11723
rect 847 11677 961 11723
rect 1007 11677 1121 11723
rect 1167 11677 1282 11723
rect 1328 11677 1444 11723
rect 1490 11677 1607 11723
rect 1653 11677 1696 11723
rect 597 11644 1696 11677
rect 597 10823 1696 10856
rect 597 10777 640 10823
rect 686 10777 801 10823
rect 847 10777 961 10823
rect 1007 10777 1121 10823
rect 1167 10777 1282 10823
rect 1328 10777 1444 10823
rect 1490 10777 1607 10823
rect 1653 10777 1696 10823
rect 597 10744 1696 10777
rect 597 9923 1696 9956
rect 597 9877 640 9923
rect 686 9877 801 9923
rect 847 9877 961 9923
rect 1007 9877 1121 9923
rect 1167 9877 1282 9923
rect 1328 9877 1444 9923
rect 1490 9877 1607 9923
rect 1653 9877 1696 9923
rect 597 9844 1696 9877
rect 597 9023 1696 9056
rect 597 8977 640 9023
rect 686 8977 801 9023
rect 847 8977 961 9023
rect 1007 8977 1121 9023
rect 1167 8977 1282 9023
rect 1328 8977 1444 9023
rect 1490 8977 1607 9023
rect 1653 8977 1696 9023
rect 597 8944 1696 8977
rect 597 8123 1696 8156
rect 597 8077 640 8123
rect 686 8077 801 8123
rect 847 8077 961 8123
rect 1007 8077 1121 8123
rect 1167 8077 1282 8123
rect 1328 8077 1444 8123
rect 1490 8077 1607 8123
rect 1653 8077 1696 8123
rect 597 8044 1696 8077
rect 597 7223 1696 7256
rect 597 7177 640 7223
rect 686 7177 801 7223
rect 847 7177 961 7223
rect 1007 7177 1121 7223
rect 1167 7177 1282 7223
rect 1328 7177 1444 7223
rect 1490 7177 1607 7223
rect 1653 7177 1696 7223
rect 597 7144 1696 7177
rect 597 6323 1696 6356
rect 597 6277 640 6323
rect 686 6277 801 6323
rect 847 6277 961 6323
rect 1007 6277 1121 6323
rect 1167 6277 1282 6323
rect 1328 6277 1444 6323
rect 1490 6277 1607 6323
rect 1653 6277 1696 6323
rect 597 6244 1696 6277
rect 597 5423 1696 5456
rect 597 5377 640 5423
rect 686 5377 801 5423
rect 847 5377 961 5423
rect 1007 5377 1121 5423
rect 1167 5377 1282 5423
rect 1328 5377 1444 5423
rect 1490 5377 1607 5423
rect 1653 5377 1696 5423
rect 597 5344 1696 5377
rect 597 4523 1696 4556
rect 597 4477 640 4523
rect 686 4477 801 4523
rect 847 4477 961 4523
rect 1007 4477 1121 4523
rect 1167 4477 1282 4523
rect 1328 4477 1444 4523
rect 1490 4477 1607 4523
rect 1653 4477 1696 4523
rect 597 4444 1696 4477
rect 597 3623 1696 3656
rect 597 3577 640 3623
rect 686 3577 801 3623
rect 847 3577 961 3623
rect 1007 3577 1121 3623
rect 1167 3577 1282 3623
rect 1328 3577 1444 3623
rect 1490 3577 1607 3623
rect 1653 3577 1696 3623
rect 597 3544 1696 3577
rect 597 2723 1696 2756
rect 597 2677 640 2723
rect 686 2677 801 2723
rect 847 2677 961 2723
rect 1007 2677 1121 2723
rect 1167 2677 1282 2723
rect 1328 2677 1444 2723
rect 1490 2677 1607 2723
rect 1653 2677 1696 2723
rect 597 2644 1696 2677
rect 597 1823 1696 1856
rect 597 1777 640 1823
rect 686 1777 801 1823
rect 847 1777 961 1823
rect 1007 1777 1121 1823
rect 1167 1777 1282 1823
rect 1328 1777 1444 1823
rect 1490 1777 1607 1823
rect 1653 1777 1696 1823
rect 597 1744 1696 1777
rect 597 923 1696 956
rect 597 877 640 923
rect 686 877 801 923
rect 847 877 961 923
rect 1007 877 1121 923
rect 1167 877 1282 923
rect 1328 877 1444 923
rect 1490 877 1607 923
rect 1653 877 1696 923
rect 597 844 1696 877
rect 597 23 1696 56
rect 597 -23 640 23
rect 686 -23 801 23
rect 847 -23 961 23
rect 1007 -23 1121 23
rect 1167 -23 1282 23
rect 1328 -23 1444 23
rect 1490 -23 1607 23
rect 1653 -23 1696 23
rect 597 -69 1696 -23
rect 26073 14423 27172 14456
rect 26073 14377 26116 14423
rect 26162 14377 26279 14423
rect 26325 14377 26441 14423
rect 26487 14377 26602 14423
rect 26648 14377 26762 14423
rect 26808 14377 26922 14423
rect 26968 14377 27083 14423
rect 27129 14377 27172 14423
rect 26073 14344 27172 14377
rect 26073 13523 27172 13556
rect 26073 13477 26116 13523
rect 26162 13477 26279 13523
rect 26325 13477 26441 13523
rect 26487 13477 26602 13523
rect 26648 13477 26762 13523
rect 26808 13477 26922 13523
rect 26968 13477 27083 13523
rect 27129 13477 27172 13523
rect 26073 13444 27172 13477
rect 26073 12623 27172 12656
rect 26073 12577 26116 12623
rect 26162 12577 26279 12623
rect 26325 12577 26441 12623
rect 26487 12577 26602 12623
rect 26648 12577 26762 12623
rect 26808 12577 26922 12623
rect 26968 12577 27083 12623
rect 27129 12577 27172 12623
rect 26073 12544 27172 12577
rect 26073 11723 27172 11756
rect 26073 11677 26116 11723
rect 26162 11677 26279 11723
rect 26325 11677 26441 11723
rect 26487 11677 26602 11723
rect 26648 11677 26762 11723
rect 26808 11677 26922 11723
rect 26968 11677 27083 11723
rect 27129 11677 27172 11723
rect 26073 11644 27172 11677
rect 26073 10823 27172 10856
rect 26073 10777 26116 10823
rect 26162 10777 26279 10823
rect 26325 10777 26441 10823
rect 26487 10777 26602 10823
rect 26648 10777 26762 10823
rect 26808 10777 26922 10823
rect 26968 10777 27083 10823
rect 27129 10777 27172 10823
rect 26073 10744 27172 10777
rect 26073 9923 27172 9956
rect 26073 9877 26116 9923
rect 26162 9877 26279 9923
rect 26325 9877 26441 9923
rect 26487 9877 26602 9923
rect 26648 9877 26762 9923
rect 26808 9877 26922 9923
rect 26968 9877 27083 9923
rect 27129 9877 27172 9923
rect 26073 9844 27172 9877
rect 26073 9023 27172 9056
rect 26073 8977 26116 9023
rect 26162 8977 26279 9023
rect 26325 8977 26441 9023
rect 26487 8977 26602 9023
rect 26648 8977 26762 9023
rect 26808 8977 26922 9023
rect 26968 8977 27083 9023
rect 27129 8977 27172 9023
rect 26073 8944 27172 8977
rect 26073 8123 27172 8156
rect 26073 8077 26116 8123
rect 26162 8077 26279 8123
rect 26325 8077 26441 8123
rect 26487 8077 26602 8123
rect 26648 8077 26762 8123
rect 26808 8077 26922 8123
rect 26968 8077 27083 8123
rect 27129 8077 27172 8123
rect 26073 8044 27172 8077
rect 26073 7223 27172 7256
rect 26073 7177 26116 7223
rect 26162 7177 26279 7223
rect 26325 7177 26441 7223
rect 26487 7177 26602 7223
rect 26648 7177 26762 7223
rect 26808 7177 26922 7223
rect 26968 7177 27083 7223
rect 27129 7177 27172 7223
rect 26073 7144 27172 7177
rect 26073 6323 27172 6356
rect 26073 6277 26116 6323
rect 26162 6277 26279 6323
rect 26325 6277 26441 6323
rect 26487 6277 26602 6323
rect 26648 6277 26762 6323
rect 26808 6277 26922 6323
rect 26968 6277 27083 6323
rect 27129 6277 27172 6323
rect 26073 6244 27172 6277
rect 26073 5423 27172 5456
rect 26073 5377 26116 5423
rect 26162 5377 26279 5423
rect 26325 5377 26441 5423
rect 26487 5377 26602 5423
rect 26648 5377 26762 5423
rect 26808 5377 26922 5423
rect 26968 5377 27083 5423
rect 27129 5377 27172 5423
rect 26073 5344 27172 5377
rect 26073 4523 27172 4556
rect 26073 4477 26116 4523
rect 26162 4477 26279 4523
rect 26325 4477 26441 4523
rect 26487 4477 26602 4523
rect 26648 4477 26762 4523
rect 26808 4477 26922 4523
rect 26968 4477 27083 4523
rect 27129 4477 27172 4523
rect 26073 4444 27172 4477
rect 26073 3623 27172 3656
rect 26073 3577 26116 3623
rect 26162 3577 26279 3623
rect 26325 3577 26441 3623
rect 26487 3577 26602 3623
rect 26648 3577 26762 3623
rect 26808 3577 26922 3623
rect 26968 3577 27083 3623
rect 27129 3577 27172 3623
rect 26073 3544 27172 3577
rect 26073 2723 27172 2756
rect 26073 2677 26116 2723
rect 26162 2677 26279 2723
rect 26325 2677 26441 2723
rect 26487 2677 26602 2723
rect 26648 2677 26762 2723
rect 26808 2677 26922 2723
rect 26968 2677 27083 2723
rect 27129 2677 27172 2723
rect 26073 2644 27172 2677
rect 26073 1823 27172 1856
rect 26073 1777 26116 1823
rect 26162 1777 26279 1823
rect 26325 1777 26441 1823
rect 26487 1777 26602 1823
rect 26648 1777 26762 1823
rect 26808 1777 26922 1823
rect 26968 1777 27083 1823
rect 27129 1777 27172 1823
rect 26073 1744 27172 1777
rect 26073 923 27172 956
rect 26073 877 26116 923
rect 26162 877 26279 923
rect 26325 877 26441 923
rect 26487 877 26602 923
rect 26648 877 26762 923
rect 26808 877 26922 923
rect 26968 877 27083 923
rect 27129 877 27172 923
rect 26073 844 27172 877
rect 26073 23 27172 56
rect 26073 -23 26116 23
rect 26162 -23 26279 23
rect 26325 -23 26441 23
rect 26487 -23 26602 23
rect 26648 -23 26762 23
rect 26808 -23 26922 23
rect 26968 -23 27083 23
rect 27129 -23 27172 23
rect 26073 -69 27172 -23
<< mvndiffc >>
rect 4337 15021 5097 15067
rect 5154 15021 5200 15067
rect 5257 15021 5303 15067
rect 5360 15021 5406 15067
rect 5463 15021 5509 15067
rect 5566 15021 5612 15067
rect 5669 15021 5715 15067
rect 5772 15021 5818 15067
rect 5875 15021 5921 15067
rect 5978 15021 6024 15067
rect 6081 15021 6127 15067
rect 6184 15021 6230 15067
rect 6287 15021 6333 15067
rect 11398 15021 11444 15067
rect 11512 15021 11558 15067
rect 11626 15021 11672 15067
rect 11740 15021 11786 15067
rect 11854 15021 11900 15067
rect 12299 15022 12345 15068
rect 12402 15022 12448 15068
rect 12505 15022 12551 15068
rect 12609 15022 12655 15068
rect 12713 15022 12759 15068
rect 12817 15022 12863 15068
rect 12921 15022 12967 15068
rect 13025 15022 13071 15068
rect 13129 15022 13175 15068
rect 13233 15022 13279 15068
rect 13337 15022 13383 15068
rect 13441 15022 13487 15068
rect 13545 15022 13591 15068
rect 4337 14797 5097 14843
rect 5154 14797 5200 14843
rect 5257 14797 5303 14843
rect 5360 14797 5406 14843
rect 5463 14797 5509 14843
rect 5566 14797 5612 14843
rect 5669 14797 5715 14843
rect 5772 14797 5818 14843
rect 5875 14797 5921 14843
rect 5978 14797 6024 14843
rect 6081 14797 6127 14843
rect 6184 14797 6230 14843
rect 6287 14797 6333 14843
rect 11398 14797 11444 14843
rect 11512 14797 11558 14843
rect 11626 14797 11672 14843
rect 11740 14797 11786 14843
rect 11854 14797 11900 14843
rect 15768 15021 15814 15067
rect 15882 15021 15928 15067
rect 15996 15021 16042 15067
rect 16110 15021 16156 15067
rect 16224 15021 16270 15067
rect 21337 15021 22097 15067
rect 22154 15021 22200 15067
rect 22257 15021 22303 15067
rect 22360 15021 22406 15067
rect 22463 15021 22509 15067
rect 22566 15021 22612 15067
rect 22669 15021 22715 15067
rect 22772 15021 22818 15067
rect 22875 15021 22921 15067
rect 22978 15021 23024 15067
rect 23081 15021 23127 15067
rect 23184 15021 23230 15067
rect 23287 15021 23333 15067
rect 12299 14798 12345 14844
rect 12402 14798 12448 14844
rect 12505 14798 12551 14844
rect 12609 14798 12655 14844
rect 12713 14798 12759 14844
rect 12817 14798 12863 14844
rect 12921 14798 12967 14844
rect 13025 14798 13071 14844
rect 13129 14798 13175 14844
rect 13233 14798 13279 14844
rect 13337 14798 13383 14844
rect 13441 14798 13487 14844
rect 13545 14798 13591 14844
rect 15768 14797 15814 14843
rect 15882 14797 15928 14843
rect 15996 14797 16042 14843
rect 16110 14797 16156 14843
rect 16224 14797 16270 14843
rect 21337 14797 22097 14843
rect 22154 14797 22200 14843
rect 22257 14797 22303 14843
rect 22360 14797 22406 14843
rect 22463 14797 22509 14843
rect 22566 14797 22612 14843
rect 22669 14797 22715 14843
rect 22772 14797 22818 14843
rect 22875 14797 22921 14843
rect 22978 14797 23024 14843
rect 23081 14797 23127 14843
rect 23184 14797 23230 14843
rect 23287 14797 23333 14843
<< mvpdiffc >>
rect 640 15277 686 15323
rect 801 15277 847 15323
rect 961 15277 1007 15323
rect 1121 15277 1167 15323
rect 1282 15277 1328 15323
rect 1444 15277 1490 15323
rect 1607 15277 1653 15323
rect 6732 15245 8614 15291
rect 8671 15245 8717 15291
rect 8774 15245 8820 15291
rect 8877 15245 8923 15291
rect 8980 15245 9026 15291
rect 9083 15245 9129 15291
rect 9186 15245 9232 15291
rect 6732 15021 8614 15067
rect 8671 15021 8717 15067
rect 8774 15021 8820 15067
rect 8877 15021 8923 15067
rect 8980 15021 9026 15067
rect 9083 15021 9129 15067
rect 9186 15021 9232 15067
rect 9699 15021 9745 15067
rect 9802 15021 9848 15067
rect 9905 15021 9951 15067
rect 10009 15021 10055 15067
rect 10113 15021 10159 15067
rect 10217 15021 10263 15067
rect 10321 15021 10367 15067
rect 10425 15021 10471 15067
rect 10529 15021 10575 15067
rect 10633 15021 10679 15067
rect 10737 15021 10783 15067
rect 10841 15021 10887 15067
rect 10945 15021 10991 15067
rect 13999 15021 14045 15067
rect 14102 15021 14148 15067
rect 14205 15021 14251 15067
rect 14309 15021 14355 15067
rect 14413 15021 14459 15067
rect 14517 15021 14563 15067
rect 14621 15021 14667 15067
rect 14725 15021 14771 15067
rect 14829 15021 14875 15067
rect 14933 15021 14979 15067
rect 15037 15021 15083 15067
rect 15141 15021 15187 15067
rect 15245 15021 15291 15067
rect 18437 15245 20319 15291
rect 20376 15245 20422 15291
rect 20479 15245 20525 15291
rect 20582 15245 20628 15291
rect 20685 15245 20731 15291
rect 20788 15245 20834 15291
rect 20891 15245 20937 15291
rect 6732 14797 8614 14843
rect 8671 14797 8717 14843
rect 8774 14797 8820 14843
rect 8877 14797 8923 14843
rect 8980 14797 9026 14843
rect 9083 14797 9129 14843
rect 9186 14797 9232 14843
rect 9699 14797 9745 14843
rect 9802 14797 9848 14843
rect 9905 14797 9951 14843
rect 10009 14797 10055 14843
rect 10113 14797 10159 14843
rect 10217 14797 10263 14843
rect 10321 14797 10367 14843
rect 10425 14797 10471 14843
rect 10529 14797 10575 14843
rect 10633 14797 10679 14843
rect 10737 14797 10783 14843
rect 10841 14797 10887 14843
rect 10945 14797 10991 14843
rect 16669 15021 16715 15067
rect 16772 15021 16818 15067
rect 16875 15021 16921 15067
rect 16979 15021 17025 15067
rect 17083 15021 17129 15067
rect 17187 15021 17233 15067
rect 17291 15021 17337 15067
rect 17395 15021 17441 15067
rect 17499 15021 17545 15067
rect 17603 15021 17649 15067
rect 17707 15021 17753 15067
rect 17811 15021 17857 15067
rect 17915 15021 17961 15067
rect 18437 15021 20319 15067
rect 20376 15021 20422 15067
rect 20479 15021 20525 15067
rect 20582 15021 20628 15067
rect 20685 15021 20731 15067
rect 20788 15021 20834 15067
rect 20891 15021 20937 15067
rect 26116 15277 26162 15323
rect 26279 15277 26325 15323
rect 26441 15277 26487 15323
rect 26602 15277 26648 15323
rect 26762 15277 26808 15323
rect 26922 15277 26968 15323
rect 27083 15277 27129 15323
rect 13999 14797 14045 14843
rect 14102 14797 14148 14843
rect 14205 14797 14251 14843
rect 14309 14797 14355 14843
rect 14413 14797 14459 14843
rect 14517 14797 14563 14843
rect 14621 14797 14667 14843
rect 14725 14797 14771 14843
rect 14829 14797 14875 14843
rect 14933 14797 14979 14843
rect 15037 14797 15083 14843
rect 15141 14797 15187 14843
rect 15245 14797 15291 14843
rect 16669 14797 16715 14843
rect 16772 14797 16818 14843
rect 16875 14797 16921 14843
rect 16979 14797 17025 14843
rect 17083 14797 17129 14843
rect 17187 14797 17233 14843
rect 17291 14797 17337 14843
rect 17395 14797 17441 14843
rect 17499 14797 17545 14843
rect 17603 14797 17649 14843
rect 17707 14797 17753 14843
rect 17811 14797 17857 14843
rect 17915 14797 17961 14843
rect 18437 14797 20319 14843
rect 20376 14797 20422 14843
rect 20479 14797 20525 14843
rect 20582 14797 20628 14843
rect 20685 14797 20731 14843
rect 20788 14797 20834 14843
rect 20891 14797 20937 14843
rect 640 14377 686 14423
rect 801 14377 847 14423
rect 961 14377 1007 14423
rect 1121 14377 1167 14423
rect 1282 14377 1328 14423
rect 1444 14377 1490 14423
rect 1607 14377 1653 14423
rect 640 13477 686 13523
rect 801 13477 847 13523
rect 961 13477 1007 13523
rect 1121 13477 1167 13523
rect 1282 13477 1328 13523
rect 1444 13477 1490 13523
rect 1607 13477 1653 13523
rect 640 12577 686 12623
rect 801 12577 847 12623
rect 961 12577 1007 12623
rect 1121 12577 1167 12623
rect 1282 12577 1328 12623
rect 1444 12577 1490 12623
rect 1607 12577 1653 12623
rect 640 11677 686 11723
rect 801 11677 847 11723
rect 961 11677 1007 11723
rect 1121 11677 1167 11723
rect 1282 11677 1328 11723
rect 1444 11677 1490 11723
rect 1607 11677 1653 11723
rect 640 10777 686 10823
rect 801 10777 847 10823
rect 961 10777 1007 10823
rect 1121 10777 1167 10823
rect 1282 10777 1328 10823
rect 1444 10777 1490 10823
rect 1607 10777 1653 10823
rect 640 9877 686 9923
rect 801 9877 847 9923
rect 961 9877 1007 9923
rect 1121 9877 1167 9923
rect 1282 9877 1328 9923
rect 1444 9877 1490 9923
rect 1607 9877 1653 9923
rect 640 8977 686 9023
rect 801 8977 847 9023
rect 961 8977 1007 9023
rect 1121 8977 1167 9023
rect 1282 8977 1328 9023
rect 1444 8977 1490 9023
rect 1607 8977 1653 9023
rect 640 8077 686 8123
rect 801 8077 847 8123
rect 961 8077 1007 8123
rect 1121 8077 1167 8123
rect 1282 8077 1328 8123
rect 1444 8077 1490 8123
rect 1607 8077 1653 8123
rect 640 7177 686 7223
rect 801 7177 847 7223
rect 961 7177 1007 7223
rect 1121 7177 1167 7223
rect 1282 7177 1328 7223
rect 1444 7177 1490 7223
rect 1607 7177 1653 7223
rect 640 6277 686 6323
rect 801 6277 847 6323
rect 961 6277 1007 6323
rect 1121 6277 1167 6323
rect 1282 6277 1328 6323
rect 1444 6277 1490 6323
rect 1607 6277 1653 6323
rect 640 5377 686 5423
rect 801 5377 847 5423
rect 961 5377 1007 5423
rect 1121 5377 1167 5423
rect 1282 5377 1328 5423
rect 1444 5377 1490 5423
rect 1607 5377 1653 5423
rect 640 4477 686 4523
rect 801 4477 847 4523
rect 961 4477 1007 4523
rect 1121 4477 1167 4523
rect 1282 4477 1328 4523
rect 1444 4477 1490 4523
rect 1607 4477 1653 4523
rect 640 3577 686 3623
rect 801 3577 847 3623
rect 961 3577 1007 3623
rect 1121 3577 1167 3623
rect 1282 3577 1328 3623
rect 1444 3577 1490 3623
rect 1607 3577 1653 3623
rect 640 2677 686 2723
rect 801 2677 847 2723
rect 961 2677 1007 2723
rect 1121 2677 1167 2723
rect 1282 2677 1328 2723
rect 1444 2677 1490 2723
rect 1607 2677 1653 2723
rect 640 1777 686 1823
rect 801 1777 847 1823
rect 961 1777 1007 1823
rect 1121 1777 1167 1823
rect 1282 1777 1328 1823
rect 1444 1777 1490 1823
rect 1607 1777 1653 1823
rect 640 877 686 923
rect 801 877 847 923
rect 961 877 1007 923
rect 1121 877 1167 923
rect 1282 877 1328 923
rect 1444 877 1490 923
rect 1607 877 1653 923
rect 640 -23 686 23
rect 801 -23 847 23
rect 961 -23 1007 23
rect 1121 -23 1167 23
rect 1282 -23 1328 23
rect 1444 -23 1490 23
rect 1607 -23 1653 23
rect 26116 14377 26162 14423
rect 26279 14377 26325 14423
rect 26441 14377 26487 14423
rect 26602 14377 26648 14423
rect 26762 14377 26808 14423
rect 26922 14377 26968 14423
rect 27083 14377 27129 14423
rect 26116 13477 26162 13523
rect 26279 13477 26325 13523
rect 26441 13477 26487 13523
rect 26602 13477 26648 13523
rect 26762 13477 26808 13523
rect 26922 13477 26968 13523
rect 27083 13477 27129 13523
rect 26116 12577 26162 12623
rect 26279 12577 26325 12623
rect 26441 12577 26487 12623
rect 26602 12577 26648 12623
rect 26762 12577 26808 12623
rect 26922 12577 26968 12623
rect 27083 12577 27129 12623
rect 26116 11677 26162 11723
rect 26279 11677 26325 11723
rect 26441 11677 26487 11723
rect 26602 11677 26648 11723
rect 26762 11677 26808 11723
rect 26922 11677 26968 11723
rect 27083 11677 27129 11723
rect 26116 10777 26162 10823
rect 26279 10777 26325 10823
rect 26441 10777 26487 10823
rect 26602 10777 26648 10823
rect 26762 10777 26808 10823
rect 26922 10777 26968 10823
rect 27083 10777 27129 10823
rect 26116 9877 26162 9923
rect 26279 9877 26325 9923
rect 26441 9877 26487 9923
rect 26602 9877 26648 9923
rect 26762 9877 26808 9923
rect 26922 9877 26968 9923
rect 27083 9877 27129 9923
rect 26116 8977 26162 9023
rect 26279 8977 26325 9023
rect 26441 8977 26487 9023
rect 26602 8977 26648 9023
rect 26762 8977 26808 9023
rect 26922 8977 26968 9023
rect 27083 8977 27129 9023
rect 26116 8077 26162 8123
rect 26279 8077 26325 8123
rect 26441 8077 26487 8123
rect 26602 8077 26648 8123
rect 26762 8077 26808 8123
rect 26922 8077 26968 8123
rect 27083 8077 27129 8123
rect 26116 7177 26162 7223
rect 26279 7177 26325 7223
rect 26441 7177 26487 7223
rect 26602 7177 26648 7223
rect 26762 7177 26808 7223
rect 26922 7177 26968 7223
rect 27083 7177 27129 7223
rect 26116 6277 26162 6323
rect 26279 6277 26325 6323
rect 26441 6277 26487 6323
rect 26602 6277 26648 6323
rect 26762 6277 26808 6323
rect 26922 6277 26968 6323
rect 27083 6277 27129 6323
rect 26116 5377 26162 5423
rect 26279 5377 26325 5423
rect 26441 5377 26487 5423
rect 26602 5377 26648 5423
rect 26762 5377 26808 5423
rect 26922 5377 26968 5423
rect 27083 5377 27129 5423
rect 26116 4477 26162 4523
rect 26279 4477 26325 4523
rect 26441 4477 26487 4523
rect 26602 4477 26648 4523
rect 26762 4477 26808 4523
rect 26922 4477 26968 4523
rect 27083 4477 27129 4523
rect 26116 3577 26162 3623
rect 26279 3577 26325 3623
rect 26441 3577 26487 3623
rect 26602 3577 26648 3623
rect 26762 3577 26808 3623
rect 26922 3577 26968 3623
rect 27083 3577 27129 3623
rect 26116 2677 26162 2723
rect 26279 2677 26325 2723
rect 26441 2677 26487 2723
rect 26602 2677 26648 2723
rect 26762 2677 26808 2723
rect 26922 2677 26968 2723
rect 27083 2677 27129 2723
rect 26116 1777 26162 1823
rect 26279 1777 26325 1823
rect 26441 1777 26487 1823
rect 26602 1777 26648 1823
rect 26762 1777 26808 1823
rect 26922 1777 26968 1823
rect 27083 1777 27129 1823
rect 26116 877 26162 923
rect 26279 877 26325 923
rect 26441 877 26487 923
rect 26602 877 26648 923
rect 26762 877 26808 923
rect 26922 877 26968 923
rect 27083 877 27129 923
rect 26116 -23 26162 23
rect 26279 -23 26325 23
rect 26441 -23 26487 23
rect 26602 -23 26648 23
rect 26762 -23 26808 23
rect 26922 -23 26968 23
rect 27083 -23 27129 23
<< mvpsubdiff >>
rect 79 15195 234 15401
rect 4312 15382 6207 15439
rect 4312 15336 4367 15382
rect 4413 15336 4525 15382
rect 4571 15336 4683 15382
rect 4729 15336 4841 15382
rect 4887 15336 5000 15382
rect 5046 15336 5158 15382
rect 5204 15336 5316 15382
rect 5362 15336 5474 15382
rect 5520 15336 5632 15382
rect 5678 15336 5790 15382
rect 5836 15336 5948 15382
rect 5994 15336 6106 15382
rect 6152 15336 6207 15382
rect 4312 15279 6207 15336
rect 11385 15382 13280 15439
rect 11385 15336 11440 15382
rect 11486 15336 11598 15382
rect 11644 15336 11756 15382
rect 11802 15336 11914 15382
rect 11960 15336 12073 15382
rect 12119 15336 12231 15382
rect 12277 15336 12389 15382
rect 12435 15336 12547 15382
rect 12593 15336 12705 15382
rect 12751 15336 12863 15382
rect 12909 15336 13021 15382
rect 13067 15336 13179 15382
rect 13225 15336 13280 15382
rect 79 15149 133 15195
rect 179 15149 234 15195
rect 79 15031 234 15149
rect 79 14985 133 15031
rect 179 14985 234 15031
rect 79 14868 234 14985
rect 79 14822 133 14868
rect 179 14822 234 14868
rect 79 14705 234 14822
rect 79 14659 133 14705
rect 179 14659 234 14705
rect 79 14541 234 14659
rect 79 14495 133 14541
rect 179 14495 234 14541
rect 79 14339 234 14495
rect 11385 15279 13280 15336
rect 15782 15382 16254 15439
rect 15782 15336 15837 15382
rect 15883 15336 15995 15382
rect 16041 15336 16153 15382
rect 16199 15336 16254 15382
rect 15782 15279 16254 15336
rect 21397 15382 23292 15439
rect 21397 15336 21452 15382
rect 21498 15336 21610 15382
rect 21656 15336 21768 15382
rect 21814 15336 21926 15382
rect 21972 15336 22085 15382
rect 22131 15336 22243 15382
rect 22289 15336 22401 15382
rect 22447 15336 22559 15382
rect 22605 15336 22717 15382
rect 22763 15336 22875 15382
rect 22921 15336 23033 15382
rect 23079 15336 23191 15382
rect 23237 15336 23292 15382
rect 21397 15279 23292 15336
rect 79 14293 133 14339
rect 179 14293 234 14339
rect 79 14176 234 14293
rect 79 14130 133 14176
rect 179 14130 234 14176
rect 79 14013 234 14130
rect 79 13967 133 14013
rect 179 13967 234 14013
rect 79 13850 234 13967
rect 79 13804 133 13850
rect 179 13804 234 13850
rect 79 13686 234 13804
rect 79 13640 133 13686
rect 179 13640 234 13686
rect 79 13523 234 13640
rect 79 13477 133 13523
rect 179 13477 234 13523
rect 79 13360 234 13477
rect 79 13314 133 13360
rect 179 13314 234 13360
rect 79 13196 234 13314
rect 79 13150 133 13196
rect 179 13150 234 13196
rect 79 13033 234 13150
rect 79 12987 133 13033
rect 179 12987 234 13033
rect 79 12870 234 12987
rect 79 12824 133 12870
rect 179 12824 234 12870
rect 79 12707 234 12824
rect 79 12661 133 12707
rect 179 12661 234 12707
rect 79 12539 234 12661
rect 79 12493 133 12539
rect 179 12493 234 12539
rect 79 12376 234 12493
rect 79 12330 133 12376
rect 179 12330 234 12376
rect 79 12213 234 12330
rect 79 12167 133 12213
rect 179 12167 234 12213
rect 79 12050 234 12167
rect 79 12004 133 12050
rect 179 12004 234 12050
rect 79 11886 234 12004
rect 79 11840 133 11886
rect 179 11840 234 11886
rect 79 11723 234 11840
rect 79 11677 133 11723
rect 179 11677 234 11723
rect 79 11560 234 11677
rect 79 11514 133 11560
rect 179 11514 234 11560
rect 79 11396 234 11514
rect 79 11350 133 11396
rect 179 11350 234 11396
rect 79 11233 234 11350
rect 79 11187 133 11233
rect 179 11187 234 11233
rect 79 11070 234 11187
rect 79 11024 133 11070
rect 179 11024 234 11070
rect 79 10907 234 11024
rect 79 10861 133 10907
rect 179 10861 234 10907
rect 79 10739 234 10861
rect 79 10693 133 10739
rect 179 10693 234 10739
rect 79 10576 234 10693
rect 79 10530 133 10576
rect 179 10530 234 10576
rect 79 10413 234 10530
rect 79 10367 133 10413
rect 179 10367 234 10413
rect 79 10250 234 10367
rect 79 10204 133 10250
rect 179 10204 234 10250
rect 79 10086 234 10204
rect 79 10040 133 10086
rect 179 10040 234 10086
rect 79 9923 234 10040
rect 79 9877 133 9923
rect 179 9877 234 9923
rect 79 9760 234 9877
rect 79 9714 133 9760
rect 179 9714 234 9760
rect 79 9596 234 9714
rect 79 9550 133 9596
rect 179 9550 234 9596
rect 79 9433 234 9550
rect 79 9387 133 9433
rect 179 9387 234 9433
rect 79 9270 234 9387
rect 79 9224 133 9270
rect 179 9224 234 9270
rect 79 9107 234 9224
rect 79 9061 133 9107
rect 179 9061 234 9107
rect 79 8939 234 9061
rect 79 8893 133 8939
rect 179 8893 234 8939
rect 79 8776 234 8893
rect 79 8730 133 8776
rect 179 8730 234 8776
rect 79 8613 234 8730
rect 79 8567 133 8613
rect 179 8567 234 8613
rect 79 8450 234 8567
rect 79 8404 133 8450
rect 179 8404 234 8450
rect 79 8286 234 8404
rect 79 8240 133 8286
rect 179 8240 234 8286
rect 79 8123 234 8240
rect 79 8077 133 8123
rect 179 8077 234 8123
rect 79 7960 234 8077
rect 79 7914 133 7960
rect 179 7914 234 7960
rect 79 7796 234 7914
rect 79 7750 133 7796
rect 179 7750 234 7796
rect 79 7633 234 7750
rect 79 7587 133 7633
rect 179 7587 234 7633
rect 79 7470 234 7587
rect 79 7424 133 7470
rect 179 7424 234 7470
rect 79 7307 234 7424
rect 79 7261 133 7307
rect 179 7261 234 7307
rect 79 7139 234 7261
rect 79 7093 133 7139
rect 179 7093 234 7139
rect 79 6976 234 7093
rect 79 6930 133 6976
rect 179 6930 234 6976
rect 79 6813 234 6930
rect 79 6767 133 6813
rect 179 6767 234 6813
rect 79 6650 234 6767
rect 79 6604 133 6650
rect 179 6604 234 6650
rect 79 6486 234 6604
rect 79 6440 133 6486
rect 179 6440 234 6486
rect 79 6323 234 6440
rect 79 6277 133 6323
rect 179 6277 234 6323
rect 79 6160 234 6277
rect 79 6114 133 6160
rect 179 6114 234 6160
rect 79 5996 234 6114
rect 79 5950 133 5996
rect 179 5950 234 5996
rect 79 5833 234 5950
rect 79 5787 133 5833
rect 179 5787 234 5833
rect 79 5670 234 5787
rect 79 5624 133 5670
rect 179 5624 234 5670
rect 79 5507 234 5624
rect 79 5461 133 5507
rect 179 5461 234 5507
rect 79 5339 234 5461
rect 79 5293 133 5339
rect 179 5293 234 5339
rect 79 5176 234 5293
rect 79 5130 133 5176
rect 179 5130 234 5176
rect 79 5013 234 5130
rect 79 4967 133 5013
rect 179 4967 234 5013
rect 79 4850 234 4967
rect 79 4804 133 4850
rect 179 4804 234 4850
rect 79 4686 234 4804
rect 79 4640 133 4686
rect 179 4640 234 4686
rect 79 4523 234 4640
rect 79 4477 133 4523
rect 179 4477 234 4523
rect 79 4360 234 4477
rect 79 4314 133 4360
rect 179 4314 234 4360
rect 79 4196 234 4314
rect 79 4150 133 4196
rect 179 4150 234 4196
rect 79 4033 234 4150
rect 79 3987 133 4033
rect 179 3987 234 4033
rect 79 3870 234 3987
rect 79 3824 133 3870
rect 179 3824 234 3870
rect 79 3707 234 3824
rect 79 3661 133 3707
rect 179 3661 234 3707
rect 79 3539 234 3661
rect 79 3493 133 3539
rect 179 3493 234 3539
rect 79 3376 234 3493
rect 79 3330 133 3376
rect 179 3330 234 3376
rect 79 3213 234 3330
rect 79 3167 133 3213
rect 179 3167 234 3213
rect 79 3050 234 3167
rect 79 3004 133 3050
rect 179 3004 234 3050
rect 79 2886 234 3004
rect 79 2840 133 2886
rect 179 2840 234 2886
rect 79 2723 234 2840
rect 79 2677 133 2723
rect 179 2677 234 2723
rect 79 2560 234 2677
rect 79 2514 133 2560
rect 179 2514 234 2560
rect 79 2396 234 2514
rect 79 2350 133 2396
rect 179 2350 234 2396
rect 79 2233 234 2350
rect 79 2187 133 2233
rect 179 2187 234 2233
rect 79 2070 234 2187
rect 79 2024 133 2070
rect 179 2024 234 2070
rect 79 1907 234 2024
rect 79 1861 133 1907
rect 179 1861 234 1907
rect 79 1739 234 1861
rect 79 1693 133 1739
rect 179 1693 234 1739
rect 79 1576 234 1693
rect 79 1530 133 1576
rect 179 1530 234 1576
rect 79 1413 234 1530
rect 79 1367 133 1413
rect 179 1367 234 1413
rect 79 1250 234 1367
rect 79 1204 133 1250
rect 179 1204 234 1250
rect 79 1086 234 1204
rect 79 1040 133 1086
rect 179 1040 234 1086
rect 79 923 234 1040
rect 79 877 133 923
rect 179 877 234 923
rect 79 760 234 877
rect 79 714 133 760
rect 179 714 234 760
rect 79 596 234 714
rect 79 550 133 596
rect 179 550 234 596
rect 79 433 234 550
rect 79 387 133 433
rect 179 387 234 433
rect 79 270 234 387
rect 79 224 133 270
rect 179 224 234 270
rect 79 107 234 224
rect 79 61 133 107
rect 179 61 234 107
rect 79 -100 234 61
rect 27535 15195 27690 15401
rect 27535 15149 27590 15195
rect 27636 15149 27690 15195
rect 27535 15031 27690 15149
rect 27535 14985 27590 15031
rect 27636 14985 27690 15031
rect 27535 14868 27690 14985
rect 27535 14822 27590 14868
rect 27636 14822 27690 14868
rect 27535 14705 27690 14822
rect 27535 14659 27590 14705
rect 27636 14659 27690 14705
rect 27535 14541 27690 14659
rect 27535 14495 27590 14541
rect 27636 14495 27690 14541
rect 27535 14339 27690 14495
rect 27535 14293 27590 14339
rect 27636 14293 27690 14339
rect 27535 14176 27690 14293
rect 27535 14130 27590 14176
rect 27636 14130 27690 14176
rect 27535 14013 27690 14130
rect 27535 13967 27590 14013
rect 27636 13967 27690 14013
rect 27535 13850 27690 13967
rect 27535 13804 27590 13850
rect 27636 13804 27690 13850
rect 27535 13686 27690 13804
rect 27535 13640 27590 13686
rect 27636 13640 27690 13686
rect 27535 13523 27690 13640
rect 27535 13477 27590 13523
rect 27636 13477 27690 13523
rect 27535 13360 27690 13477
rect 27535 13314 27590 13360
rect 27636 13314 27690 13360
rect 27535 13196 27690 13314
rect 27535 13150 27590 13196
rect 27636 13150 27690 13196
rect 27535 13033 27690 13150
rect 27535 12987 27590 13033
rect 27636 12987 27690 13033
rect 27535 12870 27690 12987
rect 27535 12824 27590 12870
rect 27636 12824 27690 12870
rect 27535 12707 27690 12824
rect 27535 12661 27590 12707
rect 27636 12661 27690 12707
rect 27535 12539 27690 12661
rect 27535 12493 27590 12539
rect 27636 12493 27690 12539
rect 27535 12376 27690 12493
rect 27535 12330 27590 12376
rect 27636 12330 27690 12376
rect 27535 12213 27690 12330
rect 27535 12167 27590 12213
rect 27636 12167 27690 12213
rect 27535 12050 27690 12167
rect 27535 12004 27590 12050
rect 27636 12004 27690 12050
rect 27535 11886 27690 12004
rect 27535 11840 27590 11886
rect 27636 11840 27690 11886
rect 27535 11723 27690 11840
rect 27535 11677 27590 11723
rect 27636 11677 27690 11723
rect 27535 11560 27690 11677
rect 27535 11514 27590 11560
rect 27636 11514 27690 11560
rect 27535 11396 27690 11514
rect 27535 11350 27590 11396
rect 27636 11350 27690 11396
rect 27535 11233 27690 11350
rect 27535 11187 27590 11233
rect 27636 11187 27690 11233
rect 27535 11070 27690 11187
rect 27535 11024 27590 11070
rect 27636 11024 27690 11070
rect 27535 10907 27690 11024
rect 27535 10861 27590 10907
rect 27636 10861 27690 10907
rect 27535 10739 27690 10861
rect 27535 10693 27590 10739
rect 27636 10693 27690 10739
rect 27535 10576 27690 10693
rect 27535 10530 27590 10576
rect 27636 10530 27690 10576
rect 27535 10413 27690 10530
rect 27535 10367 27590 10413
rect 27636 10367 27690 10413
rect 27535 10250 27690 10367
rect 27535 10204 27590 10250
rect 27636 10204 27690 10250
rect 27535 10086 27690 10204
rect 27535 10040 27590 10086
rect 27636 10040 27690 10086
rect 27535 9923 27690 10040
rect 27535 9877 27590 9923
rect 27636 9877 27690 9923
rect 27535 9760 27690 9877
rect 27535 9714 27590 9760
rect 27636 9714 27690 9760
rect 27535 9596 27690 9714
rect 27535 9550 27590 9596
rect 27636 9550 27690 9596
rect 27535 9433 27690 9550
rect 27535 9387 27590 9433
rect 27636 9387 27690 9433
rect 27535 9270 27690 9387
rect 27535 9224 27590 9270
rect 27636 9224 27690 9270
rect 27535 9107 27690 9224
rect 27535 9061 27590 9107
rect 27636 9061 27690 9107
rect 27535 8939 27690 9061
rect 27535 8893 27590 8939
rect 27636 8893 27690 8939
rect 27535 8776 27690 8893
rect 27535 8730 27590 8776
rect 27636 8730 27690 8776
rect 27535 8613 27690 8730
rect 27535 8567 27590 8613
rect 27636 8567 27690 8613
rect 27535 8450 27690 8567
rect 27535 8404 27590 8450
rect 27636 8404 27690 8450
rect 27535 8286 27690 8404
rect 27535 8240 27590 8286
rect 27636 8240 27690 8286
rect 27535 8123 27690 8240
rect 27535 8077 27590 8123
rect 27636 8077 27690 8123
rect 27535 7960 27690 8077
rect 27535 7914 27590 7960
rect 27636 7914 27690 7960
rect 27535 7796 27690 7914
rect 27535 7750 27590 7796
rect 27636 7750 27690 7796
rect 27535 7633 27690 7750
rect 27535 7587 27590 7633
rect 27636 7587 27690 7633
rect 27535 7470 27690 7587
rect 27535 7424 27590 7470
rect 27636 7424 27690 7470
rect 27535 7307 27690 7424
rect 27535 7261 27590 7307
rect 27636 7261 27690 7307
rect 27535 7139 27690 7261
rect 27535 7093 27590 7139
rect 27636 7093 27690 7139
rect 27535 6976 27690 7093
rect 27535 6930 27590 6976
rect 27636 6930 27690 6976
rect 27535 6813 27690 6930
rect 27535 6767 27590 6813
rect 27636 6767 27690 6813
rect 27535 6650 27690 6767
rect 27535 6604 27590 6650
rect 27636 6604 27690 6650
rect 27535 6486 27690 6604
rect 27535 6440 27590 6486
rect 27636 6440 27690 6486
rect 27535 6323 27690 6440
rect 27535 6277 27590 6323
rect 27636 6277 27690 6323
rect 27535 6160 27690 6277
rect 27535 6114 27590 6160
rect 27636 6114 27690 6160
rect 27535 5996 27690 6114
rect 27535 5950 27590 5996
rect 27636 5950 27690 5996
rect 27535 5833 27690 5950
rect 27535 5787 27590 5833
rect 27636 5787 27690 5833
rect 27535 5670 27690 5787
rect 27535 5624 27590 5670
rect 27636 5624 27690 5670
rect 27535 5507 27690 5624
rect 27535 5461 27590 5507
rect 27636 5461 27690 5507
rect 27535 5339 27690 5461
rect 27535 5293 27590 5339
rect 27636 5293 27690 5339
rect 27535 5176 27690 5293
rect 27535 5130 27590 5176
rect 27636 5130 27690 5176
rect 27535 5013 27690 5130
rect 27535 4967 27590 5013
rect 27636 4967 27690 5013
rect 27535 4850 27690 4967
rect 27535 4804 27590 4850
rect 27636 4804 27690 4850
rect 27535 4686 27690 4804
rect 27535 4640 27590 4686
rect 27636 4640 27690 4686
rect 27535 4523 27690 4640
rect 27535 4477 27590 4523
rect 27636 4477 27690 4523
rect 27535 4360 27690 4477
rect 27535 4314 27590 4360
rect 27636 4314 27690 4360
rect 27535 4196 27690 4314
rect 27535 4150 27590 4196
rect 27636 4150 27690 4196
rect 27535 4033 27690 4150
rect 27535 3987 27590 4033
rect 27636 3987 27690 4033
rect 27535 3870 27690 3987
rect 27535 3824 27590 3870
rect 27636 3824 27690 3870
rect 27535 3707 27690 3824
rect 27535 3661 27590 3707
rect 27636 3661 27690 3707
rect 27535 3539 27690 3661
rect 27535 3493 27590 3539
rect 27636 3493 27690 3539
rect 27535 3376 27690 3493
rect 27535 3330 27590 3376
rect 27636 3330 27690 3376
rect 27535 3213 27690 3330
rect 27535 3167 27590 3213
rect 27636 3167 27690 3213
rect 27535 3050 27690 3167
rect 27535 3004 27590 3050
rect 27636 3004 27690 3050
rect 27535 2886 27690 3004
rect 27535 2840 27590 2886
rect 27636 2840 27690 2886
rect 27535 2723 27690 2840
rect 27535 2677 27590 2723
rect 27636 2677 27690 2723
rect 27535 2560 27690 2677
rect 27535 2514 27590 2560
rect 27636 2514 27690 2560
rect 27535 2396 27690 2514
rect 27535 2350 27590 2396
rect 27636 2350 27690 2396
rect 27535 2233 27690 2350
rect 27535 2187 27590 2233
rect 27636 2187 27690 2233
rect 27535 2070 27690 2187
rect 27535 2024 27590 2070
rect 27636 2024 27690 2070
rect 27535 1907 27690 2024
rect 27535 1861 27590 1907
rect 27636 1861 27690 1907
rect 27535 1739 27690 1861
rect 27535 1693 27590 1739
rect 27636 1693 27690 1739
rect 27535 1576 27690 1693
rect 27535 1530 27590 1576
rect 27636 1530 27690 1576
rect 27535 1413 27690 1530
rect 27535 1367 27590 1413
rect 27636 1367 27690 1413
rect 27535 1250 27690 1367
rect 27535 1204 27590 1250
rect 27636 1204 27690 1250
rect 27535 1086 27690 1204
rect 27535 1040 27590 1086
rect 27636 1040 27690 1086
rect 27535 923 27690 1040
rect 27535 877 27590 923
rect 27636 877 27690 923
rect 27535 760 27690 877
rect 27535 714 27590 760
rect 27636 714 27690 760
rect 27535 596 27690 714
rect 27535 550 27590 596
rect 27636 550 27690 596
rect 27535 433 27690 550
rect 27535 387 27590 433
rect 27636 387 27690 433
rect 27535 270 27690 387
rect 27535 224 27590 270
rect 27636 224 27690 270
rect 27535 107 27690 224
rect 27535 61 27590 107
rect 27636 61 27690 107
rect 27535 -100 27690 61
<< mvnsubdiff >>
rect 1906 15366 2125 15367
rect 1906 15309 4017 15366
rect 1906 15263 2177 15309
rect 2223 15263 2335 15309
rect 2381 15263 2493 15309
rect 2539 15263 2651 15309
rect 2697 15263 2810 15309
rect 2856 15263 2968 15309
rect 3014 15263 3126 15309
rect 3172 15263 3284 15309
rect 3330 15263 3442 15309
rect 3488 15263 3600 15309
rect 3646 15263 3758 15309
rect 3804 15263 3916 15309
rect 3962 15263 4017 15309
rect 1906 15195 4017 15263
rect 13985 15382 14931 15439
rect 13985 15336 14040 15382
rect 14086 15336 14198 15382
rect 14244 15336 14356 15382
rect 14402 15336 14514 15382
rect 14560 15336 14673 15382
rect 14719 15336 14831 15382
rect 14877 15336 14931 15382
rect 13985 15279 14931 15336
rect 1906 15149 1960 15195
rect 2006 15149 4017 15195
rect 1906 15146 4017 15149
rect 1906 15100 2177 15146
rect 2223 15100 2335 15146
rect 2381 15100 2493 15146
rect 2539 15100 2651 15146
rect 2697 15100 2810 15146
rect 2856 15100 2968 15146
rect 3014 15100 3126 15146
rect 3172 15100 3284 15146
rect 3330 15100 3442 15146
rect 3488 15100 3600 15146
rect 3646 15100 3758 15146
rect 3804 15100 3916 15146
rect 3962 15100 4017 15146
rect 1906 15031 4017 15100
rect 1906 14985 1960 15031
rect 2006 14985 4017 15031
rect 1906 14982 4017 14985
rect 1906 14936 2177 14982
rect 2223 14936 2335 14982
rect 2381 14936 2493 14982
rect 2539 14936 2651 14982
rect 2697 14936 2810 14982
rect 2856 14936 2968 14982
rect 3014 14936 3126 14982
rect 3172 14936 3284 14982
rect 3330 14936 3442 14982
rect 3488 14936 3600 14982
rect 3646 14936 3758 14982
rect 3804 14936 3916 14982
rect 3962 14936 4017 14982
rect 1906 14868 4017 14936
rect 25644 15366 25863 15367
rect 23751 15309 25863 15366
rect 23751 15263 23806 15309
rect 23852 15263 23964 15309
rect 24010 15263 24122 15309
rect 24168 15263 24280 15309
rect 24326 15263 24438 15309
rect 24484 15263 24596 15309
rect 24642 15263 24754 15309
rect 24800 15263 24912 15309
rect 24958 15263 25071 15309
rect 25117 15263 25229 15309
rect 25275 15263 25387 15309
rect 25433 15263 25545 15309
rect 25591 15263 25863 15309
rect 1906 14822 1960 14868
rect 2006 14822 4017 14868
rect 1906 14819 4017 14822
rect 1906 14773 2177 14819
rect 2223 14773 2335 14819
rect 2381 14773 2493 14819
rect 2539 14773 2651 14819
rect 2697 14773 2810 14819
rect 2856 14773 2968 14819
rect 3014 14773 3126 14819
rect 3172 14773 3284 14819
rect 3330 14773 3442 14819
rect 3488 14773 3600 14819
rect 3646 14773 3758 14819
rect 3804 14773 3916 14819
rect 3962 14773 4017 14819
rect 23751 15195 25863 15263
rect 23751 15149 25763 15195
rect 25809 15149 25863 15195
rect 23751 15146 25863 15149
rect 23751 15100 23806 15146
rect 23852 15100 23964 15146
rect 24010 15100 24122 15146
rect 24168 15100 24280 15146
rect 24326 15100 24438 15146
rect 24484 15100 24596 15146
rect 24642 15100 24754 15146
rect 24800 15100 24912 15146
rect 24958 15100 25071 15146
rect 25117 15100 25229 15146
rect 25275 15100 25387 15146
rect 25433 15100 25545 15146
rect 25591 15100 25863 15146
rect 23751 15031 25863 15100
rect 23751 14985 25763 15031
rect 25809 14985 25863 15031
rect 23751 14982 25863 14985
rect 23751 14936 23806 14982
rect 23852 14936 23964 14982
rect 24010 14936 24122 14982
rect 24168 14936 24280 14982
rect 24326 14936 24438 14982
rect 24484 14936 24596 14982
rect 24642 14936 24754 14982
rect 24800 14936 24912 14982
rect 24958 14936 25071 14982
rect 25117 14936 25229 14982
rect 25275 14936 25387 14982
rect 25433 14936 25545 14982
rect 25591 14936 25863 14982
rect 23751 14868 25863 14936
rect 23751 14822 25763 14868
rect 25809 14822 25863 14868
rect 23751 14819 25863 14822
rect 1906 14716 4017 14773
rect 23751 14773 23806 14819
rect 23852 14773 23964 14819
rect 24010 14773 24122 14819
rect 24168 14773 24280 14819
rect 24326 14773 24438 14819
rect 24484 14773 24596 14819
rect 24642 14773 24754 14819
rect 24800 14773 24912 14819
rect 24958 14773 25071 14819
rect 25117 14773 25229 14819
rect 25275 14773 25387 14819
rect 25433 14773 25545 14819
rect 25591 14773 25863 14819
rect 23751 14716 25863 14773
rect 1906 14705 2278 14716
rect 1906 14659 1960 14705
rect 2006 14659 2278 14705
rect 1906 14541 2278 14659
rect 1906 14495 1960 14541
rect 2006 14495 2278 14541
rect 1906 14460 2278 14495
rect 25490 14705 25863 14716
rect 25490 14659 25763 14705
rect 25809 14659 25863 14705
rect 25490 14541 25863 14659
rect 25490 14495 25763 14541
rect 25809 14495 25863 14541
rect 25490 14460 25863 14495
rect 1906 14339 2125 14460
rect 1906 14293 1960 14339
rect 2006 14293 2125 14339
rect 1906 14176 2125 14293
rect 1906 14130 1960 14176
rect 2006 14130 2125 14176
rect 1906 14013 2125 14130
rect 1906 13967 1960 14013
rect 2006 13967 2125 14013
rect 1906 13850 2125 13967
rect 1906 13804 1960 13850
rect 2006 13804 2125 13850
rect 1906 13686 2125 13804
rect 1906 13640 1960 13686
rect 2006 13640 2125 13686
rect 1906 13523 2125 13640
rect 1906 13477 1960 13523
rect 2006 13477 2125 13523
rect 1906 13360 2125 13477
rect 1906 13314 1960 13360
rect 2006 13314 2125 13360
rect 1906 13196 2125 13314
rect 1906 13150 1960 13196
rect 2006 13150 2125 13196
rect 1906 13033 2125 13150
rect 1906 12987 1960 13033
rect 2006 12987 2125 13033
rect 1906 12870 2125 12987
rect 1906 12824 1960 12870
rect 2006 12824 2125 12870
rect 1906 12707 2125 12824
rect 1906 12661 1960 12707
rect 2006 12661 2125 12707
rect 1906 12539 2125 12661
rect 1906 12493 1960 12539
rect 2006 12493 2125 12539
rect 1906 12376 2125 12493
rect 1906 12330 1960 12376
rect 2006 12330 2125 12376
rect 1906 12213 2125 12330
rect 1906 12167 1960 12213
rect 2006 12167 2125 12213
rect 1906 12050 2125 12167
rect 1906 12004 1960 12050
rect 2006 12004 2125 12050
rect 1906 11886 2125 12004
rect 1906 11840 1960 11886
rect 2006 11840 2125 11886
rect 1906 11723 2125 11840
rect 1906 11677 1960 11723
rect 2006 11677 2125 11723
rect 1906 11560 2125 11677
rect 1906 11514 1960 11560
rect 2006 11514 2125 11560
rect 1906 11396 2125 11514
rect 1906 11350 1960 11396
rect 2006 11350 2125 11396
rect 1906 11233 2125 11350
rect 1906 11187 1960 11233
rect 2006 11187 2125 11233
rect 1906 11070 2125 11187
rect 1906 11024 1960 11070
rect 2006 11024 2125 11070
rect 1906 10907 2125 11024
rect 1906 10861 1960 10907
rect 2006 10861 2125 10907
rect 1906 10739 2125 10861
rect 1906 10693 1960 10739
rect 2006 10693 2125 10739
rect 1906 10576 2125 10693
rect 1906 10530 1960 10576
rect 2006 10530 2125 10576
rect 1906 10413 2125 10530
rect 1906 10367 1960 10413
rect 2006 10367 2125 10413
rect 1906 10250 2125 10367
rect 1906 10204 1960 10250
rect 2006 10204 2125 10250
rect 1906 10086 2125 10204
rect 1906 10040 1960 10086
rect 2006 10040 2125 10086
rect 1906 9923 2125 10040
rect 1906 9877 1960 9923
rect 2006 9877 2125 9923
rect 1906 9760 2125 9877
rect 1906 9714 1960 9760
rect 2006 9714 2125 9760
rect 1906 9596 2125 9714
rect 1906 9550 1960 9596
rect 2006 9550 2125 9596
rect 1906 9433 2125 9550
rect 1906 9387 1960 9433
rect 2006 9387 2125 9433
rect 1906 9270 2125 9387
rect 1906 9224 1960 9270
rect 2006 9224 2125 9270
rect 1906 9107 2125 9224
rect 1906 9061 1960 9107
rect 2006 9061 2125 9107
rect 1906 8939 2125 9061
rect 1906 8893 1960 8939
rect 2006 8893 2125 8939
rect 1906 8776 2125 8893
rect 1906 8730 1960 8776
rect 2006 8730 2125 8776
rect 1906 8613 2125 8730
rect 1906 8567 1960 8613
rect 2006 8567 2125 8613
rect 1906 8450 2125 8567
rect 1906 8404 1960 8450
rect 2006 8404 2125 8450
rect 1906 8286 2125 8404
rect 1906 8240 1960 8286
rect 2006 8240 2125 8286
rect 1906 8123 2125 8240
rect 1906 8077 1960 8123
rect 2006 8077 2125 8123
rect 1906 7960 2125 8077
rect 1906 7914 1960 7960
rect 2006 7914 2125 7960
rect 1906 7796 2125 7914
rect 1906 7750 1960 7796
rect 2006 7750 2125 7796
rect 1906 7633 2125 7750
rect 1906 7587 1960 7633
rect 2006 7587 2125 7633
rect 1906 7470 2125 7587
rect 1906 7424 1960 7470
rect 2006 7424 2125 7470
rect 1906 7307 2125 7424
rect 1906 7261 1960 7307
rect 2006 7261 2125 7307
rect 1906 7139 2125 7261
rect 1906 7093 1960 7139
rect 2006 7093 2125 7139
rect 1906 6976 2125 7093
rect 1906 6930 1960 6976
rect 2006 6930 2125 6976
rect 1906 6813 2125 6930
rect 1906 6767 1960 6813
rect 2006 6767 2125 6813
rect 1906 6650 2125 6767
rect 1906 6604 1960 6650
rect 2006 6604 2125 6650
rect 1906 6486 2125 6604
rect 1906 6440 1960 6486
rect 2006 6440 2125 6486
rect 1906 6323 2125 6440
rect 1906 6277 1960 6323
rect 2006 6277 2125 6323
rect 1906 6160 2125 6277
rect 1906 6114 1960 6160
rect 2006 6114 2125 6160
rect 1906 5996 2125 6114
rect 1906 5950 1960 5996
rect 2006 5950 2125 5996
rect 1906 5833 2125 5950
rect 1906 5787 1960 5833
rect 2006 5787 2125 5833
rect 1906 5670 2125 5787
rect 1906 5624 1960 5670
rect 2006 5624 2125 5670
rect 1906 5507 2125 5624
rect 1906 5461 1960 5507
rect 2006 5461 2125 5507
rect 1906 5339 2125 5461
rect 1906 5293 1960 5339
rect 2006 5293 2125 5339
rect 1906 5176 2125 5293
rect 1906 5130 1960 5176
rect 2006 5130 2125 5176
rect 1906 5013 2125 5130
rect 1906 4967 1960 5013
rect 2006 4967 2125 5013
rect 1906 4850 2125 4967
rect 1906 4804 1960 4850
rect 2006 4804 2125 4850
rect 1906 4686 2125 4804
rect 1906 4640 1960 4686
rect 2006 4640 2125 4686
rect 1906 4523 2125 4640
rect 1906 4477 1960 4523
rect 2006 4477 2125 4523
rect 1906 4360 2125 4477
rect 1906 4314 1960 4360
rect 2006 4314 2125 4360
rect 1906 4196 2125 4314
rect 1906 4150 1960 4196
rect 2006 4150 2125 4196
rect 1906 4033 2125 4150
rect 1906 3987 1960 4033
rect 2006 3987 2125 4033
rect 1906 3870 2125 3987
rect 1906 3824 1960 3870
rect 2006 3824 2125 3870
rect 1906 3707 2125 3824
rect 1906 3661 1960 3707
rect 2006 3661 2125 3707
rect 1906 3539 2125 3661
rect 1906 3493 1960 3539
rect 2006 3493 2125 3539
rect 1906 3376 2125 3493
rect 1906 3330 1960 3376
rect 2006 3330 2125 3376
rect 1906 3213 2125 3330
rect 1906 3167 1960 3213
rect 2006 3167 2125 3213
rect 1906 3050 2125 3167
rect 1906 3004 1960 3050
rect 2006 3004 2125 3050
rect 1906 2886 2125 3004
rect 1906 2840 1960 2886
rect 2006 2840 2125 2886
rect 1906 2723 2125 2840
rect 1906 2677 1960 2723
rect 2006 2677 2125 2723
rect 1906 2560 2125 2677
rect 1906 2514 1960 2560
rect 2006 2514 2125 2560
rect 1906 2396 2125 2514
rect 1906 2350 1960 2396
rect 2006 2350 2125 2396
rect 1906 2233 2125 2350
rect 1906 2187 1960 2233
rect 2006 2187 2125 2233
rect 1906 2070 2125 2187
rect 1906 2024 1960 2070
rect 2006 2024 2125 2070
rect 1906 1907 2125 2024
rect 1906 1861 1960 1907
rect 2006 1861 2125 1907
rect 1906 1739 2125 1861
rect 1906 1693 1960 1739
rect 2006 1693 2125 1739
rect 1906 1576 2125 1693
rect 1906 1530 1960 1576
rect 2006 1530 2125 1576
rect 1906 1413 2125 1530
rect 1906 1367 1960 1413
rect 2006 1367 2125 1413
rect 1906 1250 2125 1367
rect 1906 1204 1960 1250
rect 2006 1204 2125 1250
rect 1906 1086 2125 1204
rect 1906 1040 1960 1086
rect 2006 1040 2125 1086
rect 1906 923 2125 1040
rect 1906 877 1960 923
rect 2006 877 2125 923
rect 1906 760 2125 877
rect 1906 714 1960 760
rect 2006 714 2125 760
rect 1906 596 2125 714
rect 1906 550 1960 596
rect 2006 550 2125 596
rect 1906 433 2125 550
rect 1906 387 1960 433
rect 2006 387 2125 433
rect 1906 270 2125 387
rect 1906 224 1960 270
rect 2006 224 2125 270
rect 1906 107 2125 224
rect 1906 61 1960 107
rect 2006 61 2125 107
rect 1906 -66 2125 61
rect 25644 14339 25863 14460
rect 25644 14293 25763 14339
rect 25809 14293 25863 14339
rect 25644 14176 25863 14293
rect 25644 14130 25763 14176
rect 25809 14130 25863 14176
rect 25644 14013 25863 14130
rect 25644 13967 25763 14013
rect 25809 13967 25863 14013
rect 25644 13850 25863 13967
rect 25644 13804 25763 13850
rect 25809 13804 25863 13850
rect 25644 13686 25863 13804
rect 25644 13640 25763 13686
rect 25809 13640 25863 13686
rect 25644 13523 25863 13640
rect 25644 13477 25763 13523
rect 25809 13477 25863 13523
rect 25644 13360 25863 13477
rect 25644 13314 25763 13360
rect 25809 13314 25863 13360
rect 25644 13196 25863 13314
rect 25644 13150 25763 13196
rect 25809 13150 25863 13196
rect 25644 13033 25863 13150
rect 25644 12987 25763 13033
rect 25809 12987 25863 13033
rect 25644 12870 25863 12987
rect 25644 12824 25763 12870
rect 25809 12824 25863 12870
rect 25644 12707 25863 12824
rect 25644 12661 25763 12707
rect 25809 12661 25863 12707
rect 25644 12539 25863 12661
rect 25644 12493 25763 12539
rect 25809 12493 25863 12539
rect 25644 12376 25863 12493
rect 25644 12330 25763 12376
rect 25809 12330 25863 12376
rect 25644 12213 25863 12330
rect 25644 12167 25763 12213
rect 25809 12167 25863 12213
rect 25644 12050 25863 12167
rect 25644 12004 25763 12050
rect 25809 12004 25863 12050
rect 25644 11886 25863 12004
rect 25644 11840 25763 11886
rect 25809 11840 25863 11886
rect 25644 11723 25863 11840
rect 25644 11677 25763 11723
rect 25809 11677 25863 11723
rect 25644 11560 25863 11677
rect 25644 11514 25763 11560
rect 25809 11514 25863 11560
rect 25644 11396 25863 11514
rect 25644 11350 25763 11396
rect 25809 11350 25863 11396
rect 25644 11233 25863 11350
rect 25644 11187 25763 11233
rect 25809 11187 25863 11233
rect 25644 11070 25863 11187
rect 25644 11024 25763 11070
rect 25809 11024 25863 11070
rect 25644 10907 25863 11024
rect 25644 10861 25763 10907
rect 25809 10861 25863 10907
rect 25644 10739 25863 10861
rect 25644 10693 25763 10739
rect 25809 10693 25863 10739
rect 25644 10576 25863 10693
rect 25644 10530 25763 10576
rect 25809 10530 25863 10576
rect 25644 10413 25863 10530
rect 25644 10367 25763 10413
rect 25809 10367 25863 10413
rect 25644 10250 25863 10367
rect 25644 10204 25763 10250
rect 25809 10204 25863 10250
rect 25644 10086 25863 10204
rect 25644 10040 25763 10086
rect 25809 10040 25863 10086
rect 25644 9923 25863 10040
rect 25644 9877 25763 9923
rect 25809 9877 25863 9923
rect 25644 9760 25863 9877
rect 25644 9714 25763 9760
rect 25809 9714 25863 9760
rect 25644 9596 25863 9714
rect 25644 9550 25763 9596
rect 25809 9550 25863 9596
rect 25644 9433 25863 9550
rect 25644 9387 25763 9433
rect 25809 9387 25863 9433
rect 25644 9270 25863 9387
rect 25644 9224 25763 9270
rect 25809 9224 25863 9270
rect 25644 9107 25863 9224
rect 25644 9061 25763 9107
rect 25809 9061 25863 9107
rect 25644 8939 25863 9061
rect 25644 8893 25763 8939
rect 25809 8893 25863 8939
rect 25644 8776 25863 8893
rect 25644 8730 25763 8776
rect 25809 8730 25863 8776
rect 25644 8613 25863 8730
rect 25644 8567 25763 8613
rect 25809 8567 25863 8613
rect 25644 8450 25863 8567
rect 25644 8404 25763 8450
rect 25809 8404 25863 8450
rect 25644 8286 25863 8404
rect 25644 8240 25763 8286
rect 25809 8240 25863 8286
rect 25644 8123 25863 8240
rect 25644 8077 25763 8123
rect 25809 8077 25863 8123
rect 25644 7960 25863 8077
rect 25644 7914 25763 7960
rect 25809 7914 25863 7960
rect 25644 7796 25863 7914
rect 25644 7750 25763 7796
rect 25809 7750 25863 7796
rect 25644 7633 25863 7750
rect 25644 7587 25763 7633
rect 25809 7587 25863 7633
rect 25644 7470 25863 7587
rect 25644 7424 25763 7470
rect 25809 7424 25863 7470
rect 25644 7307 25863 7424
rect 25644 7261 25763 7307
rect 25809 7261 25863 7307
rect 25644 7139 25863 7261
rect 25644 7093 25763 7139
rect 25809 7093 25863 7139
rect 25644 6976 25863 7093
rect 25644 6930 25763 6976
rect 25809 6930 25863 6976
rect 25644 6813 25863 6930
rect 25644 6767 25763 6813
rect 25809 6767 25863 6813
rect 25644 6650 25863 6767
rect 25644 6604 25763 6650
rect 25809 6604 25863 6650
rect 25644 6486 25863 6604
rect 25644 6440 25763 6486
rect 25809 6440 25863 6486
rect 25644 6323 25863 6440
rect 25644 6277 25763 6323
rect 25809 6277 25863 6323
rect 25644 6160 25863 6277
rect 25644 6114 25763 6160
rect 25809 6114 25863 6160
rect 25644 5996 25863 6114
rect 25644 5950 25763 5996
rect 25809 5950 25863 5996
rect 25644 5833 25863 5950
rect 25644 5787 25763 5833
rect 25809 5787 25863 5833
rect 25644 5670 25863 5787
rect 25644 5624 25763 5670
rect 25809 5624 25863 5670
rect 25644 5507 25863 5624
rect 25644 5461 25763 5507
rect 25809 5461 25863 5507
rect 25644 5339 25863 5461
rect 25644 5293 25763 5339
rect 25809 5293 25863 5339
rect 25644 5176 25863 5293
rect 25644 5130 25763 5176
rect 25809 5130 25863 5176
rect 25644 5013 25863 5130
rect 25644 4967 25763 5013
rect 25809 4967 25863 5013
rect 25644 4850 25863 4967
rect 25644 4804 25763 4850
rect 25809 4804 25863 4850
rect 25644 4686 25863 4804
rect 25644 4640 25763 4686
rect 25809 4640 25863 4686
rect 25644 4523 25863 4640
rect 25644 4477 25763 4523
rect 25809 4477 25863 4523
rect 25644 4360 25863 4477
rect 25644 4314 25763 4360
rect 25809 4314 25863 4360
rect 25644 4196 25863 4314
rect 25644 4150 25763 4196
rect 25809 4150 25863 4196
rect 25644 4033 25863 4150
rect 25644 3987 25763 4033
rect 25809 3987 25863 4033
rect 25644 3870 25863 3987
rect 25644 3824 25763 3870
rect 25809 3824 25863 3870
rect 25644 3707 25863 3824
rect 25644 3661 25763 3707
rect 25809 3661 25863 3707
rect 25644 3539 25863 3661
rect 25644 3493 25763 3539
rect 25809 3493 25863 3539
rect 25644 3376 25863 3493
rect 25644 3330 25763 3376
rect 25809 3330 25863 3376
rect 25644 3213 25863 3330
rect 25644 3167 25763 3213
rect 25809 3167 25863 3213
rect 25644 3050 25863 3167
rect 25644 3004 25763 3050
rect 25809 3004 25863 3050
rect 25644 2886 25863 3004
rect 25644 2840 25763 2886
rect 25809 2840 25863 2886
rect 25644 2723 25863 2840
rect 25644 2677 25763 2723
rect 25809 2677 25863 2723
rect 25644 2560 25863 2677
rect 25644 2514 25763 2560
rect 25809 2514 25863 2560
rect 25644 2396 25863 2514
rect 25644 2350 25763 2396
rect 25809 2350 25863 2396
rect 25644 2233 25863 2350
rect 25644 2187 25763 2233
rect 25809 2187 25863 2233
rect 25644 2070 25863 2187
rect 25644 2024 25763 2070
rect 25809 2024 25863 2070
rect 25644 1907 25863 2024
rect 25644 1861 25763 1907
rect 25809 1861 25863 1907
rect 25644 1739 25863 1861
rect 25644 1693 25763 1739
rect 25809 1693 25863 1739
rect 25644 1576 25863 1693
rect 25644 1530 25763 1576
rect 25809 1530 25863 1576
rect 25644 1413 25863 1530
rect 25644 1367 25763 1413
rect 25809 1367 25863 1413
rect 25644 1250 25863 1367
rect 25644 1204 25763 1250
rect 25809 1204 25863 1250
rect 25644 1086 25863 1204
rect 25644 1040 25763 1086
rect 25809 1040 25863 1086
rect 25644 923 25863 1040
rect 25644 877 25763 923
rect 25809 877 25863 923
rect 25644 760 25863 877
rect 25644 714 25763 760
rect 25809 714 25863 760
rect 25644 596 25863 714
rect 25644 550 25763 596
rect 25809 550 25863 596
rect 25644 433 25863 550
rect 25644 387 25763 433
rect 25809 387 25863 433
rect 25644 270 25863 387
rect 25644 224 25763 270
rect 25809 224 25863 270
rect 25644 107 25863 224
rect 25644 61 25763 107
rect 25809 61 25863 107
rect 25644 -66 25863 61
<< mvpsubdiffcont >>
rect 4367 15336 4413 15382
rect 4525 15336 4571 15382
rect 4683 15336 4729 15382
rect 4841 15336 4887 15382
rect 5000 15336 5046 15382
rect 5158 15336 5204 15382
rect 5316 15336 5362 15382
rect 5474 15336 5520 15382
rect 5632 15336 5678 15382
rect 5790 15336 5836 15382
rect 5948 15336 5994 15382
rect 6106 15336 6152 15382
rect 11440 15336 11486 15382
rect 11598 15336 11644 15382
rect 11756 15336 11802 15382
rect 11914 15336 11960 15382
rect 12073 15336 12119 15382
rect 12231 15336 12277 15382
rect 12389 15336 12435 15382
rect 12547 15336 12593 15382
rect 12705 15336 12751 15382
rect 12863 15336 12909 15382
rect 13021 15336 13067 15382
rect 13179 15336 13225 15382
rect 133 15149 179 15195
rect 133 14985 179 15031
rect 133 14822 179 14868
rect 133 14659 179 14705
rect 133 14495 179 14541
rect 15837 15336 15883 15382
rect 15995 15336 16041 15382
rect 16153 15336 16199 15382
rect 21452 15336 21498 15382
rect 21610 15336 21656 15382
rect 21768 15336 21814 15382
rect 21926 15336 21972 15382
rect 22085 15336 22131 15382
rect 22243 15336 22289 15382
rect 22401 15336 22447 15382
rect 22559 15336 22605 15382
rect 22717 15336 22763 15382
rect 22875 15336 22921 15382
rect 23033 15336 23079 15382
rect 23191 15336 23237 15382
rect 133 14293 179 14339
rect 133 14130 179 14176
rect 133 13967 179 14013
rect 133 13804 179 13850
rect 133 13640 179 13686
rect 133 13477 179 13523
rect 133 13314 179 13360
rect 133 13150 179 13196
rect 133 12987 179 13033
rect 133 12824 179 12870
rect 133 12661 179 12707
rect 133 12493 179 12539
rect 133 12330 179 12376
rect 133 12167 179 12213
rect 133 12004 179 12050
rect 133 11840 179 11886
rect 133 11677 179 11723
rect 133 11514 179 11560
rect 133 11350 179 11396
rect 133 11187 179 11233
rect 133 11024 179 11070
rect 133 10861 179 10907
rect 133 10693 179 10739
rect 133 10530 179 10576
rect 133 10367 179 10413
rect 133 10204 179 10250
rect 133 10040 179 10086
rect 133 9877 179 9923
rect 133 9714 179 9760
rect 133 9550 179 9596
rect 133 9387 179 9433
rect 133 9224 179 9270
rect 133 9061 179 9107
rect 133 8893 179 8939
rect 133 8730 179 8776
rect 133 8567 179 8613
rect 133 8404 179 8450
rect 133 8240 179 8286
rect 133 8077 179 8123
rect 133 7914 179 7960
rect 133 7750 179 7796
rect 133 7587 179 7633
rect 133 7424 179 7470
rect 133 7261 179 7307
rect 133 7093 179 7139
rect 133 6930 179 6976
rect 133 6767 179 6813
rect 133 6604 179 6650
rect 133 6440 179 6486
rect 133 6277 179 6323
rect 133 6114 179 6160
rect 133 5950 179 5996
rect 133 5787 179 5833
rect 133 5624 179 5670
rect 133 5461 179 5507
rect 133 5293 179 5339
rect 133 5130 179 5176
rect 133 4967 179 5013
rect 133 4804 179 4850
rect 133 4640 179 4686
rect 133 4477 179 4523
rect 133 4314 179 4360
rect 133 4150 179 4196
rect 133 3987 179 4033
rect 133 3824 179 3870
rect 133 3661 179 3707
rect 133 3493 179 3539
rect 133 3330 179 3376
rect 133 3167 179 3213
rect 133 3004 179 3050
rect 133 2840 179 2886
rect 133 2677 179 2723
rect 133 2514 179 2560
rect 133 2350 179 2396
rect 133 2187 179 2233
rect 133 2024 179 2070
rect 133 1861 179 1907
rect 133 1693 179 1739
rect 133 1530 179 1576
rect 133 1367 179 1413
rect 133 1204 179 1250
rect 133 1040 179 1086
rect 133 877 179 923
rect 133 714 179 760
rect 133 550 179 596
rect 133 387 179 433
rect 133 224 179 270
rect 133 61 179 107
rect 27590 15149 27636 15195
rect 27590 14985 27636 15031
rect 27590 14822 27636 14868
rect 27590 14659 27636 14705
rect 27590 14495 27636 14541
rect 27590 14293 27636 14339
rect 27590 14130 27636 14176
rect 27590 13967 27636 14013
rect 27590 13804 27636 13850
rect 27590 13640 27636 13686
rect 27590 13477 27636 13523
rect 27590 13314 27636 13360
rect 27590 13150 27636 13196
rect 27590 12987 27636 13033
rect 27590 12824 27636 12870
rect 27590 12661 27636 12707
rect 27590 12493 27636 12539
rect 27590 12330 27636 12376
rect 27590 12167 27636 12213
rect 27590 12004 27636 12050
rect 27590 11840 27636 11886
rect 27590 11677 27636 11723
rect 27590 11514 27636 11560
rect 27590 11350 27636 11396
rect 27590 11187 27636 11233
rect 27590 11024 27636 11070
rect 27590 10861 27636 10907
rect 27590 10693 27636 10739
rect 27590 10530 27636 10576
rect 27590 10367 27636 10413
rect 27590 10204 27636 10250
rect 27590 10040 27636 10086
rect 27590 9877 27636 9923
rect 27590 9714 27636 9760
rect 27590 9550 27636 9596
rect 27590 9387 27636 9433
rect 27590 9224 27636 9270
rect 27590 9061 27636 9107
rect 27590 8893 27636 8939
rect 27590 8730 27636 8776
rect 27590 8567 27636 8613
rect 27590 8404 27636 8450
rect 27590 8240 27636 8286
rect 27590 8077 27636 8123
rect 27590 7914 27636 7960
rect 27590 7750 27636 7796
rect 27590 7587 27636 7633
rect 27590 7424 27636 7470
rect 27590 7261 27636 7307
rect 27590 7093 27636 7139
rect 27590 6930 27636 6976
rect 27590 6767 27636 6813
rect 27590 6604 27636 6650
rect 27590 6440 27636 6486
rect 27590 6277 27636 6323
rect 27590 6114 27636 6160
rect 27590 5950 27636 5996
rect 27590 5787 27636 5833
rect 27590 5624 27636 5670
rect 27590 5461 27636 5507
rect 27590 5293 27636 5339
rect 27590 5130 27636 5176
rect 27590 4967 27636 5013
rect 27590 4804 27636 4850
rect 27590 4640 27636 4686
rect 27590 4477 27636 4523
rect 27590 4314 27636 4360
rect 27590 4150 27636 4196
rect 27590 3987 27636 4033
rect 27590 3824 27636 3870
rect 27590 3661 27636 3707
rect 27590 3493 27636 3539
rect 27590 3330 27636 3376
rect 27590 3167 27636 3213
rect 27590 3004 27636 3050
rect 27590 2840 27636 2886
rect 27590 2677 27636 2723
rect 27590 2514 27636 2560
rect 27590 2350 27636 2396
rect 27590 2187 27636 2233
rect 27590 2024 27636 2070
rect 27590 1861 27636 1907
rect 27590 1693 27636 1739
rect 27590 1530 27636 1576
rect 27590 1367 27636 1413
rect 27590 1204 27636 1250
rect 27590 1040 27636 1086
rect 27590 877 27636 923
rect 27590 714 27636 760
rect 27590 550 27636 596
rect 27590 387 27636 433
rect 27590 224 27636 270
rect 27590 61 27636 107
<< mvnsubdiffcont >>
rect 2177 15263 2223 15309
rect 2335 15263 2381 15309
rect 2493 15263 2539 15309
rect 2651 15263 2697 15309
rect 2810 15263 2856 15309
rect 2968 15263 3014 15309
rect 3126 15263 3172 15309
rect 3284 15263 3330 15309
rect 3442 15263 3488 15309
rect 3600 15263 3646 15309
rect 3758 15263 3804 15309
rect 3916 15263 3962 15309
rect 14040 15336 14086 15382
rect 14198 15336 14244 15382
rect 14356 15336 14402 15382
rect 14514 15336 14560 15382
rect 14673 15336 14719 15382
rect 14831 15336 14877 15382
rect 1960 15149 2006 15195
rect 2177 15100 2223 15146
rect 2335 15100 2381 15146
rect 2493 15100 2539 15146
rect 2651 15100 2697 15146
rect 2810 15100 2856 15146
rect 2968 15100 3014 15146
rect 3126 15100 3172 15146
rect 3284 15100 3330 15146
rect 3442 15100 3488 15146
rect 3600 15100 3646 15146
rect 3758 15100 3804 15146
rect 3916 15100 3962 15146
rect 1960 14985 2006 15031
rect 2177 14936 2223 14982
rect 2335 14936 2381 14982
rect 2493 14936 2539 14982
rect 2651 14936 2697 14982
rect 2810 14936 2856 14982
rect 2968 14936 3014 14982
rect 3126 14936 3172 14982
rect 3284 14936 3330 14982
rect 3442 14936 3488 14982
rect 3600 14936 3646 14982
rect 3758 14936 3804 14982
rect 3916 14936 3962 14982
rect 23806 15263 23852 15309
rect 23964 15263 24010 15309
rect 24122 15263 24168 15309
rect 24280 15263 24326 15309
rect 24438 15263 24484 15309
rect 24596 15263 24642 15309
rect 24754 15263 24800 15309
rect 24912 15263 24958 15309
rect 25071 15263 25117 15309
rect 25229 15263 25275 15309
rect 25387 15263 25433 15309
rect 25545 15263 25591 15309
rect 1960 14822 2006 14868
rect 2177 14773 2223 14819
rect 2335 14773 2381 14819
rect 2493 14773 2539 14819
rect 2651 14773 2697 14819
rect 2810 14773 2856 14819
rect 2968 14773 3014 14819
rect 3126 14773 3172 14819
rect 3284 14773 3330 14819
rect 3442 14773 3488 14819
rect 3600 14773 3646 14819
rect 3758 14773 3804 14819
rect 3916 14773 3962 14819
rect 25763 15149 25809 15195
rect 23806 15100 23852 15146
rect 23964 15100 24010 15146
rect 24122 15100 24168 15146
rect 24280 15100 24326 15146
rect 24438 15100 24484 15146
rect 24596 15100 24642 15146
rect 24754 15100 24800 15146
rect 24912 15100 24958 15146
rect 25071 15100 25117 15146
rect 25229 15100 25275 15146
rect 25387 15100 25433 15146
rect 25545 15100 25591 15146
rect 25763 14985 25809 15031
rect 23806 14936 23852 14982
rect 23964 14936 24010 14982
rect 24122 14936 24168 14982
rect 24280 14936 24326 14982
rect 24438 14936 24484 14982
rect 24596 14936 24642 14982
rect 24754 14936 24800 14982
rect 24912 14936 24958 14982
rect 25071 14936 25117 14982
rect 25229 14936 25275 14982
rect 25387 14936 25433 14982
rect 25545 14936 25591 14982
rect 25763 14822 25809 14868
rect 23806 14773 23852 14819
rect 23964 14773 24010 14819
rect 24122 14773 24168 14819
rect 24280 14773 24326 14819
rect 24438 14773 24484 14819
rect 24596 14773 24642 14819
rect 24754 14773 24800 14819
rect 24912 14773 24958 14819
rect 25071 14773 25117 14819
rect 25229 14773 25275 14819
rect 25387 14773 25433 14819
rect 25545 14773 25591 14819
rect 1960 14659 2006 14705
rect 1960 14495 2006 14541
rect 25763 14659 25809 14705
rect 25763 14495 25809 14541
rect 1960 14293 2006 14339
rect 1960 14130 2006 14176
rect 1960 13967 2006 14013
rect 1960 13804 2006 13850
rect 1960 13640 2006 13686
rect 1960 13477 2006 13523
rect 1960 13314 2006 13360
rect 1960 13150 2006 13196
rect 1960 12987 2006 13033
rect 1960 12824 2006 12870
rect 1960 12661 2006 12707
rect 1960 12493 2006 12539
rect 1960 12330 2006 12376
rect 1960 12167 2006 12213
rect 1960 12004 2006 12050
rect 1960 11840 2006 11886
rect 1960 11677 2006 11723
rect 1960 11514 2006 11560
rect 1960 11350 2006 11396
rect 1960 11187 2006 11233
rect 1960 11024 2006 11070
rect 1960 10861 2006 10907
rect 1960 10693 2006 10739
rect 1960 10530 2006 10576
rect 1960 10367 2006 10413
rect 1960 10204 2006 10250
rect 1960 10040 2006 10086
rect 1960 9877 2006 9923
rect 1960 9714 2006 9760
rect 1960 9550 2006 9596
rect 1960 9387 2006 9433
rect 1960 9224 2006 9270
rect 1960 9061 2006 9107
rect 1960 8893 2006 8939
rect 1960 8730 2006 8776
rect 1960 8567 2006 8613
rect 1960 8404 2006 8450
rect 1960 8240 2006 8286
rect 1960 8077 2006 8123
rect 1960 7914 2006 7960
rect 1960 7750 2006 7796
rect 1960 7587 2006 7633
rect 1960 7424 2006 7470
rect 1960 7261 2006 7307
rect 1960 7093 2006 7139
rect 1960 6930 2006 6976
rect 1960 6767 2006 6813
rect 1960 6604 2006 6650
rect 1960 6440 2006 6486
rect 1960 6277 2006 6323
rect 1960 6114 2006 6160
rect 1960 5950 2006 5996
rect 1960 5787 2006 5833
rect 1960 5624 2006 5670
rect 1960 5461 2006 5507
rect 1960 5293 2006 5339
rect 1960 5130 2006 5176
rect 1960 4967 2006 5013
rect 1960 4804 2006 4850
rect 1960 4640 2006 4686
rect 1960 4477 2006 4523
rect 1960 4314 2006 4360
rect 1960 4150 2006 4196
rect 1960 3987 2006 4033
rect 1960 3824 2006 3870
rect 1960 3661 2006 3707
rect 1960 3493 2006 3539
rect 1960 3330 2006 3376
rect 1960 3167 2006 3213
rect 1960 3004 2006 3050
rect 1960 2840 2006 2886
rect 1960 2677 2006 2723
rect 1960 2514 2006 2560
rect 1960 2350 2006 2396
rect 1960 2187 2006 2233
rect 1960 2024 2006 2070
rect 1960 1861 2006 1907
rect 1960 1693 2006 1739
rect 1960 1530 2006 1576
rect 1960 1367 2006 1413
rect 1960 1204 2006 1250
rect 1960 1040 2006 1086
rect 1960 877 2006 923
rect 1960 714 2006 760
rect 1960 550 2006 596
rect 1960 387 2006 433
rect 1960 224 2006 270
rect 1960 61 2006 107
rect 25763 14293 25809 14339
rect 25763 14130 25809 14176
rect 25763 13967 25809 14013
rect 25763 13804 25809 13850
rect 25763 13640 25809 13686
rect 25763 13477 25809 13523
rect 25763 13314 25809 13360
rect 25763 13150 25809 13196
rect 25763 12987 25809 13033
rect 25763 12824 25809 12870
rect 25763 12661 25809 12707
rect 25763 12493 25809 12539
rect 25763 12330 25809 12376
rect 25763 12167 25809 12213
rect 25763 12004 25809 12050
rect 25763 11840 25809 11886
rect 25763 11677 25809 11723
rect 25763 11514 25809 11560
rect 25763 11350 25809 11396
rect 25763 11187 25809 11233
rect 25763 11024 25809 11070
rect 25763 10861 25809 10907
rect 25763 10693 25809 10739
rect 25763 10530 25809 10576
rect 25763 10367 25809 10413
rect 25763 10204 25809 10250
rect 25763 10040 25809 10086
rect 25763 9877 25809 9923
rect 25763 9714 25809 9760
rect 25763 9550 25809 9596
rect 25763 9387 25809 9433
rect 25763 9224 25809 9270
rect 25763 9061 25809 9107
rect 25763 8893 25809 8939
rect 25763 8730 25809 8776
rect 25763 8567 25809 8613
rect 25763 8404 25809 8450
rect 25763 8240 25809 8286
rect 25763 8077 25809 8123
rect 25763 7914 25809 7960
rect 25763 7750 25809 7796
rect 25763 7587 25809 7633
rect 25763 7424 25809 7470
rect 25763 7261 25809 7307
rect 25763 7093 25809 7139
rect 25763 6930 25809 6976
rect 25763 6767 25809 6813
rect 25763 6604 25809 6650
rect 25763 6440 25809 6486
rect 25763 6277 25809 6323
rect 25763 6114 25809 6160
rect 25763 5950 25809 5996
rect 25763 5787 25809 5833
rect 25763 5624 25809 5670
rect 25763 5461 25809 5507
rect 25763 5293 25809 5339
rect 25763 5130 25809 5176
rect 25763 4967 25809 5013
rect 25763 4804 25809 4850
rect 25763 4640 25809 4686
rect 25763 4477 25809 4523
rect 25763 4314 25809 4360
rect 25763 4150 25809 4196
rect 25763 3987 25809 4033
rect 25763 3824 25809 3870
rect 25763 3661 25809 3707
rect 25763 3493 25809 3539
rect 25763 3330 25809 3376
rect 25763 3167 25809 3213
rect 25763 3004 25809 3050
rect 25763 2840 25809 2886
rect 25763 2677 25809 2723
rect 25763 2514 25809 2560
rect 25763 2350 25809 2396
rect 25763 2187 25809 2233
rect 25763 2024 25809 2070
rect 25763 1861 25809 1907
rect 25763 1693 25809 1739
rect 25763 1530 25809 1576
rect 25763 1367 25809 1413
rect 25763 1204 25809 1250
rect 25763 1040 25809 1086
rect 25763 877 25809 923
rect 25763 714 25809 760
rect 25763 550 25809 596
rect 25763 387 25809 433
rect 25763 224 25809 270
rect 25763 61 25809 107
<< polysilicon >>
rect 395 15117 597 15244
rect 395 15071 439 15117
rect 485 15071 597 15117
rect 395 14954 597 15071
rect 395 14908 439 14954
rect 485 14908 597 14954
rect 395 14790 597 14908
rect 395 14744 439 14790
rect 485 14744 597 14790
rect 395 14627 597 14744
rect 395 14581 439 14627
rect 485 14581 597 14627
rect 395 14456 597 14581
rect 1696 14456 1767 15244
rect 13623 15316 13801 15335
rect 13623 15270 13642 15316
rect 13782 15270 13801 15316
rect 15364 15364 15467 15383
rect 15364 15318 15390 15364
rect 15436 15318 15467 15364
rect 13623 15251 13801 15270
rect 9314 15216 9448 15223
rect 6556 15096 6719 15216
rect 9245 15118 9448 15216
rect 9245 15096 9358 15118
rect 6556 14992 6659 15096
rect 9314 14992 9358 15096
rect 4255 14872 4324 14992
rect 6346 14872 6719 14992
rect 9245 14978 9358 14992
rect 9404 14978 9448 15118
rect 11998 15031 12082 15050
rect 11998 14992 12017 15031
rect 9245 14873 9448 14978
rect 9245 14872 9316 14873
rect 9615 14872 9686 14992
rect 11004 14872 11385 14992
rect 11913 14891 12017 14992
rect 12063 14891 12082 15031
rect 13664 14993 13768 15251
rect 11913 14872 12082 14891
rect 12215 14873 12286 14993
rect 13604 14873 13768 14993
rect 15364 14992 15467 15318
rect 18271 15106 18424 15216
rect 13915 14872 13986 14992
rect 15304 14872 15467 14992
rect 15583 15071 15667 15090
rect 15583 14931 15602 15071
rect 15648 14992 15667 15071
rect 15648 14931 15755 14992
rect 15583 14872 15755 14931
rect 16283 14872 16656 14992
rect 17974 14872 18045 14992
rect 18271 14966 18290 15106
rect 18336 15096 18424 15106
rect 20950 15096 21113 15216
rect 18336 14992 18355 15096
rect 21010 14992 21113 15096
rect 18336 14966 18424 14992
rect 18271 14872 18424 14966
rect 20950 14872 21324 14992
rect 23346 14872 23417 14992
rect 395 14217 597 14344
rect 395 14171 439 14217
rect 485 14171 597 14217
rect 395 14054 597 14171
rect 395 14008 439 14054
rect 485 14008 597 14054
rect 395 13890 597 14008
rect 395 13844 439 13890
rect 485 13844 597 13890
rect 395 13727 597 13844
rect 395 13681 439 13727
rect 485 13681 597 13727
rect 395 13556 597 13681
rect 1696 13556 1767 14344
rect 395 13317 597 13444
rect 395 13271 439 13317
rect 485 13271 597 13317
rect 395 13154 597 13271
rect 395 13108 439 13154
rect 485 13108 597 13154
rect 395 12990 597 13108
rect 395 12944 439 12990
rect 485 12944 597 12990
rect 395 12827 597 12944
rect 395 12781 439 12827
rect 485 12781 597 12827
rect 395 12656 597 12781
rect 1696 12656 1767 13444
rect 395 12417 597 12544
rect 395 12371 439 12417
rect 485 12371 597 12417
rect 395 12254 597 12371
rect 395 12208 439 12254
rect 485 12208 597 12254
rect 395 12090 597 12208
rect 395 12044 439 12090
rect 485 12044 597 12090
rect 395 11927 597 12044
rect 395 11881 439 11927
rect 485 11881 597 11927
rect 395 11756 597 11881
rect 1696 11756 1767 12544
rect 395 11517 597 11644
rect 395 11471 439 11517
rect 485 11471 597 11517
rect 395 11354 597 11471
rect 395 11308 439 11354
rect 485 11308 597 11354
rect 395 11190 597 11308
rect 395 11144 439 11190
rect 485 11144 597 11190
rect 395 11027 597 11144
rect 395 10981 439 11027
rect 485 10981 597 11027
rect 395 10856 597 10981
rect 1696 10856 1767 11644
rect 395 10617 597 10744
rect 395 10571 439 10617
rect 485 10571 597 10617
rect 395 10454 597 10571
rect 395 10408 439 10454
rect 485 10408 597 10454
rect 395 10290 597 10408
rect 395 10244 439 10290
rect 485 10244 597 10290
rect 395 10127 597 10244
rect 395 10081 439 10127
rect 485 10081 597 10127
rect 395 9956 597 10081
rect 1696 9956 1767 10744
rect 395 9717 597 9844
rect 395 9671 439 9717
rect 485 9671 597 9717
rect 395 9554 597 9671
rect 395 9508 439 9554
rect 485 9508 597 9554
rect 395 9390 597 9508
rect 395 9344 439 9390
rect 485 9344 597 9390
rect 395 9227 597 9344
rect 395 9181 439 9227
rect 485 9181 597 9227
rect 395 9056 597 9181
rect 1696 9056 1767 9844
rect 395 8817 597 8944
rect 395 8771 439 8817
rect 485 8771 597 8817
rect 395 8654 597 8771
rect 395 8608 439 8654
rect 485 8608 597 8654
rect 395 8490 597 8608
rect 395 8444 439 8490
rect 485 8444 597 8490
rect 395 8327 597 8444
rect 395 8281 439 8327
rect 485 8281 597 8327
rect 395 8156 597 8281
rect 1696 8156 1767 8944
rect 395 7917 597 8044
rect 395 7871 439 7917
rect 485 7871 597 7917
rect 395 7754 597 7871
rect 395 7708 439 7754
rect 485 7708 597 7754
rect 395 7590 597 7708
rect 395 7544 439 7590
rect 485 7544 597 7590
rect 395 7427 597 7544
rect 395 7381 439 7427
rect 485 7381 597 7427
rect 395 7256 597 7381
rect 1696 7256 1767 8044
rect 395 7017 597 7144
rect 395 6971 439 7017
rect 485 6971 597 7017
rect 395 6854 597 6971
rect 395 6808 439 6854
rect 485 6808 597 6854
rect 395 6690 597 6808
rect 395 6644 439 6690
rect 485 6644 597 6690
rect 395 6527 597 6644
rect 395 6481 439 6527
rect 485 6481 597 6527
rect 395 6356 597 6481
rect 1696 6356 1767 7144
rect 395 6117 597 6244
rect 395 6071 439 6117
rect 485 6071 597 6117
rect 395 5954 597 6071
rect 395 5908 439 5954
rect 485 5908 597 5954
rect 395 5790 597 5908
rect 395 5744 439 5790
rect 485 5744 597 5790
rect 395 5627 597 5744
rect 395 5581 439 5627
rect 485 5581 597 5627
rect 395 5456 597 5581
rect 1696 5456 1767 6244
rect 395 5217 597 5344
rect 395 5171 439 5217
rect 485 5171 597 5217
rect 395 5054 597 5171
rect 395 5008 439 5054
rect 485 5008 597 5054
rect 395 4890 597 5008
rect 395 4844 439 4890
rect 485 4844 597 4890
rect 395 4727 597 4844
rect 395 4681 439 4727
rect 485 4681 597 4727
rect 395 4556 597 4681
rect 1696 4556 1767 5344
rect 395 4317 597 4444
rect 395 4271 439 4317
rect 485 4271 597 4317
rect 395 4154 597 4271
rect 395 4108 439 4154
rect 485 4108 597 4154
rect 395 3990 597 4108
rect 395 3944 439 3990
rect 485 3944 597 3990
rect 395 3827 597 3944
rect 395 3781 439 3827
rect 485 3781 597 3827
rect 395 3656 597 3781
rect 1696 3656 1767 4444
rect 395 3417 597 3544
rect 395 3371 439 3417
rect 485 3371 597 3417
rect 395 3254 597 3371
rect 395 3208 439 3254
rect 485 3208 597 3254
rect 395 3090 597 3208
rect 395 3044 439 3090
rect 485 3044 597 3090
rect 395 2927 597 3044
rect 395 2881 439 2927
rect 485 2881 597 2927
rect 395 2756 597 2881
rect 1696 2756 1767 3544
rect 395 2517 597 2644
rect 395 2471 439 2517
rect 485 2471 597 2517
rect 395 2354 597 2471
rect 395 2308 439 2354
rect 485 2308 597 2354
rect 395 2190 597 2308
rect 395 2144 439 2190
rect 485 2144 597 2190
rect 395 2027 597 2144
rect 395 1981 439 2027
rect 485 1981 597 2027
rect 395 1856 597 1981
rect 1696 1856 1767 2644
rect 395 1617 597 1744
rect 395 1571 439 1617
rect 485 1571 597 1617
rect 395 1454 597 1571
rect 395 1408 439 1454
rect 485 1408 597 1454
rect 395 1290 597 1408
rect 395 1244 439 1290
rect 485 1244 597 1290
rect 395 1127 597 1244
rect 395 1081 439 1127
rect 485 1081 597 1127
rect 395 956 597 1081
rect 1696 956 1767 1744
rect 395 717 597 844
rect 395 671 439 717
rect 485 671 597 717
rect 395 554 597 671
rect 395 508 439 554
rect 485 508 597 554
rect 395 390 597 508
rect 395 344 439 390
rect 485 344 597 390
rect 395 227 597 344
rect 395 181 439 227
rect 485 181 597 227
rect 395 56 597 181
rect 1696 56 1767 844
rect 26002 14456 26073 15244
rect 27172 15117 27374 15244
rect 27172 15071 27284 15117
rect 27330 15071 27374 15117
rect 27172 14954 27374 15071
rect 27172 14908 27284 14954
rect 27330 14908 27374 14954
rect 27172 14790 27374 14908
rect 27172 14744 27284 14790
rect 27330 14744 27374 14790
rect 27172 14627 27374 14744
rect 27172 14581 27284 14627
rect 27330 14581 27374 14627
rect 27172 14456 27374 14581
rect 26002 13556 26073 14344
rect 27172 14217 27374 14344
rect 27172 14171 27284 14217
rect 27330 14171 27374 14217
rect 27172 14054 27374 14171
rect 27172 14008 27284 14054
rect 27330 14008 27374 14054
rect 27172 13890 27374 14008
rect 27172 13844 27284 13890
rect 27330 13844 27374 13890
rect 27172 13727 27374 13844
rect 27172 13681 27284 13727
rect 27330 13681 27374 13727
rect 27172 13556 27374 13681
rect 26002 12656 26073 13444
rect 27172 13317 27374 13444
rect 27172 13271 27284 13317
rect 27330 13271 27374 13317
rect 27172 13154 27374 13271
rect 27172 13108 27284 13154
rect 27330 13108 27374 13154
rect 27172 12990 27374 13108
rect 27172 12944 27284 12990
rect 27330 12944 27374 12990
rect 27172 12827 27374 12944
rect 27172 12781 27284 12827
rect 27330 12781 27374 12827
rect 27172 12656 27374 12781
rect 26002 11756 26073 12544
rect 27172 12417 27374 12544
rect 27172 12371 27284 12417
rect 27330 12371 27374 12417
rect 27172 12254 27374 12371
rect 27172 12208 27284 12254
rect 27330 12208 27374 12254
rect 27172 12090 27374 12208
rect 27172 12044 27284 12090
rect 27330 12044 27374 12090
rect 27172 11927 27374 12044
rect 27172 11881 27284 11927
rect 27330 11881 27374 11927
rect 27172 11756 27374 11881
rect 26002 10856 26073 11644
rect 27172 11517 27374 11644
rect 27172 11471 27284 11517
rect 27330 11471 27374 11517
rect 27172 11354 27374 11471
rect 27172 11308 27284 11354
rect 27330 11308 27374 11354
rect 27172 11190 27374 11308
rect 27172 11144 27284 11190
rect 27330 11144 27374 11190
rect 27172 11027 27374 11144
rect 27172 10981 27284 11027
rect 27330 10981 27374 11027
rect 27172 10856 27374 10981
rect 26002 9956 26073 10744
rect 27172 10617 27374 10744
rect 27172 10571 27284 10617
rect 27330 10571 27374 10617
rect 27172 10454 27374 10571
rect 27172 10408 27284 10454
rect 27330 10408 27374 10454
rect 27172 10290 27374 10408
rect 27172 10244 27284 10290
rect 27330 10244 27374 10290
rect 27172 10127 27374 10244
rect 27172 10081 27284 10127
rect 27330 10081 27374 10127
rect 27172 9956 27374 10081
rect 26002 9056 26073 9844
rect 27172 9717 27374 9844
rect 27172 9671 27284 9717
rect 27330 9671 27374 9717
rect 27172 9554 27374 9671
rect 27172 9508 27284 9554
rect 27330 9508 27374 9554
rect 27172 9390 27374 9508
rect 27172 9344 27284 9390
rect 27330 9344 27374 9390
rect 27172 9227 27374 9344
rect 27172 9181 27284 9227
rect 27330 9181 27374 9227
rect 27172 9056 27374 9181
rect 26002 8156 26073 8944
rect 27172 8817 27374 8944
rect 27172 8771 27284 8817
rect 27330 8771 27374 8817
rect 27172 8654 27374 8771
rect 27172 8608 27284 8654
rect 27330 8608 27374 8654
rect 27172 8490 27374 8608
rect 27172 8444 27284 8490
rect 27330 8444 27374 8490
rect 27172 8327 27374 8444
rect 27172 8281 27284 8327
rect 27330 8281 27374 8327
rect 27172 8156 27374 8281
rect 26002 7256 26073 8044
rect 27172 7917 27374 8044
rect 27172 7871 27284 7917
rect 27330 7871 27374 7917
rect 27172 7754 27374 7871
rect 27172 7708 27284 7754
rect 27330 7708 27374 7754
rect 27172 7590 27374 7708
rect 27172 7544 27284 7590
rect 27330 7544 27374 7590
rect 27172 7427 27374 7544
rect 27172 7381 27284 7427
rect 27330 7381 27374 7427
rect 27172 7256 27374 7381
rect 26002 6356 26073 7144
rect 27172 7017 27374 7144
rect 27172 6971 27284 7017
rect 27330 6971 27374 7017
rect 27172 6854 27374 6971
rect 27172 6808 27284 6854
rect 27330 6808 27374 6854
rect 27172 6690 27374 6808
rect 27172 6644 27284 6690
rect 27330 6644 27374 6690
rect 27172 6527 27374 6644
rect 27172 6481 27284 6527
rect 27330 6481 27374 6527
rect 27172 6356 27374 6481
rect 26002 5456 26073 6244
rect 27172 6117 27374 6244
rect 27172 6071 27284 6117
rect 27330 6071 27374 6117
rect 27172 5954 27374 6071
rect 27172 5908 27284 5954
rect 27330 5908 27374 5954
rect 27172 5790 27374 5908
rect 27172 5744 27284 5790
rect 27330 5744 27374 5790
rect 27172 5627 27374 5744
rect 27172 5581 27284 5627
rect 27330 5581 27374 5627
rect 27172 5456 27374 5581
rect 26002 4556 26073 5344
rect 27172 5217 27374 5344
rect 27172 5171 27284 5217
rect 27330 5171 27374 5217
rect 27172 5054 27374 5171
rect 27172 5008 27284 5054
rect 27330 5008 27374 5054
rect 27172 4890 27374 5008
rect 27172 4844 27284 4890
rect 27330 4844 27374 4890
rect 27172 4727 27374 4844
rect 27172 4681 27284 4727
rect 27330 4681 27374 4727
rect 27172 4556 27374 4681
rect 26002 3656 26073 4444
rect 27172 4317 27374 4444
rect 27172 4271 27284 4317
rect 27330 4271 27374 4317
rect 27172 4154 27374 4271
rect 27172 4108 27284 4154
rect 27330 4108 27374 4154
rect 27172 3990 27374 4108
rect 27172 3944 27284 3990
rect 27330 3944 27374 3990
rect 27172 3827 27374 3944
rect 27172 3781 27284 3827
rect 27330 3781 27374 3827
rect 27172 3656 27374 3781
rect 26002 2756 26073 3544
rect 27172 3417 27374 3544
rect 27172 3371 27284 3417
rect 27330 3371 27374 3417
rect 27172 3254 27374 3371
rect 27172 3208 27284 3254
rect 27330 3208 27374 3254
rect 27172 3090 27374 3208
rect 27172 3044 27284 3090
rect 27330 3044 27374 3090
rect 27172 2927 27374 3044
rect 27172 2881 27284 2927
rect 27330 2881 27374 2927
rect 27172 2756 27374 2881
rect 26002 1856 26073 2644
rect 27172 2517 27374 2644
rect 27172 2471 27284 2517
rect 27330 2471 27374 2517
rect 27172 2354 27374 2471
rect 27172 2308 27284 2354
rect 27330 2308 27374 2354
rect 27172 2190 27374 2308
rect 27172 2144 27284 2190
rect 27330 2144 27374 2190
rect 27172 2027 27374 2144
rect 27172 1981 27284 2027
rect 27330 1981 27374 2027
rect 27172 1856 27374 1981
rect 26002 956 26073 1744
rect 27172 1617 27374 1744
rect 27172 1571 27284 1617
rect 27330 1571 27374 1617
rect 27172 1454 27374 1571
rect 27172 1408 27284 1454
rect 27330 1408 27374 1454
rect 27172 1290 27374 1408
rect 27172 1244 27284 1290
rect 27330 1244 27374 1290
rect 27172 1127 27374 1244
rect 27172 1081 27284 1127
rect 27330 1081 27374 1127
rect 27172 956 27374 1081
rect 26002 56 26073 844
rect 27172 717 27374 844
rect 27172 671 27284 717
rect 27330 671 27374 717
rect 27172 554 27374 671
rect 27172 508 27284 554
rect 27330 508 27374 554
rect 27172 390 27374 508
rect 27172 344 27284 390
rect 27330 344 27374 390
rect 27172 227 27374 344
rect 27172 181 27284 227
rect 27330 181 27374 227
rect 27172 56 27374 181
<< polycontact >>
rect 439 15071 485 15117
rect 439 14908 485 14954
rect 439 14744 485 14790
rect 439 14581 485 14627
rect 13642 15270 13782 15316
rect 15390 15318 15436 15364
rect 9358 14978 9404 15118
rect 12017 14891 12063 15031
rect 15602 14931 15648 15071
rect 18290 14966 18336 15106
rect 439 14171 485 14217
rect 439 14008 485 14054
rect 439 13844 485 13890
rect 439 13681 485 13727
rect 439 13271 485 13317
rect 439 13108 485 13154
rect 439 12944 485 12990
rect 439 12781 485 12827
rect 439 12371 485 12417
rect 439 12208 485 12254
rect 439 12044 485 12090
rect 439 11881 485 11927
rect 439 11471 485 11517
rect 439 11308 485 11354
rect 439 11144 485 11190
rect 439 10981 485 11027
rect 439 10571 485 10617
rect 439 10408 485 10454
rect 439 10244 485 10290
rect 439 10081 485 10127
rect 439 9671 485 9717
rect 439 9508 485 9554
rect 439 9344 485 9390
rect 439 9181 485 9227
rect 439 8771 485 8817
rect 439 8608 485 8654
rect 439 8444 485 8490
rect 439 8281 485 8327
rect 439 7871 485 7917
rect 439 7708 485 7754
rect 439 7544 485 7590
rect 439 7381 485 7427
rect 439 6971 485 7017
rect 439 6808 485 6854
rect 439 6644 485 6690
rect 439 6481 485 6527
rect 439 6071 485 6117
rect 439 5908 485 5954
rect 439 5744 485 5790
rect 439 5581 485 5627
rect 439 5171 485 5217
rect 439 5008 485 5054
rect 439 4844 485 4890
rect 439 4681 485 4727
rect 439 4271 485 4317
rect 439 4108 485 4154
rect 439 3944 485 3990
rect 439 3781 485 3827
rect 439 3371 485 3417
rect 439 3208 485 3254
rect 439 3044 485 3090
rect 439 2881 485 2927
rect 439 2471 485 2517
rect 439 2308 485 2354
rect 439 2144 485 2190
rect 439 1981 485 2027
rect 439 1571 485 1617
rect 439 1408 485 1454
rect 439 1244 485 1290
rect 439 1081 485 1127
rect 439 671 485 717
rect 439 508 485 554
rect 439 344 485 390
rect 439 181 485 227
rect 27284 15071 27330 15117
rect 27284 14908 27330 14954
rect 27284 14744 27330 14790
rect 27284 14581 27330 14627
rect 27284 14171 27330 14217
rect 27284 14008 27330 14054
rect 27284 13844 27330 13890
rect 27284 13681 27330 13727
rect 27284 13271 27330 13317
rect 27284 13108 27330 13154
rect 27284 12944 27330 12990
rect 27284 12781 27330 12827
rect 27284 12371 27330 12417
rect 27284 12208 27330 12254
rect 27284 12044 27330 12090
rect 27284 11881 27330 11927
rect 27284 11471 27330 11517
rect 27284 11308 27330 11354
rect 27284 11144 27330 11190
rect 27284 10981 27330 11027
rect 27284 10571 27330 10617
rect 27284 10408 27330 10454
rect 27284 10244 27330 10290
rect 27284 10081 27330 10127
rect 27284 9671 27330 9717
rect 27284 9508 27330 9554
rect 27284 9344 27330 9390
rect 27284 9181 27330 9227
rect 27284 8771 27330 8817
rect 27284 8608 27330 8654
rect 27284 8444 27330 8490
rect 27284 8281 27330 8327
rect 27284 7871 27330 7917
rect 27284 7708 27330 7754
rect 27284 7544 27330 7590
rect 27284 7381 27330 7427
rect 27284 6971 27330 7017
rect 27284 6808 27330 6854
rect 27284 6644 27330 6690
rect 27284 6481 27330 6527
rect 27284 6071 27330 6117
rect 27284 5908 27330 5954
rect 27284 5744 27330 5790
rect 27284 5581 27330 5627
rect 27284 5171 27330 5217
rect 27284 5008 27330 5054
rect 27284 4844 27330 4890
rect 27284 4681 27330 4727
rect 27284 4271 27330 4317
rect 27284 4108 27330 4154
rect 27284 3944 27330 3990
rect 27284 3781 27330 3827
rect 27284 3371 27330 3417
rect 27284 3208 27330 3254
rect 27284 3044 27330 3090
rect 27284 2881 27330 2927
rect 27284 2471 27330 2517
rect 27284 2308 27330 2354
rect 27284 2144 27330 2190
rect 27284 1981 27330 2027
rect 27284 1571 27330 1617
rect 27284 1408 27330 1454
rect 27284 1244 27330 1290
rect 27284 1081 27330 1127
rect 27284 671 27330 717
rect 27284 508 27330 554
rect 27284 344 27330 390
rect 27284 181 27330 227
<< metal1 >>
rect 79 15326 519 15401
rect 4324 15382 6336 15439
rect 79 15274 168 15326
rect 220 15274 379 15326
rect 431 15274 519 15326
rect 79 15195 519 15274
rect 606 15326 1688 15367
rect 606 15323 905 15326
rect 606 15277 640 15323
rect 686 15277 801 15323
rect 847 15277 905 15323
rect 606 15274 905 15277
rect 957 15323 1116 15326
rect 1168 15323 1328 15326
rect 957 15277 961 15323
rect 1007 15277 1116 15323
rect 1168 15277 1282 15323
rect 957 15274 1116 15277
rect 1168 15274 1328 15277
rect 1380 15323 1539 15326
rect 1380 15277 1444 15323
rect 1490 15277 1539 15323
rect 1380 15274 1539 15277
rect 1591 15323 1688 15326
rect 1591 15277 1607 15323
rect 1653 15277 1688 15323
rect 1591 15274 1688 15277
rect 606 15234 1688 15274
rect 1906 15326 4017 15367
rect 1906 15274 2130 15326
rect 2182 15309 2341 15326
rect 2393 15309 2552 15326
rect 1906 15263 2177 15274
rect 2223 15263 2335 15309
rect 2393 15274 2493 15309
rect 2381 15263 2493 15274
rect 2539 15274 2552 15309
rect 2604 15309 2763 15326
rect 2815 15309 2974 15326
rect 3026 15309 3184 15326
rect 2604 15274 2651 15309
rect 2539 15263 2651 15274
rect 2697 15274 2763 15309
rect 2697 15263 2810 15274
rect 2856 15263 2968 15309
rect 3026 15274 3126 15309
rect 3014 15263 3126 15274
rect 3172 15274 3184 15309
rect 3236 15309 3395 15326
rect 3447 15309 3606 15326
rect 3658 15309 3817 15326
rect 3236 15274 3284 15309
rect 3172 15263 3284 15274
rect 3330 15274 3395 15309
rect 3330 15263 3442 15274
rect 3488 15263 3600 15309
rect 3658 15274 3758 15309
rect 3646 15263 3758 15274
rect 3804 15274 3817 15309
rect 3869 15309 4017 15326
rect 3869 15274 3916 15309
rect 3804 15263 3916 15274
rect 3962 15263 4017 15309
rect 867 15233 1629 15234
rect 79 15149 133 15195
rect 179 15149 519 15195
rect 79 15117 519 15149
rect 79 15071 439 15117
rect 485 15071 519 15117
rect 79 15031 519 15071
rect 79 14985 133 15031
rect 179 14985 519 15031
rect 79 14954 519 14985
rect 79 14908 439 14954
rect 485 14908 519 14954
rect 79 14868 519 14908
rect 79 14822 133 14868
rect 179 14822 519 14868
rect 79 14790 519 14822
rect 79 14744 439 14790
rect 485 14744 519 14790
rect 79 14705 519 14744
rect 79 14659 133 14705
rect 179 14659 519 14705
rect 79 14627 519 14659
rect 79 14581 439 14627
rect 485 14581 519 14627
rect 79 14541 519 14581
rect 79 14495 133 14541
rect 179 14495 519 14541
rect 79 14339 519 14495
rect 1906 15195 4017 15263
rect 1906 15149 1960 15195
rect 2006 15149 4017 15195
rect 1906 15146 4017 15149
rect 1906 15108 2177 15146
rect 1906 15056 2130 15108
rect 2223 15100 2335 15146
rect 2381 15108 2493 15146
rect 2393 15100 2493 15108
rect 2539 15108 2651 15146
rect 2539 15100 2552 15108
rect 2182 15056 2341 15100
rect 2393 15056 2552 15100
rect 2604 15100 2651 15108
rect 2697 15108 2810 15146
rect 2697 15100 2763 15108
rect 2856 15100 2968 15146
rect 3014 15108 3126 15146
rect 3026 15100 3126 15108
rect 3172 15108 3284 15146
rect 3172 15100 3184 15108
rect 2604 15056 2763 15100
rect 2815 15056 2974 15100
rect 3026 15056 3184 15100
rect 3236 15100 3284 15108
rect 3330 15108 3442 15146
rect 3330 15100 3395 15108
rect 3488 15100 3600 15146
rect 3646 15108 3758 15146
rect 3658 15100 3758 15108
rect 3804 15108 3916 15146
rect 3804 15100 3817 15108
rect 3236 15056 3395 15100
rect 3447 15056 3606 15100
rect 3658 15056 3817 15100
rect 3869 15100 3916 15108
rect 3962 15100 4017 15146
rect 3869 15056 4017 15100
rect 1906 15031 4017 15056
rect 1906 14985 1960 15031
rect 2006 14985 4017 15031
rect 4324 15336 4367 15382
rect 4413 15336 4525 15382
rect 4571 15336 4683 15382
rect 4729 15336 4841 15382
rect 4887 15336 5000 15382
rect 5046 15336 5158 15382
rect 5204 15336 5316 15382
rect 5362 15336 5474 15382
rect 5520 15336 5632 15382
rect 5678 15336 5790 15382
rect 5836 15336 5948 15382
rect 5994 15336 6106 15382
rect 6152 15336 6336 15382
rect 11385 15382 13260 15419
rect 4324 15326 6336 15336
rect 4324 15274 5613 15326
rect 5665 15274 5824 15326
rect 5876 15274 6035 15326
rect 6087 15274 6246 15326
rect 6298 15274 6336 15326
rect 6728 15306 7700 15346
rect 6728 15291 6766 15306
rect 6818 15291 6977 15306
rect 7029 15291 7188 15306
rect 7240 15291 7399 15306
rect 7451 15291 7610 15306
rect 7662 15291 7700 15306
rect 11385 15336 11440 15382
rect 11486 15336 11598 15382
rect 11644 15336 11756 15382
rect 11802 15336 11914 15382
rect 11960 15336 12073 15382
rect 12119 15336 12231 15382
rect 12277 15336 12389 15382
rect 12435 15336 12547 15382
rect 12593 15336 12705 15382
rect 12751 15336 12863 15382
rect 12909 15336 13021 15382
rect 13067 15336 13179 15382
rect 13225 15336 13260 15382
rect 11385 15331 13260 15336
rect 4324 15108 6336 15274
rect 6719 15245 6732 15291
rect 8614 15245 8671 15291
rect 8717 15245 8774 15291
rect 8820 15245 8877 15291
rect 8923 15245 8980 15291
rect 9026 15245 9083 15291
rect 9129 15245 9186 15291
rect 9232 15245 9245 15291
rect 11385 15279 11575 15331
rect 11627 15279 11755 15331
rect 11807 15299 13260 15331
rect 13531 15382 14912 15419
rect 15755 15418 16283 15419
rect 13531 15378 14040 15382
rect 13531 15326 14033 15378
rect 14086 15336 14198 15382
rect 14244 15378 14356 15382
rect 14085 15326 14244 15336
rect 14296 15336 14356 15378
rect 14402 15378 14514 15382
rect 14402 15336 14455 15378
rect 14296 15326 14455 15336
rect 14507 15336 14514 15378
rect 14560 15336 14673 15382
rect 14719 15336 14831 15382
rect 14877 15336 14912 15382
rect 14507 15326 14912 15336
rect 13531 15317 14912 15326
rect 11807 15279 11913 15299
rect 6728 15214 7700 15245
rect 9323 15118 9439 15185
rect 4324 15067 5613 15108
rect 4324 15021 4337 15067
rect 5097 15021 5154 15067
rect 5200 15021 5257 15067
rect 5303 15021 5360 15067
rect 5406 15021 5463 15067
rect 5509 15021 5566 15067
rect 5612 15056 5613 15067
rect 5665 15067 5824 15108
rect 5876 15067 6035 15108
rect 6087 15067 6246 15108
rect 6298 15067 6336 15108
rect 6482 15067 6767 15108
rect 5665 15056 5669 15067
rect 5612 15021 5669 15056
rect 5715 15021 5772 15067
rect 5818 15056 5824 15067
rect 5818 15021 5875 15056
rect 5921 15021 5978 15067
rect 6024 15056 6035 15067
rect 6024 15021 6081 15056
rect 6127 15021 6184 15067
rect 6230 15056 6246 15067
rect 6230 15021 6287 15056
rect 6333 15021 6346 15067
rect 6482 15021 6732 15067
rect 8614 15021 8671 15067
rect 8717 15021 8774 15067
rect 8820 15021 8877 15067
rect 8923 15021 8980 15067
rect 9026 15021 9083 15067
rect 9129 15021 9186 15067
rect 9232 15021 9245 15067
rect 5574 15016 6336 15021
rect 1906 14982 4017 14985
rect 1906 14936 2177 14982
rect 2223 14936 2335 14982
rect 2381 14936 2493 14982
rect 2539 14936 2651 14982
rect 2697 14936 2810 14982
rect 2856 14936 2968 14982
rect 3014 14936 3126 14982
rect 3172 14936 3284 14982
rect 3330 14936 3442 14982
rect 3488 14936 3600 14982
rect 3646 14936 3758 14982
rect 3804 14936 3916 14982
rect 3962 14936 4017 14982
rect 1906 14891 4017 14936
rect 1906 14868 2130 14891
rect 1906 14822 1960 14868
rect 2006 14839 2130 14868
rect 2182 14839 2341 14891
rect 2393 14839 2552 14891
rect 2604 14839 2763 14891
rect 2815 14839 2974 14891
rect 3026 14839 3184 14891
rect 3236 14839 3395 14891
rect 3447 14839 3606 14891
rect 3658 14839 3817 14891
rect 3869 14839 4017 14891
rect 6482 14988 6767 15021
rect 4335 14845 5307 14885
rect 6482 14877 6598 14988
rect 9323 14978 9358 15118
rect 9404 14978 9439 15118
rect 10338 15108 10888 15115
rect 10337 15074 10888 15108
rect 10337 15067 10376 15074
rect 10428 15067 10587 15074
rect 10639 15067 10798 15074
rect 10850 15067 10888 15074
rect 11385 15113 11913 15279
rect 13531 15265 13569 15317
rect 13621 15316 13781 15317
rect 13621 15270 13642 15316
rect 13833 15299 14912 15317
rect 15061 15382 16283 15418
rect 15061 15378 15837 15382
rect 15061 15326 15100 15378
rect 15152 15326 15311 15378
rect 15363 15364 15522 15378
rect 15363 15326 15390 15364
rect 15061 15318 15390 15326
rect 15436 15326 15522 15364
rect 15574 15326 15733 15378
rect 15785 15336 15837 15378
rect 15883 15336 15995 15382
rect 16041 15336 16153 15382
rect 16199 15336 16283 15382
rect 21324 15382 23346 15419
rect 20112 15340 20874 15346
rect 15785 15326 16283 15336
rect 15436 15318 16283 15326
rect 13833 15286 14545 15299
rect 13833 15285 14040 15286
rect 15061 15285 16283 15318
rect 13621 15265 13781 15270
rect 13833 15265 13871 15285
rect 13531 15224 13871 15265
rect 11385 15067 11575 15113
rect 11627 15067 11755 15113
rect 11807 15067 11913 15113
rect 15591 15071 15659 15082
rect 9686 15021 9699 15067
rect 9745 15021 9802 15067
rect 9848 15021 9905 15067
rect 9951 15021 10009 15067
rect 10055 15021 10113 15067
rect 10159 15021 10217 15067
rect 10263 15021 10321 15067
rect 10367 15022 10376 15067
rect 10367 15021 10425 15022
rect 10471 15021 10529 15067
rect 10575 15022 10587 15067
rect 10575 15021 10633 15022
rect 10679 15021 10737 15067
rect 10783 15022 10798 15067
rect 10783 15021 10841 15022
rect 10887 15021 10945 15067
rect 10991 15021 11004 15067
rect 11385 15021 11398 15067
rect 11444 15021 11512 15067
rect 11558 15061 11575 15067
rect 11558 15021 11626 15061
rect 11672 15021 11740 15067
rect 11807 15061 11854 15067
rect 11786 15021 11854 15061
rect 11900 15021 11913 15067
rect 12006 15031 12299 15068
rect 10337 14988 10888 15021
rect 10338 14982 10888 14988
rect 4335 14843 4373 14845
rect 4425 14843 4584 14845
rect 4636 14843 4795 14845
rect 4847 14843 5006 14845
rect 5058 14843 5217 14845
rect 5269 14843 5307 14845
rect 6240 14843 6598 14877
rect 6728 14843 7700 14883
rect 9323 14877 9439 14978
rect 12006 14891 12017 15031
rect 12063 15022 12299 15031
rect 12345 15022 12402 15068
rect 12448 15022 12505 15068
rect 12551 15022 12609 15068
rect 12655 15022 12713 15068
rect 12759 15022 12817 15068
rect 12863 15022 12921 15068
rect 12967 15022 13025 15068
rect 13071 15022 13129 15068
rect 13175 15022 13233 15068
rect 13279 15022 13337 15068
rect 13383 15022 13441 15068
rect 13487 15022 13545 15068
rect 13591 15067 14174 15068
rect 15591 15067 15602 15071
rect 13591 15022 13999 15067
rect 12063 14891 12074 15022
rect 13986 15021 13999 15022
rect 14045 15021 14102 15067
rect 14148 15021 14205 15067
rect 14251 15021 14309 15067
rect 14355 15021 14413 15067
rect 14459 15021 14517 15067
rect 14563 15021 14621 15067
rect 14667 15021 14725 15067
rect 14771 15021 14829 15067
rect 14875 15021 14933 15067
rect 14979 15021 15037 15067
rect 15083 15021 15141 15067
rect 15187 15021 15245 15067
rect 15291 15021 15602 15067
rect 15591 14931 15602 15021
rect 15648 14931 15659 15071
rect 15755 15067 16283 15285
rect 15755 15021 15768 15067
rect 15814 15021 15882 15067
rect 15928 15021 15996 15067
rect 16042 15021 16110 15067
rect 16156 15021 16224 15067
rect 16270 15021 16283 15067
rect 16656 15306 20942 15340
rect 16656 15291 20151 15306
rect 20203 15291 20362 15306
rect 20414 15291 20573 15306
rect 20625 15291 20784 15306
rect 20836 15291 20942 15306
rect 21324 15336 21452 15382
rect 21498 15336 21610 15382
rect 21656 15336 21768 15382
rect 21814 15336 21926 15382
rect 21972 15336 22085 15382
rect 22131 15336 22243 15382
rect 22289 15336 22401 15382
rect 22447 15336 22559 15382
rect 22605 15336 22717 15382
rect 22763 15336 22875 15382
rect 22921 15336 23033 15382
rect 23079 15336 23191 15382
rect 23237 15336 23346 15382
rect 21324 15326 23346 15336
rect 16656 15245 18437 15291
rect 20319 15254 20362 15291
rect 20319 15245 20376 15254
rect 20422 15245 20479 15291
rect 20525 15254 20573 15291
rect 20525 15245 20582 15254
rect 20628 15245 20685 15291
rect 20731 15254 20784 15291
rect 20836 15254 20891 15291
rect 20731 15245 20788 15254
rect 20834 15245 20891 15254
rect 20937 15245 20950 15291
rect 21324 15274 21460 15326
rect 21512 15274 21671 15326
rect 21723 15274 21882 15326
rect 21934 15274 22093 15326
rect 22145 15274 23346 15326
rect 16656 15220 20942 15245
rect 16656 15067 17974 15220
rect 20112 15213 20874 15220
rect 16656 15021 16669 15067
rect 16715 15021 16772 15067
rect 16818 15021 16875 15067
rect 16921 15021 16979 15067
rect 17025 15021 17083 15067
rect 17129 15021 17187 15067
rect 17233 15021 17291 15067
rect 17337 15021 17395 15067
rect 17441 15021 17499 15067
rect 17545 15021 17603 15067
rect 17649 15021 17707 15067
rect 17753 15021 17811 15067
rect 17857 15021 17915 15067
rect 17961 15021 17974 15067
rect 18279 15106 18347 15117
rect 15755 14988 16283 15021
rect 15591 14920 15659 14931
rect 18279 14966 18290 15106
rect 18336 14966 18347 15106
rect 21324 15108 23346 15274
rect 21324 15067 21460 15108
rect 21512 15067 21671 15108
rect 21723 15067 21882 15108
rect 21934 15067 22093 15108
rect 22145 15067 23346 15108
rect 18424 15021 18437 15067
rect 20319 15021 20376 15067
rect 20422 15021 20479 15067
rect 20525 15021 20582 15067
rect 20628 15021 20685 15067
rect 20731 15021 20788 15067
rect 20834 15021 20891 15067
rect 20937 15021 21184 15067
rect 18279 14955 18347 14966
rect 12006 14880 12074 14891
rect 9323 14843 11913 14877
rect 12294 14844 13478 14884
rect 18279 14877 18346 14955
rect 2006 14822 4017 14839
rect 1906 14819 4017 14822
rect 1906 14773 2177 14819
rect 2223 14773 2335 14819
rect 2381 14773 2493 14819
rect 2539 14773 2651 14819
rect 2697 14773 2810 14819
rect 2856 14773 2968 14819
rect 3014 14773 3126 14819
rect 3172 14773 3284 14819
rect 3330 14773 3442 14819
rect 3488 14773 3600 14819
rect 3646 14773 3758 14819
rect 3804 14773 3916 14819
rect 3962 14773 4017 14819
rect 4324 14797 4337 14843
rect 5097 14797 5154 14843
rect 5200 14797 5217 14843
rect 5303 14797 5360 14843
rect 5406 14797 5463 14843
rect 5509 14797 5566 14843
rect 5612 14797 5669 14843
rect 5715 14797 5772 14843
rect 5818 14797 5875 14843
rect 5921 14797 5978 14843
rect 6024 14797 6081 14843
rect 6127 14797 6184 14843
rect 6230 14797 6287 14843
rect 6333 14797 6598 14843
rect 6719 14797 6732 14843
rect 8614 14797 8671 14843
rect 8717 14797 8774 14843
rect 8820 14797 8877 14843
rect 8923 14797 8980 14843
rect 9026 14797 9083 14843
rect 9129 14797 9186 14843
rect 9232 14797 9245 14843
rect 9323 14797 9699 14843
rect 9745 14797 9802 14843
rect 9848 14797 9905 14843
rect 9951 14797 10009 14843
rect 10055 14797 10113 14843
rect 10159 14797 10217 14843
rect 10263 14797 10321 14843
rect 10367 14797 10425 14843
rect 10471 14797 10529 14843
rect 10575 14797 10633 14843
rect 10679 14797 10737 14843
rect 10783 14797 10841 14843
rect 10887 14797 10945 14843
rect 10991 14797 11398 14843
rect 11444 14797 11512 14843
rect 11558 14797 11626 14843
rect 11672 14797 11740 14843
rect 11786 14797 11854 14843
rect 11900 14797 11913 14843
rect 12286 14798 12299 14844
rect 12345 14843 12402 14844
rect 12385 14798 12402 14843
rect 12448 14798 12505 14844
rect 12551 14843 12609 14844
rect 12596 14798 12609 14843
rect 12655 14798 12713 14844
rect 12759 14843 12817 14844
rect 12807 14798 12817 14843
rect 12863 14798 12921 14844
rect 12967 14843 13025 14844
rect 13018 14798 13025 14843
rect 13071 14798 13129 14844
rect 13175 14843 13233 14844
rect 13175 14798 13177 14843
rect 1906 14716 4017 14773
rect 4335 14793 4373 14797
rect 4425 14793 4584 14797
rect 4636 14793 4795 14797
rect 4847 14793 5006 14797
rect 5058 14793 5217 14797
rect 5269 14793 5307 14797
rect 4335 14753 5307 14793
rect 6240 14757 6598 14797
rect 6728 14791 6766 14797
rect 6818 14791 6977 14797
rect 7029 14791 7188 14797
rect 7240 14791 7399 14797
rect 7451 14791 7610 14797
rect 7662 14791 7700 14797
rect 6728 14751 7700 14791
rect 9323 14757 11913 14797
rect 12294 14791 12333 14798
rect 12385 14791 12544 14798
rect 12596 14791 12755 14798
rect 12807 14791 12966 14798
rect 13018 14791 13177 14798
rect 13229 14798 13233 14843
rect 13279 14798 13337 14844
rect 13383 14843 13441 14844
rect 13383 14798 13387 14843
rect 13229 14791 13387 14798
rect 13439 14798 13441 14843
rect 13487 14798 13545 14844
rect 13591 14843 14174 14844
rect 15755 14843 18346 14877
rect 20112 14843 20874 14883
rect 21067 14843 21184 15021
rect 21324 15021 21337 15067
rect 22145 15056 22154 15067
rect 22097 15021 22154 15056
rect 22200 15021 22257 15067
rect 22303 15021 22360 15067
rect 22406 15021 22463 15067
rect 22509 15021 22566 15067
rect 22612 15021 22669 15067
rect 22715 15021 22772 15067
rect 22818 15021 22875 15067
rect 22921 15021 22978 15067
rect 23024 15021 23081 15067
rect 23127 15021 23184 15067
rect 23230 15021 23287 15067
rect 23333 15021 23346 15067
rect 21324 15002 23346 15021
rect 23751 15326 25863 15367
rect 23751 15309 23899 15326
rect 23751 15263 23806 15309
rect 23852 15274 23899 15309
rect 23951 15309 24110 15326
rect 24162 15309 24321 15326
rect 24373 15309 24532 15326
rect 23951 15274 23964 15309
rect 23852 15263 23964 15274
rect 24010 15274 24110 15309
rect 24010 15263 24122 15274
rect 24168 15263 24280 15309
rect 24373 15274 24438 15309
rect 24326 15263 24438 15274
rect 24484 15274 24532 15309
rect 24584 15309 24742 15326
rect 24794 15309 24953 15326
rect 25005 15309 25164 15326
rect 24584 15274 24596 15309
rect 24484 15263 24596 15274
rect 24642 15274 24742 15309
rect 24642 15263 24754 15274
rect 24800 15263 24912 15309
rect 25005 15274 25071 15309
rect 24958 15263 25071 15274
rect 25117 15274 25164 15309
rect 25216 15309 25375 15326
rect 25427 15309 25586 15326
rect 25216 15274 25229 15309
rect 25117 15263 25229 15274
rect 25275 15274 25375 15309
rect 25275 15263 25387 15274
rect 25433 15263 25545 15309
rect 25638 15274 25863 15326
rect 25591 15263 25863 15274
rect 23751 15195 25863 15263
rect 26081 15326 27163 15367
rect 26081 15323 26178 15326
rect 26081 15277 26116 15323
rect 26162 15277 26178 15323
rect 26081 15274 26178 15277
rect 26230 15323 26389 15326
rect 26230 15277 26279 15323
rect 26325 15277 26389 15323
rect 26230 15274 26389 15277
rect 26441 15323 26601 15326
rect 26653 15323 26812 15326
rect 26487 15277 26601 15323
rect 26653 15277 26762 15323
rect 26808 15277 26812 15323
rect 26441 15274 26601 15277
rect 26653 15274 26812 15277
rect 26864 15323 27163 15326
rect 26864 15277 26922 15323
rect 26968 15277 27083 15323
rect 27129 15277 27163 15323
rect 26864 15274 27163 15277
rect 26081 15234 27163 15274
rect 27250 15326 27690 15401
rect 27250 15274 27338 15326
rect 27390 15274 27549 15326
rect 27601 15274 27690 15326
rect 26140 15233 26902 15234
rect 23751 15149 25763 15195
rect 25809 15149 25863 15195
rect 23751 15146 25863 15149
rect 23751 15100 23806 15146
rect 23852 15108 23964 15146
rect 23852 15100 23899 15108
rect 23751 15056 23899 15100
rect 23951 15100 23964 15108
rect 24010 15108 24122 15146
rect 24010 15100 24110 15108
rect 24168 15100 24280 15146
rect 24326 15108 24438 15146
rect 24373 15100 24438 15108
rect 24484 15108 24596 15146
rect 24484 15100 24532 15108
rect 23951 15056 24110 15100
rect 24162 15056 24321 15100
rect 24373 15056 24532 15100
rect 24584 15100 24596 15108
rect 24642 15108 24754 15146
rect 24642 15100 24742 15108
rect 24800 15100 24912 15146
rect 24958 15108 25071 15146
rect 25005 15100 25071 15108
rect 25117 15108 25229 15146
rect 25117 15100 25164 15108
rect 24584 15056 24742 15100
rect 24794 15056 24953 15100
rect 25005 15056 25164 15100
rect 25216 15100 25229 15108
rect 25275 15108 25387 15146
rect 25275 15100 25375 15108
rect 25433 15100 25545 15146
rect 25591 15108 25863 15146
rect 25216 15056 25375 15100
rect 25427 15056 25586 15100
rect 25638 15056 25863 15108
rect 23751 15031 25863 15056
rect 23751 14985 25763 15031
rect 25809 14985 25863 15031
rect 23751 14982 25863 14985
rect 23751 14936 23806 14982
rect 23852 14936 23964 14982
rect 24010 14936 24122 14982
rect 24168 14936 24280 14982
rect 24326 14936 24438 14982
rect 24484 14936 24596 14982
rect 24642 14936 24754 14982
rect 24800 14936 24912 14982
rect 24958 14936 25071 14982
rect 25117 14936 25229 14982
rect 25275 14936 25387 14982
rect 25433 14936 25545 14982
rect 25591 14936 25863 14982
rect 23751 14891 25863 14936
rect 22366 14843 23338 14883
rect 13591 14798 13999 14843
rect 13439 14791 13478 14798
rect 13986 14797 13999 14798
rect 14045 14797 14102 14843
rect 14148 14797 14205 14843
rect 14251 14797 14309 14843
rect 14355 14797 14413 14843
rect 14459 14797 14517 14843
rect 14563 14797 14621 14843
rect 14667 14797 14725 14843
rect 14771 14797 14829 14843
rect 14875 14797 14933 14843
rect 14979 14797 15037 14843
rect 15083 14797 15141 14843
rect 15187 14797 15245 14843
rect 15291 14797 15304 14843
rect 15755 14797 15768 14843
rect 15814 14797 15882 14843
rect 15928 14797 15996 14843
rect 16042 14797 16110 14843
rect 16156 14797 16224 14843
rect 16270 14797 16669 14843
rect 16715 14797 16772 14843
rect 16818 14797 16875 14843
rect 16921 14797 16979 14843
rect 17025 14797 17083 14843
rect 17129 14797 17187 14843
rect 17233 14797 17291 14843
rect 17337 14797 17395 14843
rect 17441 14797 17499 14843
rect 17545 14797 17603 14843
rect 17649 14797 17707 14843
rect 17753 14797 17811 14843
rect 17857 14797 17915 14843
rect 17961 14797 18346 14843
rect 18424 14797 18437 14843
rect 20319 14797 20362 14843
rect 20422 14797 20479 14843
rect 20525 14797 20573 14843
rect 20628 14797 20685 14843
rect 20731 14797 20784 14843
rect 20836 14797 20891 14843
rect 20937 14797 20950 14843
rect 21067 14797 21337 14843
rect 22097 14797 22154 14843
rect 22200 14797 22257 14843
rect 22303 14797 22360 14843
rect 22456 14797 22463 14843
rect 22509 14797 22566 14843
rect 22612 14797 22615 14843
rect 12294 14750 13478 14791
rect 15755 14757 18346 14797
rect 20112 14791 20151 14797
rect 20203 14791 20362 14797
rect 20414 14791 20573 14797
rect 20625 14791 20784 14797
rect 20836 14791 20874 14797
rect 20112 14750 20874 14791
rect 22366 14791 22404 14797
rect 22456 14791 22615 14797
rect 22667 14797 22669 14843
rect 22715 14797 22772 14843
rect 22818 14797 22826 14843
rect 22921 14797 22978 14843
rect 23024 14797 23037 14843
rect 23127 14797 23184 14843
rect 23230 14797 23248 14843
rect 23333 14797 23346 14843
rect 23751 14839 23899 14891
rect 23951 14839 24110 14891
rect 24162 14839 24321 14891
rect 24373 14839 24532 14891
rect 24584 14839 24742 14891
rect 24794 14839 24953 14891
rect 25005 14839 25164 14891
rect 25216 14839 25375 14891
rect 25427 14839 25586 14891
rect 25638 14868 25863 14891
rect 25638 14839 25763 14868
rect 23751 14822 25763 14839
rect 25809 14822 25863 14868
rect 23751 14819 25863 14822
rect 22667 14791 22826 14797
rect 22878 14791 23037 14797
rect 23089 14791 23248 14797
rect 23300 14791 23338 14797
rect 22366 14751 23338 14791
rect 23751 14773 23806 14819
rect 23852 14773 23964 14819
rect 24010 14773 24122 14819
rect 24168 14773 24280 14819
rect 24326 14773 24438 14819
rect 24484 14773 24596 14819
rect 24642 14773 24754 14819
rect 24800 14773 24912 14819
rect 24958 14773 25071 14819
rect 25117 14773 25229 14819
rect 25275 14773 25387 14819
rect 25433 14773 25545 14819
rect 25591 14773 25863 14819
rect 23751 14716 25863 14773
rect 1906 14705 2278 14716
rect 1906 14659 1960 14705
rect 2006 14659 2278 14705
rect 1906 14541 2278 14659
rect 1906 14495 1960 14541
rect 2006 14495 2278 14541
rect 79 14293 133 14339
rect 179 14293 519 14339
rect 606 14426 1688 14467
rect 606 14423 905 14426
rect 606 14377 640 14423
rect 686 14377 801 14423
rect 847 14377 905 14423
rect 606 14374 905 14377
rect 957 14423 1116 14426
rect 1168 14423 1328 14426
rect 957 14377 961 14423
rect 1007 14377 1116 14423
rect 1168 14377 1282 14423
rect 957 14374 1116 14377
rect 1168 14374 1328 14377
rect 1380 14423 1539 14426
rect 1380 14377 1444 14423
rect 1490 14377 1539 14423
rect 1380 14374 1539 14377
rect 1591 14423 1688 14426
rect 1591 14377 1607 14423
rect 1653 14377 1688 14423
rect 1591 14374 1688 14377
rect 606 14334 1688 14374
rect 1906 14465 2278 14495
rect 25490 14705 25863 14716
rect 25490 14659 25763 14705
rect 25809 14659 25863 14705
rect 25490 14541 25863 14659
rect 25490 14495 25763 14541
rect 25809 14495 25863 14541
rect 25490 14465 25863 14495
rect 27250 15195 27690 15274
rect 27250 15149 27590 15195
rect 27636 15149 27690 15195
rect 27250 15117 27690 15149
rect 27250 15071 27284 15117
rect 27330 15071 27690 15117
rect 27250 15031 27690 15071
rect 27250 14985 27590 15031
rect 27636 14985 27690 15031
rect 27250 14954 27690 14985
rect 27250 14908 27284 14954
rect 27330 14908 27690 14954
rect 27250 14868 27690 14908
rect 27250 14822 27590 14868
rect 27636 14822 27690 14868
rect 27250 14790 27690 14822
rect 27250 14744 27284 14790
rect 27330 14744 27690 14790
rect 27250 14705 27690 14744
rect 27250 14659 27590 14705
rect 27636 14659 27690 14705
rect 27250 14627 27690 14659
rect 27250 14581 27284 14627
rect 27330 14581 27690 14627
rect 27250 14541 27690 14581
rect 27250 14495 27590 14541
rect 27636 14495 27690 14541
rect 1906 14339 2125 14465
rect 867 14333 1629 14334
rect 79 14217 519 14293
rect 79 14176 439 14217
rect 79 14130 133 14176
rect 179 14171 439 14176
rect 485 14171 519 14217
rect 179 14130 519 14171
rect 79 14054 519 14130
rect 79 14013 439 14054
rect 79 13967 133 14013
rect 179 14008 439 14013
rect 485 14008 519 14054
rect 179 13967 519 14008
rect 79 13890 519 13967
rect 79 13850 439 13890
rect 79 13804 133 13850
rect 179 13844 439 13850
rect 485 13844 519 13890
rect 179 13804 519 13844
rect 79 13727 519 13804
rect 79 13686 439 13727
rect 79 13640 133 13686
rect 179 13681 439 13686
rect 485 13681 519 13727
rect 179 13640 519 13681
rect 79 13526 519 13640
rect 1906 14293 1960 14339
rect 2006 14293 2125 14339
rect 1906 14176 2125 14293
rect 1906 14130 1960 14176
rect 2006 14130 2125 14176
rect 1906 14013 2125 14130
rect 1906 13967 1960 14013
rect 2006 13967 2125 14013
rect 1906 13850 2125 13967
rect 1906 13804 1960 13850
rect 2006 13804 2125 13850
rect 1906 13686 2125 13804
rect 1906 13640 1960 13686
rect 2006 13640 2125 13686
rect 79 13523 168 13526
rect 79 13477 133 13523
rect 79 13474 168 13477
rect 220 13474 379 13526
rect 431 13474 519 13526
rect 79 13360 519 13474
rect 606 13526 1688 13567
rect 606 13523 905 13526
rect 606 13477 640 13523
rect 686 13477 801 13523
rect 847 13477 905 13523
rect 606 13474 905 13477
rect 957 13523 1116 13526
rect 1168 13523 1328 13526
rect 957 13477 961 13523
rect 1007 13477 1116 13523
rect 1168 13477 1282 13523
rect 957 13474 1116 13477
rect 1168 13474 1328 13477
rect 1380 13523 1539 13526
rect 1380 13477 1444 13523
rect 1490 13477 1539 13523
rect 1380 13474 1539 13477
rect 1591 13523 1688 13526
rect 1591 13477 1607 13523
rect 1653 13477 1688 13523
rect 1591 13474 1688 13477
rect 606 13434 1688 13474
rect 1906 13523 2125 13640
rect 1906 13477 1960 13523
rect 2006 13477 2125 13523
rect 867 13433 1629 13434
rect 79 13314 133 13360
rect 179 13317 519 13360
rect 179 13314 439 13317
rect 79 13271 439 13314
rect 485 13271 519 13317
rect 79 13196 519 13271
rect 79 13150 133 13196
rect 179 13154 519 13196
rect 179 13150 439 13154
rect 79 13108 439 13150
rect 485 13108 519 13154
rect 79 13033 519 13108
rect 79 12987 133 13033
rect 179 12990 519 13033
rect 179 12987 439 12990
rect 79 12944 439 12987
rect 485 12944 519 12990
rect 79 12870 519 12944
rect 79 12824 133 12870
rect 179 12827 519 12870
rect 179 12824 439 12827
rect 79 12781 439 12824
rect 485 12781 519 12827
rect 79 12707 519 12781
rect 79 12661 133 12707
rect 179 12661 519 12707
rect 1906 13360 2125 13477
rect 1906 13314 1960 13360
rect 2006 13314 2125 13360
rect 1906 13196 2125 13314
rect 1906 13150 1960 13196
rect 2006 13150 2125 13196
rect 1906 13033 2125 13150
rect 1906 12987 1960 13033
rect 2006 12987 2125 13033
rect 1906 12870 2125 12987
rect 1906 12824 1960 12870
rect 2006 12824 2125 12870
rect 1906 12707 2125 12824
rect 79 12539 519 12661
rect 79 12493 133 12539
rect 179 12493 519 12539
rect 606 12626 1688 12667
rect 606 12623 905 12626
rect 606 12577 640 12623
rect 686 12577 801 12623
rect 847 12577 905 12623
rect 606 12574 905 12577
rect 957 12623 1116 12626
rect 1168 12623 1328 12626
rect 957 12577 961 12623
rect 1007 12577 1116 12623
rect 1168 12577 1282 12623
rect 957 12574 1116 12577
rect 1168 12574 1328 12577
rect 1380 12623 1539 12626
rect 1380 12577 1444 12623
rect 1490 12577 1539 12623
rect 1380 12574 1539 12577
rect 1591 12623 1688 12626
rect 1591 12577 1607 12623
rect 1653 12577 1688 12623
rect 1591 12574 1688 12577
rect 606 12534 1688 12574
rect 1906 12661 1960 12707
rect 2006 12661 2125 12707
rect 1906 12539 2125 12661
rect 867 12533 1629 12534
rect 79 12417 519 12493
rect 79 12376 439 12417
rect 79 12330 133 12376
rect 179 12371 439 12376
rect 485 12371 519 12417
rect 179 12330 519 12371
rect 79 12254 519 12330
rect 79 12213 439 12254
rect 79 12167 133 12213
rect 179 12208 439 12213
rect 485 12208 519 12254
rect 179 12167 519 12208
rect 79 12090 519 12167
rect 79 12050 439 12090
rect 79 12004 133 12050
rect 179 12044 439 12050
rect 485 12044 519 12090
rect 179 12004 519 12044
rect 79 11927 519 12004
rect 79 11886 439 11927
rect 79 11840 133 11886
rect 179 11881 439 11886
rect 485 11881 519 11927
rect 179 11840 519 11881
rect 79 11726 519 11840
rect 1906 12493 1960 12539
rect 2006 12493 2125 12539
rect 1906 12376 2125 12493
rect 1906 12330 1960 12376
rect 2006 12330 2125 12376
rect 1906 12213 2125 12330
rect 1906 12167 1960 12213
rect 2006 12167 2125 12213
rect 1906 12050 2125 12167
rect 1906 12004 1960 12050
rect 2006 12004 2125 12050
rect 1906 11886 2125 12004
rect 1906 11840 1960 11886
rect 2006 11840 2125 11886
rect 79 11723 168 11726
rect 79 11677 133 11723
rect 79 11674 168 11677
rect 220 11674 379 11726
rect 431 11674 519 11726
rect 79 11560 519 11674
rect 606 11726 1688 11767
rect 606 11723 905 11726
rect 606 11677 640 11723
rect 686 11677 801 11723
rect 847 11677 905 11723
rect 606 11674 905 11677
rect 957 11723 1116 11726
rect 1168 11723 1328 11726
rect 957 11677 961 11723
rect 1007 11677 1116 11723
rect 1168 11677 1282 11723
rect 957 11674 1116 11677
rect 1168 11674 1328 11677
rect 1380 11723 1539 11726
rect 1380 11677 1444 11723
rect 1490 11677 1539 11723
rect 1380 11674 1539 11677
rect 1591 11723 1688 11726
rect 1591 11677 1607 11723
rect 1653 11677 1688 11723
rect 1591 11674 1688 11677
rect 606 11634 1688 11674
rect 1906 11723 2125 11840
rect 1906 11677 1960 11723
rect 2006 11677 2125 11723
rect 867 11633 1629 11634
rect 79 11514 133 11560
rect 179 11517 519 11560
rect 179 11514 439 11517
rect 79 11471 439 11514
rect 485 11471 519 11517
rect 79 11396 519 11471
rect 79 11350 133 11396
rect 179 11354 519 11396
rect 179 11350 439 11354
rect 79 11308 439 11350
rect 485 11308 519 11354
rect 79 11233 519 11308
rect 79 11187 133 11233
rect 179 11190 519 11233
rect 179 11187 439 11190
rect 79 11144 439 11187
rect 485 11144 519 11190
rect 79 11070 519 11144
rect 79 11024 133 11070
rect 179 11027 519 11070
rect 179 11024 439 11027
rect 79 10981 439 11024
rect 485 10981 519 11027
rect 79 10907 519 10981
rect 79 10861 133 10907
rect 179 10861 519 10907
rect 1906 11560 2125 11677
rect 1906 11514 1960 11560
rect 2006 11514 2125 11560
rect 1906 11396 2125 11514
rect 1906 11350 1960 11396
rect 2006 11350 2125 11396
rect 1906 11233 2125 11350
rect 1906 11187 1960 11233
rect 2006 11187 2125 11233
rect 1906 11070 2125 11187
rect 1906 11024 1960 11070
rect 2006 11024 2125 11070
rect 1906 10907 2125 11024
rect 79 10739 519 10861
rect 79 10693 133 10739
rect 179 10693 519 10739
rect 606 10826 1688 10867
rect 606 10823 905 10826
rect 606 10777 640 10823
rect 686 10777 801 10823
rect 847 10777 905 10823
rect 606 10774 905 10777
rect 957 10823 1116 10826
rect 1168 10823 1328 10826
rect 957 10777 961 10823
rect 1007 10777 1116 10823
rect 1168 10777 1282 10823
rect 957 10774 1116 10777
rect 1168 10774 1328 10777
rect 1380 10823 1539 10826
rect 1380 10777 1444 10823
rect 1490 10777 1539 10823
rect 1380 10774 1539 10777
rect 1591 10823 1688 10826
rect 1591 10777 1607 10823
rect 1653 10777 1688 10823
rect 1591 10774 1688 10777
rect 606 10734 1688 10774
rect 1906 10861 1960 10907
rect 2006 10861 2125 10907
rect 1906 10739 2125 10861
rect 867 10733 1629 10734
rect 79 10617 519 10693
rect 79 10576 439 10617
rect 79 10530 133 10576
rect 179 10571 439 10576
rect 485 10571 519 10617
rect 179 10530 519 10571
rect 79 10454 519 10530
rect 79 10413 439 10454
rect 79 10367 133 10413
rect 179 10408 439 10413
rect 485 10408 519 10454
rect 179 10367 519 10408
rect 79 10290 519 10367
rect 79 10250 439 10290
rect 79 10204 133 10250
rect 179 10244 439 10250
rect 485 10244 519 10290
rect 179 10204 519 10244
rect 79 10127 519 10204
rect 79 10086 439 10127
rect 79 10040 133 10086
rect 179 10081 439 10086
rect 485 10081 519 10127
rect 179 10040 519 10081
rect 79 9926 519 10040
rect 1906 10693 1960 10739
rect 2006 10693 2125 10739
rect 1906 10576 2125 10693
rect 1906 10530 1960 10576
rect 2006 10530 2125 10576
rect 1906 10413 2125 10530
rect 1906 10367 1960 10413
rect 2006 10367 2125 10413
rect 1906 10250 2125 10367
rect 1906 10204 1960 10250
rect 2006 10204 2125 10250
rect 1906 10086 2125 10204
rect 1906 10040 1960 10086
rect 2006 10040 2125 10086
rect 79 9923 168 9926
rect 79 9877 133 9923
rect 79 9874 168 9877
rect 220 9874 379 9926
rect 431 9874 519 9926
rect 79 9760 519 9874
rect 606 9926 1688 9967
rect 606 9923 905 9926
rect 606 9877 640 9923
rect 686 9877 801 9923
rect 847 9877 905 9923
rect 606 9874 905 9877
rect 957 9923 1116 9926
rect 1168 9923 1328 9926
rect 957 9877 961 9923
rect 1007 9877 1116 9923
rect 1168 9877 1282 9923
rect 957 9874 1116 9877
rect 1168 9874 1328 9877
rect 1380 9923 1539 9926
rect 1380 9877 1444 9923
rect 1490 9877 1539 9923
rect 1380 9874 1539 9877
rect 1591 9923 1688 9926
rect 1591 9877 1607 9923
rect 1653 9877 1688 9923
rect 1591 9874 1688 9877
rect 606 9834 1688 9874
rect 1906 9923 2125 10040
rect 1906 9877 1960 9923
rect 2006 9877 2125 9923
rect 867 9833 1629 9834
rect 79 9714 133 9760
rect 179 9717 519 9760
rect 179 9714 439 9717
rect 79 9671 439 9714
rect 485 9671 519 9717
rect 79 9596 519 9671
rect 79 9550 133 9596
rect 179 9554 519 9596
rect 179 9550 439 9554
rect 79 9508 439 9550
rect 485 9508 519 9554
rect 79 9433 519 9508
rect 79 9387 133 9433
rect 179 9390 519 9433
rect 179 9387 439 9390
rect 79 9344 439 9387
rect 485 9344 519 9390
rect 79 9270 519 9344
rect 79 9224 133 9270
rect 179 9227 519 9270
rect 179 9224 439 9227
rect 79 9181 439 9224
rect 485 9181 519 9227
rect 79 9107 519 9181
rect 79 9061 133 9107
rect 179 9061 519 9107
rect 1906 9760 2125 9877
rect 1906 9714 1960 9760
rect 2006 9714 2125 9760
rect 1906 9596 2125 9714
rect 1906 9550 1960 9596
rect 2006 9550 2125 9596
rect 1906 9433 2125 9550
rect 1906 9387 1960 9433
rect 2006 9387 2125 9433
rect 1906 9270 2125 9387
rect 1906 9224 1960 9270
rect 2006 9224 2125 9270
rect 1906 9107 2125 9224
rect 79 8939 519 9061
rect 79 8893 133 8939
rect 179 8893 519 8939
rect 606 9026 1688 9067
rect 606 9023 905 9026
rect 606 8977 640 9023
rect 686 8977 801 9023
rect 847 8977 905 9023
rect 606 8974 905 8977
rect 957 9023 1116 9026
rect 1168 9023 1328 9026
rect 957 8977 961 9023
rect 1007 8977 1116 9023
rect 1168 8977 1282 9023
rect 957 8974 1116 8977
rect 1168 8974 1328 8977
rect 1380 9023 1539 9026
rect 1380 8977 1444 9023
rect 1490 8977 1539 9023
rect 1380 8974 1539 8977
rect 1591 9023 1688 9026
rect 1591 8977 1607 9023
rect 1653 8977 1688 9023
rect 1591 8974 1688 8977
rect 606 8934 1688 8974
rect 1906 9061 1960 9107
rect 2006 9061 2125 9107
rect 1906 8939 2125 9061
rect 867 8933 1629 8934
rect 79 8817 519 8893
rect 79 8776 439 8817
rect 79 8730 133 8776
rect 179 8771 439 8776
rect 485 8771 519 8817
rect 179 8730 519 8771
rect 79 8654 519 8730
rect 79 8613 439 8654
rect 79 8567 133 8613
rect 179 8608 439 8613
rect 485 8608 519 8654
rect 179 8567 519 8608
rect 79 8490 519 8567
rect 79 8450 439 8490
rect 79 8404 133 8450
rect 179 8444 439 8450
rect 485 8444 519 8490
rect 179 8404 519 8444
rect 79 8327 519 8404
rect 79 8286 439 8327
rect 79 8240 133 8286
rect 179 8281 439 8286
rect 485 8281 519 8327
rect 179 8240 519 8281
rect 79 8126 519 8240
rect 1906 8893 1960 8939
rect 2006 8893 2125 8939
rect 1906 8776 2125 8893
rect 1906 8730 1960 8776
rect 2006 8730 2125 8776
rect 1906 8613 2125 8730
rect 1906 8567 1960 8613
rect 2006 8567 2125 8613
rect 1906 8450 2125 8567
rect 1906 8404 1960 8450
rect 2006 8404 2125 8450
rect 1906 8286 2125 8404
rect 1906 8240 1960 8286
rect 2006 8240 2125 8286
rect 79 8123 168 8126
rect 79 8077 133 8123
rect 79 8074 168 8077
rect 220 8074 379 8126
rect 431 8074 519 8126
rect 79 7960 519 8074
rect 606 8126 1688 8167
rect 606 8123 905 8126
rect 606 8077 640 8123
rect 686 8077 801 8123
rect 847 8077 905 8123
rect 606 8074 905 8077
rect 957 8123 1116 8126
rect 1168 8123 1328 8126
rect 957 8077 961 8123
rect 1007 8077 1116 8123
rect 1168 8077 1282 8123
rect 957 8074 1116 8077
rect 1168 8074 1328 8077
rect 1380 8123 1539 8126
rect 1380 8077 1444 8123
rect 1490 8077 1539 8123
rect 1380 8074 1539 8077
rect 1591 8123 1688 8126
rect 1591 8077 1607 8123
rect 1653 8077 1688 8123
rect 1591 8074 1688 8077
rect 606 8034 1688 8074
rect 1906 8123 2125 8240
rect 1906 8077 1960 8123
rect 2006 8077 2125 8123
rect 867 8033 1629 8034
rect 79 7914 133 7960
rect 179 7917 519 7960
rect 179 7914 439 7917
rect 79 7871 439 7914
rect 485 7871 519 7917
rect 79 7796 519 7871
rect 79 7750 133 7796
rect 179 7754 519 7796
rect 179 7750 439 7754
rect 79 7708 439 7750
rect 485 7708 519 7754
rect 79 7633 519 7708
rect 79 7587 133 7633
rect 179 7590 519 7633
rect 179 7587 439 7590
rect 79 7544 439 7587
rect 485 7544 519 7590
rect 79 7470 519 7544
rect 79 7424 133 7470
rect 179 7427 519 7470
rect 179 7424 439 7427
rect 79 7381 439 7424
rect 485 7381 519 7427
rect 79 7307 519 7381
rect 79 7261 133 7307
rect 179 7261 519 7307
rect 1906 7960 2125 8077
rect 1906 7914 1960 7960
rect 2006 7914 2125 7960
rect 1906 7796 2125 7914
rect 1906 7750 1960 7796
rect 2006 7750 2125 7796
rect 1906 7633 2125 7750
rect 1906 7587 1960 7633
rect 2006 7587 2125 7633
rect 1906 7470 2125 7587
rect 1906 7424 1960 7470
rect 2006 7424 2125 7470
rect 1906 7307 2125 7424
rect 79 7139 519 7261
rect 79 7093 133 7139
rect 179 7093 519 7139
rect 606 7226 1688 7267
rect 606 7223 905 7226
rect 606 7177 640 7223
rect 686 7177 801 7223
rect 847 7177 905 7223
rect 606 7174 905 7177
rect 957 7223 1116 7226
rect 1168 7223 1328 7226
rect 957 7177 961 7223
rect 1007 7177 1116 7223
rect 1168 7177 1282 7223
rect 957 7174 1116 7177
rect 1168 7174 1328 7177
rect 1380 7223 1539 7226
rect 1380 7177 1444 7223
rect 1490 7177 1539 7223
rect 1380 7174 1539 7177
rect 1591 7223 1688 7226
rect 1591 7177 1607 7223
rect 1653 7177 1688 7223
rect 1591 7174 1688 7177
rect 606 7134 1688 7174
rect 1906 7261 1960 7307
rect 2006 7261 2125 7307
rect 1906 7139 2125 7261
rect 867 7133 1629 7134
rect 79 7017 519 7093
rect 79 6976 439 7017
rect 79 6930 133 6976
rect 179 6971 439 6976
rect 485 6971 519 7017
rect 179 6930 519 6971
rect 79 6854 519 6930
rect 79 6813 439 6854
rect 79 6767 133 6813
rect 179 6808 439 6813
rect 485 6808 519 6854
rect 179 6767 519 6808
rect 79 6690 519 6767
rect 79 6650 439 6690
rect 79 6604 133 6650
rect 179 6644 439 6650
rect 485 6644 519 6690
rect 179 6604 519 6644
rect 79 6527 519 6604
rect 79 6486 439 6527
rect 79 6440 133 6486
rect 179 6481 439 6486
rect 485 6481 519 6527
rect 179 6440 519 6481
rect 79 6326 519 6440
rect 1906 7093 1960 7139
rect 2006 7093 2125 7139
rect 1906 6976 2125 7093
rect 1906 6930 1960 6976
rect 2006 6930 2125 6976
rect 1906 6813 2125 6930
rect 1906 6767 1960 6813
rect 2006 6767 2125 6813
rect 1906 6650 2125 6767
rect 1906 6604 1960 6650
rect 2006 6604 2125 6650
rect 1906 6486 2125 6604
rect 1906 6440 1960 6486
rect 2006 6440 2125 6486
rect 79 6323 168 6326
rect 79 6277 133 6323
rect 79 6274 168 6277
rect 220 6274 379 6326
rect 431 6274 519 6326
rect 79 6160 519 6274
rect 606 6326 1688 6367
rect 606 6323 905 6326
rect 606 6277 640 6323
rect 686 6277 801 6323
rect 847 6277 905 6323
rect 606 6274 905 6277
rect 957 6323 1116 6326
rect 1168 6323 1328 6326
rect 957 6277 961 6323
rect 1007 6277 1116 6323
rect 1168 6277 1282 6323
rect 957 6274 1116 6277
rect 1168 6274 1328 6277
rect 1380 6323 1539 6326
rect 1380 6277 1444 6323
rect 1490 6277 1539 6323
rect 1380 6274 1539 6277
rect 1591 6323 1688 6326
rect 1591 6277 1607 6323
rect 1653 6277 1688 6323
rect 1591 6274 1688 6277
rect 606 6234 1688 6274
rect 1906 6323 2125 6440
rect 1906 6277 1960 6323
rect 2006 6277 2125 6323
rect 867 6233 1629 6234
rect 79 6114 133 6160
rect 179 6117 519 6160
rect 179 6114 439 6117
rect 79 6071 439 6114
rect 485 6071 519 6117
rect 79 5996 519 6071
rect 79 5950 133 5996
rect 179 5954 519 5996
rect 179 5950 439 5954
rect 79 5908 439 5950
rect 485 5908 519 5954
rect 79 5833 519 5908
rect 79 5787 133 5833
rect 179 5790 519 5833
rect 179 5787 439 5790
rect 79 5744 439 5787
rect 485 5744 519 5790
rect 79 5670 519 5744
rect 79 5624 133 5670
rect 179 5627 519 5670
rect 179 5624 439 5627
rect 79 5581 439 5624
rect 485 5581 519 5627
rect 79 5507 519 5581
rect 79 5461 133 5507
rect 179 5461 519 5507
rect 1906 6160 2125 6277
rect 1906 6114 1960 6160
rect 2006 6114 2125 6160
rect 1906 5996 2125 6114
rect 1906 5950 1960 5996
rect 2006 5950 2125 5996
rect 1906 5833 2125 5950
rect 1906 5787 1960 5833
rect 2006 5787 2125 5833
rect 1906 5670 2125 5787
rect 1906 5624 1960 5670
rect 2006 5624 2125 5670
rect 1906 5507 2125 5624
rect 79 5339 519 5461
rect 79 5293 133 5339
rect 179 5293 519 5339
rect 606 5426 1688 5467
rect 606 5423 905 5426
rect 606 5377 640 5423
rect 686 5377 801 5423
rect 847 5377 905 5423
rect 606 5374 905 5377
rect 957 5423 1116 5426
rect 1168 5423 1328 5426
rect 957 5377 961 5423
rect 1007 5377 1116 5423
rect 1168 5377 1282 5423
rect 957 5374 1116 5377
rect 1168 5374 1328 5377
rect 1380 5423 1539 5426
rect 1380 5377 1444 5423
rect 1490 5377 1539 5423
rect 1380 5374 1539 5377
rect 1591 5423 1688 5426
rect 1591 5377 1607 5423
rect 1653 5377 1688 5423
rect 1591 5374 1688 5377
rect 606 5334 1688 5374
rect 1906 5461 1960 5507
rect 2006 5461 2125 5507
rect 1906 5339 2125 5461
rect 867 5333 1629 5334
rect 79 5217 519 5293
rect 79 5176 439 5217
rect 79 5130 133 5176
rect 179 5171 439 5176
rect 485 5171 519 5217
rect 179 5130 519 5171
rect 79 5054 519 5130
rect 79 5013 439 5054
rect 79 4967 133 5013
rect 179 5008 439 5013
rect 485 5008 519 5054
rect 179 4967 519 5008
rect 79 4890 519 4967
rect 79 4850 439 4890
rect 79 4804 133 4850
rect 179 4844 439 4850
rect 485 4844 519 4890
rect 179 4804 519 4844
rect 79 4727 519 4804
rect 79 4686 439 4727
rect 79 4640 133 4686
rect 179 4681 439 4686
rect 485 4681 519 4727
rect 179 4640 519 4681
rect 79 4526 519 4640
rect 1906 5293 1960 5339
rect 2006 5293 2125 5339
rect 1906 5176 2125 5293
rect 1906 5130 1960 5176
rect 2006 5130 2125 5176
rect 1906 5013 2125 5130
rect 1906 4967 1960 5013
rect 2006 4967 2125 5013
rect 1906 4850 2125 4967
rect 1906 4804 1960 4850
rect 2006 4804 2125 4850
rect 1906 4686 2125 4804
rect 1906 4640 1960 4686
rect 2006 4640 2125 4686
rect 79 4523 168 4526
rect 79 4477 133 4523
rect 79 4474 168 4477
rect 220 4474 379 4526
rect 431 4474 519 4526
rect 79 4360 519 4474
rect 606 4526 1688 4567
rect 606 4523 905 4526
rect 606 4477 640 4523
rect 686 4477 801 4523
rect 847 4477 905 4523
rect 606 4474 905 4477
rect 957 4523 1116 4526
rect 1168 4523 1328 4526
rect 957 4477 961 4523
rect 1007 4477 1116 4523
rect 1168 4477 1282 4523
rect 957 4474 1116 4477
rect 1168 4474 1328 4477
rect 1380 4523 1539 4526
rect 1380 4477 1444 4523
rect 1490 4477 1539 4523
rect 1380 4474 1539 4477
rect 1591 4523 1688 4526
rect 1591 4477 1607 4523
rect 1653 4477 1688 4523
rect 1591 4474 1688 4477
rect 606 4434 1688 4474
rect 1906 4523 2125 4640
rect 1906 4477 1960 4523
rect 2006 4477 2125 4523
rect 867 4433 1629 4434
rect 79 4314 133 4360
rect 179 4317 519 4360
rect 179 4314 439 4317
rect 79 4271 439 4314
rect 485 4271 519 4317
rect 79 4196 519 4271
rect 79 4150 133 4196
rect 179 4154 519 4196
rect 179 4150 439 4154
rect 79 4108 439 4150
rect 485 4108 519 4154
rect 79 4033 519 4108
rect 79 3987 133 4033
rect 179 3990 519 4033
rect 179 3987 439 3990
rect 79 3944 439 3987
rect 485 3944 519 3990
rect 79 3870 519 3944
rect 79 3824 133 3870
rect 179 3827 519 3870
rect 179 3824 439 3827
rect 79 3781 439 3824
rect 485 3781 519 3827
rect 79 3707 519 3781
rect 79 3661 133 3707
rect 179 3661 519 3707
rect 1906 4360 2125 4477
rect 1906 4314 1960 4360
rect 2006 4314 2125 4360
rect 1906 4196 2125 4314
rect 1906 4150 1960 4196
rect 2006 4150 2125 4196
rect 1906 4033 2125 4150
rect 1906 3987 1960 4033
rect 2006 3987 2125 4033
rect 1906 3870 2125 3987
rect 1906 3824 1960 3870
rect 2006 3824 2125 3870
rect 1906 3707 2125 3824
rect 79 3539 519 3661
rect 79 3493 133 3539
rect 179 3493 519 3539
rect 606 3626 1688 3667
rect 606 3623 905 3626
rect 606 3577 640 3623
rect 686 3577 801 3623
rect 847 3577 905 3623
rect 606 3574 905 3577
rect 957 3623 1116 3626
rect 1168 3623 1328 3626
rect 957 3577 961 3623
rect 1007 3577 1116 3623
rect 1168 3577 1282 3623
rect 957 3574 1116 3577
rect 1168 3574 1328 3577
rect 1380 3623 1539 3626
rect 1380 3577 1444 3623
rect 1490 3577 1539 3623
rect 1380 3574 1539 3577
rect 1591 3623 1688 3626
rect 1591 3577 1607 3623
rect 1653 3577 1688 3623
rect 1591 3574 1688 3577
rect 606 3534 1688 3574
rect 1906 3661 1960 3707
rect 2006 3661 2125 3707
rect 1906 3539 2125 3661
rect 867 3533 1629 3534
rect 79 3417 519 3493
rect 79 3376 439 3417
rect 79 3330 133 3376
rect 179 3371 439 3376
rect 485 3371 519 3417
rect 179 3330 519 3371
rect 79 3254 519 3330
rect 79 3213 439 3254
rect 79 3167 133 3213
rect 179 3208 439 3213
rect 485 3208 519 3254
rect 179 3167 519 3208
rect 79 3090 519 3167
rect 79 3050 439 3090
rect 79 3004 133 3050
rect 179 3044 439 3050
rect 485 3044 519 3090
rect 179 3004 519 3044
rect 79 2927 519 3004
rect 79 2886 439 2927
rect 79 2840 133 2886
rect 179 2881 439 2886
rect 485 2881 519 2927
rect 179 2840 519 2881
rect 79 2726 519 2840
rect 1906 3493 1960 3539
rect 2006 3493 2125 3539
rect 1906 3376 2125 3493
rect 1906 3330 1960 3376
rect 2006 3330 2125 3376
rect 1906 3213 2125 3330
rect 1906 3167 1960 3213
rect 2006 3167 2125 3213
rect 1906 3050 2125 3167
rect 1906 3004 1960 3050
rect 2006 3004 2125 3050
rect 1906 2886 2125 3004
rect 1906 2840 1960 2886
rect 2006 2840 2125 2886
rect 79 2723 168 2726
rect 79 2677 133 2723
rect 79 2674 168 2677
rect 220 2674 379 2726
rect 431 2674 519 2726
rect 79 2560 519 2674
rect 606 2726 1688 2767
rect 606 2723 905 2726
rect 606 2677 640 2723
rect 686 2677 801 2723
rect 847 2677 905 2723
rect 606 2674 905 2677
rect 957 2723 1116 2726
rect 1168 2723 1328 2726
rect 957 2677 961 2723
rect 1007 2677 1116 2723
rect 1168 2677 1282 2723
rect 957 2674 1116 2677
rect 1168 2674 1328 2677
rect 1380 2723 1539 2726
rect 1380 2677 1444 2723
rect 1490 2677 1539 2723
rect 1380 2674 1539 2677
rect 1591 2723 1688 2726
rect 1591 2677 1607 2723
rect 1653 2677 1688 2723
rect 1591 2674 1688 2677
rect 606 2634 1688 2674
rect 1906 2723 2125 2840
rect 1906 2677 1960 2723
rect 2006 2677 2125 2723
rect 867 2633 1629 2634
rect 79 2514 133 2560
rect 179 2517 519 2560
rect 179 2514 439 2517
rect 79 2471 439 2514
rect 485 2471 519 2517
rect 79 2396 519 2471
rect 79 2350 133 2396
rect 179 2354 519 2396
rect 179 2350 439 2354
rect 79 2308 439 2350
rect 485 2308 519 2354
rect 79 2233 519 2308
rect 79 2187 133 2233
rect 179 2190 519 2233
rect 179 2187 439 2190
rect 79 2144 439 2187
rect 485 2144 519 2190
rect 79 2070 519 2144
rect 79 2024 133 2070
rect 179 2027 519 2070
rect 179 2024 439 2027
rect 79 1981 439 2024
rect 485 1981 519 2027
rect 79 1907 519 1981
rect 79 1861 133 1907
rect 179 1861 519 1907
rect 1906 2560 2125 2677
rect 1906 2514 1960 2560
rect 2006 2514 2125 2560
rect 1906 2396 2125 2514
rect 1906 2350 1960 2396
rect 2006 2350 2125 2396
rect 1906 2233 2125 2350
rect 1906 2187 1960 2233
rect 2006 2187 2125 2233
rect 1906 2070 2125 2187
rect 1906 2024 1960 2070
rect 2006 2024 2125 2070
rect 1906 1907 2125 2024
rect 79 1739 519 1861
rect 79 1693 133 1739
rect 179 1693 519 1739
rect 606 1826 1688 1867
rect 606 1823 905 1826
rect 606 1777 640 1823
rect 686 1777 801 1823
rect 847 1777 905 1823
rect 606 1774 905 1777
rect 957 1823 1116 1826
rect 1168 1823 1328 1826
rect 957 1777 961 1823
rect 1007 1777 1116 1823
rect 1168 1777 1282 1823
rect 957 1774 1116 1777
rect 1168 1774 1328 1777
rect 1380 1823 1539 1826
rect 1380 1777 1444 1823
rect 1490 1777 1539 1823
rect 1380 1774 1539 1777
rect 1591 1823 1688 1826
rect 1591 1777 1607 1823
rect 1653 1777 1688 1823
rect 1591 1774 1688 1777
rect 606 1734 1688 1774
rect 1906 1861 1960 1907
rect 2006 1861 2125 1907
rect 1906 1739 2125 1861
rect 867 1733 1629 1734
rect 79 1617 519 1693
rect 79 1576 439 1617
rect 79 1530 133 1576
rect 179 1571 439 1576
rect 485 1571 519 1617
rect 179 1530 519 1571
rect 79 1454 519 1530
rect 79 1413 439 1454
rect 79 1367 133 1413
rect 179 1408 439 1413
rect 485 1408 519 1454
rect 179 1367 519 1408
rect 79 1290 519 1367
rect 79 1250 439 1290
rect 79 1204 133 1250
rect 179 1244 439 1250
rect 485 1244 519 1290
rect 179 1204 519 1244
rect 79 1127 519 1204
rect 79 1086 439 1127
rect 79 1040 133 1086
rect 179 1081 439 1086
rect 485 1081 519 1127
rect 179 1040 519 1081
rect 79 926 519 1040
rect 1906 1693 1960 1739
rect 2006 1693 2125 1739
rect 1906 1576 2125 1693
rect 1906 1530 1960 1576
rect 2006 1530 2125 1576
rect 1906 1413 2125 1530
rect 1906 1367 1960 1413
rect 2006 1367 2125 1413
rect 1906 1250 2125 1367
rect 1906 1204 1960 1250
rect 2006 1204 2125 1250
rect 1906 1086 2125 1204
rect 1906 1040 1960 1086
rect 2006 1040 2125 1086
rect 79 923 168 926
rect 79 877 133 923
rect 79 874 168 877
rect 220 874 379 926
rect 431 874 519 926
rect 79 760 519 874
rect 606 926 1688 967
rect 606 923 905 926
rect 606 877 640 923
rect 686 877 801 923
rect 847 877 905 923
rect 606 874 905 877
rect 957 923 1116 926
rect 1168 923 1328 926
rect 957 877 961 923
rect 1007 877 1116 923
rect 1168 877 1282 923
rect 957 874 1116 877
rect 1168 874 1328 877
rect 1380 923 1539 926
rect 1380 877 1444 923
rect 1490 877 1539 923
rect 1380 874 1539 877
rect 1591 923 1688 926
rect 1591 877 1607 923
rect 1653 877 1688 923
rect 1591 874 1688 877
rect 606 834 1688 874
rect 1906 923 2125 1040
rect 1906 877 1960 923
rect 2006 877 2125 923
rect 867 833 1629 834
rect 79 714 133 760
rect 179 717 519 760
rect 179 714 439 717
rect 79 671 439 714
rect 485 671 519 717
rect 79 596 519 671
rect 79 550 133 596
rect 179 554 519 596
rect 179 550 439 554
rect 79 508 439 550
rect 485 508 519 554
rect 79 433 519 508
rect 79 387 133 433
rect 179 390 519 433
rect 179 387 439 390
rect 79 344 439 387
rect 485 344 519 390
rect 79 270 519 344
rect 79 224 133 270
rect 179 227 519 270
rect 179 224 439 227
rect 79 181 439 224
rect 485 181 519 227
rect 79 107 519 181
rect 79 61 133 107
rect 179 61 519 107
rect 1906 760 2125 877
rect 1906 714 1960 760
rect 2006 714 2125 760
rect 1906 596 2125 714
rect 1906 550 1960 596
rect 2006 550 2125 596
rect 1906 433 2125 550
rect 1906 387 1960 433
rect 2006 387 2125 433
rect 1906 270 2125 387
rect 1906 224 1960 270
rect 2006 224 2125 270
rect 1906 107 2125 224
rect 79 -100 519 61
rect 606 26 1688 67
rect 606 23 905 26
rect 606 -23 640 23
rect 686 -23 801 23
rect 847 -23 905 23
rect 606 -26 905 -23
rect 957 23 1116 26
rect 1168 23 1328 26
rect 957 -23 961 23
rect 1007 -23 1116 23
rect 1168 -23 1282 23
rect 957 -26 1116 -23
rect 1168 -26 1328 -23
rect 1380 23 1539 26
rect 1380 -23 1444 23
rect 1490 -23 1539 23
rect 1380 -26 1539 -23
rect 1591 23 1688 26
rect 1591 -23 1607 23
rect 1653 -23 1688 23
rect 1591 -26 1688 -23
rect 606 -66 1688 -26
rect 1906 61 1960 107
rect 2006 61 2125 107
rect 1906 -66 2125 61
rect 25644 14339 25863 14465
rect 25644 14293 25763 14339
rect 25809 14293 25863 14339
rect 26081 14426 27163 14467
rect 26081 14423 26178 14426
rect 26081 14377 26116 14423
rect 26162 14377 26178 14423
rect 26081 14374 26178 14377
rect 26230 14423 26389 14426
rect 26230 14377 26279 14423
rect 26325 14377 26389 14423
rect 26230 14374 26389 14377
rect 26441 14423 26601 14426
rect 26653 14423 26812 14426
rect 26487 14377 26601 14423
rect 26653 14377 26762 14423
rect 26808 14377 26812 14423
rect 26441 14374 26601 14377
rect 26653 14374 26812 14377
rect 26864 14423 27163 14426
rect 26864 14377 26922 14423
rect 26968 14377 27083 14423
rect 27129 14377 27163 14423
rect 26864 14374 27163 14377
rect 26081 14334 27163 14374
rect 27250 14339 27690 14495
rect 26140 14333 26902 14334
rect 25644 14176 25863 14293
rect 25644 14130 25763 14176
rect 25809 14130 25863 14176
rect 25644 14013 25863 14130
rect 25644 13967 25763 14013
rect 25809 13967 25863 14013
rect 25644 13850 25863 13967
rect 25644 13804 25763 13850
rect 25809 13804 25863 13850
rect 25644 13686 25863 13804
rect 25644 13640 25763 13686
rect 25809 13640 25863 13686
rect 25644 13523 25863 13640
rect 27250 14293 27590 14339
rect 27636 14293 27690 14339
rect 27250 14217 27690 14293
rect 27250 14171 27284 14217
rect 27330 14176 27690 14217
rect 27330 14171 27590 14176
rect 27250 14130 27590 14171
rect 27636 14130 27690 14176
rect 27250 14054 27690 14130
rect 27250 14008 27284 14054
rect 27330 14013 27690 14054
rect 27330 14008 27590 14013
rect 27250 13967 27590 14008
rect 27636 13967 27690 14013
rect 27250 13890 27690 13967
rect 27250 13844 27284 13890
rect 27330 13850 27690 13890
rect 27330 13844 27590 13850
rect 27250 13804 27590 13844
rect 27636 13804 27690 13850
rect 27250 13727 27690 13804
rect 27250 13681 27284 13727
rect 27330 13686 27690 13727
rect 27330 13681 27590 13686
rect 27250 13640 27590 13681
rect 27636 13640 27690 13686
rect 25644 13477 25763 13523
rect 25809 13477 25863 13523
rect 25644 13360 25863 13477
rect 26081 13526 27163 13567
rect 26081 13523 26178 13526
rect 26081 13477 26116 13523
rect 26162 13477 26178 13523
rect 26081 13474 26178 13477
rect 26230 13523 26389 13526
rect 26230 13477 26279 13523
rect 26325 13477 26389 13523
rect 26230 13474 26389 13477
rect 26441 13523 26601 13526
rect 26653 13523 26812 13526
rect 26487 13477 26601 13523
rect 26653 13477 26762 13523
rect 26808 13477 26812 13523
rect 26441 13474 26601 13477
rect 26653 13474 26812 13477
rect 26864 13523 27163 13526
rect 26864 13477 26922 13523
rect 26968 13477 27083 13523
rect 27129 13477 27163 13523
rect 26864 13474 27163 13477
rect 26081 13434 27163 13474
rect 27250 13526 27690 13640
rect 27250 13474 27338 13526
rect 27390 13474 27549 13526
rect 27601 13523 27690 13526
rect 27636 13477 27690 13523
rect 27601 13474 27690 13477
rect 26140 13433 26902 13434
rect 25644 13314 25763 13360
rect 25809 13314 25863 13360
rect 25644 13196 25863 13314
rect 25644 13150 25763 13196
rect 25809 13150 25863 13196
rect 25644 13033 25863 13150
rect 25644 12987 25763 13033
rect 25809 12987 25863 13033
rect 25644 12870 25863 12987
rect 25644 12824 25763 12870
rect 25809 12824 25863 12870
rect 25644 12707 25863 12824
rect 25644 12661 25763 12707
rect 25809 12661 25863 12707
rect 27250 13360 27690 13474
rect 27250 13317 27590 13360
rect 27250 13271 27284 13317
rect 27330 13314 27590 13317
rect 27636 13314 27690 13360
rect 27330 13271 27690 13314
rect 27250 13196 27690 13271
rect 27250 13154 27590 13196
rect 27250 13108 27284 13154
rect 27330 13150 27590 13154
rect 27636 13150 27690 13196
rect 27330 13108 27690 13150
rect 27250 13033 27690 13108
rect 27250 12990 27590 13033
rect 27250 12944 27284 12990
rect 27330 12987 27590 12990
rect 27636 12987 27690 13033
rect 27330 12944 27690 12987
rect 27250 12870 27690 12944
rect 27250 12827 27590 12870
rect 27250 12781 27284 12827
rect 27330 12824 27590 12827
rect 27636 12824 27690 12870
rect 27330 12781 27690 12824
rect 27250 12707 27690 12781
rect 25644 12539 25863 12661
rect 25644 12493 25763 12539
rect 25809 12493 25863 12539
rect 26081 12626 27163 12667
rect 26081 12623 26178 12626
rect 26081 12577 26116 12623
rect 26162 12577 26178 12623
rect 26081 12574 26178 12577
rect 26230 12623 26389 12626
rect 26230 12577 26279 12623
rect 26325 12577 26389 12623
rect 26230 12574 26389 12577
rect 26441 12623 26601 12626
rect 26653 12623 26812 12626
rect 26487 12577 26601 12623
rect 26653 12577 26762 12623
rect 26808 12577 26812 12623
rect 26441 12574 26601 12577
rect 26653 12574 26812 12577
rect 26864 12623 27163 12626
rect 26864 12577 26922 12623
rect 26968 12577 27083 12623
rect 27129 12577 27163 12623
rect 26864 12574 27163 12577
rect 26081 12534 27163 12574
rect 27250 12661 27590 12707
rect 27636 12661 27690 12707
rect 27250 12539 27690 12661
rect 26140 12533 26902 12534
rect 25644 12376 25863 12493
rect 25644 12330 25763 12376
rect 25809 12330 25863 12376
rect 25644 12213 25863 12330
rect 25644 12167 25763 12213
rect 25809 12167 25863 12213
rect 25644 12050 25863 12167
rect 25644 12004 25763 12050
rect 25809 12004 25863 12050
rect 25644 11886 25863 12004
rect 25644 11840 25763 11886
rect 25809 11840 25863 11886
rect 25644 11723 25863 11840
rect 27250 12493 27590 12539
rect 27636 12493 27690 12539
rect 27250 12417 27690 12493
rect 27250 12371 27284 12417
rect 27330 12376 27690 12417
rect 27330 12371 27590 12376
rect 27250 12330 27590 12371
rect 27636 12330 27690 12376
rect 27250 12254 27690 12330
rect 27250 12208 27284 12254
rect 27330 12213 27690 12254
rect 27330 12208 27590 12213
rect 27250 12167 27590 12208
rect 27636 12167 27690 12213
rect 27250 12090 27690 12167
rect 27250 12044 27284 12090
rect 27330 12050 27690 12090
rect 27330 12044 27590 12050
rect 27250 12004 27590 12044
rect 27636 12004 27690 12050
rect 27250 11927 27690 12004
rect 27250 11881 27284 11927
rect 27330 11886 27690 11927
rect 27330 11881 27590 11886
rect 27250 11840 27590 11881
rect 27636 11840 27690 11886
rect 25644 11677 25763 11723
rect 25809 11677 25863 11723
rect 25644 11560 25863 11677
rect 26081 11726 27163 11767
rect 26081 11723 26178 11726
rect 26081 11677 26116 11723
rect 26162 11677 26178 11723
rect 26081 11674 26178 11677
rect 26230 11723 26389 11726
rect 26230 11677 26279 11723
rect 26325 11677 26389 11723
rect 26230 11674 26389 11677
rect 26441 11723 26601 11726
rect 26653 11723 26812 11726
rect 26487 11677 26601 11723
rect 26653 11677 26762 11723
rect 26808 11677 26812 11723
rect 26441 11674 26601 11677
rect 26653 11674 26812 11677
rect 26864 11723 27163 11726
rect 26864 11677 26922 11723
rect 26968 11677 27083 11723
rect 27129 11677 27163 11723
rect 26864 11674 27163 11677
rect 26081 11634 27163 11674
rect 27250 11726 27690 11840
rect 27250 11674 27338 11726
rect 27390 11674 27549 11726
rect 27601 11723 27690 11726
rect 27636 11677 27690 11723
rect 27601 11674 27690 11677
rect 26140 11633 26902 11634
rect 25644 11514 25763 11560
rect 25809 11514 25863 11560
rect 25644 11396 25863 11514
rect 25644 11350 25763 11396
rect 25809 11350 25863 11396
rect 25644 11233 25863 11350
rect 25644 11187 25763 11233
rect 25809 11187 25863 11233
rect 25644 11070 25863 11187
rect 25644 11024 25763 11070
rect 25809 11024 25863 11070
rect 25644 10907 25863 11024
rect 25644 10861 25763 10907
rect 25809 10861 25863 10907
rect 27250 11560 27690 11674
rect 27250 11517 27590 11560
rect 27250 11471 27284 11517
rect 27330 11514 27590 11517
rect 27636 11514 27690 11560
rect 27330 11471 27690 11514
rect 27250 11396 27690 11471
rect 27250 11354 27590 11396
rect 27250 11308 27284 11354
rect 27330 11350 27590 11354
rect 27636 11350 27690 11396
rect 27330 11308 27690 11350
rect 27250 11233 27690 11308
rect 27250 11190 27590 11233
rect 27250 11144 27284 11190
rect 27330 11187 27590 11190
rect 27636 11187 27690 11233
rect 27330 11144 27690 11187
rect 27250 11070 27690 11144
rect 27250 11027 27590 11070
rect 27250 10981 27284 11027
rect 27330 11024 27590 11027
rect 27636 11024 27690 11070
rect 27330 10981 27690 11024
rect 27250 10907 27690 10981
rect 25644 10739 25863 10861
rect 25644 10693 25763 10739
rect 25809 10693 25863 10739
rect 26081 10826 27163 10867
rect 26081 10823 26178 10826
rect 26081 10777 26116 10823
rect 26162 10777 26178 10823
rect 26081 10774 26178 10777
rect 26230 10823 26389 10826
rect 26230 10777 26279 10823
rect 26325 10777 26389 10823
rect 26230 10774 26389 10777
rect 26441 10823 26601 10826
rect 26653 10823 26812 10826
rect 26487 10777 26601 10823
rect 26653 10777 26762 10823
rect 26808 10777 26812 10823
rect 26441 10774 26601 10777
rect 26653 10774 26812 10777
rect 26864 10823 27163 10826
rect 26864 10777 26922 10823
rect 26968 10777 27083 10823
rect 27129 10777 27163 10823
rect 26864 10774 27163 10777
rect 26081 10734 27163 10774
rect 27250 10861 27590 10907
rect 27636 10861 27690 10907
rect 27250 10739 27690 10861
rect 26140 10733 26902 10734
rect 25644 10576 25863 10693
rect 25644 10530 25763 10576
rect 25809 10530 25863 10576
rect 25644 10413 25863 10530
rect 25644 10367 25763 10413
rect 25809 10367 25863 10413
rect 25644 10250 25863 10367
rect 25644 10204 25763 10250
rect 25809 10204 25863 10250
rect 25644 10086 25863 10204
rect 25644 10040 25763 10086
rect 25809 10040 25863 10086
rect 25644 9923 25863 10040
rect 27250 10693 27590 10739
rect 27636 10693 27690 10739
rect 27250 10617 27690 10693
rect 27250 10571 27284 10617
rect 27330 10576 27690 10617
rect 27330 10571 27590 10576
rect 27250 10530 27590 10571
rect 27636 10530 27690 10576
rect 27250 10454 27690 10530
rect 27250 10408 27284 10454
rect 27330 10413 27690 10454
rect 27330 10408 27590 10413
rect 27250 10367 27590 10408
rect 27636 10367 27690 10413
rect 27250 10290 27690 10367
rect 27250 10244 27284 10290
rect 27330 10250 27690 10290
rect 27330 10244 27590 10250
rect 27250 10204 27590 10244
rect 27636 10204 27690 10250
rect 27250 10127 27690 10204
rect 27250 10081 27284 10127
rect 27330 10086 27690 10127
rect 27330 10081 27590 10086
rect 27250 10040 27590 10081
rect 27636 10040 27690 10086
rect 25644 9877 25763 9923
rect 25809 9877 25863 9923
rect 25644 9760 25863 9877
rect 26081 9926 27163 9967
rect 26081 9923 26178 9926
rect 26081 9877 26116 9923
rect 26162 9877 26178 9923
rect 26081 9874 26178 9877
rect 26230 9923 26389 9926
rect 26230 9877 26279 9923
rect 26325 9877 26389 9923
rect 26230 9874 26389 9877
rect 26441 9923 26601 9926
rect 26653 9923 26812 9926
rect 26487 9877 26601 9923
rect 26653 9877 26762 9923
rect 26808 9877 26812 9923
rect 26441 9874 26601 9877
rect 26653 9874 26812 9877
rect 26864 9923 27163 9926
rect 26864 9877 26922 9923
rect 26968 9877 27083 9923
rect 27129 9877 27163 9923
rect 26864 9874 27163 9877
rect 26081 9834 27163 9874
rect 27250 9926 27690 10040
rect 27250 9874 27338 9926
rect 27390 9874 27549 9926
rect 27601 9923 27690 9926
rect 27636 9877 27690 9923
rect 27601 9874 27690 9877
rect 26140 9833 26902 9834
rect 25644 9714 25763 9760
rect 25809 9714 25863 9760
rect 25644 9596 25863 9714
rect 25644 9550 25763 9596
rect 25809 9550 25863 9596
rect 25644 9433 25863 9550
rect 25644 9387 25763 9433
rect 25809 9387 25863 9433
rect 25644 9270 25863 9387
rect 25644 9224 25763 9270
rect 25809 9224 25863 9270
rect 25644 9107 25863 9224
rect 25644 9061 25763 9107
rect 25809 9061 25863 9107
rect 27250 9760 27690 9874
rect 27250 9717 27590 9760
rect 27250 9671 27284 9717
rect 27330 9714 27590 9717
rect 27636 9714 27690 9760
rect 27330 9671 27690 9714
rect 27250 9596 27690 9671
rect 27250 9554 27590 9596
rect 27250 9508 27284 9554
rect 27330 9550 27590 9554
rect 27636 9550 27690 9596
rect 27330 9508 27690 9550
rect 27250 9433 27690 9508
rect 27250 9390 27590 9433
rect 27250 9344 27284 9390
rect 27330 9387 27590 9390
rect 27636 9387 27690 9433
rect 27330 9344 27690 9387
rect 27250 9270 27690 9344
rect 27250 9227 27590 9270
rect 27250 9181 27284 9227
rect 27330 9224 27590 9227
rect 27636 9224 27690 9270
rect 27330 9181 27690 9224
rect 27250 9107 27690 9181
rect 25644 8939 25863 9061
rect 25644 8893 25763 8939
rect 25809 8893 25863 8939
rect 26081 9026 27163 9067
rect 26081 9023 26178 9026
rect 26081 8977 26116 9023
rect 26162 8977 26178 9023
rect 26081 8974 26178 8977
rect 26230 9023 26389 9026
rect 26230 8977 26279 9023
rect 26325 8977 26389 9023
rect 26230 8974 26389 8977
rect 26441 9023 26601 9026
rect 26653 9023 26812 9026
rect 26487 8977 26601 9023
rect 26653 8977 26762 9023
rect 26808 8977 26812 9023
rect 26441 8974 26601 8977
rect 26653 8974 26812 8977
rect 26864 9023 27163 9026
rect 26864 8977 26922 9023
rect 26968 8977 27083 9023
rect 27129 8977 27163 9023
rect 26864 8974 27163 8977
rect 26081 8934 27163 8974
rect 27250 9061 27590 9107
rect 27636 9061 27690 9107
rect 27250 8939 27690 9061
rect 26140 8933 26902 8934
rect 25644 8776 25863 8893
rect 25644 8730 25763 8776
rect 25809 8730 25863 8776
rect 25644 8613 25863 8730
rect 25644 8567 25763 8613
rect 25809 8567 25863 8613
rect 25644 8450 25863 8567
rect 25644 8404 25763 8450
rect 25809 8404 25863 8450
rect 25644 8286 25863 8404
rect 25644 8240 25763 8286
rect 25809 8240 25863 8286
rect 25644 8123 25863 8240
rect 27250 8893 27590 8939
rect 27636 8893 27690 8939
rect 27250 8817 27690 8893
rect 27250 8771 27284 8817
rect 27330 8776 27690 8817
rect 27330 8771 27590 8776
rect 27250 8730 27590 8771
rect 27636 8730 27690 8776
rect 27250 8654 27690 8730
rect 27250 8608 27284 8654
rect 27330 8613 27690 8654
rect 27330 8608 27590 8613
rect 27250 8567 27590 8608
rect 27636 8567 27690 8613
rect 27250 8490 27690 8567
rect 27250 8444 27284 8490
rect 27330 8450 27690 8490
rect 27330 8444 27590 8450
rect 27250 8404 27590 8444
rect 27636 8404 27690 8450
rect 27250 8327 27690 8404
rect 27250 8281 27284 8327
rect 27330 8286 27690 8327
rect 27330 8281 27590 8286
rect 27250 8240 27590 8281
rect 27636 8240 27690 8286
rect 25644 8077 25763 8123
rect 25809 8077 25863 8123
rect 25644 7960 25863 8077
rect 26081 8126 27163 8167
rect 26081 8123 26178 8126
rect 26081 8077 26116 8123
rect 26162 8077 26178 8123
rect 26081 8074 26178 8077
rect 26230 8123 26389 8126
rect 26230 8077 26279 8123
rect 26325 8077 26389 8123
rect 26230 8074 26389 8077
rect 26441 8123 26601 8126
rect 26653 8123 26812 8126
rect 26487 8077 26601 8123
rect 26653 8077 26762 8123
rect 26808 8077 26812 8123
rect 26441 8074 26601 8077
rect 26653 8074 26812 8077
rect 26864 8123 27163 8126
rect 26864 8077 26922 8123
rect 26968 8077 27083 8123
rect 27129 8077 27163 8123
rect 26864 8074 27163 8077
rect 26081 8034 27163 8074
rect 27250 8126 27690 8240
rect 27250 8074 27338 8126
rect 27390 8074 27549 8126
rect 27601 8123 27690 8126
rect 27636 8077 27690 8123
rect 27601 8074 27690 8077
rect 26140 8033 26902 8034
rect 25644 7914 25763 7960
rect 25809 7914 25863 7960
rect 25644 7796 25863 7914
rect 25644 7750 25763 7796
rect 25809 7750 25863 7796
rect 25644 7633 25863 7750
rect 25644 7587 25763 7633
rect 25809 7587 25863 7633
rect 25644 7470 25863 7587
rect 25644 7424 25763 7470
rect 25809 7424 25863 7470
rect 25644 7307 25863 7424
rect 25644 7261 25763 7307
rect 25809 7261 25863 7307
rect 27250 7960 27690 8074
rect 27250 7917 27590 7960
rect 27250 7871 27284 7917
rect 27330 7914 27590 7917
rect 27636 7914 27690 7960
rect 27330 7871 27690 7914
rect 27250 7796 27690 7871
rect 27250 7754 27590 7796
rect 27250 7708 27284 7754
rect 27330 7750 27590 7754
rect 27636 7750 27690 7796
rect 27330 7708 27690 7750
rect 27250 7633 27690 7708
rect 27250 7590 27590 7633
rect 27250 7544 27284 7590
rect 27330 7587 27590 7590
rect 27636 7587 27690 7633
rect 27330 7544 27690 7587
rect 27250 7470 27690 7544
rect 27250 7427 27590 7470
rect 27250 7381 27284 7427
rect 27330 7424 27590 7427
rect 27636 7424 27690 7470
rect 27330 7381 27690 7424
rect 27250 7307 27690 7381
rect 25644 7139 25863 7261
rect 25644 7093 25763 7139
rect 25809 7093 25863 7139
rect 26081 7226 27163 7267
rect 26081 7223 26178 7226
rect 26081 7177 26116 7223
rect 26162 7177 26178 7223
rect 26081 7174 26178 7177
rect 26230 7223 26389 7226
rect 26230 7177 26279 7223
rect 26325 7177 26389 7223
rect 26230 7174 26389 7177
rect 26441 7223 26601 7226
rect 26653 7223 26812 7226
rect 26487 7177 26601 7223
rect 26653 7177 26762 7223
rect 26808 7177 26812 7223
rect 26441 7174 26601 7177
rect 26653 7174 26812 7177
rect 26864 7223 27163 7226
rect 26864 7177 26922 7223
rect 26968 7177 27083 7223
rect 27129 7177 27163 7223
rect 26864 7174 27163 7177
rect 26081 7134 27163 7174
rect 27250 7261 27590 7307
rect 27636 7261 27690 7307
rect 27250 7139 27690 7261
rect 26140 7133 26902 7134
rect 25644 6976 25863 7093
rect 25644 6930 25763 6976
rect 25809 6930 25863 6976
rect 25644 6813 25863 6930
rect 25644 6767 25763 6813
rect 25809 6767 25863 6813
rect 25644 6650 25863 6767
rect 25644 6604 25763 6650
rect 25809 6604 25863 6650
rect 25644 6486 25863 6604
rect 25644 6440 25763 6486
rect 25809 6440 25863 6486
rect 25644 6323 25863 6440
rect 27250 7093 27590 7139
rect 27636 7093 27690 7139
rect 27250 7017 27690 7093
rect 27250 6971 27284 7017
rect 27330 6976 27690 7017
rect 27330 6971 27590 6976
rect 27250 6930 27590 6971
rect 27636 6930 27690 6976
rect 27250 6854 27690 6930
rect 27250 6808 27284 6854
rect 27330 6813 27690 6854
rect 27330 6808 27590 6813
rect 27250 6767 27590 6808
rect 27636 6767 27690 6813
rect 27250 6690 27690 6767
rect 27250 6644 27284 6690
rect 27330 6650 27690 6690
rect 27330 6644 27590 6650
rect 27250 6604 27590 6644
rect 27636 6604 27690 6650
rect 27250 6527 27690 6604
rect 27250 6481 27284 6527
rect 27330 6486 27690 6527
rect 27330 6481 27590 6486
rect 27250 6440 27590 6481
rect 27636 6440 27690 6486
rect 25644 6277 25763 6323
rect 25809 6277 25863 6323
rect 25644 6160 25863 6277
rect 26081 6326 27163 6367
rect 26081 6323 26178 6326
rect 26081 6277 26116 6323
rect 26162 6277 26178 6323
rect 26081 6274 26178 6277
rect 26230 6323 26389 6326
rect 26230 6277 26279 6323
rect 26325 6277 26389 6323
rect 26230 6274 26389 6277
rect 26441 6323 26601 6326
rect 26653 6323 26812 6326
rect 26487 6277 26601 6323
rect 26653 6277 26762 6323
rect 26808 6277 26812 6323
rect 26441 6274 26601 6277
rect 26653 6274 26812 6277
rect 26864 6323 27163 6326
rect 26864 6277 26922 6323
rect 26968 6277 27083 6323
rect 27129 6277 27163 6323
rect 26864 6274 27163 6277
rect 26081 6234 27163 6274
rect 27250 6326 27690 6440
rect 27250 6274 27338 6326
rect 27390 6274 27549 6326
rect 27601 6323 27690 6326
rect 27636 6277 27690 6323
rect 27601 6274 27690 6277
rect 26140 6233 26902 6234
rect 25644 6114 25763 6160
rect 25809 6114 25863 6160
rect 25644 5996 25863 6114
rect 25644 5950 25763 5996
rect 25809 5950 25863 5996
rect 25644 5833 25863 5950
rect 25644 5787 25763 5833
rect 25809 5787 25863 5833
rect 25644 5670 25863 5787
rect 25644 5624 25763 5670
rect 25809 5624 25863 5670
rect 25644 5507 25863 5624
rect 25644 5461 25763 5507
rect 25809 5461 25863 5507
rect 27250 6160 27690 6274
rect 27250 6117 27590 6160
rect 27250 6071 27284 6117
rect 27330 6114 27590 6117
rect 27636 6114 27690 6160
rect 27330 6071 27690 6114
rect 27250 5996 27690 6071
rect 27250 5954 27590 5996
rect 27250 5908 27284 5954
rect 27330 5950 27590 5954
rect 27636 5950 27690 5996
rect 27330 5908 27690 5950
rect 27250 5833 27690 5908
rect 27250 5790 27590 5833
rect 27250 5744 27284 5790
rect 27330 5787 27590 5790
rect 27636 5787 27690 5833
rect 27330 5744 27690 5787
rect 27250 5670 27690 5744
rect 27250 5627 27590 5670
rect 27250 5581 27284 5627
rect 27330 5624 27590 5627
rect 27636 5624 27690 5670
rect 27330 5581 27690 5624
rect 27250 5507 27690 5581
rect 25644 5339 25863 5461
rect 25644 5293 25763 5339
rect 25809 5293 25863 5339
rect 26081 5426 27163 5467
rect 26081 5423 26178 5426
rect 26081 5377 26116 5423
rect 26162 5377 26178 5423
rect 26081 5374 26178 5377
rect 26230 5423 26389 5426
rect 26230 5377 26279 5423
rect 26325 5377 26389 5423
rect 26230 5374 26389 5377
rect 26441 5423 26601 5426
rect 26653 5423 26812 5426
rect 26487 5377 26601 5423
rect 26653 5377 26762 5423
rect 26808 5377 26812 5423
rect 26441 5374 26601 5377
rect 26653 5374 26812 5377
rect 26864 5423 27163 5426
rect 26864 5377 26922 5423
rect 26968 5377 27083 5423
rect 27129 5377 27163 5423
rect 26864 5374 27163 5377
rect 26081 5334 27163 5374
rect 27250 5461 27590 5507
rect 27636 5461 27690 5507
rect 27250 5339 27690 5461
rect 26140 5333 26902 5334
rect 25644 5176 25863 5293
rect 25644 5130 25763 5176
rect 25809 5130 25863 5176
rect 25644 5013 25863 5130
rect 25644 4967 25763 5013
rect 25809 4967 25863 5013
rect 25644 4850 25863 4967
rect 25644 4804 25763 4850
rect 25809 4804 25863 4850
rect 25644 4686 25863 4804
rect 25644 4640 25763 4686
rect 25809 4640 25863 4686
rect 25644 4523 25863 4640
rect 27250 5293 27590 5339
rect 27636 5293 27690 5339
rect 27250 5217 27690 5293
rect 27250 5171 27284 5217
rect 27330 5176 27690 5217
rect 27330 5171 27590 5176
rect 27250 5130 27590 5171
rect 27636 5130 27690 5176
rect 27250 5054 27690 5130
rect 27250 5008 27284 5054
rect 27330 5013 27690 5054
rect 27330 5008 27590 5013
rect 27250 4967 27590 5008
rect 27636 4967 27690 5013
rect 27250 4890 27690 4967
rect 27250 4844 27284 4890
rect 27330 4850 27690 4890
rect 27330 4844 27590 4850
rect 27250 4804 27590 4844
rect 27636 4804 27690 4850
rect 27250 4727 27690 4804
rect 27250 4681 27284 4727
rect 27330 4686 27690 4727
rect 27330 4681 27590 4686
rect 27250 4640 27590 4681
rect 27636 4640 27690 4686
rect 25644 4477 25763 4523
rect 25809 4477 25863 4523
rect 25644 4360 25863 4477
rect 26081 4526 27163 4567
rect 26081 4523 26178 4526
rect 26081 4477 26116 4523
rect 26162 4477 26178 4523
rect 26081 4474 26178 4477
rect 26230 4523 26389 4526
rect 26230 4477 26279 4523
rect 26325 4477 26389 4523
rect 26230 4474 26389 4477
rect 26441 4523 26601 4526
rect 26653 4523 26812 4526
rect 26487 4477 26601 4523
rect 26653 4477 26762 4523
rect 26808 4477 26812 4523
rect 26441 4474 26601 4477
rect 26653 4474 26812 4477
rect 26864 4523 27163 4526
rect 26864 4477 26922 4523
rect 26968 4477 27083 4523
rect 27129 4477 27163 4523
rect 26864 4474 27163 4477
rect 26081 4434 27163 4474
rect 27250 4526 27690 4640
rect 27250 4474 27338 4526
rect 27390 4474 27549 4526
rect 27601 4523 27690 4526
rect 27636 4477 27690 4523
rect 27601 4474 27690 4477
rect 26140 4433 26902 4434
rect 25644 4314 25763 4360
rect 25809 4314 25863 4360
rect 25644 4196 25863 4314
rect 25644 4150 25763 4196
rect 25809 4150 25863 4196
rect 25644 4033 25863 4150
rect 25644 3987 25763 4033
rect 25809 3987 25863 4033
rect 25644 3870 25863 3987
rect 25644 3824 25763 3870
rect 25809 3824 25863 3870
rect 25644 3707 25863 3824
rect 25644 3661 25763 3707
rect 25809 3661 25863 3707
rect 27250 4360 27690 4474
rect 27250 4317 27590 4360
rect 27250 4271 27284 4317
rect 27330 4314 27590 4317
rect 27636 4314 27690 4360
rect 27330 4271 27690 4314
rect 27250 4196 27690 4271
rect 27250 4154 27590 4196
rect 27250 4108 27284 4154
rect 27330 4150 27590 4154
rect 27636 4150 27690 4196
rect 27330 4108 27690 4150
rect 27250 4033 27690 4108
rect 27250 3990 27590 4033
rect 27250 3944 27284 3990
rect 27330 3987 27590 3990
rect 27636 3987 27690 4033
rect 27330 3944 27690 3987
rect 27250 3870 27690 3944
rect 27250 3827 27590 3870
rect 27250 3781 27284 3827
rect 27330 3824 27590 3827
rect 27636 3824 27690 3870
rect 27330 3781 27690 3824
rect 27250 3707 27690 3781
rect 25644 3539 25863 3661
rect 25644 3493 25763 3539
rect 25809 3493 25863 3539
rect 26081 3626 27163 3667
rect 26081 3623 26178 3626
rect 26081 3577 26116 3623
rect 26162 3577 26178 3623
rect 26081 3574 26178 3577
rect 26230 3623 26389 3626
rect 26230 3577 26279 3623
rect 26325 3577 26389 3623
rect 26230 3574 26389 3577
rect 26441 3623 26601 3626
rect 26653 3623 26812 3626
rect 26487 3577 26601 3623
rect 26653 3577 26762 3623
rect 26808 3577 26812 3623
rect 26441 3574 26601 3577
rect 26653 3574 26812 3577
rect 26864 3623 27163 3626
rect 26864 3577 26922 3623
rect 26968 3577 27083 3623
rect 27129 3577 27163 3623
rect 26864 3574 27163 3577
rect 26081 3534 27163 3574
rect 27250 3661 27590 3707
rect 27636 3661 27690 3707
rect 27250 3539 27690 3661
rect 26140 3533 26902 3534
rect 25644 3376 25863 3493
rect 25644 3330 25763 3376
rect 25809 3330 25863 3376
rect 25644 3213 25863 3330
rect 25644 3167 25763 3213
rect 25809 3167 25863 3213
rect 25644 3050 25863 3167
rect 25644 3004 25763 3050
rect 25809 3004 25863 3050
rect 25644 2886 25863 3004
rect 25644 2840 25763 2886
rect 25809 2840 25863 2886
rect 25644 2723 25863 2840
rect 27250 3493 27590 3539
rect 27636 3493 27690 3539
rect 27250 3417 27690 3493
rect 27250 3371 27284 3417
rect 27330 3376 27690 3417
rect 27330 3371 27590 3376
rect 27250 3330 27590 3371
rect 27636 3330 27690 3376
rect 27250 3254 27690 3330
rect 27250 3208 27284 3254
rect 27330 3213 27690 3254
rect 27330 3208 27590 3213
rect 27250 3167 27590 3208
rect 27636 3167 27690 3213
rect 27250 3090 27690 3167
rect 27250 3044 27284 3090
rect 27330 3050 27690 3090
rect 27330 3044 27590 3050
rect 27250 3004 27590 3044
rect 27636 3004 27690 3050
rect 27250 2927 27690 3004
rect 27250 2881 27284 2927
rect 27330 2886 27690 2927
rect 27330 2881 27590 2886
rect 27250 2840 27590 2881
rect 27636 2840 27690 2886
rect 25644 2677 25763 2723
rect 25809 2677 25863 2723
rect 25644 2560 25863 2677
rect 26081 2726 27163 2767
rect 26081 2723 26178 2726
rect 26081 2677 26116 2723
rect 26162 2677 26178 2723
rect 26081 2674 26178 2677
rect 26230 2723 26389 2726
rect 26230 2677 26279 2723
rect 26325 2677 26389 2723
rect 26230 2674 26389 2677
rect 26441 2723 26601 2726
rect 26653 2723 26812 2726
rect 26487 2677 26601 2723
rect 26653 2677 26762 2723
rect 26808 2677 26812 2723
rect 26441 2674 26601 2677
rect 26653 2674 26812 2677
rect 26864 2723 27163 2726
rect 26864 2677 26922 2723
rect 26968 2677 27083 2723
rect 27129 2677 27163 2723
rect 26864 2674 27163 2677
rect 26081 2634 27163 2674
rect 27250 2726 27690 2840
rect 27250 2674 27338 2726
rect 27390 2674 27549 2726
rect 27601 2723 27690 2726
rect 27636 2677 27690 2723
rect 27601 2674 27690 2677
rect 26140 2633 26902 2634
rect 25644 2514 25763 2560
rect 25809 2514 25863 2560
rect 25644 2396 25863 2514
rect 25644 2350 25763 2396
rect 25809 2350 25863 2396
rect 25644 2233 25863 2350
rect 25644 2187 25763 2233
rect 25809 2187 25863 2233
rect 25644 2070 25863 2187
rect 25644 2024 25763 2070
rect 25809 2024 25863 2070
rect 25644 1907 25863 2024
rect 25644 1861 25763 1907
rect 25809 1861 25863 1907
rect 27250 2560 27690 2674
rect 27250 2517 27590 2560
rect 27250 2471 27284 2517
rect 27330 2514 27590 2517
rect 27636 2514 27690 2560
rect 27330 2471 27690 2514
rect 27250 2396 27690 2471
rect 27250 2354 27590 2396
rect 27250 2308 27284 2354
rect 27330 2350 27590 2354
rect 27636 2350 27690 2396
rect 27330 2308 27690 2350
rect 27250 2233 27690 2308
rect 27250 2190 27590 2233
rect 27250 2144 27284 2190
rect 27330 2187 27590 2190
rect 27636 2187 27690 2233
rect 27330 2144 27690 2187
rect 27250 2070 27690 2144
rect 27250 2027 27590 2070
rect 27250 1981 27284 2027
rect 27330 2024 27590 2027
rect 27636 2024 27690 2070
rect 27330 1981 27690 2024
rect 27250 1907 27690 1981
rect 25644 1739 25863 1861
rect 25644 1693 25763 1739
rect 25809 1693 25863 1739
rect 26081 1826 27163 1867
rect 26081 1823 26178 1826
rect 26081 1777 26116 1823
rect 26162 1777 26178 1823
rect 26081 1774 26178 1777
rect 26230 1823 26389 1826
rect 26230 1777 26279 1823
rect 26325 1777 26389 1823
rect 26230 1774 26389 1777
rect 26441 1823 26601 1826
rect 26653 1823 26812 1826
rect 26487 1777 26601 1823
rect 26653 1777 26762 1823
rect 26808 1777 26812 1823
rect 26441 1774 26601 1777
rect 26653 1774 26812 1777
rect 26864 1823 27163 1826
rect 26864 1777 26922 1823
rect 26968 1777 27083 1823
rect 27129 1777 27163 1823
rect 26864 1774 27163 1777
rect 26081 1734 27163 1774
rect 27250 1861 27590 1907
rect 27636 1861 27690 1907
rect 27250 1739 27690 1861
rect 26140 1733 26902 1734
rect 25644 1576 25863 1693
rect 25644 1530 25763 1576
rect 25809 1530 25863 1576
rect 25644 1413 25863 1530
rect 25644 1367 25763 1413
rect 25809 1367 25863 1413
rect 25644 1250 25863 1367
rect 25644 1204 25763 1250
rect 25809 1204 25863 1250
rect 25644 1086 25863 1204
rect 25644 1040 25763 1086
rect 25809 1040 25863 1086
rect 25644 923 25863 1040
rect 27250 1693 27590 1739
rect 27636 1693 27690 1739
rect 27250 1617 27690 1693
rect 27250 1571 27284 1617
rect 27330 1576 27690 1617
rect 27330 1571 27590 1576
rect 27250 1530 27590 1571
rect 27636 1530 27690 1576
rect 27250 1454 27690 1530
rect 27250 1408 27284 1454
rect 27330 1413 27690 1454
rect 27330 1408 27590 1413
rect 27250 1367 27590 1408
rect 27636 1367 27690 1413
rect 27250 1290 27690 1367
rect 27250 1244 27284 1290
rect 27330 1250 27690 1290
rect 27330 1244 27590 1250
rect 27250 1204 27590 1244
rect 27636 1204 27690 1250
rect 27250 1127 27690 1204
rect 27250 1081 27284 1127
rect 27330 1086 27690 1127
rect 27330 1081 27590 1086
rect 27250 1040 27590 1081
rect 27636 1040 27690 1086
rect 25644 877 25763 923
rect 25809 877 25863 923
rect 25644 760 25863 877
rect 26081 926 27163 967
rect 26081 923 26178 926
rect 26081 877 26116 923
rect 26162 877 26178 923
rect 26081 874 26178 877
rect 26230 923 26389 926
rect 26230 877 26279 923
rect 26325 877 26389 923
rect 26230 874 26389 877
rect 26441 923 26601 926
rect 26653 923 26812 926
rect 26487 877 26601 923
rect 26653 877 26762 923
rect 26808 877 26812 923
rect 26441 874 26601 877
rect 26653 874 26812 877
rect 26864 923 27163 926
rect 26864 877 26922 923
rect 26968 877 27083 923
rect 27129 877 27163 923
rect 26864 874 27163 877
rect 26081 834 27163 874
rect 27250 926 27690 1040
rect 27250 874 27338 926
rect 27390 874 27549 926
rect 27601 923 27690 926
rect 27636 877 27690 923
rect 27601 874 27690 877
rect 26140 833 26902 834
rect 25644 714 25763 760
rect 25809 714 25863 760
rect 25644 596 25863 714
rect 25644 550 25763 596
rect 25809 550 25863 596
rect 25644 433 25863 550
rect 25644 387 25763 433
rect 25809 387 25863 433
rect 25644 270 25863 387
rect 25644 224 25763 270
rect 25809 224 25863 270
rect 25644 107 25863 224
rect 25644 61 25763 107
rect 25809 61 25863 107
rect 27250 760 27690 874
rect 27250 717 27590 760
rect 27250 671 27284 717
rect 27330 714 27590 717
rect 27636 714 27690 760
rect 27330 671 27690 714
rect 27250 596 27690 671
rect 27250 554 27590 596
rect 27250 508 27284 554
rect 27330 550 27590 554
rect 27636 550 27690 596
rect 27330 508 27690 550
rect 27250 433 27690 508
rect 27250 390 27590 433
rect 27250 344 27284 390
rect 27330 387 27590 390
rect 27636 387 27690 433
rect 27330 344 27690 387
rect 27250 270 27690 344
rect 27250 227 27590 270
rect 27250 181 27284 227
rect 27330 224 27590 227
rect 27636 224 27690 270
rect 27330 181 27690 224
rect 27250 107 27690 181
rect 25644 -66 25863 61
rect 26081 26 27163 67
rect 26081 23 26178 26
rect 26081 -23 26116 23
rect 26162 -23 26178 23
rect 26081 -26 26178 -23
rect 26230 23 26389 26
rect 26230 -23 26279 23
rect 26325 -23 26389 23
rect 26230 -26 26389 -23
rect 26441 23 26601 26
rect 26653 23 26812 26
rect 26487 -23 26601 23
rect 26653 -23 26762 23
rect 26808 -23 26812 23
rect 26441 -26 26601 -23
rect 26653 -26 26812 -23
rect 26864 23 27163 26
rect 26864 -23 26922 23
rect 26968 -23 27083 23
rect 27129 -23 27163 23
rect 26864 -26 27163 -23
rect 26081 -66 27163 -26
rect 27250 61 27590 107
rect 27636 61 27690 107
rect 867 -67 1629 -66
rect 26140 -67 26902 -66
rect 27250 -100 27690 61
<< via1 >>
rect 168 15274 220 15326
rect 379 15274 431 15326
rect 905 15274 957 15326
rect 1116 15323 1168 15326
rect 1116 15277 1121 15323
rect 1121 15277 1167 15323
rect 1167 15277 1168 15323
rect 1116 15274 1168 15277
rect 1328 15274 1380 15326
rect 1539 15274 1591 15326
rect 2130 15309 2182 15326
rect 2341 15309 2393 15326
rect 2130 15274 2177 15309
rect 2177 15274 2182 15309
rect 2341 15274 2381 15309
rect 2381 15274 2393 15309
rect 2552 15274 2604 15326
rect 2763 15309 2815 15326
rect 2974 15309 3026 15326
rect 2763 15274 2810 15309
rect 2810 15274 2815 15309
rect 2974 15274 3014 15309
rect 3014 15274 3026 15309
rect 3184 15274 3236 15326
rect 3395 15309 3447 15326
rect 3606 15309 3658 15326
rect 3395 15274 3442 15309
rect 3442 15274 3447 15309
rect 3606 15274 3646 15309
rect 3646 15274 3658 15309
rect 3817 15274 3869 15326
rect 2130 15100 2177 15108
rect 2177 15100 2182 15108
rect 2341 15100 2381 15108
rect 2381 15100 2393 15108
rect 2130 15056 2182 15100
rect 2341 15056 2393 15100
rect 2552 15056 2604 15108
rect 2763 15100 2810 15108
rect 2810 15100 2815 15108
rect 2974 15100 3014 15108
rect 3014 15100 3026 15108
rect 2763 15056 2815 15100
rect 2974 15056 3026 15100
rect 3184 15056 3236 15108
rect 3395 15100 3442 15108
rect 3442 15100 3447 15108
rect 3606 15100 3646 15108
rect 3646 15100 3658 15108
rect 3395 15056 3447 15100
rect 3606 15056 3658 15100
rect 3817 15056 3869 15108
rect 5613 15274 5665 15326
rect 5824 15274 5876 15326
rect 6035 15274 6087 15326
rect 6246 15274 6298 15326
rect 6766 15291 6818 15306
rect 6977 15291 7029 15306
rect 7188 15291 7240 15306
rect 7399 15291 7451 15306
rect 7610 15291 7662 15306
rect 6766 15254 6818 15291
rect 6977 15254 7029 15291
rect 7188 15254 7240 15291
rect 7399 15254 7451 15291
rect 7610 15254 7662 15291
rect 11575 15279 11627 15331
rect 11755 15279 11807 15331
rect 14033 15336 14040 15378
rect 14040 15336 14085 15378
rect 14033 15326 14085 15336
rect 14244 15326 14296 15378
rect 14455 15326 14507 15378
rect 5613 15056 5665 15108
rect 5824 15067 5876 15108
rect 6035 15067 6087 15108
rect 6246 15067 6298 15108
rect 5824 15056 5875 15067
rect 5875 15056 5876 15067
rect 6035 15056 6081 15067
rect 6081 15056 6087 15067
rect 6246 15056 6287 15067
rect 6287 15056 6298 15067
rect 2130 14839 2182 14891
rect 2341 14839 2393 14891
rect 2552 14839 2604 14891
rect 2763 14839 2815 14891
rect 2974 14839 3026 14891
rect 3184 14839 3236 14891
rect 3395 14839 3447 14891
rect 3606 14839 3658 14891
rect 3817 14839 3869 14891
rect 10376 15067 10428 15074
rect 10587 15067 10639 15074
rect 10798 15067 10850 15074
rect 13569 15265 13621 15317
rect 13781 15316 13833 15317
rect 13781 15270 13782 15316
rect 13782 15270 13833 15316
rect 15100 15326 15152 15378
rect 15311 15326 15363 15378
rect 15522 15326 15574 15378
rect 15733 15326 15785 15378
rect 13781 15265 13833 15270
rect 11575 15067 11627 15113
rect 11755 15067 11807 15113
rect 10376 15022 10425 15067
rect 10425 15022 10428 15067
rect 10587 15022 10633 15067
rect 10633 15022 10639 15067
rect 10798 15022 10841 15067
rect 10841 15022 10850 15067
rect 11575 15061 11626 15067
rect 11626 15061 11627 15067
rect 11755 15061 11786 15067
rect 11786 15061 11807 15067
rect 4373 14843 4425 14845
rect 4584 14843 4636 14845
rect 4795 14843 4847 14845
rect 5006 14843 5058 14845
rect 5217 14843 5269 14845
rect 20151 15291 20203 15306
rect 20362 15291 20414 15306
rect 20573 15291 20625 15306
rect 20784 15291 20836 15306
rect 20151 15254 20203 15291
rect 20362 15254 20376 15291
rect 20376 15254 20414 15291
rect 20573 15254 20582 15291
rect 20582 15254 20625 15291
rect 20784 15254 20788 15291
rect 20788 15254 20834 15291
rect 20834 15254 20836 15291
rect 21460 15274 21512 15326
rect 21671 15274 21723 15326
rect 21882 15274 21934 15326
rect 22093 15274 22145 15326
rect 21460 15067 21512 15108
rect 21671 15067 21723 15108
rect 21882 15067 21934 15108
rect 22093 15067 22145 15108
rect 4373 14797 4425 14843
rect 4584 14797 4636 14843
rect 4795 14797 4847 14843
rect 5006 14797 5058 14843
rect 5217 14797 5257 14843
rect 5257 14797 5269 14843
rect 6766 14797 6818 14843
rect 6977 14797 7029 14843
rect 7188 14797 7240 14843
rect 7399 14797 7451 14843
rect 7610 14797 7662 14843
rect 12333 14798 12345 14843
rect 12345 14798 12385 14843
rect 12544 14798 12551 14843
rect 12551 14798 12596 14843
rect 12755 14798 12759 14843
rect 12759 14798 12807 14843
rect 12966 14798 12967 14843
rect 12967 14798 13018 14843
rect 4373 14793 4425 14797
rect 4584 14793 4636 14797
rect 4795 14793 4847 14797
rect 5006 14793 5058 14797
rect 5217 14793 5269 14797
rect 6766 14791 6818 14797
rect 6977 14791 7029 14797
rect 7188 14791 7240 14797
rect 7399 14791 7451 14797
rect 7610 14791 7662 14797
rect 12333 14791 12385 14798
rect 12544 14791 12596 14798
rect 12755 14791 12807 14798
rect 12966 14791 13018 14798
rect 13177 14791 13229 14843
rect 13387 14791 13439 14843
rect 21460 15056 21512 15067
rect 21671 15056 21723 15067
rect 21882 15056 21934 15067
rect 22093 15056 22097 15067
rect 22097 15056 22145 15067
rect 23899 15274 23951 15326
rect 24110 15309 24162 15326
rect 24321 15309 24373 15326
rect 24110 15274 24122 15309
rect 24122 15274 24162 15309
rect 24321 15274 24326 15309
rect 24326 15274 24373 15309
rect 24532 15274 24584 15326
rect 24742 15309 24794 15326
rect 24953 15309 25005 15326
rect 24742 15274 24754 15309
rect 24754 15274 24794 15309
rect 24953 15274 24958 15309
rect 24958 15274 25005 15309
rect 25164 15274 25216 15326
rect 25375 15309 25427 15326
rect 25586 15309 25638 15326
rect 25375 15274 25387 15309
rect 25387 15274 25427 15309
rect 25586 15274 25591 15309
rect 25591 15274 25638 15309
rect 26178 15274 26230 15326
rect 26389 15274 26441 15326
rect 26601 15323 26653 15326
rect 26601 15277 26602 15323
rect 26602 15277 26648 15323
rect 26648 15277 26653 15323
rect 26601 15274 26653 15277
rect 26812 15274 26864 15326
rect 27338 15274 27390 15326
rect 27549 15274 27601 15326
rect 23899 15056 23951 15108
rect 24110 15100 24122 15108
rect 24122 15100 24162 15108
rect 24321 15100 24326 15108
rect 24326 15100 24373 15108
rect 24110 15056 24162 15100
rect 24321 15056 24373 15100
rect 24532 15056 24584 15108
rect 24742 15100 24754 15108
rect 24754 15100 24794 15108
rect 24953 15100 24958 15108
rect 24958 15100 25005 15108
rect 24742 15056 24794 15100
rect 24953 15056 25005 15100
rect 25164 15056 25216 15108
rect 25375 15100 25387 15108
rect 25387 15100 25427 15108
rect 25586 15100 25591 15108
rect 25591 15100 25638 15108
rect 25375 15056 25427 15100
rect 25586 15056 25638 15100
rect 20151 14797 20203 14843
rect 20362 14797 20376 14843
rect 20376 14797 20414 14843
rect 20573 14797 20582 14843
rect 20582 14797 20625 14843
rect 20784 14797 20788 14843
rect 20788 14797 20834 14843
rect 20834 14797 20836 14843
rect 22404 14797 22406 14843
rect 22406 14797 22456 14843
rect 20151 14791 20203 14797
rect 20362 14791 20414 14797
rect 20573 14791 20625 14797
rect 20784 14791 20836 14797
rect 22404 14791 22456 14797
rect 22615 14791 22667 14843
rect 22826 14797 22875 14843
rect 22875 14797 22878 14843
rect 23037 14797 23081 14843
rect 23081 14797 23089 14843
rect 23248 14797 23287 14843
rect 23287 14797 23300 14843
rect 23899 14839 23951 14891
rect 24110 14839 24162 14891
rect 24321 14839 24373 14891
rect 24532 14839 24584 14891
rect 24742 14839 24794 14891
rect 24953 14839 25005 14891
rect 25164 14839 25216 14891
rect 25375 14839 25427 14891
rect 25586 14839 25638 14891
rect 22826 14791 22878 14797
rect 23037 14791 23089 14797
rect 23248 14791 23300 14797
rect 905 14374 957 14426
rect 1116 14423 1168 14426
rect 1116 14377 1121 14423
rect 1121 14377 1167 14423
rect 1167 14377 1168 14423
rect 1116 14374 1168 14377
rect 1328 14374 1380 14426
rect 1539 14374 1591 14426
rect 168 13523 220 13526
rect 168 13477 179 13523
rect 179 13477 220 13523
rect 168 13474 220 13477
rect 379 13474 431 13526
rect 905 13474 957 13526
rect 1116 13523 1168 13526
rect 1116 13477 1121 13523
rect 1121 13477 1167 13523
rect 1167 13477 1168 13523
rect 1116 13474 1168 13477
rect 1328 13474 1380 13526
rect 1539 13474 1591 13526
rect 905 12574 957 12626
rect 1116 12623 1168 12626
rect 1116 12577 1121 12623
rect 1121 12577 1167 12623
rect 1167 12577 1168 12623
rect 1116 12574 1168 12577
rect 1328 12574 1380 12626
rect 1539 12574 1591 12626
rect 168 11723 220 11726
rect 168 11677 179 11723
rect 179 11677 220 11723
rect 168 11674 220 11677
rect 379 11674 431 11726
rect 905 11674 957 11726
rect 1116 11723 1168 11726
rect 1116 11677 1121 11723
rect 1121 11677 1167 11723
rect 1167 11677 1168 11723
rect 1116 11674 1168 11677
rect 1328 11674 1380 11726
rect 1539 11674 1591 11726
rect 905 10774 957 10826
rect 1116 10823 1168 10826
rect 1116 10777 1121 10823
rect 1121 10777 1167 10823
rect 1167 10777 1168 10823
rect 1116 10774 1168 10777
rect 1328 10774 1380 10826
rect 1539 10774 1591 10826
rect 168 9923 220 9926
rect 168 9877 179 9923
rect 179 9877 220 9923
rect 168 9874 220 9877
rect 379 9874 431 9926
rect 905 9874 957 9926
rect 1116 9923 1168 9926
rect 1116 9877 1121 9923
rect 1121 9877 1167 9923
rect 1167 9877 1168 9923
rect 1116 9874 1168 9877
rect 1328 9874 1380 9926
rect 1539 9874 1591 9926
rect 905 8974 957 9026
rect 1116 9023 1168 9026
rect 1116 8977 1121 9023
rect 1121 8977 1167 9023
rect 1167 8977 1168 9023
rect 1116 8974 1168 8977
rect 1328 8974 1380 9026
rect 1539 8974 1591 9026
rect 168 8123 220 8126
rect 168 8077 179 8123
rect 179 8077 220 8123
rect 168 8074 220 8077
rect 379 8074 431 8126
rect 905 8074 957 8126
rect 1116 8123 1168 8126
rect 1116 8077 1121 8123
rect 1121 8077 1167 8123
rect 1167 8077 1168 8123
rect 1116 8074 1168 8077
rect 1328 8074 1380 8126
rect 1539 8074 1591 8126
rect 905 7174 957 7226
rect 1116 7223 1168 7226
rect 1116 7177 1121 7223
rect 1121 7177 1167 7223
rect 1167 7177 1168 7223
rect 1116 7174 1168 7177
rect 1328 7174 1380 7226
rect 1539 7174 1591 7226
rect 168 6323 220 6326
rect 168 6277 179 6323
rect 179 6277 220 6323
rect 168 6274 220 6277
rect 379 6274 431 6326
rect 905 6274 957 6326
rect 1116 6323 1168 6326
rect 1116 6277 1121 6323
rect 1121 6277 1167 6323
rect 1167 6277 1168 6323
rect 1116 6274 1168 6277
rect 1328 6274 1380 6326
rect 1539 6274 1591 6326
rect 905 5374 957 5426
rect 1116 5423 1168 5426
rect 1116 5377 1121 5423
rect 1121 5377 1167 5423
rect 1167 5377 1168 5423
rect 1116 5374 1168 5377
rect 1328 5374 1380 5426
rect 1539 5374 1591 5426
rect 168 4523 220 4526
rect 168 4477 179 4523
rect 179 4477 220 4523
rect 168 4474 220 4477
rect 379 4474 431 4526
rect 905 4474 957 4526
rect 1116 4523 1168 4526
rect 1116 4477 1121 4523
rect 1121 4477 1167 4523
rect 1167 4477 1168 4523
rect 1116 4474 1168 4477
rect 1328 4474 1380 4526
rect 1539 4474 1591 4526
rect 905 3574 957 3626
rect 1116 3623 1168 3626
rect 1116 3577 1121 3623
rect 1121 3577 1167 3623
rect 1167 3577 1168 3623
rect 1116 3574 1168 3577
rect 1328 3574 1380 3626
rect 1539 3574 1591 3626
rect 168 2723 220 2726
rect 168 2677 179 2723
rect 179 2677 220 2723
rect 168 2674 220 2677
rect 379 2674 431 2726
rect 905 2674 957 2726
rect 1116 2723 1168 2726
rect 1116 2677 1121 2723
rect 1121 2677 1167 2723
rect 1167 2677 1168 2723
rect 1116 2674 1168 2677
rect 1328 2674 1380 2726
rect 1539 2674 1591 2726
rect 905 1774 957 1826
rect 1116 1823 1168 1826
rect 1116 1777 1121 1823
rect 1121 1777 1167 1823
rect 1167 1777 1168 1823
rect 1116 1774 1168 1777
rect 1328 1774 1380 1826
rect 1539 1774 1591 1826
rect 168 923 220 926
rect 168 877 179 923
rect 179 877 220 923
rect 168 874 220 877
rect 379 874 431 926
rect 905 874 957 926
rect 1116 923 1168 926
rect 1116 877 1121 923
rect 1121 877 1167 923
rect 1167 877 1168 923
rect 1116 874 1168 877
rect 1328 874 1380 926
rect 1539 874 1591 926
rect 905 -26 957 26
rect 1116 23 1168 26
rect 1116 -23 1121 23
rect 1121 -23 1167 23
rect 1167 -23 1168 23
rect 1116 -26 1168 -23
rect 1328 -26 1380 26
rect 1539 -26 1591 26
rect 26178 14374 26230 14426
rect 26389 14374 26441 14426
rect 26601 14423 26653 14426
rect 26601 14377 26602 14423
rect 26602 14377 26648 14423
rect 26648 14377 26653 14423
rect 26601 14374 26653 14377
rect 26812 14374 26864 14426
rect 26178 13474 26230 13526
rect 26389 13474 26441 13526
rect 26601 13523 26653 13526
rect 26601 13477 26602 13523
rect 26602 13477 26648 13523
rect 26648 13477 26653 13523
rect 26601 13474 26653 13477
rect 26812 13474 26864 13526
rect 27338 13474 27390 13526
rect 27549 13523 27601 13526
rect 27549 13477 27590 13523
rect 27590 13477 27601 13523
rect 27549 13474 27601 13477
rect 26178 12574 26230 12626
rect 26389 12574 26441 12626
rect 26601 12623 26653 12626
rect 26601 12577 26602 12623
rect 26602 12577 26648 12623
rect 26648 12577 26653 12623
rect 26601 12574 26653 12577
rect 26812 12574 26864 12626
rect 26178 11674 26230 11726
rect 26389 11674 26441 11726
rect 26601 11723 26653 11726
rect 26601 11677 26602 11723
rect 26602 11677 26648 11723
rect 26648 11677 26653 11723
rect 26601 11674 26653 11677
rect 26812 11674 26864 11726
rect 27338 11674 27390 11726
rect 27549 11723 27601 11726
rect 27549 11677 27590 11723
rect 27590 11677 27601 11723
rect 27549 11674 27601 11677
rect 26178 10774 26230 10826
rect 26389 10774 26441 10826
rect 26601 10823 26653 10826
rect 26601 10777 26602 10823
rect 26602 10777 26648 10823
rect 26648 10777 26653 10823
rect 26601 10774 26653 10777
rect 26812 10774 26864 10826
rect 26178 9874 26230 9926
rect 26389 9874 26441 9926
rect 26601 9923 26653 9926
rect 26601 9877 26602 9923
rect 26602 9877 26648 9923
rect 26648 9877 26653 9923
rect 26601 9874 26653 9877
rect 26812 9874 26864 9926
rect 27338 9874 27390 9926
rect 27549 9923 27601 9926
rect 27549 9877 27590 9923
rect 27590 9877 27601 9923
rect 27549 9874 27601 9877
rect 26178 8974 26230 9026
rect 26389 8974 26441 9026
rect 26601 9023 26653 9026
rect 26601 8977 26602 9023
rect 26602 8977 26648 9023
rect 26648 8977 26653 9023
rect 26601 8974 26653 8977
rect 26812 8974 26864 9026
rect 26178 8074 26230 8126
rect 26389 8074 26441 8126
rect 26601 8123 26653 8126
rect 26601 8077 26602 8123
rect 26602 8077 26648 8123
rect 26648 8077 26653 8123
rect 26601 8074 26653 8077
rect 26812 8074 26864 8126
rect 27338 8074 27390 8126
rect 27549 8123 27601 8126
rect 27549 8077 27590 8123
rect 27590 8077 27601 8123
rect 27549 8074 27601 8077
rect 26178 7174 26230 7226
rect 26389 7174 26441 7226
rect 26601 7223 26653 7226
rect 26601 7177 26602 7223
rect 26602 7177 26648 7223
rect 26648 7177 26653 7223
rect 26601 7174 26653 7177
rect 26812 7174 26864 7226
rect 26178 6274 26230 6326
rect 26389 6274 26441 6326
rect 26601 6323 26653 6326
rect 26601 6277 26602 6323
rect 26602 6277 26648 6323
rect 26648 6277 26653 6323
rect 26601 6274 26653 6277
rect 26812 6274 26864 6326
rect 27338 6274 27390 6326
rect 27549 6323 27601 6326
rect 27549 6277 27590 6323
rect 27590 6277 27601 6323
rect 27549 6274 27601 6277
rect 26178 5374 26230 5426
rect 26389 5374 26441 5426
rect 26601 5423 26653 5426
rect 26601 5377 26602 5423
rect 26602 5377 26648 5423
rect 26648 5377 26653 5423
rect 26601 5374 26653 5377
rect 26812 5374 26864 5426
rect 26178 4474 26230 4526
rect 26389 4474 26441 4526
rect 26601 4523 26653 4526
rect 26601 4477 26602 4523
rect 26602 4477 26648 4523
rect 26648 4477 26653 4523
rect 26601 4474 26653 4477
rect 26812 4474 26864 4526
rect 27338 4474 27390 4526
rect 27549 4523 27601 4526
rect 27549 4477 27590 4523
rect 27590 4477 27601 4523
rect 27549 4474 27601 4477
rect 26178 3574 26230 3626
rect 26389 3574 26441 3626
rect 26601 3623 26653 3626
rect 26601 3577 26602 3623
rect 26602 3577 26648 3623
rect 26648 3577 26653 3623
rect 26601 3574 26653 3577
rect 26812 3574 26864 3626
rect 26178 2674 26230 2726
rect 26389 2674 26441 2726
rect 26601 2723 26653 2726
rect 26601 2677 26602 2723
rect 26602 2677 26648 2723
rect 26648 2677 26653 2723
rect 26601 2674 26653 2677
rect 26812 2674 26864 2726
rect 27338 2674 27390 2726
rect 27549 2723 27601 2726
rect 27549 2677 27590 2723
rect 27590 2677 27601 2723
rect 27549 2674 27601 2677
rect 26178 1774 26230 1826
rect 26389 1774 26441 1826
rect 26601 1823 26653 1826
rect 26601 1777 26602 1823
rect 26602 1777 26648 1823
rect 26648 1777 26653 1823
rect 26601 1774 26653 1777
rect 26812 1774 26864 1826
rect 26178 874 26230 926
rect 26389 874 26441 926
rect 26601 923 26653 926
rect 26601 877 26602 923
rect 26602 877 26648 923
rect 26648 877 26653 923
rect 26601 874 26653 877
rect 26812 874 26864 926
rect 27338 874 27390 926
rect 27549 923 27601 926
rect 27549 877 27590 923
rect 27590 877 27601 923
rect 27549 874 27601 877
rect 26178 -26 26230 26
rect 26389 -26 26441 26
rect 26601 23 26653 26
rect 26601 -23 26602 23
rect 26602 -23 26648 23
rect 26648 -23 26653 23
rect 26601 -26 26653 -23
rect 26812 -26 26864 26
<< metal2 >>
rect 129 15328 469 15367
rect 129 15272 166 15328
rect 222 15272 377 15328
rect 433 15272 469 15328
rect 129 15233 469 15272
rect 808 15326 1688 15401
rect 808 15274 905 15326
rect 957 15274 1116 15326
rect 1168 15274 1328 15326
rect 1380 15274 1539 15326
rect 1591 15274 1688 15326
rect 808 14428 1688 15274
rect 808 14372 903 14428
rect 959 14372 1114 14428
rect 1170 14372 1326 14428
rect 1382 14372 1537 14428
rect 1593 14372 1688 14428
rect 2092 15326 4211 15476
rect 2092 15274 2130 15326
rect 2182 15274 2341 15326
rect 2393 15274 2552 15326
rect 2604 15274 2763 15326
rect 2815 15274 2974 15326
rect 3026 15274 3184 15326
rect 3236 15274 3395 15326
rect 3447 15274 3606 15326
rect 3658 15274 3817 15326
rect 3869 15274 4211 15326
rect 2092 15108 4211 15274
rect 2092 15056 2130 15108
rect 2182 15056 2341 15108
rect 2393 15056 2552 15108
rect 2604 15056 2763 15108
rect 2815 15056 2974 15108
rect 3026 15056 3184 15108
rect 3236 15056 3395 15108
rect 3447 15056 3606 15108
rect 3658 15056 3817 15108
rect 3869 15056 4211 15108
rect 2092 14891 4211 15056
rect 2092 14839 2130 14891
rect 2182 14839 2341 14891
rect 2393 14839 2552 14891
rect 2604 14839 2763 14891
rect 2815 14839 2974 14891
rect 3026 14839 3184 14891
rect 3236 14839 3395 14891
rect 3447 14839 3606 14891
rect 3658 14839 3817 14891
rect 3869 14839 4211 14891
rect 5550 15328 6347 15401
rect 5550 15272 5611 15328
rect 5667 15272 5822 15328
rect 5878 15272 6033 15328
rect 6089 15272 6244 15328
rect 6300 15272 6347 15328
rect 5550 15108 6347 15272
rect 5550 15056 5613 15108
rect 5665 15056 5824 15108
rect 5876 15056 6035 15108
rect 6087 15056 6246 15108
rect 6298 15056 6347 15108
rect 2092 14413 4211 14839
rect 4334 14847 5307 14886
rect 4334 14791 4371 14847
rect 4427 14791 4582 14847
rect 4638 14791 4793 14847
rect 4849 14791 5004 14847
rect 5060 14791 5215 14847
rect 5271 14791 5307 14847
rect 4334 14753 5307 14791
rect 5550 14413 6347 15056
rect 6451 15306 7738 15401
rect 6451 15254 6766 15306
rect 6818 15254 6977 15306
rect 7029 15254 7188 15306
rect 7240 15254 7399 15306
rect 7451 15254 7610 15306
rect 7662 15254 7738 15306
rect 6451 14843 7738 15254
rect 6451 14791 6766 14843
rect 6818 14791 6977 14843
rect 7029 14791 7188 14843
rect 7240 14791 7399 14843
rect 7451 14791 7610 14843
rect 7662 14791 7738 14843
rect 6451 14413 7738 14791
rect 8186 14845 9066 14884
rect 8186 14789 8222 14845
rect 8278 14789 8433 14845
rect 8489 14789 8644 14845
rect 8700 14789 8855 14845
rect 8911 14789 9066 14845
rect 8186 14413 9066 14789
rect 9591 14413 10186 15401
rect 10276 15074 10941 15401
rect 10276 15022 10376 15074
rect 10428 15022 10587 15074
rect 10639 15022 10798 15074
rect 10850 15022 10941 15074
rect 10276 14413 10941 15022
rect 11537 15331 11846 15401
rect 13994 15378 14545 15419
rect 11537 15328 11575 15331
rect 11627 15328 11755 15331
rect 11807 15328 11846 15331
rect 11537 15272 11573 15328
rect 11629 15272 11753 15328
rect 11809 15272 11846 15328
rect 11537 15113 11846 15272
rect 13531 15317 13871 15358
rect 13531 15265 13569 15317
rect 13621 15265 13781 15317
rect 13833 15265 13871 15317
rect 13531 15224 13871 15265
rect 13994 15326 14033 15378
rect 14085 15326 14244 15378
rect 14296 15326 14455 15378
rect 14507 15326 14545 15378
rect 11537 15061 11575 15113
rect 11627 15061 11755 15113
rect 11807 15061 11846 15113
rect 11537 14413 11846 15061
rect 12294 14845 13478 14884
rect 12294 14789 12331 14845
rect 12387 14789 12542 14845
rect 12598 14789 12753 14845
rect 12809 14789 12964 14845
rect 13020 14789 13175 14845
rect 13231 14789 13385 14845
rect 13441 14789 13478 14845
rect 12294 14750 13478 14789
rect 13994 14838 14545 15326
rect 13994 14782 14031 14838
rect 14087 14782 14242 14838
rect 14298 14782 14453 14838
rect 14509 14782 14545 14838
rect 13994 14744 14545 14782
rect 15026 15378 15887 15419
rect 15026 15326 15100 15378
rect 15152 15326 15311 15378
rect 15363 15326 15522 15378
rect 15574 15326 15733 15378
rect 15785 15326 15887 15378
rect 12040 14428 12639 14564
rect 129 13528 469 13567
rect 129 13526 377 13528
rect 129 13474 168 13526
rect 220 13474 377 13526
rect 129 13472 377 13474
rect 433 13472 469 13528
rect 129 13433 469 13472
rect 808 13526 1688 14372
rect 12040 14372 12100 14428
rect 12156 14372 12311 14428
rect 12367 14372 12522 14428
rect 12578 14372 12639 14428
rect 15026 14413 15887 15326
rect 20112 15306 21313 15401
rect 20112 15254 20151 15306
rect 20203 15254 20362 15306
rect 20414 15254 20573 15306
rect 20625 15254 20784 15306
rect 20836 15254 21313 15306
rect 20112 14843 21313 15254
rect 20112 14791 20151 14843
rect 20203 14791 20362 14843
rect 20414 14791 20573 14843
rect 20625 14791 20784 14843
rect 20836 14791 21313 14843
rect 20112 14413 21313 14791
rect 21421 15328 22236 15419
rect 21421 15272 21458 15328
rect 21514 15272 21669 15328
rect 21725 15272 21880 15328
rect 21936 15272 22091 15328
rect 22147 15272 22236 15328
rect 21421 15108 22236 15272
rect 21421 15056 21460 15108
rect 21512 15056 21671 15108
rect 21723 15056 21882 15108
rect 21934 15056 22093 15108
rect 22145 15056 22236 15108
rect 21421 14413 22236 15056
rect 23549 15326 25677 15476
rect 23549 15274 23899 15326
rect 23951 15274 24110 15326
rect 24162 15274 24321 15326
rect 24373 15274 24532 15326
rect 24584 15274 24742 15326
rect 24794 15274 24953 15326
rect 25005 15274 25164 15326
rect 25216 15274 25375 15326
rect 25427 15274 25586 15326
rect 25638 15274 25677 15326
rect 23549 15108 25677 15274
rect 23549 15056 23899 15108
rect 23951 15056 24110 15108
rect 24162 15056 24321 15108
rect 24373 15056 24532 15108
rect 24584 15056 24742 15108
rect 24794 15056 24953 15108
rect 25005 15056 25164 15108
rect 25216 15056 25375 15108
rect 25427 15056 25586 15108
rect 25638 15056 25677 15108
rect 23549 14891 25677 15056
rect 22365 14845 23338 14884
rect 22365 14789 22402 14845
rect 22458 14789 22613 14845
rect 22669 14789 22824 14845
rect 22880 14789 23035 14845
rect 23091 14789 23246 14845
rect 23302 14789 23338 14845
rect 22365 14751 23338 14789
rect 23549 14839 23899 14891
rect 23951 14839 24110 14891
rect 24162 14839 24321 14891
rect 24373 14839 24532 14891
rect 24584 14839 24742 14891
rect 24794 14839 24953 14891
rect 25005 14839 25164 14891
rect 25216 14839 25375 14891
rect 25427 14839 25586 14891
rect 25638 14839 25677 14891
rect 23549 14413 25677 14839
rect 26081 15326 26961 15401
rect 26081 15274 26178 15326
rect 26230 15274 26389 15326
rect 26441 15274 26601 15326
rect 26653 15274 26812 15326
rect 26864 15274 26961 15326
rect 26081 14428 26961 15274
rect 27300 15328 27640 15367
rect 27300 15272 27336 15328
rect 27392 15272 27547 15328
rect 27603 15272 27640 15328
rect 27300 15233 27640 15272
rect 12040 14299 12639 14372
rect 26081 14372 26176 14428
rect 26232 14372 26387 14428
rect 26443 14372 26599 14428
rect 26655 14372 26810 14428
rect 26866 14372 26961 14428
rect 808 13474 905 13526
rect 957 13474 1116 13526
rect 1168 13474 1328 13526
rect 1380 13474 1539 13526
rect 1591 13474 1688 13526
rect 808 12628 1688 13474
rect 808 12572 903 12628
rect 959 12572 1114 12628
rect 1170 12572 1326 12628
rect 1382 12572 1537 12628
rect 1593 12572 1688 12628
rect 129 11728 469 11767
rect 129 11726 377 11728
rect 129 11674 168 11726
rect 220 11674 377 11726
rect 129 11672 377 11674
rect 433 11672 469 11728
rect 129 11633 469 11672
rect 808 11726 1688 12572
rect 808 11674 905 11726
rect 957 11674 1116 11726
rect 1168 11674 1328 11726
rect 1380 11674 1539 11726
rect 1591 11674 1688 11726
rect 808 10828 1688 11674
rect 808 10772 903 10828
rect 959 10772 1114 10828
rect 1170 10772 1326 10828
rect 1382 10772 1537 10828
rect 1593 10772 1688 10828
rect 129 9928 469 9967
rect 129 9926 377 9928
rect 129 9874 168 9926
rect 220 9874 377 9926
rect 129 9872 377 9874
rect 433 9872 469 9928
rect 129 9833 469 9872
rect 808 9926 1688 10772
rect 808 9874 905 9926
rect 957 9874 1116 9926
rect 1168 9874 1328 9926
rect 1380 9874 1539 9926
rect 1591 9874 1688 9926
rect 808 9028 1688 9874
rect 808 8972 903 9028
rect 959 8972 1114 9028
rect 1170 8972 1326 9028
rect 1382 8972 1537 9028
rect 1593 8972 1688 9028
rect 129 8128 469 8167
rect 129 8126 377 8128
rect 129 8074 168 8126
rect 220 8074 377 8126
rect 129 8072 377 8074
rect 433 8072 469 8128
rect 129 8033 469 8072
rect 808 8126 1688 8972
rect 808 8074 905 8126
rect 957 8074 1116 8126
rect 1168 8074 1328 8126
rect 1380 8074 1539 8126
rect 1591 8074 1688 8126
rect 808 7228 1688 8074
rect 808 7172 903 7228
rect 959 7172 1114 7228
rect 1170 7172 1326 7228
rect 1382 7172 1537 7228
rect 1593 7172 1688 7228
rect 129 6328 469 6367
rect 129 6326 377 6328
rect 129 6274 168 6326
rect 220 6274 377 6326
rect 129 6272 377 6274
rect 433 6272 469 6328
rect 129 6233 469 6272
rect 808 6326 1688 7172
rect 808 6274 905 6326
rect 957 6274 1116 6326
rect 1168 6274 1328 6326
rect 1380 6274 1539 6326
rect 1591 6274 1688 6326
rect 808 5428 1688 6274
rect 808 5372 903 5428
rect 959 5372 1114 5428
rect 1170 5372 1326 5428
rect 1382 5372 1537 5428
rect 1593 5372 1688 5428
rect 129 4528 469 4567
rect 129 4526 377 4528
rect 129 4474 168 4526
rect 220 4474 377 4526
rect 129 4472 377 4474
rect 433 4472 469 4528
rect 129 4433 469 4472
rect 808 4526 1688 5372
rect 808 4474 905 4526
rect 957 4474 1116 4526
rect 1168 4474 1328 4526
rect 1380 4474 1539 4526
rect 1591 4474 1688 4526
rect 808 3628 1688 4474
rect 808 3572 903 3628
rect 959 3572 1114 3628
rect 1170 3572 1326 3628
rect 1382 3572 1537 3628
rect 1593 3572 1688 3628
rect 129 2728 469 2767
rect 129 2726 377 2728
rect 129 2674 168 2726
rect 220 2674 377 2726
rect 129 2672 377 2674
rect 433 2672 469 2728
rect 129 2633 469 2672
rect 808 2726 1688 3572
rect 808 2674 905 2726
rect 957 2674 1116 2726
rect 1168 2674 1328 2726
rect 1380 2674 1539 2726
rect 1591 2674 1688 2726
rect 808 1828 1688 2674
rect 808 1772 903 1828
rect 959 1772 1114 1828
rect 1170 1772 1326 1828
rect 1382 1772 1537 1828
rect 1593 1772 1688 1828
rect 129 928 469 967
rect 129 926 377 928
rect 129 874 168 926
rect 220 874 377 926
rect 129 872 377 874
rect 433 872 469 928
rect 129 833 469 872
rect 808 926 1688 1772
rect 808 874 905 926
rect 957 874 1116 926
rect 1168 874 1328 926
rect 1380 874 1539 926
rect 1591 874 1688 926
rect 808 28 1688 874
rect 26081 13526 26961 14372
rect 26081 13474 26178 13526
rect 26230 13474 26389 13526
rect 26441 13474 26601 13526
rect 26653 13474 26812 13526
rect 26864 13474 26961 13526
rect 26081 12628 26961 13474
rect 27300 13528 27640 13567
rect 27300 13472 27336 13528
rect 27392 13526 27640 13528
rect 27392 13474 27549 13526
rect 27601 13474 27640 13526
rect 27392 13472 27640 13474
rect 27300 13433 27640 13472
rect 26081 12572 26176 12628
rect 26232 12572 26387 12628
rect 26443 12572 26599 12628
rect 26655 12572 26810 12628
rect 26866 12572 26961 12628
rect 26081 11726 26961 12572
rect 26081 11674 26178 11726
rect 26230 11674 26389 11726
rect 26441 11674 26601 11726
rect 26653 11674 26812 11726
rect 26864 11674 26961 11726
rect 26081 10828 26961 11674
rect 27300 11728 27640 11767
rect 27300 11672 27336 11728
rect 27392 11726 27640 11728
rect 27392 11674 27549 11726
rect 27601 11674 27640 11726
rect 27392 11672 27640 11674
rect 27300 11633 27640 11672
rect 26081 10772 26176 10828
rect 26232 10772 26387 10828
rect 26443 10772 26599 10828
rect 26655 10772 26810 10828
rect 26866 10772 26961 10828
rect 26081 9926 26961 10772
rect 26081 9874 26178 9926
rect 26230 9874 26389 9926
rect 26441 9874 26601 9926
rect 26653 9874 26812 9926
rect 26864 9874 26961 9926
rect 26081 9028 26961 9874
rect 27300 9928 27640 9967
rect 27300 9872 27336 9928
rect 27392 9926 27640 9928
rect 27392 9874 27549 9926
rect 27601 9874 27640 9926
rect 27392 9872 27640 9874
rect 27300 9833 27640 9872
rect 26081 8972 26176 9028
rect 26232 8972 26387 9028
rect 26443 8972 26599 9028
rect 26655 8972 26810 9028
rect 26866 8972 26961 9028
rect 26081 8126 26961 8972
rect 26081 8074 26178 8126
rect 26230 8074 26389 8126
rect 26441 8074 26601 8126
rect 26653 8074 26812 8126
rect 26864 8074 26961 8126
rect 26081 7228 26961 8074
rect 27300 8128 27640 8167
rect 27300 8072 27336 8128
rect 27392 8126 27640 8128
rect 27392 8074 27549 8126
rect 27601 8074 27640 8126
rect 27392 8072 27640 8074
rect 27300 8033 27640 8072
rect 26081 7172 26176 7228
rect 26232 7172 26387 7228
rect 26443 7172 26599 7228
rect 26655 7172 26810 7228
rect 26866 7172 26961 7228
rect 26081 6326 26961 7172
rect 26081 6274 26178 6326
rect 26230 6274 26389 6326
rect 26441 6274 26601 6326
rect 26653 6274 26812 6326
rect 26864 6274 26961 6326
rect 26081 5428 26961 6274
rect 27300 6328 27640 6367
rect 27300 6272 27336 6328
rect 27392 6326 27640 6328
rect 27392 6274 27549 6326
rect 27601 6274 27640 6326
rect 27392 6272 27640 6274
rect 27300 6233 27640 6272
rect 26081 5372 26176 5428
rect 26232 5372 26387 5428
rect 26443 5372 26599 5428
rect 26655 5372 26810 5428
rect 26866 5372 26961 5428
rect 26081 4526 26961 5372
rect 26081 4474 26178 4526
rect 26230 4474 26389 4526
rect 26441 4474 26601 4526
rect 26653 4474 26812 4526
rect 26864 4474 26961 4526
rect 26081 3628 26961 4474
rect 27300 4528 27640 4567
rect 27300 4472 27336 4528
rect 27392 4526 27640 4528
rect 27392 4474 27549 4526
rect 27601 4474 27640 4526
rect 27392 4472 27640 4474
rect 27300 4433 27640 4472
rect 26081 3572 26176 3628
rect 26232 3572 26387 3628
rect 26443 3572 26599 3628
rect 26655 3572 26810 3628
rect 26866 3572 26961 3628
rect 26081 2726 26961 3572
rect 26081 2674 26178 2726
rect 26230 2674 26389 2726
rect 26441 2674 26601 2726
rect 26653 2674 26812 2726
rect 26864 2674 26961 2726
rect 26081 1828 26961 2674
rect 27300 2728 27640 2767
rect 27300 2672 27336 2728
rect 27392 2726 27640 2728
rect 27392 2674 27549 2726
rect 27601 2674 27640 2726
rect 27392 2672 27640 2674
rect 27300 2633 27640 2672
rect 26081 1772 26176 1828
rect 26232 1772 26387 1828
rect 26443 1772 26599 1828
rect 26655 1772 26810 1828
rect 26866 1772 26961 1828
rect 26081 926 26961 1772
rect 26081 874 26178 926
rect 26230 874 26389 926
rect 26441 874 26601 926
rect 26653 874 26812 926
rect 26864 874 26961 926
rect 808 -28 903 28
rect 959 -28 1114 28
rect 1170 -28 1326 28
rect 1382 -28 1537 28
rect 1593 -28 1688 28
rect 8561 -21 8691 112
rect 26081 28 26961 874
rect 27300 928 27640 967
rect 27300 872 27336 928
rect 27392 926 27640 928
rect 27392 874 27549 926
rect 27601 874 27640 926
rect 27392 872 27640 874
rect 27300 833 27640 872
rect 808 -100 1688 -28
rect 26081 -28 26176 28
rect 26232 -28 26387 28
rect 26443 -28 26599 28
rect 26655 -28 26810 28
rect 26866 -28 26961 28
rect 12841 -164 12971 -31
rect 13219 -164 13348 -31
rect 13597 -164 13726 -31
rect 13974 -164 14104 -31
rect 14352 -164 14481 -31
rect 14730 -164 14859 -31
rect 16882 -164 17011 -31
rect 17260 -164 17389 -31
rect 17637 -164 17767 -31
rect 18015 -164 18144 -31
rect 18393 -164 18522 -31
rect 18770 -164 18900 -31
rect 19148 -164 19277 -31
rect 19526 -164 19655 -31
rect 26081 -100 26961 -28
<< via2 >>
rect 166 15326 222 15328
rect 166 15274 168 15326
rect 168 15274 220 15326
rect 220 15274 222 15326
rect 166 15272 222 15274
rect 377 15326 433 15328
rect 377 15274 379 15326
rect 379 15274 431 15326
rect 431 15274 433 15326
rect 377 15272 433 15274
rect 903 14426 959 14428
rect 903 14374 905 14426
rect 905 14374 957 14426
rect 957 14374 959 14426
rect 903 14372 959 14374
rect 1114 14426 1170 14428
rect 1114 14374 1116 14426
rect 1116 14374 1168 14426
rect 1168 14374 1170 14426
rect 1114 14372 1170 14374
rect 1326 14426 1382 14428
rect 1326 14374 1328 14426
rect 1328 14374 1380 14426
rect 1380 14374 1382 14426
rect 1326 14372 1382 14374
rect 1537 14426 1593 14428
rect 1537 14374 1539 14426
rect 1539 14374 1591 14426
rect 1591 14374 1593 14426
rect 1537 14372 1593 14374
rect 5611 15326 5667 15328
rect 5611 15274 5613 15326
rect 5613 15274 5665 15326
rect 5665 15274 5667 15326
rect 5611 15272 5667 15274
rect 5822 15326 5878 15328
rect 5822 15274 5824 15326
rect 5824 15274 5876 15326
rect 5876 15274 5878 15326
rect 5822 15272 5878 15274
rect 6033 15326 6089 15328
rect 6033 15274 6035 15326
rect 6035 15274 6087 15326
rect 6087 15274 6089 15326
rect 6033 15272 6089 15274
rect 6244 15326 6300 15328
rect 6244 15274 6246 15326
rect 6246 15274 6298 15326
rect 6298 15274 6300 15326
rect 6244 15272 6300 15274
rect 4371 14845 4427 14847
rect 4371 14793 4373 14845
rect 4373 14793 4425 14845
rect 4425 14793 4427 14845
rect 4371 14791 4427 14793
rect 4582 14845 4638 14847
rect 4582 14793 4584 14845
rect 4584 14793 4636 14845
rect 4636 14793 4638 14845
rect 4582 14791 4638 14793
rect 4793 14845 4849 14847
rect 4793 14793 4795 14845
rect 4795 14793 4847 14845
rect 4847 14793 4849 14845
rect 4793 14791 4849 14793
rect 5004 14845 5060 14847
rect 5004 14793 5006 14845
rect 5006 14793 5058 14845
rect 5058 14793 5060 14845
rect 5004 14791 5060 14793
rect 5215 14845 5271 14847
rect 5215 14793 5217 14845
rect 5217 14793 5269 14845
rect 5269 14793 5271 14845
rect 5215 14791 5271 14793
rect 8222 14789 8278 14845
rect 8433 14789 8489 14845
rect 8644 14789 8700 14845
rect 8855 14789 8911 14845
rect 11573 15279 11575 15328
rect 11575 15279 11627 15328
rect 11627 15279 11629 15328
rect 11573 15272 11629 15279
rect 11753 15279 11755 15328
rect 11755 15279 11807 15328
rect 11807 15279 11809 15328
rect 11753 15272 11809 15279
rect 12331 14843 12387 14845
rect 12331 14791 12333 14843
rect 12333 14791 12385 14843
rect 12385 14791 12387 14843
rect 12331 14789 12387 14791
rect 12542 14843 12598 14845
rect 12542 14791 12544 14843
rect 12544 14791 12596 14843
rect 12596 14791 12598 14843
rect 12542 14789 12598 14791
rect 12753 14843 12809 14845
rect 12753 14791 12755 14843
rect 12755 14791 12807 14843
rect 12807 14791 12809 14843
rect 12753 14789 12809 14791
rect 12964 14843 13020 14845
rect 12964 14791 12966 14843
rect 12966 14791 13018 14843
rect 13018 14791 13020 14843
rect 12964 14789 13020 14791
rect 13175 14843 13231 14845
rect 13175 14791 13177 14843
rect 13177 14791 13229 14843
rect 13229 14791 13231 14843
rect 13175 14789 13231 14791
rect 13385 14843 13441 14845
rect 13385 14791 13387 14843
rect 13387 14791 13439 14843
rect 13439 14791 13441 14843
rect 13385 14789 13441 14791
rect 14031 14782 14087 14838
rect 14242 14782 14298 14838
rect 14453 14782 14509 14838
rect 377 13526 433 13528
rect 377 13474 379 13526
rect 379 13474 431 13526
rect 431 13474 433 13526
rect 377 13472 433 13474
rect 12100 14372 12156 14428
rect 12311 14372 12367 14428
rect 12522 14372 12578 14428
rect 21458 15326 21514 15328
rect 21458 15274 21460 15326
rect 21460 15274 21512 15326
rect 21512 15274 21514 15326
rect 21458 15272 21514 15274
rect 21669 15326 21725 15328
rect 21669 15274 21671 15326
rect 21671 15274 21723 15326
rect 21723 15274 21725 15326
rect 21669 15272 21725 15274
rect 21880 15326 21936 15328
rect 21880 15274 21882 15326
rect 21882 15274 21934 15326
rect 21934 15274 21936 15326
rect 21880 15272 21936 15274
rect 22091 15326 22147 15328
rect 22091 15274 22093 15326
rect 22093 15274 22145 15326
rect 22145 15274 22147 15326
rect 22091 15272 22147 15274
rect 22402 14843 22458 14845
rect 22402 14791 22404 14843
rect 22404 14791 22456 14843
rect 22456 14791 22458 14843
rect 22402 14789 22458 14791
rect 22613 14843 22669 14845
rect 22613 14791 22615 14843
rect 22615 14791 22667 14843
rect 22667 14791 22669 14843
rect 22613 14789 22669 14791
rect 22824 14843 22880 14845
rect 22824 14791 22826 14843
rect 22826 14791 22878 14843
rect 22878 14791 22880 14843
rect 22824 14789 22880 14791
rect 23035 14843 23091 14845
rect 23035 14791 23037 14843
rect 23037 14791 23089 14843
rect 23089 14791 23091 14843
rect 23035 14789 23091 14791
rect 23246 14843 23302 14845
rect 23246 14791 23248 14843
rect 23248 14791 23300 14843
rect 23300 14791 23302 14843
rect 23246 14789 23302 14791
rect 27336 15326 27392 15328
rect 27336 15274 27338 15326
rect 27338 15274 27390 15326
rect 27390 15274 27392 15326
rect 27336 15272 27392 15274
rect 27547 15326 27603 15328
rect 27547 15274 27549 15326
rect 27549 15274 27601 15326
rect 27601 15274 27603 15326
rect 27547 15272 27603 15274
rect 26176 14426 26232 14428
rect 26176 14374 26178 14426
rect 26178 14374 26230 14426
rect 26230 14374 26232 14426
rect 26176 14372 26232 14374
rect 26387 14426 26443 14428
rect 26387 14374 26389 14426
rect 26389 14374 26441 14426
rect 26441 14374 26443 14426
rect 26387 14372 26443 14374
rect 26599 14426 26655 14428
rect 26599 14374 26601 14426
rect 26601 14374 26653 14426
rect 26653 14374 26655 14426
rect 26599 14372 26655 14374
rect 26810 14426 26866 14428
rect 26810 14374 26812 14426
rect 26812 14374 26864 14426
rect 26864 14374 26866 14426
rect 26810 14372 26866 14374
rect 903 12626 959 12628
rect 903 12574 905 12626
rect 905 12574 957 12626
rect 957 12574 959 12626
rect 903 12572 959 12574
rect 1114 12626 1170 12628
rect 1114 12574 1116 12626
rect 1116 12574 1168 12626
rect 1168 12574 1170 12626
rect 1114 12572 1170 12574
rect 1326 12626 1382 12628
rect 1326 12574 1328 12626
rect 1328 12574 1380 12626
rect 1380 12574 1382 12626
rect 1326 12572 1382 12574
rect 1537 12626 1593 12628
rect 1537 12574 1539 12626
rect 1539 12574 1591 12626
rect 1591 12574 1593 12626
rect 1537 12572 1593 12574
rect 377 11726 433 11728
rect 377 11674 379 11726
rect 379 11674 431 11726
rect 431 11674 433 11726
rect 377 11672 433 11674
rect 903 10826 959 10828
rect 903 10774 905 10826
rect 905 10774 957 10826
rect 957 10774 959 10826
rect 903 10772 959 10774
rect 1114 10826 1170 10828
rect 1114 10774 1116 10826
rect 1116 10774 1168 10826
rect 1168 10774 1170 10826
rect 1114 10772 1170 10774
rect 1326 10826 1382 10828
rect 1326 10774 1328 10826
rect 1328 10774 1380 10826
rect 1380 10774 1382 10826
rect 1326 10772 1382 10774
rect 1537 10826 1593 10828
rect 1537 10774 1539 10826
rect 1539 10774 1591 10826
rect 1591 10774 1593 10826
rect 1537 10772 1593 10774
rect 377 9926 433 9928
rect 377 9874 379 9926
rect 379 9874 431 9926
rect 431 9874 433 9926
rect 377 9872 433 9874
rect 903 9026 959 9028
rect 903 8974 905 9026
rect 905 8974 957 9026
rect 957 8974 959 9026
rect 903 8972 959 8974
rect 1114 9026 1170 9028
rect 1114 8974 1116 9026
rect 1116 8974 1168 9026
rect 1168 8974 1170 9026
rect 1114 8972 1170 8974
rect 1326 9026 1382 9028
rect 1326 8974 1328 9026
rect 1328 8974 1380 9026
rect 1380 8974 1382 9026
rect 1326 8972 1382 8974
rect 1537 9026 1593 9028
rect 1537 8974 1539 9026
rect 1539 8974 1591 9026
rect 1591 8974 1593 9026
rect 1537 8972 1593 8974
rect 377 8126 433 8128
rect 377 8074 379 8126
rect 379 8074 431 8126
rect 431 8074 433 8126
rect 377 8072 433 8074
rect 903 7226 959 7228
rect 903 7174 905 7226
rect 905 7174 957 7226
rect 957 7174 959 7226
rect 903 7172 959 7174
rect 1114 7226 1170 7228
rect 1114 7174 1116 7226
rect 1116 7174 1168 7226
rect 1168 7174 1170 7226
rect 1114 7172 1170 7174
rect 1326 7226 1382 7228
rect 1326 7174 1328 7226
rect 1328 7174 1380 7226
rect 1380 7174 1382 7226
rect 1326 7172 1382 7174
rect 1537 7226 1593 7228
rect 1537 7174 1539 7226
rect 1539 7174 1591 7226
rect 1591 7174 1593 7226
rect 1537 7172 1593 7174
rect 377 6326 433 6328
rect 377 6274 379 6326
rect 379 6274 431 6326
rect 431 6274 433 6326
rect 377 6272 433 6274
rect 903 5426 959 5428
rect 903 5374 905 5426
rect 905 5374 957 5426
rect 957 5374 959 5426
rect 903 5372 959 5374
rect 1114 5426 1170 5428
rect 1114 5374 1116 5426
rect 1116 5374 1168 5426
rect 1168 5374 1170 5426
rect 1114 5372 1170 5374
rect 1326 5426 1382 5428
rect 1326 5374 1328 5426
rect 1328 5374 1380 5426
rect 1380 5374 1382 5426
rect 1326 5372 1382 5374
rect 1537 5426 1593 5428
rect 1537 5374 1539 5426
rect 1539 5374 1591 5426
rect 1591 5374 1593 5426
rect 1537 5372 1593 5374
rect 377 4526 433 4528
rect 377 4474 379 4526
rect 379 4474 431 4526
rect 431 4474 433 4526
rect 377 4472 433 4474
rect 903 3626 959 3628
rect 903 3574 905 3626
rect 905 3574 957 3626
rect 957 3574 959 3626
rect 903 3572 959 3574
rect 1114 3626 1170 3628
rect 1114 3574 1116 3626
rect 1116 3574 1168 3626
rect 1168 3574 1170 3626
rect 1114 3572 1170 3574
rect 1326 3626 1382 3628
rect 1326 3574 1328 3626
rect 1328 3574 1380 3626
rect 1380 3574 1382 3626
rect 1326 3572 1382 3574
rect 1537 3626 1593 3628
rect 1537 3574 1539 3626
rect 1539 3574 1591 3626
rect 1591 3574 1593 3626
rect 1537 3572 1593 3574
rect 377 2726 433 2728
rect 377 2674 379 2726
rect 379 2674 431 2726
rect 431 2674 433 2726
rect 377 2672 433 2674
rect 903 1826 959 1828
rect 903 1774 905 1826
rect 905 1774 957 1826
rect 957 1774 959 1826
rect 903 1772 959 1774
rect 1114 1826 1170 1828
rect 1114 1774 1116 1826
rect 1116 1774 1168 1826
rect 1168 1774 1170 1826
rect 1114 1772 1170 1774
rect 1326 1826 1382 1828
rect 1326 1774 1328 1826
rect 1328 1774 1380 1826
rect 1380 1774 1382 1826
rect 1326 1772 1382 1774
rect 1537 1826 1593 1828
rect 1537 1774 1539 1826
rect 1539 1774 1591 1826
rect 1591 1774 1593 1826
rect 1537 1772 1593 1774
rect 377 926 433 928
rect 377 874 379 926
rect 379 874 431 926
rect 431 874 433 926
rect 377 872 433 874
rect 27336 13526 27392 13528
rect 27336 13474 27338 13526
rect 27338 13474 27390 13526
rect 27390 13474 27392 13526
rect 27336 13472 27392 13474
rect 26176 12626 26232 12628
rect 26176 12574 26178 12626
rect 26178 12574 26230 12626
rect 26230 12574 26232 12626
rect 26176 12572 26232 12574
rect 26387 12626 26443 12628
rect 26387 12574 26389 12626
rect 26389 12574 26441 12626
rect 26441 12574 26443 12626
rect 26387 12572 26443 12574
rect 26599 12626 26655 12628
rect 26599 12574 26601 12626
rect 26601 12574 26653 12626
rect 26653 12574 26655 12626
rect 26599 12572 26655 12574
rect 26810 12626 26866 12628
rect 26810 12574 26812 12626
rect 26812 12574 26864 12626
rect 26864 12574 26866 12626
rect 26810 12572 26866 12574
rect 27336 11726 27392 11728
rect 27336 11674 27338 11726
rect 27338 11674 27390 11726
rect 27390 11674 27392 11726
rect 27336 11672 27392 11674
rect 26176 10826 26232 10828
rect 26176 10774 26178 10826
rect 26178 10774 26230 10826
rect 26230 10774 26232 10826
rect 26176 10772 26232 10774
rect 26387 10826 26443 10828
rect 26387 10774 26389 10826
rect 26389 10774 26441 10826
rect 26441 10774 26443 10826
rect 26387 10772 26443 10774
rect 26599 10826 26655 10828
rect 26599 10774 26601 10826
rect 26601 10774 26653 10826
rect 26653 10774 26655 10826
rect 26599 10772 26655 10774
rect 26810 10826 26866 10828
rect 26810 10774 26812 10826
rect 26812 10774 26864 10826
rect 26864 10774 26866 10826
rect 26810 10772 26866 10774
rect 27336 9926 27392 9928
rect 27336 9874 27338 9926
rect 27338 9874 27390 9926
rect 27390 9874 27392 9926
rect 27336 9872 27392 9874
rect 26176 9026 26232 9028
rect 26176 8974 26178 9026
rect 26178 8974 26230 9026
rect 26230 8974 26232 9026
rect 26176 8972 26232 8974
rect 26387 9026 26443 9028
rect 26387 8974 26389 9026
rect 26389 8974 26441 9026
rect 26441 8974 26443 9026
rect 26387 8972 26443 8974
rect 26599 9026 26655 9028
rect 26599 8974 26601 9026
rect 26601 8974 26653 9026
rect 26653 8974 26655 9026
rect 26599 8972 26655 8974
rect 26810 9026 26866 9028
rect 26810 8974 26812 9026
rect 26812 8974 26864 9026
rect 26864 8974 26866 9026
rect 26810 8972 26866 8974
rect 27336 8126 27392 8128
rect 27336 8074 27338 8126
rect 27338 8074 27390 8126
rect 27390 8074 27392 8126
rect 27336 8072 27392 8074
rect 26176 7226 26232 7228
rect 26176 7174 26178 7226
rect 26178 7174 26230 7226
rect 26230 7174 26232 7226
rect 26176 7172 26232 7174
rect 26387 7226 26443 7228
rect 26387 7174 26389 7226
rect 26389 7174 26441 7226
rect 26441 7174 26443 7226
rect 26387 7172 26443 7174
rect 26599 7226 26655 7228
rect 26599 7174 26601 7226
rect 26601 7174 26653 7226
rect 26653 7174 26655 7226
rect 26599 7172 26655 7174
rect 26810 7226 26866 7228
rect 26810 7174 26812 7226
rect 26812 7174 26864 7226
rect 26864 7174 26866 7226
rect 26810 7172 26866 7174
rect 27336 6326 27392 6328
rect 27336 6274 27338 6326
rect 27338 6274 27390 6326
rect 27390 6274 27392 6326
rect 27336 6272 27392 6274
rect 26176 5426 26232 5428
rect 26176 5374 26178 5426
rect 26178 5374 26230 5426
rect 26230 5374 26232 5426
rect 26176 5372 26232 5374
rect 26387 5426 26443 5428
rect 26387 5374 26389 5426
rect 26389 5374 26441 5426
rect 26441 5374 26443 5426
rect 26387 5372 26443 5374
rect 26599 5426 26655 5428
rect 26599 5374 26601 5426
rect 26601 5374 26653 5426
rect 26653 5374 26655 5426
rect 26599 5372 26655 5374
rect 26810 5426 26866 5428
rect 26810 5374 26812 5426
rect 26812 5374 26864 5426
rect 26864 5374 26866 5426
rect 26810 5372 26866 5374
rect 27336 4526 27392 4528
rect 27336 4474 27338 4526
rect 27338 4474 27390 4526
rect 27390 4474 27392 4526
rect 27336 4472 27392 4474
rect 26176 3626 26232 3628
rect 26176 3574 26178 3626
rect 26178 3574 26230 3626
rect 26230 3574 26232 3626
rect 26176 3572 26232 3574
rect 26387 3626 26443 3628
rect 26387 3574 26389 3626
rect 26389 3574 26441 3626
rect 26441 3574 26443 3626
rect 26387 3572 26443 3574
rect 26599 3626 26655 3628
rect 26599 3574 26601 3626
rect 26601 3574 26653 3626
rect 26653 3574 26655 3626
rect 26599 3572 26655 3574
rect 26810 3626 26866 3628
rect 26810 3574 26812 3626
rect 26812 3574 26864 3626
rect 26864 3574 26866 3626
rect 26810 3572 26866 3574
rect 27336 2726 27392 2728
rect 27336 2674 27338 2726
rect 27338 2674 27390 2726
rect 27390 2674 27392 2726
rect 27336 2672 27392 2674
rect 26176 1826 26232 1828
rect 26176 1774 26178 1826
rect 26178 1774 26230 1826
rect 26230 1774 26232 1826
rect 26176 1772 26232 1774
rect 26387 1826 26443 1828
rect 26387 1774 26389 1826
rect 26389 1774 26441 1826
rect 26441 1774 26443 1826
rect 26387 1772 26443 1774
rect 26599 1826 26655 1828
rect 26599 1774 26601 1826
rect 26601 1774 26653 1826
rect 26653 1774 26655 1826
rect 26599 1772 26655 1774
rect 26810 1826 26866 1828
rect 26810 1774 26812 1826
rect 26812 1774 26864 1826
rect 26864 1774 26866 1826
rect 26810 1772 26866 1774
rect 903 26 959 28
rect 903 -26 905 26
rect 905 -26 957 26
rect 957 -26 959 26
rect 903 -28 959 -26
rect 1114 26 1170 28
rect 1114 -26 1116 26
rect 1116 -26 1168 26
rect 1168 -26 1170 26
rect 1114 -28 1170 -26
rect 1326 26 1382 28
rect 1326 -26 1328 26
rect 1328 -26 1380 26
rect 1380 -26 1382 26
rect 1326 -28 1382 -26
rect 1537 26 1593 28
rect 1537 -26 1539 26
rect 1539 -26 1591 26
rect 1591 -26 1593 26
rect 1537 -28 1593 -26
rect 27336 926 27392 928
rect 27336 874 27338 926
rect 27338 874 27390 926
rect 27390 874 27392 926
rect 27336 872 27392 874
rect 26176 26 26232 28
rect 26176 -26 26178 26
rect 26178 -26 26230 26
rect 26230 -26 26232 26
rect 26176 -28 26232 -26
rect 26387 26 26443 28
rect 26387 -26 26389 26
rect 26389 -26 26441 26
rect 26441 -26 26443 26
rect 26387 -28 26443 -26
rect 26599 26 26655 28
rect 26599 -26 26601 26
rect 26601 -26 26653 26
rect 26653 -26 26655 26
rect 26599 -28 26655 -26
rect 26810 26 26866 28
rect 26810 -26 26812 26
rect 26812 -26 26864 26
rect 26864 -26 26866 26
rect 26810 -28 26866 -26
<< metal3 >>
rect -1048 15328 28817 15401
rect -1048 15272 166 15328
rect 222 15272 377 15328
rect 433 15272 5611 15328
rect 5667 15272 5822 15328
rect 5878 15272 6033 15328
rect 6089 15272 6244 15328
rect 6300 15272 11573 15328
rect 11629 15272 11753 15328
rect 11809 15272 21458 15328
rect 21514 15272 21669 15328
rect 21725 15272 21880 15328
rect 21936 15272 22091 15328
rect 22147 15272 27336 15328
rect 27392 15272 27547 15328
rect 27603 15272 28817 15328
rect -1048 15200 28817 15272
rect 1725 15199 25945 15200
rect 0 14907 5307 14941
rect -1 14847 5307 14907
rect -1 14791 4371 14847
rect 4427 14791 4582 14847
rect 4638 14791 4793 14847
rect 4849 14791 5004 14847
rect 5060 14791 5215 14847
rect 5271 14791 5307 14847
rect -1 14773 5307 14791
rect 0 14739 5307 14773
rect 8186 14845 13478 14884
rect 8186 14789 8222 14845
rect 8278 14789 8433 14845
rect 8489 14789 8644 14845
rect 8700 14789 8855 14845
rect 8911 14789 12331 14845
rect 12387 14789 12542 14845
rect 12598 14789 12753 14845
rect 12809 14789 12964 14845
rect 13020 14789 13175 14845
rect 13231 14789 13385 14845
rect 13441 14789 13478 14845
rect 13994 14838 14545 14877
rect 13994 14803 14031 14838
rect 8186 14750 13478 14789
rect 13993 14782 14031 14803
rect 14087 14782 14242 14838
rect 14298 14782 14453 14838
rect 14509 14782 14545 14838
rect 13993 14744 14545 14782
rect 22365 14845 27769 14941
rect 22365 14789 22402 14845
rect 22458 14789 22613 14845
rect 22669 14789 22824 14845
rect 22880 14789 23035 14845
rect 23091 14789 23246 14845
rect 23302 14789 27769 14845
rect -1 14500 2204 14501
rect -3364 14428 2204 14500
rect -3364 14372 903 14428
rect 959 14372 1114 14428
rect 1170 14372 1326 14428
rect 1382 14372 1537 14428
rect 1593 14372 2204 14428
rect -3364 14300 2204 14372
rect 12063 14428 12615 14467
rect 13993 14432 14092 14744
rect 22365 14739 27769 14789
rect 25565 14500 27770 14501
rect 12063 14372 12100 14428
rect 12156 14372 12311 14428
rect 12367 14372 12522 14428
rect 12578 14372 12615 14428
rect 12063 14333 12615 14372
rect 25565 14428 31133 14500
rect 25565 14372 26176 14428
rect 26232 14372 26387 14428
rect 26443 14372 26599 14428
rect 26655 14372 26810 14428
rect 26866 14372 31133 14428
rect 25565 14300 31133 14372
rect -3364 13859 2204 14061
rect 25565 13859 31133 14061
rect -3364 13528 2204 13599
rect -3364 13472 377 13528
rect 433 13472 2204 13528
rect -3364 13399 2204 13472
rect 25565 13528 31133 13599
rect 25565 13472 27336 13528
rect 27392 13472 31133 13528
rect 25565 13399 31133 13472
rect -3364 12939 2204 13141
rect 25565 12939 31133 13141
rect -3364 12628 2204 12700
rect -3364 12572 903 12628
rect 959 12572 1114 12628
rect 1170 12572 1326 12628
rect 1382 12572 1537 12628
rect 1593 12572 2204 12628
rect -3364 12500 2204 12572
rect 25565 12628 31133 12700
rect 25565 12572 26176 12628
rect 26232 12572 26387 12628
rect 26443 12572 26599 12628
rect 26655 12572 26810 12628
rect 26866 12572 31133 12628
rect 25565 12500 31133 12572
rect -3364 12059 2204 12261
rect 25565 12059 31133 12261
rect -3364 11728 2204 11799
rect -3364 11672 377 11728
rect 433 11672 2204 11728
rect -3364 11599 2204 11672
rect 25565 11728 31133 11799
rect 25565 11672 27336 11728
rect 27392 11672 31133 11728
rect 25565 11599 31133 11672
rect -3364 11139 2204 11341
rect 25565 11139 31133 11341
rect -3364 10828 2204 10900
rect -3364 10772 903 10828
rect 959 10772 1114 10828
rect 1170 10772 1326 10828
rect 1382 10772 1537 10828
rect 1593 10772 2204 10828
rect -3364 10700 2204 10772
rect 25565 10828 31133 10900
rect 25565 10772 26176 10828
rect 26232 10772 26387 10828
rect 26443 10772 26599 10828
rect 26655 10772 26810 10828
rect 26866 10772 31133 10828
rect 25565 10700 31133 10772
rect -3364 10259 2204 10461
rect 25565 10259 31133 10461
rect -3364 9928 2204 9999
rect -3364 9872 377 9928
rect 433 9872 2204 9928
rect -3364 9799 2204 9872
rect 25565 9928 31133 9999
rect 25565 9872 27336 9928
rect 27392 9872 31133 9928
rect 25565 9799 31133 9872
rect -3364 9339 2204 9541
rect 25565 9339 31133 9541
rect -3364 9028 2204 9100
rect -3364 8972 903 9028
rect 959 8972 1114 9028
rect 1170 8972 1326 9028
rect 1382 8972 1537 9028
rect 1593 8972 2204 9028
rect -3364 8900 2204 8972
rect 25565 9028 31133 9100
rect 25565 8972 26176 9028
rect 26232 8972 26387 9028
rect 26443 8972 26599 9028
rect 26655 8972 26810 9028
rect 26866 8972 31133 9028
rect 25565 8900 31133 8972
rect -3364 8459 2204 8661
rect 25565 8459 31133 8661
rect -3364 8128 2204 8199
rect -3364 8072 377 8128
rect 433 8072 2204 8128
rect -3364 7999 2204 8072
rect 25565 8128 31133 8199
rect 25565 8072 27336 8128
rect 27392 8072 31133 8128
rect 25565 7999 31133 8072
rect -3364 7539 2204 7741
rect 25565 7539 31133 7741
rect -3364 7228 2204 7300
rect -3364 7172 903 7228
rect 959 7172 1114 7228
rect 1170 7172 1326 7228
rect 1382 7172 1537 7228
rect 1593 7172 2204 7228
rect -3364 7100 2204 7172
rect 25565 7228 31133 7300
rect 25565 7172 26176 7228
rect 26232 7172 26387 7228
rect 26443 7172 26599 7228
rect 26655 7172 26810 7228
rect 26866 7172 31133 7228
rect 25565 7100 31133 7172
rect -3364 6659 2204 6861
rect 25565 6659 31133 6861
rect -3364 6328 2204 6399
rect -3364 6272 377 6328
rect 433 6272 2204 6328
rect -3364 6199 2204 6272
rect 25565 6328 31133 6399
rect 25565 6272 27336 6328
rect 27392 6272 31133 6328
rect 25565 6199 31133 6272
rect -3364 5739 2204 5941
rect 25565 5739 31133 5941
rect -3364 5428 2204 5500
rect -3364 5372 903 5428
rect 959 5372 1114 5428
rect 1170 5372 1326 5428
rect 1382 5372 1537 5428
rect 1593 5372 2204 5428
rect -3364 5300 2204 5372
rect 25565 5428 31133 5500
rect 25565 5372 26176 5428
rect 26232 5372 26387 5428
rect 26443 5372 26599 5428
rect 26655 5372 26810 5428
rect 26866 5372 31133 5428
rect 25565 5300 31133 5372
rect -3364 4859 2204 5061
rect 25565 4859 31133 5061
rect -3364 4528 2204 4599
rect -3364 4472 377 4528
rect 433 4472 2204 4528
rect -3364 4399 2204 4472
rect 25565 4528 31133 4599
rect 25565 4472 27336 4528
rect 27392 4472 31133 4528
rect 25565 4399 31133 4472
rect -3364 3939 2204 4141
rect 25565 3939 31133 4141
rect -3364 3628 2204 3700
rect -3364 3572 903 3628
rect 959 3572 1114 3628
rect 1170 3572 1326 3628
rect 1382 3572 1537 3628
rect 1593 3572 2204 3628
rect -3364 3500 2204 3572
rect 25565 3628 31133 3700
rect 25565 3572 26176 3628
rect 26232 3572 26387 3628
rect 26443 3572 26599 3628
rect 26655 3572 26810 3628
rect 26866 3572 31133 3628
rect 25565 3500 31133 3572
rect -3364 3059 2204 3261
rect 25565 3059 31133 3261
rect -3364 2728 2204 2799
rect -3364 2672 377 2728
rect 433 2672 2204 2728
rect -3364 2599 2204 2672
rect 25565 2728 31133 2799
rect 25565 2672 27336 2728
rect 27392 2672 31133 2728
rect 25565 2599 31133 2672
rect -3364 2139 2204 2341
rect 25565 2139 31133 2341
rect -3364 1828 2204 1900
rect -3364 1772 903 1828
rect 959 1772 1114 1828
rect 1170 1772 1326 1828
rect 1382 1772 1537 1828
rect 1593 1772 2204 1828
rect -3364 1700 2204 1772
rect 25565 1828 31133 1900
rect 25565 1772 26176 1828
rect 26232 1772 26387 1828
rect 26443 1772 26599 1828
rect 26655 1772 26810 1828
rect 26866 1772 31133 1828
rect 25565 1700 31133 1772
rect -3364 1259 2204 1461
rect 25565 1259 31133 1461
rect -3364 928 2204 999
rect -3364 872 377 928
rect 433 872 2204 928
rect -3364 799 2204 872
rect 25565 928 31133 999
rect 25565 872 27336 928
rect 27392 872 31133 928
rect 25565 799 31133 872
rect -3364 339 2204 541
rect 25565 339 31133 541
rect -3364 28 2204 100
rect -3364 -28 903 28
rect 959 -28 1114 28
rect 1170 -28 1326 28
rect 1382 -28 1537 28
rect 1593 -28 2204 28
rect -3364 -100 2204 -28
rect 25565 28 31133 100
rect 25565 -28 26176 28
rect 26232 -28 26387 28
rect 26443 -28 26599 28
rect 26655 -28 26810 28
rect 26866 -28 31133 28
rect 25565 -100 31133 -28
use M1_NACTIVE$$203393068_128x8m81  M1_NACTIVE$$203393068_128x8m81_0
timestamp 1698431365
transform 1 0 14063 0 1 15359
box 0 0 1 1
use M1_NWELL$$204218412_128x8m81  M1_NWELL$$204218412_128x8m81_0
timestamp 1698431365
transform -1 0 25568 0 1 15286
box 0 0 1 1
use M1_NWELL$$204218412_128x8m81  M1_NWELL$$204218412_128x8m81_1
timestamp 1698431365
transform 1 0 2200 0 1 15286
box 0 0 1 1
use M1_PACTIVE$$204148780_128x8m81  M1_PACTIVE$$204148780_128x8m81_0
timestamp 1698431365
transform 1 0 11463 0 1 15359
box 0 0 1 1
use M1_PACTIVE$$204148780_128x8m81  M1_PACTIVE$$204148780_128x8m81_1
timestamp 1698431365
transform 1 0 21475 0 1 15359
box 0 0 1 1
use M1_PACTIVE$$204148780_128x8m81  M1_PACTIVE$$204148780_128x8m81_2
timestamp 1698431365
transform 1 0 4390 0 1 15359
box 0 0 1 1
use M1_PACTIVE$$204149804_128x8m81  M1_PACTIVE$$204149804_128x8m81_0
timestamp 1698431365
transform 1 0 15860 0 1 15359
box 0 0 1 1
use M1_POLY2$$204150828_128x8m81  M1_POLY2$$204150828_128x8m81_0
timestamp 1698431365
transform 1 0 9381 0 1 15048
box 0 0 1 1
use M1_POLY24310590548732_128x8m81  M1_POLY24310590548732_128x8m81_0
timestamp 1698431365
transform 1 0 15413 0 1 15341
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_0
timestamp 1698431365
transform 0 -1 13712 1 0 15293
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_1
timestamp 1698431365
transform 1 0 15625 0 1 15001
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_2
timestamp 1698431365
transform 1 0 18313 0 1 15036
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_3
timestamp 1698431365
transform 1 0 12040 0 1 14961
box 0 0 1 1
use M2_M1$$201262124_128x8m81  M2_M1$$201262124_128x8m81_0
timestamp 1698431365
transform 1 0 13701 0 1 15291
box 0 0 1 1
use M2_M1$$204138540_128x8m81  M2_M1$$204138540_128x8m81_0
timestamp 1698431365
transform 1 0 10402 0 1 15048
box 0 0 1 1
use M2_M1$$204138540_128x8m81  M2_M1$$204138540_128x8m81_1
timestamp 1698431365
transform 1 0 14059 0 1 15352
box 0 0 1 1
use M2_M1$$204139564_128x8m81  M2_M1$$204139564_128x8m81_0
timestamp 1698431365
transform 1 0 11601 0 1 15305
box 0 0 1 1
use M2_M1$$204140588_128x8m81  M2_M1$$204140588_128x8m81_0
timestamp 1698431365
transform 1 0 12359 0 1 14817
box 0 0 1 1
use M2_M1$$204141612_128x8m81  M2_M1$$204141612_128x8m81_0
timestamp 1698431365
transform 1 0 15126 0 1 15352
box 0 0 1 1
use M2_M1$$204141612_128x8m81  M2_M1$$204141612_128x8m81_1
timestamp 1698431365
transform 1 0 20177 0 1 15280
box 0 0 1 1
use M2_M1$$204141612_128x8m81  M2_M1$$204141612_128x8m81_2
timestamp 1698431365
transform 1 0 20177 0 1 14817
box 0 0 1 1
use M2_M1$$204220460_128x8m81  M2_M1$$204220460_128x8m81_0
timestamp 1698431365
transform 1 0 6792 0 1 14817
box 0 0 1 1
use M2_M1$$204220460_128x8m81  M2_M1$$204220460_128x8m81_1
timestamp 1698431365
transform 1 0 22430 0 1 14817
box 0 0 1 1
use M2_M1$$204220460_128x8m81  M2_M1$$204220460_128x8m81_2
timestamp 1698431365
transform 1 0 4399 0 1 14819
box 0 0 1 1
use M2_M1$$204220460_128x8m81  M2_M1$$204220460_128x8m81_3
timestamp 1698431365
transform 1 0 6792 0 1 15280
box 0 0 1 1
use M2_M1$$204221484_128x8m81  M2_M1$$204221484_128x8m81_0
timestamp 1698431365
transform -1 0 25612 0 1 15300
box 0 0 1 1
use M2_M1$$204221484_128x8m81  M2_M1$$204221484_128x8m81_1
timestamp 1698431365
transform 1 0 2156 0 1 15300
box 0 0 1 1
use M2_M1$$204222508_128x8m81  M2_M1$$204222508_128x8m81_0
timestamp 1698431365
transform 1 0 21486 0 1 15300
box 0 0 1 1
use M2_M1$$204222508_128x8m81  M2_M1$$204222508_128x8m81_1
timestamp 1698431365
transform 1 0 5639 0 1 15300
box 0 0 1 1
use M3_M2$$204142636_128x8m81  M3_M2$$204142636_128x8m81_0
timestamp 1698431365
transform 1 0 5639 0 1 15300
box 0 0 1 1
use M3_M2$$204142636_128x8m81  M3_M2$$204142636_128x8m81_1
timestamp 1698431365
transform 1 0 8250 0 1 14817
box 0 0 1 1
use M3_M2$$204142636_128x8m81  M3_M2$$204142636_128x8m81_2
timestamp 1698431365
transform 1 0 21486 0 1 15300
box 0 0 1 1
use M3_M2$$204143660_128x8m81  M3_M2$$204143660_128x8m81_0
timestamp 1698431365
transform 1 0 11601 0 1 15300
box 0 0 1 1
use M3_M2$$204144684_128x8m81  M3_M2$$204144684_128x8m81_0
timestamp 1698431365
transform 1 0 22430 0 1 14817
box 0 0 1 1
use M3_M2$$204144684_128x8m81  M3_M2$$204144684_128x8m81_1
timestamp 1698431365
transform 1 0 4399 0 1 14819
box 0 0 1 1
use M3_M2$$204145708_128x8m81  M3_M2$$204145708_128x8m81_0
timestamp 1698431365
transform 1 0 12359 0 1 14817
box 0 0 1 1
use M3_M2$$204146732_128x8m81  M3_M2$$204146732_128x8m81_0
timestamp 1698431365
transform 1 0 14059 0 1 14810
box 0 0 1 1
use M3_M2$$204147756_128x8m81  M3_M2$$204147756_128x8m81_0
timestamp 1698431365
transform 1 0 12339 0 1 14400
box 0 0 1 1
use nmos_1p2$$204213292_R90_128x8m81  nmos_1p2$$204213292_R90_128x8m81_0
timestamp 1698431365
transform 0 -1 6346 1 0 14903
box -31 0 -30 1
use nmos_1p2$$204215340_128x8m81  nmos_1p2$$204215340_128x8m81_0
timestamp 1698431365
transform 0 -1 13604 -1 0 14962
box -31 0 -30 1
use nmos_5p04310590548799_128x8m81  nmos_5p04310590548799_128x8m81_0
timestamp 1698431365
transform 0 -1 23346 1 0 14872
box 0 0 1 1
use nmos_5p043105905487111_128x8m81  nmos_5p043105905487111_128x8m81_0
timestamp 1698431365
transform 0 -1 16283 1 0 14872
box 0 0 1 1
use nmos_5p043105905487111_128x8m81  nmos_5p043105905487111_128x8m81_1
timestamp 1698431365
transform 0 -1 11913 1 0 14872
box 0 0 1 1
use pmos_1p2$$204216364_128x8m81  pmos_1p2$$204216364_128x8m81_0
timestamp 1698431365
transform 0 -1 20950 1 0 14903
box -31 0 -30 1
use pmos_1p2$$204216364_128x8m81  pmos_1p2$$204216364_128x8m81_1
timestamp 1698431365
transform 0 -1 9245 1 0 14903
box -31 0 -30 1
use pmos_1p2$$204217388_R90_128x8m81  pmos_1p2$$204217388_R90_128x8m81_0
timestamp 1698431365
transform 0 -1 11004 1 0 14903
box -31 0 -30 1
use pmos_5p043105905487100_128x8m81  pmos_5p043105905487100_128x8m81_0
timestamp 1698431365
transform 0 -1 15304 1 0 14872
box 0 0 1 1
use pmos_5p043105905487100_128x8m81  pmos_5p043105905487100_128x8m81_1
timestamp 1698431365
transform 0 -1 17974 1 0 14872
box 0 0 1 1
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_0
timestamp 1698431365
transform 0 -1 2203 -1 0 14550
box 0 0 1 1
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_1
timestamp 1698431365
transform 0 -1 2203 -1 0 12750
box 0 0 1 1
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_2
timestamp 1698431365
transform 0 -1 2203 -1 0 10950
box 0 0 1 1
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_3
timestamp 1698431365
transform 0 -1 2203 -1 0 9150
box 0 0 1 1
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_4
timestamp 1698431365
transform 0 -1 2203 -1 0 7350
box 0 0 1 1
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_5
timestamp 1698431365
transform 0 -1 2203 -1 0 5550
box 0 0 1 1
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_6
timestamp 1698431365
transform 0 -1 2203 -1 0 3750
box 0 0 1 1
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_7
timestamp 1698431365
transform 0 -1 2203 -1 0 1950
box 0 0 1 1
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_8
timestamp 1698431365
transform 0 1 25566 -1 0 14550
box 0 0 1 1
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_9
timestamp 1698431365
transform 0 1 25566 -1 0 12750
box 0 0 1 1
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_10
timestamp 1698431365
transform 0 1 25566 -1 0 10950
box 0 0 1 1
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_11
timestamp 1698431365
transform 0 1 25566 -1 0 9150
box 0 0 1 1
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_12
timestamp 1698431365
transform 0 1 25566 -1 0 7350
box 0 0 1 1
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_13
timestamp 1698431365
transform 0 1 25566 -1 0 5550
box 0 0 1 1
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_14
timestamp 1698431365
transform 0 1 25566 -1 0 3750
box 0 0 1 1
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_15
timestamp 1698431365
transform 0 1 25566 -1 0 1950
box 0 0 1 1
use pmoscap_W2_5_R270_128x8m81  pmoscap_W2_5_R270_128x8m81_0
timestamp 1698431365
transform 0 -1 2203 -1 0 15450
box 150 220 1051 2048
use pmoscap_W2_5_R270_128x8m81  pmoscap_W2_5_R270_128x8m81_1
timestamp 1698431365
transform 0 1 25566 -1 0 15450
box 150 220 1051 2048
use xdec16_128x8_128x8m81  xdec16_128x8_128x8m81_0
timestamp 1698431365
transform 1 0 1726 0 1 0
box 0 -228 24219 14628
<< labels >>
rlabel metal3 s 27705 14840 27705 14840 4 DRWL
port 1 nsew
rlabel metal3 s 27705 5860 27705 5860 4 RWL[6]
port 2 nsew
rlabel metal3 s 27705 4060 27705 4060 4 RWL[4]
port 3 nsew
rlabel metal3 s 27705 2260 27705 2260 4 RWL[2]
port 4 nsew
rlabel metal3 s 27705 460 27705 460 4 RWL[0]
port 5 nsew
rlabel metal3 s 27705 1340 27705 1340 4 RWL[1]
port 6 nsew
rlabel metal3 s 27705 3140 27705 3140 4 RWL[3]
port 7 nsew
rlabel metal3 s 27705 4940 27705 4940 4 RWL[5]
port 8 nsew
rlabel metal3 s 27705 6740 27705 6740 4 RWL[7]
port 9 nsew
rlabel metal3 s 27705 7660 27705 7660 4 RWL[8]
port 10 nsew
rlabel metal3 s 27705 8540 27705 8540 4 RWL[9]
port 11 nsew
rlabel metal3 s 27705 9460 27705 9460 4 RWL[10]
port 12 nsew
rlabel metal3 s 27705 10340 27705 10340 4 RWL[11]
port 13 nsew
rlabel metal3 s 27705 11260 27705 11260 4 RWL[12]
port 14 nsew
rlabel metal3 s 27705 12140 27705 12140 4 RWL[13]
port 15 nsew
rlabel metal3 s 27705 13060 27705 13060 4 RWL[14]
port 16 nsew
rlabel metal3 s 27705 13940 27705 13940 4 RWL[15]
port 17 nsew
rlabel metal3 s 64 9460 64 9460 4 LWL[10]
port 18 nsew
rlabel metal3 s 64 10340 64 10340 4 LWL[11]
port 19 nsew
rlabel metal3 s 64 11260 64 11260 4 LWL[12]
port 20 nsew
rlabel metal3 s 64 12140 64 12140 4 LWL[13]
port 21 nsew
rlabel metal3 s 64 13060 64 13060 4 LWL[14]
port 22 nsew
rlabel metal3 s 64 13940 64 13940 4 LWL[15]
port 23 nsew
rlabel metal3 s 64 4940 64 4940 4 LWL[5]
port 24 nsew
rlabel metal3 s 64 4060 64 4060 4 LWL[4]
port 25 nsew
rlabel metal3 s 64 3140 64 3140 4 LWL[3]
port 26 nsew
rlabel metal3 s 64 2260 64 2260 4 LWL[2]
port 27 nsew
rlabel metal3 s 64 1340 64 1340 4 LWL[1]
port 28 nsew
rlabel metal3 s 64 460 64 460 4 LWL[0]
port 29 nsew
rlabel metal3 s 64 7660 64 7660 4 LWL[8]
port 30 nsew
rlabel metal3 s 64 8540 64 8540 4 LWL[9]
port 31 nsew
rlabel metal3 s 64 5860 64 5860 4 LWL[6]
port 32 nsew
rlabel metal3 s 64 6740 64 6740 4 LWL[7]
port 33 nsew
rlabel metal3 s 134 15300 134 15300 4 vss
port 34 nsew
rlabel metal3 s 134 14400 134 14400 4 vdd
port 35 nsew
rlabel metal3 s 64 14840 64 14840 4 DLWL
port 36 nsew
rlabel metal2 s 14794 -97 14794 -97 4 xb[0]
port 37 nsew
rlabel metal2 s 14417 -97 14417 -97 4 xb[1]
port 38 nsew
rlabel metal2 s 14039 -97 14039 -97 4 xb[2]
port 39 nsew
rlabel metal2 s 13661 -97 13661 -97 4 xb[3]
port 40 nsew
rlabel metal2 s 16947 -97 16947 -97 4 xa[7]
port 41 nsew
rlabel metal2 s 17324 -97 17324 -97 4 xa[6]
port 42 nsew
rlabel metal2 s 17702 -97 17702 -97 4 xa[5]
port 43 nsew
rlabel metal2 s 18080 -97 18080 -97 4 xa[4]
port 44 nsew
rlabel metal2 s 19591 -97 19591 -97 4 xa[0]
port 45 nsew
rlabel metal2 s 8626 45 8626 45 4 men
port 46 nsew
rlabel metal2 s 18457 -97 18457 -97 4 xa[3]
port 47 nsew
rlabel metal2 s 18835 -97 18835 -97 4 xa[2]
port 48 nsew
rlabel metal2 s 19213 -97 19213 -97 4 xa[1]
port 49 nsew
rlabel metal2 s 13284 -97 13284 -97 4 xc[0]
port 50 nsew
rlabel metal2 s 12906 -97 12906 -97 4 xc[1]
port 51 nsew
<< properties >>
string GDS_END 2206704
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 2192594
<< end >>
