magic
tech gf180mcuA
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 453 4118 1094
<< pwell >>
rect -86 -86 4118 453
<< mvnmos >>
rect 124 156 244 296
rect 348 156 468 296
rect 575 156 695 296
rect 799 156 919 296
rect 967 156 1087 296
rect 1191 156 1311 296
rect 1567 156 1687 296
rect 1791 156 1911 296
rect 2247 156 2367 316
rect 2471 156 2591 316
rect 2695 156 2815 316
rect 3067 133 3187 333
rect 3291 133 3411 333
rect 3515 133 3635 333
rect 3739 133 3859 333
<< mvpmos >>
rect 340 576 440 852
rect 488 576 588 852
rect 683 576 783 852
rect 887 576 987 852
rect 1035 576 1135 852
rect 1239 576 1339 852
rect 1587 573 1687 849
rect 1791 573 1891 849
rect 2287 585 2387 921
rect 2491 585 2591 921
rect 2639 585 2739 921
rect 3077 573 3177 939
rect 3281 573 3381 939
rect 3485 573 3585 939
rect 3689 573 3789 939
<< mvndiff >>
rect 36 215 124 296
rect 36 169 49 215
rect 95 169 124 215
rect 36 156 124 169
rect 244 215 348 296
rect 244 169 273 215
rect 319 169 348 215
rect 244 156 348 169
rect 468 215 575 296
rect 468 169 497 215
rect 543 169 575 215
rect 468 156 575 169
rect 695 215 799 296
rect 695 169 724 215
rect 770 169 799 215
rect 695 156 799 169
rect 919 156 967 296
rect 1087 215 1191 296
rect 1087 169 1116 215
rect 1162 169 1191 215
rect 1087 156 1191 169
rect 1311 215 1399 296
rect 1311 169 1340 215
rect 1386 169 1399 215
rect 1311 156 1399 169
rect 1479 215 1567 296
rect 1479 169 1492 215
rect 1538 169 1567 215
rect 1479 156 1567 169
rect 1687 215 1791 296
rect 1687 169 1716 215
rect 1762 169 1791 215
rect 1687 156 1791 169
rect 1911 215 1999 296
rect 1911 169 1940 215
rect 1986 169 1999 215
rect 1911 156 1999 169
rect 2159 303 2247 316
rect 2159 257 2172 303
rect 2218 257 2247 303
rect 2159 156 2247 257
rect 2367 215 2471 316
rect 2367 169 2396 215
rect 2442 169 2471 215
rect 2367 156 2471 169
rect 2591 303 2695 316
rect 2591 257 2620 303
rect 2666 257 2695 303
rect 2591 156 2695 257
rect 2815 215 2903 316
rect 2815 169 2844 215
rect 2890 169 2903 215
rect 2815 156 2903 169
rect 2979 309 3067 333
rect 2979 169 2992 309
rect 3038 169 3067 309
rect 2979 133 3067 169
rect 3187 309 3291 333
rect 3187 169 3216 309
rect 3262 169 3291 309
rect 3187 133 3291 169
rect 3411 203 3515 333
rect 3411 157 3440 203
rect 3486 157 3515 203
rect 3411 133 3515 157
rect 3635 309 3739 333
rect 3635 169 3664 309
rect 3710 169 3739 309
rect 3635 133 3739 169
rect 3859 309 3947 333
rect 3859 169 3888 309
rect 3934 169 3947 309
rect 3859 133 3947 169
<< mvpdiff >>
rect 252 781 340 852
rect 252 641 265 781
rect 311 641 340 781
rect 252 576 340 641
rect 440 576 488 852
rect 588 576 683 852
rect 783 781 887 852
rect 783 641 812 781
rect 858 641 887 781
rect 783 576 887 641
rect 987 576 1035 852
rect 1135 781 1239 852
rect 1135 641 1164 781
rect 1210 641 1239 781
rect 1135 576 1239 641
rect 1339 769 1427 852
rect 1339 629 1368 769
rect 1414 629 1427 769
rect 1339 576 1427 629
rect 1499 769 1587 849
rect 1499 629 1512 769
rect 1558 629 1587 769
rect 1499 573 1587 629
rect 1687 781 1791 849
rect 1687 641 1716 781
rect 1762 641 1791 781
rect 1687 573 1791 641
rect 1891 781 1979 849
rect 1891 641 1920 781
rect 1966 641 1979 781
rect 1891 573 1979 641
rect 2199 644 2287 921
rect 2199 598 2212 644
rect 2258 598 2287 644
rect 2199 585 2287 598
rect 2387 908 2491 921
rect 2387 768 2416 908
rect 2462 768 2491 908
rect 2387 585 2491 768
rect 2591 585 2639 921
rect 2739 781 2827 921
rect 2739 641 2768 781
rect 2814 641 2827 781
rect 2739 585 2827 641
rect 2989 781 3077 939
rect 2989 641 3002 781
rect 3048 641 3077 781
rect 2989 573 3077 641
rect 3177 781 3281 939
rect 3177 641 3206 781
rect 3252 641 3281 781
rect 3177 573 3281 641
rect 3381 781 3485 939
rect 3381 641 3410 781
rect 3456 641 3485 781
rect 3381 573 3485 641
rect 3585 781 3689 939
rect 3585 641 3614 781
rect 3660 641 3689 781
rect 3585 573 3689 641
rect 3789 781 3877 939
rect 3789 641 3818 781
rect 3864 641 3877 781
rect 3789 573 3877 641
<< mvndiffc >>
rect 49 169 95 215
rect 273 169 319 215
rect 497 169 543 215
rect 724 169 770 215
rect 1116 169 1162 215
rect 1340 169 1386 215
rect 1492 169 1538 215
rect 1716 169 1762 215
rect 1940 169 1986 215
rect 2172 257 2218 303
rect 2396 169 2442 215
rect 2620 257 2666 303
rect 2844 169 2890 215
rect 2992 169 3038 309
rect 3216 169 3262 309
rect 3440 157 3486 203
rect 3664 169 3710 309
rect 3888 169 3934 309
<< mvpdiffc >>
rect 265 641 311 781
rect 812 641 858 781
rect 1164 641 1210 781
rect 1368 629 1414 769
rect 1512 629 1558 769
rect 1716 641 1762 781
rect 1920 641 1966 781
rect 2212 598 2258 644
rect 2416 768 2462 908
rect 2768 641 2814 781
rect 3002 641 3048 781
rect 3206 641 3252 781
rect 3410 641 3456 781
rect 3614 641 3660 781
rect 3818 641 3864 781
<< polysilicon >>
rect 1035 944 1891 984
rect 340 852 440 896
rect 488 852 588 896
rect 683 852 783 896
rect 887 852 987 896
rect 1035 852 1135 944
rect 1239 852 1339 896
rect 1587 849 1687 893
rect 1791 849 1891 944
rect 2287 921 2387 965
rect 2491 921 2591 965
rect 2639 921 2739 965
rect 3077 939 3177 983
rect 3281 939 3381 983
rect 3485 939 3585 983
rect 3689 939 3789 983
rect 340 532 440 576
rect 488 532 588 576
rect 683 532 783 576
rect 340 434 380 532
rect 488 434 528 532
rect 743 516 783 532
rect 743 476 839 516
rect 124 421 380 434
rect 124 375 148 421
rect 194 394 380 421
rect 428 421 528 434
rect 194 375 244 394
rect 124 296 244 375
rect 428 375 469 421
rect 515 375 528 421
rect 428 362 528 375
rect 655 415 751 428
rect 655 369 692 415
rect 738 369 751 415
rect 428 340 468 362
rect 655 356 751 369
rect 655 340 695 356
rect 348 296 468 340
rect 575 296 695 340
rect 799 340 839 476
rect 887 492 987 576
rect 887 446 905 492
rect 951 446 987 492
rect 887 433 987 446
rect 1035 532 1135 576
rect 1239 532 1339 576
rect 1035 340 1087 532
rect 1239 340 1311 532
rect 1587 421 1687 573
rect 1587 375 1604 421
rect 1650 375 1687 421
rect 1587 340 1687 375
rect 799 296 919 340
rect 967 296 1087 340
rect 1191 296 1311 340
rect 1567 296 1687 340
rect 1791 421 1891 573
rect 2287 541 2387 585
rect 2491 552 2591 585
rect 1791 375 1804 421
rect 1850 375 1891 421
rect 1791 340 1891 375
rect 2059 429 2131 442
rect 2287 434 2367 541
rect 2059 383 2072 429
rect 2118 383 2131 429
rect 2059 370 2131 383
rect 2247 421 2367 434
rect 2247 375 2276 421
rect 2322 375 2367 421
rect 1791 296 1911 340
rect 124 112 244 156
rect 348 112 468 156
rect 575 112 695 156
rect 799 64 919 156
rect 967 112 1087 156
rect 1191 64 1311 156
rect 1567 112 1687 156
rect 1791 112 1911 156
rect 2059 64 2099 370
rect 2247 316 2367 375
rect 2491 506 2504 552
rect 2550 506 2591 552
rect 2639 541 2739 585
rect 2491 360 2591 506
rect 2471 316 2591 360
rect 2695 360 2739 541
rect 3077 466 3177 573
rect 3281 466 3381 573
rect 3485 466 3585 573
rect 3689 466 3789 573
rect 3067 453 3859 466
rect 3067 407 3080 453
rect 3502 407 3859 453
rect 3067 394 3859 407
rect 2695 316 2815 360
rect 3067 333 3187 394
rect 3291 393 3859 394
rect 3291 333 3411 393
rect 3515 333 3635 393
rect 3739 333 3859 393
rect 799 24 2099 64
rect 2247 64 2367 156
rect 2471 112 2591 156
rect 2695 64 2815 156
rect 3067 89 3187 133
rect 3291 89 3411 133
rect 3515 89 3635 133
rect 3739 89 3859 133
rect 2247 24 2815 64
<< polycontact >>
rect 148 375 194 421
rect 469 375 515 421
rect 692 369 738 415
rect 905 446 951 492
rect 1604 375 1650 421
rect 1804 375 1850 421
rect 2072 383 2118 429
rect 2276 375 2322 421
rect 2504 506 2550 552
rect 3080 407 3502 453
<< metal1 >>
rect 0 918 4032 1098
rect 265 781 311 918
rect 812 781 858 792
rect 265 630 311 641
rect 142 421 194 542
rect 142 375 148 421
rect 142 354 194 375
rect 469 421 530 654
rect 812 584 858 641
rect 1164 781 1210 918
rect 1164 630 1210 641
rect 1256 826 1650 872
rect 1256 584 1302 826
rect 812 559 1302 584
rect 515 375 530 421
rect 469 364 530 375
rect 589 538 1302 559
rect 1368 769 1414 780
rect 589 513 853 538
rect 589 323 635 513
rect 894 446 905 492
rect 951 446 962 492
rect 894 415 962 446
rect 1368 415 1414 629
rect 681 369 692 415
rect 738 369 1414 415
rect 49 261 543 307
rect 589 277 770 323
rect 49 215 95 261
rect 497 215 543 261
rect 49 158 95 169
rect 262 169 273 215
rect 319 169 330 215
rect 262 90 330 169
rect 497 158 543 169
rect 724 215 770 277
rect 724 158 770 169
rect 1116 215 1162 226
rect 1116 90 1162 169
rect 1340 215 1414 369
rect 1386 169 1414 215
rect 1340 158 1414 169
rect 1492 769 1558 780
rect 1492 629 1512 769
rect 1492 318 1558 629
rect 1604 421 1650 826
rect 1716 781 1762 918
rect 2416 908 2462 918
rect 1716 630 1762 641
rect 1920 781 1966 792
rect 2416 757 2462 768
rect 2768 781 2814 792
rect 1966 711 2371 747
rect 1966 701 2550 711
rect 1966 641 1986 701
rect 2326 665 2550 701
rect 1604 364 1650 375
rect 1696 375 1804 421
rect 1850 375 1861 421
rect 1696 318 1742 375
rect 1492 272 1742 318
rect 1492 215 1538 272
rect 1492 158 1538 169
rect 1716 215 1762 226
rect 1716 90 1762 169
rect 1920 215 1986 641
rect 2172 644 2258 655
rect 2172 598 2212 644
rect 2172 587 2258 598
rect 2072 429 2118 440
rect 2072 292 2118 383
rect 2172 303 2218 587
rect 2504 552 2550 665
rect 2270 421 2322 542
rect 2504 495 2550 506
rect 2270 375 2276 421
rect 2270 354 2322 375
rect 2768 464 2814 641
rect 3002 781 3048 918
rect 3002 630 3048 641
rect 3206 781 3252 792
rect 3206 584 3252 641
rect 3410 781 3456 918
rect 3410 630 3456 641
rect 3614 781 3710 792
rect 3660 641 3710 781
rect 3614 584 3710 641
rect 3818 781 3864 918
rect 3818 630 3864 641
rect 3206 538 3710 584
rect 2768 453 3502 464
rect 2768 407 3080 453
rect 2768 396 3502 407
rect 2768 307 2814 396
rect 3614 320 3710 538
rect 2072 257 2172 292
rect 2609 303 2814 307
rect 2609 257 2620 303
rect 2666 261 2814 303
rect 2992 309 3038 320
rect 2666 257 2677 261
rect 2072 246 2218 257
rect 1920 169 1940 215
rect 1920 158 1986 169
rect 2396 215 2442 226
rect 2396 90 2442 169
rect 2844 215 2890 226
rect 2844 90 2890 169
rect 2992 90 3038 169
rect 3206 309 3710 320
rect 3206 169 3216 309
rect 3262 260 3664 309
rect 3206 158 3262 169
rect 3440 203 3486 214
rect 3664 158 3710 169
rect 3888 309 3934 320
rect 3440 90 3486 157
rect 3888 90 3934 169
rect 0 -90 4032 90
<< labels >>
flabel metal1 s 2270 354 2322 542 0 FreeSans 200 0 0 0 CLKN
port 1 nsew clock input
flabel metal1 s 469 364 530 654 0 FreeSans 200 0 0 0 E
port 2 nsew default input
flabel metal1 s 3614 584 3710 792 0 FreeSans 200 0 0 0 Q
port 4 nsew default output
flabel metal1 s 142 354 194 542 0 FreeSans 200 0 0 0 TE
port 3 nsew default input
flabel metal1 s 0 918 4032 1098 0 FreeSans 200 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 3888 226 3934 320 0 FreeSans 200 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 6 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 3206 584 3252 792 1 Q
port 4 nsew default output
rlabel metal1 s 3206 538 3710 584 1 Q
port 4 nsew default output
rlabel metal1 s 3614 320 3710 538 1 Q
port 4 nsew default output
rlabel metal1 s 3206 260 3710 320 1 Q
port 4 nsew default output
rlabel metal1 s 3664 158 3710 260 1 Q
port 4 nsew default output
rlabel metal1 s 3206 158 3262 260 1 Q
port 4 nsew default output
rlabel metal1 s 3818 757 3864 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3410 757 3456 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3002 757 3048 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2416 757 2462 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1716 757 1762 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1164 757 1210 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 265 757 311 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3818 630 3864 757 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3410 630 3456 757 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3002 630 3048 757 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1716 630 1762 757 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1164 630 1210 757 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 265 630 311 757 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2992 226 3038 320 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3888 215 3934 226 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2992 215 3038 226 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2844 215 2890 226 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2396 215 2442 226 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1716 215 1762 226 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1116 215 1162 226 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3888 214 3934 215 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2992 214 3038 215 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2844 214 2890 215 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2396 214 2442 215 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1716 214 1762 215 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1116 214 1162 215 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 262 214 330 215 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3888 90 3934 214 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3440 90 3486 214 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2992 90 3038 214 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2844 90 2890 214 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2396 90 2442 214 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1716 90 1762 214 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1116 90 1162 214 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 262 90 330 214 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 4032 90 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4032 1008
string GDS_END 845240
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 835988
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
