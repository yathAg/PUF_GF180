VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_fd_sc_mcu9t5v0__addf_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__addf_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.800 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.265 2.330 3.455 2.710 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 13.525 2.265 13.850 2.710 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.547000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.890 2.115 12.550 2.345 ;
        RECT 11.910 1.770 12.170 2.115 ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 15.830 2.890 16.475 3.685 ;
        RECT 16.145 0.845 16.475 2.890 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.324400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 0.845 0.575 3.830 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 16.800 5.490 ;
        RECT 1.365 3.875 1.595 4.590 ;
        RECT 6.625 3.610 6.855 4.590 ;
        RECT 8.665 3.140 8.895 4.590 ;
        RECT 10.705 3.505 10.935 4.590 ;
        RECT 15.125 3.875 15.355 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 17.230 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 17.230 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.305 ;
        RECT 6.625 0.450 6.855 1.425 ;
        RECT 8.865 0.450 9.095 1.425 ;
        RECT 10.705 0.450 10.935 1.425 ;
        RECT 15.125 0.450 15.355 1.165 ;
        RECT 0.000 -0.450 16.800 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 4.385 3.170 4.615 3.790 ;
        RECT 1.805 2.940 4.615 3.170 ;
        RECT 5.605 3.265 5.835 3.845 ;
        RECT 9.685 3.265 9.915 3.845 ;
        RECT 11.725 3.265 11.955 3.845 ;
        RECT 5.605 3.035 7.930 3.265 ;
        RECT 9.685 3.035 11.955 3.265 ;
        RECT 12.845 3.170 13.075 3.685 ;
        RECT 12.845 2.940 14.310 3.170 ;
        RECT 1.805 2.060 2.035 2.940 ;
        RECT 12.845 2.805 13.075 2.940 ;
        RECT 5.010 2.575 13.075 2.805 ;
        RECT 0.870 1.885 2.035 2.060 ;
        RECT 14.080 2.115 14.310 2.940 ;
        RECT 14.080 2.005 15.795 2.115 ;
        RECT 0.870 1.655 4.615 1.885 ;
        RECT 4.385 1.315 4.615 1.655 ;
        RECT 5.505 1.655 7.975 1.885 ;
        RECT 5.505 1.315 5.735 1.655 ;
        RECT 7.745 1.315 7.975 1.655 ;
        RECT 9.585 1.655 11.680 1.885 ;
        RECT 9.585 1.315 9.815 1.655 ;
        RECT 11.450 1.540 11.680 1.655 ;
        RECT 12.945 1.775 15.795 2.005 ;
        RECT 11.450 1.310 12.110 1.540 ;
        RECT 12.945 1.315 13.175 1.775 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__addf_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__addf_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__addf_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.040 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.700000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.425 2.330 4.605 2.710 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.700000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.710 2.150 16.110 2.710 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.525000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.050 1.920 13.850 2.150 ;
        RECT 13.590 1.770 13.850 1.920 ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.622400 ;
    PORT
      LAYER Metal1 ;
        RECT 17.165 2.710 17.395 3.685 ;
        RECT 17.165 0.845 17.770 2.710 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.622400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 0.845 1.855 3.830 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 19.040 5.490 ;
        RECT 0.605 3.845 0.835 4.590 ;
        RECT 2.645 3.845 2.875 4.590 ;
        RECT 7.785 3.905 8.015 4.590 ;
        RECT 10.025 3.435 10.255 4.590 ;
        RECT 11.765 3.435 11.995 4.590 ;
        RECT 15.965 3.905 16.195 4.590 ;
        RECT 18.185 3.845 18.415 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 19.470 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 19.470 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.285 0.450 0.515 1.165 ;
        RECT 2.525 0.450 2.755 1.165 ;
        RECT 7.785 0.450 8.015 1.215 ;
        RECT 10.025 0.450 10.255 1.215 ;
        RECT 11.865 0.450 12.095 1.215 ;
        RECT 16.265 0.450 16.495 1.195 ;
        RECT 18.505 0.450 18.735 1.165 ;
        RECT 0.000 -0.450 19.040 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 5.545 3.170 5.775 3.685 ;
        RECT 2.965 2.940 5.775 3.170 ;
        RECT 8.805 3.160 9.035 3.740 ;
        RECT 2.965 2.115 3.195 2.940 ;
        RECT 5.545 2.875 5.775 2.940 ;
        RECT 6.710 2.930 9.035 3.160 ;
        RECT 10.745 3.160 10.975 3.740 ;
        RECT 12.885 3.160 13.115 3.740 ;
        RECT 10.745 2.930 13.115 3.160 ;
        RECT 14.105 2.985 16.935 3.215 ;
        RECT 14.105 2.700 14.335 2.985 ;
        RECT 6.070 2.470 14.335 2.700 ;
        RECT 2.085 1.775 3.195 2.115 ;
        RECT 2.965 1.600 3.195 1.775 ;
        RECT 2.965 1.370 5.830 1.600 ;
        RECT 6.665 1.445 9.135 1.675 ;
        RECT 6.665 1.315 6.895 1.445 ;
        RECT 8.905 1.315 9.135 1.445 ;
        RECT 10.745 1.445 13.215 1.675 ;
        RECT 16.705 1.655 16.935 2.985 ;
        RECT 10.745 1.315 10.975 1.445 ;
        RECT 12.985 1.315 13.215 1.445 ;
        RECT 14.050 1.425 16.935 1.655 ;
        RECT 14.050 1.370 14.390 1.425 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__addf_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__addf_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__addf_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.700000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.705 1.860 6.785 2.710 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.700000 ;
    PORT
      LAYER Metal1 ;
        RECT 16.965 2.330 18.530 2.710 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.525000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.330 1.920 15.990 2.150 ;
        RECT 11.910 1.770 12.170 1.920 ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.642000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.635 3.105 19.865 3.685 ;
        RECT 21.875 3.105 22.105 3.685 ;
        RECT 19.635 2.875 22.105 3.105 ;
        RECT 20.725 1.655 21.185 2.875 ;
        RECT 19.685 1.425 22.155 1.655 ;
        RECT 19.685 0.845 19.915 1.425 ;
        RECT 21.925 0.845 22.155 1.425 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.815850 ;
    PORT
      LAYER Metal1 ;
        RECT 1.445 3.105 1.675 3.685 ;
        RECT 3.785 3.105 4.015 3.685 ;
        RECT 1.445 2.875 4.015 3.105 ;
        RECT 2.380 1.655 2.840 2.875 ;
        RECT 1.445 1.425 3.915 1.655 ;
        RECT 1.445 0.845 1.675 1.425 ;
        RECT 3.685 0.845 3.915 1.425 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 23.520 5.490 ;
        RECT 0.325 3.875 0.555 4.590 ;
        RECT 2.555 3.875 2.785 4.590 ;
        RECT 4.905 3.875 5.135 4.590 ;
        RECT 10.065 3.905 10.295 4.590 ;
        RECT 12.205 3.435 12.435 4.590 ;
        RECT 14.145 3.435 14.375 4.590 ;
        RECT 18.465 3.875 18.695 4.590 ;
        RECT 20.750 3.875 20.980 4.590 ;
        RECT 22.945 3.875 23.175 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 23.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 23.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.325 0.450 0.555 1.165 ;
        RECT 2.565 0.450 2.795 1.165 ;
        RECT 4.805 0.450 5.035 1.165 ;
        RECT 10.065 0.450 10.295 1.215 ;
        RECT 12.305 0.450 12.535 1.215 ;
        RECT 14.145 0.450 14.375 1.215 ;
        RECT 18.565 0.450 18.795 1.165 ;
        RECT 20.805 0.450 21.035 1.165 ;
        RECT 23.045 0.450 23.275 1.165 ;
        RECT 0.000 -0.450 23.520 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 7.825 3.170 8.055 3.685 ;
        RECT 5.245 2.940 8.055 3.170 ;
        RECT 4.310 2.060 4.595 2.585 ;
        RECT 5.245 2.060 5.475 2.940 ;
        RECT 7.825 2.875 8.055 2.940 ;
        RECT 9.045 3.160 9.275 3.740 ;
        RECT 13.125 3.160 13.355 3.740 ;
        RECT 15.165 3.160 15.395 3.740 ;
        RECT 16.285 3.170 16.515 3.750 ;
        RECT 9.045 2.930 11.370 3.160 ;
        RECT 13.125 2.930 15.395 3.160 ;
        RECT 15.625 2.940 19.235 3.170 ;
        RECT 15.625 2.700 15.855 2.940 ;
        RECT 8.450 2.470 15.855 2.700 ;
        RECT 4.310 1.830 5.475 2.060 ;
        RECT 19.005 2.005 19.235 2.940 ;
        RECT 5.245 1.545 5.475 1.830 ;
        RECT 16.385 1.775 19.235 2.005 ;
        RECT 5.245 1.315 8.110 1.545 ;
        RECT 8.945 1.445 11.415 1.675 ;
        RECT 8.945 1.315 9.175 1.445 ;
        RECT 11.185 1.315 11.415 1.445 ;
        RECT 13.025 1.445 15.495 1.675 ;
        RECT 13.025 1.315 13.255 1.445 ;
        RECT 15.265 1.315 15.495 1.445 ;
        RECT 16.385 1.315 16.615 1.775 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__addf_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__addh_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__addh_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.285 2.950 6.075 3.270 ;
        RECT 2.285 2.215 2.515 2.950 ;
        RECT 5.845 2.215 6.075 2.950 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 2.270 5.195 2.650 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 0.845 0.575 4.360 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.845 1.590 9.175 4.360 ;
        RECT 8.550 1.210 9.175 1.590 ;
        RECT 8.945 0.845 9.175 1.210 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 9.520 5.490 ;
        RECT 1.365 3.550 1.595 4.590 ;
        RECT 3.645 3.960 3.875 4.590 ;
        RECT 4.385 3.960 4.615 4.590 ;
        RECT 7.645 3.550 7.875 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 9.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.350 ;
        RECT 7.645 0.450 7.875 1.355 ;
        RECT 0.000 -0.450 9.520 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 2.625 3.730 2.855 4.360 ;
        RECT 6.570 3.960 7.415 4.190 ;
        RECT 1.825 3.500 6.955 3.730 ;
        RECT 1.825 2.555 2.055 3.500 ;
        RECT 0.925 2.215 2.055 2.555 ;
        RECT 6.725 2.500 6.955 3.500 ;
        RECT 7.185 3.320 7.415 3.960 ;
        RECT 7.185 3.090 7.810 3.320 ;
        RECT 7.580 2.555 7.810 3.090 ;
        RECT 6.725 2.270 7.350 2.500 ;
        RECT 1.825 1.300 2.055 2.215 ;
        RECT 7.580 2.215 8.495 2.555 ;
        RECT 7.580 1.985 7.810 2.215 ;
        RECT 5.405 1.755 7.810 1.985 ;
        RECT 1.825 1.070 3.850 1.300 ;
        RECT 4.285 0.910 4.515 1.355 ;
        RECT 5.405 1.140 5.635 1.755 ;
        RECT 6.525 0.910 6.755 1.355 ;
        RECT 4.285 0.680 6.755 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__addh_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__addh_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__addh_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.760 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.610 2.940 6.010 3.170 ;
        RECT 3.610 2.500 3.840 2.940 ;
        RECT 3.030 2.270 3.840 2.500 ;
        RECT 5.750 2.500 6.010 2.940 ;
        RECT 5.750 2.270 7.160 2.500 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.070 2.150 4.330 2.710 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.821000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 0.770 1.615 4.355 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.729500 ;
    PORT
      LAYER Metal1 ;
        RECT 9.985 1.590 10.215 4.355 ;
        RECT 9.985 0.770 10.490 1.590 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 11.760 5.490 ;
        RECT 0.315 3.875 0.545 4.590 ;
        RECT 2.455 3.875 2.685 4.590 ;
        RECT 4.545 3.875 4.775 4.590 ;
        RECT 5.365 3.875 5.595 4.590 ;
        RECT 8.865 3.875 9.095 4.590 ;
        RECT 11.055 3.875 11.285 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 12.190 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.190 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.265 0.450 0.495 1.580 ;
        RECT 2.505 0.450 2.735 1.580 ;
        RECT 8.865 0.450 9.095 1.580 ;
        RECT 11.105 0.450 11.335 1.580 ;
        RECT 0.000 -0.450 11.760 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.525 3.630 3.755 4.325 ;
        RECT 7.505 3.875 8.635 4.215 ;
        RECT 2.570 3.400 8.175 3.630 ;
        RECT 2.570 2.665 2.800 3.400 ;
        RECT 2.015 2.385 2.800 2.665 ;
        RECT 2.015 1.855 2.245 2.385 ;
        RECT 7.945 2.040 8.175 3.400 ;
        RECT 4.545 1.810 8.175 2.040 ;
        RECT 8.405 2.645 8.635 3.875 ;
        RECT 8.405 2.270 9.635 2.645 ;
        RECT 4.545 0.770 4.775 1.810 ;
        RECT 5.265 0.910 5.495 1.580 ;
        RECT 8.405 1.570 8.635 2.270 ;
        RECT 9.400 1.835 9.635 2.270 ;
        RECT 6.385 1.340 8.635 1.570 ;
        RECT 6.385 1.140 6.615 1.340 ;
        RECT 7.505 0.910 7.735 1.110 ;
        RECT 5.265 0.680 7.735 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__addh_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__addh_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__addh_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.300000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.100 2.630 8.080 2.860 ;
        RECT 1.100 2.215 1.330 2.630 ;
        RECT 3.930 2.285 6.450 2.630 ;
        RECT 7.850 2.500 8.080 2.630 ;
        RECT 7.850 2.270 9.860 2.500 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.300000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.770 2.055 3.050 2.400 ;
        RECT 6.680 2.170 7.620 2.400 ;
        RECT 6.680 2.055 6.910 2.170 ;
        RECT 1.770 1.825 6.910 2.055 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.550500 ;
    PORT
      LAYER Metal1 ;
        RECT 12.470 2.985 15.100 3.215 ;
        RECT 12.470 1.595 12.805 2.985 ;
        RECT 12.470 1.365 15.150 1.595 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.660300 ;
    PORT
      LAYER Metal1 ;
        RECT 16.950 3.320 17.235 4.360 ;
        RECT 19.205 3.320 19.435 4.360 ;
        RECT 16.950 2.960 19.435 3.320 ;
        RECT 19.075 1.790 19.435 2.960 ;
        RECT 16.950 1.430 19.575 1.790 ;
        RECT 16.950 0.695 17.335 1.430 ;
        RECT 19.345 0.695 19.575 1.430 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 21.280 5.490 ;
        RECT 0.295 3.550 0.525 4.590 ;
        RECT 2.335 3.550 2.565 4.590 ;
        RECT 4.425 3.550 4.655 4.590 ;
        RECT 7.915 4.010 8.145 4.590 ;
        RECT 11.275 4.010 11.505 4.590 ;
        RECT 13.695 4.010 13.925 4.590 ;
        RECT 15.885 3.550 16.115 4.590 ;
        RECT 18.125 3.550 18.355 4.590 ;
        RECT 20.335 3.550 20.565 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 21.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 21.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.200 ;
        RECT 4.425 0.450 4.655 1.595 ;
        RECT 11.505 0.675 11.735 1.125 ;
        RECT 15.985 0.675 16.215 1.200 ;
        RECT 11.505 0.450 16.215 0.675 ;
        RECT 18.225 0.450 18.455 1.200 ;
        RECT 20.465 0.450 20.695 1.200 ;
        RECT 0.000 -0.450 21.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.315 3.320 1.545 4.360 ;
        RECT 3.405 3.320 3.635 4.360 ;
        RECT 5.725 3.780 5.955 4.360 ;
        RECT 10.155 3.780 10.385 4.360 ;
        RECT 5.725 3.550 15.610 3.780 ;
        RECT 0.640 3.090 10.320 3.320 ;
        RECT 0.640 1.595 0.870 3.090 ;
        RECT 10.090 2.500 10.320 3.090 ;
        RECT 15.380 2.555 15.610 3.550 ;
        RECT 10.090 2.270 12.230 2.500 ;
        RECT 15.380 2.215 18.590 2.555 ;
        RECT 0.640 1.365 2.615 1.595 ;
        RECT 2.385 0.695 2.615 1.365 ;
        RECT 6.790 1.355 12.195 1.585 ;
        RECT 11.965 1.135 12.195 1.355 ;
        RECT 15.380 1.135 15.610 2.215 ;
        RECT 5.670 0.845 10.490 1.075 ;
        RECT 11.965 0.905 15.610 1.135 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__addh_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__and2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.806000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.710 0.970 2.960 ;
        RECT 0.115 2.150 0.970 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.806000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 2.710 2.060 2.960 ;
        RECT 1.830 2.150 2.715 2.710 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 0.845 3.855 3.685 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 4.480 5.490 ;
        RECT 0.245 4.345 0.475 4.590 ;
        RECT 2.285 4.345 2.515 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 4.910 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.505 0.450 2.735 1.165 ;
        RECT 0.000 -0.450 4.480 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.210 4.115 1.550 4.170 ;
        RECT 1.210 3.885 3.175 4.115 ;
        RECT 2.945 1.625 3.175 3.885 ;
        RECT 0.190 1.395 3.175 1.625 ;
        RECT 0.190 1.370 0.530 1.395 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and2_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__and2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.040 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.612000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.330 0.970 2.715 ;
        RECT 0.710 1.905 0.970 2.330 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.612000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 2.330 2.090 2.710 ;
        RECT 1.830 1.900 2.090 2.330 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.420 0.845 3.770 3.685 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.040 5.490 ;
        RECT 0.260 3.685 0.490 4.590 ;
        RECT 2.520 3.875 2.750 4.590 ;
        RECT 4.560 3.875 4.790 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 5.470 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 5.470 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.300 0.450 2.530 1.165 ;
        RECT 4.540 0.450 4.770 1.165 ;
        RECT 0.000 -0.450 5.040 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.280 3.170 1.510 3.750 ;
        RECT 1.280 2.940 2.970 3.170 ;
        RECT 2.740 1.655 2.970 2.940 ;
        RECT 0.260 1.425 2.970 1.655 ;
        RECT 0.260 0.845 0.490 1.425 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and2_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__and2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.224000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.205 1.210 2.090 2.060 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.224000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.355 2.290 4.030 2.715 ;
        RECT 0.355 1.770 0.970 2.290 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.445 2.790 8.085 3.685 ;
        RECT 7.485 1.600 8.085 2.790 ;
        RECT 5.390 0.900 8.085 1.600 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 9.520 5.490 ;
        RECT 0.245 3.875 0.475 4.590 ;
        RECT 2.285 3.875 2.515 4.590 ;
        RECT 4.325 3.875 4.555 4.590 ;
        RECT 6.545 4.230 6.775 4.590 ;
        RECT 8.585 4.225 8.815 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 9.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.165 ;
        RECT 4.325 0.450 4.555 1.165 ;
        RECT 6.510 0.450 6.850 0.640 ;
        RECT 8.805 0.450 9.035 1.165 ;
        RECT 0.000 -0.450 9.520 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.265 3.180 1.495 3.875 ;
        RECT 3.305 3.180 3.535 3.875 ;
        RECT 1.265 2.950 4.995 3.180 ;
        RECT 4.765 2.315 4.995 2.950 ;
        RECT 4.765 1.975 6.465 2.315 ;
        RECT 4.765 1.655 4.995 1.975 ;
        RECT 2.320 1.425 4.995 1.655 ;
        RECT 2.320 0.845 2.550 1.425 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and2_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__and3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.761000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 2.740 1.145 3.345 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.761000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.820 2.740 2.725 3.375 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.761000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.565 1.770 2.955 2.150 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.630 0.845 4.995 3.830 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.600 5.490 ;
        RECT 1.265 4.345 1.495 4.590 ;
        RECT 3.645 4.345 3.875 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 3.645 0.450 3.875 1.350 ;
        RECT 0.000 -0.450 5.600 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 4.115 0.475 4.315 ;
        RECT 2.285 4.115 3.415 4.315 ;
        RECT 0.245 3.885 3.415 4.115 ;
        RECT 3.185 2.115 3.415 3.885 ;
        RECT 3.185 1.775 4.315 2.115 ;
        RECT 0.245 0.980 0.475 1.355 ;
        RECT 3.185 0.980 3.415 1.775 ;
        RECT 0.245 0.750 3.415 0.980 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and3_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__and3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.160 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.115 2.150 0.970 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.210 2.150 2.090 2.710 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.390 2.290 3.210 2.710 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.480 0.845 4.890 3.685 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 6.160 5.490 ;
        RECT 1.320 3.875 1.550 4.590 ;
        RECT 3.360 3.875 3.590 4.590 ;
        RECT 5.580 3.875 5.810 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.590 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.590 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 3.360 0.450 3.590 1.165 ;
        RECT 5.600 0.450 5.830 1.165 ;
        RECT 0.000 -0.450 6.160 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 2.340 3.530 2.570 4.110 ;
        RECT 0.245 3.300 4.210 3.530 ;
        RECT 3.980 1.920 4.210 3.300 ;
        RECT 0.300 1.690 4.210 1.920 ;
        RECT 0.300 0.845 0.530 1.690 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and3_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__and3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.200 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.245 1.730 3.115 2.150 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.790 2.380 5.000 2.610 ;
        RECT 3.995 1.770 5.000 2.380 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.840 6.020 3.070 ;
        RECT 0.150 2.330 0.995 2.840 ;
        RECT 5.785 2.415 6.020 2.840 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.550 2.925 9.930 3.630 ;
        RECT 9.580 1.600 9.930 2.925 ;
        RECT 7.250 0.895 9.930 1.600 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 11.200 5.490 ;
        RECT 0.245 3.505 0.475 4.590 ;
        RECT 2.285 3.975 2.515 4.590 ;
        RECT 4.325 3.975 4.555 4.590 ;
        RECT 6.585 3.875 6.815 4.590 ;
        RECT 8.625 3.875 8.855 4.590 ;
        RECT 10.665 3.875 10.895 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 11.630 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 11.630 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.325 0.450 0.555 0.695 ;
        RECT 6.185 0.450 6.415 1.165 ;
        RECT 8.370 0.450 8.710 0.640 ;
        RECT 10.665 0.450 10.895 1.165 ;
        RECT 0.000 -0.450 11.200 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.265 3.530 1.495 4.110 ;
        RECT 3.305 3.530 3.535 4.110 ;
        RECT 5.345 3.530 5.575 4.110 ;
        RECT 1.265 3.300 6.855 3.530 ;
        RECT 6.625 2.310 6.855 3.300 ;
        RECT 6.625 1.970 9.260 2.310 ;
        RECT 6.625 1.625 6.855 1.970 ;
        RECT 5.500 1.520 6.855 1.625 ;
        RECT 3.305 1.395 6.855 1.520 ;
        RECT 3.305 1.290 5.755 1.395 ;
        RECT 3.305 0.710 3.535 1.290 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and3_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__and4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.160 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.716000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.115 2.165 0.975 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.716000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.230 1.210 2.090 2.115 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.716000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.320 1.210 3.210 2.115 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.716000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.830 2.330 4.500 2.710 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.190 2.890 6.045 3.685 ;
        RECT 5.585 0.845 6.045 2.890 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 6.160 5.490 ;
        RECT 0.305 3.155 0.535 4.590 ;
        RECT 2.345 3.155 2.575 4.590 ;
        RECT 4.565 4.345 4.795 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.590 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.590 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 4.565 0.450 4.795 1.350 ;
        RECT 0.000 -0.450 6.160 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.325 2.925 1.555 3.215 ;
        RECT 3.365 2.985 4.960 3.215 ;
        RECT 3.365 2.925 3.595 2.985 ;
        RECT 1.325 2.695 3.595 2.925 ;
        RECT 4.730 2.115 4.960 2.985 ;
        RECT 4.730 2.005 5.235 2.115 ;
        RECT 3.440 1.775 5.235 2.005 ;
        RECT 0.305 0.980 0.535 1.355 ;
        RECT 3.440 0.980 3.670 1.775 ;
        RECT 0.305 0.750 3.670 0.980 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and4_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__and4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.115 2.150 0.970 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.200 2.150 2.090 2.710 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.320 2.290 3.210 2.710 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.440 2.330 4.330 2.710 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.580 1.725 6.100 3.685 ;
        RECT 5.190 0.845 6.100 1.725 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.280 5.490 ;
        RECT 0.300 3.875 0.530 4.590 ;
        RECT 2.340 4.345 2.570 4.590 ;
        RECT 4.380 3.875 4.610 4.590 ;
        RECT 6.600 3.875 6.830 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 7.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 4.380 0.450 4.610 0.695 ;
        RECT 6.620 0.450 6.850 1.165 ;
        RECT 0.000 -0.450 7.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.360 3.765 3.590 4.235 ;
        RECT 1.320 3.645 3.590 3.765 ;
        RECT 1.320 3.415 4.790 3.645 ;
        RECT 4.560 2.720 4.790 3.415 ;
        RECT 4.560 2.380 5.230 2.720 ;
        RECT 4.560 1.600 4.790 2.380 ;
        RECT 0.245 1.370 4.790 1.600 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and4_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__and4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and4_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.440 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.790 1.770 3.890 2.150 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.825 2.380 4.750 2.610 ;
        RECT 4.520 2.150 4.750 2.380 ;
        RECT 4.520 1.770 6.030 2.150 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.975 1.540 2.145 2.060 ;
        RECT 6.260 1.830 7.105 2.060 ;
        RECT 6.260 1.540 6.490 1.830 ;
        RECT 0.975 1.310 6.490 1.540 ;
        RECT 0.975 1.210 2.090 1.310 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.115 2.840 5.210 3.070 ;
        RECT 0.115 2.330 0.970 2.840 ;
        RECT 4.980 2.700 5.210 2.840 ;
        RECT 4.980 2.470 8.125 2.700 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.540 2.920 12.210 3.640 ;
        RECT 11.770 1.600 12.210 2.920 ;
        RECT 9.485 0.900 12.210 1.600 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 13.440 5.490 ;
        RECT 0.260 3.325 0.490 4.590 ;
        RECT 2.300 3.795 2.530 4.590 ;
        RECT 4.340 3.795 4.570 4.590 ;
        RECT 6.380 3.795 6.610 4.590 ;
        RECT 8.420 3.795 8.650 4.590 ;
        RECT 10.640 3.875 10.870 4.590 ;
        RECT 12.680 3.875 12.910 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 13.870 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 13.870 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.260 0.450 0.490 1.165 ;
        RECT 8.420 0.450 8.650 0.695 ;
        RECT 10.605 0.450 10.945 0.640 ;
        RECT 12.900 0.450 13.130 1.165 ;
        RECT 0.000 -0.450 13.440 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.280 3.530 1.510 4.110 ;
        RECT 3.320 3.530 3.550 4.110 ;
        RECT 5.360 3.530 5.590 4.110 ;
        RECT 1.280 3.430 5.590 3.530 ;
        RECT 7.400 3.430 7.630 4.010 ;
        RECT 1.280 3.300 9.090 3.430 ;
        RECT 5.400 3.200 9.090 3.300 ;
        RECT 8.860 2.315 9.090 3.200 ;
        RECT 8.860 1.975 10.550 2.315 ;
        RECT 8.860 1.260 9.090 1.975 ;
        RECT 6.715 1.080 9.090 1.260 ;
        RECT 4.285 1.030 9.090 1.080 ;
        RECT 4.285 0.850 6.940 1.030 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and4_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__antenna
  CLASS core ANTENNACELL ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__antenna ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.120 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNADIFFAREA 0.406800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 1.315 0.475 3.215 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 1.120 5.490 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 1.550 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 1.550 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.450 1.120 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__antenna

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi21_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi21_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 2.415 2.655 3.270 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.115 2.285 0.970 2.710 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.467000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 1.805 3.780 2.815 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.755600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 2.150 1.495 3.685 ;
        RECT 1.265 1.770 2.515 2.150 ;
        RECT 2.285 0.845 2.515 1.770 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 4.480 5.490 ;
        RECT 3.485 3.875 3.715 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 4.910 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.165 ;
        RECT 3.585 0.450 3.815 1.565 ;
        RECT 0.000 -0.450 4.480 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 4.130 2.515 4.360 ;
        RECT 0.245 3.550 0.475 4.130 ;
        RECT 2.285 3.550 2.515 4.130 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi21_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi21_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi21_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.000 1.755 5.120 2.300 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.410 2.560 6.605 2.790 ;
        RECT 3.410 1.770 3.660 2.560 ;
        RECT 5.690 2.155 6.605 2.560 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.934000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.115 1.665 0.980 2.150 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.287600 ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 3.250 3.700 3.830 ;
        RECT 5.630 3.250 5.860 3.830 ;
        RECT 2.330 3.020 5.860 3.250 ;
        RECT 2.330 1.490 2.715 3.020 ;
        RECT 2.330 1.155 4.920 1.490 ;
        RECT 1.375 0.925 4.920 1.155 ;
        RECT 3.010 0.680 4.920 0.925 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.280 5.490 ;
        RECT 1.330 4.345 1.560 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 7.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.310 0.450 0.540 1.165 ;
        RECT 2.550 0.450 2.780 0.695 ;
        RECT 6.650 0.450 6.880 1.165 ;
        RECT 0.000 -0.450 7.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.310 3.765 0.540 4.360 ;
        RECT 2.445 4.060 6.880 4.290 ;
        RECT 2.445 3.765 2.680 4.060 ;
        RECT 0.310 3.480 2.680 3.765 ;
        RECT 4.610 3.480 4.840 4.060 ;
        RECT 6.650 3.480 6.880 4.060 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi21_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi21_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi21_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.440 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.615 2.135 2.845 ;
        RECT 0.710 1.570 0.970 2.615 ;
        RECT 1.905 2.420 2.135 2.615 ;
        RECT 5.665 1.570 5.895 2.110 ;
        RECT 0.710 1.325 5.895 1.570 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.430 2.475 8.310 2.710 ;
        RECT 1.200 2.190 1.430 2.385 ;
        RECT 3.430 2.190 4.365 2.475 ;
        RECT 1.200 1.960 4.365 2.190 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.868000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.630 2.330 12.735 2.750 ;
        RECT 12.470 2.150 12.730 2.330 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.136000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.410 3.305 1.695 3.835 ;
        RECT 3.505 3.305 3.735 3.835 ;
        RECT 5.545 3.305 5.775 3.885 ;
        RECT 7.585 3.305 7.815 3.885 ;
        RECT 1.410 3.245 7.815 3.305 ;
        RECT 1.410 3.075 8.830 3.245 ;
        RECT 7.580 3.015 8.830 3.075 ;
        RECT 8.550 2.020 8.830 3.015 ;
        RECT 8.550 2.000 12.075 2.020 ;
        RECT 6.345 1.790 12.075 2.000 ;
        RECT 6.345 1.770 9.835 1.790 ;
        RECT 6.345 1.095 6.575 1.770 ;
        RECT 2.370 0.865 6.575 1.095 ;
        RECT 9.605 0.840 9.835 1.770 ;
        RECT 11.845 0.840 12.075 1.790 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 13.440 5.490 ;
        RECT 9.850 3.935 10.190 4.590 ;
        RECT 11.890 3.935 12.230 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 13.870 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 13.870 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.465 0.450 0.695 0.690 ;
        RECT 4.330 0.450 4.670 0.635 ;
        RECT 8.305 0.450 8.535 1.085 ;
        RECT 10.725 0.450 10.955 1.560 ;
        RECT 12.965 0.450 13.195 1.560 ;
        RECT 0.000 -0.450 13.440 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.445 4.115 8.880 4.345 ;
        RECT 0.445 3.535 0.675 4.115 ;
        RECT 2.485 3.535 2.715 4.115 ;
        RECT 4.525 3.535 4.755 4.115 ;
        RECT 6.565 3.535 6.795 4.115 ;
        RECT 8.550 3.705 8.880 4.115 ;
        RECT 10.870 3.705 11.210 4.230 ;
        RECT 12.910 3.705 13.250 4.230 ;
        RECT 8.550 3.475 13.250 3.705 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi21_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi22_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi22_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.040 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.930 1.210 3.830 2.115 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.950 2.330 4.915 2.710 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.250 1.210 2.090 2.115 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.130 2.175 0.980 2.710 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.365 3.355 3.600 3.830 ;
        RECT 2.350 2.855 3.600 3.355 ;
        RECT 2.350 0.845 2.580 2.855 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.040 5.490 ;
        RECT 1.330 3.875 1.560 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 5.470 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 5.470 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.310 0.450 0.540 1.165 ;
        RECT 4.390 0.450 4.620 1.165 ;
        RECT 0.000 -0.450 5.040 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.310 3.645 0.540 4.360 ;
        RECT 1.820 4.060 4.620 4.290 ;
        RECT 1.820 3.645 2.050 4.060 ;
        RECT 0.310 3.410 2.050 3.645 ;
        RECT 4.390 3.480 4.620 4.060 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi22_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi22_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi22_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.960 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 1.720 7.210 2.315 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.950 2.560 8.270 2.790 ;
        RECT 4.950 1.830 5.510 2.560 ;
        RECT 7.860 2.180 8.270 2.560 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.650 1.630 2.090 2.060 ;
        RECT 1.220 1.210 2.090 1.630 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.690 2.290 4.030 2.520 ;
        RECT 0.690 1.770 0.970 2.290 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.322200 ;
    PORT
      LAYER Metal1 ;
        RECT 4.345 3.250 5.575 3.830 ;
        RECT 7.385 3.250 7.615 3.830 ;
        RECT 4.345 3.020 7.615 3.250 ;
        RECT 4.345 1.490 4.720 3.020 ;
        RECT 2.320 1.105 2.550 1.490 ;
        RECT 4.340 1.105 4.720 1.490 ;
        RECT 6.365 1.105 6.595 1.490 ;
        RECT 2.320 0.875 6.595 1.105 ;
        RECT 2.320 0.680 2.550 0.875 ;
        RECT 6.365 0.680 6.595 0.875 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 8.960 5.490 ;
        RECT 1.265 3.875 1.495 4.590 ;
        RECT 3.305 3.875 3.535 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 9.390 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.390 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.165 ;
        RECT 4.270 0.450 4.610 0.640 ;
        RECT 8.405 0.450 8.635 1.165 ;
        RECT 0.000 -0.450 8.960 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.645 0.475 4.225 ;
        RECT 2.285 3.645 2.515 4.225 ;
        RECT 3.795 4.060 8.635 4.290 ;
        RECT 3.795 3.645 4.025 4.060 ;
        RECT 0.245 3.415 4.025 3.645 ;
        RECT 6.365 3.480 6.595 4.060 ;
        RECT 8.405 3.480 8.635 4.060 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi22_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi22_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi22_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.360 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 11.440 2.710 14.415 2.860 ;
        RECT 11.210 2.630 14.415 2.710 ;
        RECT 11.210 2.270 11.660 2.630 ;
        RECT 14.185 2.215 14.415 2.630 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.325 2.000 9.555 2.555 ;
        RECT 12.470 2.000 13.415 2.400 ;
        RECT 9.325 1.770 13.415 2.000 ;
        RECT 13.185 0.910 13.415 1.770 ;
        RECT 16.125 0.910 16.355 2.555 ;
        RECT 13.185 0.680 16.355 0.910 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.810 2.785 4.435 3.015 ;
        RECT 2.810 2.270 3.210 2.785 ;
        RECT 4.205 2.500 4.435 2.785 ;
        RECT 4.205 2.270 6.070 2.500 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.000 0.915 2.555 ;
        RECT 3.745 2.000 3.975 2.555 ;
        RECT 7.485 2.215 7.955 2.555 ;
        RECT 7.485 2.000 7.715 2.215 ;
        RECT 0.150 1.770 7.715 2.000 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.552000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.865 3.310 9.895 3.900 ;
        RECT 11.705 3.320 11.935 3.900 ;
        RECT 13.745 3.320 13.975 3.900 ;
        RECT 15.270 3.320 16.015 3.900 ;
        RECT 11.195 3.315 16.015 3.320 ;
        RECT 10.965 3.310 16.015 3.315 ;
        RECT 8.865 3.090 16.015 3.310 ;
        RECT 8.865 3.080 11.245 3.090 ;
        RECT 8.865 1.985 9.095 3.080 ;
        RECT 7.945 1.755 9.095 1.985 ;
        RECT 7.945 1.540 8.175 1.755 ;
        RECT 2.285 1.310 8.175 1.540 ;
        RECT 8.865 1.540 9.095 1.755 ;
        RECT 2.285 0.730 2.515 1.310 ;
        RECT 6.365 0.730 6.595 1.310 ;
        RECT 8.865 0.730 10.915 1.540 ;
        RECT 14.765 1.140 14.995 3.090 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.360 5.490 ;
        RECT 1.265 3.245 1.495 4.590 ;
        RECT 3.305 3.705 3.535 4.590 ;
        RECT 5.345 3.705 5.575 4.590 ;
        RECT 7.385 3.705 7.615 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 17.790 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 17.790 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.540 ;
        RECT 4.325 0.450 4.555 1.070 ;
        RECT 8.405 0.450 8.635 1.525 ;
        RECT 12.725 0.450 12.955 1.540 ;
        RECT 16.805 0.450 17.035 1.540 ;
        RECT 0.000 -0.450 17.360 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 8.405 4.130 17.035 4.360 ;
        RECT 0.245 3.015 0.475 4.055 ;
        RECT 2.150 3.475 2.515 4.055 ;
        RECT 4.325 3.475 4.555 4.055 ;
        RECT 6.365 3.475 6.595 4.055 ;
        RECT 8.405 3.475 8.635 4.130 ;
        RECT 10.685 3.540 10.915 4.130 ;
        RECT 12.725 3.550 12.955 4.130 ;
        RECT 14.765 3.550 14.995 4.130 ;
        RECT 2.150 3.245 8.635 3.475 ;
        RECT 16.805 3.245 17.035 4.130 ;
        RECT 2.150 3.015 2.380 3.245 ;
        RECT 0.245 2.785 2.380 3.015 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi22_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi211_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi211_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.626000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.770 1.210 2.695 2.115 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.626000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.115 1.705 0.970 2.595 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.925 1.615 3.815 2.150 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.045 1.615 4.915 2.150 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.010200 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 0.980 1.530 3.830 ;
        RECT 3.050 1.060 4.860 1.290 ;
        RECT 3.050 0.980 3.280 1.060 ;
        RECT 1.270 0.750 3.280 0.980 ;
        RECT 4.630 0.920 4.860 1.060 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.600 5.490 ;
        RECT 4.530 3.875 4.760 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 0.450 0.480 1.300 ;
        RECT 3.510 0.450 3.740 0.830 ;
        RECT 0.000 -0.450 5.600 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.250 4.130 2.520 4.360 ;
        RECT 0.250 3.550 0.480 4.130 ;
        RECT 2.290 3.550 2.520 4.130 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi211_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi211_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi211_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.252000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.765 1.770 2.955 2.215 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.252000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 2.445 3.770 2.775 ;
        RECT 0.630 2.305 1.155 2.445 ;
        RECT 3.510 1.770 3.770 2.445 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.560 2.470 8.430 2.700 ;
        RECT 4.560 1.725 5.450 2.470 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 1.770 7.295 2.150 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.341000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.210 3.400 4.330 3.630 ;
        RECT 4.070 1.525 4.330 3.400 ;
        RECT 2.205 1.495 4.330 1.525 ;
        RECT 2.205 1.265 4.960 1.495 ;
        RECT 2.205 0.715 2.435 1.265 ;
        RECT 4.730 1.160 4.960 1.265 ;
        RECT 4.730 0.930 7.935 1.160 ;
        RECT 5.465 0.695 5.695 0.930 ;
        RECT 7.705 0.790 7.935 0.930 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 9.520 5.490 ;
        RECT 6.505 4.345 6.735 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 9.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.170 ;
        RECT 4.165 0.450 4.395 0.700 ;
        RECT 6.585 0.450 6.815 0.700 ;
        RECT 8.825 0.450 9.055 0.700 ;
        RECT 0.000 -0.450 9.520 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.860 8.815 4.090 ;
        RECT 0.245 3.280 0.475 3.860 ;
        RECT 8.585 3.280 8.815 3.860 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi211_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi211_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi211_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.160 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.504000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 2.150 3.850 2.400 ;
        RECT 5.575 2.170 6.640 2.400 ;
        RECT 3.510 1.985 4.890 2.150 ;
        RECT 5.575 1.985 5.805 2.170 ;
        RECT 3.510 1.755 5.805 1.985 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.504000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.545 2.630 8.725 2.860 ;
        RECT 1.545 2.215 1.775 2.630 ;
        RECT 5.115 2.215 5.345 2.630 ;
        RECT 6.870 2.215 8.725 2.630 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.556000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.860 2.730 19.450 2.960 ;
        RECT 9.860 2.270 10.200 2.730 ;
        RECT 13.505 2.215 13.735 2.730 ;
        RECT 18.960 2.270 19.450 2.730 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.556000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.520 1.985 12.860 2.500 ;
        RECT 14.190 2.270 16.500 2.500 ;
        RECT 14.190 2.150 14.420 2.270 ;
        RECT 13.960 1.985 14.420 2.150 ;
        RECT 12.520 1.755 14.420 1.985 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.682000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.935 3.320 2.165 3.900 ;
        RECT 3.975 3.320 4.205 3.900 ;
        RECT 5.750 3.320 6.245 3.900 ;
        RECT 8.055 3.320 8.285 3.900 ;
        RECT 1.085 3.090 8.285 3.320 ;
        RECT 1.085 1.540 1.315 3.090 ;
        RECT 1.085 1.525 3.040 1.540 ;
        RECT 1.085 1.310 18.670 1.525 ;
        RECT 2.955 1.180 18.670 1.310 ;
        RECT 2.955 0.680 3.185 1.180 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 20.160 5.490 ;
        RECT 11.475 3.650 11.705 4.590 ;
        RECT 16.795 3.650 17.025 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 20.590 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 20.590 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.675 0.450 0.905 1.165 ;
        RECT 4.995 0.450 5.225 0.695 ;
        RECT 9.020 0.450 9.360 0.950 ;
        RECT 11.680 0.450 12.020 0.950 ;
        RECT 14.340 0.450 14.680 0.950 ;
        RECT 17.000 0.450 17.340 0.950 ;
        RECT 19.505 0.450 19.735 1.035 ;
        RECT 0.000 -0.450 20.160 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.915 4.130 9.305 4.360 ;
        RECT 0.915 3.550 1.145 4.130 ;
        RECT 2.955 3.550 3.185 4.130 ;
        RECT 4.995 3.550 5.225 4.130 ;
        RECT 7.035 3.550 7.265 4.130 ;
        RECT 9.075 3.420 9.305 4.130 ;
        RECT 14.135 3.420 14.365 4.360 ;
        RECT 19.455 3.420 19.685 4.360 ;
        RECT 9.075 3.190 19.685 3.420 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi211_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi221_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi221_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.160 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.626000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.145 2.865 6.040 3.270 ;
        RECT 5.145 2.415 5.375 2.865 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.626000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 2.165 4.330 2.710 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.626000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.255 1.210 2.090 2.065 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.626000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 2.255 1.015 2.710 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.360 1.670 3.210 2.230 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.184000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.565 1.590 4.795 3.685 ;
        RECT 4.565 1.440 5.915 1.590 ;
        RECT 2.425 1.210 5.915 1.440 ;
        RECT 2.425 1.075 2.655 1.210 ;
        RECT 5.685 0.680 5.915 1.210 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 6.160 5.490 ;
        RECT 1.365 3.875 1.595 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.590 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.590 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.285 0.450 0.515 1.300 ;
        RECT 3.725 0.450 3.955 0.980 ;
        RECT 0.000 -0.450 6.160 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.545 4.130 5.815 4.360 ;
        RECT 0.345 3.170 0.575 3.750 ;
        RECT 2.385 3.170 2.615 3.685 ;
        RECT 3.545 3.550 3.775 4.130 ;
        RECT 5.585 3.550 5.815 4.130 ;
        RECT 0.345 2.940 2.615 3.170 ;
        RECT 2.385 2.875 2.615 2.940 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi221_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi221_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi221_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.760 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.252000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.225 2.470 10.490 2.700 ;
        RECT 10.165 1.210 10.490 2.470 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.252000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.240 1.590 8.470 2.115 ;
        RECT 7.300 1.210 8.470 1.590 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.252000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.945 1.665 3.845 2.180 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.252000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.890 2.440 5.480 2.670 ;
        RECT 4.490 2.205 5.480 2.440 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.715 2.145 1.010 2.785 ;
        RECT 0.715 1.915 2.715 2.145 ;
        RECT 2.485 1.435 2.715 1.915 ;
        RECT 4.630 1.520 6.370 1.750 ;
        RECT 4.630 1.435 4.890 1.520 ;
        RECT 2.485 1.205 4.890 1.435 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.111250 ;
    PORT
      LAYER Metal1 ;
        RECT 7.720 3.250 7.950 3.830 ;
        RECT 9.760 3.250 11.110 3.830 ;
        RECT 6.765 3.020 11.110 3.250 ;
        RECT 0.245 1.455 2.255 1.685 ;
        RECT 0.245 1.315 0.475 1.455 ;
        RECT 2.025 0.975 2.255 1.455 ;
        RECT 6.765 1.290 6.995 3.020 ;
        RECT 5.120 1.060 6.995 1.290 ;
        RECT 5.120 0.975 5.350 1.060 ;
        RECT 2.025 0.745 5.350 0.975 ;
        RECT 6.765 0.920 6.995 1.060 ;
        RECT 10.880 0.845 11.110 3.020 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 11.760 5.490 ;
        RECT 2.330 4.400 2.670 4.590 ;
        RECT 4.390 4.400 4.730 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 12.190 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.190 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 5.580 0.450 5.810 0.830 ;
        RECT 8.920 0.450 9.150 1.300 ;
        RECT 0.000 -0.450 11.760 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 6.665 4.170 11.065 4.290 ;
        RECT 0.345 4.060 11.065 4.170 ;
        RECT 0.345 3.940 6.895 4.060 ;
        RECT 0.345 3.360 0.575 3.940 ;
        RECT 1.365 3.480 5.695 3.710 ;
        RECT 6.665 3.480 6.895 3.940 ;
        RECT 8.740 3.480 8.970 4.060 ;
        RECT 1.365 2.900 1.595 3.480 ;
        RECT 3.405 2.900 3.635 3.480 ;
        RECT 5.465 2.900 5.695 3.480 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi221_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi221_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi221_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.400 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.504000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.210 2.140 14.550 2.500 ;
        RECT 16.930 2.140 17.270 2.400 ;
        RECT 14.210 1.910 17.270 2.140 ;
        RECT 19.540 2.370 21.450 2.600 ;
        RECT 19.540 1.950 19.770 2.370 ;
        RECT 16.950 1.440 17.270 1.910 ;
        RECT 18.000 1.720 19.770 1.950 ;
        RECT 18.000 1.440 18.230 1.720 ;
        RECT 16.950 1.210 18.230 1.440 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.504000 ;
    PORT
      LAYER Metal1 ;
        RECT 16.470 2.630 17.740 2.860 ;
        RECT 16.470 2.600 16.700 2.630 ;
        RECT 16.150 2.370 16.700 2.600 ;
        RECT 17.510 2.500 17.740 2.630 ;
        RECT 17.510 2.270 19.310 2.500 ;
        RECT 17.510 1.770 17.770 2.270 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.504000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.700 2.085 1.040 2.600 ;
        RECT 3.695 2.085 3.925 2.400 ;
        RECT 0.700 1.985 3.925 2.085 ;
        RECT 6.195 2.370 8.160 2.600 ;
        RECT 6.195 1.985 6.425 2.370 ;
        RECT 0.700 1.855 6.425 1.985 ;
        RECT 3.510 1.755 6.425 1.855 ;
        RECT 3.510 1.210 3.770 1.755 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.504000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 2.630 5.965 2.860 ;
        RECT 1.270 2.315 1.985 2.630 ;
        RECT 5.735 2.215 5.965 2.630 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.556000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.110 2.270 9.650 2.710 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 8.064500 ;
    PORT
      LAYER Metal1 ;
        RECT 14.605 3.320 14.835 3.900 ;
        RECT 16.645 3.320 16.875 3.900 ;
        RECT 18.685 3.320 18.915 3.900 ;
        RECT 20.725 3.320 20.955 3.900 ;
        RECT 13.590 3.090 20.955 3.320 ;
        RECT 0.245 1.395 3.280 1.625 ;
        RECT 13.590 1.480 13.850 3.090 ;
        RECT 0.245 0.680 0.475 1.395 ;
        RECT 3.050 0.965 3.280 1.395 ;
        RECT 4.430 1.250 16.720 1.480 ;
        RECT 4.430 0.965 4.660 1.250 ;
        RECT 3.050 0.735 4.660 0.965 ;
        RECT 8.555 0.680 8.785 1.250 ;
        RECT 11.165 0.680 11.395 1.250 ;
        RECT 13.405 0.680 13.635 1.250 ;
        RECT 16.490 0.965 16.720 1.250 ;
        RECT 18.460 1.260 21.975 1.490 ;
        RECT 18.460 0.965 18.690 1.260 ;
        RECT 16.490 0.735 18.690 0.965 ;
        RECT 21.745 0.680 21.975 1.260 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 22.400 5.490 ;
        RECT 0.295 3.090 0.525 4.590 ;
        RECT 2.335 3.550 2.565 4.590 ;
        RECT 4.375 3.550 4.605 4.590 ;
        RECT 6.415 3.550 6.645 4.590 ;
        RECT 8.455 3.550 8.685 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 22.830 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 22.830 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.335 0.450 2.565 1.165 ;
        RECT 6.415 0.450 6.645 1.020 ;
        RECT 10.045 0.450 10.275 1.020 ;
        RECT 12.285 0.450 12.515 1.020 ;
        RECT 15.625 0.450 15.855 1.020 ;
        RECT 19.705 0.450 19.935 1.020 ;
        RECT 0.000 -0.450 22.400 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 9.175 4.130 21.975 4.360 ;
        RECT 1.315 3.320 1.545 3.900 ;
        RECT 3.355 3.320 3.585 3.900 ;
        RECT 5.395 3.320 5.625 3.900 ;
        RECT 7.435 3.320 7.665 3.900 ;
        RECT 9.175 3.550 9.405 4.130 ;
        RECT 10.195 3.320 10.425 3.900 ;
        RECT 11.215 3.535 11.445 4.130 ;
        RECT 1.315 3.305 10.425 3.320 ;
        RECT 12.235 3.305 12.465 3.900 ;
        RECT 13.305 3.545 13.535 4.130 ;
        RECT 15.625 3.550 15.855 4.130 ;
        RECT 17.665 3.550 17.895 4.130 ;
        RECT 19.705 3.550 19.935 4.130 ;
        RECT 1.315 3.090 12.465 3.305 ;
        RECT 21.745 3.090 21.975 4.130 ;
        RECT 10.340 3.075 12.465 3.090 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi221_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi222_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi222_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.800 2.415 7.725 3.270 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.145 1.770 6.010 2.150 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.670 1.770 3.830 2.150 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.050 2.255 4.910 2.710 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.220 1.210 2.145 2.060 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.115 2.235 1.070 2.710 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.169200 ;
    PORT
      LAYER Metal1 ;
        RECT 6.220 2.875 6.470 3.215 ;
        RECT 6.240 1.590 6.470 2.875 ;
        RECT 6.240 1.490 7.470 1.590 ;
        RECT 3.160 1.210 7.470 1.490 ;
        RECT 3.160 0.680 3.390 1.210 ;
        RECT 7.240 0.680 7.470 1.210 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.840 5.490 ;
        RECT 0.400 3.875 0.630 4.590 ;
        RECT 2.440 3.875 2.670 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 8.270 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.270 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.480 0.450 0.710 1.165 ;
        RECT 5.200 0.450 5.430 0.695 ;
        RECT 0.000 -0.450 7.840 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.160 4.130 7.470 4.360 ;
        RECT 1.365 3.170 1.710 3.700 ;
        RECT 3.160 3.550 3.390 4.130 ;
        RECT 4.125 3.170 4.465 3.810 ;
        RECT 5.200 3.550 7.470 4.130 ;
        RECT 1.365 2.940 4.465 3.170 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi222_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi222_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi222_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.000 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.700 2.345 12.960 2.575 ;
        RECT 11.775 1.210 12.960 2.345 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.945 1.210 11.050 2.115 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.605 2.380 8.810 2.610 ;
        RECT 7.605 1.770 8.810 2.380 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.255 1.770 6.770 2.150 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.115 2.645 0.970 3.270 ;
        RECT 0.115 2.415 4.065 2.645 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.825 1.770 2.090 2.150 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 5.275800 ;
    PORT
      LAYER Metal1 ;
        RECT 10.195 3.105 10.425 3.685 ;
        RECT 12.235 3.105 12.465 3.685 ;
        RECT 9.040 2.875 13.485 3.105 ;
        RECT 9.040 1.490 9.470 2.875 ;
        RECT 0.280 0.925 9.470 1.490 ;
        RECT 0.280 0.680 0.510 0.925 ;
        RECT 4.980 0.680 5.210 0.925 ;
        RECT 9.160 0.845 9.470 0.925 ;
        RECT 13.255 0.845 13.485 2.875 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 14.000 5.490 ;
        RECT 0.280 3.875 0.510 4.590 ;
        RECT 2.320 3.875 2.550 4.590 ;
        RECT 4.360 3.875 4.590 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 14.430 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.430 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.320 0.450 2.550 0.695 ;
        RECT 7.120 0.450 7.350 0.695 ;
        RECT 11.215 0.450 11.445 0.695 ;
        RECT 0.000 -0.450 14.000 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 5.080 3.915 13.485 4.145 ;
        RECT 1.300 3.105 1.530 3.685 ;
        RECT 3.340 3.105 3.570 3.685 ;
        RECT 5.080 3.335 5.310 3.915 ;
        RECT 6.100 3.105 6.330 3.685 ;
        RECT 7.120 3.335 7.350 3.915 ;
        RECT 8.140 3.105 8.370 3.685 ;
        RECT 9.160 3.335 9.390 3.915 ;
        RECT 11.215 3.335 11.445 3.915 ;
        RECT 13.255 3.335 13.485 3.915 ;
        RECT 1.300 2.875 8.370 3.105 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi222_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi222_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi222_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.320 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 17.865 2.150 18.095 2.555 ;
        RECT 17.865 1.985 19.450 2.150 ;
        RECT 20.785 1.985 21.015 2.400 ;
        RECT 24.865 1.985 25.095 2.555 ;
        RECT 17.865 1.755 25.095 1.985 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 20.135 2.770 22.780 2.860 ;
        RECT 19.750 2.630 23.055 2.770 ;
        RECT 19.750 2.270 20.320 2.630 ;
        RECT 22.595 2.215 23.055 2.630 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.670 1.600 9.930 2.555 ;
        RECT 12.625 1.655 12.855 2.400 ;
        RECT 16.605 1.655 16.835 2.555 ;
        RECT 12.625 1.600 16.835 1.655 ;
        RECT 9.670 1.425 16.835 1.600 ;
        RECT 9.670 1.370 12.775 1.425 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.100 2.770 14.140 2.860 ;
        RECT 12.100 2.630 14.895 2.770 ;
        RECT 12.100 2.500 12.330 2.630 ;
        RECT 13.955 2.540 14.895 2.630 ;
        RECT 11.690 1.830 12.330 2.500 ;
        RECT 14.665 2.215 14.895 2.540 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.825 1.985 1.055 2.555 ;
        RECT 3.745 1.985 3.975 2.555 ;
        RECT 7.825 2.150 8.055 2.555 ;
        RECT 6.310 1.985 8.055 2.150 ;
        RECT 0.825 1.755 8.055 1.985 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.285 2.855 5.710 3.015 ;
        RECT 3.285 2.785 6.015 2.855 ;
        RECT 1.830 2.445 2.090 2.710 ;
        RECT 3.285 2.445 3.515 2.785 ;
        RECT 5.490 2.625 6.015 2.785 ;
        RECT 1.830 2.215 3.515 2.445 ;
        RECT 5.785 2.215 6.015 2.625 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 9.284400 ;
    PORT
      LAYER Metal1 ;
        RECT 18.305 3.230 18.535 3.900 ;
        RECT 20.345 3.320 20.575 3.900 ;
        RECT 22.385 3.320 22.615 3.900 ;
        RECT 19.740 3.230 23.220 3.320 ;
        RECT 24.425 3.230 24.655 3.900 ;
        RECT 17.665 3.090 24.655 3.230 ;
        RECT 17.665 3.015 19.925 3.090 ;
        RECT 17.285 3.000 19.925 3.015 ;
        RECT 23.035 3.000 24.655 3.090 ;
        RECT 17.285 2.785 17.895 3.000 ;
        RECT 17.285 1.195 17.515 2.785 ;
        RECT 0.190 1.140 8.690 1.195 ;
        RECT 17.285 1.155 25.730 1.195 ;
        RECT 13.405 1.140 25.730 1.155 ;
        RECT 0.190 0.925 25.730 1.140 ;
        RECT 0.190 0.910 13.490 0.925 ;
        RECT 24.730 0.710 25.730 0.925 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 26.320 5.490 ;
        RECT 0.245 3.245 0.475 4.590 ;
        RECT 2.285 3.705 2.515 4.590 ;
        RECT 4.325 3.705 4.555 4.590 ;
        RECT 6.365 3.560 6.595 4.590 ;
        RECT 8.405 3.545 8.635 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 26.750 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 26.750 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.230 0.450 2.570 0.680 ;
        RECT 6.310 0.450 6.650 0.680 ;
        RECT 11.110 0.450 11.450 0.680 ;
        RECT 15.245 0.450 15.475 0.695 ;
        RECT 19.325 0.450 19.555 0.695 ;
        RECT 23.405 0.450 23.635 0.695 ;
        RECT 0.000 -0.450 26.320 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 9.125 4.130 25.675 4.360 ;
        RECT 1.265 3.475 1.495 4.055 ;
        RECT 3.305 3.475 3.535 4.055 ;
        RECT 5.345 3.475 5.575 4.055 ;
        RECT 1.265 3.315 6.150 3.475 ;
        RECT 7.385 3.315 7.615 4.055 ;
        RECT 9.125 3.545 9.355 4.130 ;
        RECT 10.145 3.320 10.375 3.900 ;
        RECT 11.165 3.550 11.395 4.130 ;
        RECT 12.185 3.320 12.415 3.900 ;
        RECT 13.205 3.550 13.435 4.130 ;
        RECT 14.225 3.320 14.510 3.900 ;
        RECT 15.245 3.460 15.475 4.130 ;
        RECT 9.405 3.315 14.510 3.320 ;
        RECT 1.265 3.245 14.510 3.315 ;
        RECT 5.930 3.230 14.510 3.245 ;
        RECT 16.265 3.230 16.495 3.900 ;
        RECT 17.285 3.405 17.515 4.130 ;
        RECT 19.325 3.460 19.555 4.130 ;
        RECT 21.365 3.550 21.595 4.130 ;
        RECT 23.405 3.460 23.635 4.130 ;
        RECT 25.445 3.245 25.675 4.130 ;
        RECT 5.930 3.090 16.495 3.230 ;
        RECT 5.930 3.085 9.455 3.090 ;
        RECT 14.325 3.000 16.495 3.090 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi222_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__buf_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__buf_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.853500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 1.015 2.710 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.390 2.890 2.895 3.775 ;
        RECT 2.665 1.590 2.895 2.890 ;
        RECT 2.390 0.740 2.895 1.590 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 3.360 5.490 ;
        RECT 1.365 3.400 1.595 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 3.790 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 3.790 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.080 ;
        RECT 0.000 -0.450 3.360 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 3.170 0.575 3.775 ;
        RECT 0.345 2.940 2.160 3.170 ;
        RECT 1.930 2.585 2.160 2.940 ;
        RECT 1.930 1.775 2.215 2.585 ;
        RECT 1.930 1.540 2.160 1.775 ;
        RECT 0.245 1.310 2.160 1.540 ;
        RECT 0.245 0.740 0.475 1.310 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__buf_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__buf_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__buf_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.330 0.970 2.710 ;
        RECT 0.630 2.000 0.970 2.330 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.821000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.485 3.015 2.715 4.360 ;
        RECT 2.485 2.730 3.280 3.015 ;
        RECT 2.980 1.590 3.280 2.730 ;
        RECT 2.330 1.210 3.280 1.590 ;
        RECT 2.330 0.710 2.715 1.210 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 4.480 5.490 ;
        RECT 1.265 3.550 1.495 4.590 ;
        RECT 3.505 3.550 3.735 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 4.910 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.165 ;
        RECT 3.605 0.450 3.835 1.520 ;
        RECT 0.000 -0.450 4.480 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.320 0.475 4.360 ;
        RECT 0.245 3.090 1.430 3.320 ;
        RECT 1.200 2.500 1.430 3.090 ;
        RECT 1.200 2.270 2.750 2.500 ;
        RECT 1.200 1.625 1.430 2.270 ;
        RECT 0.245 1.395 1.430 1.625 ;
        RECT 0.245 0.710 0.475 1.395 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__buf_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__buf_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__buf_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.585 0.410 2.710 ;
        RECT 0.150 1.770 0.915 2.585 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.207000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.675 3.105 2.905 4.360 ;
        RECT 4.815 3.105 5.045 3.685 ;
        RECT 2.675 2.875 5.045 3.105 ;
        RECT 3.510 2.000 4.005 2.875 ;
        RECT 2.675 1.770 5.145 2.000 ;
        RECT 2.675 0.730 2.905 1.770 ;
        RECT 4.915 0.730 5.145 1.770 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.600 5.490 ;
        RECT 1.265 3.550 1.495 4.590 ;
        RECT 3.695 3.550 3.925 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.555 0.450 1.785 1.165 ;
        RECT 3.795 0.450 4.025 1.540 ;
        RECT 0.000 -0.450 5.600 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.320 0.475 4.360 ;
        RECT 0.245 3.090 1.375 3.320 ;
        RECT 1.145 2.500 1.375 3.090 ;
        RECT 1.145 2.270 3.220 2.500 ;
        RECT 1.145 1.540 1.375 2.270 ;
        RECT 0.245 1.310 1.375 1.540 ;
        RECT 0.245 0.730 0.475 1.310 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__buf_3

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__buf_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__buf_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 2.270 1.910 2.650 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.642000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.605 3.320 3.835 4.360 ;
        RECT 5.745 3.320 6.075 4.360 ;
        RECT 3.605 3.090 6.075 3.320 ;
        RECT 5.575 1.950 6.075 3.090 ;
        RECT 3.605 1.720 6.075 1.950 ;
        RECT 3.605 0.680 3.865 1.720 ;
        RECT 5.845 0.680 6.075 1.720 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.840 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 8.270 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.270 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 4.725 0.450 4.955 1.490 ;
        RECT 6.965 0.450 7.195 1.490 ;
        RECT 0.000 -0.450 7.840 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 1.365 3.090 2.370 3.320 ;
        RECT 2.140 2.500 2.370 3.090 ;
        RECT 2.140 2.270 4.620 2.500 ;
        RECT 2.140 1.920 2.370 2.270 ;
        RECT 1.365 1.690 2.370 1.920 ;
        RECT 1.365 0.680 1.595 1.690 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__buf_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__buf_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__buf_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.560 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.685 2.215 4.205 2.650 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 7.284000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.845 3.320 6.075 4.360 ;
        RECT 7.985 3.320 8.215 4.360 ;
        RECT 10.225 3.320 10.455 4.360 ;
        RECT 12.465 3.320 12.695 4.360 ;
        RECT 5.845 2.880 12.695 3.320 ;
        RECT 8.970 2.040 9.470 2.880 ;
        RECT 5.845 1.985 9.470 2.040 ;
        RECT 5.845 1.720 12.795 1.985 ;
        RECT 5.845 0.680 6.075 1.720 ;
        RECT 8.055 0.680 8.315 1.720 ;
        RECT 10.325 0.680 10.555 1.720 ;
        RECT 12.565 0.680 12.795 1.720 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 14.560 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
        RECT 9.105 3.550 9.335 4.590 ;
        RECT 11.345 3.550 11.575 4.590 ;
        RECT 13.585 3.550 13.815 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 14.990 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.990 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 4.725 0.450 4.955 1.490 ;
        RECT 6.965 0.450 7.195 1.490 ;
        RECT 9.205 0.450 9.435 1.165 ;
        RECT 11.445 0.450 11.675 1.490 ;
        RECT 13.685 0.450 13.915 1.490 ;
        RECT 0.000 -0.450 14.560 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 3.205 1.595 4.360 ;
        RECT 3.505 3.205 3.735 4.360 ;
        RECT 1.365 2.975 4.665 3.205 ;
        RECT 4.435 2.650 4.665 2.975 ;
        RECT 4.435 2.270 8.740 2.650 ;
        RECT 4.435 1.985 4.665 2.270 ;
        RECT 9.700 2.215 13.220 2.650 ;
        RECT 1.365 1.755 4.665 1.985 ;
        RECT 1.365 0.680 1.595 1.755 ;
        RECT 3.605 0.680 3.835 1.755 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__buf_8

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__buf_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__buf_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 10.242000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.130 2.270 5.640 2.650 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 10.926000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.135 3.320 8.365 4.360 ;
        RECT 10.275 3.320 10.505 4.360 ;
        RECT 12.515 3.320 12.745 4.360 ;
        RECT 14.755 3.320 14.985 4.360 ;
        RECT 16.995 3.320 17.225 4.360 ;
        RECT 19.235 3.320 19.465 4.360 ;
        RECT 8.135 2.840 19.465 3.320 ;
        RECT 13.500 2.040 14.000 2.840 ;
        RECT 8.135 1.985 14.000 2.040 ;
        RECT 8.135 1.755 19.565 1.985 ;
        RECT 8.135 0.680 8.365 1.755 ;
        RECT 10.375 0.680 10.605 1.755 ;
        RECT 12.385 0.680 12.845 1.755 ;
        RECT 14.855 0.680 15.085 1.755 ;
        RECT 17.095 0.680 17.325 1.755 ;
        RECT 19.335 0.680 19.565 1.755 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 21.280 5.490 ;
        RECT 0.295 3.550 0.525 4.590 ;
        RECT 2.435 3.550 2.665 4.590 ;
        RECT 4.675 3.550 4.905 4.590 ;
        RECT 6.915 3.550 7.145 4.590 ;
        RECT 9.155 3.875 9.385 4.590 ;
        RECT 11.395 3.550 11.625 4.590 ;
        RECT 13.635 3.550 13.865 4.590 ;
        RECT 15.875 3.550 16.105 4.590 ;
        RECT 18.115 3.550 18.345 4.590 ;
        RECT 20.355 3.550 20.585 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 21.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 21.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.295 0.450 0.525 1.490 ;
        RECT 2.535 0.450 2.765 1.490 ;
        RECT 4.775 0.450 5.005 1.490 ;
        RECT 7.015 0.450 7.245 1.490 ;
        RECT 9.255 0.450 9.485 1.490 ;
        RECT 11.495 0.450 11.725 1.490 ;
        RECT 13.735 0.450 13.965 1.490 ;
        RECT 15.975 0.450 16.205 1.490 ;
        RECT 18.215 0.450 18.445 1.490 ;
        RECT 20.455 0.450 20.685 1.490 ;
        RECT 0.000 -0.450 21.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.415 3.320 1.645 4.360 ;
        RECT 3.555 3.320 3.785 4.360 ;
        RECT 5.820 3.320 6.225 4.360 ;
        RECT 1.415 2.880 6.225 3.320 ;
        RECT 5.895 2.500 6.225 2.880 ;
        RECT 5.895 2.270 12.910 2.500 ;
        RECT 5.895 2.040 6.225 2.270 ;
        RECT 14.230 2.215 19.630 2.555 ;
        RECT 1.415 1.720 6.225 2.040 ;
        RECT 1.415 0.680 1.645 1.720 ;
        RECT 3.655 0.680 3.885 1.720 ;
        RECT 5.895 0.680 6.225 1.720 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__buf_12

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__buf_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__buf_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.000 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 13.655999 ;
    PORT
      LAYER Metal1 ;
        RECT 0.440 2.270 7.830 2.650 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 14.568000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.325 3.320 10.555 4.360 ;
        RECT 12.465 3.320 12.695 4.360 ;
        RECT 14.705 3.320 14.935 4.360 ;
        RECT 16.945 3.320 17.175 4.360 ;
        RECT 19.185 3.320 19.415 4.360 ;
        RECT 21.425 3.320 21.655 4.360 ;
        RECT 23.665 3.320 23.895 4.360 ;
        RECT 25.905 3.320 26.135 4.360 ;
        RECT 10.325 2.960 26.135 3.320 ;
        RECT 17.805 2.040 18.555 2.960 ;
        RECT 10.325 1.985 18.555 2.040 ;
        RECT 10.325 1.720 26.235 1.985 ;
        RECT 10.325 0.680 10.555 1.720 ;
        RECT 12.565 0.680 12.795 1.720 ;
        RECT 14.805 0.680 15.035 1.720 ;
        RECT 17.045 0.680 17.305 1.720 ;
        RECT 19.285 0.680 19.515 1.720 ;
        RECT 21.525 0.680 21.755 1.720 ;
        RECT 23.765 0.680 23.995 1.720 ;
        RECT 26.005 0.680 26.235 1.720 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 28.000 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
        RECT 9.105 3.550 9.335 4.590 ;
        RECT 11.345 3.550 11.575 4.590 ;
        RECT 13.585 3.550 13.815 4.590 ;
        RECT 15.825 3.550 16.055 4.590 ;
        RECT 18.065 3.550 18.295 4.590 ;
        RECT 20.305 3.550 20.535 4.590 ;
        RECT 22.545 3.550 22.775 4.590 ;
        RECT 24.785 3.550 25.015 4.590 ;
        RECT 27.025 3.550 27.255 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 28.430 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 28.430 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 4.725 0.450 4.955 1.490 ;
        RECT 6.965 0.450 7.195 1.490 ;
        RECT 9.205 0.450 9.435 1.490 ;
        RECT 11.445 0.450 11.675 1.490 ;
        RECT 13.685 0.450 13.915 1.490 ;
        RECT 15.925 0.450 16.155 1.490 ;
        RECT 18.165 0.450 18.395 1.490 ;
        RECT 20.405 0.450 20.635 1.490 ;
        RECT 22.645 0.450 22.875 1.490 ;
        RECT 24.885 0.450 25.115 1.490 ;
        RECT 27.125 0.450 27.355 1.490 ;
        RECT 0.000 -0.450 28.000 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.505 3.320 3.735 4.360 ;
        RECT 5.745 3.320 5.975 4.360 ;
        RECT 8.060 3.320 8.425 4.360 ;
        RECT 1.365 2.880 8.425 3.320 ;
        RECT 8.060 2.630 8.425 2.880 ;
        RECT 8.060 2.270 16.980 2.630 ;
        RECT 8.060 2.040 8.425 2.270 ;
        RECT 18.785 2.215 26.065 2.555 ;
        RECT 1.365 1.720 8.425 2.040 ;
        RECT 1.365 0.680 1.595 1.720 ;
        RECT 3.605 0.680 3.835 1.720 ;
        RECT 5.845 0.680 6.075 1.720 ;
        RECT 8.085 0.680 8.425 1.720 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__buf_16

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__buf_20
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__buf_20 ;
  ORIGIN 0.000 0.000 ;
  SIZE 34.720 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 17.070000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.685 2.215 9.845 2.650 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 18.209999 ;
    PORT
      LAYER Metal1 ;
        RECT 12.565 3.320 12.795 4.360 ;
        RECT 14.705 3.320 14.935 4.360 ;
        RECT 16.945 3.320 17.175 4.360 ;
        RECT 19.185 3.320 19.415 4.360 ;
        RECT 21.425 3.320 21.655 4.360 ;
        RECT 23.665 3.320 23.895 4.360 ;
        RECT 25.905 3.320 26.135 4.360 ;
        RECT 28.145 3.320 28.375 4.360 ;
        RECT 30.385 3.320 30.615 4.360 ;
        RECT 32.625 3.320 32.855 4.360 ;
        RECT 12.565 2.885 32.855 3.320 ;
        RECT 22.285 2.880 32.855 2.885 ;
        RECT 22.285 2.030 23.035 2.880 ;
        RECT 12.565 1.980 23.035 2.030 ;
        RECT 12.565 1.720 32.955 1.980 ;
        RECT 12.565 0.680 12.825 1.720 ;
        RECT 14.805 0.680 15.035 1.720 ;
        RECT 17.045 0.680 17.275 1.720 ;
        RECT 19.285 0.680 19.515 1.720 ;
        RECT 21.525 0.680 21.755 1.720 ;
        RECT 23.765 0.680 23.995 1.720 ;
        RECT 26.005 0.680 26.235 1.720 ;
        RECT 28.245 0.680 28.475 1.720 ;
        RECT 30.485 0.680 30.715 1.720 ;
        RECT 32.725 0.680 32.955 1.720 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 34.720 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
        RECT 9.105 3.550 9.335 4.590 ;
        RECT 11.345 3.875 11.575 4.590 ;
        RECT 13.585 3.550 13.815 4.590 ;
        RECT 15.825 3.550 16.055 4.590 ;
        RECT 18.065 3.550 18.295 4.590 ;
        RECT 20.305 3.550 20.535 4.590 ;
        RECT 22.545 3.550 22.775 4.590 ;
        RECT 24.785 3.550 25.015 4.590 ;
        RECT 27.025 3.550 27.255 4.590 ;
        RECT 29.265 3.550 29.495 4.590 ;
        RECT 31.505 3.550 31.735 4.590 ;
        RECT 33.745 3.550 33.975 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 35.150 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 35.150 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 4.725 0.450 4.955 1.490 ;
        RECT 6.965 0.450 7.195 1.490 ;
        RECT 9.205 0.450 9.435 1.490 ;
        RECT 11.445 0.450 11.675 1.490 ;
        RECT 13.685 0.450 13.915 1.490 ;
        RECT 15.925 0.450 16.155 1.490 ;
        RECT 18.165 0.450 18.395 1.490 ;
        RECT 20.405 0.450 20.635 1.490 ;
        RECT 22.645 0.450 22.875 1.490 ;
        RECT 24.885 0.450 25.115 1.490 ;
        RECT 27.125 0.450 27.355 1.490 ;
        RECT 29.365 0.450 29.595 1.490 ;
        RECT 31.605 0.450 31.835 1.490 ;
        RECT 33.845 0.450 34.075 1.490 ;
        RECT 0.000 -0.450 34.720 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.505 3.320 3.735 4.360 ;
        RECT 5.745 3.320 5.975 4.360 ;
        RECT 7.985 3.320 8.215 4.360 ;
        RECT 10.225 3.320 10.555 4.360 ;
        RECT 1.365 2.900 10.555 3.320 ;
        RECT 10.225 2.650 10.555 2.900 ;
        RECT 10.225 2.270 21.100 2.650 ;
        RECT 10.225 1.975 10.555 2.270 ;
        RECT 23.265 2.215 32.425 2.650 ;
        RECT 1.365 1.720 10.555 1.975 ;
        RECT 1.365 0.680 1.595 1.720 ;
        RECT 3.605 0.680 3.835 1.720 ;
        RECT 5.845 0.680 6.075 1.720 ;
        RECT 8.085 0.680 8.315 1.720 ;
        RECT 10.325 0.680 10.555 1.720 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__buf_20

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__bufz_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__bufz_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.698000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.870 2.330 2.090 2.710 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.849000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.630 1.745 4.990 2.150 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.640 1.650 6.870 3.685 ;
        RECT 6.640 0.840 7.130 1.650 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.280 5.490 ;
        RECT 1.365 3.635 1.595 4.590 ;
        RECT 5.440 3.875 5.670 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 7.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.425 ;
        RECT 5.660 0.450 5.890 0.690 ;
        RECT 0.000 -0.450 7.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.060 0.575 4.285 ;
        RECT 2.385 4.055 4.650 4.285 ;
        RECT 2.385 3.475 2.615 4.055 ;
        RECT 2.630 2.815 2.895 3.155 ;
        RECT 2.630 2.060 2.860 2.815 ;
        RECT 3.405 2.060 3.635 3.815 ;
        RECT 0.245 1.830 2.860 2.060 ;
        RECT 3.090 1.830 3.635 2.060 ;
        RECT 4.170 2.700 4.650 4.055 ;
        RECT 4.170 2.470 6.345 2.700 ;
        RECT 0.245 1.315 0.475 1.830 ;
        RECT 2.485 0.950 2.715 1.425 ;
        RECT 3.090 1.115 3.320 1.830 ;
        RECT 4.170 1.600 4.400 2.470 ;
        RECT 3.550 1.370 4.400 1.600 ;
        RECT 5.305 1.115 6.385 2.055 ;
        RECT 3.090 0.950 6.385 1.115 ;
        RECT 2.485 0.920 6.385 0.950 ;
        RECT 2.485 0.720 5.430 0.920 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__bufz_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__bufz_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__bufz_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.400 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.880 2.330 2.090 2.715 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.692000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.125 2.285 5.465 2.710 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.622400 ;
    PORT
      LAYER Metal1 ;
        RECT 6.705 0.840 7.130 3.720 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 8.400 5.490 ;
        RECT 1.375 3.845 1.605 4.590 ;
        RECT 5.685 3.880 5.915 4.590 ;
        RECT 7.725 3.880 7.955 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 8.830 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.830 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.375 0.450 1.605 1.165 ;
        RECT 5.685 0.450 5.915 1.160 ;
        RECT 7.925 0.450 8.155 1.160 ;
        RECT 0.000 -0.450 8.400 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.255 2.060 0.585 3.685 ;
        RECT 2.925 3.505 4.890 3.685 ;
        RECT 2.925 3.455 6.355 3.505 ;
        RECT 2.925 2.875 3.155 3.455 ;
        RECT 4.665 3.275 6.355 3.455 ;
        RECT 2.320 2.415 3.715 2.645 ;
        RECT 2.320 2.060 2.550 2.415 ;
        RECT 3.945 2.185 4.175 3.215 ;
        RECT 0.255 1.830 2.550 2.060 ;
        RECT 3.155 1.955 4.175 2.185 ;
        RECT 0.255 0.845 0.485 1.830 ;
        RECT 3.155 1.490 3.385 1.955 ;
        RECT 4.665 1.655 4.895 3.275 ;
        RECT 6.125 2.450 6.355 3.275 ;
        RECT 2.495 1.085 3.385 1.490 ;
        RECT 3.615 1.315 4.895 1.655 ;
        RECT 5.125 1.825 6.410 2.055 ;
        RECT 5.125 1.085 5.355 1.825 ;
        RECT 2.495 0.680 5.355 1.085 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__bufz_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__bufz_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__bufz_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.640 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.870 2.330 2.090 2.710 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.547000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 1.750 6.115 2.150 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.995200 ;
    PORT
      LAYER Metal1 ;
        RECT 7.895 3.140 8.125 3.720 ;
        RECT 9.935 3.140 10.165 3.720 ;
        RECT 7.895 2.910 10.165 3.140 ;
        RECT 9.045 1.650 9.390 2.910 ;
        RECT 7.865 1.390 10.335 1.650 ;
        RECT 7.865 0.840 8.095 1.390 ;
        RECT 10.105 0.840 10.335 1.390 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 10.640 5.490 ;
        RECT 1.365 3.845 1.595 4.590 ;
        RECT 4.655 4.035 4.885 4.590 ;
        RECT 6.695 3.565 6.925 4.590 ;
        RECT 8.915 3.880 9.145 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 11.070 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 11.070 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.165 ;
        RECT 4.270 0.450 4.610 0.680 ;
        RECT 6.510 0.450 6.850 0.680 ;
        RECT 8.985 0.450 9.215 1.160 ;
        RECT 0.000 -0.450 10.640 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.060 0.575 3.685 ;
        RECT 2.915 3.510 5.905 3.740 ;
        RECT 2.915 2.930 3.145 3.510 ;
        RECT 2.320 2.470 3.650 2.700 ;
        RECT 2.320 2.060 2.550 2.470 ;
        RECT 3.935 2.060 4.165 3.215 ;
        RECT 5.675 2.695 5.905 3.510 ;
        RECT 0.245 1.830 2.550 2.060 ;
        RECT 3.090 1.830 4.165 2.060 ;
        RECT 5.290 2.465 7.665 2.695 ;
        RECT 0.245 0.845 0.475 1.830 ;
        RECT 3.090 1.490 3.320 1.830 ;
        RECT 5.290 1.600 5.520 2.465 ;
        RECT 2.485 1.140 3.320 1.490 ;
        RECT 3.550 1.370 5.520 1.600 ;
        RECT 6.345 1.825 7.665 2.055 ;
        RECT 6.345 1.140 6.575 1.825 ;
        RECT 2.485 0.910 6.575 1.140 ;
        RECT 2.485 0.680 2.715 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__bufz_3

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__bufz_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__bufz_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.760 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.870 2.330 2.090 2.710 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.735 1.770 6.115 2.150 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.244800 ;
    PORT
      LAYER Metal1 ;
        RECT 7.785 3.200 8.015 3.780 ;
        RECT 9.825 3.200 10.055 3.780 ;
        RECT 7.785 2.970 10.055 3.200 ;
        RECT 8.960 1.620 9.420 2.970 ;
        RECT 7.685 1.390 10.155 1.620 ;
        RECT 7.685 0.680 7.915 1.390 ;
        RECT 9.925 0.680 10.155 1.390 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 11.760 5.490 ;
        RECT 1.365 3.845 1.595 4.590 ;
        RECT 4.725 4.350 4.955 4.590 ;
        RECT 6.765 3.880 6.995 4.590 ;
        RECT 8.805 3.880 9.035 4.590 ;
        RECT 10.845 3.880 11.075 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 12.190 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.190 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.165 ;
        RECT 4.270 0.450 4.610 0.635 ;
        RECT 6.510 0.450 6.850 0.635 ;
        RECT 8.805 0.450 9.035 1.160 ;
        RECT 11.045 0.450 11.275 1.160 ;
        RECT 0.000 -0.450 11.760 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.060 0.575 3.685 ;
        RECT 2.915 3.510 4.625 3.740 ;
        RECT 2.915 2.930 3.145 3.510 ;
        RECT 2.320 2.470 3.650 2.700 ;
        RECT 2.320 2.060 2.550 2.470 ;
        RECT 3.935 2.060 4.165 3.215 ;
        RECT 0.245 1.830 2.550 2.060 ;
        RECT 3.090 1.830 4.165 2.060 ;
        RECT 4.395 2.735 4.625 3.510 ;
        RECT 5.745 2.735 5.975 3.720 ;
        RECT 4.395 2.505 8.560 2.735 ;
        RECT 0.245 0.845 0.475 1.830 ;
        RECT 3.090 1.490 3.320 1.830 ;
        RECT 4.395 1.600 4.625 2.505 ;
        RECT 2.485 1.140 3.320 1.490 ;
        RECT 3.550 1.370 4.625 1.600 ;
        RECT 6.345 1.850 8.560 2.080 ;
        RECT 6.345 1.140 6.575 1.850 ;
        RECT 2.485 0.910 6.575 1.140 ;
        RECT 2.485 0.680 2.715 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__bufz_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__bufz_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__bufz_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.480 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.150 1.530 2.710 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.768000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.175 1.770 8.810 2.150 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.489600 ;
    PORT
      LAYER Metal1 ;
        RECT 10.015 3.080 16.365 3.835 ;
        RECT 15.760 1.650 16.365 3.080 ;
        RECT 15.760 1.595 17.065 1.650 ;
        RECT 10.115 0.865 17.065 1.595 ;
        RECT 16.835 0.840 17.065 0.865 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 18.480 5.490 ;
        RECT 1.265 3.845 1.495 4.590 ;
        RECT 4.915 3.880 5.145 4.590 ;
        RECT 6.955 3.880 7.185 4.590 ;
        RECT 8.995 3.880 9.225 4.590 ;
        RECT 11.035 4.350 11.265 4.590 ;
        RECT 13.075 4.350 13.305 4.590 ;
        RECT 15.115 4.350 15.345 4.590 ;
        RECT 17.155 3.880 17.385 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 18.910 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 18.910 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 0.695 ;
        RECT 4.270 0.450 4.610 0.625 ;
        RECT 6.755 0.450 6.985 0.690 ;
        RECT 8.995 0.450 9.225 0.690 ;
        RECT 11.180 0.450 11.520 0.635 ;
        RECT 13.420 0.450 13.760 0.635 ;
        RECT 15.660 0.450 16.000 0.635 ;
        RECT 17.955 0.450 18.185 1.160 ;
        RECT 0.000 -0.450 18.480 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 2.925 3.915 4.635 4.145 ;
        RECT 0.245 1.545 0.475 3.685 ;
        RECT 2.925 3.335 3.155 3.915 ;
        RECT 1.805 2.470 3.650 2.700 ;
        RECT 1.805 1.545 2.035 2.470 ;
        RECT 3.945 2.240 4.175 3.685 ;
        RECT 0.245 1.315 2.035 1.545 ;
        RECT 3.145 2.010 4.175 2.240 ;
        RECT 4.405 3.250 4.635 3.915 ;
        RECT 7.975 3.250 8.205 3.830 ;
        RECT 4.405 3.140 8.205 3.250 ;
        RECT 4.405 2.910 9.665 3.140 ;
        RECT 3.145 1.490 3.375 2.010 ;
        RECT 4.405 1.780 4.635 2.910 ;
        RECT 9.435 2.750 9.665 2.910 ;
        RECT 9.435 2.410 14.895 2.750 ;
        RECT 2.485 1.085 3.375 1.490 ;
        RECT 3.605 1.550 4.635 1.780 ;
        RECT 9.435 1.825 14.325 2.150 ;
        RECT 3.605 1.315 3.835 1.550 ;
        RECT 9.435 1.490 9.665 1.825 ;
        RECT 5.635 1.260 9.665 1.490 ;
        RECT 5.635 1.085 5.865 1.260 ;
        RECT 2.485 0.855 5.865 1.085 ;
        RECT 2.485 0.680 2.715 0.855 ;
        RECT 7.875 0.680 8.105 1.260 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__bufz_8

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__bufz_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__bufz_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.200 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.330 1.575 2.710 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 10.151999 ;
    PORT
      LAYER Metal1 ;
        RECT 6.040 1.770 11.050 2.150 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 9.734400 ;
    PORT
      LAYER Metal1 ;
        RECT 12.255 3.365 22.685 4.175 ;
        RECT 22.080 1.650 22.685 3.365 ;
        RECT 22.080 1.600 23.785 1.650 ;
        RECT 12.355 0.865 23.785 1.600 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 25.200 5.490 ;
        RECT 1.505 3.845 1.735 4.590 ;
        RECT 5.115 3.880 5.345 4.590 ;
        RECT 7.155 3.880 7.385 4.590 ;
        RECT 9.195 3.880 9.425 4.590 ;
        RECT 11.235 3.880 11.465 4.590 ;
        RECT 13.220 4.405 13.560 4.590 ;
        RECT 15.260 4.405 15.600 4.590 ;
        RECT 17.300 4.405 17.640 4.590 ;
        RECT 19.340 4.405 19.680 4.590 ;
        RECT 21.380 4.405 21.720 4.590 ;
        RECT 23.475 3.880 23.705 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 25.630 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 25.630 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 0.695 ;
        RECT 4.270 0.450 4.610 0.625 ;
        RECT 6.700 0.450 7.040 0.635 ;
        RECT 8.940 0.450 9.280 0.635 ;
        RECT 11.180 0.450 11.520 0.635 ;
        RECT 13.420 0.450 13.760 0.635 ;
        RECT 15.660 0.450 16.000 0.635 ;
        RECT 17.900 0.450 18.240 0.635 ;
        RECT 20.140 0.450 20.480 0.635 ;
        RECT 22.380 0.450 22.720 0.635 ;
        RECT 24.675 0.450 24.905 1.160 ;
        RECT 0.000 -0.450 25.200 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.485 3.170 0.715 3.750 ;
        RECT 2.925 3.675 3.155 4.255 ;
        RECT 2.925 3.445 4.635 3.675 ;
        RECT 4.405 3.360 4.635 3.445 ;
        RECT 10.215 3.360 10.445 3.940 ;
        RECT 0.485 2.940 3.595 3.170 ;
        RECT 1.805 1.600 2.035 2.940 ;
        RECT 3.365 2.415 3.595 2.940 ;
        RECT 3.945 2.185 4.175 3.215 ;
        RECT 0.190 1.370 2.035 1.600 ;
        RECT 3.145 1.955 4.175 2.185 ;
        RECT 4.405 3.140 10.445 3.360 ;
        RECT 4.405 2.910 11.695 3.140 ;
        RECT 3.145 1.490 3.375 1.955 ;
        RECT 4.405 1.655 4.635 2.910 ;
        RECT 11.465 2.790 11.695 2.910 ;
        RECT 11.465 2.450 21.210 2.790 ;
        RECT 2.485 1.085 3.375 1.490 ;
        RECT 3.605 1.315 4.635 1.655 ;
        RECT 11.675 1.830 21.035 2.150 ;
        RECT 11.675 1.490 11.905 1.830 ;
        RECT 5.635 1.260 11.905 1.490 ;
        RECT 5.635 1.085 8.105 1.260 ;
        RECT 2.485 0.865 8.105 1.085 ;
        RECT 2.485 0.855 5.865 0.865 ;
        RECT 2.485 0.680 2.715 0.855 ;
        RECT 7.875 0.680 8.105 0.865 ;
        RECT 10.115 0.680 10.345 1.260 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__bufz_12

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__bufz_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__bufz_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 31.920 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.545 2.330 1.575 2.710 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 13.535999 ;
    PORT
      LAYER Metal1 ;
        RECT 5.300 2.150 12.125 2.710 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 12.979199 ;
    PORT
      LAYER Metal1 ;
        RECT 14.520 3.365 29.090 4.175 ;
        RECT 28.530 1.650 29.090 3.365 ;
        RECT 28.530 1.635 30.505 1.650 ;
        RECT 14.595 0.865 30.505 1.635 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 31.920 5.490 ;
        RECT 1.505 3.845 1.735 4.590 ;
        RECT 4.860 4.370 5.200 4.590 ;
        RECT 6.900 4.370 7.240 4.590 ;
        RECT 8.940 4.370 9.280 4.590 ;
        RECT 11.280 4.370 11.620 4.590 ;
        RECT 13.500 4.405 13.840 4.590 ;
        RECT 15.540 4.405 15.880 4.590 ;
        RECT 17.580 4.405 17.920 4.590 ;
        RECT 19.620 4.405 19.960 4.590 ;
        RECT 21.660 4.405 22.000 4.590 ;
        RECT 23.700 4.405 24.040 4.590 ;
        RECT 25.740 4.405 26.080 4.590 ;
        RECT 27.780 4.405 28.120 4.590 ;
        RECT 29.875 3.880 30.105 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 32.350 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 32.350 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 0.695 ;
        RECT 4.270 0.450 4.610 0.625 ;
        RECT 6.700 0.450 7.040 0.635 ;
        RECT 8.940 0.450 9.280 0.635 ;
        RECT 11.180 0.450 11.520 0.635 ;
        RECT 13.405 0.450 13.780 0.635 ;
        RECT 15.660 0.450 16.000 0.635 ;
        RECT 17.900 0.450 18.240 0.635 ;
        RECT 20.140 0.450 20.480 0.635 ;
        RECT 22.380 0.450 22.720 0.635 ;
        RECT 24.620 0.450 24.960 0.635 ;
        RECT 26.860 0.450 27.200 0.635 ;
        RECT 29.100 0.450 29.440 0.635 ;
        RECT 31.395 0.450 31.625 1.160 ;
        RECT 0.000 -0.450 31.920 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.485 3.170 0.715 3.750 ;
        RECT 2.925 3.445 12.700 4.140 ;
        RECT 4.405 3.330 12.700 3.445 ;
        RECT 0.485 2.940 3.595 3.170 ;
        RECT 1.805 1.600 2.035 2.940 ;
        RECT 3.365 2.415 3.595 2.940 ;
        RECT 3.945 2.185 4.175 3.215 ;
        RECT 0.190 1.370 2.035 1.600 ;
        RECT 3.145 1.955 4.175 2.185 ;
        RECT 3.145 1.490 3.375 1.955 ;
        RECT 4.405 1.655 4.635 3.330 ;
        RECT 12.355 2.755 12.700 3.330 ;
        RECT 12.355 2.470 27.620 2.755 ;
        RECT 2.485 1.085 3.375 1.490 ;
        RECT 3.605 1.315 4.635 1.655 ;
        RECT 13.855 1.865 27.775 2.160 ;
        RECT 13.855 1.650 14.145 1.865 ;
        RECT 5.635 1.085 14.145 1.650 ;
        RECT 2.485 0.865 14.145 1.085 ;
        RECT 2.485 0.855 5.865 0.865 ;
        RECT 2.485 0.680 2.715 0.855 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__bufz_16

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.676500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.740 1.015 2.550 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.157200 ;
    PORT
      LAYER Metal1 ;
        RECT 2.565 1.590 2.895 3.775 ;
        RECT 2.390 1.210 2.895 1.590 ;
        RECT 2.665 0.710 2.895 1.210 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 3.360 5.490 ;
        RECT 1.365 3.240 1.595 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 3.790 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 3.790 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.050 ;
        RECT 0.000 -0.450 3.360 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 3.010 0.575 3.775 ;
        RECT 0.345 2.780 2.215 3.010 ;
        RECT 1.930 1.740 2.215 2.780 ;
        RECT 1.930 1.510 2.160 1.740 ;
        RECT 0.245 1.280 2.160 1.510 ;
        RECT 0.245 0.710 0.475 1.280 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.353000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 2.000 0.970 3.270 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.550600 ;
    PORT
      LAYER Metal1 ;
        RECT 2.665 3.960 3.110 4.300 ;
        RECT 2.880 1.215 3.110 3.960 ;
        RECT 2.330 0.710 3.110 1.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 4.480 5.490 ;
        RECT 1.265 3.960 1.495 4.590 ;
        RECT 3.685 3.550 3.915 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 4.910 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.215 ;
        RECT 3.785 0.450 4.015 1.215 ;
        RECT 0.000 -0.450 4.480 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.730 0.475 4.360 ;
        RECT 0.245 3.500 1.600 3.730 ;
        RECT 1.370 2.500 1.600 3.500 ;
        RECT 1.370 2.270 2.650 2.500 ;
        RECT 1.370 1.770 1.600 2.270 ;
        RECT 0.245 1.540 1.600 1.770 ;
        RECT 0.245 0.875 0.475 1.540 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.035000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.805 2.215 1.975 2.555 ;
        RECT 0.805 1.770 1.530 2.215 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.329000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.785 3.190 4.015 4.230 ;
        RECT 5.925 3.190 6.255 4.230 ;
        RECT 3.785 2.960 6.255 3.190 ;
        RECT 5.750 1.875 6.255 2.960 ;
        RECT 3.785 1.645 6.255 1.875 ;
        RECT 3.785 1.075 4.015 1.645 ;
        RECT 5.750 1.075 6.255 1.645 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.840 5.490 ;
        RECT 0.245 3.420 0.475 4.590 ;
        RECT 2.385 3.420 2.615 4.590 ;
        RECT 4.805 3.420 5.035 4.590 ;
        RECT 7.045 3.420 7.275 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 8.270 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.270 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.415 ;
        RECT 2.665 0.450 2.895 1.415 ;
        RECT 4.905 0.450 5.135 1.415 ;
        RECT 7.145 0.450 7.375 1.415 ;
        RECT 0.000 -0.450 7.840 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 3.190 1.595 4.230 ;
        RECT 1.365 2.960 2.435 3.190 ;
        RECT 2.205 2.555 2.435 2.960 ;
        RECT 2.205 2.215 4.745 2.555 ;
        RECT 2.205 1.360 2.435 2.215 ;
        RECT 1.310 1.130 2.435 1.360 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_3

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.706000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.805 2.215 1.975 2.555 ;
        RECT 0.805 1.770 1.530 2.215 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.101200 ;
    PORT
      LAYER Metal1 ;
        RECT 3.785 3.320 4.015 4.360 ;
        RECT 5.925 3.320 6.155 4.360 ;
        RECT 3.785 3.090 6.155 3.320 ;
        RECT 5.750 1.875 6.155 3.090 ;
        RECT 5.750 1.675 6.255 1.875 ;
        RECT 3.785 1.445 6.255 1.675 ;
        RECT 3.785 0.875 4.015 1.445 ;
        RECT 5.750 0.875 6.255 1.445 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.840 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.805 3.550 5.035 4.590 ;
        RECT 7.045 3.550 7.275 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 8.270 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.270 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.215 ;
        RECT 2.665 0.450 2.895 1.215 ;
        RECT 4.905 0.450 5.135 1.215 ;
        RECT 7.145 0.450 7.375 1.215 ;
        RECT 0.000 -0.450 7.840 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 1.365 3.090 2.435 3.320 ;
        RECT 2.205 2.555 2.435 3.090 ;
        RECT 2.205 2.215 4.745 2.555 ;
        RECT 2.205 1.160 2.435 2.215 ;
        RECT 1.310 0.930 2.435 1.160 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.560 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.412000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 2.215 4.205 2.650 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.202400 ;
    PORT
      LAYER Metal1 ;
        RECT 6.025 3.320 6.255 4.360 ;
        RECT 8.165 3.320 8.395 4.360 ;
        RECT 10.230 3.320 10.635 4.360 ;
        RECT 12.645 3.320 12.875 4.360 ;
        RECT 6.025 3.090 12.875 3.320 ;
        RECT 9.150 1.745 9.650 3.090 ;
        RECT 6.025 1.515 12.975 1.745 ;
        RECT 6.025 0.945 6.255 1.515 ;
        RECT 8.265 0.945 8.495 1.515 ;
        RECT 10.505 0.945 10.735 1.515 ;
        RECT 12.745 0.945 12.975 1.515 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 14.560 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.875 4.855 4.590 ;
        RECT 7.045 3.550 7.275 4.590 ;
        RECT 9.285 3.550 9.515 4.590 ;
        RECT 11.525 3.550 11.755 4.590 ;
        RECT 13.765 3.550 13.995 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 14.990 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.990 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.285 ;
        RECT 2.485 0.450 2.715 1.285 ;
        RECT 4.725 0.450 4.955 1.285 ;
        RECT 7.145 0.450 7.375 1.285 ;
        RECT 9.385 0.450 9.615 1.215 ;
        RECT 11.625 0.450 11.855 1.215 ;
        RECT 13.865 0.450 14.095 1.285 ;
        RECT 0.000 -0.450 14.560 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.505 3.320 3.735 4.360 ;
        RECT 1.365 3.090 4.665 3.320 ;
        RECT 4.435 2.650 4.665 3.090 ;
        RECT 4.435 2.270 8.920 2.650 ;
        RECT 9.880 2.270 13.510 2.650 ;
        RECT 4.435 1.745 4.665 2.270 ;
        RECT 1.365 1.515 4.665 1.745 ;
        RECT 1.365 0.945 1.595 1.515 ;
        RECT 3.605 0.945 3.835 1.515 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_8

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 8.118000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.275 2.215 6.675 2.555 ;
        RECT 1.275 1.770 6.010 2.215 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 9.303599 ;
    PORT
      LAYER Metal1 ;
        RECT 8.485 3.320 8.715 4.360 ;
        RECT 10.625 3.320 10.855 4.360 ;
        RECT 12.865 3.320 13.095 4.360 ;
        RECT 14.710 3.320 15.335 4.360 ;
        RECT 17.345 3.320 17.575 4.360 ;
        RECT 19.585 3.320 19.815 4.360 ;
        RECT 8.485 3.090 19.815 3.320 ;
        RECT 13.465 1.540 14.350 3.090 ;
        RECT 8.485 1.310 19.915 1.540 ;
        RECT 8.485 1.180 8.715 1.310 ;
        RECT 10.725 0.740 10.955 1.310 ;
        RECT 12.965 0.740 13.195 1.310 ;
        RECT 15.205 0.740 15.435 1.310 ;
        RECT 17.445 0.740 17.675 1.310 ;
        RECT 19.685 1.180 19.915 1.310 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 21.280 5.490 ;
        RECT 0.465 3.550 0.695 4.590 ;
        RECT 2.605 3.550 2.835 4.590 ;
        RECT 4.845 3.550 5.075 4.590 ;
        RECT 7.365 3.875 7.595 4.590 ;
        RECT 9.505 3.550 9.735 4.590 ;
        RECT 11.745 3.550 11.975 4.590 ;
        RECT 13.985 3.550 14.215 4.590 ;
        RECT 16.225 3.550 16.455 4.590 ;
        RECT 18.465 3.550 18.695 4.590 ;
        RECT 20.705 3.550 20.935 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 21.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 21.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.315 ;
        RECT 2.705 0.450 2.935 1.080 ;
        RECT 4.945 0.450 5.175 1.080 ;
        RECT 7.185 0.450 7.415 1.080 ;
        RECT 9.605 0.450 9.835 1.080 ;
        RECT 11.845 0.450 12.075 1.080 ;
        RECT 14.085 0.450 14.315 1.080 ;
        RECT 16.325 0.450 16.555 1.080 ;
        RECT 18.565 0.450 18.795 1.080 ;
        RECT 20.805 0.450 21.035 1.080 ;
        RECT 0.000 -0.450 21.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.585 3.320 1.815 4.360 ;
        RECT 3.725 3.320 3.955 4.360 ;
        RECT 5.965 3.320 6.195 4.360 ;
        RECT 1.585 3.090 7.135 3.320 ;
        RECT 6.905 2.555 7.135 3.090 ;
        RECT 6.905 2.215 13.205 2.555 ;
        RECT 14.580 2.215 19.980 2.555 ;
        RECT 6.905 1.540 7.135 2.215 ;
        RECT 1.585 1.310 7.135 1.540 ;
        RECT 1.585 1.110 1.815 1.310 ;
        RECT 3.825 1.110 4.055 1.310 ;
        RECT 6.065 1.110 6.295 1.310 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_12

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.000 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 10.823999 ;
    PORT
      LAYER Metal1 ;
        RECT 0.685 2.125 7.965 2.840 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 12.404799 ;
    PORT
      LAYER Metal1 ;
        RECT 10.505 3.320 10.735 4.360 ;
        RECT 12.645 3.320 12.875 4.360 ;
        RECT 14.885 3.320 15.115 4.360 ;
        RECT 17.125 3.320 17.355 4.360 ;
        RECT 19.365 3.320 19.595 4.360 ;
        RECT 21.605 3.320 21.835 4.360 ;
        RECT 23.845 3.320 24.075 4.360 ;
        RECT 26.085 3.320 26.315 4.360 ;
        RECT 10.505 3.090 26.315 3.320 ;
        RECT 17.985 1.895 18.735 3.090 ;
        RECT 10.505 1.745 18.735 1.895 ;
        RECT 10.505 1.665 26.415 1.745 ;
        RECT 10.505 1.515 12.975 1.665 ;
        RECT 10.505 0.945 10.735 1.515 ;
        RECT 12.745 0.945 12.975 1.515 ;
        RECT 14.985 0.945 15.215 1.665 ;
        RECT 17.225 1.515 26.415 1.665 ;
        RECT 17.225 0.945 17.455 1.515 ;
        RECT 19.465 0.945 19.695 1.515 ;
        RECT 21.705 0.945 21.935 1.515 ;
        RECT 23.945 0.945 24.175 1.515 ;
        RECT 26.185 0.945 26.415 1.515 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 28.000 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
        RECT 9.105 3.875 9.335 4.590 ;
        RECT 11.525 3.550 11.755 4.590 ;
        RECT 13.765 3.550 13.995 4.590 ;
        RECT 16.005 3.550 16.235 4.590 ;
        RECT 18.245 3.550 18.475 4.590 ;
        RECT 20.485 3.550 20.715 4.590 ;
        RECT 22.725 3.550 22.955 4.590 ;
        RECT 24.965 3.550 25.195 4.590 ;
        RECT 27.205 3.550 27.435 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 28.430 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 28.430 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.285 ;
        RECT 2.485 0.450 2.715 1.285 ;
        RECT 4.725 0.450 4.955 1.285 ;
        RECT 6.965 0.450 7.195 1.285 ;
        RECT 9.205 0.450 9.435 1.285 ;
        RECT 11.625 0.450 11.855 1.285 ;
        RECT 13.865 0.450 14.095 1.285 ;
        RECT 16.105 0.450 16.335 1.215 ;
        RECT 18.345 0.450 18.575 1.215 ;
        RECT 20.585 0.450 20.815 1.285 ;
        RECT 22.825 0.450 23.055 1.215 ;
        RECT 25.065 0.450 25.295 1.215 ;
        RECT 27.305 0.450 27.535 1.285 ;
        RECT 0.000 -0.450 28.000 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.505 3.320 3.735 4.360 ;
        RECT 5.745 3.320 5.975 4.360 ;
        RECT 8.085 3.320 8.550 4.360 ;
        RECT 1.365 3.090 8.550 3.320 ;
        RECT 8.320 2.555 8.550 3.090 ;
        RECT 8.320 2.215 17.105 2.555 ;
        RECT 18.965 2.215 26.245 2.555 ;
        RECT 8.320 1.745 8.550 2.215 ;
        RECT 1.365 1.515 8.550 1.745 ;
        RECT 1.365 0.945 1.595 1.515 ;
        RECT 3.605 0.945 3.835 1.515 ;
        RECT 5.845 0.945 6.075 1.515 ;
        RECT 8.085 0.945 8.550 1.515 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_16

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_20
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 ;
  ORIGIN 0.000 0.000 ;
  SIZE 34.720 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 13.530000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.685 2.215 9.845 2.650 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 15.506000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.745 3.320 12.975 4.360 ;
        RECT 14.885 3.320 15.115 4.360 ;
        RECT 17.125 3.320 17.355 4.360 ;
        RECT 19.365 3.320 19.595 4.360 ;
        RECT 21.605 3.320 21.835 4.360 ;
        RECT 23.845 3.320 24.075 4.360 ;
        RECT 26.085 3.320 26.315 4.360 ;
        RECT 28.325 3.320 28.555 4.360 ;
        RECT 30.565 3.320 30.795 4.360 ;
        RECT 32.805 3.320 33.035 4.360 ;
        RECT 12.745 3.090 33.035 3.320 ;
        RECT 22.465 1.745 23.215 3.090 ;
        RECT 12.745 1.675 23.215 1.745 ;
        RECT 12.745 1.515 33.135 1.675 ;
        RECT 12.745 0.945 13.005 1.515 ;
        RECT 14.985 0.945 15.215 1.515 ;
        RECT 17.225 0.945 17.455 1.515 ;
        RECT 19.465 0.945 19.695 1.515 ;
        RECT 21.705 1.445 33.135 1.515 ;
        RECT 21.705 0.945 21.935 1.445 ;
        RECT 23.945 0.945 24.175 1.445 ;
        RECT 26.185 0.945 26.415 1.445 ;
        RECT 28.425 0.945 28.655 1.445 ;
        RECT 30.665 0.945 30.895 1.445 ;
        RECT 32.905 0.945 33.135 1.445 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 34.720 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
        RECT 9.105 3.550 9.335 4.590 ;
        RECT 11.345 3.875 11.575 4.590 ;
        RECT 13.765 3.550 13.995 4.590 ;
        RECT 16.005 3.550 16.235 4.590 ;
        RECT 18.245 3.550 18.475 4.590 ;
        RECT 20.485 3.550 20.715 4.590 ;
        RECT 22.725 3.550 22.955 4.590 ;
        RECT 24.965 3.550 25.195 4.590 ;
        RECT 27.205 3.550 27.435 4.590 ;
        RECT 29.445 3.550 29.675 4.590 ;
        RECT 31.685 3.550 31.915 4.590 ;
        RECT 33.925 3.550 34.155 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 35.150 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 35.150 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.285 ;
        RECT 2.485 0.450 2.715 1.285 ;
        RECT 4.725 0.450 4.955 1.285 ;
        RECT 6.965 0.450 7.195 1.285 ;
        RECT 9.205 0.450 9.435 1.285 ;
        RECT 11.445 0.450 11.675 1.285 ;
        RECT 13.865 0.450 14.095 1.285 ;
        RECT 16.105 0.450 16.335 1.285 ;
        RECT 18.345 0.450 18.575 1.285 ;
        RECT 20.585 0.450 20.815 1.215 ;
        RECT 22.825 0.450 23.055 1.215 ;
        RECT 25.065 0.450 25.295 1.215 ;
        RECT 27.305 0.450 27.535 1.215 ;
        RECT 29.545 0.450 29.775 1.215 ;
        RECT 31.785 0.450 32.015 1.215 ;
        RECT 34.025 0.450 34.255 1.285 ;
        RECT 0.000 -0.450 34.720 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.505 3.320 3.735 4.360 ;
        RECT 5.745 3.320 5.975 4.360 ;
        RECT 7.985 3.320 8.215 4.360 ;
        RECT 10.225 3.320 10.455 4.360 ;
        RECT 1.365 3.090 10.455 3.320 ;
        RECT 10.225 2.650 10.455 3.090 ;
        RECT 10.225 2.215 21.225 2.650 ;
        RECT 23.445 2.215 32.605 2.650 ;
        RECT 10.225 1.745 10.555 2.215 ;
        RECT 1.365 1.515 10.555 1.745 ;
        RECT 1.365 0.945 1.595 1.515 ;
        RECT 3.605 0.945 3.835 1.515 ;
        RECT 5.845 0.945 6.075 1.515 ;
        RECT 8.085 0.945 8.315 1.515 ;
        RECT 10.325 0.945 10.555 1.515 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_20

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkinv_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkinv_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.240 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.353000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 1.830 0.970 2.530 ;
        RECT 0.710 1.210 0.970 1.830 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.126400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 0.945 1.595 4.360 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 2.240 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 2.670 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 2.670 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.285 ;
        RECT 0.000 -0.450 2.240 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__clkinv_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkinv_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkinv_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.706000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.360 2.270 1.640 2.710 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.514200 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.830 1.595 4.360 ;
        RECT 1.365 3.550 2.100 3.830 ;
        RECT 1.830 2.890 2.100 3.550 ;
        RECT 1.870 2.040 2.100 2.890 ;
        RECT 1.365 1.810 2.100 2.040 ;
        RECT 1.365 0.945 1.595 1.810 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 3.360 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 3.790 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 3.790 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.285 ;
        RECT 2.485 0.450 2.715 1.285 ;
        RECT 0.000 -0.450 3.360 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__clkinv_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkinv_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkinv_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.059000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.685 2.215 2.325 2.710 ;
        RECT 1.830 1.770 2.090 2.215 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.640600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.505 3.320 3.835 4.360 ;
        RECT 1.365 3.090 3.835 3.320 ;
        RECT 3.510 1.440 3.835 3.090 ;
        RECT 1.365 1.210 3.835 1.440 ;
        RECT 1.365 0.680 1.595 1.210 ;
        RECT 3.605 0.680 3.835 1.210 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 4.480 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 4.910 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.020 ;
        RECT 2.485 0.450 2.715 0.980 ;
        RECT 0.000 -0.450 4.480 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__clkinv_3

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkinv_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkinv_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.412000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 2.270 2.380 2.650 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.028400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.500 3.320 3.835 4.360 ;
        RECT 1.365 3.090 3.835 3.320 ;
        RECT 2.950 1.745 3.835 3.090 ;
        RECT 1.365 1.515 3.835 1.745 ;
        RECT 1.365 0.945 1.595 1.515 ;
        RECT 3.600 0.945 3.835 1.515 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.600 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.285 ;
        RECT 2.485 0.450 2.715 1.285 ;
        RECT 4.725 0.450 4.955 1.285 ;
        RECT 0.000 -0.450 5.600 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__clkinv_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkinv_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkinv_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 10.823999 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 2.265 4.260 2.645 ;
        RECT 5.360 2.215 8.880 2.650 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.056800 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.505 3.320 3.735 4.360 ;
        RECT 5.745 3.320 5.975 4.360 ;
        RECT 7.985 3.320 8.215 4.360 ;
        RECT 1.365 3.090 8.215 3.320 ;
        RECT 4.630 1.745 5.130 3.090 ;
        RECT 1.365 1.515 8.315 1.745 ;
        RECT 1.365 0.945 1.625 1.515 ;
        RECT 3.605 0.945 3.835 1.515 ;
        RECT 5.845 0.945 6.075 1.515 ;
        RECT 8.085 0.945 8.315 1.515 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 10.080 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
        RECT 9.105 3.550 9.335 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 10.510 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 10.510 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.285 ;
        RECT 2.485 0.450 2.715 1.285 ;
        RECT 4.725 0.450 4.955 1.285 ;
        RECT 6.965 0.450 7.195 1.285 ;
        RECT 9.205 0.450 9.435 1.285 ;
        RECT 0.000 -0.450 10.080 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__clkinv_8

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkinv_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkinv_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.560 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 16.236000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 2.270 6.140 2.650 ;
        RECT 7.660 2.270 13.170 2.650 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 9.085199 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.505 3.320 3.735 4.360 ;
        RECT 5.745 3.320 5.975 4.360 ;
        RECT 7.985 3.320 8.215 4.360 ;
        RECT 10.225 3.320 10.455 4.360 ;
        RECT 12.465 3.320 12.695 4.360 ;
        RECT 1.365 3.090 12.695 3.320 ;
        RECT 6.370 1.745 7.120 3.090 ;
        RECT 1.365 1.515 12.795 1.745 ;
        RECT 1.365 0.945 1.595 1.515 ;
        RECT 3.605 0.945 3.835 1.515 ;
        RECT 5.845 0.945 6.075 1.515 ;
        RECT 8.085 0.945 8.315 1.515 ;
        RECT 10.325 0.945 10.555 1.515 ;
        RECT 12.565 0.945 12.795 1.515 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 14.560 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
        RECT 9.105 3.550 9.335 4.590 ;
        RECT 11.345 3.550 11.575 4.590 ;
        RECT 13.585 3.550 13.815 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 14.990 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.990 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.285 ;
        RECT 2.485 0.450 2.715 1.285 ;
        RECT 4.725 0.450 4.955 1.285 ;
        RECT 6.965 0.450 7.195 1.285 ;
        RECT 9.205 0.450 9.435 1.285 ;
        RECT 11.445 0.450 11.675 1.285 ;
        RECT 13.685 0.450 13.915 1.285 ;
        RECT 0.000 -0.450 14.560 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__clkinv_12

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkinv_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkinv_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.040 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 21.647999 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 2.270 8.020 2.650 ;
        RECT 9.295 2.270 16.685 2.650 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 12.113600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.505 3.320 3.735 4.360 ;
        RECT 5.745 3.320 5.975 4.360 ;
        RECT 7.985 3.320 8.215 4.360 ;
        RECT 10.225 3.320 10.455 4.360 ;
        RECT 12.465 3.320 12.695 4.360 ;
        RECT 14.705 3.320 14.935 4.360 ;
        RECT 16.945 3.320 17.175 4.360 ;
        RECT 1.365 3.090 17.175 3.320 ;
        RECT 8.265 1.745 9.065 3.090 ;
        RECT 1.365 1.515 17.275 1.745 ;
        RECT 1.365 0.945 1.625 1.515 ;
        RECT 3.605 0.945 3.835 1.515 ;
        RECT 5.845 0.945 6.075 1.515 ;
        RECT 8.085 0.945 8.315 1.515 ;
        RECT 10.325 0.945 10.555 1.515 ;
        RECT 12.565 0.945 12.795 1.515 ;
        RECT 14.805 0.945 15.035 1.515 ;
        RECT 17.045 0.945 17.275 1.515 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 19.040 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
        RECT 9.105 3.550 9.335 4.590 ;
        RECT 11.345 3.550 11.575 4.590 ;
        RECT 13.585 3.550 13.815 4.590 ;
        RECT 15.825 3.550 16.055 4.590 ;
        RECT 18.065 3.550 18.295 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 19.470 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 19.470 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.285 ;
        RECT 2.485 0.450 2.715 1.285 ;
        RECT 4.725 0.450 4.955 1.285 ;
        RECT 6.965 0.450 7.195 1.285 ;
        RECT 9.205 0.450 9.435 1.285 ;
        RECT 11.445 0.450 11.675 1.285 ;
        RECT 13.685 0.450 13.915 1.285 ;
        RECT 15.925 0.450 16.155 1.285 ;
        RECT 18.165 0.450 18.395 1.285 ;
        RECT 0.000 -0.450 19.040 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__clkinv_16

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkinv_20
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkinv_20 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 27.059999 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 2.270 9.900 2.650 ;
        RECT 11.110 2.270 20.380 2.650 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 15.141999 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.505 3.320 3.735 4.360 ;
        RECT 5.745 3.320 5.975 4.360 ;
        RECT 7.985 3.320 8.215 4.360 ;
        RECT 10.225 3.320 10.455 4.360 ;
        RECT 12.465 3.320 12.695 4.360 ;
        RECT 14.705 3.320 14.935 4.360 ;
        RECT 16.945 3.320 17.175 4.360 ;
        RECT 19.185 3.320 19.415 4.360 ;
        RECT 21.425 3.320 21.655 4.360 ;
        RECT 1.365 3.090 21.655 3.320 ;
        RECT 10.130 1.745 10.880 3.090 ;
        RECT 1.365 1.515 21.755 1.745 ;
        RECT 1.365 0.945 1.625 1.515 ;
        RECT 3.605 0.945 3.835 1.515 ;
        RECT 5.845 0.945 6.075 1.515 ;
        RECT 8.085 0.945 8.315 1.515 ;
        RECT 10.325 0.945 10.555 1.515 ;
        RECT 12.565 0.945 12.795 1.515 ;
        RECT 14.805 0.945 15.035 1.515 ;
        RECT 17.045 0.945 17.275 1.515 ;
        RECT 19.285 0.945 19.515 1.515 ;
        RECT 21.525 0.945 21.755 1.515 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 23.520 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
        RECT 9.105 3.550 9.335 4.590 ;
        RECT 11.345 3.550 11.575 4.590 ;
        RECT 13.585 3.550 13.815 4.590 ;
        RECT 15.825 3.550 16.055 4.590 ;
        RECT 18.065 3.550 18.295 4.590 ;
        RECT 20.305 3.550 20.535 4.590 ;
        RECT 22.545 3.550 22.775 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 23.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 23.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.285 ;
        RECT 2.485 0.450 2.715 1.285 ;
        RECT 4.725 0.450 4.955 1.285 ;
        RECT 6.965 0.450 7.195 1.285 ;
        RECT 9.205 0.450 9.435 1.285 ;
        RECT 11.445 0.450 11.675 1.285 ;
        RECT 13.685 0.450 13.915 1.285 ;
        RECT 15.925 0.450 16.155 1.285 ;
        RECT 18.165 0.450 18.395 1.285 ;
        RECT 20.405 0.450 20.635 1.285 ;
        RECT 22.645 0.450 22.875 1.285 ;
        RECT 0.000 -0.450 23.520 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__clkinv_20

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.800 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 2.330 4.330 2.710 ;
    END
  END D
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.235 1.570 2.710 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.710 1.315 15.055 3.215 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 16.800 5.490 ;
        RECT 1.365 3.425 1.595 4.590 ;
        RECT 3.305 3.610 3.535 4.590 ;
        RECT 7.405 3.140 7.635 4.590 ;
        RECT 12.545 3.905 12.775 4.590 ;
        RECT 15.845 3.875 16.075 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 17.230 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 17.230 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.205 0.450 3.435 1.130 ;
        RECT 7.625 0.450 7.855 0.625 ;
        RECT 12.765 0.450 12.995 0.625 ;
        RECT 15.945 0.450 16.175 1.165 ;
        RECT 0.000 -0.450 16.800 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.765 4.125 6.170 4.355 ;
        RECT 0.345 3.170 0.575 3.750 ;
        RECT 3.765 3.220 3.995 4.125 ;
        RECT 0.345 2.940 2.035 3.170 ;
        RECT 1.805 1.740 2.035 2.940 ;
        RECT 0.245 1.510 2.035 1.740 ;
        RECT 2.385 2.990 3.995 3.220 ;
        RECT 0.245 1.315 0.475 1.510 ;
        RECT 2.385 1.315 2.715 2.990 ;
        RECT 4.425 2.970 4.790 3.780 ;
        RECT 4.560 1.360 4.790 2.970 ;
        RECT 4.325 1.020 4.790 1.360 ;
        RECT 5.445 2.280 5.675 3.780 ;
        RECT 8.965 2.850 9.195 3.780 ;
        RECT 6.965 2.510 9.195 2.850 ;
        RECT 5.445 2.050 8.515 2.280 ;
        RECT 5.445 1.020 5.675 2.050 ;
        RECT 8.285 1.940 8.515 2.050 ;
        RECT 6.125 1.085 6.355 1.820 ;
        RECT 8.965 1.315 9.195 2.510 ;
        RECT 10.085 2.990 10.315 3.780 ;
        RECT 11.470 3.445 15.515 3.675 ;
        RECT 10.085 2.760 13.410 2.990 ;
        RECT 10.085 1.315 10.315 2.760 ;
        RECT 10.545 2.300 11.250 2.530 ;
        RECT 13.925 2.460 14.155 3.215 ;
        RECT 12.050 2.455 14.155 2.460 ;
        RECT 10.545 1.085 10.775 2.300 ;
        RECT 12.050 2.230 14.480 2.455 ;
        RECT 14.105 1.315 14.480 2.230 ;
        RECT 6.125 0.855 10.775 1.085 ;
        RECT 11.425 1.085 11.655 1.225 ;
        RECT 15.285 1.085 15.515 3.445 ;
        RECT 11.425 0.855 15.515 1.085 ;
        RECT 9.350 0.680 10.775 0.855 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnq_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.360 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 1.690 4.325 2.235 ;
    END
  END D
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.330 1.865 2.710 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 15.820 1.600 16.090 3.270 ;
        RECT 15.710 1.370 16.090 1.600 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.360 5.490 ;
        RECT 1.655 3.425 1.885 4.590 ;
        RECT 3.495 3.615 3.725 4.590 ;
        RECT 7.925 3.145 8.155 4.590 ;
        RECT 12.805 4.345 13.035 4.590 ;
        RECT 14.800 4.345 15.030 4.590 ;
        RECT 16.840 3.875 17.070 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 17.790 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 17.790 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.555 0.450 1.785 1.225 ;
        RECT 3.395 0.450 3.625 1.190 ;
        RECT 7.925 0.450 8.155 1.190 ;
        RECT 12.805 0.450 13.035 1.165 ;
        RECT 14.590 0.450 14.930 0.640 ;
        RECT 16.885 0.450 17.115 1.165 ;
        RECT 0.000 -0.450 17.360 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.955 4.130 6.690 4.360 ;
        RECT 0.635 3.170 0.865 3.750 ;
        RECT 3.955 3.215 4.185 4.130 ;
        RECT 0.635 2.940 2.325 3.170 ;
        RECT 2.095 1.740 2.325 2.940 ;
        RECT 0.435 1.510 2.325 1.740 ;
        RECT 2.675 2.985 4.185 3.215 ;
        RECT 0.435 1.315 0.665 1.510 ;
        RECT 2.675 1.315 2.905 2.985 ;
        RECT 4.515 2.975 4.790 3.785 ;
        RECT 4.560 1.080 4.790 2.975 ;
        RECT 5.965 2.285 6.195 3.785 ;
        RECT 8.945 2.855 9.175 3.785 ;
        RECT 7.485 2.625 9.175 2.855 ;
        RECT 7.485 2.515 7.715 2.625 ;
        RECT 8.365 2.285 8.595 2.395 ;
        RECT 5.965 2.055 8.595 2.285 ;
        RECT 8.945 2.285 9.175 2.625 ;
        RECT 10.385 2.880 10.615 3.785 ;
        RECT 11.785 3.690 16.550 3.920 ;
        RECT 11.785 3.110 12.015 3.690 ;
        RECT 10.385 2.650 13.530 2.880 ;
        RECT 8.945 2.055 9.495 2.285 ;
        RECT 5.965 1.080 6.195 2.055 ;
        RECT 6.590 1.595 9.035 1.825 ;
        RECT 8.805 0.910 9.035 1.595 ;
        RECT 9.265 1.315 9.495 2.055 ;
        RECT 10.385 1.315 10.615 2.650 ;
        RECT 13.190 2.470 13.530 2.650 ;
        RECT 11.170 2.190 11.550 2.420 ;
        RECT 11.170 0.910 11.400 2.190 ;
        RECT 13.825 2.150 14.055 3.215 ;
        RECT 12.310 2.060 14.055 2.150 ;
        RECT 12.310 1.920 15.525 2.060 ;
        RECT 13.870 1.830 15.525 1.920 ;
        RECT 11.630 1.395 13.640 1.625 ;
        RECT 11.630 1.370 11.970 1.395 ;
        RECT 13.410 1.140 13.640 1.395 ;
        RECT 13.870 1.370 14.210 1.830 ;
        RECT 16.320 1.140 16.550 3.690 ;
        RECT 13.410 0.910 16.550 1.140 ;
        RECT 8.805 0.680 11.400 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnq_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.430 2.330 4.330 2.710 ;
    END
  END D
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.330 1.705 2.710 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 15.710 2.890 18.290 3.230 ;
        RECT 17.785 1.640 18.290 2.890 ;
        RECT 15.710 1.370 18.290 1.640 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 19.600 5.490 ;
        RECT 1.495 3.425 1.725 4.590 ;
        RECT 3.435 3.515 3.665 4.590 ;
        RECT 7.535 3.045 7.765 4.590 ;
        RECT 12.805 4.345 13.035 4.590 ;
        RECT 14.745 4.345 14.975 4.590 ;
        RECT 16.785 4.345 17.015 4.590 ;
        RECT 18.825 4.345 19.055 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 20.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 20.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.495 0.450 1.725 1.225 ;
        RECT 3.335 0.450 3.565 1.145 ;
        RECT 7.755 0.450 7.985 0.625 ;
        RECT 12.750 0.450 13.090 0.640 ;
        RECT 14.590 0.450 14.930 0.640 ;
        RECT 16.830 0.450 17.170 0.640 ;
        RECT 19.125 0.450 19.355 1.165 ;
        RECT 0.000 -0.450 19.600 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.895 4.030 6.300 4.260 ;
        RECT 0.475 3.170 0.705 3.750 ;
        RECT 3.895 3.215 4.125 4.030 ;
        RECT 0.475 2.940 2.165 3.170 ;
        RECT 1.935 2.005 2.165 2.940 ;
        RECT 0.375 1.775 2.165 2.005 ;
        RECT 2.515 2.985 4.125 3.215 ;
        RECT 0.375 1.315 0.605 1.775 ;
        RECT 2.515 1.315 2.845 2.985 ;
        RECT 4.555 2.875 4.790 3.685 ;
        RECT 4.560 1.375 4.790 2.875 ;
        RECT 4.455 1.035 4.790 1.375 ;
        RECT 5.575 2.240 5.805 3.685 ;
        RECT 9.030 2.700 9.265 3.685 ;
        RECT 7.040 2.470 9.265 2.700 ;
        RECT 5.575 2.010 8.585 2.240 ;
        RECT 5.575 1.035 5.805 2.010 ;
        RECT 8.355 1.900 8.585 2.010 ;
        RECT 6.200 1.085 6.540 1.780 ;
        RECT 9.035 1.315 9.265 2.470 ;
        RECT 10.155 3.215 10.385 3.685 ;
        RECT 11.730 3.500 18.750 3.730 ;
        RECT 10.155 2.985 11.855 3.215 ;
        RECT 10.155 1.315 10.385 2.985 ;
        RECT 11.165 1.085 11.395 2.755 ;
        RECT 11.625 2.700 11.855 2.985 ;
        RECT 11.625 2.470 13.530 2.700 ;
        RECT 13.825 2.210 14.055 3.215 ;
        RECT 13.825 2.150 17.555 2.210 ;
        RECT 12.310 1.920 17.555 2.150 ;
        RECT 13.870 1.870 17.555 1.920 ;
        RECT 6.200 0.855 11.395 1.085 ;
        RECT 9.420 0.680 11.395 0.855 ;
        RECT 11.685 1.140 11.915 1.490 ;
        RECT 13.870 1.370 14.210 1.870 ;
        RECT 18.520 1.140 18.750 3.500 ;
        RECT 11.685 0.910 18.750 1.140 ;
        RECT 11.685 0.680 11.915 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnq_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnrnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnrnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.920 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.945 2.310 3.770 2.710 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.030000 ;
    PORT
      LAYER Metal1 ;
        RECT 13.590 1.210 13.910 2.025 ;
    END
  END RN
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.665 2.235 1.575 2.710 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 15.830 3.450 16.390 3.830 ;
        RECT 16.160 0.845 16.390 3.450 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.920 5.490 ;
        RECT 1.305 3.425 1.535 4.590 ;
        RECT 3.045 3.515 3.275 4.590 ;
        RECT 7.125 3.515 7.355 4.590 ;
        RECT 8.865 3.355 9.095 4.590 ;
        RECT 13.185 4.260 13.525 4.590 ;
        RECT 15.280 3.735 15.510 4.590 ;
        RECT 17.180 3.875 17.410 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 18.350 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 18.350 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.205 0.450 3.435 1.225 ;
        RECT 8.245 0.450 8.475 1.225 ;
        RECT 13.020 0.450 13.250 1.225 ;
        RECT 17.280 0.450 17.510 1.165 ;
        RECT 0.000 -0.450 17.920 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.505 3.975 5.755 4.315 ;
        RECT 0.285 3.170 0.515 3.750 ;
        RECT 2.325 3.285 2.555 3.685 ;
        RECT 3.505 3.285 3.735 3.975 ;
        RECT 0.285 2.940 2.035 3.170 ;
        RECT 1.805 1.740 2.035 2.940 ;
        RECT 0.245 1.510 2.035 1.740 ;
        RECT 2.325 3.055 3.735 3.285 ;
        RECT 0.245 1.315 0.475 1.510 ;
        RECT 2.325 1.315 2.715 3.055 ;
        RECT 4.065 1.510 4.295 3.685 ;
        RECT 5.085 2.995 5.315 3.685 ;
        RECT 6.105 3.275 6.335 3.855 ;
        RECT 8.145 3.275 8.375 3.855 ;
        RECT 6.105 3.045 8.375 3.275 ;
        RECT 5.085 2.815 5.670 2.995 ;
        RECT 5.085 2.765 9.590 2.815 ;
        RECT 5.445 2.585 9.590 2.765 ;
        RECT 4.065 1.280 4.610 1.510 ;
        RECT 5.445 1.225 5.675 2.585 ;
        RECT 9.885 2.360 10.115 3.995 ;
        RECT 9.640 2.180 10.115 2.360 ;
        RECT 6.670 2.130 10.115 2.180 ;
        RECT 10.780 3.765 14.950 3.995 ;
        RECT 10.780 3.185 11.135 3.765 ;
        RECT 6.125 1.685 6.355 2.025 ;
        RECT 6.670 1.950 9.865 2.130 ;
        RECT 6.125 1.455 9.405 1.685 ;
        RECT 9.175 0.995 9.405 1.455 ;
        RECT 9.635 1.225 9.865 1.950 ;
        RECT 10.320 0.995 10.550 2.025 ;
        RECT 10.780 1.225 11.010 3.185 ;
        RECT 11.345 0.995 11.575 3.065 ;
        RECT 11.900 1.225 12.155 3.525 ;
        RECT 12.580 3.295 14.490 3.525 ;
        RECT 12.580 2.725 12.810 3.295 ;
        RECT 14.260 2.495 14.490 3.295 ;
        RECT 14.720 2.725 14.950 3.765 ;
        RECT 14.260 2.265 15.930 2.495 ;
        RECT 15.440 1.975 15.930 2.265 ;
        RECT 15.440 1.315 15.670 1.975 ;
        RECT 9.175 0.765 11.575 0.995 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnrnq_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.945 1.770 3.895 2.150 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.255000 ;
    PORT
      LAYER Metal1 ;
        RECT 13.380 1.675 14.410 2.150 ;
    END
  END RN
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 1.575 2.245 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 17.510 3.450 17.915 3.830 ;
        RECT 17.685 0.845 17.915 3.450 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 19.600 5.490 ;
        RECT 1.365 3.425 1.595 4.590 ;
        RECT 3.225 3.045 3.455 4.590 ;
        RECT 7.305 3.515 7.535 4.590 ;
        RECT 9.045 3.440 9.275 4.590 ;
        RECT 13.525 4.345 13.755 4.590 ;
        RECT 15.845 3.875 16.075 4.590 ;
        RECT 16.665 3.875 16.895 4.590 ;
        RECT 18.705 3.875 18.935 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 20.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 20.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.450 1.650 1.080 ;
        RECT 3.205 0.450 3.435 1.310 ;
        RECT 8.425 0.450 8.655 1.310 ;
        RECT 13.425 0.450 13.655 1.310 ;
        RECT 16.565 0.450 16.795 1.165 ;
        RECT 18.805 0.450 19.035 1.165 ;
        RECT 0.000 -0.450 19.600 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.685 4.030 5.990 4.260 ;
        RECT 0.345 3.105 0.575 3.685 ;
        RECT 0.345 2.875 2.035 3.105 ;
        RECT 1.805 1.540 2.035 2.875 ;
        RECT 0.245 1.310 2.035 1.540 ;
        RECT 2.385 2.815 2.615 3.685 ;
        RECT 3.685 2.815 3.915 4.030 ;
        RECT 2.385 2.585 3.915 2.815 ;
        RECT 0.245 1.190 0.475 1.310 ;
        RECT 2.385 1.190 2.715 2.585 ;
        RECT 4.245 1.310 4.555 3.685 ;
        RECT 5.265 2.690 5.495 3.685 ;
        RECT 6.285 3.150 6.515 3.730 ;
        RECT 8.325 3.150 8.555 3.730 ;
        RECT 6.285 2.920 8.555 3.150 ;
        RECT 5.265 2.460 9.770 2.690 ;
        RECT 5.265 1.310 5.675 2.460 ;
        RECT 10.065 2.230 10.295 4.080 ;
        RECT 6.070 1.825 6.580 2.055 ;
        RECT 6.810 2.000 10.295 2.230 ;
        RECT 11.185 3.850 15.495 4.080 ;
        RECT 11.185 3.270 11.420 3.850 ;
        RECT 6.350 1.770 6.580 1.825 ;
        RECT 6.350 1.540 9.835 1.770 ;
        RECT 9.605 1.080 9.835 1.540 ;
        RECT 10.065 1.310 10.295 2.000 ;
        RECT 10.525 1.080 10.755 2.110 ;
        RECT 11.185 1.310 11.415 3.270 ;
        RECT 11.645 1.080 11.875 3.150 ;
        RECT 12.285 1.310 12.535 3.610 ;
        RECT 14.545 2.610 14.775 3.215 ;
        RECT 12.810 2.380 15.035 2.610 ;
        RECT 15.265 2.415 15.495 3.850 ;
        RECT 14.805 2.185 15.035 2.380 ;
        RECT 14.805 1.955 17.390 2.185 ;
        RECT 15.845 1.830 17.390 1.955 ;
        RECT 9.605 0.850 11.875 1.080 ;
        RECT 15.845 0.845 16.075 1.830 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnrnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnrnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.840 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.945 2.330 3.895 2.710 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.255000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.105 1.590 14.335 2.050 ;
        RECT 14.105 1.210 14.410 1.590 ;
    END
  END RN
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.235 1.575 2.710 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 17.685 3.295 17.915 3.685 ;
        RECT 19.725 3.295 20.175 3.685 ;
        RECT 17.685 2.875 20.175 3.295 ;
        RECT 19.715 1.655 20.175 2.875 ;
        RECT 17.685 1.395 20.175 1.655 ;
        RECT 17.685 0.845 17.915 1.395 ;
        RECT 19.750 0.815 20.175 1.395 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 21.840 5.490 ;
        RECT 1.365 3.425 1.595 4.590 ;
        RECT 3.225 3.615 3.455 4.590 ;
        RECT 7.305 3.615 7.535 4.590 ;
        RECT 9.045 3.380 9.275 4.590 ;
        RECT 13.525 4.345 13.755 4.590 ;
        RECT 15.845 3.875 16.075 4.590 ;
        RECT 16.665 3.875 16.895 4.590 ;
        RECT 18.705 3.875 18.935 4.590 ;
        RECT 20.745 3.875 20.975 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 22.270 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 22.270 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.205 0.450 3.435 1.250 ;
        RECT 8.725 0.450 8.955 1.250 ;
        RECT 13.425 0.450 13.655 1.250 ;
        RECT 16.565 0.450 16.795 1.165 ;
        RECT 18.805 0.450 19.035 1.165 ;
        RECT 21.045 0.450 21.275 1.165 ;
        RECT 0.000 -0.450 21.840 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.685 4.130 5.990 4.360 ;
        RECT 0.345 3.170 0.575 3.750 ;
        RECT 2.385 3.385 2.615 3.685 ;
        RECT 3.685 3.385 3.915 4.130 ;
        RECT 0.345 2.940 2.035 3.170 ;
        RECT 1.805 2.005 2.035 2.940 ;
        RECT 0.245 1.775 2.035 2.005 ;
        RECT 2.385 3.155 3.915 3.385 ;
        RECT 0.245 1.315 0.475 1.775 ;
        RECT 2.385 1.315 2.715 3.155 ;
        RECT 4.245 1.250 4.555 3.785 ;
        RECT 5.265 2.915 5.495 3.785 ;
        RECT 6.285 3.375 6.515 3.955 ;
        RECT 8.325 3.375 8.555 3.955 ;
        RECT 6.285 3.145 8.555 3.375 ;
        RECT 5.265 2.685 9.770 2.915 ;
        RECT 5.265 1.250 5.675 2.685 ;
        RECT 10.065 2.455 10.295 4.020 ;
        RECT 6.810 2.225 10.295 2.455 ;
        RECT 6.070 1.765 9.835 1.995 ;
        RECT 9.605 1.020 9.835 1.765 ;
        RECT 10.065 1.250 10.295 2.225 ;
        RECT 11.185 3.790 15.300 4.020 ;
        RECT 11.185 3.210 11.420 3.790 ;
        RECT 10.525 1.020 10.755 2.050 ;
        RECT 11.185 1.250 11.415 3.210 ;
        RECT 11.645 1.020 11.875 3.090 ;
        RECT 12.285 1.250 12.535 3.550 ;
        RECT 14.555 2.550 14.840 3.215 ;
        RECT 12.810 2.320 14.840 2.550 ;
        RECT 15.070 2.700 15.300 3.790 ;
        RECT 15.070 2.470 15.550 2.700 ;
        RECT 14.610 2.240 14.840 2.320 ;
        RECT 15.845 2.240 19.485 2.275 ;
        RECT 14.610 2.015 19.485 2.240 ;
        RECT 14.610 2.010 16.075 2.015 ;
        RECT 9.605 0.790 11.875 1.020 ;
        RECT 15.845 0.845 16.075 2.010 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnrnq_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.945 2.330 3.975 2.710 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018000 ;
    PORT
      LAYER Metal1 ;
        RECT 16.965 2.200 17.770 2.760 ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.545 2.330 15.575 2.805 ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.235 1.575 2.710 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.705 1.655 20.010 3.685 ;
        RECT 19.685 0.845 20.010 1.655 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 21.280 5.490 ;
        RECT 1.365 3.425 1.595 4.590 ;
        RECT 3.305 3.515 3.535 4.590 ;
        RECT 7.605 4.375 7.835 4.590 ;
        RECT 10.805 4.375 11.035 4.590 ;
        RECT 14.850 3.950 15.190 4.590 ;
        RECT 16.890 3.950 17.230 4.590 ;
        RECT 18.985 3.425 19.215 4.590 ;
        RECT 20.725 3.875 20.955 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 21.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 21.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.205 0.450 3.435 1.425 ;
        RECT 8.945 0.450 9.175 1.425 ;
        RECT 16.945 0.450 17.175 1.225 ;
        RECT 20.805 0.450 21.035 1.165 ;
        RECT 0.000 -0.450 21.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.765 4.145 6.070 4.260 ;
        RECT 12.485 4.145 12.715 4.315 ;
        RECT 3.765 3.915 12.715 4.145 ;
        RECT 0.345 3.170 0.575 3.750 ;
        RECT 2.385 3.285 2.615 3.685 ;
        RECT 3.765 3.285 3.995 3.915 ;
        RECT 0.345 2.940 2.035 3.170 ;
        RECT 1.805 1.740 2.035 2.940 ;
        RECT 0.245 1.510 2.035 1.740 ;
        RECT 2.385 3.055 3.995 3.285 ;
        RECT 0.245 1.315 0.655 1.510 ;
        RECT 2.385 1.315 2.715 3.055 ;
        RECT 4.325 1.315 4.555 3.685 ;
        RECT 5.345 2.915 5.575 3.685 ;
        RECT 6.365 3.345 9.075 3.685 ;
        RECT 9.565 3.445 12.275 3.685 ;
        RECT 9.565 3.345 11.655 3.445 ;
        RECT 5.345 2.685 10.235 2.915 ;
        RECT 5.825 1.315 6.055 2.685 ;
        RECT 10.005 2.575 10.235 2.685 ;
        RECT 7.105 2.345 7.335 2.455 ;
        RECT 11.390 2.345 11.655 3.345 ;
        RECT 12.045 2.875 12.275 3.445 ;
        RECT 13.065 3.455 18.690 3.685 ;
        RECT 7.105 2.115 11.655 2.345 ;
        RECT 6.285 1.885 6.515 2.115 ;
        RECT 6.285 1.655 11.195 1.885 ;
        RECT 10.965 0.910 11.195 1.655 ;
        RECT 11.425 1.315 11.655 2.115 ;
        RECT 13.065 1.655 13.295 3.455 ;
        RECT 14.085 2.115 14.315 3.215 ;
        RECT 12.545 1.315 13.295 1.655 ;
        RECT 13.665 2.100 14.315 2.115 ;
        RECT 15.925 2.100 16.155 3.215 ;
        RECT 17.965 2.885 18.230 3.225 ;
        RECT 13.665 1.870 16.155 2.100 ;
        RECT 16.505 1.970 16.735 2.115 ;
        RECT 18.000 2.025 18.230 2.885 ;
        RECT 18.460 2.415 18.690 3.455 ;
        RECT 18.910 2.025 19.475 2.315 ;
        RECT 18.000 1.975 19.475 2.025 ;
        RECT 18.000 1.970 19.135 1.975 ;
        RECT 13.665 1.315 13.895 1.870 ;
        RECT 14.325 0.910 14.555 1.640 ;
        RECT 14.985 1.315 15.215 1.870 ;
        RECT 16.505 1.740 19.135 1.970 ;
        RECT 18.905 1.315 19.135 1.740 ;
        RECT 10.965 0.680 14.555 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.400 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.390 1.770 4.330 2.150 ;
        RECT 3.990 1.210 4.330 1.770 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018000 ;
    PORT
      LAYER Metal1 ;
        RECT 16.755 2.320 17.770 2.710 ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018000 ;
    PORT
      LAYER Metal1 ;
        RECT 15.270 1.210 15.610 2.060 ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 1.580 2.150 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 20.670 0.845 21.130 3.830 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 22.400 5.490 ;
        RECT 1.470 3.425 1.700 4.590 ;
        RECT 3.210 3.595 3.440 4.590 ;
        RECT 7.690 4.480 7.920 4.590 ;
        RECT 10.830 4.480 11.060 4.590 ;
        RECT 14.775 3.960 15.115 4.590 ;
        RECT 16.815 3.960 17.155 4.590 ;
        RECT 18.910 3.905 19.140 4.590 ;
        RECT 19.650 3.875 19.880 4.590 ;
        RECT 21.690 3.875 21.920 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 22.830 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 22.830 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.415 0.450 1.755 1.045 ;
        RECT 3.440 0.450 3.670 1.425 ;
        RECT 8.875 0.450 9.215 1.370 ;
        RECT 16.870 0.450 17.100 1.225 ;
        RECT 19.550 0.450 19.780 1.165 ;
        RECT 21.790 0.450 22.020 1.165 ;
        RECT 0.000 -0.450 22.400 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.670 4.250 5.975 4.340 ;
        RECT 12.455 4.250 12.795 4.350 ;
        RECT 3.670 4.020 12.795 4.250 ;
        RECT 0.450 3.105 0.680 3.685 ;
        RECT 3.670 3.215 3.900 4.020 ;
        RECT 0.450 2.875 2.140 3.105 ;
        RECT 1.910 1.540 2.140 2.875 ;
        RECT 0.350 1.310 2.140 1.540 ;
        RECT 2.490 2.985 3.900 3.215 ;
        RECT 4.230 3.185 4.460 3.765 ;
        RECT 0.350 1.190 0.580 1.310 ;
        RECT 2.490 1.190 2.820 2.985 ;
        RECT 4.230 2.955 4.790 3.185 ;
        RECT 4.560 1.315 4.790 2.955 ;
        RECT 5.250 2.750 5.480 3.765 ;
        RECT 6.520 3.450 9.160 3.790 ;
        RECT 6.520 2.980 6.750 3.450 ;
        RECT 9.650 3.305 9.880 3.790 ;
        RECT 9.650 3.075 10.780 3.305 ;
        RECT 9.650 2.980 9.880 3.075 ;
        RECT 10.090 2.750 10.320 2.845 ;
        RECT 5.250 2.520 10.320 2.750 ;
        RECT 5.680 1.315 5.910 2.520 ;
        RECT 10.090 2.505 10.320 2.520 ;
        RECT 10.550 2.455 10.780 3.075 ;
        RECT 12.070 2.455 12.300 3.775 ;
        RECT 7.100 2.275 10.005 2.290 ;
        RECT 10.550 2.275 12.300 2.455 ;
        RECT 7.100 2.225 12.300 2.275 ;
        RECT 13.090 3.730 14.635 3.775 ;
        RECT 13.090 3.545 18.690 3.730 ;
        RECT 6.360 1.720 6.590 2.115 ;
        RECT 7.100 2.060 11.440 2.225 ;
        RECT 7.100 1.950 7.330 2.060 ;
        RECT 9.920 2.045 11.440 2.060 ;
        RECT 7.530 1.720 9.835 1.830 ;
        RECT 6.360 1.600 9.835 1.720 ;
        RECT 6.360 1.490 7.730 1.600 ;
        RECT 9.605 0.910 9.835 1.600 ;
        RECT 11.210 1.315 11.440 2.045 ;
        RECT 13.090 1.900 13.320 3.545 ;
        RECT 14.495 3.500 18.690 3.545 ;
        RECT 12.330 1.670 13.320 1.900 ;
        RECT 12.330 1.315 12.560 1.670 ;
        RECT 14.110 1.480 14.340 3.305 ;
        RECT 13.450 1.370 14.340 1.480 ;
        RECT 13.450 1.140 15.040 1.370 ;
        RECT 14.810 0.980 15.040 1.140 ;
        RECT 15.850 0.980 16.080 3.225 ;
        RECT 17.890 2.910 18.230 3.250 ;
        RECT 18.000 2.115 18.230 2.910 ;
        RECT 18.460 2.425 18.690 3.500 ;
        RECT 18.000 2.090 20.320 2.115 ;
        RECT 16.375 1.860 20.320 2.090 ;
        RECT 18.830 1.775 20.320 1.860 ;
        RECT 18.830 1.315 19.060 1.775 ;
        RECT 9.605 0.680 14.380 0.910 ;
        RECT 14.810 0.750 16.080 0.980 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 24.640 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.055 2.330 3.890 2.710 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018000 ;
    PORT
      LAYER Metal1 ;
        RECT 16.950 2.710 17.210 3.270 ;
        RECT 16.950 2.480 17.515 2.710 ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018000 ;
    PORT
      LAYER Metal1 ;
        RECT 15.270 1.770 15.530 2.765 ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.295 1.570 2.710 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 20.590 3.105 20.820 3.685 ;
        RECT 22.630 3.105 23.060 3.685 ;
        RECT 20.590 2.875 23.060 3.105 ;
        RECT 22.665 1.655 23.060 2.875 ;
        RECT 20.590 1.395 23.060 1.655 ;
        RECT 20.590 0.845 20.820 1.395 ;
        RECT 22.550 0.815 23.060 1.395 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 24.640 5.490 ;
        RECT 1.365 3.425 1.595 4.590 ;
        RECT 3.205 3.515 3.435 4.590 ;
        RECT 7.465 4.490 7.695 4.590 ;
        RECT 10.665 4.490 10.895 4.590 ;
        RECT 14.695 3.960 15.035 4.590 ;
        RECT 16.735 3.960 17.075 4.590 ;
        RECT 18.830 3.435 19.060 4.590 ;
        RECT 19.570 3.875 19.800 4.590 ;
        RECT 21.610 3.875 21.840 4.590 ;
        RECT 23.650 3.875 23.880 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 25.070 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 25.070 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.205 0.450 3.435 1.425 ;
        RECT 8.405 0.450 8.635 1.425 ;
        RECT 16.790 0.450 17.020 1.225 ;
        RECT 19.470 0.450 19.700 1.165 ;
        RECT 21.710 0.450 21.940 1.165 ;
        RECT 23.950 0.450 24.180 1.165 ;
        RECT 0.000 -0.450 24.640 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.665 4.030 12.630 4.260 ;
        RECT 0.345 3.170 0.575 3.750 ;
        RECT 2.385 3.285 2.615 3.685 ;
        RECT 3.665 3.285 3.895 4.030 ;
        RECT 0.345 2.940 2.035 3.170 ;
        RECT 1.805 2.005 2.035 2.940 ;
        RECT 0.245 1.775 2.035 2.005 ;
        RECT 2.385 3.055 3.895 3.285 ;
        RECT 0.245 1.315 0.475 1.775 ;
        RECT 2.385 1.315 2.715 3.055 ;
        RECT 4.225 1.315 4.555 3.685 ;
        RECT 5.245 2.915 5.475 3.685 ;
        RECT 6.285 3.350 8.935 3.800 ;
        RECT 9.425 3.570 12.135 3.800 ;
        RECT 9.425 3.460 11.515 3.570 ;
        RECT 5.245 2.685 10.095 2.915 ;
        RECT 5.245 1.315 5.675 2.685 ;
        RECT 9.865 2.575 10.095 2.685 ;
        RECT 6.865 2.345 7.095 2.455 ;
        RECT 11.285 2.345 11.515 3.460 ;
        RECT 11.905 2.875 12.135 3.570 ;
        RECT 12.925 3.500 18.500 3.730 ;
        RECT 6.865 2.115 11.515 2.345 ;
        RECT 6.125 1.885 6.355 2.115 ;
        RECT 6.125 1.655 11.055 1.885 ;
        RECT 10.825 0.910 11.055 1.655 ;
        RECT 11.285 1.315 11.515 2.115 ;
        RECT 12.925 1.655 13.155 3.500 ;
        RECT 13.945 1.655 14.175 3.215 ;
        RECT 12.405 1.315 13.155 1.655 ;
        RECT 13.525 1.540 14.175 1.655 ;
        RECT 15.770 1.540 16.000 3.225 ;
        RECT 17.810 2.115 18.040 3.225 ;
        RECT 18.270 2.425 18.500 3.500 ;
        RECT 20.010 2.115 22.435 2.290 ;
        RECT 17.810 2.060 22.435 2.115 ;
        RECT 16.295 2.005 22.435 2.060 ;
        RECT 16.295 1.830 20.240 2.005 ;
        RECT 13.525 1.310 16.000 1.540 ;
        RECT 18.750 1.775 20.240 1.830 ;
        RECT 18.750 1.315 18.980 1.775 ;
        RECT 10.825 0.680 14.455 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnsnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.160 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 2.330 4.550 2.710 ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.150 2.265 14.975 2.710 ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 1.770 1.530 2.150 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 18.145 1.590 18.375 3.685 ;
        RECT 18.070 0.845 18.375 1.590 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 20.160 5.490 ;
        RECT 1.265 3.425 1.495 4.590 ;
        RECT 3.005 3.905 3.235 4.590 ;
        RECT 7.245 3.905 7.475 4.590 ;
        RECT 9.725 3.905 9.955 4.590 ;
        RECT 13.805 3.915 14.035 4.590 ;
        RECT 16.345 3.175 16.575 4.590 ;
        RECT 19.165 3.875 19.395 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 20.590 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 20.590 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.080 ;
        RECT 3.225 0.450 3.455 1.425 ;
        RECT 7.425 0.450 7.655 1.425 ;
        RECT 16.305 0.450 16.535 1.420 ;
        RECT 19.265 0.450 19.495 1.165 ;
        RECT 0.000 -0.450 20.160 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.105 0.475 3.685 ;
        RECT 2.285 3.675 2.515 3.685 ;
        RECT 5.650 3.675 5.990 4.260 ;
        RECT 11.305 3.675 11.535 4.315 ;
        RECT 14.130 3.685 16.115 3.705 ;
        RECT 2.285 3.445 11.535 3.675 ;
        RECT 11.885 3.475 16.115 3.685 ;
        RECT 11.885 3.455 14.225 3.475 ;
        RECT 0.245 2.875 2.035 3.105 ;
        RECT 1.805 1.540 2.035 2.875 ;
        RECT 0.245 1.310 2.035 1.540 ;
        RECT 0.245 1.170 0.475 1.310 ;
        RECT 2.285 1.170 2.715 3.445 ;
        RECT 3.050 2.985 4.530 3.215 ;
        RECT 3.050 2.100 3.280 2.985 ;
        RECT 3.050 1.870 3.915 2.100 ;
        RECT 3.685 1.655 3.915 1.870 ;
        RECT 5.265 2.060 5.495 3.215 ;
        RECT 8.485 2.700 8.715 3.215 ;
        RECT 10.865 2.700 11.095 3.215 ;
        RECT 6.530 2.470 11.095 2.700 ;
        RECT 5.265 1.830 8.190 2.060 ;
        RECT 3.685 1.315 4.575 1.655 ;
        RECT 5.265 1.315 5.695 1.830 ;
        RECT 9.425 1.315 9.655 2.470 ;
        RECT 11.885 2.005 12.115 3.455 ;
        RECT 15.105 3.215 15.335 3.245 ;
        RECT 13.085 2.985 15.335 3.215 ;
        RECT 13.085 2.875 13.920 2.985 ;
        RECT 15.105 2.905 15.335 2.985 ;
        RECT 10.725 1.775 12.115 2.005 ;
        RECT 10.725 1.315 10.955 1.775 ;
        RECT 13.690 1.545 13.920 2.875 ;
        RECT 15.885 2.730 16.115 3.475 ;
        RECT 15.885 2.500 17.070 2.730 ;
        RECT 17.365 2.315 17.595 3.715 ;
        RECT 17.365 2.270 17.915 2.315 ;
        RECT 15.685 1.975 17.915 2.270 ;
        RECT 15.685 1.930 17.655 1.975 ;
        RECT 11.845 1.205 13.920 1.545 ;
        RECT 17.425 1.315 17.655 1.930 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnsnq_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnsnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.830 1.960 4.890 2.190 ;
        RECT 4.630 1.770 4.890 1.960 ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 13.655 2.165 14.860 2.710 ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.235 1.575 2.710 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.120 0.845 19.450 3.685 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 21.280 5.490 ;
        RECT 1.365 3.425 1.595 4.590 ;
        RECT 3.305 3.580 3.535 4.590 ;
        RECT 7.305 3.110 7.535 4.590 ;
        RECT 9.365 3.110 9.595 4.590 ;
        RECT 13.745 3.970 13.975 4.590 ;
        RECT 16.345 3.210 16.575 4.590 ;
        RECT 18.100 3.875 18.330 4.590 ;
        RECT 20.140 3.875 20.370 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 21.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 21.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.150 0.450 3.490 1.270 ;
        RECT 7.405 0.450 7.635 1.325 ;
        RECT 16.245 0.450 16.475 1.420 ;
        RECT 18.100 0.450 18.330 1.165 ;
        RECT 20.340 0.450 20.570 1.165 ;
        RECT 0.000 -0.450 21.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.765 4.095 7.075 4.325 ;
        RECT 0.345 3.170 0.575 3.710 ;
        RECT 3.765 3.215 3.995 4.095 ;
        RECT 0.345 2.940 2.035 3.170 ;
        RECT 0.345 2.900 0.575 2.940 ;
        RECT 1.805 2.005 2.035 2.940 ;
        RECT 0.245 1.775 2.035 2.005 ;
        RECT 2.385 2.985 3.995 3.215 ;
        RECT 0.245 1.315 0.475 1.775 ;
        RECT 2.385 1.315 2.715 2.985 ;
        RECT 4.325 2.650 4.555 3.750 ;
        RECT 3.370 2.420 4.555 2.650 ;
        RECT 3.370 1.730 3.600 2.420 ;
        RECT 5.445 1.960 5.675 3.750 ;
        RECT 6.845 2.880 7.075 4.095 ;
        RECT 7.765 3.980 9.135 4.210 ;
        RECT 7.765 2.880 7.995 3.980 ;
        RECT 6.845 2.650 7.995 2.880 ;
        RECT 8.325 2.420 8.555 3.750 ;
        RECT 8.905 2.880 9.135 3.980 ;
        RECT 9.825 3.975 11.435 4.315 ;
        RECT 9.825 2.880 10.055 3.975 ;
        RECT 8.905 2.650 10.055 2.880 ;
        RECT 10.765 2.420 10.995 3.685 ;
        RECT 6.810 2.190 10.995 2.420 ;
        RECT 11.785 3.510 16.115 3.740 ;
        RECT 5.445 1.730 8.130 1.960 ;
        RECT 3.370 1.550 3.940 1.730 ;
        RECT 3.370 1.500 4.555 1.550 ;
        RECT 3.715 1.320 4.555 1.500 ;
        RECT 4.325 1.210 4.555 1.320 ;
        RECT 5.445 1.215 5.675 1.730 ;
        RECT 9.365 1.215 9.595 2.190 ;
        RECT 11.785 1.960 12.015 3.510 ;
        RECT 10.665 1.730 12.015 1.960 ;
        RECT 13.025 2.940 15.275 3.280 ;
        RECT 10.665 1.215 10.895 1.730 ;
        RECT 13.025 1.500 13.255 2.940 ;
        RECT 15.885 2.765 16.115 3.510 ;
        RECT 15.885 2.535 17.070 2.765 ;
        RECT 17.365 2.115 17.595 3.750 ;
        RECT 15.625 1.775 18.770 2.115 ;
        RECT 11.785 1.160 13.875 1.500 ;
        RECT 17.365 1.315 17.595 1.775 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnsnq_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnsnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 2.330 4.525 2.710 ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.710 2.150 15.530 2.710 ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.240 1.575 2.710 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.665 3.105 19.895 3.685 ;
        RECT 21.705 3.105 22.135 3.685 ;
        RECT 19.665 2.875 22.135 3.105 ;
        RECT 21.655 1.655 22.135 2.875 ;
        RECT 19.665 1.395 22.135 1.655 ;
        RECT 19.665 0.845 19.895 1.395 ;
        RECT 21.430 0.815 22.135 1.395 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 23.520 5.490 ;
        RECT 1.365 3.425 1.595 4.590 ;
        RECT 3.105 3.860 3.335 4.590 ;
        RECT 7.345 3.905 7.575 4.590 ;
        RECT 9.825 3.905 10.055 4.590 ;
        RECT 14.205 3.915 14.435 4.590 ;
        RECT 16.745 3.155 16.975 4.590 ;
        RECT 18.645 3.875 18.875 4.590 ;
        RECT 20.685 3.875 20.915 4.590 ;
        RECT 22.725 3.875 22.955 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 23.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 23.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.225 0.450 3.455 1.425 ;
        RECT 7.525 0.450 7.755 1.425 ;
        RECT 16.525 0.450 16.755 1.425 ;
        RECT 18.545 0.450 18.775 1.165 ;
        RECT 20.785 0.450 21.015 1.165 ;
        RECT 23.025 0.450 23.255 1.165 ;
        RECT 0.000 -0.450 23.520 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 3.170 0.575 3.750 ;
        RECT 5.805 3.720 6.035 4.360 ;
        RECT 2.385 3.630 2.615 3.685 ;
        RECT 3.520 3.675 6.035 3.720 ;
        RECT 11.565 3.675 11.795 4.315 ;
        RECT 3.520 3.630 11.795 3.675 ;
        RECT 2.385 3.490 11.795 3.630 ;
        RECT 2.385 3.400 3.705 3.490 ;
        RECT 5.895 3.445 11.795 3.490 ;
        RECT 12.145 3.455 16.515 3.685 ;
        RECT 0.345 2.940 2.035 3.170 ;
        RECT 1.805 1.685 2.035 2.940 ;
        RECT 0.245 1.455 2.035 1.685 ;
        RECT 0.245 1.315 0.475 1.455 ;
        RECT 2.385 1.315 2.715 3.400 ;
        RECT 4.290 3.170 4.630 3.205 ;
        RECT 3.050 2.940 4.630 3.170 ;
        RECT 3.050 2.100 3.280 2.940 ;
        RECT 3.050 1.870 4.575 2.100 ;
        RECT 4.345 1.315 4.575 1.870 ;
        RECT 5.365 2.060 5.595 3.260 ;
        RECT 8.585 2.745 8.815 3.215 ;
        RECT 11.125 2.745 11.355 3.215 ;
        RECT 6.630 2.515 11.355 2.745 ;
        RECT 5.365 1.830 8.290 2.060 ;
        RECT 5.365 1.315 5.795 1.830 ;
        RECT 9.825 1.315 10.055 2.515 ;
        RECT 12.145 2.005 12.375 3.455 ;
        RECT 13.485 2.995 15.790 3.225 ;
        RECT 13.485 2.875 14.335 2.995 ;
        RECT 11.125 1.775 12.375 2.005 ;
        RECT 11.125 1.315 11.355 1.775 ;
        RECT 14.105 1.545 14.335 2.875 ;
        RECT 16.285 2.710 16.515 3.455 ;
        RECT 16.285 2.480 17.470 2.710 ;
        RECT 17.765 2.320 17.995 3.695 ;
        RECT 17.765 2.115 21.425 2.320 ;
        RECT 16.085 1.960 21.425 2.115 ;
        RECT 16.085 1.775 18.055 1.960 ;
        RECT 12.245 1.205 14.335 1.545 ;
        RECT 17.825 1.315 18.055 1.775 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnsnq_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.680 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.630 1.210 4.890 2.115 ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.235 1.575 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.710 2.330 15.115 3.685 ;
        RECT 14.885 0.845 15.115 2.330 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 15.680 5.490 ;
        RECT 1.365 3.895 1.595 4.590 ;
        RECT 3.185 3.905 3.415 4.590 ;
        RECT 7.205 3.045 7.435 4.590 ;
        RECT 12.025 3.145 12.255 4.590 ;
        RECT 13.765 3.875 13.995 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 16.110 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 16.110 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.205 0.450 3.435 1.435 ;
        RECT 7.295 0.450 7.525 0.625 ;
        RECT 11.925 0.450 12.155 1.265 ;
        RECT 13.765 0.450 13.995 1.165 ;
        RECT 0.000 -0.450 15.680 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 3.655 0.575 4.235 ;
        RECT 5.885 3.675 6.115 4.315 ;
        RECT 1.940 3.655 6.115 3.675 ;
        RECT 0.345 3.445 6.115 3.655 ;
        RECT 0.345 3.425 2.035 3.445 ;
        RECT 1.805 2.005 2.035 3.425 ;
        RECT 2.385 2.755 2.615 3.215 ;
        RECT 5.165 2.755 5.395 3.215 ;
        RECT 2.385 2.525 4.075 2.755 ;
        RECT 0.245 1.775 2.035 2.005 ;
        RECT 3.845 1.895 4.075 2.525 ;
        RECT 0.245 1.315 0.475 1.775 ;
        RECT 2.485 1.665 4.075 1.895 ;
        RECT 2.485 1.315 2.715 1.665 ;
        RECT 3.845 0.920 4.075 1.665 ;
        RECT 5.165 2.415 7.875 2.755 ;
        RECT 5.165 1.315 5.395 2.415 ;
        RECT 8.225 2.115 8.455 3.685 ;
        RECT 6.685 1.775 8.455 2.115 ;
        RECT 8.225 1.655 8.455 1.775 ;
        RECT 9.745 3.455 11.795 3.685 ;
        RECT 8.225 1.315 8.855 1.655 ;
        RECT 9.745 1.315 9.975 3.455 ;
        RECT 10.505 1.085 10.735 2.755 ;
        RECT 11.565 2.700 11.795 3.455 ;
        RECT 11.565 2.470 12.750 2.700 ;
        RECT 13.045 2.115 13.275 3.685 ;
        RECT 11.265 2.060 13.275 2.115 ;
        RECT 11.265 1.830 14.490 2.060 ;
        RECT 11.265 1.775 13.275 1.830 ;
        RECT 13.045 1.315 13.275 1.775 ;
        RECT 5.665 0.920 10.735 1.085 ;
        RECT 3.845 0.855 10.735 0.920 ;
        RECT 3.845 0.690 5.890 0.855 ;
        RECT 9.010 0.690 10.735 0.855 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffq_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.800 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.630 1.210 5.080 2.050 ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 1.770 1.490 2.150 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.995 1.590 15.325 3.685 ;
        RECT 14.710 1.210 15.325 1.590 ;
        RECT 15.095 0.845 15.325 1.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 16.800 5.490 ;
        RECT 1.210 3.950 1.550 4.590 ;
        RECT 3.395 3.885 3.625 4.590 ;
        RECT 7.235 3.090 7.465 4.590 ;
        RECT 12.235 3.875 12.465 4.590 ;
        RECT 13.975 3.875 14.205 4.590 ;
        RECT 16.015 3.875 16.245 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 17.230 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 17.230 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.665 1.595 1.080 ;
        RECT 1.365 0.450 3.425 0.665 ;
        RECT 7.555 0.450 7.785 0.545 ;
        RECT 12.135 0.450 12.365 1.160 ;
        RECT 13.975 0.450 14.205 1.165 ;
        RECT 16.215 0.450 16.445 1.165 ;
        RECT 0.000 -0.450 16.800 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.675 0.475 4.235 ;
        RECT 3.855 4.020 6.145 4.360 ;
        RECT 0.245 3.655 3.300 3.675 ;
        RECT 3.855 3.655 4.085 4.020 ;
        RECT 0.245 3.445 4.085 3.655 ;
        RECT 0.245 3.425 2.035 3.445 ;
        RECT 3.205 3.425 4.085 3.445 ;
        RECT 1.805 1.540 2.035 3.425 ;
        RECT 0.245 1.310 2.035 1.540 ;
        RECT 2.385 2.800 2.615 3.215 ;
        RECT 5.375 2.800 5.605 3.730 ;
        RECT 2.385 2.570 4.285 2.800 ;
        RECT 0.245 1.170 0.475 1.310 ;
        RECT 2.385 1.170 2.715 2.570 ;
        RECT 4.055 0.980 4.285 2.570 ;
        RECT 5.375 2.460 8.085 2.800 ;
        RECT 5.375 1.305 5.605 2.460 ;
        RECT 8.835 2.105 9.065 3.730 ;
        RECT 6.655 1.765 9.065 2.105 ;
        RECT 8.835 1.310 9.065 1.765 ;
        RECT 9.955 3.500 12.055 3.730 ;
        RECT 9.955 1.310 10.185 3.500 ;
        RECT 10.715 1.005 10.945 2.800 ;
        RECT 11.825 2.700 12.055 3.500 ;
        RECT 11.825 2.470 12.960 2.700 ;
        RECT 13.255 2.110 13.485 3.685 ;
        RECT 11.475 2.060 13.485 2.110 ;
        RECT 11.475 1.830 14.700 2.060 ;
        RECT 11.475 1.770 13.485 1.830 ;
        RECT 5.995 0.980 10.945 1.005 ;
        RECT 4.055 0.775 10.945 0.980 ;
        RECT 13.255 0.840 13.485 1.770 ;
        RECT 4.055 0.680 6.100 0.775 ;
        RECT 9.220 0.685 10.945 0.775 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffq_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.630 1.210 4.890 2.115 ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.235 1.505 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 15.125 3.105 15.355 3.685 ;
        RECT 17.165 3.105 17.770 3.685 ;
        RECT 15.125 2.875 17.770 3.105 ;
        RECT 17.115 1.655 17.770 2.875 ;
        RECT 15.285 1.395 17.770 1.655 ;
        RECT 15.285 0.845 15.515 1.395 ;
        RECT 17.510 0.815 17.770 1.395 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 19.600 5.490 ;
        RECT 1.310 3.950 1.650 4.590 ;
        RECT 3.185 3.905 3.415 4.590 ;
        RECT 7.125 3.045 7.355 4.590 ;
        RECT 12.065 3.875 12.295 4.590 ;
        RECT 14.105 3.875 14.335 4.590 ;
        RECT 16.145 3.875 16.375 4.590 ;
        RECT 18.185 3.875 18.415 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 20.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 20.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.205 0.450 3.435 1.435 ;
        RECT 7.290 0.450 7.520 0.625 ;
        RECT 11.925 0.450 12.155 1.165 ;
        RECT 14.165 0.450 14.395 1.165 ;
        RECT 16.405 0.450 16.635 1.165 ;
        RECT 18.645 0.450 18.875 1.165 ;
        RECT 0.000 -0.450 19.600 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 3.675 0.575 4.235 ;
        RECT 5.805 3.675 6.035 4.315 ;
        RECT 0.345 3.445 6.035 3.675 ;
        RECT 0.345 3.425 2.035 3.445 ;
        RECT 1.805 2.005 2.035 3.425 ;
        RECT 2.385 2.755 2.615 3.215 ;
        RECT 5.165 2.755 5.395 3.215 ;
        RECT 2.385 2.525 4.075 2.755 ;
        RECT 0.245 1.775 2.035 2.005 ;
        RECT 3.845 1.895 4.075 2.525 ;
        RECT 0.245 1.315 0.475 1.775 ;
        RECT 2.485 1.665 4.075 1.895 ;
        RECT 2.485 1.315 2.715 1.665 ;
        RECT 3.845 0.920 4.075 1.665 ;
        RECT 5.165 2.415 8.175 2.755 ;
        RECT 5.165 1.315 5.395 2.415 ;
        RECT 8.620 2.115 8.855 3.685 ;
        RECT 6.685 1.775 8.855 2.115 ;
        RECT 8.625 1.315 8.855 1.775 ;
        RECT 9.745 3.455 11.935 3.685 ;
        RECT 9.745 1.315 9.975 3.455 ;
        RECT 10.625 1.085 10.855 2.755 ;
        RECT 11.705 2.700 11.935 3.455 ;
        RECT 11.705 2.470 12.790 2.700 ;
        RECT 13.085 2.315 13.315 3.685 ;
        RECT 13.085 2.115 16.885 2.315 ;
        RECT 11.265 1.975 16.885 2.115 ;
        RECT 11.265 1.775 13.310 1.975 ;
        RECT 5.665 0.920 10.855 1.085 ;
        RECT 3.845 0.855 10.855 0.920 ;
        RECT 3.845 0.690 5.890 0.855 ;
        RECT 9.010 0.690 10.855 0.855 ;
        RECT 13.045 0.845 13.310 1.775 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffq_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.920 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.280 2.330 3.915 2.710 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.830000 ;
    PORT
      LAYER Metal1 ;
        RECT 13.865 1.660 14.380 2.000 ;
        RECT 14.150 1.590 14.380 1.660 ;
        RECT 14.150 1.210 15.070 1.590 ;
    END
  END RN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.660 2.150 0.970 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 16.345 2.190 16.650 3.685 ;
        RECT 16.325 0.845 16.650 2.190 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.920 5.490 ;
        RECT 1.285 3.425 1.515 4.590 ;
        RECT 3.245 3.615 3.475 4.590 ;
        RECT 7.325 3.615 7.555 4.590 ;
        RECT 9.065 3.330 9.295 4.590 ;
        RECT 13.365 4.190 13.595 4.590 ;
        RECT 15.625 3.310 15.855 4.590 ;
        RECT 17.365 3.875 17.595 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 18.350 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 18.350 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.385 0.450 1.615 1.225 ;
        RECT 3.225 0.450 3.455 1.200 ;
        RECT 8.705 0.450 8.935 1.200 ;
        RECT 13.185 0.450 13.415 1.200 ;
        RECT 17.445 0.450 17.675 1.165 ;
        RECT 0.000 -0.450 17.920 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.705 4.130 4.990 4.360 ;
        RECT 0.265 3.170 0.495 3.685 ;
        RECT 2.305 3.385 2.535 3.685 ;
        RECT 3.705 3.385 3.935 4.130 ;
        RECT 0.265 2.940 1.430 3.170 ;
        RECT 0.265 2.875 0.495 2.940 ;
        RECT 1.200 2.260 1.430 2.940 ;
        RECT 2.305 3.155 3.935 3.385 ;
        RECT 1.200 2.030 2.010 2.260 ;
        RECT 1.200 1.685 1.430 2.030 ;
        RECT 0.210 1.455 1.430 1.685 ;
        RECT 0.210 1.370 1.085 1.455 ;
        RECT 2.305 1.315 2.735 3.155 ;
        RECT 4.265 1.200 4.575 3.785 ;
        RECT 5.285 2.915 5.515 3.785 ;
        RECT 6.305 3.375 6.535 3.955 ;
        RECT 8.345 3.375 8.575 3.955 ;
        RECT 6.305 3.145 8.575 3.375 ;
        RECT 5.285 2.685 9.790 2.915 ;
        RECT 5.285 1.540 5.520 2.685 ;
        RECT 10.085 2.460 10.315 3.970 ;
        RECT 9.855 2.405 10.315 2.460 ;
        RECT 6.830 2.230 10.315 2.405 ;
        RECT 10.945 3.960 11.335 3.970 ;
        RECT 10.945 3.730 15.295 3.960 ;
        RECT 10.945 3.160 11.335 3.730 ;
        RECT 6.830 2.175 10.055 2.230 ;
        RECT 5.850 1.715 9.595 1.945 ;
        RECT 5.285 1.200 5.695 1.540 ;
        RECT 9.365 0.970 9.595 1.715 ;
        RECT 9.825 1.200 10.055 2.175 ;
        RECT 10.285 0.970 10.515 2.000 ;
        RECT 10.945 1.200 11.175 3.160 ;
        RECT 11.485 0.970 11.830 2.985 ;
        RECT 12.065 1.200 12.355 3.500 ;
        RECT 14.605 2.650 14.835 3.500 ;
        RECT 15.065 2.700 15.295 3.730 ;
        RECT 12.650 2.470 14.835 2.650 ;
        RECT 12.650 2.240 16.100 2.470 ;
        RECT 15.605 1.290 15.835 2.240 ;
        RECT 9.365 0.740 11.830 0.970 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffrnq_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffrnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.040 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.960 2.330 3.895 2.710 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.255000 ;
    PORT
      LAYER Metal1 ;
        RECT 13.590 2.330 14.015 2.710 ;
    END
  END RN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.265 1.590 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.601600 ;
    PORT
      LAYER Metal1 ;
        RECT 17.445 0.845 17.770 3.685 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 19.040 5.490 ;
        RECT 1.365 3.425 1.595 4.590 ;
        RECT 3.225 3.615 3.455 4.590 ;
        RECT 7.305 3.615 7.535 4.590 ;
        RECT 9.045 3.320 9.275 4.590 ;
        RECT 13.345 4.345 13.575 4.590 ;
        RECT 15.385 3.875 15.615 4.590 ;
        RECT 16.425 3.875 16.655 4.590 ;
        RECT 18.465 3.875 18.695 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 19.470 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 19.470 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.200 ;
        RECT 3.205 0.450 3.435 1.195 ;
        RECT 8.425 0.450 8.655 1.195 ;
        RECT 13.135 0.450 13.365 1.195 ;
        RECT 16.325 0.450 16.555 1.235 ;
        RECT 18.565 0.450 18.795 1.235 ;
        RECT 0.000 -0.450 19.040 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.685 4.130 4.970 4.360 ;
        RECT 0.345 3.195 0.575 3.735 ;
        RECT 2.385 3.385 2.615 3.685 ;
        RECT 3.685 3.385 3.915 4.130 ;
        RECT 0.345 2.965 2.090 3.195 ;
        RECT 0.345 2.925 0.575 2.965 ;
        RECT 1.860 2.035 2.090 2.965 ;
        RECT 0.245 1.805 2.090 2.035 ;
        RECT 2.385 3.155 3.915 3.385 ;
        RECT 0.245 1.290 0.475 1.805 ;
        RECT 2.385 1.290 2.715 3.155 ;
        RECT 4.245 1.195 4.555 3.785 ;
        RECT 5.265 2.915 5.495 3.785 ;
        RECT 6.285 3.375 6.515 3.955 ;
        RECT 8.325 3.375 8.555 3.955 ;
        RECT 6.285 3.145 8.555 3.375 ;
        RECT 5.265 2.685 9.770 2.915 ;
        RECT 5.265 1.525 5.495 2.685 ;
        RECT 10.065 2.455 10.295 3.960 ;
        RECT 6.810 2.225 10.295 2.455 ;
        RECT 10.895 3.730 15.155 3.960 ;
        RECT 5.855 1.710 9.535 1.940 ;
        RECT 5.265 1.185 5.675 1.525 ;
        RECT 9.305 0.965 9.535 1.710 ;
        RECT 9.765 1.195 9.995 2.225 ;
        RECT 10.225 0.965 10.455 1.995 ;
        RECT 10.895 1.195 11.315 3.730 ;
        RECT 11.555 2.690 11.815 3.030 ;
        RECT 11.555 0.965 11.785 2.690 ;
        RECT 12.105 1.535 12.335 3.490 ;
        RECT 12.630 2.940 14.695 3.170 ;
        RECT 12.630 2.745 12.970 2.940 ;
        RECT 14.465 2.185 14.695 2.940 ;
        RECT 14.925 2.415 15.155 3.730 ;
        RECT 14.465 1.955 17.050 2.185 ;
        RECT 12.015 1.195 12.335 1.535 ;
        RECT 15.555 1.830 17.050 1.955 ;
        RECT 9.305 0.735 11.785 0.965 ;
        RECT 15.555 0.725 15.785 1.830 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffrnq_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffrnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.890 1.750 3.895 2.090 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.123000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.970 1.750 13.780 2.090 ;
    END
  END RN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.330 1.570 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 17.370 3.215 17.605 3.685 ;
        RECT 19.410 3.215 19.840 3.685 ;
        RECT 17.370 2.875 19.840 3.215 ;
        RECT 19.595 1.625 19.840 2.875 ;
        RECT 17.370 1.395 19.840 1.625 ;
        RECT 17.370 0.815 17.600 1.395 ;
        RECT 19.610 0.815 19.840 1.395 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 21.280 5.490 ;
        RECT 1.365 3.425 1.595 4.590 ;
        RECT 3.105 3.090 3.335 4.590 ;
        RECT 7.185 3.560 7.415 4.590 ;
        RECT 8.925 3.390 9.155 4.590 ;
        RECT 13.330 4.345 13.560 4.590 ;
        RECT 15.370 3.875 15.605 4.590 ;
        RECT 16.345 3.875 16.580 4.590 ;
        RECT 18.390 4.585 20.660 4.590 ;
        RECT 18.390 3.875 18.620 4.585 ;
        RECT 20.430 3.875 20.660 4.585 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 21.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 21.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.225 0.450 3.455 1.370 ;
        RECT 8.305 0.450 8.535 1.370 ;
        RECT 13.110 0.640 13.340 1.370 ;
        RECT 13.110 0.450 16.535 0.640 ;
        RECT 18.490 0.450 18.720 1.165 ;
        RECT 20.730 0.450 20.960 1.165 ;
        RECT 0.000 -0.450 21.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.665 4.020 4.795 4.360 ;
        RECT 0.345 3.170 0.575 3.750 ;
        RECT 0.345 2.940 2.035 3.170 ;
        RECT 1.805 1.685 2.035 2.940 ;
        RECT 0.245 1.455 2.035 1.685 ;
        RECT 2.385 2.860 2.615 3.685 ;
        RECT 3.665 2.860 3.895 4.020 ;
        RECT 2.385 2.630 3.895 2.860 ;
        RECT 2.385 1.600 2.615 2.630 ;
        RECT 0.245 1.315 0.475 1.455 ;
        RECT 2.385 1.260 2.715 1.600 ;
        RECT 4.125 1.260 4.575 3.730 ;
        RECT 5.145 2.860 5.375 3.730 ;
        RECT 6.165 3.320 6.395 3.900 ;
        RECT 8.205 3.320 8.435 3.900 ;
        RECT 6.165 3.090 8.435 3.320 ;
        RECT 5.145 2.630 9.650 2.860 ;
        RECT 5.145 1.600 5.375 2.630 ;
        RECT 9.995 2.430 10.225 4.030 ;
        RECT 9.765 2.290 10.225 2.430 ;
        RECT 6.690 2.200 10.225 2.290 ;
        RECT 10.870 3.800 15.060 4.030 ;
        RECT 10.870 3.220 11.245 3.800 ;
        RECT 6.690 2.060 9.980 2.200 ;
        RECT 6.145 1.830 6.375 2.060 ;
        RECT 6.145 1.600 9.520 1.830 ;
        RECT 5.145 1.260 5.695 1.600 ;
        RECT 9.290 1.030 9.520 1.600 ;
        RECT 9.750 1.260 9.980 2.060 ;
        RECT 10.410 1.030 10.640 2.060 ;
        RECT 10.870 1.260 11.100 3.220 ;
        RECT 11.455 1.030 11.685 3.100 ;
        RECT 11.990 1.260 12.265 3.560 ;
        RECT 12.670 2.760 14.580 3.215 ;
        RECT 14.350 2.185 14.580 2.760 ;
        RECT 14.830 2.415 15.060 3.800 ;
        RECT 14.350 1.955 19.365 2.185 ;
        RECT 15.530 1.315 15.760 1.955 ;
        RECT 9.290 0.800 11.685 1.030 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffrnq_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffrsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffrsnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.720 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.965 2.545 3.770 2.710 ;
        RECT 2.965 2.315 4.010 2.545 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018000 ;
    PORT
      LAYER Metal1 ;
        RECT 16.300 2.330 17.210 2.890 ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.710 2.890 15.055 3.270 ;
        RECT 14.825 2.470 15.055 2.890 ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.480 1.580 3.270 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.125 0.845 19.450 3.685 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 20.720 5.490 ;
        RECT 1.265 3.960 1.495 4.590 ;
        RECT 3.005 3.560 3.235 4.590 ;
        RECT 7.245 4.490 7.475 4.590 ;
        RECT 10.445 4.490 10.675 4.590 ;
        RECT 14.330 4.005 14.670 4.590 ;
        RECT 16.370 4.005 16.710 4.590 ;
        RECT 18.465 3.480 18.695 4.590 ;
        RECT 20.205 3.875 20.435 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 21.150 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 21.150 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.385 0.450 1.615 1.225 ;
        RECT 3.285 0.450 3.515 1.425 ;
        RECT 8.585 0.450 8.815 1.425 ;
        RECT 16.360 0.450 16.590 1.225 ;
        RECT 20.245 0.450 20.475 1.165 ;
        RECT 0.000 -0.450 20.720 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.465 4.020 4.835 4.360 ;
        RECT 5.570 4.260 5.910 4.305 ;
        RECT 5.570 4.030 12.490 4.260 ;
        RECT 0.245 3.500 2.055 3.730 ;
        RECT 0.245 3.390 0.475 3.500 ;
        RECT 1.825 1.740 2.055 3.500 ;
        RECT 0.265 1.510 2.055 1.740 ;
        RECT 2.285 3.330 2.515 3.750 ;
        RECT 3.465 3.330 3.695 4.020 ;
        RECT 2.285 3.100 3.695 3.330 ;
        RECT 0.265 1.315 0.495 1.510 ;
        RECT 2.285 1.315 2.735 3.100 ;
        RECT 4.025 3.005 4.255 3.730 ;
        RECT 4.025 2.775 4.635 3.005 ;
        RECT 4.405 1.315 4.635 2.775 ;
        RECT 5.045 2.915 5.275 3.730 ;
        RECT 6.065 3.350 8.715 3.800 ;
        RECT 9.205 3.570 11.855 3.800 ;
        RECT 9.205 3.460 9.955 3.570 ;
        RECT 5.045 2.685 9.495 2.915 ;
        RECT 5.525 1.315 5.755 2.685 ;
        RECT 9.265 2.575 9.495 2.685 ;
        RECT 6.805 2.345 7.035 2.455 ;
        RECT 9.725 2.345 9.955 3.460 ;
        RECT 11.625 2.875 11.855 3.570 ;
        RECT 12.645 3.545 18.135 3.775 ;
        RECT 12.645 3.195 12.875 3.545 ;
        RECT 12.085 2.965 12.875 3.195 ;
        RECT 12.085 2.645 12.315 2.965 ;
        RECT 13.665 2.735 13.895 3.215 ;
        RECT 11.665 2.415 12.315 2.645 ;
        RECT 12.785 2.505 14.495 2.735 ;
        RECT 6.805 2.115 10.775 2.345 ;
        RECT 5.985 1.885 6.215 2.115 ;
        RECT 5.985 1.655 10.315 1.885 ;
        RECT 10.085 0.910 10.315 1.655 ;
        RECT 10.545 1.315 10.775 2.115 ;
        RECT 11.665 1.315 11.895 2.415 ;
        RECT 12.785 1.315 13.015 2.505 ;
        RECT 13.295 0.910 13.525 2.275 ;
        RECT 14.265 2.240 14.495 2.505 ;
        RECT 15.405 2.240 15.635 3.270 ;
        RECT 14.265 2.010 15.635 2.240 ;
        RECT 17.445 2.060 17.675 3.270 ;
        RECT 17.905 2.470 18.135 3.545 ;
        RECT 18.320 2.060 18.895 2.315 ;
        RECT 14.265 1.315 14.630 2.010 ;
        RECT 15.865 1.975 18.895 2.060 ;
        RECT 15.865 1.830 18.550 1.975 ;
        RECT 18.320 1.315 18.550 1.830 ;
        RECT 10.085 0.680 13.525 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffrsnq_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffrsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffrsnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.840 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.945 2.500 3.770 2.710 ;
        RECT 2.945 2.270 4.010 2.500 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018000 ;
    PORT
      LAYER Metal1 ;
        RECT 16.040 2.330 17.275 2.710 ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.220 1.770 15.115 2.150 ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.685 2.200 1.575 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 20.245 0.845 20.570 3.685 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 21.840 5.490 ;
        RECT 1.265 3.425 1.495 4.590 ;
        RECT 3.005 3.515 3.235 4.590 ;
        RECT 7.305 4.490 7.535 4.590 ;
        RECT 10.505 4.490 10.735 4.590 ;
        RECT 14.390 3.950 14.730 4.590 ;
        RECT 16.430 3.950 16.770 4.590 ;
        RECT 18.525 3.425 18.755 4.590 ;
        RECT 19.245 3.875 19.475 4.590 ;
        RECT 21.285 3.875 21.515 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 22.270 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 22.270 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.285 0.450 3.515 1.425 ;
        RECT 8.645 0.450 8.875 1.425 ;
        RECT 16.405 0.450 16.635 1.225 ;
        RECT 19.125 0.450 19.355 1.165 ;
        RECT 21.365 0.450 21.595 1.165 ;
        RECT 0.000 -0.450 21.840 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.465 3.975 4.835 4.315 ;
        RECT 5.570 4.030 12.550 4.260 ;
        RECT 0.245 3.170 0.475 3.750 ;
        RECT 2.285 3.285 2.515 3.685 ;
        RECT 3.465 3.285 3.695 3.975 ;
        RECT 0.245 2.940 2.035 3.170 ;
        RECT 1.805 1.740 2.035 2.940 ;
        RECT 0.245 1.510 2.035 1.740 ;
        RECT 2.285 3.055 3.695 3.285 ;
        RECT 0.245 1.315 0.475 1.510 ;
        RECT 2.285 1.315 2.715 3.055 ;
        RECT 4.025 2.960 4.255 3.685 ;
        RECT 5.045 3.105 5.275 3.685 ;
        RECT 6.065 3.350 8.775 3.800 ;
        RECT 9.265 3.570 11.915 3.800 ;
        RECT 9.265 3.460 10.835 3.570 ;
        RECT 4.025 2.730 4.635 2.960 ;
        RECT 5.045 2.875 9.555 3.105 ;
        RECT 4.405 1.315 4.635 2.730 ;
        RECT 5.525 1.315 5.755 2.875 ;
        RECT 9.325 2.575 9.555 2.875 ;
        RECT 6.805 2.345 7.035 2.455 ;
        RECT 10.605 2.345 10.835 3.460 ;
        RECT 11.685 2.875 11.915 3.570 ;
        RECT 12.705 3.455 18.195 3.685 ;
        RECT 6.805 2.115 10.835 2.345 ;
        RECT 5.985 1.885 6.215 2.115 ;
        RECT 5.985 1.655 10.375 1.885 ;
        RECT 10.145 0.910 10.375 1.655 ;
        RECT 10.605 1.315 10.835 2.115 ;
        RECT 12.705 2.110 12.935 3.455 ;
        RECT 11.725 1.880 12.935 2.110 ;
        RECT 11.725 1.315 11.955 1.880 ;
        RECT 13.725 1.650 13.955 3.215 ;
        RECT 12.845 1.540 13.955 1.650 ;
        RECT 15.450 2.875 15.695 3.215 ;
        RECT 15.450 1.540 15.680 2.875 ;
        RECT 17.505 2.115 17.735 3.215 ;
        RECT 17.965 2.415 18.195 3.455 ;
        RECT 17.505 2.100 19.795 2.115 ;
        RECT 15.910 1.870 19.795 2.100 ;
        RECT 12.845 1.200 15.680 1.540 ;
        RECT 18.365 1.775 19.795 1.870 ;
        RECT 18.365 1.315 18.595 1.775 ;
        RECT 10.145 0.680 13.790 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffrsnq_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffrsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffrsnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 24.080 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.945 2.500 3.770 2.710 ;
        RECT 2.945 2.270 4.010 2.500 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018000 ;
    PORT
      LAYER Metal1 ;
        RECT 16.185 2.330 17.275 2.710 ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.260 1.770 15.115 2.150 ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.685 2.200 1.575 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 20.205 3.105 20.495 3.685 ;
        RECT 22.305 3.105 22.885 3.685 ;
        RECT 20.205 2.875 22.885 3.105 ;
        RECT 22.300 1.655 22.885 2.875 ;
        RECT 20.205 1.395 22.885 1.655 ;
        RECT 20.205 0.845 20.435 1.395 ;
        RECT 22.445 0.845 22.885 1.395 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 24.080 5.490 ;
        RECT 1.265 3.425 1.495 4.590 ;
        RECT 3.005 3.515 3.235 4.590 ;
        RECT 7.305 4.490 7.535 4.590 ;
        RECT 10.505 4.490 10.735 4.590 ;
        RECT 14.390 3.950 14.730 4.590 ;
        RECT 16.430 3.950 16.770 4.590 ;
        RECT 18.525 3.425 18.755 4.590 ;
        RECT 19.245 3.875 19.475 4.590 ;
        RECT 21.285 3.875 21.515 4.590 ;
        RECT 23.325 3.875 23.555 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 24.510 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 24.510 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.285 0.450 3.515 1.425 ;
        RECT 8.645 0.450 8.875 1.425 ;
        RECT 16.405 0.450 16.635 1.225 ;
        RECT 19.085 0.450 19.315 1.165 ;
        RECT 21.325 0.450 21.555 1.165 ;
        RECT 23.565 0.450 23.795 1.165 ;
        RECT 0.000 -0.450 24.080 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.465 3.975 4.835 4.315 ;
        RECT 5.570 4.030 12.550 4.260 ;
        RECT 0.245 3.170 0.475 3.750 ;
        RECT 2.285 3.285 2.515 3.685 ;
        RECT 3.465 3.285 3.695 3.975 ;
        RECT 0.245 2.940 2.035 3.170 ;
        RECT 1.805 1.740 2.035 2.940 ;
        RECT 0.245 1.510 2.035 1.740 ;
        RECT 2.285 3.055 3.695 3.285 ;
        RECT 0.245 1.315 0.475 1.510 ;
        RECT 2.285 1.315 2.715 3.055 ;
        RECT 4.025 2.960 4.255 3.685 ;
        RECT 5.045 3.105 5.275 3.685 ;
        RECT 6.065 3.350 8.775 3.800 ;
        RECT 9.265 3.570 11.915 3.800 ;
        RECT 9.265 3.460 10.835 3.570 ;
        RECT 4.025 2.730 4.635 2.960 ;
        RECT 5.045 2.875 9.555 3.105 ;
        RECT 4.405 1.315 4.635 2.730 ;
        RECT 5.525 1.315 5.755 2.875 ;
        RECT 9.325 2.575 9.555 2.875 ;
        RECT 6.805 2.345 7.035 2.455 ;
        RECT 10.605 2.345 10.835 3.460 ;
        RECT 11.685 2.875 11.915 3.570 ;
        RECT 12.705 3.455 18.195 3.685 ;
        RECT 6.805 2.115 10.835 2.345 ;
        RECT 5.985 1.885 6.215 2.115 ;
        RECT 5.985 1.655 10.375 1.885 ;
        RECT 10.145 0.910 10.375 1.655 ;
        RECT 10.605 1.315 10.835 2.115 ;
        RECT 12.705 2.110 12.935 3.455 ;
        RECT 11.725 1.880 12.935 2.110 ;
        RECT 11.725 1.315 11.955 1.880 ;
        RECT 13.725 1.650 13.955 3.215 ;
        RECT 12.845 1.540 13.955 1.650 ;
        RECT 15.450 2.875 15.695 3.215 ;
        RECT 15.450 1.540 15.680 2.875 ;
        RECT 17.505 2.115 17.735 3.215 ;
        RECT 17.965 2.415 18.195 3.455 ;
        RECT 19.520 2.115 22.070 2.315 ;
        RECT 17.505 2.100 22.070 2.115 ;
        RECT 15.910 1.975 22.070 2.100 ;
        RECT 15.910 1.870 19.755 1.975 ;
        RECT 12.845 1.200 15.680 1.540 ;
        RECT 18.365 1.865 19.755 1.870 ;
        RECT 18.365 1.315 18.595 1.865 ;
        RECT 10.145 0.680 13.790 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffrsnq_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffsnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.160 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 1.770 4.030 2.150 ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.970 1.830 14.655 2.170 ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.330 1.530 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.190 0.845 19.450 3.685 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 20.160 5.490 ;
        RECT 1.365 3.425 1.595 4.590 ;
        RECT 3.305 3.145 3.535 4.590 ;
        RECT 7.525 3.960 7.755 4.590 ;
        RECT 10.005 4.005 10.235 4.590 ;
        RECT 13.985 3.145 14.215 4.590 ;
        RECT 16.025 3.615 16.255 4.590 ;
        RECT 18.185 3.875 18.415 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 20.590 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 20.590 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.205 0.450 3.435 1.245 ;
        RECT 7.405 0.450 7.635 1.245 ;
        RECT 16.245 0.450 16.475 1.265 ;
        RECT 18.085 0.450 18.315 1.165 ;
        RECT 0.000 -0.450 20.160 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.765 4.130 5.150 4.360 ;
        RECT 0.345 3.170 0.575 3.750 ;
        RECT 0.345 2.940 2.035 3.170 ;
        RECT 1.805 2.005 2.035 2.940 ;
        RECT 0.245 1.775 2.035 2.005 ;
        RECT 2.385 2.915 2.615 3.685 ;
        RECT 3.765 2.915 3.995 4.130 ;
        RECT 2.385 2.685 3.995 2.915 ;
        RECT 0.245 1.315 0.475 1.775 ;
        RECT 2.385 1.315 2.715 2.685 ;
        RECT 4.325 1.135 4.555 3.785 ;
        RECT 5.445 2.340 5.675 3.785 ;
        RECT 5.970 3.730 6.310 4.360 ;
        RECT 11.345 3.775 11.575 4.315 ;
        RECT 7.895 3.730 11.575 3.775 ;
        RECT 5.970 3.545 11.575 3.730 ;
        RECT 5.970 3.500 8.035 3.545 ;
        RECT 8.765 2.975 11.135 3.315 ;
        RECT 8.765 2.800 10.015 2.975 ;
        RECT 6.810 2.570 10.015 2.800 ;
        RECT 5.445 2.110 8.470 2.340 ;
        RECT 5.445 1.135 5.675 2.110 ;
        RECT 6.070 1.650 8.095 1.880 ;
        RECT 7.865 0.910 8.095 1.650 ;
        RECT 9.785 1.315 10.015 2.570 ;
        RECT 11.925 2.115 12.155 3.685 ;
        RECT 13.265 2.915 13.495 3.685 ;
        RECT 15.005 2.915 15.235 3.785 ;
        RECT 13.265 2.685 15.235 2.915 ;
        RECT 15.585 2.730 17.455 3.215 ;
        RECT 13.265 2.630 13.495 2.685 ;
        RECT 10.905 1.885 12.155 2.115 ;
        RECT 12.510 2.400 13.495 2.630 ;
        RECT 15.585 2.515 18.855 2.730 ;
        RECT 10.905 1.030 11.135 1.885 ;
        RECT 12.510 1.655 12.740 2.400 ;
        RECT 17.365 2.390 18.855 2.515 ;
        RECT 12.025 1.600 12.740 1.655 ;
        RECT 14.885 1.830 16.970 2.060 ;
        RECT 12.025 1.260 14.215 1.600 ;
        RECT 14.885 1.030 15.115 1.830 ;
        RECT 17.365 1.315 17.595 2.390 ;
        RECT 7.865 0.680 10.510 0.910 ;
        RECT 10.905 0.800 15.115 1.030 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffsnq_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.720 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.075 1.770 3.975 2.150 ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.435 1.590 14.665 2.115 ;
        RECT 14.435 1.210 14.970 1.590 ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.240 1.390 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.125 0.845 19.450 3.685 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 20.720 5.490 ;
        RECT 1.365 3.895 1.595 4.590 ;
        RECT 3.305 3.615 3.535 4.590 ;
        RECT 7.475 3.615 7.705 4.590 ;
        RECT 9.875 3.830 10.105 4.590 ;
        RECT 13.855 3.515 14.085 4.590 ;
        RECT 15.895 3.045 16.125 4.590 ;
        RECT 18.105 3.875 18.335 4.590 ;
        RECT 20.145 3.875 20.375 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 21.150 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 21.150 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.205 0.450 3.435 1.320 ;
        RECT 7.475 0.450 7.705 1.320 ;
        RECT 16.115 0.450 16.345 1.165 ;
        RECT 18.005 0.450 18.235 1.165 ;
        RECT 20.245 0.450 20.475 1.165 ;
        RECT 0.000 -0.450 20.720 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.765 4.130 5.295 4.360 ;
        RECT 0.345 3.010 2.035 3.240 ;
        RECT 3.765 3.215 3.995 4.130 ;
        RECT 0.345 2.900 0.575 3.010 ;
        RECT 1.805 1.740 2.035 3.010 ;
        RECT 0.245 1.510 2.035 1.740 ;
        RECT 2.385 2.985 3.995 3.215 ;
        RECT 0.245 1.315 0.475 1.510 ;
        RECT 2.385 1.315 2.715 2.985 ;
        RECT 4.325 1.210 4.555 3.785 ;
        RECT 5.445 2.415 5.820 3.785 ;
        RECT 6.115 3.385 6.455 4.360 ;
        RECT 7.935 3.600 9.650 3.775 ;
        RECT 11.215 3.675 11.445 4.315 ;
        RECT 10.275 3.600 11.445 3.675 ;
        RECT 7.935 3.545 11.445 3.600 ;
        RECT 7.935 3.385 8.165 3.545 ;
        RECT 6.115 3.155 8.165 3.385 ;
        RECT 9.425 3.445 11.445 3.545 ;
        RECT 9.425 3.370 10.445 3.445 ;
        RECT 8.575 2.800 8.805 3.315 ;
        RECT 10.775 2.800 11.005 3.215 ;
        RECT 6.980 2.570 11.005 2.800 ;
        RECT 5.445 2.340 6.810 2.415 ;
        RECT 5.445 2.185 8.420 2.340 ;
        RECT 5.445 1.210 5.675 2.185 ;
        RECT 6.640 2.110 8.420 2.185 ;
        RECT 6.130 1.880 6.470 1.955 ;
        RECT 6.130 1.650 8.165 1.880 ;
        RECT 7.935 0.910 8.165 1.650 ;
        RECT 9.655 1.315 9.885 2.570 ;
        RECT 11.795 2.115 12.025 3.685 ;
        RECT 14.875 3.215 15.105 3.795 ;
        RECT 11.435 1.885 12.025 2.115 ;
        RECT 13.135 2.985 15.105 3.215 ;
        RECT 10.775 0.980 11.005 1.425 ;
        RECT 11.435 0.980 11.665 1.885 ;
        RECT 13.135 1.655 13.365 2.985 ;
        RECT 17.135 2.630 17.445 3.685 ;
        RECT 15.455 2.290 17.445 2.630 ;
        RECT 17.215 2.115 17.445 2.290 ;
        RECT 11.895 1.550 13.365 1.655 ;
        RECT 15.200 1.830 16.840 2.060 ;
        RECT 11.895 1.210 14.165 1.550 ;
        RECT 15.200 0.980 15.430 1.830 ;
        RECT 7.935 0.680 10.380 0.910 ;
        RECT 10.775 0.750 15.430 0.980 ;
        RECT 17.215 1.775 18.775 2.115 ;
        RECT 17.215 0.845 17.465 1.775 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffsnq_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffsnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.945 2.330 4.030 2.710 ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 13.530 2.220 14.515 2.710 ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.240 1.570 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.110 3.105 19.340 3.685 ;
        RECT 21.150 3.105 21.880 3.685 ;
        RECT 19.110 2.875 21.880 3.105 ;
        RECT 21.590 1.655 21.880 2.875 ;
        RECT 19.405 1.395 21.880 1.655 ;
        RECT 19.405 0.845 19.640 1.395 ;
        RECT 21.590 0.845 21.880 1.395 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 23.520 5.490 ;
        RECT 1.365 3.425 1.595 4.590 ;
        RECT 3.305 3.615 3.535 4.590 ;
        RECT 7.510 3.615 7.740 4.590 ;
        RECT 9.715 3.885 10.055 4.590 ;
        RECT 13.790 3.515 14.020 4.590 ;
        RECT 15.830 3.045 16.060 4.590 ;
        RECT 18.090 3.875 18.320 4.590 ;
        RECT 20.130 3.875 20.360 4.590 ;
        RECT 22.170 3.875 22.400 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 23.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 23.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.205 0.450 3.435 1.425 ;
        RECT 7.455 0.450 7.795 1.370 ;
        RECT 15.995 0.450 16.335 0.640 ;
        RECT 18.290 0.450 18.520 1.165 ;
        RECT 20.530 0.450 20.760 1.165 ;
        RECT 22.770 0.450 23.000 1.165 ;
        RECT 0.000 -0.450 23.520 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.765 4.130 5.295 4.360 ;
        RECT 0.345 3.170 0.575 3.750 ;
        RECT 2.385 3.385 2.615 3.685 ;
        RECT 3.765 3.385 3.995 4.130 ;
        RECT 0.345 2.940 2.090 3.170 ;
        RECT 1.860 1.685 2.090 2.940 ;
        RECT 0.245 1.455 2.090 1.685 ;
        RECT 2.385 3.155 3.995 3.385 ;
        RECT 0.245 1.315 0.475 1.455 ;
        RECT 2.385 1.315 2.715 3.155 ;
        RECT 4.325 1.315 4.555 3.785 ;
        RECT 5.445 2.520 5.820 3.785 ;
        RECT 6.115 3.385 6.455 4.360 ;
        RECT 7.970 3.655 9.545 3.720 ;
        RECT 11.150 3.655 11.380 4.315 ;
        RECT 7.970 3.490 11.380 3.655 ;
        RECT 7.970 3.385 8.200 3.490 ;
        RECT 9.320 3.425 11.380 3.490 ;
        RECT 6.115 3.155 8.200 3.385 ;
        RECT 8.475 2.800 8.815 3.260 ;
        RECT 10.655 2.800 10.995 3.160 ;
        RECT 7.015 2.570 10.995 2.800 ;
        RECT 5.445 2.340 6.790 2.520 ;
        RECT 5.445 2.290 8.235 2.340 ;
        RECT 5.445 1.315 5.675 2.290 ;
        RECT 6.565 2.110 8.235 2.290 ;
        RECT 6.000 1.880 6.340 2.060 ;
        RECT 6.000 1.650 9.320 1.880 ;
        RECT 9.090 0.910 9.320 1.650 ;
        RECT 9.550 1.315 9.780 2.570 ;
        RECT 11.730 2.115 11.960 3.685 ;
        RECT 14.810 3.215 15.040 3.685 ;
        RECT 11.370 1.885 11.960 2.115 ;
        RECT 13.070 2.985 15.040 3.215 ;
        RECT 11.370 1.425 11.600 1.885 ;
        RECT 13.070 1.655 13.300 2.985 ;
        RECT 14.810 2.875 15.040 2.985 ;
        RECT 17.070 2.520 17.305 3.685 ;
        RECT 15.250 2.325 17.305 2.520 ;
        RECT 15.250 2.290 20.920 2.325 ;
        RECT 15.250 2.180 15.480 2.290 ;
        RECT 15.680 1.830 16.775 2.060 ;
        RECT 17.075 2.030 20.920 2.290 ;
        RECT 10.710 1.085 11.600 1.425 ;
        RECT 11.830 1.315 14.100 1.655 ;
        RECT 15.680 1.085 15.910 1.830 ;
        RECT 9.090 0.680 10.315 0.910 ;
        RECT 10.710 0.855 15.910 1.085 ;
        RECT 17.075 0.845 17.400 2.030 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffsnq_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dlya_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlya_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.160 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 1.770 1.045 2.495 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.130 4.070 5.865 4.330 ;
        RECT 5.535 0.845 5.865 4.070 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 6.160 5.490 ;
        RECT 1.265 3.240 1.495 4.590 ;
        RECT 4.125 3.240 4.355 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.590 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.590 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.620 ;
        RECT 4.515 0.450 4.745 0.695 ;
        RECT 0.000 -0.450 6.160 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.955 0.475 3.580 ;
        RECT 0.245 2.725 2.035 2.955 ;
        RECT 0.245 1.280 0.475 2.725 ;
        RECT 1.805 1.740 2.035 2.725 ;
        RECT 2.385 2.495 2.615 3.580 ;
        RECT 3.105 3.010 3.335 3.580 ;
        RECT 3.105 2.780 4.290 3.010 ;
        RECT 4.060 2.585 4.290 2.780 ;
        RECT 2.385 1.795 3.830 2.495 ;
        RECT 2.385 1.280 2.715 1.795 ;
        RECT 4.060 1.745 5.185 2.585 ;
        RECT 4.055 1.695 5.185 1.745 ;
        RECT 4.055 0.910 4.285 1.695 ;
        RECT 3.000 0.680 4.285 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlya_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dlya_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlya_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.210 0.970 2.795 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.821000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.130 3.265 5.615 4.330 ;
        RECT 5.130 3.035 6.435 3.265 ;
        RECT 6.205 1.990 6.435 3.035 ;
        RECT 5.485 1.760 6.435 1.990 ;
        RECT 5.485 0.845 5.715 1.760 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.280 5.490 ;
        RECT 1.265 3.485 1.495 4.590 ;
        RECT 4.130 3.485 4.360 4.590 ;
        RECT 6.505 3.485 6.735 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 7.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.645 ;
        RECT 4.365 0.450 4.595 0.960 ;
        RECT 6.625 0.450 6.855 1.630 ;
        RECT 0.000 -0.450 7.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.255 0.475 3.825 ;
        RECT 0.245 3.025 2.035 3.255 ;
        RECT 0.245 1.305 0.475 3.025 ;
        RECT 1.805 1.985 2.035 3.025 ;
        RECT 2.385 2.270 2.615 3.825 ;
        RECT 3.110 3.255 3.340 3.825 ;
        RECT 3.110 3.025 4.295 3.255 ;
        RECT 3.550 2.270 3.835 2.795 ;
        RECT 2.385 2.040 3.835 2.270 ;
        RECT 4.065 2.560 4.295 3.025 ;
        RECT 4.065 2.220 5.975 2.560 ;
        RECT 2.385 1.305 2.715 2.040 ;
        RECT 4.065 1.410 4.295 2.220 ;
        RECT 2.955 1.180 4.295 1.410 ;
        RECT 2.955 0.680 3.295 1.180 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlya_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dlya_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlya_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.035 1.050 2.735 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.642000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.680 3.210 5.910 4.250 ;
        RECT 7.820 3.210 8.050 4.250 ;
        RECT 5.680 2.980 8.050 3.210 ;
        RECT 5.680 2.950 7.575 2.980 ;
        RECT 7.345 2.040 7.575 2.950 ;
        RECT 5.630 1.810 8.100 2.040 ;
        RECT 5.630 0.770 5.860 1.810 ;
        RECT 7.870 0.770 8.100 1.810 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 9.520 5.490 ;
        RECT 1.270 3.440 1.500 4.590 ;
        RECT 4.280 3.440 4.510 4.590 ;
        RECT 6.700 3.440 6.930 4.590 ;
        RECT 8.890 3.440 9.120 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 9.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.370 0.450 1.600 1.110 ;
        RECT 4.330 0.450 4.560 1.110 ;
        RECT 6.750 0.450 6.980 1.580 ;
        RECT 8.990 0.450 9.220 1.580 ;
        RECT 0.000 -0.450 9.520 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.250 3.195 0.480 3.780 ;
        RECT 0.250 2.965 2.095 3.195 ;
        RECT 0.250 0.770 0.480 2.965 ;
        RECT 1.755 2.035 2.095 2.965 ;
        RECT 2.390 2.735 2.620 3.780 ;
        RECT 3.260 3.210 3.490 3.780 ;
        RECT 3.260 2.980 4.445 3.210 ;
        RECT 2.390 2.505 3.985 2.735 ;
        RECT 3.700 2.030 3.985 2.505 ;
        RECT 2.490 1.800 3.985 2.030 ;
        RECT 4.215 2.500 4.445 2.980 ;
        RECT 4.215 2.270 7.115 2.500 ;
        RECT 2.490 0.770 2.720 1.800 ;
        RECT 4.215 1.570 4.445 2.270 ;
        RECT 3.210 1.340 4.445 1.570 ;
        RECT 3.210 0.770 3.440 1.340 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlya_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dlyb_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyb_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 1.770 0.990 2.560 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.535 3.270 6.865 4.340 ;
        RECT 5.190 2.890 6.865 3.270 ;
        RECT 6.635 0.680 6.865 2.890 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.280 5.490 ;
        RECT 1.265 4.020 1.495 4.590 ;
        RECT 4.735 4.040 4.965 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.295 7.710 5.470 ;
        RECT -0.430 2.265 0.430 2.295 ;
        RECT 5.300 2.265 7.710 2.295 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 0.430 2.265 5.300 2.295 ;
        RECT -0.430 -0.430 7.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 0.965 ;
        RECT 4.835 0.450 5.065 0.695 ;
        RECT 0.000 -0.450 7.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.190 3.020 0.475 4.360 ;
        RECT 1.555 3.300 2.740 3.640 ;
        RECT 0.190 2.790 2.280 3.020 ;
        RECT 0.190 0.910 0.420 2.790 ;
        RECT 1.940 1.860 2.280 2.790 ;
        RECT 2.510 1.630 2.740 3.300 ;
        RECT 4.730 3.320 4.965 3.660 ;
        RECT 4.155 1.630 4.385 2.615 ;
        RECT 1.500 1.400 4.385 1.630 ;
        RECT 4.730 2.090 4.960 3.320 ;
        RECT 5.900 2.090 6.240 2.560 ;
        RECT 4.730 1.860 6.240 2.090 ;
        RECT 4.730 1.075 5.065 1.860 ;
        RECT 0.190 0.680 0.530 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyb_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dlyb_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyb_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.400 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 1.770 0.990 2.560 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.912500 ;
    PORT
      LAYER Metal1 ;
        RECT 6.635 3.270 6.865 4.360 ;
        RECT 6.310 2.890 6.865 3.270 ;
        RECT 6.635 0.680 6.865 2.890 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 8.400 5.490 ;
        RECT 1.265 3.915 1.495 4.590 ;
        RECT 4.735 3.915 4.965 4.590 ;
        RECT 7.705 3.880 7.935 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.295 8.830 5.470 ;
        RECT -0.430 2.265 0.430 2.295 ;
        RECT 5.315 2.265 8.830 2.295 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 0.430 2.265 5.315 2.295 ;
        RECT -0.430 -0.430 8.830 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 0.965 ;
        RECT 4.835 0.450 5.065 0.695 ;
        RECT 7.755 0.450 7.985 1.435 ;
        RECT 0.000 -0.450 8.400 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.190 3.020 0.475 4.255 ;
        RECT 1.500 3.250 2.740 3.480 ;
        RECT 0.190 2.790 2.280 3.020 ;
        RECT 0.190 0.910 0.420 2.790 ;
        RECT 1.940 1.860 2.280 2.790 ;
        RECT 2.510 2.035 2.740 3.250 ;
        RECT 4.155 2.035 4.385 2.615 ;
        RECT 2.510 1.805 4.385 2.035 ;
        RECT 4.735 2.325 4.965 3.535 ;
        RECT 4.735 2.095 6.380 2.325 ;
        RECT 2.510 1.630 2.740 1.805 ;
        RECT 1.500 1.400 2.740 1.630 ;
        RECT 4.735 1.075 5.065 2.095 ;
        RECT 0.190 0.680 0.530 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyb_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dlyb_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyb_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.640 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.900 0.970 2.710 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.825000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.740 3.650 6.970 4.360 ;
        RECT 8.930 3.650 9.160 4.360 ;
        RECT 6.740 3.420 9.160 3.650 ;
        RECT 8.930 1.590 9.160 3.420 ;
        RECT 6.690 1.210 9.160 1.590 ;
        RECT 6.690 0.680 6.920 1.210 ;
        RECT 8.930 0.680 9.160 1.210 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 10.640 5.490 ;
        RECT 1.320 4.060 1.550 4.590 ;
        RECT 4.790 4.060 5.020 4.590 ;
        RECT 7.760 3.880 7.990 4.590 ;
        RECT 9.950 3.880 10.180 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.295 11.070 5.470 ;
        RECT -0.430 2.265 0.430 2.295 ;
        RECT 5.370 2.265 11.070 2.295 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 0.430 2.265 5.370 2.295 ;
        RECT -0.430 -0.430 11.070 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.420 0.450 1.650 0.965 ;
        RECT 4.890 0.450 5.120 0.695 ;
        RECT 7.810 0.450 8.040 0.965 ;
        RECT 10.050 0.450 10.280 1.435 ;
        RECT 0.000 -0.450 10.640 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.170 0.585 4.345 ;
        RECT 1.555 3.395 2.795 3.625 ;
        RECT 0.245 2.940 1.505 3.170 ;
        RECT 0.245 0.910 0.475 2.940 ;
        RECT 1.275 2.655 1.505 2.940 ;
        RECT 1.275 2.425 2.335 2.655 ;
        RECT 2.050 1.900 2.335 2.425 ;
        RECT 2.565 1.630 2.795 3.395 ;
        RECT 4.210 1.630 4.440 2.710 ;
        RECT 1.555 1.400 4.440 1.630 ;
        RECT 4.790 2.420 5.020 3.680 ;
        RECT 4.790 2.190 8.175 2.420 ;
        RECT 4.790 1.075 5.120 2.190 ;
        RECT 0.245 0.680 0.585 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyb_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dlyc_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyc_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.200 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 1.770 0.970 2.560 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.590 3.270 10.920 4.360 ;
        RECT 10.230 2.890 10.920 3.270 ;
        RECT 10.690 0.680 10.920 2.890 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 11.200 5.490 ;
        RECT 1.610 4.220 1.840 4.590 ;
        RECT 1.610 3.880 9.020 4.220 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.295 11.630 5.470 ;
        RECT -0.430 2.265 0.430 2.295 ;
        RECT 9.355 2.265 11.630 2.295 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 0.430 2.265 9.355 2.295 ;
        RECT -0.430 -0.430 11.630 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 0.965 ;
        RECT 4.890 0.450 5.120 0.690 ;
        RECT 8.890 0.450 9.120 0.695 ;
        RECT 0.000 -0.450 11.200 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.170 3.020 0.475 4.220 ;
        RECT 1.555 3.215 4.440 3.445 ;
        RECT 0.170 2.790 1.430 3.020 ;
        RECT 0.170 0.910 0.400 2.790 ;
        RECT 1.200 2.560 1.430 2.790 ;
        RECT 1.200 2.330 2.335 2.560 ;
        RECT 1.995 1.860 2.335 2.330 ;
        RECT 4.210 1.630 4.440 3.215 ;
        RECT 1.555 1.400 4.440 1.630 ;
        RECT 4.790 2.090 5.020 3.500 ;
        RECT 5.610 3.020 5.840 3.500 ;
        RECT 5.610 2.790 6.795 3.020 ;
        RECT 5.995 2.090 6.335 2.560 ;
        RECT 4.790 1.860 6.335 2.090 ;
        RECT 4.790 1.070 5.120 1.860 ;
        RECT 6.565 1.630 6.795 2.790 ;
        RECT 8.210 1.630 8.440 2.615 ;
        RECT 5.610 1.400 8.440 1.630 ;
        RECT 8.790 2.090 9.020 3.500 ;
        RECT 9.955 2.090 10.295 2.560 ;
        RECT 8.790 1.860 10.295 2.090 ;
        RECT 5.610 1.070 5.840 1.400 ;
        RECT 8.790 1.075 9.120 1.860 ;
        RECT 0.170 0.680 0.530 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyc_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dlyc_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyc_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.320 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 1.770 0.990 2.560 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.912500 ;
    PORT
      LAYER Metal1 ;
        RECT 10.635 1.590 10.865 4.360 ;
        RECT 10.230 1.210 10.865 1.590 ;
        RECT 10.635 0.680 10.865 1.210 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 12.320 5.490 ;
        RECT 1.265 3.915 1.495 4.590 ;
        RECT 4.735 3.915 4.965 4.590 ;
        RECT 8.735 3.915 8.965 4.590 ;
        RECT 11.705 3.880 11.935 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.295 12.750 5.470 ;
        RECT -0.430 2.265 0.430 2.295 ;
        RECT 9.315 2.265 12.750 2.295 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 0.430 2.265 9.315 2.295 ;
        RECT -0.430 -0.430 12.750 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 0.965 ;
        RECT 4.835 0.450 5.065 0.690 ;
        RECT 8.835 0.450 9.065 0.695 ;
        RECT 11.755 0.450 11.985 1.435 ;
        RECT 0.000 -0.450 12.320 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.190 3.020 0.475 4.255 ;
        RECT 1.500 3.250 2.740 3.480 ;
        RECT 0.190 2.790 2.280 3.020 ;
        RECT 0.190 0.910 0.420 2.790 ;
        RECT 1.940 1.860 2.280 2.790 ;
        RECT 2.510 1.630 2.740 3.250 ;
        RECT 4.155 1.630 4.385 2.615 ;
        RECT 1.500 1.400 4.385 1.630 ;
        RECT 4.735 2.090 4.965 3.535 ;
        RECT 5.555 3.020 5.785 3.535 ;
        RECT 5.555 2.790 6.740 3.020 ;
        RECT 5.940 2.090 6.280 2.560 ;
        RECT 4.735 1.860 6.280 2.090 ;
        RECT 4.735 1.070 5.065 1.860 ;
        RECT 6.510 1.630 6.740 2.790 ;
        RECT 8.155 1.630 8.385 2.615 ;
        RECT 5.555 1.400 8.385 1.630 ;
        RECT 8.735 2.325 8.965 3.535 ;
        RECT 8.735 2.095 10.380 2.325 ;
        RECT 5.555 1.070 5.785 1.400 ;
        RECT 8.735 1.075 9.065 2.095 ;
        RECT 0.190 0.680 0.530 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyc_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dlyc_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyc_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.560 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 1.140 0.990 1.840 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.642000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.565 3.105 10.795 3.685 ;
        RECT 12.705 3.105 12.935 3.685 ;
        RECT 10.565 2.875 12.935 3.105 ;
        RECT 12.225 1.655 12.455 2.875 ;
        RECT 10.565 1.425 13.035 1.655 ;
        RECT 10.565 0.845 10.795 1.425 ;
        RECT 12.470 0.845 13.035 1.425 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 14.560 5.490 ;
        RECT 1.265 3.710 1.495 4.590 ;
        RECT 4.665 3.710 4.895 4.590 ;
        RECT 8.665 3.710 8.895 4.590 ;
        RECT 11.585 3.875 11.815 4.590 ;
        RECT 13.825 3.875 14.055 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.380 14.990 5.470 ;
        RECT -0.430 2.265 0.430 2.380 ;
        RECT 9.065 2.265 14.990 2.380 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 0.430 2.265 9.065 2.380 ;
        RECT -0.430 -0.430 14.990 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 0.965 ;
        RECT 4.765 0.450 4.995 0.935 ;
        RECT 8.765 0.450 8.995 0.935 ;
        RECT 11.685 0.450 11.915 1.165 ;
        RECT 13.925 0.450 14.155 1.165 ;
        RECT 0.000 -0.450 14.560 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.190 2.760 0.475 4.050 ;
        RECT 1.485 2.990 4.315 3.330 ;
        RECT 0.190 2.530 2.210 2.760 ;
        RECT 0.190 0.910 0.420 2.530 ;
        RECT 1.870 2.060 2.210 2.530 ;
        RECT 4.085 1.715 4.315 2.990 ;
        RECT 1.430 1.485 4.315 1.715 ;
        RECT 4.665 2.060 4.895 3.330 ;
        RECT 5.485 2.990 5.715 3.330 ;
        RECT 5.485 2.760 8.315 2.990 ;
        RECT 5.870 2.060 6.210 2.530 ;
        RECT 4.665 1.830 6.210 2.060 ;
        RECT 4.665 1.315 4.995 1.830 ;
        RECT 8.085 1.600 8.315 2.760 ;
        RECT 5.430 1.370 8.315 1.600 ;
        RECT 8.665 2.315 8.895 3.330 ;
        RECT 8.665 1.975 11.995 2.315 ;
        RECT 8.665 1.315 8.995 1.975 ;
        RECT 0.190 0.680 0.530 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyc_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dlyd_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyd_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.120 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 0.970 2.580 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.545 0.840 14.970 4.360 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 15.120 5.490 ;
        RECT 1.270 3.895 1.500 4.590 ;
        RECT 4.740 3.895 4.970 4.590 ;
        RECT 8.740 3.895 8.970 4.590 ;
        RECT 12.745 3.895 12.975 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.295 15.550 5.470 ;
        RECT -0.430 2.265 0.430 2.295 ;
        RECT 13.310 2.265 15.550 2.295 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 0.430 2.265 13.310 2.295 ;
        RECT -0.430 -0.430 15.550 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.370 0.450 1.600 0.965 ;
        RECT 4.840 0.450 5.070 0.930 ;
        RECT 8.840 0.450 9.070 0.930 ;
        RECT 12.845 0.450 13.075 0.690 ;
        RECT 0.000 -0.450 15.120 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.195 3.040 0.480 4.235 ;
        RECT 1.505 3.230 2.690 3.460 ;
        RECT 0.195 3.000 1.375 3.040 ;
        RECT 0.195 2.810 2.230 3.000 ;
        RECT 0.195 0.910 0.425 2.810 ;
        RECT 1.245 2.770 2.230 2.810 ;
        RECT 2.000 2.190 2.230 2.770 ;
        RECT 2.460 1.630 2.690 3.230 ;
        RECT 4.740 2.580 4.970 3.515 ;
        RECT 5.560 3.040 5.790 3.515 ;
        RECT 5.560 2.810 6.690 3.040 ;
        RECT 4.160 1.630 4.390 2.580 ;
        RECT 1.505 1.400 4.390 1.630 ;
        RECT 4.740 2.350 6.230 2.580 ;
        RECT 4.740 1.310 5.070 2.350 ;
        RECT 6.000 1.770 6.230 2.350 ;
        RECT 5.505 1.540 5.845 1.595 ;
        RECT 6.460 1.540 6.690 2.810 ;
        RECT 8.740 2.580 8.970 3.515 ;
        RECT 9.560 3.040 9.790 3.515 ;
        RECT 9.560 2.810 10.690 3.040 ;
        RECT 8.160 1.540 8.390 2.580 ;
        RECT 5.505 1.310 8.390 1.540 ;
        RECT 8.740 2.350 10.230 2.580 ;
        RECT 8.740 1.310 9.070 2.350 ;
        RECT 10.000 1.770 10.230 2.350 ;
        RECT 9.505 1.540 9.845 1.595 ;
        RECT 10.460 1.540 10.690 2.810 ;
        RECT 12.165 1.540 12.395 2.580 ;
        RECT 9.505 1.310 12.395 1.540 ;
        RECT 12.745 2.000 12.975 3.515 ;
        RECT 13.965 2.000 14.195 2.580 ;
        RECT 12.745 1.770 14.195 2.000 ;
        RECT 12.745 1.070 13.075 1.770 ;
        RECT 0.195 0.680 0.535 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyd_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dlyd_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyd_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.240 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 1.770 0.990 2.570 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.821000 ;
    PORT
      LAYER Metal1 ;
        RECT 13.530 4.070 14.765 4.360 ;
        RECT 14.535 3.365 14.765 4.070 ;
        RECT 14.535 3.135 15.585 3.365 ;
        RECT 15.355 1.820 15.585 3.135 ;
        RECT 14.635 1.590 15.585 1.820 ;
        RECT 14.635 0.845 14.865 1.590 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 16.240 5.490 ;
        RECT 1.265 3.925 1.495 4.590 ;
        RECT 4.735 3.925 4.965 4.590 ;
        RECT 8.735 3.925 8.965 4.590 ;
        RECT 12.735 3.925 12.965 4.590 ;
        RECT 15.655 3.585 15.885 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.295 16.670 5.470 ;
        RECT -0.430 2.265 0.430 2.295 ;
        RECT 13.315 2.265 16.670 2.295 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 0.430 2.265 13.315 2.295 ;
        RECT -0.430 -0.430 16.670 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 0.965 ;
        RECT 4.835 0.450 5.065 0.690 ;
        RECT 8.835 0.450 9.065 0.920 ;
        RECT 12.835 0.450 13.065 0.695 ;
        RECT 15.755 0.450 15.985 1.435 ;
        RECT 0.000 -0.450 16.240 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.190 3.030 0.475 4.265 ;
        RECT 1.500 3.260 4.385 3.490 ;
        RECT 0.190 2.800 2.225 3.030 ;
        RECT 0.190 0.910 0.420 2.800 ;
        RECT 1.995 2.220 2.225 2.800 ;
        RECT 4.155 1.630 4.385 3.260 ;
        RECT 1.500 1.400 4.385 1.630 ;
        RECT 4.735 2.625 4.965 3.545 ;
        RECT 5.555 3.085 5.785 3.545 ;
        RECT 5.555 2.855 8.385 3.085 ;
        RECT 4.735 1.815 6.225 2.625 ;
        RECT 4.735 1.070 5.065 1.815 ;
        RECT 8.155 1.585 8.385 2.855 ;
        RECT 5.555 1.355 8.385 1.585 ;
        RECT 8.735 2.625 8.965 3.545 ;
        RECT 9.555 3.085 9.785 3.545 ;
        RECT 9.555 2.855 12.385 3.085 ;
        RECT 8.735 1.815 10.225 2.625 ;
        RECT 5.555 1.070 5.785 1.355 ;
        RECT 8.735 1.300 9.065 1.815 ;
        RECT 12.155 1.585 12.385 2.855 ;
        RECT 9.500 1.355 12.385 1.585 ;
        RECT 12.735 2.390 12.965 3.545 ;
        RECT 12.735 2.050 15.125 2.390 ;
        RECT 12.735 1.075 13.065 2.050 ;
        RECT 0.190 0.680 0.530 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyd_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dlyd_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyd_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.480 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.660 1.770 1.000 2.595 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.825000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.695 3.120 14.970 4.360 ;
        RECT 16.735 3.120 16.965 4.360 ;
        RECT 14.695 2.890 16.965 3.120 ;
        RECT 16.360 1.900 16.590 2.890 ;
        RECT 14.645 1.670 17.115 1.900 ;
        RECT 14.645 0.680 14.875 1.670 ;
        RECT 16.885 0.680 17.115 1.670 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 18.480 5.490 ;
        RECT 1.275 3.930 1.505 4.590 ;
        RECT 4.745 3.930 4.975 4.590 ;
        RECT 8.745 3.930 8.975 4.590 ;
        RECT 12.745 3.930 12.975 4.590 ;
        RECT 15.715 3.880 15.945 4.590 ;
        RECT 17.905 3.880 18.135 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.300 18.910 5.470 ;
        RECT -0.430 2.265 0.430 2.300 ;
        RECT 13.310 2.265 18.910 2.300 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 0.430 2.265 13.310 2.300 ;
        RECT -0.430 -0.430 18.910 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.375 0.450 1.605 0.970 ;
        RECT 4.845 0.450 5.075 0.970 ;
        RECT 8.845 0.450 9.075 0.965 ;
        RECT 12.845 0.450 13.075 0.695 ;
        RECT 15.765 0.450 15.995 1.440 ;
        RECT 18.005 0.450 18.235 1.440 ;
        RECT 0.000 -0.450 18.480 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.200 3.055 0.485 4.270 ;
        RECT 1.510 3.265 2.750 3.495 ;
        RECT 0.200 3.035 1.415 3.055 ;
        RECT 0.200 2.825 2.290 3.035 ;
        RECT 0.200 0.915 0.430 2.825 ;
        RECT 1.320 2.805 2.290 2.825 ;
        RECT 1.950 1.895 2.290 2.805 ;
        RECT 2.520 1.635 2.750 3.265 ;
        RECT 4.165 1.635 4.395 2.650 ;
        RECT 1.510 1.405 4.395 1.635 ;
        RECT 4.745 2.125 4.975 3.550 ;
        RECT 5.565 3.055 5.795 3.550 ;
        RECT 5.565 2.825 6.750 3.055 ;
        RECT 5.950 2.125 6.290 2.595 ;
        RECT 4.745 1.895 6.290 2.125 ;
        RECT 4.745 1.350 5.075 1.895 ;
        RECT 6.520 1.635 6.750 2.825 ;
        RECT 8.165 1.635 8.395 2.650 ;
        RECT 5.510 1.405 8.395 1.635 ;
        RECT 8.745 2.125 8.975 3.550 ;
        RECT 9.565 3.055 9.795 3.550 ;
        RECT 9.565 2.825 10.750 3.055 ;
        RECT 9.950 2.125 10.290 2.595 ;
        RECT 8.745 1.895 10.290 2.125 ;
        RECT 10.520 2.070 10.750 2.825 ;
        RECT 12.165 2.070 12.395 2.650 ;
        RECT 8.745 1.345 9.075 1.895 ;
        RECT 10.520 1.840 12.395 2.070 ;
        RECT 12.745 2.360 12.975 3.550 ;
        RECT 12.745 2.130 16.130 2.360 ;
        RECT 10.520 1.630 10.750 1.840 ;
        RECT 9.510 1.400 10.750 1.630 ;
        RECT 12.745 1.075 13.075 2.130 ;
        RECT 0.200 0.685 0.540 0.915 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyd_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__endcap
  CLASS ENDCAP PRE ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__endcap ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.120 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Nwell ;
        RECT -2.930 2.265 1.550 5.470 ;
      LAYER Metal1 ;
        RECT 0.000 4.590 1.120 5.490 ;
        RECT 0.230 2.340 0.850 4.590 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Pwell ;
        RECT -2.930 -0.430 1.550 2.265 ;
      LAYER Metal1 ;
        RECT 0.230 0.450 0.850 1.530 ;
        RECT 0.000 -0.450 1.120 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__endcap

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__fill_1
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fill_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.560 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 0.560 5.490 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 0.990 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 0.990 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.450 0.560 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__fill_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__fill_2
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fill_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.120 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 1.120 5.490 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 1.550 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 1.550 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.450 1.120 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__fill_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__fill_4
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fill_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.240 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 2.240 5.490 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 2.670 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 2.670 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.450 2.240 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__fill_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__fill_8
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fill_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 4.480 5.490 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 4.910 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.450 4.480 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__fill_8

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__fill_16
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fill_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.960 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 8.960 5.490 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 9.390 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.390 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.450 8.960 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__fill_16

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__fill_32
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fill_32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.920 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.920 5.490 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 18.350 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 18.350 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.450 17.920 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__fill_32

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__fill_64
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fill_64 ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.840 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 35.840 5.490 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 36.270 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 36.270 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.450 35.840 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__fill_64

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__fillcap_4
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fillcap_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.240 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 2.240 5.490 ;
        RECT 1.765 3.550 1.995 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 2.670 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 2.670 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 0.000 -0.450 2.240 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.060 0.475 4.360 ;
        RECT 1.270 2.470 1.995 2.700 ;
        RECT 0.245 1.830 0.970 2.060 ;
        RECT 1.765 0.680 1.995 2.470 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__fillcap_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__fillcap_8
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fillcap_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 4.480 5.490 ;
        RECT 1.765 3.550 1.995 4.590 ;
        RECT 4.005 3.550 4.235 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 4.910 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 0.000 -0.450 4.480 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.060 0.475 4.360 ;
        RECT 1.270 2.470 1.995 2.700 ;
        RECT 0.245 1.830 0.970 2.060 ;
        RECT 1.765 0.680 1.995 2.470 ;
        RECT 2.485 2.060 2.715 4.360 ;
        RECT 3.510 2.470 4.235 2.700 ;
        RECT 2.485 1.830 3.210 2.060 ;
        RECT 4.005 0.680 4.235 2.470 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__fillcap_8

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__fillcap_16
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fillcap_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.960 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 8.960 5.490 ;
        RECT 1.765 3.550 1.995 4.590 ;
        RECT 4.005 3.550 4.235 4.590 ;
        RECT 6.245 3.550 6.475 4.590 ;
        RECT 8.485 3.550 8.715 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 9.390 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.390 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 4.725 0.450 4.955 1.490 ;
        RECT 6.965 0.450 7.195 1.490 ;
        RECT 0.000 -0.450 8.960 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.060 0.475 4.360 ;
        RECT 1.270 2.470 1.995 2.700 ;
        RECT 0.245 1.830 0.970 2.060 ;
        RECT 1.765 0.680 1.995 2.470 ;
        RECT 2.485 2.060 2.715 4.360 ;
        RECT 3.510 2.470 4.235 2.700 ;
        RECT 2.485 1.830 3.210 2.060 ;
        RECT 4.005 0.680 4.235 2.470 ;
        RECT 4.725 2.060 4.955 4.360 ;
        RECT 5.750 2.470 6.475 2.700 ;
        RECT 4.725 1.830 5.450 2.060 ;
        RECT 6.245 0.680 6.475 2.470 ;
        RECT 6.965 2.060 7.195 4.360 ;
        RECT 7.990 2.470 8.715 2.700 ;
        RECT 6.965 1.830 7.690 2.060 ;
        RECT 8.485 0.680 8.715 2.470 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__fillcap_16

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__fillcap_32
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fillcap_32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.920 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.920 5.490 ;
        RECT 1.765 3.550 1.995 4.590 ;
        RECT 4.005 3.550 4.235 4.590 ;
        RECT 6.245 3.550 6.475 4.590 ;
        RECT 8.485 3.550 8.715 4.590 ;
        RECT 10.725 3.550 10.955 4.590 ;
        RECT 12.965 3.550 13.195 4.590 ;
        RECT 15.205 3.550 15.435 4.590 ;
        RECT 17.445 3.550 17.675 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 18.350 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 18.350 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 4.725 0.450 4.955 1.490 ;
        RECT 6.965 0.450 7.195 1.490 ;
        RECT 9.205 0.450 9.435 1.490 ;
        RECT 11.445 0.450 11.675 1.490 ;
        RECT 13.685 0.450 13.915 1.490 ;
        RECT 15.925 0.450 16.155 1.490 ;
        RECT 0.000 -0.450 17.920 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.060 0.475 4.360 ;
        RECT 0.245 1.830 0.970 2.060 ;
        RECT 1.325 1.490 1.555 2.755 ;
        RECT 2.485 2.060 2.715 4.360 ;
        RECT 2.485 1.830 3.210 2.060 ;
        RECT 3.565 1.490 3.795 2.755 ;
        RECT 4.725 2.060 4.955 4.360 ;
        RECT 4.725 1.830 5.450 2.060 ;
        RECT 5.805 1.490 6.035 2.755 ;
        RECT 6.965 2.060 7.195 4.360 ;
        RECT 6.965 1.830 7.690 2.060 ;
        RECT 8.045 1.490 8.275 2.755 ;
        RECT 9.205 2.060 9.435 4.360 ;
        RECT 9.205 1.830 9.930 2.060 ;
        RECT 10.285 1.490 10.515 2.755 ;
        RECT 11.445 2.060 11.675 4.360 ;
        RECT 11.445 1.830 12.170 2.060 ;
        RECT 12.525 1.490 12.755 2.755 ;
        RECT 13.685 2.060 13.915 4.360 ;
        RECT 13.685 1.830 14.410 2.060 ;
        RECT 14.765 1.490 14.995 2.755 ;
        RECT 15.925 2.060 16.155 4.360 ;
        RECT 15.925 1.830 16.650 2.060 ;
        RECT 17.005 1.490 17.235 2.755 ;
        RECT 1.325 1.260 1.995 1.490 ;
        RECT 3.565 1.260 4.235 1.490 ;
        RECT 5.805 1.260 6.475 1.490 ;
        RECT 8.045 1.260 8.715 1.490 ;
        RECT 10.285 1.260 10.955 1.490 ;
        RECT 12.525 1.260 13.195 1.490 ;
        RECT 14.765 1.260 15.435 1.490 ;
        RECT 17.005 1.260 17.675 1.490 ;
        RECT 1.765 0.680 1.995 1.260 ;
        RECT 4.005 0.680 4.235 1.260 ;
        RECT 6.245 0.680 6.475 1.260 ;
        RECT 8.485 0.680 8.715 1.260 ;
        RECT 10.725 0.680 10.955 1.260 ;
        RECT 12.965 0.680 13.195 1.260 ;
        RECT 15.205 0.680 15.435 1.260 ;
        RECT 17.445 0.680 17.675 1.260 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__fillcap_32

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__fillcap_64
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fillcap_64 ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.840 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 35.840 5.490 ;
        RECT 1.765 3.550 1.995 4.590 ;
        RECT 4.005 3.550 4.235 4.590 ;
        RECT 6.245 3.550 6.475 4.590 ;
        RECT 8.485 3.550 8.715 4.590 ;
        RECT 10.725 3.550 10.955 4.590 ;
        RECT 12.965 3.550 13.195 4.590 ;
        RECT 15.205 3.550 15.435 4.590 ;
        RECT 17.445 3.550 17.675 4.590 ;
        RECT 19.685 3.550 19.915 4.590 ;
        RECT 21.925 3.550 22.155 4.590 ;
        RECT 24.165 3.550 24.395 4.590 ;
        RECT 26.405 3.550 26.635 4.590 ;
        RECT 28.645 3.550 28.875 4.590 ;
        RECT 30.885 3.550 31.115 4.590 ;
        RECT 33.125 3.550 33.355 4.590 ;
        RECT 35.365 3.550 35.595 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 36.270 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 36.270 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 4.725 0.450 4.955 1.490 ;
        RECT 6.965 0.450 7.195 1.490 ;
        RECT 9.205 0.450 9.435 1.490 ;
        RECT 11.445 0.450 11.675 1.490 ;
        RECT 13.685 0.450 13.915 1.490 ;
        RECT 15.925 0.450 16.155 1.490 ;
        RECT 18.165 0.450 18.395 1.490 ;
        RECT 20.405 0.450 20.635 1.490 ;
        RECT 22.645 0.450 22.875 1.490 ;
        RECT 24.885 0.450 25.115 1.490 ;
        RECT 27.125 0.450 27.355 1.490 ;
        RECT 29.365 0.450 29.595 1.490 ;
        RECT 31.605 0.450 31.835 1.490 ;
        RECT 33.845 0.450 34.075 1.490 ;
        RECT 0.000 -0.450 35.840 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.060 0.475 4.360 ;
        RECT 0.245 1.830 0.970 2.060 ;
        RECT 1.325 1.490 1.555 2.755 ;
        RECT 2.485 2.060 2.715 4.360 ;
        RECT 2.485 1.830 3.210 2.060 ;
        RECT 3.565 1.490 3.795 2.755 ;
        RECT 4.725 2.060 4.955 4.360 ;
        RECT 4.725 1.830 5.450 2.060 ;
        RECT 5.805 1.490 6.035 2.755 ;
        RECT 6.965 2.060 7.195 4.360 ;
        RECT 6.965 1.830 7.690 2.060 ;
        RECT 8.045 1.490 8.275 2.755 ;
        RECT 9.205 2.060 9.435 4.360 ;
        RECT 9.205 1.830 9.930 2.060 ;
        RECT 10.285 1.490 10.515 2.755 ;
        RECT 11.445 2.060 11.675 4.360 ;
        RECT 11.445 1.830 12.170 2.060 ;
        RECT 12.525 1.490 12.755 2.755 ;
        RECT 13.685 2.060 13.915 4.360 ;
        RECT 13.685 1.830 14.410 2.060 ;
        RECT 14.765 1.490 14.995 2.755 ;
        RECT 15.925 2.060 16.155 4.360 ;
        RECT 15.925 1.830 16.650 2.060 ;
        RECT 17.005 1.490 17.235 2.755 ;
        RECT 18.165 2.060 18.395 4.360 ;
        RECT 18.165 1.830 18.890 2.060 ;
        RECT 19.245 1.490 19.475 2.755 ;
        RECT 20.405 2.060 20.635 4.360 ;
        RECT 20.405 1.830 21.130 2.060 ;
        RECT 21.485 1.490 21.715 2.755 ;
        RECT 22.645 2.060 22.875 4.360 ;
        RECT 22.645 1.830 23.370 2.060 ;
        RECT 23.725 1.490 23.955 2.755 ;
        RECT 24.885 2.060 25.115 4.360 ;
        RECT 24.885 1.830 25.610 2.060 ;
        RECT 25.965 1.490 26.195 2.755 ;
        RECT 27.125 2.060 27.355 4.360 ;
        RECT 27.125 1.830 27.850 2.060 ;
        RECT 28.205 1.490 28.435 2.755 ;
        RECT 29.365 2.060 29.595 4.360 ;
        RECT 29.365 1.830 30.090 2.060 ;
        RECT 30.445 1.490 30.675 2.755 ;
        RECT 31.605 2.060 31.835 4.360 ;
        RECT 31.605 1.830 32.330 2.060 ;
        RECT 32.685 1.490 32.915 2.755 ;
        RECT 33.845 2.060 34.075 4.360 ;
        RECT 33.845 1.830 34.570 2.060 ;
        RECT 34.925 1.490 35.155 2.755 ;
        RECT 1.325 1.260 1.995 1.490 ;
        RECT 3.565 1.260 4.235 1.490 ;
        RECT 5.805 1.260 6.475 1.490 ;
        RECT 8.045 1.260 8.715 1.490 ;
        RECT 10.285 1.260 10.955 1.490 ;
        RECT 12.525 1.260 13.195 1.490 ;
        RECT 14.765 1.260 15.435 1.490 ;
        RECT 17.005 1.260 17.675 1.490 ;
        RECT 19.245 1.260 19.915 1.490 ;
        RECT 21.485 1.260 22.155 1.490 ;
        RECT 23.725 1.260 24.395 1.490 ;
        RECT 25.965 1.260 26.635 1.490 ;
        RECT 28.205 1.260 28.875 1.490 ;
        RECT 30.445 1.260 31.115 1.490 ;
        RECT 32.685 1.260 33.355 1.490 ;
        RECT 34.925 1.260 35.595 1.490 ;
        RECT 1.765 0.680 1.995 1.260 ;
        RECT 4.005 0.680 4.235 1.260 ;
        RECT 6.245 0.680 6.475 1.260 ;
        RECT 8.485 0.680 8.715 1.260 ;
        RECT 10.725 0.680 10.955 1.260 ;
        RECT 12.965 0.680 13.195 1.260 ;
        RECT 15.205 0.680 15.435 1.260 ;
        RECT 17.445 0.680 17.675 1.260 ;
        RECT 19.685 0.680 19.915 1.260 ;
        RECT 21.925 0.680 22.155 1.260 ;
        RECT 24.165 0.680 24.395 1.260 ;
        RECT 26.405 0.680 26.635 1.260 ;
        RECT 28.645 0.680 28.875 1.260 ;
        RECT 30.885 0.680 31.115 1.260 ;
        RECT 33.125 0.680 33.355 1.260 ;
        RECT 35.365 0.680 35.595 1.260 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__fillcap_64

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__filltie
  CLASS core WELLTAP ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__filltie ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.120 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 1.550 5.470 ;
      LAYER Metal1 ;
        RECT 0.000 4.590 1.120 5.490 ;
        RECT 0.330 2.340 0.710 4.590 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 1.550 2.265 ;
      LAYER Metal1 ;
        RECT 0.330 0.450 0.710 1.910 ;
        RECT 0.000 -0.450 1.120 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__filltie

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__hold
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__hold ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.040 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN Z
    DIRECTION INOUT ;
    ANTENNAGATEAREA 1.707000 ;
    ANTENNADIFFAREA 0.489600 ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 1.645 0.575 3.605 ;
        RECT 3.510 1.645 3.950 2.575 ;
        RECT 0.245 1.415 3.950 1.645 ;
        RECT 0.245 0.845 0.475 1.415 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.040 5.490 ;
        RECT 3.225 3.265 3.455 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 5.470 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 5.470 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 3.225 0.450 3.455 1.185 ;
        RECT 0.000 -0.450 5.040 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 4.245 3.035 4.575 4.075 ;
        RECT 2.510 2.805 4.575 3.035 ;
        RECT 2.510 1.875 2.850 2.805 ;
        RECT 4.345 0.845 4.575 2.805 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__hold

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__icgtn_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__icgtn_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.800 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.220000 ;
    PORT
      LAYER Metal1 ;
        RECT 11.350 1.770 11.715 2.710 ;
    END
  END CLKN
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.210 1.770 2.090 2.265 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.265 0.410 2.710 ;
        RECT 0.150 1.770 0.915 2.265 ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.245200 ;
    PORT
      LAYER Metal1 ;
        RECT 16.195 3.830 16.475 4.200 ;
        RECT 15.830 3.390 16.475 3.830 ;
        RECT 16.245 1.590 16.475 3.390 ;
        RECT 15.830 1.210 16.475 1.590 ;
        RECT 16.245 0.795 16.475 1.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 16.800 5.490 ;
        RECT 0.675 3.390 0.905 4.590 ;
        RECT 5.805 3.390 6.035 4.590 ;
        RECT 8.665 3.390 8.895 4.590 ;
        RECT 12.245 3.390 12.475 4.590 ;
        RECT 15.175 3.390 15.405 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 17.230 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 17.230 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.450 1.650 1.080 ;
        RECT 5.805 0.450 6.035 1.135 ;
        RECT 8.765 0.450 8.995 1.135 ;
        RECT 12.165 0.450 12.395 1.135 ;
        RECT 14.405 0.450 14.635 1.135 ;
        RECT 15.125 0.450 15.355 1.605 ;
        RECT 0.000 -0.450 16.800 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.555 3.160 3.785 4.200 ;
        RECT 6.265 4.130 8.335 4.360 ;
        RECT 6.265 3.160 6.495 4.130 ;
        RECT 2.985 2.930 6.495 3.160 ;
        RECT 0.245 1.310 2.715 1.540 ;
        RECT 0.245 0.795 0.475 1.310 ;
        RECT 2.485 0.795 2.715 1.310 ;
        RECT 2.985 1.080 3.215 2.930 ;
        RECT 6.825 2.700 7.155 3.900 ;
        RECT 3.445 2.470 7.155 2.700 ;
        RECT 3.445 1.790 3.675 2.470 ;
        RECT 2.985 0.850 3.890 1.080 ;
        RECT 6.925 0.795 7.155 2.470 ;
        RECT 7.645 1.695 7.875 3.900 ;
        RECT 8.105 1.925 8.335 4.130 ;
        RECT 9.685 4.130 12.015 4.360 ;
        RECT 8.565 1.980 9.390 2.210 ;
        RECT 8.565 1.695 8.795 1.980 ;
        RECT 7.645 1.465 8.795 1.695 ;
        RECT 7.645 0.795 7.875 1.465 ;
        RECT 9.685 0.795 10.115 4.130 ;
        RECT 11.225 3.170 11.455 3.900 ;
        RECT 10.385 2.940 11.455 3.170 ;
        RECT 11.785 3.160 12.015 4.130 ;
        RECT 10.385 1.080 10.615 2.940 ;
        RECT 11.785 2.930 12.915 3.160 ;
        RECT 12.685 1.925 12.915 2.930 ;
        RECT 14.005 2.210 14.235 4.200 ;
        RECT 14.005 1.980 15.740 2.210 ;
        RECT 14.005 1.520 14.235 1.980 ;
        RECT 13.285 1.290 14.235 1.520 ;
        RECT 10.385 0.850 11.330 1.080 ;
        RECT 13.285 0.795 13.515 1.290 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__icgtn_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__icgtn_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__icgtn_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.920 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.640000 ;
    PORT
      LAYER Metal1 ;
        RECT 11.350 1.770 11.675 2.710 ;
    END
  END CLKN
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.390 1.770 2.650 2.710 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 0.970 2.710 ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.471600 ;
    PORT
      LAYER Metal1 ;
        RECT 16.275 0.815 16.650 4.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.920 5.490 ;
        RECT 1.435 3.400 1.665 4.590 ;
        RECT 5.805 3.400 6.035 4.590 ;
        RECT 8.625 3.400 8.855 4.590 ;
        RECT 12.025 3.400 12.255 4.590 ;
        RECT 15.255 3.400 15.485 4.590 ;
        RECT 17.295 3.400 17.525 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 18.350 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 18.350 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.450 1.650 1.100 ;
        RECT 5.565 0.450 5.795 1.155 ;
        RECT 8.525 0.450 8.755 1.155 ;
        RECT 11.925 0.450 12.155 1.155 ;
        RECT 14.165 0.450 14.395 1.155 ;
        RECT 15.205 0.450 15.435 1.625 ;
        RECT 17.445 0.450 17.675 1.625 ;
        RECT 0.000 -0.450 17.920 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 4.045 3.170 4.275 4.210 ;
        RECT 6.265 4.130 8.345 4.360 ;
        RECT 6.265 3.170 6.495 4.130 ;
        RECT 4.045 3.065 6.495 3.170 ;
        RECT 2.930 2.940 6.495 3.065 ;
        RECT 2.930 2.835 4.240 2.940 ;
        RECT 2.930 1.615 3.160 2.835 ;
        RECT 4.435 2.075 4.775 2.710 ;
        RECT 6.825 2.075 7.055 3.900 ;
        RECT 3.390 1.845 7.055 2.075 ;
        RECT 1.065 1.540 2.295 1.560 ;
        RECT 0.245 1.330 2.295 1.540 ;
        RECT 2.930 1.385 3.835 1.615 ;
        RECT 0.245 1.310 1.160 1.330 ;
        RECT 0.245 0.815 0.475 1.310 ;
        RECT 2.065 1.155 2.295 1.330 ;
        RECT 2.065 0.815 2.715 1.155 ;
        RECT 3.605 0.815 3.835 1.385 ;
        RECT 6.685 0.815 7.055 1.845 ;
        RECT 7.405 1.655 7.835 3.900 ;
        RECT 8.115 1.885 8.345 4.130 ;
        RECT 9.645 3.980 11.795 4.210 ;
        RECT 8.575 1.940 9.350 2.170 ;
        RECT 8.575 1.655 8.805 1.940 ;
        RECT 7.405 1.425 8.805 1.655 ;
        RECT 7.405 0.815 7.635 1.425 ;
        RECT 9.645 0.815 9.875 3.980 ;
        RECT 11.005 3.140 11.235 3.720 ;
        RECT 10.305 2.910 11.235 3.140 ;
        RECT 11.565 3.170 11.795 3.980 ;
        RECT 11.565 2.940 12.695 3.170 ;
        RECT 10.305 1.540 10.535 2.910 ;
        RECT 12.465 2.415 12.695 2.940 ;
        RECT 13.785 2.170 14.015 4.210 ;
        RECT 13.785 1.940 15.980 2.170 ;
        RECT 13.785 1.560 14.015 1.940 ;
        RECT 10.305 1.310 11.090 1.540 ;
        RECT 12.990 1.330 14.015 1.560 ;
        RECT 12.990 1.310 13.330 1.330 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__icgtn_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__icgtn_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__icgtn_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.160 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.640000 ;
    PORT
      LAYER Metal1 ;
        RECT 11.350 1.770 11.610 2.710 ;
    END
  END CLKN
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.345 1.820 2.650 3.270 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 0.970 2.710 ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.943200 ;
    PORT
      LAYER Metal1 ;
        RECT 16.030 2.920 16.260 3.960 ;
        RECT 18.070 2.920 18.550 3.960 ;
        RECT 16.030 2.690 18.550 2.920 ;
        RECT 18.070 1.600 18.550 2.690 ;
        RECT 16.030 1.300 18.550 1.600 ;
        RECT 16.030 0.790 16.310 1.300 ;
        RECT 18.320 0.790 18.550 1.300 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 20.160 5.490 ;
        RECT 1.325 3.150 1.555 4.590 ;
        RECT 5.820 3.150 6.050 4.590 ;
        RECT 8.580 3.150 8.810 4.590 ;
        RECT 12.080 3.785 12.310 4.590 ;
        RECT 15.010 3.150 15.240 4.590 ;
        RECT 17.050 3.150 17.280 4.590 ;
        RECT 19.090 3.150 19.320 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 20.590 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 20.590 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.450 1.650 1.075 ;
        RECT 5.580 0.450 5.810 1.130 ;
        RECT 8.580 0.450 8.810 1.130 ;
        RECT 11.980 0.450 12.210 1.130 ;
        RECT 14.220 0.450 14.450 1.130 ;
        RECT 14.960 0.450 15.190 1.600 ;
        RECT 17.200 0.450 17.430 1.070 ;
        RECT 19.440 0.450 19.670 1.600 ;
        RECT 0.000 -0.450 20.160 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 6.280 4.130 8.250 4.360 ;
        RECT 4.060 2.920 4.290 3.960 ;
        RECT 6.280 2.920 6.510 4.130 ;
        RECT 4.060 2.795 6.510 2.920 ;
        RECT 2.945 2.690 6.510 2.795 ;
        RECT 2.945 2.565 4.265 2.690 ;
        RECT 2.945 1.615 3.175 2.565 ;
        RECT 4.470 2.075 4.810 2.460 ;
        RECT 6.840 2.075 7.070 3.900 ;
        RECT 3.405 1.845 7.070 2.075 ;
        RECT 0.245 1.305 2.715 1.535 ;
        RECT 2.945 1.385 3.850 1.615 ;
        RECT 0.245 0.790 0.475 1.305 ;
        RECT 2.485 0.790 2.715 1.305 ;
        RECT 3.620 0.790 3.850 1.385 ;
        RECT 6.700 0.790 7.070 1.845 ;
        RECT 7.460 1.590 7.790 3.900 ;
        RECT 8.020 1.820 8.250 4.130 ;
        RECT 9.600 3.735 9.830 3.960 ;
        RECT 9.600 3.555 11.855 3.735 ;
        RECT 9.600 3.505 12.750 3.555 ;
        RECT 8.480 1.875 9.305 2.105 ;
        RECT 8.480 1.590 8.710 1.875 ;
        RECT 7.460 1.360 8.710 1.590 ;
        RECT 7.460 0.790 7.690 1.360 ;
        RECT 9.600 0.790 9.930 3.505 ;
        RECT 11.630 3.325 12.750 3.505 ;
        RECT 10.860 2.935 11.290 3.275 ;
        RECT 10.360 1.460 10.590 2.200 ;
        RECT 10.860 1.460 11.090 2.935 ;
        RECT 12.520 2.475 12.750 3.325 ;
        RECT 13.840 2.320 14.070 3.960 ;
        RECT 13.840 1.980 17.510 2.320 ;
        RECT 13.840 1.535 14.070 1.980 ;
        RECT 10.360 1.230 11.090 1.460 ;
        RECT 13.045 1.305 14.070 1.535 ;
        RECT 13.045 1.285 13.385 1.305 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__icgtn_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__icgtp_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__icgtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.120 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.220000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.230 1.770 10.490 2.710 ;
    END
  END CLK
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.255 2.710 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.270 1.190 2.500 ;
        RECT 0.150 1.210 0.410 2.270 ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.245200 ;
    PORT
      LAYER Metal1 ;
        RECT 14.150 0.695 14.610 3.685 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 15.120 5.490 ;
        RECT 0.845 3.435 1.075 4.590 ;
        RECT 6.025 3.910 6.255 4.590 ;
        RECT 8.980 4.235 9.210 4.590 ;
        RECT 8.980 4.005 13.240 4.235 ;
        RECT 8.980 3.895 11.200 4.005 ;
        RECT 13.010 3.425 13.240 4.005 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 15.550 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 15.550 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.530 0.450 1.870 1.075 ;
        RECT 5.785 0.450 6.015 1.130 ;
        RECT 9.260 0.450 9.490 1.035 ;
        RECT 13.260 0.450 13.490 1.015 ;
        RECT 0.000 -0.450 15.120 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.205 3.175 3.595 4.245 ;
        RECT 7.045 3.640 7.275 4.245 ;
        RECT 5.680 3.410 10.975 3.640 ;
        RECT 3.205 2.945 5.450 3.175 ;
        RECT 0.640 1.305 2.935 1.535 ;
        RECT 0.640 0.980 0.870 1.305 ;
        RECT 0.190 0.750 0.870 0.980 ;
        RECT 2.705 0.790 2.935 1.305 ;
        RECT 3.205 1.075 3.435 2.945 ;
        RECT 3.665 2.485 4.990 2.715 ;
        RECT 3.665 1.790 3.895 2.485 ;
        RECT 5.220 1.985 5.450 2.945 ;
        RECT 5.680 2.215 5.910 3.410 ;
        RECT 6.140 2.270 6.750 2.500 ;
        RECT 6.140 1.985 6.370 2.270 ;
        RECT 5.220 1.755 6.370 1.985 ;
        RECT 6.980 1.130 7.210 3.410 ;
        RECT 8.135 2.605 8.475 3.180 ;
        RECT 7.565 2.375 8.475 2.605 ;
        RECT 9.770 2.950 10.515 3.180 ;
        RECT 9.770 2.500 10.000 2.950 ;
        RECT 3.205 0.845 4.110 1.075 ;
        RECT 6.905 0.790 7.210 1.130 ;
        RECT 8.140 0.695 8.475 2.375 ;
        RECT 8.715 2.270 10.000 2.500 ;
        RECT 10.745 2.500 10.975 3.410 ;
        RECT 11.990 3.105 12.220 3.685 ;
        RECT 11.990 2.875 13.015 3.105 ;
        RECT 12.785 2.500 13.015 2.875 ;
        RECT 10.745 2.270 12.555 2.500 ;
        RECT 12.785 2.270 13.915 2.500 ;
        RECT 9.770 0.980 10.000 2.270 ;
        RECT 12.785 1.035 13.015 2.270 ;
        RECT 9.770 0.750 10.665 0.980 ;
        RECT 11.100 0.695 13.015 1.035 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__icgtp_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__icgtp_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__icgtp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.680 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.625000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.230 1.210 10.490 2.405 ;
    END
  END CLK
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.210 1.770 2.090 2.350 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 0.970 2.710 ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.471600 ;
    PORT
      LAYER Metal1 ;
        RECT 13.590 2.890 14.200 3.685 ;
        RECT 13.940 1.590 14.200 2.890 ;
        RECT 13.590 1.210 14.200 1.590 ;
        RECT 13.940 0.790 14.200 1.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 15.680 5.490 ;
        RECT 0.695 3.440 0.925 4.590 ;
        RECT 5.805 3.850 6.035 4.590 ;
        RECT 8.720 4.250 8.950 4.590 ;
        RECT 8.720 4.020 15.220 4.250 ;
        RECT 8.720 3.850 11.140 4.020 ;
        RECT 12.950 3.440 13.180 4.020 ;
        RECT 14.990 3.440 15.220 4.020 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 16.110 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 16.110 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.450 1.650 1.075 ;
        RECT 5.620 0.450 5.850 1.130 ;
        RECT 9.020 0.450 9.250 1.130 ;
        RECT 12.820 0.450 13.050 1.430 ;
        RECT 15.060 0.450 15.290 1.430 ;
        RECT 0.000 -0.450 15.680 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.555 3.175 3.785 4.250 ;
        RECT 6.825 3.620 7.055 4.250 ;
        RECT 5.460 3.390 11.700 3.620 ;
        RECT 2.985 2.945 5.230 3.175 ;
        RECT 0.245 1.305 2.715 1.535 ;
        RECT 0.245 0.790 0.475 1.305 ;
        RECT 2.485 0.790 2.715 1.305 ;
        RECT 2.985 1.075 3.215 2.945 ;
        RECT 3.445 2.485 4.770 2.715 ;
        RECT 3.445 1.790 3.675 2.485 ;
        RECT 5.000 1.835 5.230 2.945 ;
        RECT 5.460 2.065 5.690 3.390 ;
        RECT 6.005 1.835 6.345 2.350 ;
        RECT 5.000 1.605 6.345 1.835 ;
        RECT 2.985 0.845 3.890 1.075 ;
        RECT 6.740 0.790 6.970 3.390 ;
        RECT 7.400 2.930 7.985 3.160 ;
        RECT 9.685 2.930 10.025 3.160 ;
        RECT 7.400 1.075 7.630 2.930 ;
        RECT 9.685 2.350 9.915 2.930 ;
        RECT 8.225 2.120 9.915 2.350 ;
        RECT 11.470 2.350 11.700 3.390 ;
        RECT 11.930 3.105 12.160 3.685 ;
        RECT 11.930 2.875 12.885 3.105 ;
        RECT 12.655 2.405 12.885 2.875 ;
        RECT 11.470 2.120 12.425 2.350 ;
        RECT 7.400 0.845 8.185 1.075 ;
        RECT 9.685 0.980 9.915 2.120 ;
        RECT 12.655 2.065 13.490 2.405 ;
        RECT 12.655 1.890 12.885 2.065 ;
        RECT 10.860 1.660 12.885 1.890 ;
        RECT 9.685 0.750 10.425 0.980 ;
        RECT 10.860 0.790 11.090 1.660 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__icgtp_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__icgtp_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__icgtp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.920 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.625000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.230 1.770 10.490 2.710 ;
    END
  END CLK
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.405 0.970 2.710 ;
        RECT 0.710 2.175 2.090 2.405 ;
        RECT 0.710 1.770 0.970 2.175 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 1.770 0.415 2.710 ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.943200 ;
    PORT
      LAYER Metal1 ;
        RECT 13.885 3.105 14.145 3.685 ;
        RECT 15.955 3.105 16.355 3.685 ;
        RECT 13.885 2.875 16.355 3.105 ;
        RECT 15.955 1.745 16.355 2.875 ;
        RECT 13.885 1.515 16.355 1.745 ;
        RECT 13.885 0.795 14.115 1.515 ;
        RECT 15.770 0.710 16.355 1.515 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.920 5.490 ;
        RECT 0.625 3.440 0.855 4.590 ;
        RECT 5.805 3.855 6.035 4.590 ;
        RECT 8.865 3.855 9.095 4.590 ;
        RECT 10.855 3.855 11.085 4.590 ;
        RECT 12.895 4.250 13.125 4.590 ;
        RECT 12.895 4.020 17.205 4.250 ;
        RECT 12.895 3.440 13.125 4.020 ;
        RECT 14.935 3.440 15.165 4.020 ;
        RECT 16.975 3.440 17.205 4.020 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 18.350 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 18.350 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.450 1.650 1.080 ;
        RECT 5.565 0.450 5.795 1.135 ;
        RECT 8.965 0.450 9.195 1.135 ;
        RECT 12.765 0.450 12.995 1.485 ;
        RECT 15.005 0.450 15.235 1.035 ;
        RECT 17.245 0.450 17.475 1.485 ;
        RECT 0.000 -0.450 17.920 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 4.035 3.230 4.265 4.250 ;
        RECT 6.825 3.625 7.055 4.250 ;
        RECT 5.405 3.395 11.645 3.625 ;
        RECT 4.035 3.050 5.175 3.230 ;
        RECT 2.985 3.000 5.175 3.050 ;
        RECT 2.985 2.820 4.260 3.000 ;
        RECT 0.245 1.310 2.715 1.540 ;
        RECT 0.245 0.795 0.475 1.310 ;
        RECT 2.485 0.795 2.715 1.310 ;
        RECT 2.985 1.080 3.215 2.820 ;
        RECT 4.485 2.130 4.715 2.770 ;
        RECT 3.445 1.790 4.715 2.130 ;
        RECT 4.945 1.890 5.175 3.000 ;
        RECT 5.405 2.120 5.635 3.395 ;
        RECT 5.865 2.175 6.530 2.405 ;
        RECT 5.865 1.890 6.095 2.175 ;
        RECT 4.945 1.660 6.095 1.890 ;
        RECT 6.760 1.135 6.990 3.395 ;
        RECT 7.790 2.460 8.130 3.160 ;
        RECT 7.345 2.120 8.130 2.460 ;
        RECT 9.770 2.935 10.170 3.165 ;
        RECT 9.770 2.405 10.000 2.935 ;
        RECT 8.370 2.175 10.000 2.405 ;
        RECT 11.415 2.405 11.645 3.395 ;
        RECT 11.875 3.105 12.105 3.685 ;
        RECT 11.875 2.875 13.060 3.105 ;
        RECT 11.415 2.175 12.600 2.405 ;
        RECT 12.830 2.315 13.060 2.875 ;
        RECT 2.985 0.850 3.890 1.080 ;
        RECT 6.685 0.795 6.990 1.135 ;
        RECT 7.845 0.795 8.130 2.120 ;
        RECT 9.770 1.540 10.000 2.175 ;
        RECT 12.830 1.975 15.370 2.315 ;
        RECT 12.830 1.945 13.060 1.975 ;
        RECT 10.805 1.715 13.060 1.945 ;
        RECT 9.770 1.310 10.315 1.540 ;
        RECT 10.085 0.795 10.315 1.310 ;
        RECT 10.805 0.795 11.035 1.715 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__icgtp_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__inv_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__inv_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.240 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.300 1.070 2.530 ;
        RECT 0.710 1.210 1.015 2.300 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 2.150 1.595 4.360 ;
        RECT 1.270 0.680 1.595 2.150 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 2.240 5.490 ;
        RECT 0.345 3.550 0.575 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 2.670 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 2.670 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 0.000 -0.450 2.240 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__inv_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__inv_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__inv_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 2.270 1.910 2.710 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.915500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.395 3.830 1.625 4.360 ;
        RECT 1.395 3.450 2.370 3.830 ;
        RECT 2.140 1.850 2.370 3.450 ;
        RECT 1.830 1.670 2.370 1.850 ;
        RECT 1.830 1.490 2.285 1.670 ;
        RECT 1.395 1.210 2.285 1.490 ;
        RECT 1.395 0.680 1.625 1.210 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 3.360 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.600 3.550 2.830 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 3.790 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 3.790 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.515 0.450 2.745 1.490 ;
        RECT 0.000 -0.450 3.360 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__inv_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__inv_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__inv_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.121000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.410 2.270 2.160 2.710 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.207000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.505 3.320 3.735 4.360 ;
        RECT 1.365 3.090 3.735 3.320 ;
        RECT 2.390 1.950 2.805 3.090 ;
        RECT 1.365 1.720 3.835 1.950 ;
        RECT 1.365 0.680 1.595 1.720 ;
        RECT 3.605 0.680 3.835 1.720 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 4.480 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 4.910 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 0.000 -0.450 4.480 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__inv_3

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__inv_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__inv_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.580 2.270 2.330 2.650 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.642000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.350 1.595 4.360 ;
        RECT 3.505 3.350 3.835 4.360 ;
        RECT 1.365 3.120 3.835 3.350 ;
        RECT 3.335 1.890 3.835 3.120 ;
        RECT 1.365 1.660 3.835 1.890 ;
        RECT 1.365 0.680 1.595 1.660 ;
        RECT 3.605 0.680 3.835 1.660 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.600 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.580 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.430 ;
        RECT 2.485 0.450 2.715 1.430 ;
        RECT 4.725 0.450 4.955 1.430 ;
        RECT 0.000 -0.450 5.600 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__inv_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__inv_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__inv_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 13.655999 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 2.265 4.260 2.645 ;
        RECT 5.360 2.215 8.880 2.650 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 7.284000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.505 3.320 3.735 4.360 ;
        RECT 5.745 3.320 5.975 4.360 ;
        RECT 7.985 3.320 8.215 4.360 ;
        RECT 1.365 3.090 8.215 3.320 ;
        RECT 4.630 1.985 5.130 3.090 ;
        RECT 1.365 1.755 8.315 1.985 ;
        RECT 1.365 0.680 1.595 1.755 ;
        RECT 3.575 0.680 3.835 1.755 ;
        RECT 5.845 0.680 6.075 1.755 ;
        RECT 8.085 0.680 8.315 1.755 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 10.080 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
        RECT 9.105 3.550 9.335 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 10.510 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 10.510 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 4.725 0.450 4.955 1.165 ;
        RECT 6.965 0.450 7.195 1.490 ;
        RECT 9.205 0.450 9.435 1.490 ;
        RECT 0.000 -0.450 10.080 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__inv_8

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__inv_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__inv_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.560 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 20.483999 ;
    PORT
      LAYER Metal1 ;
        RECT 0.180 2.270 5.690 2.650 ;
        RECT 7.600 2.215 13.000 2.650 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 10.926000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.505 3.320 3.735 4.360 ;
        RECT 5.745 3.320 5.975 4.360 ;
        RECT 7.985 3.320 8.215 4.360 ;
        RECT 10.225 3.320 10.455 4.360 ;
        RECT 12.465 3.320 12.695 4.360 ;
        RECT 1.365 3.090 12.695 3.320 ;
        RECT 6.755 1.950 7.370 3.090 ;
        RECT 1.365 1.720 12.795 1.950 ;
        RECT 1.365 0.680 1.625 1.720 ;
        RECT 3.605 0.680 3.835 1.720 ;
        RECT 5.845 0.680 6.075 1.720 ;
        RECT 8.085 0.680 8.315 1.720 ;
        RECT 10.325 0.680 10.555 1.720 ;
        RECT 12.565 0.680 12.795 1.720 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 14.560 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
        RECT 9.105 3.550 9.335 4.590 ;
        RECT 11.345 3.550 11.575 4.590 ;
        RECT 13.585 3.550 13.815 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 14.990 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.990 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 4.725 0.450 4.955 1.490 ;
        RECT 6.965 0.450 7.195 1.490 ;
        RECT 9.205 0.450 9.435 1.490 ;
        RECT 11.445 0.450 11.675 1.490 ;
        RECT 13.685 0.450 13.915 1.490 ;
        RECT 0.000 -0.450 14.560 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__inv_12

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__inv_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__inv_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.040 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 27.311998 ;
    PORT
      LAYER Metal1 ;
        RECT 0.685 2.215 7.965 2.650 ;
        RECT 9.225 2.215 16.505 2.650 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 14.568000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.210 1.595 4.360 ;
        RECT 3.505 3.210 3.735 4.360 ;
        RECT 5.745 3.210 5.975 4.360 ;
        RECT 8.080 3.210 8.310 4.360 ;
        RECT 1.365 3.180 8.310 3.210 ;
        RECT 10.225 3.180 10.455 4.360 ;
        RECT 12.465 3.180 12.695 4.360 ;
        RECT 14.705 3.180 14.935 4.360 ;
        RECT 16.945 3.180 17.175 4.360 ;
        RECT 1.365 2.980 17.175 3.180 ;
        RECT 8.195 2.950 17.175 2.980 ;
        RECT 8.195 1.950 8.995 2.950 ;
        RECT 1.365 1.720 17.275 1.950 ;
        RECT 1.365 0.680 1.625 1.720 ;
        RECT 3.605 0.680 3.835 1.720 ;
        RECT 5.845 0.680 6.075 1.720 ;
        RECT 8.085 0.680 8.315 1.720 ;
        RECT 10.325 0.680 10.555 1.720 ;
        RECT 12.565 0.680 12.795 1.720 ;
        RECT 14.805 0.680 15.035 1.720 ;
        RECT 17.045 0.680 17.275 1.720 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 19.040 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
        RECT 9.105 3.550 9.335 4.590 ;
        RECT 11.345 3.550 11.575 4.590 ;
        RECT 13.585 3.550 13.815 4.590 ;
        RECT 15.825 3.550 16.055 4.590 ;
        RECT 18.065 3.550 18.295 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 19.470 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 19.470 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 4.725 0.450 4.955 1.490 ;
        RECT 6.965 0.450 7.195 1.490 ;
        RECT 9.205 0.450 9.435 1.490 ;
        RECT 11.445 0.450 11.675 1.490 ;
        RECT 13.685 0.450 13.915 1.490 ;
        RECT 15.925 0.450 16.155 1.490 ;
        RECT 18.165 0.450 18.395 1.490 ;
        RECT 0.000 -0.450 19.040 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__inv_16

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__inv_20
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__inv_20 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 34.139999 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 2.270 9.900 2.650 ;
        RECT 11.110 2.270 20.380 2.650 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 18.209999 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.505 3.320 3.735 4.360 ;
        RECT 5.745 3.320 5.975 4.360 ;
        RECT 7.985 3.320 8.215 4.360 ;
        RECT 10.225 3.320 10.455 4.360 ;
        RECT 12.465 3.320 12.695 4.360 ;
        RECT 14.705 3.320 14.935 4.360 ;
        RECT 16.945 3.320 17.175 4.360 ;
        RECT 19.185 3.320 19.415 4.360 ;
        RECT 21.425 3.320 21.655 4.360 ;
        RECT 1.365 3.090 21.655 3.320 ;
        RECT 10.130 1.950 10.880 3.090 ;
        RECT 1.335 1.720 21.755 1.950 ;
        RECT 1.335 0.680 1.595 1.720 ;
        RECT 3.605 0.680 3.835 1.720 ;
        RECT 5.845 0.680 6.075 1.720 ;
        RECT 8.085 0.680 8.315 1.720 ;
        RECT 10.325 0.680 10.555 1.720 ;
        RECT 12.565 0.680 12.795 1.720 ;
        RECT 14.805 0.680 15.035 1.720 ;
        RECT 17.045 0.680 17.275 1.720 ;
        RECT 19.285 0.680 19.515 1.720 ;
        RECT 21.525 0.680 21.755 1.720 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 23.520 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
        RECT 9.105 3.550 9.335 4.590 ;
        RECT 11.345 3.550 11.575 4.590 ;
        RECT 13.585 3.550 13.815 4.590 ;
        RECT 15.825 3.550 16.055 4.590 ;
        RECT 18.065 3.550 18.295 4.590 ;
        RECT 20.305 3.550 20.535 4.590 ;
        RECT 22.545 3.550 22.775 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 23.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 23.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 4.725 0.450 4.955 1.490 ;
        RECT 6.965 0.450 7.195 1.490 ;
        RECT 9.205 0.450 9.435 1.490 ;
        RECT 11.445 0.450 11.675 1.490 ;
        RECT 13.685 0.450 13.915 1.490 ;
        RECT 15.925 0.450 16.155 1.490 ;
        RECT 18.165 0.450 18.395 1.490 ;
        RECT 20.405 0.450 20.635 1.490 ;
        RECT 22.645 0.450 22.875 1.490 ;
        RECT 0.000 -0.450 23.520 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__inv_20

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__invz_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__invz_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.698000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.015 0.970 2.710 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.849000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.505 1.770 8.810 2.710 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.372800 ;
    PORT
      LAYER Metal1 ;
        RECT 4.610 1.770 4.890 3.900 ;
        RECT 4.610 1.140 4.840 1.770 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 9.520 5.490 ;
        RECT 1.265 3.480 1.495 4.590 ;
        RECT 5.680 3.860 5.910 4.590 ;
        RECT 7.585 3.480 7.815 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 9.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.610 0.450 1.840 1.480 ;
        RECT 5.730 0.450 5.960 1.165 ;
        RECT 7.585 0.450 7.815 1.480 ;
        RECT 0.000 -0.450 9.520 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.250 0.475 4.290 ;
        RECT 2.335 4.130 5.350 4.360 ;
        RECT 2.335 3.480 2.565 4.130 ;
        RECT 0.245 3.020 3.060 3.250 ;
        RECT 2.105 2.245 2.335 3.020 ;
        RECT 1.200 2.015 2.335 2.245 ;
        RECT 1.200 1.820 1.430 2.015 ;
        RECT 1.095 1.625 1.430 1.820 ;
        RECT 1.095 1.425 1.325 1.625 ;
        RECT 3.355 1.425 3.585 3.820 ;
        RECT 0.190 1.195 1.325 1.425 ;
        RECT 2.675 1.195 3.585 1.425 ;
        RECT 3.355 0.910 3.585 1.195 ;
        RECT 3.850 1.140 4.080 4.130 ;
        RECT 5.120 3.630 5.350 4.130 ;
        RECT 6.565 3.630 6.795 4.290 ;
        RECT 5.120 3.400 6.795 3.630 ;
        RECT 5.120 2.430 5.415 3.400 ;
        RECT 8.945 3.380 9.175 4.290 ;
        RECT 8.045 3.150 9.175 3.380 ;
        RECT 8.045 2.245 8.275 3.150 ;
        RECT 5.145 1.625 5.375 2.170 ;
        RECT 7.090 2.015 8.275 2.245 ;
        RECT 5.145 1.565 6.695 1.625 ;
        RECT 5.070 1.395 6.695 1.565 ;
        RECT 5.070 0.910 5.300 1.395 ;
        RECT 6.465 1.140 6.695 1.395 ;
        RECT 8.045 1.425 8.275 2.015 ;
        RECT 8.045 1.195 9.330 1.425 ;
        RECT 3.355 0.680 5.300 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__invz_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__invz_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__invz_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 0.970 2.710 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.692000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.990 1.770 8.460 2.710 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.622400 ;
    PORT
      LAYER Metal1 ;
        RECT 6.770 2.710 7.000 3.750 ;
        RECT 6.770 1.490 7.130 2.710 ;
        RECT 6.620 1.210 7.130 1.490 ;
        RECT 6.620 0.680 6.850 1.210 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 9.520 5.490 ;
        RECT 1.370 3.400 1.600 4.590 ;
        RECT 5.750 4.350 5.980 4.590 ;
        RECT 7.790 3.400 8.020 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 9.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.420 0.450 1.650 1.020 ;
        RECT 5.500 0.450 5.730 1.020 ;
        RECT 7.740 0.450 7.970 1.490 ;
        RECT 0.000 -0.450 9.520 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.350 3.170 0.580 4.210 ;
        RECT 2.900 4.130 4.960 4.360 ;
        RECT 2.900 3.400 3.130 4.130 ;
        RECT 0.350 2.940 3.625 3.170 ;
        RECT 1.860 2.470 3.625 2.940 ;
        RECT 1.860 1.490 2.090 2.470 ;
        RECT 3.920 2.240 4.150 3.900 ;
        RECT 3.200 2.010 4.150 2.240 ;
        RECT 4.585 2.220 4.960 4.130 ;
        RECT 6.165 3.980 7.560 4.210 ;
        RECT 6.165 3.155 6.395 3.980 ;
        RECT 5.240 2.925 6.395 3.155 ;
        RECT 7.330 3.170 7.560 3.980 ;
        RECT 8.810 3.170 9.090 4.210 ;
        RECT 7.330 2.940 9.090 3.170 ;
        RECT 5.240 2.450 5.470 2.925 ;
        RECT 5.700 2.465 6.475 2.695 ;
        RECT 5.700 2.220 5.930 2.465 ;
        RECT 3.200 1.490 3.430 2.010 ;
        RECT 4.585 1.990 5.930 2.220 ;
        RECT 4.585 1.780 4.815 1.990 ;
        RECT 0.300 1.260 2.090 1.490 ;
        RECT 0.300 0.680 0.530 1.260 ;
        RECT 2.540 1.085 3.430 1.490 ;
        RECT 3.660 1.550 4.815 1.780 ;
        RECT 3.660 1.315 3.890 1.550 ;
        RECT 6.160 1.480 6.390 2.110 ;
        RECT 5.035 1.250 6.390 1.480 ;
        RECT 5.035 1.085 5.265 1.250 ;
        RECT 2.540 0.680 5.265 1.085 ;
        RECT 8.860 0.680 9.090 2.940 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__invz_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__invz_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__invz_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.880 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 0.970 2.710 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.692000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.190 1.770 5.645 2.710 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.995200 ;
    PORT
      LAYER Metal1 ;
        RECT 9.465 3.195 9.930 4.210 ;
        RECT 11.505 3.195 11.735 4.210 ;
        RECT 9.465 2.965 12.495 3.195 ;
        RECT 12.265 1.600 12.495 2.965 ;
        RECT 10.025 1.370 12.495 1.600 ;
        RECT 10.025 0.790 10.255 1.370 ;
        RECT 12.265 0.840 12.495 1.370 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 12.880 5.490 ;
        RECT 1.370 3.845 1.600 4.590 ;
        RECT 6.045 4.280 6.275 4.590 ;
        RECT 8.265 3.400 8.495 4.590 ;
        RECT 10.485 3.880 10.715 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 13.310 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 13.310 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.420 0.450 1.650 1.020 ;
        RECT 6.235 0.450 6.575 0.620 ;
        RECT 8.725 0.450 8.955 1.160 ;
        RECT 11.145 0.450 11.375 1.020 ;
        RECT 0.000 -0.450 12.880 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.350 3.170 0.580 4.210 ;
        RECT 2.895 4.050 5.825 4.210 ;
        RECT 2.895 3.980 7.475 4.050 ;
        RECT 2.895 3.400 3.125 3.980 ;
        RECT 0.350 2.940 3.565 3.170 ;
        RECT 3.335 2.060 3.565 2.940 ;
        RECT 1.200 1.830 3.565 2.060 ;
        RECT 3.795 2.940 4.145 3.750 ;
        RECT 1.200 1.540 1.430 1.830 ;
        RECT 0.300 1.310 1.430 1.540 ;
        RECT 3.795 1.490 4.025 2.940 ;
        RECT 4.375 1.655 4.605 3.980 ;
        RECT 5.605 3.820 7.475 3.980 ;
        RECT 5.025 3.170 5.255 3.750 ;
        RECT 5.025 2.940 6.980 3.170 ;
        RECT 0.300 0.680 0.530 1.310 ;
        RECT 2.540 1.080 4.025 1.490 ;
        RECT 4.255 1.315 4.605 1.655 ;
        RECT 6.750 2.060 6.980 2.940 ;
        RECT 7.245 2.735 7.475 3.820 ;
        RECT 7.245 2.505 11.365 2.735 ;
        RECT 6.750 1.540 7.090 2.060 ;
        RECT 4.920 1.310 7.090 1.540 ;
        RECT 7.605 1.830 12.030 2.060 ;
        RECT 7.605 1.080 7.835 1.830 ;
        RECT 2.540 0.850 7.835 1.080 ;
        RECT 2.540 0.680 2.770 0.850 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__invz_3

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__invz_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__invz_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.440 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.060 0.410 2.710 ;
        RECT 0.150 1.770 1.020 2.060 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.692000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.130 1.830 6.070 2.650 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.244800 ;
    PORT
      LAYER Metal1 ;
        RECT 9.110 3.310 9.410 3.900 ;
        RECT 11.190 3.310 11.870 3.900 ;
        RECT 9.110 2.965 11.870 3.310 ;
        RECT 11.585 1.620 11.870 2.965 ;
        RECT 9.180 1.390 11.870 1.620 ;
        RECT 9.180 0.730 9.630 1.390 ;
        RECT 11.640 0.730 11.870 1.390 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 13.440 5.490 ;
        RECT 1.315 3.845 1.545 4.590 ;
        RECT 6.040 3.800 6.270 4.590 ;
        RECT 8.130 3.880 8.360 4.590 ;
        RECT 10.170 3.880 10.400 4.590 ;
        RECT 12.210 3.090 12.440 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 13.870 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 13.870 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.070 ;
        RECT 5.985 0.450 6.325 0.635 ;
        RECT 8.280 0.450 8.510 0.690 ;
        RECT 10.520 0.450 10.750 1.160 ;
        RECT 12.760 0.450 12.990 1.540 ;
        RECT 0.000 -0.450 13.440 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 2.925 4.130 5.810 4.360 ;
        RECT 0.295 3.320 0.525 3.900 ;
        RECT 0.295 3.090 1.480 3.320 ;
        RECT 2.925 3.090 3.155 4.130 ;
        RECT 1.250 2.060 1.480 3.090 ;
        RECT 3.365 2.520 3.595 2.755 ;
        RECT 1.860 2.290 3.595 2.520 ;
        RECT 1.860 2.060 2.090 2.290 ;
        RECT 3.945 2.060 4.175 3.900 ;
        RECT 1.250 1.830 2.090 2.060 ;
        RECT 3.090 1.830 4.175 2.060 ;
        RECT 1.250 1.540 1.480 1.830 ;
        RECT 0.245 1.310 1.480 1.540 ;
        RECT 0.245 0.730 0.475 1.310 ;
        RECT 2.485 0.960 2.715 1.540 ;
        RECT 3.090 1.135 3.320 1.830 ;
        RECT 4.405 1.600 4.635 4.130 ;
        RECT 5.020 3.110 5.250 3.900 ;
        RECT 5.580 3.570 5.810 4.130 ;
        RECT 7.110 3.570 7.345 4.150 ;
        RECT 5.580 3.340 7.345 3.570 ;
        RECT 5.020 2.880 6.760 3.110 ;
        RECT 3.550 1.370 4.635 1.600 ;
        RECT 6.530 1.595 6.760 2.880 ;
        RECT 7.115 2.735 7.345 3.340 ;
        RECT 7.115 2.505 11.075 2.735 ;
        RECT 4.865 1.365 6.760 1.595 ;
        RECT 8.720 1.850 10.265 2.110 ;
        RECT 8.720 1.270 8.950 1.850 ;
        RECT 7.235 1.135 8.950 1.270 ;
        RECT 3.090 1.040 8.950 1.135 ;
        RECT 3.090 0.960 7.445 1.040 ;
        RECT 2.485 0.905 7.445 0.960 ;
        RECT 2.485 0.730 3.315 0.905 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__invz_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__invz_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__invz_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.720 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 1.770 1.555 2.710 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.165 2.330 5.450 3.270 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.669600 ;
    PORT
      LAYER Metal1 ;
        RECT 12.215 3.155 12.455 4.190 ;
        RECT 14.255 3.155 14.485 4.190 ;
        RECT 16.295 3.155 16.525 4.195 ;
        RECT 18.335 3.155 18.805 4.195 ;
        RECT 12.215 2.925 18.805 3.155 ;
        RECT 18.315 1.595 18.805 2.925 ;
        RECT 12.165 1.215 19.115 1.595 ;
        RECT 12.165 1.210 14.635 1.215 ;
        RECT 12.165 0.680 12.395 1.210 ;
        RECT 14.405 0.680 14.635 1.210 ;
        RECT 16.645 1.210 19.115 1.215 ;
        RECT 16.645 0.680 16.875 1.210 ;
        RECT 18.885 0.680 19.115 1.210 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 20.720 5.490 ;
        RECT 1.905 3.420 2.135 4.590 ;
        RECT 4.675 4.350 4.905 4.590 ;
        RECT 6.715 4.350 6.945 4.590 ;
        RECT 8.755 3.380 8.985 4.590 ;
        RECT 10.995 3.880 11.225 4.590 ;
        RECT 13.235 3.385 13.465 4.590 ;
        RECT 15.275 3.385 15.505 4.590 ;
        RECT 17.315 3.385 17.545 4.590 ;
        RECT 19.355 3.380 19.585 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 21.150 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 21.150 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.020 ;
        RECT 4.270 0.450 4.610 0.635 ;
        RECT 6.510 0.450 6.850 0.635 ;
        RECT 8.805 0.450 9.035 1.490 ;
        RECT 11.045 0.450 11.275 1.490 ;
        RECT 13.285 0.450 13.515 0.980 ;
        RECT 15.525 0.450 15.755 0.980 ;
        RECT 17.765 0.450 17.995 0.980 ;
        RECT 20.005 0.450 20.235 1.490 ;
        RECT 0.000 -0.450 20.720 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.885 3.170 1.115 4.190 ;
        RECT 7.735 4.120 7.965 4.190 ;
        RECT 2.925 3.890 7.965 4.120 ;
        RECT 2.925 3.380 3.155 3.890 ;
        RECT 0.885 3.150 2.725 3.170 ;
        RECT 0.885 2.940 3.650 3.150 ;
        RECT 2.630 2.425 3.650 2.940 ;
        RECT 2.630 2.110 2.860 2.425 ;
        RECT 1.805 1.880 2.860 2.110 ;
        RECT 3.945 2.055 4.175 3.660 ;
        RECT 1.805 1.490 2.035 1.880 ;
        RECT 3.090 1.825 4.175 2.055 ;
        RECT 3.090 1.490 3.320 1.825 ;
        RECT 4.405 1.595 4.635 3.890 ;
        RECT 5.695 2.710 5.925 3.660 ;
        RECT 5.695 2.480 7.385 2.710 ;
        RECT 7.155 1.595 7.385 2.480 ;
        RECT 7.735 2.695 7.965 3.890 ;
        RECT 9.875 2.695 10.105 4.190 ;
        RECT 7.735 2.405 17.195 2.695 ;
        RECT 0.245 1.260 2.035 1.490 ;
        RECT 0.245 0.680 0.475 1.260 ;
        RECT 2.485 1.135 3.320 1.490 ;
        RECT 3.550 1.365 4.635 1.595 ;
        RECT 5.390 1.365 7.385 1.595 ;
        RECT 7.745 1.825 17.535 2.055 ;
        RECT 7.745 1.135 7.975 1.825 ;
        RECT 2.485 0.905 7.975 1.135 ;
        RECT 2.485 0.680 2.715 0.905 ;
        RECT 7.630 0.855 7.975 0.905 ;
        RECT 9.925 0.840 10.155 1.825 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__invz_8

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__invz_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__invz_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 29.120 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 0.970 2.710 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.076000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.570 1.785 6.010 3.270 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 10.274400 ;
    PORT
      LAYER Metal1 ;
        RECT 16.140 3.490 16.370 4.280 ;
        RECT 18.280 3.490 18.510 4.280 ;
        RECT 20.520 3.490 20.750 4.280 ;
        RECT 22.660 3.490 22.890 4.280 ;
        RECT 24.700 3.490 24.930 4.280 ;
        RECT 26.735 3.490 26.970 4.280 ;
        RECT 16.140 3.010 26.970 3.490 ;
        RECT 26.450 1.595 26.980 3.010 ;
        RECT 16.090 0.895 27.520 1.595 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 29.120 5.490 ;
        RECT 1.830 3.470 2.060 4.590 ;
        RECT 6.030 4.510 6.260 4.590 ;
        RECT 8.510 4.510 8.740 4.590 ;
        RECT 10.770 3.950 11.000 4.590 ;
        RECT 12.810 3.470 13.040 4.590 ;
        RECT 14.920 3.880 15.150 4.590 ;
        RECT 17.160 3.960 17.390 4.590 ;
        RECT 19.400 3.940 19.630 4.590 ;
        RECT 21.640 3.940 21.870 4.590 ;
        RECT 23.680 3.940 23.910 4.590 ;
        RECT 25.720 3.940 25.950 4.590 ;
        RECT 27.760 3.470 27.990 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 29.550 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 29.550 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.070 ;
        RECT 5.955 0.450 6.295 0.635 ;
        RECT 8.195 0.450 8.535 0.635 ;
        RECT 10.490 0.450 10.720 1.540 ;
        RECT 12.730 0.450 12.960 1.540 ;
        RECT 14.970 0.450 15.200 1.540 ;
        RECT 17.155 0.450 17.495 0.635 ;
        RECT 19.395 0.450 19.735 0.635 ;
        RECT 21.635 0.450 21.975 0.635 ;
        RECT 23.875 0.450 24.215 0.635 ;
        RECT 26.115 0.450 26.455 0.635 ;
        RECT 28.410 0.450 28.640 1.540 ;
        RECT 0.000 -0.450 29.120 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.810 3.170 1.040 4.280 ;
        RECT 2.850 4.050 9.980 4.280 ;
        RECT 2.850 3.470 3.080 4.050 ;
        RECT 0.810 2.940 3.575 3.170 ;
        RECT 1.805 2.480 3.575 2.940 ;
        RECT 1.805 1.540 2.035 2.480 ;
        RECT 3.870 2.055 4.100 3.820 ;
        RECT 3.090 1.825 4.100 2.055 ;
        RECT 0.245 1.310 2.035 1.540 ;
        RECT 0.245 0.730 0.475 1.310 ;
        RECT 2.485 1.095 2.715 1.540 ;
        RECT 3.090 1.095 3.320 1.825 ;
        RECT 4.330 1.595 4.560 4.050 ;
        RECT 4.790 3.590 7.500 3.820 ;
        RECT 4.790 3.010 5.020 3.590 ;
        RECT 7.270 2.525 7.500 3.590 ;
        RECT 9.750 2.735 9.980 4.050 ;
        RECT 11.790 2.735 12.020 4.280 ;
        RECT 13.830 2.735 14.060 4.280 ;
        RECT 7.270 2.230 8.975 2.525 ;
        RECT 9.750 2.505 25.570 2.735 ;
        RECT 3.550 1.365 4.560 1.595 ;
        RECT 8.690 1.555 8.975 2.230 ;
        RECT 4.835 1.325 8.975 1.555 ;
        RECT 9.430 1.825 25.940 2.055 ;
        RECT 9.430 1.095 9.660 1.825 ;
        RECT 2.485 0.865 9.660 1.095 ;
        RECT 2.485 0.730 2.715 0.865 ;
        RECT 9.315 0.815 9.660 0.865 ;
        RECT 11.610 0.840 11.840 1.825 ;
        RECT 13.850 0.840 14.080 1.825 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__invz_12

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__invz_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__invz_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 36.960 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.815 1.850 1.155 2.275 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.768000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.065 2.030 7.710 2.605 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 14.329200 ;
    PORT
      LAYER Metal1 ;
        RECT 19.405 3.365 19.635 4.120 ;
        RECT 21.545 3.365 21.775 4.120 ;
        RECT 23.785 3.365 24.015 4.120 ;
        RECT 26.025 3.365 26.255 4.120 ;
        RECT 28.265 3.365 28.495 4.120 ;
        RECT 30.505 3.365 30.735 4.120 ;
        RECT 32.745 3.365 32.975 4.120 ;
        RECT 35.085 3.365 35.315 4.120 ;
        RECT 19.405 2.965 35.315 3.365 ;
        RECT 34.835 1.595 35.315 2.965 ;
        RECT 19.405 0.895 35.315 1.595 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 36.960 5.490 ;
        RECT 1.905 3.310 2.135 4.590 ;
        RECT 4.665 4.350 4.895 4.590 ;
        RECT 6.805 4.350 7.035 4.590 ;
        RECT 9.045 3.310 9.275 4.590 ;
        RECT 11.285 3.310 11.515 4.590 ;
        RECT 13.525 3.310 13.755 4.590 ;
        RECT 15.765 3.310 15.995 4.590 ;
        RECT 18.185 3.880 18.415 4.590 ;
        RECT 20.425 3.745 20.655 4.590 ;
        RECT 22.665 3.745 22.895 4.590 ;
        RECT 24.905 3.745 25.135 4.590 ;
        RECT 27.145 3.745 27.375 4.590 ;
        RECT 29.385 3.745 29.615 4.590 ;
        RECT 31.625 3.745 31.855 4.590 ;
        RECT 33.865 3.745 34.095 4.590 ;
        RECT 36.105 3.310 36.335 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 37.390 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 37.390 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.160 ;
        RECT 4.610 0.450 4.950 0.640 ;
        RECT 6.850 0.450 7.190 0.640 ;
        RECT 9.090 0.450 9.430 0.640 ;
        RECT 11.385 0.450 11.615 1.455 ;
        RECT 13.625 0.450 13.855 1.490 ;
        RECT 15.865 0.450 16.095 1.490 ;
        RECT 18.285 0.450 18.515 1.490 ;
        RECT 20.470 0.450 20.810 0.665 ;
        RECT 22.710 0.450 23.050 0.665 ;
        RECT 24.950 0.450 25.290 0.665 ;
        RECT 27.190 0.450 27.530 0.665 ;
        RECT 29.430 0.450 29.770 0.665 ;
        RECT 31.670 0.450 32.010 0.665 ;
        RECT 33.910 0.450 34.250 0.665 ;
        RECT 36.205 0.450 36.435 1.490 ;
        RECT 0.000 -0.450 36.960 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.885 2.735 1.115 4.120 ;
        RECT 2.925 3.890 8.815 4.120 ;
        RECT 2.925 3.310 3.155 3.890 ;
        RECT 0.885 2.505 3.650 2.735 ;
        RECT 1.805 1.620 2.035 2.505 ;
        RECT 3.945 2.095 4.175 3.650 ;
        RECT 0.245 1.390 2.035 1.620 ;
        RECT 3.090 1.865 4.175 2.095 ;
        RECT 3.090 1.490 3.320 1.865 ;
        RECT 4.405 1.595 4.635 3.890 ;
        RECT 5.730 3.310 8.310 3.650 ;
        RECT 8.080 2.620 8.310 3.310 ;
        RECT 8.585 3.080 8.815 3.890 ;
        RECT 10.165 3.080 10.395 4.120 ;
        RECT 12.405 3.080 12.635 4.120 ;
        RECT 14.645 3.080 14.875 4.120 ;
        RECT 17.065 3.080 17.295 4.120 ;
        RECT 8.585 2.850 17.295 3.080 ;
        RECT 17.065 2.735 17.295 2.850 ;
        RECT 8.080 2.305 16.450 2.620 ;
        RECT 17.065 2.505 33.700 2.735 ;
        RECT 8.080 1.600 8.310 2.305 ;
        RECT 18.610 2.075 33.730 2.095 ;
        RECT 0.245 0.680 0.475 1.390 ;
        RECT 2.485 1.135 3.320 1.490 ;
        RECT 3.550 1.365 4.635 1.595 ;
        RECT 5.730 1.370 8.310 1.600 ;
        RECT 10.270 1.865 33.730 2.075 ;
        RECT 10.270 1.750 18.800 1.865 ;
        RECT 10.270 1.135 10.500 1.750 ;
        RECT 2.485 0.905 10.500 1.135 ;
        RECT 2.485 0.680 2.715 0.905 ;
        RECT 10.265 0.680 10.500 0.905 ;
        RECT 12.505 0.680 12.735 1.750 ;
        RECT 14.745 0.680 14.975 1.750 ;
        RECT 17.165 0.680 17.395 1.750 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__invz_16

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__latq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.200 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.065 1.210 4.330 2.150 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.575 1.015 2.710 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.605 0.680 9.930 4.080 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 11.200 5.490 ;
        RECT 1.365 3.270 1.595 4.590 ;
        RECT 3.485 3.270 3.715 4.590 ;
        RECT 7.465 3.270 7.695 4.590 ;
        RECT 10.625 3.270 10.855 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 11.630 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 11.630 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 0.895 ;
        RECT 3.385 0.450 3.615 1.020 ;
        RECT 7.765 0.450 7.995 0.885 ;
        RECT 10.725 0.450 10.955 1.490 ;
        RECT 0.000 -0.450 11.200 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.270 0.575 4.080 ;
        RECT 0.245 1.345 0.475 3.270 ;
        RECT 2.665 2.610 2.895 4.080 ;
        RECT 5.245 3.410 5.475 4.080 ;
        RECT 5.245 3.180 6.215 3.410 ;
        RECT 5.525 2.610 5.755 2.950 ;
        RECT 2.665 2.380 5.755 2.610 ;
        RECT 2.085 1.355 2.315 1.915 ;
        RECT 1.085 1.345 2.315 1.355 ;
        RECT 0.245 1.125 2.315 1.345 ;
        RECT 0.245 1.115 1.155 1.125 ;
        RECT 0.245 0.680 0.475 1.115 ;
        RECT 2.665 0.680 2.895 2.380 ;
        RECT 4.665 1.575 4.895 2.380 ;
        RECT 5.985 1.345 6.215 3.180 ;
        RECT 8.485 2.375 8.735 4.080 ;
        RECT 7.085 2.365 8.735 2.375 ;
        RECT 7.085 2.145 9.115 2.365 ;
        RECT 7.085 1.575 7.315 2.145 ;
        RECT 8.205 1.345 8.435 1.915 ;
        RECT 5.985 1.225 8.435 1.345 ;
        RECT 5.345 1.115 8.435 1.225 ;
        RECT 5.345 0.885 6.190 1.115 ;
        RECT 8.665 0.975 9.115 2.145 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latq_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__latq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.320 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.065 1.210 4.330 2.150 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.575 1.015 2.710 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.675 1.590 11.050 4.235 ;
        RECT 10.230 1.210 11.050 1.590 ;
        RECT 10.725 0.680 11.050 1.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 12.320 5.490 ;
        RECT 1.365 3.425 1.595 4.590 ;
        RECT 3.485 3.425 3.715 4.590 ;
        RECT 7.465 3.425 7.695 4.590 ;
        RECT 9.655 3.425 9.885 4.590 ;
        RECT 11.695 3.425 11.925 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 12.750 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.750 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 0.895 ;
        RECT 3.385 0.450 3.615 1.020 ;
        RECT 7.765 0.450 7.995 0.885 ;
        RECT 9.605 0.450 9.835 1.490 ;
        RECT 11.845 0.450 12.075 1.490 ;
        RECT 0.000 -0.450 12.320 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.425 0.575 4.235 ;
        RECT 0.245 1.345 0.475 3.425 ;
        RECT 2.665 2.610 2.895 4.235 ;
        RECT 5.245 3.410 5.475 4.235 ;
        RECT 5.245 3.180 6.215 3.410 ;
        RECT 5.525 2.610 5.755 2.950 ;
        RECT 2.665 2.380 5.755 2.610 ;
        RECT 2.085 1.355 2.315 1.915 ;
        RECT 1.085 1.345 2.315 1.355 ;
        RECT 0.245 1.125 2.315 1.345 ;
        RECT 0.245 1.115 1.155 1.125 ;
        RECT 0.245 0.680 0.475 1.115 ;
        RECT 2.665 0.680 2.895 2.380 ;
        RECT 4.665 1.575 4.895 2.380 ;
        RECT 5.985 1.345 6.215 3.180 ;
        RECT 8.485 2.375 8.735 4.235 ;
        RECT 7.085 2.365 8.735 2.375 ;
        RECT 7.085 2.145 9.115 2.365 ;
        RECT 7.085 1.575 7.315 2.145 ;
        RECT 8.205 1.345 8.435 1.915 ;
        RECT 5.985 1.315 8.435 1.345 ;
        RECT 5.345 1.115 8.435 1.315 ;
        RECT 5.345 0.975 6.100 1.115 ;
        RECT 8.665 0.975 9.115 2.145 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latq_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__latq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.680 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.070 1.210 4.330 2.150 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 1.020 2.710 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 11.010 2.150 11.240 4.065 ;
        RECT 11.010 1.920 11.610 2.150 ;
        RECT 11.310 1.440 11.610 1.920 ;
        RECT 13.050 1.490 13.280 4.065 ;
        RECT 13.050 1.440 13.780 1.490 ;
        RECT 11.310 1.210 13.780 1.440 ;
        RECT 11.310 0.680 11.540 1.210 ;
        RECT 13.550 0.680 13.780 1.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 15.680 5.490 ;
        RECT 1.370 3.255 1.600 4.590 ;
        RECT 3.790 3.255 4.020 4.590 ;
        RECT 7.770 3.255 8.000 4.590 ;
        RECT 9.810 3.255 10.040 4.590 ;
        RECT 12.030 3.255 12.260 4.590 ;
        RECT 14.070 3.255 14.300 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 16.110 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 16.110 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.370 0.450 1.600 1.020 ;
        RECT 3.390 0.450 3.620 1.020 ;
        RECT 7.770 0.450 8.000 1.020 ;
        RECT 10.010 0.450 10.240 1.020 ;
        RECT 12.430 0.450 12.660 0.980 ;
        RECT 14.670 0.450 14.900 1.490 ;
        RECT 0.000 -0.450 15.680 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.250 3.255 0.580 4.065 ;
        RECT 0.250 1.540 0.480 3.255 ;
        RECT 2.570 2.720 2.800 4.065 ;
        RECT 5.550 3.180 5.780 4.065 ;
        RECT 5.550 2.950 6.520 3.180 ;
        RECT 2.570 2.380 6.060 2.720 ;
        RECT 1.990 1.540 2.220 2.150 ;
        RECT 0.250 1.310 2.220 1.540 ;
        RECT 0.250 0.680 0.480 1.310 ;
        RECT 2.570 0.680 2.900 2.380 ;
        RECT 4.670 1.810 4.900 2.380 ;
        RECT 6.290 1.020 6.520 2.950 ;
        RECT 8.790 2.610 9.120 4.065 ;
        RECT 7.330 2.380 9.120 2.610 ;
        RECT 7.330 1.810 7.560 2.380 ;
        RECT 8.210 1.480 8.440 2.150 ;
        RECT 5.350 0.910 6.520 1.020 ;
        RECT 7.310 1.250 8.440 1.480 ;
        RECT 7.310 0.910 7.540 1.250 ;
        RECT 5.350 0.680 7.540 0.910 ;
        RECT 8.890 0.680 9.120 2.380 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latq_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__latrnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latrnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.880 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 1.770 3.295 2.710 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.084000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.965 2.440 5.500 2.670 ;
        RECT 0.705 1.540 0.970 2.295 ;
        RECT 3.675 1.725 4.135 2.295 ;
        RECT 4.965 1.725 5.195 2.440 ;
        RECT 3.675 1.540 5.195 1.725 ;
        RECT 0.705 1.495 5.195 1.540 ;
        RECT 0.705 1.310 3.905 1.495 ;
        RECT 0.705 1.210 0.970 1.310 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.340000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.455 2.710 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 11.910 0.845 12.355 4.360 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 12.880 5.490 ;
        RECT 1.265 3.550 1.495 4.590 ;
        RECT 3.025 3.860 3.255 4.590 ;
        RECT 6.630 3.550 6.860 4.590 ;
        RECT 9.215 3.550 9.445 4.590 ;
        RECT 11.055 3.875 11.285 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 13.310 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 13.310 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.450 1.650 1.080 ;
        RECT 7.145 0.450 7.375 1.135 ;
        RECT 9.165 0.450 9.395 1.135 ;
        RECT 11.005 0.450 11.235 1.605 ;
        RECT 0.000 -0.450 12.880 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.170 0.475 4.360 ;
        RECT 2.005 3.630 2.235 4.360 ;
        RECT 4.785 4.130 5.960 4.360 ;
        RECT 4.785 3.630 5.015 4.130 ;
        RECT 2.005 3.400 5.015 3.630 ;
        RECT 0.245 2.940 4.735 3.170 ;
        RECT 0.245 0.795 0.475 2.940 ;
        RECT 4.505 1.955 4.735 2.940 ;
        RECT 5.730 1.725 5.960 4.130 ;
        RECT 7.830 2.755 8.240 4.360 ;
        RECT 6.190 2.525 8.240 2.755 ;
        RECT 6.190 1.955 6.420 2.525 ;
        RECT 8.010 2.295 8.240 2.525 ;
        RECT 7.550 1.765 7.780 2.295 ;
        RECT 8.010 2.065 9.835 2.295 ;
        RECT 6.550 1.725 7.780 1.765 ;
        RECT 5.730 1.535 7.780 1.725 ;
        RECT 8.445 1.955 9.835 2.065 ;
        RECT 10.235 2.260 10.465 4.360 ;
        RECT 10.235 2.030 11.620 2.260 ;
        RECT 5.730 1.495 6.680 1.535 ;
        RECT 6.450 1.135 6.680 1.495 ;
        RECT 4.345 0.795 6.680 1.135 ;
        RECT 8.445 0.795 8.675 1.955 ;
        RECT 10.235 1.225 10.515 2.030 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latrnq_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__latrnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latrnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.000 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 1.770 3.260 2.710 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.084000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.770 2.765 5.380 2.995 ;
        RECT 4.770 2.150 5.000 2.765 ;
        RECT 0.895 1.835 1.600 2.065 ;
        RECT 1.370 1.540 1.600 1.835 ;
        RECT 4.070 1.780 5.000 2.150 ;
        RECT 4.070 1.540 4.330 1.780 ;
        RECT 1.370 1.310 4.330 1.540 ;
        RECT 4.070 1.210 4.330 1.310 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.340000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 2.065 2.090 2.710 ;
        RECT 1.830 1.770 2.475 2.065 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.355 0.845 12.730 4.360 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 14.000 5.490 ;
        RECT 1.390 3.550 1.620 4.590 ;
        RECT 3.130 3.860 3.360 4.590 ;
        RECT 6.650 3.690 6.880 4.590 ;
        RECT 9.420 3.550 9.650 4.590 ;
        RECT 11.335 3.880 11.565 4.590 ;
        RECT 13.375 3.880 13.605 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 14.430 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.430 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.435 0.450 1.775 1.080 ;
        RECT 7.350 0.450 7.580 1.135 ;
        RECT 9.370 0.450 9.600 1.135 ;
        RECT 11.285 0.450 11.515 1.605 ;
        RECT 13.525 0.450 13.755 1.605 ;
        RECT 0.000 -0.450 14.000 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.370 3.170 0.600 4.360 ;
        RECT 2.110 3.630 2.340 4.030 ;
        RECT 4.890 3.800 5.840 4.030 ;
        RECT 4.890 3.630 5.120 3.800 ;
        RECT 2.110 3.400 5.120 3.630 ;
        RECT 0.370 2.940 4.540 3.170 ;
        RECT 0.370 0.795 0.600 2.940 ;
        RECT 4.310 2.380 4.540 2.940 ;
        RECT 5.610 1.135 5.840 3.800 ;
        RECT 7.895 2.580 8.440 4.360 ;
        RECT 7.290 2.350 8.440 2.580 ;
        RECT 7.290 2.120 7.520 2.350 ;
        RECT 8.210 2.120 8.440 2.350 ;
        RECT 6.070 1.890 7.520 2.120 ;
        RECT 6.070 1.780 6.300 1.890 ;
        RECT 7.750 1.595 7.980 2.120 ;
        RECT 4.550 1.025 5.840 1.135 ;
        RECT 6.440 1.365 7.980 1.595 ;
        RECT 8.210 1.780 10.040 2.120 ;
        RECT 10.440 2.065 10.670 4.360 ;
        RECT 10.440 1.835 12.010 2.065 ;
        RECT 6.440 1.025 6.670 1.365 ;
        RECT 4.550 0.795 6.670 1.025 ;
        RECT 8.210 0.795 8.880 1.780 ;
        RECT 10.440 1.225 10.720 1.835 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latrnq_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__latrnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latrnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.920 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.500 1.770 3.770 2.720 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.084000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.740 1.540 0.970 2.720 ;
        RECT 4.120 1.585 4.350 2.720 ;
        RECT 5.640 2.150 5.870 2.720 ;
        RECT 5.190 1.920 5.870 2.150 ;
        RECT 5.190 1.585 5.450 1.920 ;
        RECT 4.120 1.540 5.450 1.585 ;
        RECT 0.740 1.355 5.450 1.540 ;
        RECT 0.740 1.310 4.260 1.355 ;
        RECT 5.190 1.210 5.450 1.355 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.340000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.390 1.770 2.650 2.720 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.035 3.645 14.265 4.360 ;
        RECT 16.075 3.645 16.305 4.360 ;
        RECT 14.035 3.415 16.305 3.645 ;
        RECT 14.035 2.055 14.410 3.415 ;
        RECT 14.035 1.825 16.555 2.055 ;
        RECT 14.035 0.785 14.410 1.825 ;
        RECT 16.325 0.785 16.555 1.825 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.920 5.490 ;
        RECT 1.320 3.550 1.550 4.590 ;
        RECT 3.240 3.870 3.470 4.590 ;
        RECT 7.610 3.700 7.840 4.590 ;
        RECT 9.880 3.550 10.110 4.590 ;
        RECT 12.070 3.550 12.300 4.590 ;
        RECT 13.015 3.875 13.245 4.590 ;
        RECT 15.055 3.875 15.285 4.590 ;
        RECT 17.095 3.875 17.325 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 18.350 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 18.350 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.345 0.450 1.685 1.070 ;
        RECT 7.740 0.450 7.970 1.125 ;
        RECT 9.980 0.450 10.210 1.125 ;
        RECT 12.220 0.450 12.450 1.125 ;
        RECT 12.965 0.450 13.195 1.595 ;
        RECT 15.205 0.450 15.435 1.595 ;
        RECT 17.445 0.450 17.675 1.595 ;
        RECT 0.000 -0.450 17.920 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.280 3.180 0.530 4.360 ;
        RECT 2.220 3.640 2.450 4.040 ;
        RECT 5.320 3.810 6.330 4.040 ;
        RECT 5.320 3.640 5.550 3.810 ;
        RECT 2.220 3.410 5.550 3.640 ;
        RECT 0.280 2.950 5.270 3.180 ;
        RECT 0.280 0.785 0.510 2.950 ;
        RECT 5.040 2.380 5.270 2.950 ;
        RECT 6.100 2.150 6.330 3.810 ;
        RECT 8.810 3.180 9.040 4.360 ;
        RECT 11.050 3.550 11.325 4.360 ;
        RECT 7.170 2.950 10.840 3.180 ;
        RECT 7.170 2.380 7.400 2.950 ;
        RECT 8.230 2.150 8.460 2.720 ;
        RECT 6.100 1.920 8.460 2.150 ;
        RECT 4.580 0.980 4.810 1.125 ;
        RECT 6.100 0.980 6.330 1.920 ;
        RECT 4.580 0.750 6.330 0.980 ;
        RECT 8.860 0.785 9.090 2.950 ;
        RECT 10.610 2.380 10.840 2.950 ;
        RECT 11.095 2.665 11.325 3.550 ;
        RECT 11.095 2.435 13.740 2.665 ;
        RECT 11.095 0.785 11.330 2.435 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latrnq_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__latrsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latrsnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.440 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 1.770 3.335 2.710 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.084000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 2.275 1.600 2.505 ;
        RECT 1.370 1.540 1.600 2.275 ;
        RECT 3.945 2.150 4.175 2.560 ;
        RECT 5.265 2.150 5.495 2.560 ;
        RECT 3.945 1.770 5.495 2.150 ;
        RECT 3.945 1.540 4.175 1.770 ;
        RECT 1.370 1.310 4.175 1.540 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.340000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.495 2.710 ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.550 1.770 8.875 2.710 ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.425 0.845 12.735 4.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 13.440 5.490 ;
        RECT 1.265 3.400 1.495 4.590 ;
        RECT 3.065 3.890 3.295 4.590 ;
        RECT 6.645 3.890 6.875 4.590 ;
        RECT 8.925 3.400 9.155 4.590 ;
        RECT 11.225 3.430 11.455 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 13.870 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 13.870 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.080 ;
        RECT 7.130 0.450 7.470 1.075 ;
        RECT 11.385 0.450 11.615 1.165 ;
        RECT 0.000 -0.450 13.440 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.170 0.475 4.210 ;
        RECT 2.045 3.630 2.275 4.210 ;
        RECT 4.825 3.630 5.055 4.210 ;
        RECT 2.045 3.400 7.315 3.630 ;
        RECT 0.245 2.940 4.775 3.170 ;
        RECT 7.085 3.020 7.315 3.400 ;
        RECT 0.245 0.790 0.475 2.940 ;
        RECT 4.545 2.380 4.775 2.940 ;
        RECT 5.725 2.790 7.315 3.020 ;
        RECT 7.905 3.170 8.135 4.210 ;
        RECT 10.205 3.200 10.435 4.210 ;
        RECT 7.905 2.940 9.555 3.170 ;
        RECT 10.205 2.970 11.915 3.200 ;
        RECT 5.725 1.130 5.955 2.790 ;
        RECT 9.325 2.560 9.555 2.940 ;
        RECT 6.185 1.540 6.415 2.560 ;
        RECT 9.325 2.220 10.715 2.560 ;
        RECT 9.325 1.540 9.555 2.220 ;
        RECT 11.685 1.655 11.915 2.970 ;
        RECT 6.185 1.310 9.555 1.540 ;
        RECT 10.045 1.425 11.915 1.655 ;
        RECT 10.045 1.315 10.275 1.425 ;
        RECT 4.385 0.790 5.955 1.130 ;
        RECT 9.325 0.790 9.555 1.310 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latrsnq_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__latrsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latrsnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.560 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.020000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 2.505 3.210 3.270 ;
        RECT 2.950 2.275 3.810 2.505 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.322000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.925 1.990 1.155 2.560 ;
        RECT 4.070 1.990 4.755 2.710 ;
        RECT 5.885 1.990 6.115 2.560 ;
        RECT 0.925 1.760 6.115 1.990 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.440000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 2.275 2.650 2.710 ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.302000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.110 1.770 9.535 2.710 ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.945 2.150 13.175 4.310 ;
        RECT 12.470 1.210 13.175 2.150 ;
        RECT 12.945 0.790 13.175 1.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 14.560 5.490 ;
        RECT 1.365 3.880 1.595 4.590 ;
        RECT 3.425 4.420 3.655 4.590 ;
        RECT 7.565 3.500 7.795 4.590 ;
        RECT 9.985 3.880 10.215 4.590 ;
        RECT 11.825 3.880 12.055 4.590 ;
        RECT 14.065 3.880 14.295 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 14.990 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.990 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.585 0.450 1.815 1.130 ;
        RECT 7.605 0.450 7.835 1.130 ;
        RECT 11.825 0.450 12.055 1.530 ;
        RECT 14.065 0.450 14.295 1.600 ;
        RECT 0.000 -0.450 14.560 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.650 0.475 4.310 ;
        RECT 2.085 4.190 2.315 4.220 ;
        RECT 5.605 4.190 5.835 4.310 ;
        RECT 2.085 3.960 5.835 4.190 ;
        RECT 2.085 3.880 2.315 3.960 ;
        RECT 2.490 3.650 5.355 3.730 ;
        RECT 0.245 3.500 5.355 3.650 ;
        RECT 0.245 3.420 2.665 3.500 ;
        RECT 0.245 0.790 0.695 3.420 ;
        RECT 5.125 2.220 5.355 3.500 ;
        RECT 5.605 3.020 5.835 3.960 ;
        RECT 8.865 3.650 9.095 4.310 ;
        RECT 10.705 3.650 10.935 4.310 ;
        RECT 8.865 3.420 9.995 3.650 ;
        RECT 10.705 3.420 12.240 3.650 ;
        RECT 5.605 2.790 8.235 3.020 ;
        RECT 6.345 1.130 6.575 2.790 ;
        RECT 7.135 1.990 7.365 2.560 ;
        RECT 8.005 2.220 8.235 2.790 ;
        RECT 9.765 2.560 9.995 3.420 ;
        RECT 9.765 2.220 11.375 2.560 ;
        RECT 7.135 1.760 8.210 1.990 ;
        RECT 7.980 1.540 8.210 1.760 ;
        RECT 9.765 1.540 9.995 2.220 ;
        RECT 12.010 1.990 12.240 3.420 ;
        RECT 7.980 1.310 9.995 1.540 ;
        RECT 4.805 0.790 6.575 1.130 ;
        RECT 9.745 0.790 9.995 1.310 ;
        RECT 10.705 1.760 12.240 1.990 ;
        RECT 10.705 0.790 10.935 1.760 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latrsnq_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__latrsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latrsnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.360 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 2.195 3.210 2.710 ;
        RECT 2.950 1.770 3.500 2.195 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.084000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.525 2.875 5.370 3.105 ;
        RECT 1.830 2.195 2.090 2.710 ;
        RECT 0.970 1.965 2.090 2.195 ;
        RECT 4.525 2.120 4.755 2.875 ;
        RECT 1.830 1.540 2.090 1.965 ;
        RECT 4.055 1.890 4.755 2.120 ;
        RECT 4.055 1.540 4.285 1.890 ;
        RECT 1.830 1.310 4.285 1.540 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.340000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.375 1.770 2.650 2.710 ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.550 1.770 8.985 2.710 ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 13.265 3.650 13.495 4.290 ;
        RECT 15.305 3.650 15.535 4.290 ;
        RECT 13.265 3.420 15.535 3.650 ;
        RECT 13.515 2.150 13.745 3.420 ;
        RECT 13.515 1.920 15.530 2.150 ;
        RECT 13.515 0.845 13.745 1.920 ;
        RECT 15.270 1.655 15.530 1.920 ;
        RECT 15.270 1.210 15.985 1.655 ;
        RECT 15.755 0.845 15.985 1.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.360 5.490 ;
        RECT 1.305 3.480 1.535 4.590 ;
        RECT 3.045 4.120 3.275 4.590 ;
        RECT 6.565 3.480 6.795 4.590 ;
        RECT 8.785 3.650 9.015 4.590 ;
        RECT 10.205 3.880 10.435 4.590 ;
        RECT 12.245 3.880 12.475 4.590 ;
        RECT 14.285 3.880 14.515 4.590 ;
        RECT 16.325 3.880 16.555 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 17.790 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 17.790 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.460 0.450 1.800 1.080 ;
        RECT 7.240 0.450 7.580 1.080 ;
        RECT 10.155 0.450 10.385 1.165 ;
        RECT 12.395 0.450 12.625 1.165 ;
        RECT 14.635 0.450 14.865 1.165 ;
        RECT 16.875 0.450 17.105 1.165 ;
        RECT 0.000 -0.450 17.360 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.285 3.170 0.515 4.290 ;
        RECT 2.025 3.710 2.255 4.290 ;
        RECT 4.805 3.710 5.035 4.290 ;
        RECT 2.025 3.565 5.035 3.710 ;
        RECT 2.025 3.480 5.830 3.565 ;
        RECT 4.820 3.335 5.830 3.480 ;
        RECT 0.285 2.940 4.295 3.170 ;
        RECT 0.285 0.795 0.625 2.940 ;
        RECT 4.065 2.380 4.295 2.940 ;
        RECT 5.600 2.720 5.830 3.335 ;
        RECT 7.765 3.420 7.995 4.290 ;
        RECT 7.765 3.190 9.665 3.420 ;
        RECT 5.600 2.655 7.535 2.720 ;
        RECT 5.535 2.490 7.535 2.655 ;
        RECT 5.535 1.135 5.765 2.490 ;
        RECT 6.135 1.540 6.365 2.260 ;
        RECT 7.305 1.935 7.535 2.490 ;
        RECT 9.435 2.250 9.665 3.190 ;
        RECT 11.225 2.760 11.455 4.290 ;
        RECT 11.225 2.530 12.915 2.760 ;
        RECT 9.435 1.910 11.065 2.250 ;
        RECT 9.435 1.540 9.665 1.910 ;
        RECT 12.685 1.655 12.915 2.530 ;
        RECT 6.135 1.310 9.665 1.540 ;
        RECT 4.495 0.795 5.765 1.135 ;
        RECT 9.435 0.795 9.665 1.310 ;
        RECT 11.275 1.425 12.915 1.655 ;
        RECT 11.275 0.845 11.505 1.425 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latrsnq_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__latsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latsnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.760 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.210 2.270 2.160 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.084000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.390 3.295 2.620 ;
        RECT 0.710 1.770 1.015 2.390 ;
        RECT 3.065 2.090 3.295 2.390 ;
        RECT 3.690 2.090 4.030 3.200 ;
        RECT 3.065 1.830 4.030 2.090 ;
    END
  END E
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.870 1.210 7.210 2.160 ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.720 0.845 11.050 4.230 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 11.760 5.490 ;
        RECT 1.365 3.420 1.595 4.590 ;
        RECT 5.225 3.420 5.455 4.590 ;
        RECT 7.685 3.420 7.915 4.590 ;
        RECT 9.570 3.420 9.800 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 12.190 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.190 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.185 ;
        RECT 5.465 0.450 5.695 1.185 ;
        RECT 9.700 0.450 9.930 1.220 ;
        RECT 0.000 -0.450 11.760 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.190 0.575 4.230 ;
        RECT 3.305 4.000 4.490 4.230 ;
        RECT 3.305 3.420 3.535 4.000 ;
        RECT 0.245 2.850 2.955 3.190 ;
        RECT 0.245 0.845 0.475 2.850 ;
        RECT 4.260 1.185 4.490 4.000 ;
        RECT 6.665 2.675 6.895 4.230 ;
        RECT 8.500 3.205 8.730 4.230 ;
        RECT 8.500 2.975 9.485 3.205 ;
        RECT 5.625 2.620 6.895 2.675 ;
        RECT 5.625 2.445 7.835 2.620 ;
        RECT 5.625 2.215 5.855 2.445 ;
        RECT 6.745 2.390 7.835 2.445 ;
        RECT 7.605 2.215 7.835 2.390 ;
        RECT 4.785 1.875 5.855 2.215 ;
        RECT 6.085 1.645 6.315 2.215 ;
        RECT 3.505 1.075 4.490 1.185 ;
        RECT 5.005 1.415 6.315 1.645 ;
        RECT 7.605 1.875 9.025 2.215 ;
        RECT 9.255 1.935 9.485 2.975 ;
        RECT 10.140 1.935 10.370 2.215 ;
        RECT 5.005 1.075 5.235 1.415 ;
        RECT 3.505 0.845 5.235 1.075 ;
        RECT 7.605 0.845 7.835 1.875 ;
        RECT 9.255 1.790 10.370 1.935 ;
        RECT 9.240 1.705 10.370 1.790 ;
        RECT 9.240 1.225 9.470 1.705 ;
        RECT 8.355 0.885 9.470 1.225 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latsnq_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__latsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latsnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.320 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.210 2.090 2.335 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.084000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.235 3.090 4.080 3.320 ;
        RECT 3.235 2.795 3.465 3.090 ;
        RECT 0.925 2.565 3.465 2.795 ;
        RECT 0.925 1.995 1.155 2.565 ;
        RECT 2.950 2.050 3.465 2.565 ;
        RECT 2.950 1.770 3.210 2.050 ;
    END
  END E
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.870 1.770 7.155 2.710 ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.575 2.150 10.805 4.200 ;
        RECT 10.575 0.680 11.050 2.150 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 12.320 5.490 ;
        RECT 1.415 3.665 1.645 4.590 ;
        RECT 5.115 3.550 5.345 4.590 ;
        RECT 7.335 3.550 7.565 4.590 ;
        RECT 9.555 3.860 9.785 4.590 ;
        RECT 11.595 3.550 11.825 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 12.750 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.750 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.020 ;
        RECT 5.465 0.450 5.695 1.020 ;
        RECT 9.605 0.450 9.835 1.305 ;
        RECT 11.845 0.450 12.075 1.490 ;
        RECT 0.000 -0.450 12.320 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.365 0.625 4.360 ;
        RECT 3.355 4.130 4.540 4.360 ;
        RECT 3.355 3.550 3.585 4.130 ;
        RECT 0.245 3.025 3.005 3.365 ;
        RECT 0.245 0.680 0.475 3.025 ;
        RECT 4.310 1.765 4.540 4.130 ;
        RECT 6.315 3.170 6.545 4.200 ;
        RECT 8.535 3.630 8.765 4.210 ;
        RECT 8.535 3.400 10.225 3.630 ;
        RECT 5.025 2.940 9.205 3.170 ;
        RECT 5.025 1.995 5.255 2.940 ;
        RECT 5.735 1.765 5.965 2.335 ;
        RECT 8.975 2.225 9.205 2.940 ;
        RECT 3.505 1.535 5.965 1.765 ;
        RECT 7.605 1.995 9.205 2.225 ;
        RECT 3.505 0.680 3.735 1.535 ;
        RECT 7.605 0.680 7.835 1.995 ;
        RECT 9.995 1.765 10.225 3.400 ;
        RECT 8.485 1.535 10.225 1.765 ;
        RECT 8.485 0.680 8.715 1.535 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latsnq_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__latsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latsnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.680 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.245 1.210 2.650 2.150 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.084000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 2.945 4.195 3.270 ;
        RECT 3.510 2.610 3.770 2.945 ;
        RECT 1.785 2.380 3.770 2.610 ;
        RECT 1.785 2.150 2.015 2.380 ;
        RECT 0.945 1.920 2.015 2.150 ;
        RECT 2.880 2.330 3.770 2.380 ;
        RECT 2.880 1.920 3.220 2.330 ;
    END
  END E
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.870 1.770 7.230 2.710 ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 11.510 3.320 11.740 4.250 ;
        RECT 13.550 3.320 13.780 4.250 ;
        RECT 11.510 3.090 13.780 3.320 ;
        RECT 11.760 1.440 11.990 3.090 ;
        RECT 13.590 1.650 13.850 2.150 ;
        RECT 13.590 1.440 14.230 1.650 ;
        RECT 11.760 1.210 14.230 1.440 ;
        RECT 11.760 0.840 11.990 1.210 ;
        RECT 14.000 0.840 14.230 1.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 15.680 5.490 ;
        RECT 1.610 3.705 1.840 4.590 ;
        RECT 5.390 3.550 5.620 4.590 ;
        RECT 7.610 3.875 7.840 4.590 ;
        RECT 8.450 3.875 8.680 4.590 ;
        RECT 10.490 3.875 10.720 4.590 ;
        RECT 12.530 3.550 12.760 4.590 ;
        RECT 14.570 3.875 14.800 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 16.110 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 16.110 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.440 0.450 1.670 1.305 ;
        RECT 5.540 0.450 5.770 1.310 ;
        RECT 8.400 0.450 8.630 1.160 ;
        RECT 10.640 0.450 10.870 1.160 ;
        RECT 12.880 0.450 13.110 0.690 ;
        RECT 15.120 0.450 15.350 1.160 ;
        RECT 0.000 -0.450 15.680 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.590 3.180 0.820 4.360 ;
        RECT 3.630 4.130 4.655 4.360 ;
        RECT 3.630 3.550 3.860 4.130 ;
        RECT 0.590 2.890 3.280 3.180 ;
        RECT 0.320 2.840 3.280 2.890 ;
        RECT 0.320 2.660 0.815 2.840 ;
        RECT 0.320 0.880 0.550 2.660 ;
        RECT 4.425 1.770 4.655 4.130 ;
        RECT 6.590 3.170 6.820 4.250 ;
        RECT 6.590 3.135 9.070 3.170 ;
        RECT 5.100 2.940 9.070 3.135 ;
        RECT 5.100 2.905 6.715 2.940 ;
        RECT 5.100 2.000 5.330 2.905 ;
        RECT 6.000 1.770 6.230 2.310 ;
        RECT 3.580 1.540 6.230 1.770 ;
        RECT 8.840 1.650 9.070 2.940 ;
        RECT 3.580 0.970 3.810 1.540 ;
        RECT 7.680 1.420 9.070 1.650 ;
        RECT 9.470 2.280 9.700 4.250 ;
        RECT 9.470 1.940 11.300 2.280 ;
        RECT 7.680 0.840 7.910 1.420 ;
        RECT 9.470 0.840 9.750 1.940 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latsnq_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__mux2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__mux2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.853500 ;
    PORT
      LAYER Metal1 ;
        RECT 4.630 1.770 5.450 2.150 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.853500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.390 1.770 2.650 2.710 ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 2.705 6.035 3.270 ;
        RECT 3.225 2.475 6.035 2.705 ;
        RECT 3.225 1.380 3.455 2.475 ;
        RECT 5.750 1.770 6.035 2.475 ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 0.720 0.575 4.235 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.280 5.490 ;
        RECT 1.365 2.970 1.595 4.590 ;
        RECT 5.310 3.480 5.650 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 7.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.060 ;
        RECT 5.465 0.450 5.695 0.990 ;
        RECT 0.000 -0.450 7.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.930 3.545 3.835 3.775 ;
        RECT 1.930 2.055 2.160 3.545 ;
        RECT 3.605 2.965 3.835 3.545 ;
        RECT 0.870 1.825 2.160 2.055 ;
        RECT 1.930 1.005 2.160 1.825 ;
        RECT 3.945 1.540 4.175 2.110 ;
        RECT 6.385 1.540 6.815 3.775 ;
        RECT 3.945 1.310 6.815 1.540 ;
        RECT 1.930 0.775 3.790 1.005 ;
        RECT 6.585 0.720 6.815 1.310 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__mux2_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__mux2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__mux2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.400 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 1.770 6.570 2.150 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 1.770 3.255 2.710 ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.005 2.470 7.315 2.710 ;
        RECT 4.005 1.775 4.235 2.470 ;
        RECT 6.870 1.770 7.315 2.470 ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.729500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 0.680 1.595 4.360 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 8.400 5.490 ;
        RECT 0.295 3.550 0.525 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 6.645 3.550 6.875 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 8.830 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.830 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.020 ;
        RECT 6.645 0.450 6.875 1.020 ;
        RECT 0.000 -0.450 8.400 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 4.885 3.170 5.115 4.360 ;
        RECT 1.945 2.940 5.115 3.170 ;
        RECT 1.945 1.540 2.175 2.940 ;
        RECT 4.830 1.830 5.520 2.060 ;
        RECT 5.290 1.540 5.520 1.830 ;
        RECT 7.665 1.540 7.995 4.360 ;
        RECT 1.945 1.310 4.675 1.540 ;
        RECT 5.290 1.310 7.995 1.540 ;
        RECT 4.445 0.680 4.675 1.310 ;
        RECT 7.765 0.680 7.995 1.310 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__mux2_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__mux2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__mux2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.640 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.990 1.830 8.645 2.150 ;
        RECT 7.990 1.210 8.250 1.830 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.130 1.770 6.010 2.150 ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.300 2.470 9.430 2.700 ;
        RECT 6.300 1.775 6.530 2.470 ;
        RECT 9.050 2.060 9.430 2.470 ;
        RECT 9.050 1.830 9.665 2.060 ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.550500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.420 2.710 1.650 4.360 ;
        RECT 3.610 2.710 3.890 4.360 ;
        RECT 1.420 2.330 3.890 2.710 ;
        RECT 1.420 0.680 1.650 2.330 ;
        RECT 3.660 0.680 3.890 2.330 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 10.640 5.490 ;
        RECT 0.350 3.550 0.580 4.590 ;
        RECT 2.490 3.550 2.720 4.590 ;
        RECT 4.680 3.550 4.910 4.590 ;
        RECT 8.940 3.550 9.170 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 11.070 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 11.070 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 0.450 0.530 1.490 ;
        RECT 2.540 0.450 2.770 1.490 ;
        RECT 4.780 0.450 5.010 1.020 ;
        RECT 8.940 0.450 9.170 1.020 ;
        RECT 0.000 -0.450 10.640 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 7.180 3.160 7.410 4.360 ;
        RECT 4.670 2.930 7.410 3.160 ;
        RECT 4.670 2.115 4.900 2.930 ;
        RECT 4.240 1.775 4.900 2.115 ;
        RECT 7.125 1.830 7.760 2.060 ;
        RECT 4.670 1.540 4.900 1.775 ;
        RECT 4.670 1.310 6.970 1.540 ;
        RECT 6.740 0.680 6.970 1.310 ;
        RECT 7.530 0.980 7.760 1.830 ;
        RECT 9.960 1.480 10.290 4.360 ;
        RECT 8.480 1.250 10.290 1.480 ;
        RECT 8.480 0.980 8.710 1.250 ;
        RECT 7.530 0.750 8.710 0.980 ;
        RECT 10.060 0.680 10.290 1.250 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__mux2_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__mux4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__mux4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.360 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.853500 ;
    PORT
      LAYER Metal1 ;
        RECT 14.710 1.210 14.970 2.555 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.853500 ;
    PORT
      LAYER Metal1 ;
        RECT 11.350 1.770 11.610 2.710 ;
    END
  END I1
  PIN I2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.853500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 0.970 2.710 ;
    END
  END I2
  PIN I3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.853500 ;
    PORT
      LAYER Metal1 ;
        RECT 4.070 1.770 4.375 2.710 ;
    END
  END I3
  PIN S0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.560500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.390 1.900 2.650 2.995 ;
        RECT 2.390 1.670 3.210 1.900 ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.405 2.155 8.810 3.195 ;
        RECT 7.675 1.770 8.810 2.155 ;
    END
  END S1
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.003200 ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 2.330 6.255 3.175 ;
        RECT 6.025 1.590 6.255 2.330 ;
        RECT 5.750 1.210 6.255 1.590 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.360 5.490 ;
        RECT 0.295 3.440 0.525 4.590 ;
        RECT 4.725 3.865 4.955 4.590 ;
        RECT 10.935 3.440 11.165 4.590 ;
        RECT 15.015 3.440 15.245 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.280 17.790 5.470 ;
        RECT -0.430 2.265 0.430 2.280 ;
        RECT 16.930 2.265 17.790 2.280 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 4.745 2.265 6.455 2.280 ;
        RECT -0.430 -0.430 17.790 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.430 ;
        RECT 4.725 0.450 4.955 1.430 ;
        RECT 10.835 0.450 11.065 1.430 ;
        RECT 15.315 0.450 15.545 1.430 ;
        RECT 0.000 -0.450 17.360 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 1.090 1.595 4.170 ;
        RECT 2.665 3.940 4.495 4.170 ;
        RECT 2.665 3.455 2.895 3.940 ;
        RECT 1.930 3.225 2.895 3.455 ;
        RECT 3.605 3.355 3.915 3.695 ;
        RECT 4.265 3.635 4.495 3.940 ;
        RECT 6.805 3.635 7.035 4.170 ;
        RECT 4.265 3.405 7.035 3.635 ;
        RECT 6.755 3.360 7.035 3.405 ;
        RECT 1.930 1.375 2.160 3.225 ;
        RECT 1.930 1.145 2.770 1.375 ;
        RECT 3.605 1.090 3.835 3.355 ;
        RECT 5.290 1.790 5.575 2.130 ;
        RECT 5.290 0.925 5.520 1.790 ;
        RECT 6.755 1.155 6.985 3.360 ;
        RECT 7.825 2.615 8.055 4.170 ;
        RECT 8.845 4.005 10.705 4.235 ;
        RECT 8.845 3.425 9.270 4.005 ;
        RECT 7.215 2.385 8.055 2.615 ;
        RECT 7.215 0.925 7.445 2.385 ;
        RECT 9.040 1.430 9.270 3.425 ;
        RECT 9.915 2.315 10.145 3.695 ;
        RECT 10.475 3.210 10.705 4.005 ;
        RECT 11.395 3.940 13.305 4.170 ;
        RECT 11.395 3.210 11.625 3.940 ;
        RECT 10.475 2.980 11.625 3.210 ;
        RECT 7.875 0.925 8.105 1.345 ;
        RECT 8.995 1.090 9.270 1.430 ;
        RECT 9.500 1.090 10.145 2.315 ;
        RECT 11.955 1.090 12.185 3.695 ;
        RECT 12.975 1.090 13.305 3.940 ;
        RECT 13.995 3.475 14.225 4.250 ;
        RECT 13.675 3.245 14.225 3.475 ;
        RECT 13.675 1.375 13.905 3.245 ;
        RECT 16.035 3.015 16.265 4.170 ;
        RECT 14.135 2.785 16.665 3.015 ;
        RECT 14.135 2.215 14.365 2.785 ;
        RECT 13.675 1.145 14.480 1.375 ;
        RECT 16.435 1.090 16.665 2.785 ;
        RECT 5.290 0.695 8.105 0.925 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__mux4_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__mux4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__mux4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.040 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.120000 ;
    PORT
      LAYER Metal1 ;
        RECT 16.950 1.210 17.210 2.030 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.120000 ;
    PORT
      LAYER Metal1 ;
        RECT 13.590 1.770 13.850 2.390 ;
    END
  END I1
  PIN I2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.120000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.050 1.015 3.270 ;
    END
  END I2
  PIN I3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.120000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.625 2.050 4.890 2.710 ;
    END
  END I3
  PIN S0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.360000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.285 2.000 2.515 2.390 ;
        RECT 3.510 2.000 3.815 2.260 ;
        RECT 2.285 1.770 3.815 2.000 ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.240000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.600 2.150 10.830 2.830 ;
        RECT 9.560 1.770 10.830 2.150 ;
        RECT 9.560 1.690 9.790 1.770 ;
    END
  END S1
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.081600 ;
    PORT
      LAYER Metal1 ;
        RECT 6.310 1.200 6.755 3.380 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 19.040 5.490 ;
        RECT 0.250 3.080 0.480 4.590 ;
        RECT 5.285 4.070 5.515 4.590 ;
        RECT 7.545 3.080 7.775 4.590 ;
        RECT 13.000 3.080 13.230 4.590 ;
        RECT 17.340 3.080 17.570 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 19.470 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 19.470 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.540 ;
        RECT 5.405 0.450 5.635 1.540 ;
        RECT 7.645 0.450 7.875 1.540 ;
        RECT 12.960 0.450 13.190 1.540 ;
        RECT 17.440 0.450 17.670 1.540 ;
        RECT 0.000 -0.450 19.040 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 11.120 4.120 12.770 4.350 ;
        RECT 1.365 1.200 1.595 3.890 ;
        RECT 1.825 3.840 2.955 3.890 ;
        RECT 1.825 3.610 7.315 3.840 ;
        RECT 1.825 1.485 2.055 3.610 ;
        RECT 2.725 3.080 2.955 3.610 ;
        RECT 4.045 1.845 4.275 3.380 ;
        RECT 7.085 2.850 7.315 3.610 ;
        RECT 8.640 3.080 9.005 3.890 ;
        RECT 9.235 3.660 10.180 3.890 ;
        RECT 8.640 2.850 8.870 3.080 ;
        RECT 7.085 2.620 8.870 2.850 ;
        RECT 7.105 2.000 7.335 2.390 ;
        RECT 4.045 1.615 4.515 1.845 ;
        RECT 7.105 1.770 8.410 2.000 ;
        RECT 1.825 1.255 3.450 1.485 ;
        RECT 4.285 1.200 4.515 1.615 ;
        RECT 8.180 0.980 8.410 1.770 ;
        RECT 8.640 1.210 8.870 2.620 ;
        RECT 9.235 2.570 9.465 3.660 ;
        RECT 9.950 3.080 10.180 3.660 ;
        RECT 9.100 2.360 9.465 2.570 ;
        RECT 9.100 0.980 9.330 2.360 ;
        RECT 10.000 0.980 10.230 1.540 ;
        RECT 11.120 1.200 11.410 4.120 ;
        RECT 11.680 1.200 12.210 3.890 ;
        RECT 12.540 2.850 12.770 4.120 ;
        RECT 13.460 4.120 15.430 4.350 ;
        RECT 13.460 2.850 13.690 4.120 ;
        RECT 12.540 2.620 13.690 2.850 ;
        RECT 14.080 1.200 14.310 3.890 ;
        RECT 15.170 1.200 15.430 4.120 ;
        RECT 16.190 2.895 16.420 3.890 ;
        RECT 15.700 2.665 16.420 2.895 ;
        RECT 15.700 1.485 15.930 2.665 ;
        RECT 18.460 2.490 18.790 3.890 ;
        RECT 16.570 2.435 18.790 2.490 ;
        RECT 16.160 2.260 18.790 2.435 ;
        RECT 16.160 2.050 16.720 2.260 ;
        RECT 15.700 1.255 16.605 1.485 ;
        RECT 18.560 1.200 18.790 2.260 ;
        RECT 8.180 0.750 10.230 0.980 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__mux4_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__mux4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__mux4_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.120000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.190 1.210 19.450 2.030 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.120000 ;
    PORT
      LAYER Metal1 ;
        RECT 15.830 2.150 16.090 2.710 ;
    END
  END I1
  PIN I2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.120000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.700 2.330 1.080 2.710 ;
    END
  END I2
  PIN I3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.120000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.630 2.150 4.890 2.710 ;
    END
  END I3
  PIN S0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.360000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.350 2.220 2.580 2.710 ;
        RECT 2.350 1.770 3.885 2.220 ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.240000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.905 2.175 13.135 2.830 ;
        RECT 11.790 1.945 13.135 2.175 ;
        RECT 12.470 1.210 12.730 1.945 ;
    END
  END S1
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.163200 ;
    PORT
      LAYER Metal1 ;
        RECT 6.590 2.030 6.825 3.380 ;
        RECT 9.075 2.030 9.370 3.380 ;
        RECT 6.590 1.800 9.370 2.030 ;
        RECT 6.590 1.230 6.820 1.800 ;
        RECT 8.830 1.210 9.370 1.800 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 21.280 5.490 ;
        RECT 0.410 3.040 0.640 4.590 ;
        RECT 5.355 4.070 5.585 4.590 ;
        RECT 7.835 4.070 8.065 4.590 ;
        RECT 10.095 3.440 10.325 4.590 ;
        RECT 15.245 3.400 15.475 4.590 ;
        RECT 19.585 3.040 19.815 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 21.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 21.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.310 0.450 0.540 1.570 ;
        RECT 5.470 0.450 5.700 1.570 ;
        RECT 7.710 0.450 7.940 1.570 ;
        RECT 9.950 0.450 10.180 1.570 ;
        RECT 15.205 0.450 15.435 1.570 ;
        RECT 19.685 0.450 19.915 1.570 ;
        RECT 0.000 -0.450 21.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 13.465 4.080 15.015 4.310 ;
        RECT 1.430 1.230 1.660 3.850 ;
        RECT 1.890 3.840 3.020 3.850 ;
        RECT 1.890 3.610 9.865 3.840 ;
        RECT 1.890 1.515 2.120 3.610 ;
        RECT 2.790 3.040 3.020 3.610 ;
        RECT 4.115 1.925 4.345 3.380 ;
        RECT 9.635 3.210 9.865 3.610 ;
        RECT 11.425 3.270 11.655 3.850 ;
        RECT 10.945 3.210 11.655 3.270 ;
        RECT 9.635 3.040 11.655 3.210 ;
        RECT 9.635 2.980 11.100 3.040 ;
        RECT 9.655 2.030 9.885 2.710 ;
        RECT 4.115 1.695 4.580 1.925 ;
        RECT 9.655 1.800 10.640 2.030 ;
        RECT 1.890 1.285 3.515 1.515 ;
        RECT 4.350 1.230 4.580 1.695 ;
        RECT 10.410 1.000 10.640 1.800 ;
        RECT 10.870 1.230 11.100 2.980 ;
        RECT 12.445 2.635 12.675 3.850 ;
        RECT 11.330 2.405 12.675 2.635 ;
        RECT 11.330 1.000 11.560 2.405 ;
        RECT 13.465 1.570 13.695 4.080 ;
        RECT 12.005 1.000 12.235 1.570 ;
        RECT 13.125 1.230 13.695 1.570 ;
        RECT 13.925 1.230 14.455 3.850 ;
        RECT 14.785 3.170 15.015 4.080 ;
        RECT 15.705 4.080 17.675 4.310 ;
        RECT 15.705 3.170 15.935 4.080 ;
        RECT 14.785 2.940 15.935 3.170 ;
        RECT 16.325 1.230 16.555 3.850 ;
        RECT 17.445 1.230 17.675 4.080 ;
        RECT 18.565 2.950 18.795 3.850 ;
        RECT 17.945 2.720 18.795 2.950 ;
        RECT 17.945 1.515 18.175 2.720 ;
        RECT 20.705 2.490 21.035 3.850 ;
        RECT 18.405 2.260 21.035 2.490 ;
        RECT 18.405 2.150 18.635 2.260 ;
        RECT 17.945 1.285 18.850 1.515 ;
        RECT 20.805 1.230 21.035 2.260 ;
        RECT 10.410 0.770 12.235 1.000 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__mux4_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nand2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.800 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.614500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 2.330 2.090 3.270 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.614500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.635 1.770 0.975 2.710 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.436200 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 3.600 2.550 3.830 ;
        RECT 1.270 3.020 1.530 3.600 ;
        RECT 2.320 1.590 2.550 3.600 ;
        RECT 1.270 1.210 2.550 1.590 ;
        RECT 2.290 0.680 2.550 1.210 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 2.800 5.490 ;
        RECT 0.250 3.690 0.480 4.590 ;
        RECT 2.290 4.160 2.520 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 3.230 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 3.230 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 0.450 0.480 1.165 ;
        RECT 0.000 -0.450 2.800 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nand2_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nand2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.040 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.229000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.685 1.830 2.715 2.305 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.229000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.940 3.245 3.170 ;
        RECT 0.710 1.210 0.970 2.940 ;
        RECT 3.015 2.100 3.245 2.940 ;
        RECT 3.015 1.830 4.030 2.100 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.397200 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 3.630 1.495 4.210 ;
        RECT 3.305 3.630 3.535 4.210 ;
        RECT 1.265 3.580 3.535 3.630 ;
        RECT 1.265 3.400 4.490 3.580 ;
        RECT 3.390 3.350 4.490 3.400 ;
        RECT 4.070 2.330 4.490 3.350 ;
        RECT 4.260 1.590 4.490 2.330 ;
        RECT 2.285 1.210 4.490 1.590 ;
        RECT 2.285 0.680 2.515 1.210 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.040 5.490 ;
        RECT 0.245 3.860 0.475 4.590 ;
        RECT 2.285 3.860 2.515 4.590 ;
        RECT 4.325 3.860 4.555 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 5.470 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 5.470 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.165 ;
        RECT 4.325 0.450 4.555 0.695 ;
        RECT 0.000 -0.450 5.040 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nand2_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nand2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.960 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.458000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.670 2.950 6.070 3.210 ;
        RECT 2.670 2.470 3.010 2.950 ;
        RECT 5.730 2.470 6.070 2.950 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.458000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.770 1.830 8.110 2.150 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.853800 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 3.780 1.495 4.360 ;
        RECT 3.305 3.780 3.535 4.360 ;
        RECT 5.345 3.780 5.575 4.360 ;
        RECT 7.370 3.780 7.750 4.330 ;
        RECT 1.265 3.550 7.750 3.780 ;
        RECT 7.385 3.460 7.750 3.550 ;
        RECT 7.385 3.230 8.570 3.460 ;
        RECT 8.340 1.105 8.570 3.230 ;
        RECT 7.940 1.100 8.570 1.105 ;
        RECT 2.275 0.875 8.570 1.100 ;
        RECT 2.275 0.870 8.145 0.875 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 8.960 5.490 ;
        RECT 0.245 3.690 0.475 4.590 ;
        RECT 2.285 4.160 2.515 4.590 ;
        RECT 4.325 4.160 4.555 4.590 ;
        RECT 6.365 4.160 6.595 4.590 ;
        RECT 8.405 3.690 8.635 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 9.390 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.390 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.325 0.450 0.555 1.165 ;
        RECT 4.235 0.450 4.575 0.640 ;
        RECT 8.350 0.450 8.690 0.640 ;
        RECT 0.000 -0.450 8.960 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nand2_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nand3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.920 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 1.210 3.210 2.150 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.090 2.710 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.330 1.105 3.270 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.982400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 3.830 1.630 4.360 ;
        RECT 1.400 3.550 3.670 3.830 ;
        RECT 2.950 2.890 3.670 3.550 ;
        RECT 3.440 0.845 3.670 2.890 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 3.920 5.490 ;
        RECT 0.380 3.590 0.610 4.590 ;
        RECT 2.420 4.060 2.650 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 4.350 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.350 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.380 0.450 0.610 1.165 ;
        RECT 0.000 -0.450 3.920 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nand3_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nand3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.865 1.210 3.210 2.150 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.790 2.380 4.995 2.610 ;
        RECT 4.630 1.210 4.995 2.380 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.300 2.840 6.015 3.070 ;
        RECT 1.300 2.150 1.530 2.840 ;
        RECT 0.770 1.920 1.530 2.150 ;
        RECT 5.740 2.070 6.015 2.840 ;
        RECT 1.270 1.915 1.530 1.920 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.964000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 3.530 1.495 4.110 ;
        RECT 3.305 3.530 3.535 4.110 ;
        RECT 5.345 3.530 5.575 4.110 ;
        RECT 0.150 3.300 5.575 3.530 ;
        RECT 0.150 1.095 0.410 3.300 ;
        RECT 0.150 0.980 1.070 1.095 ;
        RECT 0.150 0.865 3.590 0.980 ;
        RECT 0.870 0.750 3.590 0.865 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.280 5.490 ;
        RECT 0.245 4.230 0.475 4.590 ;
        RECT 2.285 3.760 2.515 4.590 ;
        RECT 4.325 3.760 4.555 4.590 ;
        RECT 6.365 3.760 6.595 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 7.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.330 0.450 0.670 0.635 ;
        RECT 6.365 0.450 6.595 1.160 ;
        RECT 0.000 -0.450 7.280 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nand3_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nand3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.000 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.088000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.300 2.270 11.230 2.500 ;
        RECT 9.300 1.770 9.930 2.270 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.088000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.750 2.730 8.355 2.960 ;
        RECT 0.750 2.215 0.980 2.730 ;
        RECT 3.510 2.270 4.130 2.730 ;
        RECT 8.125 2.215 8.355 2.730 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.088000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.210 2.040 1.990 2.500 ;
        RECT 4.410 2.270 6.270 2.500 ;
        RECT 4.410 2.040 4.640 2.270 ;
        RECT 1.210 1.810 4.640 2.040 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.220000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 3.420 1.495 4.360 ;
        RECT 3.405 3.420 3.635 4.360 ;
        RECT 5.545 3.420 5.775 4.360 ;
        RECT 7.685 3.420 7.915 4.360 ;
        RECT 9.725 3.420 9.955 4.360 ;
        RECT 11.965 3.420 12.195 4.360 ;
        RECT 1.265 3.190 12.195 3.420 ;
        RECT 11.965 1.530 12.195 3.190 ;
        RECT 11.965 1.515 12.790 1.530 ;
        RECT 9.825 1.285 12.790 1.515 ;
        RECT 9.825 1.140 10.055 1.285 ;
        RECT 12.010 1.140 12.790 1.285 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 14.000 5.490 ;
        RECT 0.245 3.650 0.475 4.590 ;
        RECT 2.285 3.875 2.515 4.590 ;
        RECT 4.425 3.650 4.655 4.590 ;
        RECT 6.565 3.650 6.795 4.590 ;
        RECT 8.705 3.650 8.935 4.590 ;
        RECT 10.845 3.650 11.075 4.590 ;
        RECT 13.085 3.650 13.315 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 14.430 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.430 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.385 0.450 2.615 1.110 ;
        RECT 6.665 0.450 6.895 1.110 ;
        RECT 0.000 -0.450 14.000 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 1.350 3.075 1.580 ;
        RECT 0.245 0.770 0.475 1.350 ;
        RECT 2.845 1.000 3.075 1.350 ;
        RECT 4.525 1.350 9.170 1.580 ;
        RECT 4.525 1.000 4.755 1.350 ;
        RECT 2.845 0.770 4.755 1.000 ;
        RECT 8.940 0.910 9.170 1.350 ;
        RECT 10.890 0.910 11.230 1.055 ;
        RECT 13.185 0.910 13.415 1.580 ;
        RECT 8.940 0.680 13.415 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__nand3_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nand4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.040 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.985 2.270 4.330 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.915 2.215 3.210 2.710 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.090 2.555 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 1.125 2.500 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.912000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.420 3.490 1.650 4.360 ;
        RECT 3.460 3.490 3.770 4.360 ;
        RECT 1.420 3.260 3.770 3.490 ;
        RECT 3.540 3.255 3.770 3.260 ;
        RECT 3.540 3.025 4.790 3.255 ;
        RECT 4.560 1.490 4.790 3.025 ;
        RECT 4.480 0.680 4.790 1.490 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.040 5.490 ;
        RECT 0.400 3.720 0.630 4.590 ;
        RECT 2.440 3.720 2.670 4.590 ;
        RECT 4.480 3.485 4.710 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 5.470 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 5.470 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 0.450 0.630 1.490 ;
        RECT 0.000 -0.450 5.040 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nand4_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nand4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.960 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 2.215 3.875 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.865 2.940 4.465 3.170 ;
        RECT 2.865 2.215 3.095 2.940 ;
        RECT 4.235 2.710 4.465 2.940 ;
        RECT 4.235 2.215 6.015 2.710 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.985 2.090 2.555 ;
        RECT 6.805 1.985 7.035 2.555 ;
        RECT 1.830 1.755 7.035 1.985 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.050 3.540 4.925 3.630 ;
        RECT 1.300 3.400 4.925 3.540 ;
        RECT 1.300 3.310 2.235 3.400 ;
        RECT 1.300 2.555 1.530 3.310 ;
        RECT 4.695 3.170 4.925 3.400 ;
        RECT 4.695 2.940 8.055 3.170 ;
        RECT 0.825 2.215 1.530 2.555 ;
        RECT 7.825 2.215 8.055 2.940 ;
        RECT 1.270 1.770 1.530 2.215 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.809600 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 4.000 0.475 4.360 ;
        RECT 1.680 4.045 5.205 4.090 ;
        RECT 1.680 4.000 6.595 4.045 ;
        RECT 0.150 3.860 6.595 4.000 ;
        RECT 0.150 3.770 1.865 3.860 ;
        RECT 5.065 3.815 6.595 3.860 ;
        RECT 0.150 1.985 0.475 3.770 ;
        RECT 6.365 3.630 6.595 3.815 ;
        RECT 8.405 3.630 8.635 4.360 ;
        RECT 6.365 3.400 8.635 3.630 ;
        RECT 0.150 1.755 1.040 1.985 ;
        RECT 0.810 0.910 1.040 1.755 ;
        RECT 4.325 0.910 4.555 1.490 ;
        RECT 0.810 0.680 4.555 0.910 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 8.960 5.490 ;
        RECT 1.265 4.230 1.495 4.590 ;
        RECT 3.305 4.320 3.535 4.590 ;
        RECT 5.345 4.275 5.575 4.590 ;
        RECT 7.385 3.860 7.615 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 9.390 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.390 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 8.405 0.450 8.635 1.490 ;
        RECT 0.000 -0.450 8.960 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nand4_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nand4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand4_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.360 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.728000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.670 1.985 10.150 2.500 ;
        RECT 12.365 2.270 14.230 2.500 ;
        RECT 12.365 1.985 12.595 2.270 ;
        RECT 9.670 1.755 12.595 1.985 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.728000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.930 2.730 15.935 2.960 ;
        RECT 8.930 2.270 9.270 2.730 ;
        RECT 11.350 2.215 12.135 2.730 ;
        RECT 15.705 2.215 15.935 2.730 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.728000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.730 6.530 2.960 ;
        RECT 0.710 2.270 1.050 2.730 ;
        RECT 3.745 2.215 3.975 2.730 ;
        RECT 6.300 2.500 6.530 2.730 ;
        RECT 6.300 2.270 8.110 2.500 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.728000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.985 2.170 2.500 ;
        RECT 4.205 2.270 6.070 2.500 ;
        RECT 4.205 1.985 4.435 2.270 ;
        RECT 1.830 1.755 4.435 1.985 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.697600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 3.420 1.495 4.360 ;
        RECT 2.890 3.420 3.535 4.360 ;
        RECT 5.345 3.420 5.575 4.360 ;
        RECT 7.385 3.420 7.615 4.360 ;
        RECT 9.425 3.420 9.655 4.360 ;
        RECT 11.465 3.420 11.695 4.360 ;
        RECT 13.505 3.420 13.735 4.360 ;
        RECT 15.545 3.420 15.775 4.360 ;
        RECT 1.265 3.190 16.395 3.420 ;
        RECT 16.165 1.425 16.395 3.190 ;
        RECT 10.390 1.195 16.395 1.425 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.360 5.490 ;
        RECT 0.245 3.650 0.475 4.590 ;
        RECT 2.285 3.650 2.515 4.590 ;
        RECT 4.325 3.650 4.555 4.590 ;
        RECT 6.365 3.650 6.595 4.590 ;
        RECT 8.405 3.650 8.635 4.590 ;
        RECT 10.445 3.650 10.675 4.590 ;
        RECT 12.485 3.650 12.715 4.590 ;
        RECT 14.525 3.650 14.755 4.590 ;
        RECT 16.565 3.650 16.795 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 17.790 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 17.790 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.285 0.450 2.515 1.020 ;
        RECT 6.365 0.450 6.595 1.020 ;
        RECT 0.000 -0.450 17.360 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 1.260 10.160 1.490 ;
        RECT 0.245 0.680 0.475 1.260 ;
        RECT 4.325 0.680 4.555 1.260 ;
        RECT 9.930 0.965 10.160 1.260 ;
        RECT 9.930 0.735 16.850 0.965 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__nand4_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nor2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.467000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.090 2.555 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.467000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.680 2.270 1.020 2.710 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.283600 ;
    PORT
      LAYER Metal1 ;
        RECT 2.435 3.015 2.665 4.360 ;
        RECT 1.270 2.785 2.665 3.015 ;
        RECT 1.270 0.680 1.595 2.785 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 3.360 5.490 ;
        RECT 0.295 3.550 0.525 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 3.790 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 3.790 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.400 ;
        RECT 2.485 0.450 2.715 1.400 ;
        RECT 0.000 -0.450 3.360 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nor2_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nor2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.934000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.800 2.270 2.140 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.934000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.875 2.940 3.950 3.170 ;
        RECT 0.875 2.215 1.105 2.940 ;
        RECT 3.510 2.270 3.950 2.940 ;
        RECT 3.510 1.770 3.770 2.270 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.999900 ;
    PORT
      LAYER Metal1 ;
        RECT 2.485 3.780 2.715 4.360 ;
        RECT 2.485 3.550 4.410 3.780 ;
        RECT 4.180 1.720 4.410 3.550 ;
        RECT 4.070 1.490 4.410 1.720 ;
        RECT 1.365 1.210 4.410 1.490 ;
        RECT 1.365 1.160 3.835 1.210 ;
        RECT 1.365 0.680 1.595 1.160 ;
        RECT 3.605 0.680 3.835 1.160 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.600 5.490 ;
        RECT 0.295 3.550 0.525 4.590 ;
        RECT 4.675 3.550 4.905 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.400 ;
        RECT 2.485 0.450 2.715 0.930 ;
        RECT 4.725 0.450 4.955 1.400 ;
        RECT 0.000 -0.450 5.600 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nor2_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nor2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.868000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.060 2.270 3.810 2.500 ;
        RECT 3.580 2.000 3.810 2.270 ;
        RECT 4.630 2.270 6.620 2.500 ;
        RECT 4.630 2.000 4.890 2.270 ;
        RECT 3.580 1.770 4.890 2.000 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.868000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.600 2.730 7.080 2.960 ;
        RECT 2.600 2.500 2.830 2.730 ;
        RECT 1.200 2.270 2.830 2.500 ;
        RECT 4.040 2.270 4.380 2.730 ;
        RECT 6.850 2.500 7.080 2.730 ;
        RECT 6.850 2.270 8.860 2.500 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.091300 ;
    PORT
      LAYER Metal1 ;
        RECT 2.485 3.420 2.715 4.360 ;
        RECT 6.915 3.420 7.145 4.360 ;
        RECT 0.710 3.190 7.145 3.420 ;
        RECT 0.710 1.490 0.970 3.190 ;
        RECT 0.710 1.260 8.315 1.490 ;
        RECT 1.365 0.680 1.595 1.260 ;
        RECT 3.605 0.680 3.835 1.260 ;
        RECT 5.845 0.680 6.075 1.260 ;
        RECT 8.085 0.680 8.315 1.260 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 10.080 5.490 ;
        RECT 0.295 3.650 0.525 4.590 ;
        RECT 4.675 3.650 4.905 4.590 ;
        RECT 9.155 3.650 9.385 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 10.510 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 10.510 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.020 ;
        RECT 4.725 0.450 4.955 1.020 ;
        RECT 6.965 0.450 7.195 1.020 ;
        RECT 9.205 0.450 9.435 1.400 ;
        RECT 0.000 -0.450 10.080 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nor2_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nor3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 1.770 3.210 2.555 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.800 2.270 2.140 2.710 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.215 1.015 2.710 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.563600 ;
    PORT
      LAYER Metal1 ;
        RECT 3.505 1.480 3.835 4.360 ;
        RECT 1.365 1.250 3.835 1.480 ;
        RECT 1.365 0.680 1.595 1.250 ;
        RECT 3.605 0.680 3.835 1.250 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 4.480 5.490 ;
        RECT 0.345 3.550 0.575 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 4.910 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.020 ;
        RECT 2.485 0.450 2.715 1.020 ;
        RECT 0.000 -0.450 4.480 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nor3_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nor3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.475 2.215 3.770 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 2.940 5.445 3.170 ;
        RECT 1.830 2.215 2.135 2.940 ;
        RECT 5.215 2.215 5.445 2.940 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 3.400 6.570 3.630 ;
        RECT 1.265 2.215 1.495 3.400 ;
        RECT 6.310 2.215 6.570 3.400 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.651400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.805 3.930 3.840 4.160 ;
        RECT 0.805 1.590 1.035 3.930 ;
        RECT 0.245 1.480 1.035 1.590 ;
        RECT 0.245 1.250 7.195 1.480 ;
        RECT 0.245 1.210 2.715 1.250 ;
        RECT 0.245 0.680 0.475 1.210 ;
        RECT 2.485 0.680 2.715 1.210 ;
        RECT 4.725 0.680 4.955 1.250 ;
        RECT 6.965 0.680 7.195 1.250 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.840 5.490 ;
        RECT 0.345 3.875 0.575 4.590 ;
        RECT 6.865 3.875 7.095 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 8.270 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.270 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 0.980 ;
        RECT 3.605 0.450 3.835 1.020 ;
        RECT 5.845 0.450 6.075 1.020 ;
        RECT 0.000 -0.450 7.840 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nor3_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nor3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.560 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.556000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.800 1.710 11.730 2.150 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.556000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.825 2.895 6.975 3.125 ;
        RECT 0.825 2.325 1.055 2.895 ;
        RECT 3.510 2.380 4.330 2.895 ;
        RECT 6.745 2.610 6.975 2.895 ;
        RECT 6.745 2.380 8.810 2.610 ;
        RECT 3.510 2.330 3.770 2.380 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.556000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.940 2.000 3.280 2.610 ;
        RECT 6.285 2.150 6.515 2.665 ;
        RECT 4.070 2.000 6.515 2.150 ;
        RECT 2.940 1.770 6.515 2.000 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.734000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.325 2.880 10.555 3.900 ;
        RECT 11.910 3.090 12.695 3.900 ;
        RECT 11.910 2.880 12.190 3.090 ;
        RECT 10.325 2.650 12.190 2.880 ;
        RECT 11.960 1.480 12.190 2.650 ;
        RECT 1.365 1.250 12.795 1.480 ;
        RECT 1.365 0.680 1.595 1.250 ;
        RECT 3.605 0.680 3.835 1.250 ;
        RECT 5.845 0.680 6.075 1.250 ;
        RECT 8.085 0.680 8.315 1.250 ;
        RECT 10.325 0.680 10.555 1.250 ;
        RECT 12.565 0.680 12.795 1.250 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 14.560 5.490 ;
        RECT 2.385 3.825 2.615 4.590 ;
        RECT 6.865 3.815 7.095 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 14.990 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.990 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.020 ;
        RECT 2.485 0.450 2.715 1.020 ;
        RECT 4.725 0.450 4.955 1.020 ;
        RECT 6.965 0.450 7.195 1.020 ;
        RECT 9.205 0.450 9.435 1.020 ;
        RECT 11.445 0.450 11.675 1.020 ;
        RECT 13.685 0.450 13.915 1.020 ;
        RECT 0.000 -0.450 14.560 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.585 0.475 3.920 ;
        RECT 4.625 3.585 4.855 4.165 ;
        RECT 7.375 4.130 13.815 4.360 ;
        RECT 7.375 3.585 7.605 4.130 ;
        RECT 0.245 3.355 7.605 3.585 ;
        RECT 0.245 3.110 0.475 3.355 ;
        RECT 11.345 3.110 11.575 4.130 ;
        RECT 13.585 3.110 13.815 4.130 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__nor3_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nor4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.311000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.070 1.770 4.330 2.555 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.311000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.920 2.270 3.260 2.710 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.311000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.800 2.270 2.140 2.710 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.311000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.215 1.015 2.710 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.491600 ;
    PORT
      LAYER Metal1 ;
        RECT 4.625 3.015 4.855 4.360 ;
        RECT 3.510 2.785 4.855 3.015 ;
        RECT 3.510 1.440 3.835 2.785 ;
        RECT 1.365 1.210 3.835 1.440 ;
        RECT 1.365 0.680 1.595 1.210 ;
        RECT 3.605 0.680 3.835 1.210 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.600 5.490 ;
        RECT 0.345 3.550 0.575 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.005 ;
        RECT 2.485 0.450 2.715 0.980 ;
        RECT 4.725 0.450 4.955 1.005 ;
        RECT 0.000 -0.450 5.600 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nor4_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nor4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.622000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.870 2.150 7.130 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.622000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.340 2.940 9.120 3.170 ;
        RECT 6.340 2.555 6.570 2.940 ;
        RECT 5.770 1.770 6.570 2.555 ;
        RECT 8.890 2.215 9.120 2.940 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.622000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.930 2.785 4.510 3.015 ;
        RECT 0.930 2.215 1.160 2.785 ;
        RECT 4.070 1.770 4.510 2.785 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.622000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.090 2.555 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.718200 ;
    PORT
      LAYER Metal1 ;
        RECT 7.280 3.630 7.510 3.890 ;
        RECT 5.190 3.400 7.510 3.630 ;
        RECT 5.190 1.455 5.450 3.400 ;
        RECT 1.370 1.225 8.680 1.455 ;
        RECT 1.370 0.680 1.600 1.225 ;
        RECT 3.610 1.210 6.440 1.225 ;
        RECT 3.610 0.680 3.840 1.210 ;
        RECT 6.210 0.680 6.440 1.210 ;
        RECT 8.450 0.680 8.680 1.225 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 10.080 5.490 ;
        RECT 2.440 3.705 2.670 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 10.510 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 10.510 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 0.450 0.480 1.020 ;
        RECT 2.490 0.450 2.720 0.995 ;
        RECT 4.910 0.450 5.140 0.980 ;
        RECT 7.330 0.450 7.560 0.995 ;
        RECT 9.570 0.450 9.800 0.995 ;
        RECT 0.000 -0.450 10.080 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.350 4.130 2.210 4.360 ;
        RECT 0.350 3.550 0.580 4.130 ;
        RECT 1.980 3.475 2.210 4.130 ;
        RECT 2.900 4.130 9.700 4.360 ;
        RECT 2.900 3.475 3.130 4.130 ;
        RECT 9.470 3.550 9.700 4.130 ;
        RECT 1.980 3.245 3.130 3.475 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__nor4_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nor4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor4_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.244000 ;
    PORT
      LAYER Metal1 ;
        RECT 13.465 2.215 17.460 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.244000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.870 1.985 11.100 2.555 ;
        RECT 19.550 1.985 20.010 2.555 ;
        RECT 10.870 1.755 20.010 1.985 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.244000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.100 2.785 7.700 3.015 ;
        RECT 1.100 2.150 1.330 2.785 ;
        RECT 4.590 2.215 4.820 2.785 ;
        RECT 7.470 2.500 7.700 2.785 ;
        RECT 7.470 2.270 9.715 2.500 ;
        RECT 0.710 1.770 1.330 2.150 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.244000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.480 1.985 3.710 2.555 ;
        RECT 6.780 1.985 7.240 2.555 ;
        RECT 3.480 1.755 7.240 1.985 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.389400 ;
    PORT
      LAYER Metal1 ;
        RECT 12.890 3.320 13.120 3.900 ;
        RECT 17.810 3.320 18.040 3.900 ;
        RECT 12.890 3.090 20.635 3.320 ;
        RECT 20.405 1.590 20.635 3.090 ;
        RECT 20.175 1.455 20.635 1.590 ;
        RECT 1.680 1.225 5.910 1.455 ;
        RECT 1.680 0.680 1.910 1.225 ;
        RECT 3.920 0.680 4.150 1.225 ;
        RECT 5.680 0.910 5.910 1.225 ;
        RECT 6.520 1.225 20.635 1.455 ;
        RECT 6.520 0.910 6.750 1.225 ;
        RECT 5.680 0.680 6.750 0.910 ;
        RECT 8.760 0.680 8.990 1.225 ;
        RECT 11.360 0.680 11.590 1.225 ;
        RECT 13.960 0.680 14.190 1.225 ;
        RECT 16.560 0.680 16.790 1.225 ;
        RECT 19.160 1.210 20.635 1.225 ;
        RECT 19.160 0.680 19.390 1.210 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 21.280 5.490 ;
        RECT 2.750 3.705 2.980 4.590 ;
        RECT 7.590 3.705 7.820 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 21.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 21.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.560 0.450 0.790 0.995 ;
        RECT 2.800 0.450 3.030 0.995 ;
        RECT 5.220 0.450 5.450 0.995 ;
        RECT 7.640 0.450 7.870 0.995 ;
        RECT 10.060 0.450 10.290 0.995 ;
        RECT 12.660 0.450 12.890 0.995 ;
        RECT 15.260 0.450 15.490 0.970 ;
        RECT 17.860 0.450 18.090 0.995 ;
        RECT 20.460 0.450 20.690 0.980 ;
        RECT 0.000 -0.450 21.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.660 4.130 2.520 4.360 ;
        RECT 0.660 3.550 0.890 4.130 ;
        RECT 2.290 3.475 2.520 4.130 ;
        RECT 5.170 3.475 5.400 4.360 ;
        RECT 8.050 4.130 20.590 4.360 ;
        RECT 8.050 3.475 8.280 4.130 ;
        RECT 15.210 3.550 15.440 4.130 ;
        RECT 20.360 3.550 20.590 4.130 ;
        RECT 2.290 3.245 8.280 3.475 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__nor4_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai21_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai21_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.090 2.555 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.680 2.270 1.020 2.710 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.614500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 2.270 3.290 2.710 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.911900 ;
    PORT
      LAYER Metal1 ;
        RECT 2.385 3.015 2.615 4.360 ;
        RECT 1.270 2.785 2.615 3.015 ;
        RECT 1.270 1.140 1.595 2.785 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 4.480 5.490 ;
        RECT 0.295 3.550 0.525 4.590 ;
        RECT 3.585 3.550 3.815 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 4.910 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 3.605 0.450 3.835 1.655 ;
        RECT 0.000 -0.450 4.480 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 0.910 0.475 1.655 ;
        RECT 2.485 0.910 2.715 1.655 ;
        RECT 0.245 0.680 2.715 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai21_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai21_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai21_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.035 2.215 4.330 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 2.940 6.515 3.170 ;
        RECT 2.950 2.270 3.310 2.940 ;
        RECT 6.285 2.215 6.515 2.940 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.229000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 2.270 1.070 2.650 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.362800 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.630 1.595 4.320 ;
        RECT 4.675 3.630 4.905 4.360 ;
        RECT 1.365 3.400 6.975 3.630 ;
        RECT 6.745 1.950 6.975 3.400 ;
        RECT 3.605 1.720 6.975 1.950 ;
        RECT 3.605 1.140 3.835 1.720 ;
        RECT 5.190 1.140 6.075 1.720 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.840 5.490 ;
        RECT 0.345 3.665 0.575 4.590 ;
        RECT 2.385 3.860 2.615 4.590 ;
        RECT 6.865 3.860 7.095 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 8.270 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.270 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.490 ;
        RECT 0.000 -0.450 7.840 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 1.720 2.715 1.950 ;
        RECT 0.245 0.680 0.475 1.720 ;
        RECT 2.485 0.910 2.715 1.720 ;
        RECT 4.725 0.910 4.955 1.490 ;
        RECT 6.965 0.910 7.195 1.490 ;
        RECT 2.485 0.680 7.195 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai21_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai21_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai21_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.560 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.060 2.270 3.770 2.500 ;
        RECT 3.510 2.040 3.770 2.270 ;
        RECT 4.610 2.270 6.570 2.500 ;
        RECT 4.610 2.040 4.840 2.270 ;
        RECT 3.510 1.810 4.840 2.040 ;
        RECT 3.510 1.770 3.770 1.810 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.600 2.730 7.030 2.960 ;
        RECT 2.600 2.500 2.830 2.730 ;
        RECT 1.250 2.270 2.830 2.500 ;
        RECT 4.040 2.270 4.380 2.730 ;
        RECT 6.800 2.500 7.030 2.730 ;
        RECT 6.800 2.270 8.810 2.500 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.458000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.270 2.270 12.850 2.500 ;
        RECT 11.350 1.770 11.610 2.270 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.798600 ;
    PORT
      LAYER Metal1 ;
        RECT 2.485 3.420 2.715 4.360 ;
        RECT 6.915 3.420 7.145 4.360 ;
        RECT 10.325 3.420 10.555 4.360 ;
        RECT 12.515 3.420 12.745 4.360 ;
        RECT 0.790 3.190 12.745 3.420 ;
        RECT 0.790 2.040 1.020 3.190 ;
        RECT 0.790 1.810 3.210 2.040 ;
        RECT 1.365 1.140 1.595 1.810 ;
        RECT 2.950 1.480 3.210 1.810 ;
        RECT 3.935 1.480 8.315 1.570 ;
        RECT 2.950 1.340 8.315 1.480 ;
        RECT 2.950 1.140 4.120 1.340 ;
        RECT 5.845 1.140 6.075 1.340 ;
        RECT 8.085 1.140 8.315 1.340 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 14.560 5.490 ;
        RECT 0.345 3.650 0.575 4.590 ;
        RECT 4.675 3.650 4.905 4.590 ;
        RECT 9.105 3.650 9.335 4.590 ;
        RECT 11.345 3.650 11.575 4.590 ;
        RECT 13.635 3.650 13.865 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 14.990 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.990 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 10.325 0.450 10.555 1.195 ;
        RECT 12.565 0.450 12.795 1.110 ;
        RECT 0.000 -0.450 14.560 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 0.910 0.475 1.580 ;
        RECT 2.485 0.910 2.715 1.580 ;
        RECT 9.205 1.540 11.150 1.655 ;
        RECT 11.775 1.540 13.915 1.580 ;
        RECT 9.205 1.425 13.915 1.540 ;
        RECT 4.725 0.910 4.955 1.110 ;
        RECT 6.965 0.910 7.195 1.110 ;
        RECT 9.205 0.910 9.435 1.425 ;
        RECT 10.950 1.350 13.915 1.425 ;
        RECT 10.950 1.310 11.905 1.350 ;
        RECT 0.245 0.680 9.435 0.910 ;
        RECT 11.445 0.730 11.905 1.310 ;
        RECT 13.685 0.770 13.915 1.350 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai21_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai22_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai22_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 1.770 3.210 2.555 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.070 1.770 4.330 2.555 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.800 2.270 2.140 2.710 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.215 1.015 3.270 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.821000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.535 3.015 2.765 4.360 ;
        RECT 2.535 2.785 3.835 3.015 ;
        RECT 3.510 1.140 3.835 2.785 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.600 5.490 ;
        RECT 0.345 3.550 0.575 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.525 ;
        RECT 0.000 -0.450 5.600 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 1.755 2.715 1.985 ;
        RECT 0.245 0.715 0.475 1.755 ;
        RECT 2.485 0.910 2.715 1.755 ;
        RECT 4.725 0.910 4.955 1.525 ;
        RECT 2.485 0.680 4.955 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai22_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai22_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai22_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.280 2.270 6.620 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.350 2.940 8.755 3.170 ;
        RECT 5.350 2.270 5.690 2.940 ;
        RECT 6.870 2.215 8.755 2.940 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.750 2.270 2.090 2.710 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.870 2.940 4.330 3.170 ;
        RECT 0.870 2.270 1.210 2.940 ;
        RECT 2.390 2.270 4.330 2.940 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.733500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.535 3.630 2.765 4.360 ;
        RECT 6.915 3.630 7.145 4.360 ;
        RECT 2.535 3.400 9.215 3.630 ;
        RECT 8.985 1.985 9.215 3.400 ;
        RECT 5.845 1.755 9.215 1.985 ;
        RECT 5.845 1.140 6.075 1.755 ;
        RECT 7.990 1.140 8.315 1.755 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 10.080 5.490 ;
        RECT 0.345 3.860 0.575 4.590 ;
        RECT 4.625 3.860 4.855 4.590 ;
        RECT 9.105 3.860 9.335 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 10.510 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 10.510 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.525 ;
        RECT 3.605 0.450 3.835 1.055 ;
        RECT 0.000 -0.450 10.080 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 1.755 4.955 1.985 ;
        RECT 0.245 0.715 0.475 1.755 ;
        RECT 2.485 1.285 4.955 1.755 ;
        RECT 4.725 0.910 4.955 1.285 ;
        RECT 6.965 0.910 7.195 1.525 ;
        RECT 9.205 0.910 9.435 1.525 ;
        RECT 4.725 0.680 9.435 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai22_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai22_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai22_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.040 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.730 1.985 11.340 2.500 ;
        RECT 13.515 2.270 15.530 2.500 ;
        RECT 13.515 1.985 13.745 2.270 ;
        RECT 10.730 1.755 13.745 1.985 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.885 2.730 17.715 2.960 ;
        RECT 9.885 2.215 10.115 2.730 ;
        RECT 12.470 2.215 13.285 2.730 ;
        RECT 17.485 2.215 17.715 2.730 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.110 2.040 3.450 2.500 ;
        RECT 4.810 2.270 6.570 2.500 ;
        RECT 4.810 2.150 5.040 2.270 ;
        RECT 4.580 2.040 5.040 2.150 ;
        RECT 3.110 1.770 5.040 2.040 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.875 2.730 7.030 2.960 ;
        RECT 0.875 2.215 1.105 2.730 ;
        RECT 4.040 2.270 4.380 2.730 ;
        RECT 6.800 2.500 7.030 2.730 ;
        RECT 6.800 2.270 8.810 2.500 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 7.558500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.585 3.420 2.815 4.360 ;
        RECT 6.865 3.420 7.095 4.360 ;
        RECT 11.395 3.420 11.625 4.360 ;
        RECT 15.975 3.830 16.205 4.360 ;
        RECT 15.975 3.450 18.330 3.830 ;
        RECT 15.975 3.420 18.175 3.450 ;
        RECT 2.585 3.190 18.175 3.420 ;
        RECT 17.945 1.475 18.175 3.190 ;
        RECT 10.270 1.245 18.175 1.475 ;
        RECT 10.270 1.140 10.610 1.245 ;
        RECT 12.510 1.140 15.090 1.245 ;
        RECT 16.990 1.140 18.175 1.245 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 19.040 5.490 ;
        RECT 0.295 3.550 0.525 4.590 ;
        RECT 4.675 3.650 4.905 4.590 ;
        RECT 9.105 3.650 9.335 4.590 ;
        RECT 13.635 3.650 13.865 4.590 ;
        RECT 18.065 4.060 18.295 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 19.470 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 19.470 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.070 ;
        RECT 3.605 0.450 3.835 1.070 ;
        RECT 5.845 0.450 6.075 1.070 ;
        RECT 8.085 0.450 8.315 1.070 ;
        RECT 0.000 -0.450 19.040 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 1.310 9.435 1.540 ;
        RECT 0.245 0.730 0.475 1.310 ;
        RECT 2.485 0.730 2.715 1.310 ;
        RECT 4.725 0.730 4.955 1.310 ;
        RECT 6.965 0.730 7.195 1.310 ;
        RECT 9.205 0.910 9.435 1.310 ;
        RECT 11.390 0.910 11.730 1.015 ;
        RECT 15.870 0.910 16.210 1.015 ;
        RECT 18.405 0.910 18.635 1.540 ;
        RECT 9.205 0.680 18.635 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai22_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai31_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai31_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.135 2.555 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.920 1.770 3.260 2.500 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.990 1.770 4.330 2.500 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.614500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 1.770 0.970 2.500 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.525600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.465 3.830 1.695 4.360 ;
        RECT 1.465 3.450 2.650 3.830 ;
        RECT 2.420 1.540 2.650 3.450 ;
        RECT 2.420 1.310 4.955 1.540 ;
        RECT 2.420 1.140 2.770 1.310 ;
        RECT 4.725 0.730 4.955 1.310 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.600 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.540 ;
        RECT 0.000 -0.450 5.600 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 0.910 1.595 1.540 ;
        RECT 3.605 0.910 3.835 1.070 ;
        RECT 1.365 0.680 3.835 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai31_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai31_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai31_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.630 2.270 5.500 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.040 2.150 4.380 2.500 ;
        RECT 3.510 2.040 4.380 2.150 ;
        RECT 6.045 2.215 7.685 2.555 ;
        RECT 6.045 2.040 6.275 2.215 ;
        RECT 3.510 1.810 6.275 2.040 ;
        RECT 3.510 1.770 3.770 1.810 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.055 2.940 8.220 3.170 ;
        RECT 3.055 2.215 3.285 2.940 ;
        RECT 7.990 2.710 8.220 2.940 ;
        RECT 7.990 2.215 8.755 2.710 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.229000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.675 2.215 0.970 2.710 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.131450 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.630 1.595 4.360 ;
        RECT 5.795 3.630 6.025 4.360 ;
        RECT 1.365 3.400 9.215 3.630 ;
        RECT 8.985 1.935 9.215 3.400 ;
        RECT 6.505 1.705 9.215 1.935 ;
        RECT 6.505 1.580 6.735 1.705 ;
        RECT 3.935 1.540 6.735 1.580 ;
        RECT 3.605 1.350 6.735 1.540 ;
        RECT 3.605 1.140 4.065 1.350 ;
        RECT 5.845 1.140 6.735 1.350 ;
        RECT 7.430 1.140 8.315 1.705 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 10.080 5.490 ;
        RECT 0.295 3.860 0.525 4.590 ;
        RECT 2.385 3.860 2.615 4.590 ;
        RECT 9.105 3.860 9.335 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 10.510 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 10.510 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.525 ;
        RECT 0.000 -0.450 10.080 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 1.755 2.715 1.985 ;
        RECT 0.245 0.845 0.475 1.755 ;
        RECT 2.485 0.910 2.715 1.755 ;
        RECT 4.725 0.910 4.955 1.120 ;
        RECT 6.965 0.910 7.195 1.185 ;
        RECT 9.440 0.910 9.670 1.655 ;
        RECT 2.485 0.680 9.670 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai31_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai31_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai31_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.590 2.270 8.250 2.500 ;
        RECT 7.990 2.000 8.250 2.270 ;
        RECT 10.160 2.270 11.100 2.500 ;
        RECT 10.160 2.000 10.390 2.270 ;
        RECT 7.990 1.770 10.390 2.000 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.355 2.730 13.235 2.960 ;
        RECT 5.355 2.215 5.585 2.730 ;
        RECT 9.590 2.270 9.930 2.730 ;
        RECT 13.005 2.215 13.235 2.730 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 2.270 3.890 2.500 ;
        RECT 1.270 1.770 1.530 2.270 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.458000 ;
    PORT
      LAYER Metal1 ;
        RECT 15.270 2.270 17.850 2.710 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 8.509650 ;
    PORT
      LAYER Metal1 ;
        RECT 6.960 3.605 11.625 3.890 ;
        RECT 11.395 3.420 11.625 3.605 ;
        RECT 15.325 3.420 15.555 4.360 ;
        RECT 11.395 3.320 15.555 3.420 ;
        RECT 17.515 3.320 17.745 4.360 ;
        RECT 11.395 3.190 17.745 3.320 ;
        RECT 13.465 3.090 17.745 3.190 ;
        RECT 13.465 1.985 13.695 3.090 ;
        RECT 10.620 1.755 13.695 1.985 ;
        RECT 1.695 1.540 7.825 1.605 ;
        RECT 10.620 1.540 10.850 1.755 ;
        RECT 1.365 1.375 10.850 1.540 ;
        RECT 1.365 1.140 1.860 1.375 ;
        RECT 3.550 1.140 3.890 1.375 ;
        RECT 5.190 1.140 6.130 1.375 ;
        RECT 7.660 1.310 10.850 1.375 ;
        RECT 7.660 1.140 8.370 1.310 ;
        RECT 10.270 1.140 10.850 1.310 ;
        RECT 12.565 1.140 12.795 1.755 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 19.600 5.490 ;
        RECT 1.365 3.550 1.595 4.590 ;
        RECT 3.555 3.550 3.785 4.590 ;
        RECT 14.305 3.875 14.535 4.590 ;
        RECT 16.495 3.550 16.725 4.590 ;
        RECT 18.635 3.550 18.865 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 20.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 20.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 15.325 0.450 15.555 1.580 ;
        RECT 17.565 0.450 17.795 1.580 ;
        RECT 0.000 -0.450 19.600 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 3.320 0.575 4.360 ;
        RECT 2.485 3.320 2.715 4.360 ;
        RECT 4.935 4.120 13.870 4.350 ;
        RECT 4.935 3.320 5.165 4.120 ;
        RECT 0.345 3.090 5.165 3.320 ;
        RECT 13.925 1.810 18.915 2.040 ;
        RECT 0.245 0.910 0.475 1.615 ;
        RECT 2.485 0.910 2.715 1.145 ;
        RECT 4.725 0.910 4.955 1.145 ;
        RECT 6.965 0.910 7.195 1.145 ;
        RECT 9.150 0.910 9.490 1.080 ;
        RECT 11.445 0.910 11.675 1.525 ;
        RECT 13.925 0.910 14.155 1.810 ;
        RECT 0.245 0.680 14.155 0.910 ;
        RECT 16.445 0.805 16.675 1.810 ;
        RECT 18.685 0.805 18.915 1.810 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai31_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai32_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai32_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.720 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.920 2.270 3.260 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.800 2.270 2.140 2.710 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.215 1.015 2.710 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.070 1.770 4.330 2.555 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.190 1.770 5.450 2.555 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.821000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.655 3.015 3.885 4.360 ;
        RECT 3.655 2.785 4.955 3.015 ;
        RECT 4.630 1.140 4.955 2.785 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 6.720 5.490 ;
        RECT 0.345 3.550 0.575 4.590 ;
        RECT 5.745 3.550 5.975 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 7.150 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.150 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.580 ;
        RECT 2.485 0.450 2.715 1.580 ;
        RECT 0.000 -0.450 6.720 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 1.810 3.835 2.040 ;
        RECT 1.365 0.770 1.595 1.810 ;
        RECT 3.605 0.910 3.835 1.810 ;
        RECT 5.845 0.910 6.075 1.580 ;
        RECT 3.605 0.680 6.075 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai32_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai32_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai32_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.320 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.920 2.270 3.260 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.940 2.270 2.690 2.500 ;
        RECT 2.460 2.040 2.690 2.270 ;
        RECT 4.630 2.270 5.450 2.500 ;
        RECT 4.630 2.040 4.890 2.270 ;
        RECT 2.460 1.810 4.890 2.040 ;
        RECT 4.630 1.770 4.890 1.810 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.940 5.910 3.170 ;
        RECT 0.710 2.215 1.015 2.940 ;
        RECT 5.680 2.500 5.910 2.940 ;
        RECT 5.680 2.270 6.570 2.500 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.515 2.215 8.810 2.710 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.430 2.940 10.995 3.170 ;
        RECT 7.430 2.215 7.735 2.940 ;
        RECT 10.765 2.215 10.995 2.940 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.642000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.655 3.645 3.885 4.355 ;
        RECT 9.155 3.645 9.385 4.340 ;
        RECT 3.655 3.415 11.455 3.645 ;
        RECT 11.225 1.985 11.455 3.415 ;
        RECT 7.990 1.755 11.455 1.985 ;
        RECT 7.990 1.140 8.315 1.755 ;
        RECT 10.325 1.140 10.555 1.755 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 12.320 5.490 ;
        RECT 0.345 3.875 0.575 4.590 ;
        RECT 6.865 3.875 7.095 4.590 ;
        RECT 11.345 3.875 11.575 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 12.750 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.750 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.095 ;
        RECT 3.605 0.450 3.835 1.095 ;
        RECT 5.845 0.450 6.075 1.095 ;
        RECT 0.000 -0.450 12.320 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 1.540 4.475 1.565 ;
        RECT 5.055 1.540 7.195 1.565 ;
        RECT 0.245 1.335 7.195 1.540 ;
        RECT 0.245 0.755 0.475 1.335 ;
        RECT 2.485 0.755 2.715 1.335 ;
        RECT 4.370 1.310 5.160 1.335 ;
        RECT 4.725 0.730 5.160 1.310 ;
        RECT 6.965 0.910 7.195 1.335 ;
        RECT 9.205 0.910 9.435 1.525 ;
        RECT 11.685 0.910 11.915 1.565 ;
        RECT 6.965 0.680 11.915 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai32_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai32_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai32_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 24.080 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.670 2.270 13.055 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.080 2.785 4.475 3.015 ;
        RECT 1.080 2.215 1.310 2.785 ;
        RECT 4.245 2.500 4.475 2.785 ;
        RECT 6.870 2.785 9.010 3.015 ;
        RECT 6.870 2.500 7.130 2.785 ;
        RECT 4.245 2.270 7.130 2.500 ;
        RECT 8.780 2.215 9.010 2.785 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.370 2.040 3.600 2.555 ;
        RECT 7.430 2.040 7.690 2.555 ;
        RECT 3.370 1.810 7.690 2.040 ;
        RECT 7.430 1.770 7.690 1.810 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 17.275 2.040 17.615 2.500 ;
        RECT 20.310 2.270 20.785 2.500 ;
        RECT 20.310 2.040 20.570 2.270 ;
        RECT 17.275 1.810 20.570 2.040 ;
        RECT 20.310 1.770 20.570 1.810 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 18.630 2.960 18.890 3.270 ;
        RECT 15.305 2.730 18.075 2.960 ;
        RECT 15.305 2.500 15.535 2.730 ;
        RECT 15.035 2.270 15.535 2.500 ;
        RECT 17.845 2.500 18.075 2.730 ;
        RECT 18.630 2.730 22.590 2.960 ;
        RECT 18.630 2.500 18.860 2.730 ;
        RECT 17.845 2.270 18.860 2.500 ;
        RECT 22.360 2.215 22.590 2.730 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 7.467000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.530 3.320 10.760 3.900 ;
        RECT 12.570 3.320 12.800 3.900 ;
        RECT 16.700 3.770 21.310 4.000 ;
        RECT 16.700 3.450 17.210 3.770 ;
        RECT 16.700 3.420 16.930 3.450 ;
        RECT 14.925 3.320 16.930 3.420 ;
        RECT 10.530 3.190 16.930 3.320 ;
        RECT 21.080 3.420 21.310 3.770 ;
        RECT 21.080 3.190 23.050 3.420 ;
        RECT 10.530 3.090 15.115 3.190 ;
        RECT 15.530 1.540 20.070 1.570 ;
        RECT 22.820 1.565 23.050 3.190 ;
        RECT 20.675 1.540 23.050 1.565 ;
        RECT 15.530 1.340 23.050 1.540 ;
        RECT 15.530 1.140 15.760 1.340 ;
        RECT 17.770 1.140 18.000 1.340 ;
        RECT 19.955 1.335 23.050 1.340 ;
        RECT 19.955 1.140 20.780 1.335 ;
        RECT 22.250 1.140 23.050 1.335 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 24.080 5.490 ;
        RECT 2.590 3.705 2.820 4.590 ;
        RECT 7.070 3.705 7.300 4.590 ;
        RECT 14.510 3.560 14.740 4.590 ;
        RECT 18.840 4.345 19.070 4.590 ;
        RECT 23.280 3.090 23.510 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 24.510 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 24.510 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.570 0.450 1.800 1.110 ;
        RECT 3.810 0.450 4.040 1.110 ;
        RECT 6.050 0.450 6.280 1.110 ;
        RECT 8.290 0.450 8.520 1.110 ;
        RECT 10.530 0.450 10.760 1.110 ;
        RECT 12.770 0.450 13.000 1.110 ;
        RECT 0.000 -0.450 24.080 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 7.530 4.130 14.020 4.360 ;
        RECT 0.500 3.475 0.730 3.900 ;
        RECT 4.880 3.475 5.110 3.900 ;
        RECT 7.530 3.475 7.760 4.130 ;
        RECT 11.550 3.550 11.780 4.130 ;
        RECT 13.790 3.550 14.020 4.130 ;
        RECT 0.500 3.245 7.760 3.475 ;
        RECT 0.500 3.090 0.730 3.245 ;
        RECT 4.880 3.090 5.110 3.245 ;
        RECT 0.450 1.540 7.300 1.580 ;
        RECT 7.820 1.540 14.120 1.580 ;
        RECT 0.450 1.350 14.120 1.540 ;
        RECT 0.450 0.770 0.680 1.350 ;
        RECT 2.690 0.770 2.920 1.350 ;
        RECT 4.930 0.770 5.160 1.350 ;
        RECT 7.170 1.310 7.950 1.350 ;
        RECT 7.170 0.730 7.400 1.310 ;
        RECT 9.410 0.770 9.640 1.350 ;
        RECT 11.650 0.770 11.880 1.350 ;
        RECT 13.890 0.910 14.120 1.350 ;
        RECT 16.650 0.910 16.880 1.110 ;
        RECT 18.890 0.910 19.120 1.110 ;
        RECT 21.130 0.910 21.360 1.105 ;
        RECT 23.370 0.910 23.600 1.580 ;
        RECT 13.890 0.680 23.600 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai32_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai33_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai33_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.070 1.770 4.330 2.555 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.190 2.215 5.450 3.270 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.230 2.270 6.570 2.710 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.920 2.270 3.260 2.710 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.800 2.270 2.140 2.710 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.215 1.015 2.710 ;
    END
  END B3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.401800 ;
    PORT
      LAYER Metal1 ;
        RECT 3.655 3.015 3.885 4.360 ;
        RECT 3.655 2.785 4.900 3.015 ;
        RECT 4.670 1.985 4.900 2.785 ;
        RECT 4.670 1.755 6.540 1.985 ;
        RECT 4.670 1.140 4.955 1.755 ;
        RECT 6.310 1.590 6.540 1.755 ;
        RECT 6.310 1.210 7.195 1.590 ;
        RECT 6.965 0.715 7.195 1.210 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.840 5.490 ;
        RECT 0.345 3.550 0.575 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 8.270 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.270 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.525 ;
        RECT 2.485 0.450 2.715 1.525 ;
        RECT 0.000 -0.450 7.840 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 1.755 3.175 1.985 ;
        RECT 1.365 0.715 1.595 1.755 ;
        RECT 2.945 0.910 3.175 1.755 ;
        RECT 3.605 0.910 3.835 1.525 ;
        RECT 5.845 0.910 6.075 1.525 ;
        RECT 2.945 0.680 6.075 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai33_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai33_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai33_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.560 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.590 2.280 9.930 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.550 2.050 8.890 2.500 ;
        RECT 10.160 2.270 12.220 2.500 ;
        RECT 10.160 2.050 10.390 2.270 ;
        RECT 8.550 1.820 10.390 2.050 ;
        RECT 8.550 1.770 8.810 1.820 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.430 2.940 13.235 3.170 ;
        RECT 7.430 2.215 7.735 2.940 ;
        RECT 13.005 2.215 13.235 2.940 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.920 2.270 3.260 2.710 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.990 2.270 2.650 2.500 ;
        RECT 2.390 2.000 2.650 2.270 ;
        RECT 3.490 2.270 5.500 2.500 ;
        RECT 3.490 2.000 3.720 2.270 ;
        RECT 2.390 1.770 3.720 2.000 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.940 5.960 3.170 ;
        RECT 0.710 2.215 1.015 2.940 ;
        RECT 5.730 2.500 5.960 2.940 ;
        RECT 5.730 2.270 6.620 2.500 ;
    END
  END B3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.328400 ;
    PORT
      LAYER Metal1 ;
        RECT 3.655 3.630 3.885 4.360 ;
        RECT 10.275 3.630 10.505 4.360 ;
        RECT 3.655 3.400 13.695 3.630 ;
        RECT 13.465 1.590 13.695 3.400 ;
        RECT 10.230 1.480 13.695 1.590 ;
        RECT 8.030 1.250 13.695 1.480 ;
        RECT 10.230 1.140 10.555 1.250 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 14.560 5.490 ;
        RECT 0.345 3.860 0.575 4.590 ;
        RECT 6.915 3.860 7.145 4.590 ;
        RECT 13.585 3.860 13.815 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 14.990 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.990 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.455 ;
        RECT 3.605 0.450 3.835 1.000 ;
        RECT 5.845 0.450 6.075 1.565 ;
        RECT 0.000 -0.450 14.560 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 1.685 2.160 1.915 ;
        RECT 0.245 0.845 0.475 1.685 ;
        RECT 1.930 1.540 2.160 1.685 ;
        RECT 4.725 1.795 7.195 2.025 ;
        RECT 4.725 1.540 4.955 1.795 ;
        RECT 1.930 1.310 4.955 1.540 ;
        RECT 1.930 0.730 2.715 1.310 ;
        RECT 4.725 0.730 4.955 1.310 ;
        RECT 6.965 1.020 7.195 1.795 ;
        RECT 6.965 0.910 9.435 1.020 ;
        RECT 11.445 0.910 13.915 1.020 ;
        RECT 6.965 0.680 13.915 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai33_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai33_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai33_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.560 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 15.325 2.190 17.850 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.120 2.495 27.195 2.725 ;
        RECT 19.120 2.270 19.460 2.495 ;
        RECT 21.990 2.270 22.820 2.495 ;
        RECT 26.965 2.215 27.195 2.495 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.690 2.040 20.580 2.265 ;
        RECT 24.720 2.040 25.060 2.265 ;
        RECT 19.690 1.810 25.060 2.040 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.325 2.190 12.795 2.710 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.820 2.650 7.030 2.880 ;
        RECT 0.820 2.190 1.160 2.650 ;
        RECT 4.040 2.270 4.380 2.650 ;
        RECT 6.800 2.500 7.030 2.650 ;
        RECT 6.800 2.270 8.860 2.500 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 2.000 2.170 2.420 ;
        RECT 4.610 2.190 6.570 2.420 ;
        RECT 4.610 2.000 4.840 2.190 ;
        RECT 1.830 1.770 4.840 2.000 ;
    END
  END B3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 8.382299 ;
    PORT
      LAYER Metal1 ;
        RECT 10.325 3.185 10.555 3.830 ;
        RECT 12.565 3.185 13.850 3.830 ;
        RECT 15.325 3.185 15.555 3.460 ;
        RECT 17.515 3.185 17.745 3.460 ;
        RECT 10.325 2.955 27.655 3.185 ;
        RECT 27.425 1.530 27.655 2.955 ;
        RECT 15.270 1.300 27.655 1.530 ;
        RECT 17.510 1.140 17.850 1.300 ;
        RECT 19.750 1.140 20.090 1.300 ;
        RECT 21.990 1.140 22.330 1.300 ;
        RECT 24.230 1.140 24.570 1.300 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 28.560 5.490 ;
        RECT 2.385 3.580 2.615 4.590 ;
        RECT 6.865 3.580 7.095 4.590 ;
        RECT 20.875 4.150 21.105 4.590 ;
        RECT 25.355 3.875 25.585 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 28.990 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 28.990 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.070 ;
        RECT 3.605 0.450 3.835 1.070 ;
        RECT 5.845 0.450 6.075 1.070 ;
        RECT 8.085 0.450 8.315 1.070 ;
        RECT 10.325 0.450 10.555 1.070 ;
        RECT 12.565 0.450 12.795 1.070 ;
        RECT 0.000 -0.450 28.560 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 7.325 4.060 13.870 4.290 ;
        RECT 0.295 3.350 0.525 3.930 ;
        RECT 4.675 3.350 4.905 3.930 ;
        RECT 7.325 3.350 7.555 4.060 ;
        RECT 11.345 3.480 11.575 4.060 ;
        RECT 14.305 3.690 23.345 3.920 ;
        RECT 14.305 3.480 14.535 3.690 ;
        RECT 16.445 3.480 16.675 3.690 ;
        RECT 23.115 3.645 23.345 3.690 ;
        RECT 27.545 3.645 27.775 4.225 ;
        RECT 23.115 3.415 27.775 3.645 ;
        RECT 0.295 3.120 7.555 3.350 ;
        RECT 0.245 1.310 14.430 1.540 ;
        RECT 0.245 0.730 0.475 1.310 ;
        RECT 2.485 0.730 2.715 1.310 ;
        RECT 4.725 0.730 4.955 1.310 ;
        RECT 6.965 0.730 7.195 1.310 ;
        RECT 9.205 0.730 9.435 1.310 ;
        RECT 11.445 0.730 11.675 1.310 ;
        RECT 14.200 1.070 14.430 1.310 ;
        RECT 14.200 0.910 16.675 1.070 ;
        RECT 18.630 0.910 18.970 1.015 ;
        RECT 20.870 0.910 21.210 1.015 ;
        RECT 23.110 0.910 23.450 1.015 ;
        RECT 25.405 0.910 27.875 1.070 ;
        RECT 14.200 0.680 27.875 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai33_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai211_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai211_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 2.270 2.170 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.215 1.015 2.710 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 2.270 3.290 2.710 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.990 2.270 4.330 2.710 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.498800 ;
    PORT
      LAYER Metal1 ;
        RECT 2.385 3.320 2.615 4.360 ;
        RECT 4.605 3.320 4.835 4.360 ;
        RECT 1.270 3.090 4.835 3.320 ;
        RECT 1.270 1.140 1.595 3.090 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.600 5.490 ;
        RECT 0.345 3.550 0.575 4.590 ;
        RECT 3.585 3.550 3.815 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 4.605 0.450 4.835 1.655 ;
        RECT 0.000 -0.450 5.600 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 0.910 0.475 1.655 ;
        RECT 2.485 0.910 2.715 1.655 ;
        RECT 0.245 0.680 2.715 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai211_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai211_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai211_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.795 2.215 2.090 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.200 2.940 2.620 3.170 ;
        RECT 1.200 2.270 1.540 2.940 ;
        RECT 2.390 2.710 2.620 2.940 ;
        RECT 2.390 2.270 4.330 2.710 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.330 2.940 8.535 3.170 ;
        RECT 5.330 2.270 5.670 2.940 ;
        RECT 6.870 2.215 8.535 2.940 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.230 2.270 6.570 2.710 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.025800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.865 4.070 2.665 4.360 ;
        RECT 0.865 3.580 1.095 4.070 ;
        RECT 0.740 3.375 1.095 3.580 ;
        RECT 2.435 3.630 2.665 4.070 ;
        RECT 5.825 3.630 6.055 4.360 ;
        RECT 7.865 3.630 8.095 4.360 ;
        RECT 2.435 3.400 8.095 3.630 ;
        RECT 0.740 1.570 0.970 3.375 ;
        RECT 0.740 1.340 3.890 1.570 ;
        RECT 0.740 1.140 1.595 1.340 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 9.520 5.490 ;
        RECT 0.345 3.860 0.575 4.590 ;
        RECT 4.625 3.860 4.855 4.590 ;
        RECT 6.845 3.860 7.075 4.590 ;
        RECT 8.885 3.860 9.115 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 9.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 6.845 0.450 7.075 1.525 ;
        RECT 0.000 -0.450 9.520 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 4.725 1.755 9.115 1.985 ;
        RECT 0.245 0.910 0.475 1.580 ;
        RECT 4.725 1.110 4.955 1.755 ;
        RECT 2.485 0.910 4.955 1.110 ;
        RECT 0.245 0.680 4.955 0.910 ;
        RECT 8.885 0.770 9.115 1.755 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai211_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai211_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai211_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.920 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.060 2.390 3.770 2.620 ;
        RECT 3.510 2.100 3.770 2.390 ;
        RECT 4.560 2.390 6.620 2.620 ;
        RECT 4.560 2.100 4.790 2.390 ;
        RECT 3.510 1.870 4.790 2.100 ;
        RECT 3.510 1.770 3.770 1.870 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.870 2.850 7.080 3.080 ;
        RECT 0.870 2.390 1.210 2.850 ;
        RECT 4.070 2.330 4.330 2.850 ;
        RECT 6.850 2.620 7.080 2.850 ;
        RECT 6.850 2.390 8.810 2.620 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.088000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.670 2.850 15.470 3.080 ;
        RECT 9.670 2.330 9.955 2.850 ;
        RECT 12.875 2.335 13.105 2.850 ;
        RECT 15.240 2.620 15.470 2.850 ;
        RECT 15.240 2.390 17.150 2.620 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.088000 ;
    PORT
      LAYER Metal1 ;
        RECT 11.850 2.390 12.500 2.620 ;
        RECT 12.270 2.155 12.500 2.390 ;
        RECT 13.335 2.390 15.010 2.620 ;
        RECT 12.270 2.000 12.730 2.155 ;
        RECT 13.335 2.000 13.565 2.390 ;
        RECT 12.330 1.770 13.565 2.000 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 7.960100 ;
    PORT
      LAYER Metal1 ;
        RECT 2.485 3.540 2.715 4.360 ;
        RECT 6.915 3.540 7.145 4.360 ;
        RECT 10.305 3.540 10.535 4.120 ;
        RECT 12.345 3.830 12.575 4.360 ;
        RECT 11.910 3.540 12.575 3.830 ;
        RECT 14.385 3.540 14.615 4.345 ;
        RECT 16.425 3.540 16.655 4.360 ;
        RECT 0.410 3.310 16.655 3.540 ;
        RECT 0.410 1.950 0.640 3.310 ;
        RECT 0.410 1.720 3.280 1.950 ;
        RECT 1.365 1.140 1.595 1.720 ;
        RECT 3.050 1.540 3.280 1.720 ;
        RECT 5.980 1.600 8.315 1.830 ;
        RECT 5.980 1.580 6.210 1.600 ;
        RECT 3.990 1.540 6.210 1.580 ;
        RECT 3.050 1.350 6.210 1.540 ;
        RECT 3.050 1.140 4.120 1.350 ;
        RECT 5.845 1.140 6.210 1.350 ;
        RECT 8.085 1.140 8.315 1.600 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.920 5.490 ;
        RECT 0.345 3.770 0.575 4.590 ;
        RECT 4.675 3.770 4.905 4.590 ;
        RECT 9.105 3.770 9.335 4.590 ;
        RECT 11.325 3.770 11.555 4.590 ;
        RECT 13.365 3.770 13.595 4.590 ;
        RECT 15.405 3.770 15.635 4.590 ;
        RECT 17.445 3.770 17.675 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 18.350 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 18.350 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 11.325 0.450 11.555 1.265 ;
        RECT 15.405 0.450 15.635 1.490 ;
        RECT 0.000 -0.450 17.920 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 9.205 1.540 12.100 1.725 ;
        RECT 13.795 1.720 17.675 1.950 ;
        RECT 13.795 1.540 14.025 1.720 ;
        RECT 9.205 1.495 14.025 1.540 ;
        RECT 0.245 0.910 0.475 1.490 ;
        RECT 2.430 0.910 2.770 0.965 ;
        RECT 4.670 0.910 5.010 0.965 ;
        RECT 6.910 0.910 7.250 0.965 ;
        RECT 9.205 0.910 9.435 1.495 ;
        RECT 11.870 1.310 14.025 1.495 ;
        RECT 0.245 0.680 9.435 0.910 ;
        RECT 13.365 0.680 13.595 1.310 ;
        RECT 17.445 0.680 17.675 1.720 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai211_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai221_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai221_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.720 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.190 1.770 5.455 2.555 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.070 2.215 4.435 2.710 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 2.150 2.090 2.710 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 1.015 2.555 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 2.270 3.290 2.710 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.661600 ;
    PORT
      LAYER Metal1 ;
        RECT 2.565 3.320 2.795 4.360 ;
        RECT 5.805 3.320 6.035 4.360 ;
        RECT 2.565 3.090 6.035 3.320 ;
        RECT 4.665 1.590 4.895 3.090 ;
        RECT 4.630 1.480 4.895 1.590 ;
        RECT 4.630 1.140 5.015 1.480 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 6.720 5.490 ;
        RECT 0.345 3.550 0.575 4.590 ;
        RECT 3.585 3.550 3.815 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 7.150 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.150 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.070 ;
        RECT 0.000 -0.450 6.720 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 1.310 2.715 1.540 ;
        RECT 0.245 0.730 0.475 1.310 ;
        RECT 2.485 0.730 2.715 1.310 ;
        RECT 3.665 0.910 3.895 1.540 ;
        RECT 5.905 0.910 6.135 1.540 ;
        RECT 3.665 0.680 6.135 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai221_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai221_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai221_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.320 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.530 2.890 9.305 3.270 ;
        RECT 7.530 2.215 7.760 2.890 ;
        RECT 9.075 2.500 9.305 2.890 ;
        RECT 9.075 2.270 11.140 2.500 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.990 2.215 8.845 2.555 ;
        RECT 7.990 1.770 8.250 2.215 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 2.150 3.210 2.710 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.270 2.940 4.805 3.170 ;
        RECT 2.270 2.555 2.500 2.940 ;
        RECT 1.210 2.325 2.500 2.555 ;
        RECT 4.575 2.555 4.805 2.940 ;
        RECT 1.210 1.830 2.165 2.325 ;
        RECT 4.575 2.215 5.425 2.555 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.980 3.580 5.265 3.630 ;
        RECT 0.710 3.400 5.265 3.580 ;
        RECT 0.710 3.350 2.125 3.400 ;
        RECT 0.710 1.770 0.970 3.350 ;
        RECT 5.035 3.015 5.265 3.400 ;
        RECT 5.035 2.785 6.625 3.015 ;
        RECT 6.395 2.215 6.625 2.785 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 5.216500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.295 4.040 0.525 4.360 ;
        RECT 3.535 4.090 3.765 4.360 ;
        RECT 1.690 4.040 5.725 4.090 ;
        RECT 0.295 3.860 5.725 4.040 ;
        RECT 0.295 3.810 1.835 3.860 ;
        RECT 5.495 3.780 5.725 3.860 ;
        RECT 6.975 3.780 7.205 4.360 ;
        RECT 5.495 3.550 11.665 3.780 ;
        RECT 10.790 2.890 11.665 3.550 ;
        RECT 11.435 1.985 11.665 2.890 ;
        RECT 8.480 1.755 11.665 1.985 ;
        RECT 8.480 1.540 8.710 1.755 ;
        RECT 8.120 1.310 8.710 1.540 ;
        RECT 10.415 1.140 10.645 1.755 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 12.320 5.490 ;
        RECT 1.315 4.270 1.545 4.590 ;
        RECT 5.955 4.020 6.185 4.590 ;
        RECT 9.245 4.020 9.475 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 12.750 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.750 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.460 0.450 2.800 0.640 ;
        RECT 4.700 0.450 5.040 0.640 ;
        RECT 0.000 -0.450 12.320 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 1.100 0.475 1.525 ;
        RECT 1.340 1.330 6.160 1.560 ;
        RECT 7.055 1.100 7.285 1.190 ;
        RECT 0.245 0.910 7.285 1.100 ;
        RECT 9.295 0.910 9.525 1.525 ;
        RECT 11.535 0.910 11.765 1.525 ;
        RECT 0.245 0.870 11.765 0.910 ;
        RECT 0.245 0.715 0.475 0.870 ;
        RECT 7.055 0.680 11.765 0.870 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai221_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai221_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai221_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 24.080 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 15.030 3.040 21.190 3.270 ;
        RECT 15.030 2.270 15.370 3.040 ;
        RECT 19.140 2.890 21.190 3.040 ;
        RECT 19.140 2.215 19.370 2.890 ;
        RECT 20.960 2.500 21.190 2.890 ;
        RECT 20.960 2.270 22.970 2.500 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 17.270 2.270 17.770 2.500 ;
        RECT 17.510 1.985 17.770 2.270 ;
        RECT 19.600 2.270 20.730 2.500 ;
        RECT 19.600 1.985 19.830 2.270 ;
        RECT 17.510 1.755 19.830 1.985 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.870 2.730 7.080 2.960 ;
        RECT 0.870 2.270 1.210 2.730 ;
        RECT 4.070 2.270 4.410 2.730 ;
        RECT 6.850 2.500 7.080 2.730 ;
        RECT 6.850 2.270 8.860 2.500 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.060 2.270 3.630 2.500 ;
        RECT 3.400 2.175 3.630 2.270 ;
        RECT 4.640 2.270 6.620 2.500 ;
        RECT 3.400 2.040 3.860 2.175 ;
        RECT 4.640 2.040 4.870 2.270 ;
        RECT 3.400 2.020 4.870 2.040 ;
        RECT 3.460 1.770 4.870 2.020 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.088000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.990 2.270 13.570 2.710 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 10.615000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.345 3.420 0.575 4.360 ;
        RECT 4.675 3.730 4.905 4.360 ;
        RECT 9.155 3.730 9.385 4.360 ;
        RECT 12.165 3.730 12.395 4.360 ;
        RECT 14.305 3.730 14.535 4.360 ;
        RECT 18.570 3.730 19.065 4.360 ;
        RECT 23.265 3.730 23.495 4.360 ;
        RECT 4.675 3.500 23.495 3.730 ;
        RECT 4.675 3.420 4.905 3.500 ;
        RECT 0.345 3.190 4.905 3.420 ;
        RECT 23.200 1.970 23.495 3.500 ;
        RECT 20.060 1.740 23.495 1.970 ;
        RECT 20.060 1.520 20.290 1.740 ;
        RECT 15.525 1.290 20.290 1.520 ;
        RECT 15.525 1.140 15.755 1.290 ;
        RECT 17.710 1.140 18.050 1.290 ;
        RECT 20.005 1.140 20.290 1.290 ;
        RECT 22.245 1.140 22.475 1.740 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 24.080 5.490 ;
        RECT 2.435 3.650 2.665 4.590 ;
        RECT 6.915 3.960 7.145 4.590 ;
        RECT 10.945 3.960 11.175 4.590 ;
        RECT 13.185 3.960 13.415 4.590 ;
        RECT 16.595 3.960 16.825 4.590 ;
        RECT 21.075 3.960 21.305 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 24.510 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 24.510 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.510 ;
        RECT 2.485 0.450 2.715 1.510 ;
        RECT 4.725 0.450 4.955 1.040 ;
        RECT 6.965 0.450 7.195 1.040 ;
        RECT 9.205 0.450 9.435 1.040 ;
        RECT 0.000 -0.450 24.080 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 1.740 3.175 1.970 ;
        RECT 1.365 0.700 1.595 1.740 ;
        RECT 2.945 1.510 3.175 1.740 ;
        RECT 2.945 1.280 13.515 1.510 ;
        RECT 3.605 0.700 3.835 1.280 ;
        RECT 5.845 0.700 6.075 1.280 ;
        RECT 8.085 0.700 8.315 1.280 ;
        RECT 10.990 1.140 11.330 1.280 ;
        RECT 13.285 1.140 13.515 1.280 ;
        RECT 9.925 0.910 10.155 1.040 ;
        RECT 12.110 0.910 12.450 0.985 ;
        RECT 14.350 0.910 14.690 0.985 ;
        RECT 16.590 0.910 16.930 0.985 ;
        RECT 18.830 0.910 19.170 0.985 ;
        RECT 21.125 0.910 21.355 1.510 ;
        RECT 23.365 0.910 23.595 1.510 ;
        RECT 9.925 0.680 23.595 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai221_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai222_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai222_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.400 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.870 2.270 7.290 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 2.270 6.180 2.710 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 1.770 3.980 2.500 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.630 2.270 5.050 2.710 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 2.150 2.090 2.710 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.215 1.015 2.710 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.943800 ;
    PORT
      LAYER Metal1 ;
        RECT 3.255 3.830 3.485 4.360 ;
        RECT 7.585 3.830 7.815 4.360 ;
        RECT 3.255 3.550 7.815 3.830 ;
        RECT 3.255 3.450 6.640 3.550 ;
        RECT 6.410 1.480 6.640 3.450 ;
        RECT 6.410 1.140 6.795 1.480 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 8.400 5.490 ;
        RECT 0.345 3.550 0.575 4.590 ;
        RECT 5.345 4.060 5.575 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 8.830 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.830 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.205 ;
        RECT 0.000 -0.450 8.400 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 1.540 3.305 1.665 ;
        RECT 1.365 1.435 4.555 1.540 ;
        RECT 1.365 0.680 1.595 1.435 ;
        RECT 3.100 1.310 4.555 1.435 ;
        RECT 4.325 1.140 4.555 1.310 ;
        RECT 3.150 0.910 3.490 0.965 ;
        RECT 5.445 0.910 5.675 1.490 ;
        RECT 7.685 0.910 7.915 1.490 ;
        RECT 3.150 0.680 7.915 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai222_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai222_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai222_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.120 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.605 2.940 12.500 3.170 ;
        RECT 10.605 2.215 10.835 2.940 ;
        RECT 12.270 2.710 12.500 2.940 ;
        RECT 12.270 2.215 14.005 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 11.350 2.215 11.715 2.710 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.190 3.040 9.525 3.270 ;
        RECT 5.190 2.215 6.165 3.040 ;
        RECT 9.295 2.215 9.525 3.040 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.870 2.215 7.285 2.710 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.925 2.785 4.330 3.015 ;
        RECT 0.925 2.215 1.155 2.785 ;
        RECT 4.070 1.770 4.330 2.785 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.090 2.555 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.570000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.345 3.550 0.575 4.360 ;
        RECT 4.675 3.730 4.905 4.360 ;
        RECT 8.490 4.130 10.105 4.360 ;
        RECT 8.490 3.730 8.870 4.130 ;
        RECT 4.675 3.550 8.870 3.730 ;
        RECT 0.345 3.500 8.870 3.550 ;
        RECT 9.875 3.630 10.105 4.130 ;
        RECT 14.355 3.630 14.585 4.360 ;
        RECT 0.345 3.320 4.900 3.500 ;
        RECT 9.875 3.400 14.585 3.630 ;
        RECT 14.355 1.950 14.585 3.400 ;
        RECT 11.045 1.720 14.585 1.950 ;
        RECT 11.045 1.140 11.275 1.720 ;
        RECT 13.285 1.140 13.515 1.720 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 15.120 5.490 ;
        RECT 2.435 3.780 2.665 4.590 ;
        RECT 7.635 3.960 7.865 4.590 ;
        RECT 12.115 3.860 12.345 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 15.550 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 15.550 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.655 ;
        RECT 2.485 0.450 2.715 0.695 ;
        RECT 4.725 0.450 4.955 0.695 ;
        RECT 0.000 -0.450 15.120 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 1.140 9.035 1.540 ;
        RECT 1.365 0.925 3.835 1.140 ;
        RECT 1.365 0.730 1.595 0.925 ;
        RECT 3.605 0.730 3.835 0.925 ;
        RECT 9.925 0.910 10.155 1.575 ;
        RECT 12.165 0.910 12.395 1.490 ;
        RECT 14.405 0.910 14.635 1.490 ;
        RECT 5.390 0.680 14.635 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai222_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai222_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai222_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.560 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.190 2.000 19.660 2.500 ;
        RECT 22.685 2.000 22.915 2.145 ;
        RECT 27.165 2.000 27.395 2.555 ;
        RECT 19.190 1.770 27.395 2.000 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 21.700 2.480 25.260 2.710 ;
        RECT 21.700 2.270 22.040 2.480 ;
        RECT 23.110 2.270 25.260 2.480 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.605 3.040 18.540 3.270 ;
        RECT 10.605 2.890 14.060 3.040 ;
        RECT 10.605 2.215 10.835 2.890 ;
        RECT 13.720 2.270 14.060 2.890 ;
        RECT 18.200 2.270 18.540 3.040 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.740 2.270 13.290 2.500 ;
        RECT 13.030 2.000 13.290 2.270 ;
        RECT 14.290 2.270 16.250 2.500 ;
        RECT 14.290 2.000 14.520 2.270 ;
        RECT 13.030 1.770 14.520 2.000 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.875 2.785 7.080 3.015 ;
        RECT 0.875 2.215 1.105 2.785 ;
        RECT 4.040 2.270 4.380 2.785 ;
        RECT 6.850 2.500 7.080 2.785 ;
        RECT 6.850 2.270 8.860 2.500 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.165 2.215 3.770 2.555 ;
        RECT 3.510 2.000 3.770 2.215 ;
        RECT 4.610 2.270 6.620 2.500 ;
        RECT 4.610 2.000 4.840 2.270 ;
        RECT 3.510 1.770 4.840 2.000 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 11.529600 ;
    PORT
      LAYER Metal1 ;
        RECT 0.295 3.475 0.525 4.360 ;
        RECT 4.675 3.550 4.905 4.360 ;
        RECT 9.155 3.730 9.385 4.360 ;
        RECT 12.970 3.730 14.585 4.360 ;
        RECT 18.835 3.730 19.065 4.360 ;
        RECT 9.155 3.550 19.065 3.730 ;
        RECT 4.675 3.500 19.065 3.550 ;
        RECT 4.675 3.475 9.380 3.500 ;
        RECT 0.295 3.245 9.380 3.475 ;
        RECT 18.835 3.320 19.065 3.500 ;
        RECT 23.265 3.320 23.495 4.360 ;
        RECT 27.745 3.320 27.975 4.360 ;
        RECT 18.835 3.090 27.975 3.320 ;
        RECT 27.745 1.515 27.975 3.090 ;
        RECT 20.005 1.285 27.975 1.515 ;
        RECT 20.005 1.140 20.235 1.285 ;
        RECT 22.190 1.140 22.530 1.285 ;
        RECT 24.430 1.140 24.770 1.285 ;
        RECT 26.670 1.140 27.010 1.285 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 28.560 5.490 ;
        RECT 2.435 3.705 2.665 4.590 ;
        RECT 6.915 3.780 7.145 4.590 ;
        RECT 12.115 3.960 12.345 4.590 ;
        RECT 16.595 3.960 16.825 4.590 ;
        RECT 21.075 3.550 21.305 4.590 ;
        RECT 25.555 3.550 25.785 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 28.990 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 28.990 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.525 ;
        RECT 2.485 0.450 2.715 1.525 ;
        RECT 4.725 0.450 4.955 1.055 ;
        RECT 6.965 0.450 7.195 1.525 ;
        RECT 9.205 0.450 9.435 1.525 ;
        RECT 0.000 -0.450 28.560 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 1.755 3.280 1.985 ;
        RECT 1.365 0.715 1.595 1.755 ;
        RECT 3.050 1.525 3.280 1.755 ;
        RECT 5.845 1.755 11.220 1.985 ;
        RECT 5.845 1.525 6.075 1.755 ;
        RECT 3.050 1.295 6.075 1.525 ;
        RECT 3.605 0.715 3.835 1.295 ;
        RECT 5.845 0.715 6.075 1.295 ;
        RECT 8.085 0.715 8.315 1.755 ;
        RECT 9.925 0.910 10.155 1.525 ;
        RECT 10.990 1.520 11.220 1.755 ;
        RECT 15.580 1.755 17.995 1.985 ;
        RECT 15.580 1.520 15.810 1.755 ;
        RECT 10.990 1.290 15.810 1.520 ;
        RECT 10.990 1.140 11.275 1.290 ;
        RECT 13.230 1.140 13.570 1.290 ;
        RECT 15.525 1.140 15.810 1.290 ;
        RECT 12.110 0.910 12.450 1.000 ;
        RECT 14.350 0.910 14.690 1.000 ;
        RECT 16.645 0.910 16.875 1.525 ;
        RECT 17.765 1.140 17.995 1.755 ;
        RECT 18.885 0.910 19.115 1.525 ;
        RECT 21.070 0.910 21.410 1.000 ;
        RECT 23.310 0.910 23.650 1.000 ;
        RECT 25.550 0.910 25.890 1.000 ;
        RECT 27.845 0.910 28.075 1.055 ;
        RECT 9.925 0.680 28.075 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai222_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__or2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.853500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.215 1.070 3.270 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.853500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.210 2.090 2.555 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.800 1.590 4.130 4.360 ;
        RECT 3.510 1.210 4.130 1.590 ;
        RECT 3.900 0.680 4.130 1.210 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 4.480 5.490 ;
        RECT 2.780 3.790 3.010 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 4.910 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 0.450 0.530 0.995 ;
        RECT 2.780 0.450 3.010 0.995 ;
        RECT 0.000 -0.450 4.480 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 3.845 2.550 4.075 ;
        RECT 2.320 2.500 2.550 3.845 ;
        RECT 2.320 2.270 3.505 2.500 ;
        RECT 2.320 0.940 2.550 2.270 ;
        RECT 1.365 0.710 2.550 0.940 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or2_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__or2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.270 1.070 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.795 2.215 2.090 2.710 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.729500 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 0.680 3.835 4.360 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.600 5.490 ;
        RECT 2.435 3.550 2.665 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 4.725 0.450 4.955 1.490 ;
        RECT 0.000 -0.450 5.600 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 3.320 0.575 4.360 ;
        RECT 0.345 3.090 3.205 3.320 ;
        RECT 2.975 1.950 3.205 3.090 ;
        RECT 1.365 1.720 3.205 1.950 ;
        RECT 1.365 0.680 1.595 1.720 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or2_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__or2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.800 2.270 2.140 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.870 2.940 4.275 3.170 ;
        RECT 0.870 2.270 1.210 2.940 ;
        RECT 2.390 2.215 4.275 2.940 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.550500 ;
    PORT
      LAYER Metal1 ;
        RECT 6.085 3.320 6.315 4.360 ;
        RECT 8.175 3.320 8.405 4.360 ;
        RECT 6.085 3.090 8.405 3.320 ;
        RECT 7.620 1.590 7.850 3.090 ;
        RECT 5.985 1.490 7.850 1.590 ;
        RECT 5.985 1.210 8.455 1.490 ;
        RECT 5.985 0.680 6.215 1.210 ;
        RECT 8.225 0.680 8.455 1.210 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 10.080 5.490 ;
        RECT 0.345 3.550 0.575 4.590 ;
        RECT 4.965 3.550 5.195 4.590 ;
        RECT 7.105 3.550 7.335 4.590 ;
        RECT 9.245 3.550 9.475 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 10.510 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 10.510 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 4.725 0.450 4.955 1.490 ;
        RECT 7.105 0.450 7.335 0.980 ;
        RECT 9.345 0.450 9.575 1.490 ;
        RECT 0.000 -0.450 10.080 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 2.535 3.630 2.765 4.360 ;
        RECT 2.535 3.400 4.735 3.630 ;
        RECT 4.505 2.500 4.735 3.400 ;
        RECT 4.505 2.270 7.390 2.500 ;
        RECT 4.505 1.970 4.735 2.270 ;
        RECT 1.365 1.740 4.735 1.970 ;
        RECT 1.365 0.680 1.595 1.740 ;
        RECT 3.605 0.680 3.835 1.740 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or2_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__or3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.160 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.772500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.785 2.150 1.015 2.555 ;
        RECT 0.150 1.770 1.015 2.150 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.772500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.090 2.555 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.772500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 2.215 3.335 2.710 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.045 0.680 5.450 4.360 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 6.160 5.490 ;
        RECT 4.025 3.790 4.255 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.590 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.590 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 0.860 ;
        RECT 3.785 0.450 4.015 0.860 ;
        RECT 0.000 -0.450 6.160 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.290 3.845 3.795 4.075 ;
        RECT 3.565 2.500 3.795 3.845 ;
        RECT 3.565 2.270 4.750 2.500 ;
        RECT 3.565 1.320 3.795 2.270 ;
        RECT 0.245 1.090 3.795 1.320 ;
        RECT 0.245 0.680 0.475 1.090 ;
        RECT 2.485 0.680 2.715 1.090 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or3_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__or3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.720 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.545000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.270 1.070 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.545000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.795 2.215 2.090 2.710 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.545000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.915 2.215 3.210 2.710 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.729500 ;
    PORT
      LAYER Metal1 ;
        RECT 4.630 2.890 5.135 4.360 ;
        RECT 4.905 0.680 5.135 2.890 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 6.720 5.490 ;
        RECT 3.555 3.550 3.785 4.590 ;
        RECT 5.925 3.550 6.155 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 7.150 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.150 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.385 ;
        RECT 3.605 0.450 3.835 1.385 ;
        RECT 6.025 0.450 6.255 1.490 ;
        RECT 0.000 -0.450 6.720 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 3.320 0.575 4.360 ;
        RECT 0.345 3.090 3.670 3.320 ;
        RECT 3.440 2.555 3.670 3.090 ;
        RECT 3.440 2.215 4.505 2.555 ;
        RECT 3.440 1.845 3.670 2.215 ;
        RECT 0.245 1.615 3.670 1.845 ;
        RECT 0.245 0.680 0.475 1.615 ;
        RECT 2.485 0.680 2.715 1.615 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or3_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__or3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.320 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.090000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.920 2.270 3.260 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.090000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 2.000 2.170 2.500 ;
        RECT 3.490 2.270 5.500 2.500 ;
        RECT 3.490 2.000 3.720 2.270 ;
        RECT 1.830 1.770 3.720 2.000 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.090000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.940 6.570 3.170 ;
        RECT 0.710 2.270 1.070 2.940 ;
        RECT 6.230 2.270 6.570 2.940 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.459000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.315 3.630 8.545 4.360 ;
        RECT 10.455 3.630 10.685 4.360 ;
        RECT 8.315 3.400 10.685 3.630 ;
        RECT 9.900 1.590 10.130 3.400 ;
        RECT 8.265 1.490 10.130 1.590 ;
        RECT 8.265 1.210 10.735 1.490 ;
        RECT 8.265 0.680 8.495 1.210 ;
        RECT 10.505 0.680 10.735 1.210 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 12.320 5.490 ;
        RECT 0.345 3.860 0.575 4.590 ;
        RECT 6.865 3.860 7.095 4.590 ;
        RECT 9.335 3.860 9.565 4.590 ;
        RECT 11.525 3.860 11.755 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 12.750 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.750 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.385 ;
        RECT 2.485 0.450 2.715 0.915 ;
        RECT 4.725 0.450 4.955 0.915 ;
        RECT 6.965 0.450 7.195 0.915 ;
        RECT 9.385 0.450 9.615 0.915 ;
        RECT 11.625 0.450 11.855 1.385 ;
        RECT 0.000 -0.450 12.320 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.655 3.630 3.885 4.360 ;
        RECT 3.655 3.400 7.030 3.630 ;
        RECT 6.800 2.500 7.030 3.400 ;
        RECT 6.800 2.270 9.670 2.500 ;
        RECT 6.800 1.375 7.030 2.270 ;
        RECT 1.365 1.145 7.030 1.375 ;
        RECT 1.365 0.680 1.595 1.145 ;
        RECT 3.605 0.680 3.835 1.145 ;
        RECT 5.845 0.680 6.075 1.145 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or3_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__or4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.694500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.785 2.150 1.015 2.555 ;
        RECT 0.150 1.770 1.015 2.150 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.694500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.215 2.555 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.694500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 1.770 3.385 2.555 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.694500 ;
    PORT
      LAYER Metal1 ;
        RECT 4.345 1.590 4.575 2.555 ;
        RECT 4.070 1.210 4.575 1.590 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.285 0.680 6.615 4.360 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.280 5.490 ;
        RECT 5.265 3.790 5.495 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 7.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.015 ;
        RECT 2.665 0.450 2.895 1.015 ;
        RECT 5.265 0.450 5.495 0.940 ;
        RECT 0.000 -0.450 7.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.290 3.845 5.035 4.075 ;
        RECT 4.805 2.500 5.035 3.845 ;
        RECT 4.805 2.270 5.990 2.500 ;
        RECT 1.545 1.245 3.840 1.475 ;
        RECT 1.545 0.680 1.775 1.245 ;
        RECT 3.610 0.930 3.840 1.245 ;
        RECT 4.805 0.930 5.035 2.270 ;
        RECT 3.610 0.700 5.035 0.930 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or4_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__or4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.270 1.070 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.090 2.555 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.390 2.270 3.260 2.710 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 2.270 4.380 2.710 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.729500 ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 2.890 6.255 4.360 ;
        RECT 6.025 0.680 6.255 2.890 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.840 5.490 ;
        RECT 4.675 3.550 4.905 4.590 ;
        RECT 7.045 3.550 7.275 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 8.270 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.270 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.020 ;
        RECT 2.485 0.450 2.715 1.020 ;
        RECT 4.725 0.450 4.955 1.020 ;
        RECT 7.145 0.450 7.375 1.490 ;
        RECT 0.000 -0.450 7.840 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 3.320 0.575 4.360 ;
        RECT 0.345 3.090 4.840 3.320 ;
        RECT 4.610 2.555 4.840 3.090 ;
        RECT 4.610 2.215 5.625 2.555 ;
        RECT 4.610 1.480 4.840 2.215 ;
        RECT 1.365 1.250 4.840 1.480 ;
        RECT 1.365 0.680 1.595 1.250 ;
        RECT 3.605 0.680 3.835 1.250 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or4_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__or4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or4_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.560 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.035 2.215 4.330 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.440 2.940 4.860 3.170 ;
        RECT 3.440 2.500 3.670 2.940 ;
        RECT 3.060 2.270 3.670 2.500 ;
        RECT 4.630 2.710 4.860 2.940 ;
        RECT 4.630 2.215 6.565 2.710 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.940 1.985 2.280 2.500 ;
        RECT 6.870 2.270 7.740 2.500 ;
        RECT 6.870 1.985 7.130 2.270 ;
        RECT 1.940 1.755 7.130 1.985 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.870 3.400 8.200 3.630 ;
        RECT 0.870 2.890 3.210 3.400 ;
        RECT 0.870 2.270 1.210 2.890 ;
        RECT 7.970 2.500 8.200 3.400 ;
        RECT 7.970 2.270 8.860 2.500 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.550500 ;
    PORT
      LAYER Metal1 ;
        RECT 10.170 3.525 10.735 4.360 ;
        RECT 12.645 3.525 12.875 4.360 ;
        RECT 10.170 3.295 12.875 3.525 ;
        RECT 11.280 1.950 11.835 3.295 ;
        RECT 10.505 1.720 12.975 1.950 ;
        RECT 10.505 0.680 10.735 1.720 ;
        RECT 12.745 0.680 12.975 1.720 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 14.560 5.490 ;
        RECT 0.345 3.755 0.575 4.590 ;
        RECT 9.460 4.275 9.690 4.590 ;
        RECT 11.575 3.755 11.805 4.590 ;
        RECT 13.765 3.755 13.995 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 14.990 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.990 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.020 ;
        RECT 2.485 0.450 2.715 1.020 ;
        RECT 4.725 0.450 4.955 1.020 ;
        RECT 6.965 0.450 7.195 1.020 ;
        RECT 9.205 0.450 9.435 1.020 ;
        RECT 11.625 0.450 11.855 1.490 ;
        RECT 13.865 0.450 14.095 1.490 ;
        RECT 0.000 -0.450 14.560 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 4.720 3.860 9.320 4.090 ;
        RECT 9.090 2.500 9.320 3.860 ;
        RECT 9.090 2.270 11.050 2.500 ;
        RECT 9.090 1.480 9.320 2.270 ;
        RECT 1.365 1.250 9.320 1.480 ;
        RECT 1.365 0.680 1.595 1.250 ;
        RECT 3.605 0.680 3.835 1.250 ;
        RECT 5.845 0.680 6.075 1.250 ;
        RECT 8.085 0.680 8.315 1.250 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or4_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.630 1.210 4.890 2.520 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.696000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.180 0.915 2.710 ;
        RECT 0.150 1.770 0.410 2.180 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 2.180 2.020 2.710 ;
        RECT 1.270 1.770 1.530 2.180 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.310 1.770 6.835 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.495 2.710 19.725 3.690 ;
        RECT 19.190 1.210 19.725 2.710 ;
        RECT 19.445 0.790 19.725 1.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 21.280 5.490 ;
        RECT 1.315 3.440 1.545 4.590 ;
        RECT 5.030 3.965 5.370 4.590 ;
        RECT 7.180 3.995 7.520 4.590 ;
        RECT 12.595 3.440 12.825 4.590 ;
        RECT 17.025 3.595 17.255 4.590 ;
        RECT 20.515 3.880 20.745 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.310 21.710 5.470 ;
        RECT -0.430 2.265 0.430 2.310 ;
        RECT 19.210 2.270 21.710 2.310 ;
        RECT 20.850 2.265 21.710 2.270 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 9.270 2.265 17.710 2.310 ;
        RECT -0.430 -0.430 21.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.450 1.650 1.075 ;
        RECT 5.450 0.450 5.790 0.510 ;
        RECT 7.450 0.450 7.790 0.510 ;
        RECT 12.810 0.450 13.150 0.505 ;
        RECT 17.385 0.450 17.615 0.720 ;
        RECT 20.565 0.450 20.795 1.600 ;
        RECT 0.000 -0.450 21.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.295 3.210 0.525 4.250 ;
        RECT 3.125 3.735 3.355 4.250 ;
        RECT 9.615 3.735 9.845 3.845 ;
        RECT 3.125 3.505 9.845 3.735 ;
        RECT 3.125 3.440 3.355 3.505 ;
        RECT 0.295 2.980 2.775 3.210 ;
        RECT 2.545 1.535 2.775 2.980 ;
        RECT 6.030 3.045 8.355 3.275 ;
        RECT 6.030 2.935 6.260 3.045 ;
        RECT 8.125 1.540 8.355 3.045 ;
        RECT 0.245 1.305 2.775 1.535 ;
        RECT 0.245 0.790 0.475 1.305 ;
        RECT 6.165 1.200 8.355 1.540 ;
        RECT 8.705 2.520 8.935 3.260 ;
        RECT 8.705 2.180 10.285 2.520 ;
        RECT 8.705 1.220 9.075 2.180 ;
        RECT 10.685 1.950 10.915 4.250 ;
        RECT 14.015 2.980 14.375 4.250 ;
        RECT 12.205 2.750 14.375 2.980 ;
        RECT 12.205 2.180 12.435 2.750 ;
        RECT 13.435 1.950 13.665 2.520 ;
        RECT 10.685 1.720 13.665 1.950 ;
        RECT 3.325 0.970 3.555 1.130 ;
        RECT 9.565 0.970 9.795 1.480 ;
        RECT 10.685 1.360 10.915 1.720 ;
        RECT 14.145 1.360 14.375 2.750 ;
        RECT 15.265 3.365 15.495 4.250 ;
        RECT 15.265 3.135 17.930 3.365 ;
        RECT 15.265 1.360 15.495 3.135 ;
        RECT 15.725 1.020 16.065 2.905 ;
        RECT 16.630 1.545 16.970 2.465 ;
        RECT 17.590 2.235 17.930 3.135 ;
        RECT 18.225 2.520 18.455 4.250 ;
        RECT 18.225 2.290 18.955 2.520 ;
        RECT 18.725 1.545 18.955 2.290 ;
        RECT 16.630 1.315 18.955 1.545 ;
        RECT 3.325 0.740 9.795 0.970 ;
        RECT 11.365 0.735 16.065 1.020 ;
        RECT 11.365 0.680 11.595 0.735 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffq_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.400 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.070 2.225 4.835 2.710 ;
        RECT 4.070 1.770 4.330 2.225 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.696000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.225 1.015 2.710 ;
        RECT 0.150 1.770 0.410 2.225 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.135 2.710 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.430 1.770 7.690 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.702050 ;
    PORT
      LAYER Metal1 ;
        RECT 20.790 0.845 21.130 4.250 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 22.400 5.490 ;
        RECT 1.365 3.440 1.595 4.590 ;
        RECT 5.235 3.905 5.465 4.590 ;
        RECT 7.830 3.905 8.170 4.590 ;
        RECT 13.235 3.440 13.465 4.590 ;
        RECT 17.645 3.600 17.875 4.590 ;
        RECT 19.735 3.880 19.965 4.590 ;
        RECT 21.810 3.880 22.040 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 22.830 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 22.830 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.450 1.650 1.075 ;
        RECT 5.505 0.450 5.735 0.620 ;
        RECT 7.565 0.450 7.795 0.620 ;
        RECT 12.870 0.450 13.100 0.620 ;
        RECT 17.745 0.450 17.975 1.590 ;
        RECT 19.685 0.450 19.915 1.600 ;
        RECT 21.925 0.450 22.155 1.165 ;
        RECT 0.000 -0.450 22.400 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 3.210 0.575 4.250 ;
        RECT 3.375 4.020 5.005 4.250 ;
        RECT 3.375 3.440 3.605 4.020 ;
        RECT 4.775 3.675 5.005 4.020 ;
        RECT 10.455 3.675 10.685 3.785 ;
        RECT 4.775 3.445 10.685 3.675 ;
        RECT 0.345 2.980 2.895 3.210 ;
        RECT 2.665 1.540 2.895 2.980 ;
        RECT 6.865 2.985 8.555 3.215 ;
        RECT 6.865 2.875 7.095 2.985 ;
        RECT 0.245 1.310 2.895 1.540 ;
        RECT 6.225 1.540 6.455 1.650 ;
        RECT 8.325 1.540 8.555 2.985 ;
        RECT 6.225 1.310 8.555 1.540 ;
        RECT 8.905 2.565 9.135 3.215 ;
        RECT 8.905 2.225 11.125 2.565 ;
        RECT 8.905 1.310 9.135 2.225 ;
        RECT 11.475 1.995 11.705 4.250 ;
        RECT 14.255 3.025 14.485 4.250 ;
        RECT 12.795 2.795 14.485 3.025 ;
        RECT 12.795 2.225 13.025 2.795 ;
        RECT 13.525 1.995 13.755 2.565 ;
        RECT 11.475 1.765 13.755 1.995 ;
        RECT 11.475 1.650 11.705 1.765 ;
        RECT 0.245 0.790 0.475 1.310 ;
        RECT 3.325 1.080 3.555 1.130 ;
        RECT 9.625 1.080 9.855 1.430 ;
        RECT 10.745 1.310 11.705 1.650 ;
        RECT 14.205 1.310 14.485 2.795 ;
        RECT 15.325 3.370 15.555 4.250 ;
        RECT 15.325 3.140 17.895 3.370 ;
        RECT 15.325 1.310 15.555 3.140 ;
        RECT 15.785 1.080 16.015 2.910 ;
        RECT 17.205 2.050 17.435 2.565 ;
        RECT 17.665 2.510 17.895 3.140 ;
        RECT 18.665 2.565 18.895 4.250 ;
        RECT 17.665 2.280 18.370 2.510 ;
        RECT 18.665 2.225 19.410 2.565 ;
        RECT 18.665 2.050 19.095 2.225 ;
        RECT 17.205 1.820 19.095 2.050 ;
        RECT 3.325 0.850 9.855 1.080 ;
        RECT 11.370 0.850 16.015 1.080 ;
        RECT 3.325 0.790 3.555 0.850 ;
        RECT 11.370 0.685 11.710 0.850 ;
        RECT 14.730 0.685 16.015 0.850 ;
        RECT 18.865 0.790 19.095 1.820 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffq_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 24.640 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.070 2.370 4.330 2.710 ;
        RECT 4.070 2.030 4.835 2.370 ;
        RECT 4.070 1.770 4.330 2.030 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.696000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 1.770 0.415 2.710 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.370 0.970 2.710 ;
        RECT 0.710 2.030 2.035 2.370 ;
        RECT 0.710 1.770 0.970 2.030 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.190 1.770 5.625 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.468150 ;
    PORT
      LAYER Metal1 ;
        RECT 20.705 3.645 20.985 4.250 ;
        RECT 22.805 3.645 23.035 4.250 ;
        RECT 20.705 3.415 23.035 3.645 ;
        RECT 20.705 2.150 20.935 3.415 ;
        RECT 20.705 1.920 22.810 2.150 ;
        RECT 20.705 0.845 20.935 1.920 ;
        RECT 22.550 1.655 22.810 1.920 ;
        RECT 22.550 1.210 23.175 1.655 ;
        RECT 22.945 0.845 23.175 1.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 24.640 5.490 ;
        RECT 1.645 3.440 1.875 4.590 ;
        RECT 5.235 4.135 5.465 4.590 ;
        RECT 5.235 3.905 8.170 4.135 ;
        RECT 13.085 3.440 13.315 4.590 ;
        RECT 17.645 3.550 17.875 4.590 ;
        RECT 19.735 3.875 19.965 4.590 ;
        RECT 21.775 3.875 22.005 4.590 ;
        RECT 23.930 3.875 24.160 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 25.070 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 25.070 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.450 1.650 1.075 ;
        RECT 5.505 0.450 5.735 0.625 ;
        RECT 7.565 0.450 7.795 0.625 ;
        RECT 12.920 0.450 13.150 0.625 ;
        RECT 17.745 0.450 17.975 1.395 ;
        RECT 19.585 0.450 19.815 1.600 ;
        RECT 21.825 0.450 22.055 1.165 ;
        RECT 24.065 0.450 24.295 1.165 ;
        RECT 0.000 -0.450 24.640 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.625 3.210 0.855 4.250 ;
        RECT 3.405 3.675 3.635 4.250 ;
        RECT 10.290 3.675 10.520 3.785 ;
        RECT 3.405 3.445 10.520 3.675 ;
        RECT 3.405 3.440 3.635 3.445 ;
        RECT 0.625 2.980 3.055 3.210 ;
        RECT 2.825 1.535 3.055 2.980 ;
        RECT 6.865 2.875 8.455 3.215 ;
        RECT 8.225 1.655 8.455 2.875 ;
        RECT 0.245 1.305 3.055 1.535 ;
        RECT 6.225 1.315 8.455 1.655 ;
        RECT 8.905 2.370 9.135 3.215 ;
        RECT 8.905 2.030 11.095 2.370 ;
        RECT 8.905 1.315 9.135 2.030 ;
        RECT 11.325 1.800 11.555 4.250 ;
        RECT 14.205 2.830 14.435 4.250 ;
        RECT 12.645 2.600 14.435 2.830 ;
        RECT 12.645 2.030 12.875 2.600 ;
        RECT 13.525 1.800 13.755 2.370 ;
        RECT 11.325 1.655 13.755 1.800 ;
        RECT 10.745 1.570 13.755 1.655 ;
        RECT 0.245 0.790 0.475 1.305 ;
        RECT 3.325 1.085 3.555 1.130 ;
        RECT 9.625 1.085 9.855 1.435 ;
        RECT 10.745 1.315 11.540 1.570 ;
        RECT 14.205 1.315 14.435 2.600 ;
        RECT 15.325 3.320 15.555 4.250 ;
        RECT 15.325 3.090 17.895 3.320 ;
        RECT 15.325 1.315 15.555 3.090 ;
        RECT 15.785 1.085 16.125 2.860 ;
        RECT 17.205 1.855 17.435 2.370 ;
        RECT 17.665 2.315 17.895 3.090 ;
        RECT 18.735 2.370 18.965 4.250 ;
        RECT 17.665 2.085 18.440 2.315 ;
        RECT 18.735 2.030 20.255 2.370 ;
        RECT 18.735 1.855 19.095 2.030 ;
        RECT 17.205 1.625 19.095 1.855 ;
        RECT 3.325 0.855 9.855 1.085 ;
        RECT 11.370 0.855 16.125 1.085 ;
        RECT 3.325 0.790 3.555 0.855 ;
        RECT 11.370 0.690 11.710 0.855 ;
        RECT 14.730 0.690 16.125 0.855 ;
        RECT 18.865 0.790 19.095 1.625 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffq_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffrnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffrnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.960 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 2.330 4.330 2.710 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.696000 ;
    PORT
      LAYER Metal1 ;
        RECT 18.630 1.770 18.890 2.710 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.696000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.330 0.970 2.710 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 2.330 2.090 2.710 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.310 2.330 7.130 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 20.870 0.845 21.330 4.250 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 22.960 5.490 ;
        RECT 1.315 3.440 1.545 4.590 ;
        RECT 5.085 3.440 5.315 4.590 ;
        RECT 7.180 4.030 7.520 4.590 ;
        RECT 12.155 3.910 12.385 4.590 ;
        RECT 13.955 3.440 14.185 4.590 ;
        RECT 18.200 3.910 18.430 4.590 ;
        RECT 20.240 3.440 20.470 4.590 ;
        RECT 22.120 3.440 22.350 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 23.390 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 23.390 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.285 ;
        RECT 5.450 0.450 5.680 0.530 ;
        RECT 7.285 0.450 7.515 1.180 ;
        RECT 13.265 0.450 13.495 1.440 ;
        RECT 18.200 0.450 18.430 1.275 ;
        RECT 22.170 0.450 22.400 1.655 ;
        RECT 0.000 -0.450 22.960 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.295 3.210 0.525 4.250 ;
        RECT 3.325 3.210 3.555 4.250 ;
        RECT 5.545 3.525 9.380 3.755 ;
        RECT 5.545 3.210 5.775 3.525 ;
        RECT 0.295 2.980 2.775 3.210 ;
        RECT 3.325 2.980 5.775 3.210 ;
        RECT 6.160 3.010 7.955 3.240 ;
        RECT 2.545 2.100 2.775 2.980 ;
        RECT 4.605 2.100 4.835 2.635 ;
        RECT 7.725 2.100 7.955 3.010 ;
        RECT 8.305 2.580 8.535 3.295 ;
        RECT 10.115 3.095 10.345 4.250 ;
        RECT 11.135 3.670 11.365 4.250 ;
        RECT 13.175 3.670 13.405 4.250 ;
        RECT 11.135 3.440 13.405 3.670 ;
        RECT 10.115 2.865 14.310 3.095 ;
        RECT 8.305 2.390 9.820 2.580 ;
        RECT 0.245 1.870 4.835 2.100 ;
        RECT 6.165 1.870 7.955 2.100 ;
        RECT 8.405 2.350 9.820 2.390 ;
        RECT 0.245 0.945 0.475 1.870 ;
        RECT 3.325 0.990 3.555 1.285 ;
        RECT 6.165 1.210 6.395 1.870 ;
        RECT 6.625 1.410 8.175 1.640 ;
        RECT 3.325 0.980 6.095 0.990 ;
        RECT 6.625 0.980 6.855 1.410 ;
        RECT 3.325 0.760 6.855 0.980 ;
        RECT 6.025 0.750 6.855 0.760 ;
        RECT 7.945 0.910 8.175 1.410 ;
        RECT 8.405 1.140 8.635 2.350 ;
        RECT 9.125 0.910 9.355 1.275 ;
        RECT 10.115 0.945 10.475 2.865 ;
        RECT 10.825 1.900 11.055 2.635 ;
        RECT 11.765 2.360 11.995 2.635 ;
        RECT 13.970 2.590 14.310 2.865 ;
        RECT 14.975 2.435 15.205 4.250 ;
        RECT 14.665 2.360 15.205 2.435 ;
        RECT 11.765 2.205 15.205 2.360 ;
        RECT 15.995 4.020 17.970 4.250 ;
        RECT 11.765 2.130 14.835 2.205 ;
        RECT 10.825 1.670 14.375 1.900 ;
        RECT 7.945 0.680 9.355 0.910 ;
        RECT 14.145 0.925 14.375 1.670 ;
        RECT 14.605 1.155 14.835 2.130 ;
        RECT 15.065 0.925 15.295 1.955 ;
        RECT 15.995 1.440 16.225 4.020 ;
        RECT 15.670 1.210 16.225 1.440 ;
        RECT 16.600 0.925 16.830 3.150 ;
        RECT 17.080 1.155 17.410 3.780 ;
        RECT 17.740 3.680 17.970 4.020 ;
        RECT 18.660 4.010 19.910 4.240 ;
        RECT 18.660 3.680 18.890 4.010 ;
        RECT 17.740 3.450 18.890 3.680 ;
        RECT 19.220 3.170 19.450 3.780 ;
        RECT 17.760 2.940 19.450 3.170 ;
        RECT 17.760 2.295 17.990 2.940 ;
        RECT 19.220 2.065 19.450 2.940 ;
        RECT 19.680 2.295 19.910 4.010 ;
        RECT 20.400 2.065 20.630 2.635 ;
        RECT 19.220 1.835 20.630 2.065 ;
        RECT 20.240 0.945 20.630 1.835 ;
        RECT 14.145 0.695 16.830 0.925 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffrnq_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffrnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffrnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 2.330 3.995 3.270 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.144000 ;
    PORT
      LAYER Metal1 ;
        RECT 18.070 2.890 18.890 3.270 ;
        RECT 18.610 1.770 18.890 2.890 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.330 1.530 2.735 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.770 1.830 2.150 2.750 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.310 2.330 7.130 2.735 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.674600 ;
    PORT
      LAYER Metal1 ;
        RECT 21.895 0.840 22.250 4.250 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 23.520 5.490 ;
        RECT 1.365 3.440 1.595 4.590 ;
        RECT 5.085 3.440 5.315 4.590 ;
        RECT 7.175 3.940 7.515 4.590 ;
        RECT 12.030 3.440 12.260 4.590 ;
        RECT 13.770 3.440 14.000 4.590 ;
        RECT 18.070 4.480 18.300 4.590 ;
        RECT 20.330 3.440 20.560 4.590 ;
        RECT 22.915 3.440 23.145 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 23.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 23.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.140 ;
        RECT 5.505 0.450 5.735 0.605 ;
        RECT 7.330 0.450 7.560 1.180 ;
        RECT 13.130 0.450 13.360 1.325 ;
        RECT 17.850 0.450 18.080 1.325 ;
        RECT 20.805 0.450 21.035 1.160 ;
        RECT 23.045 0.450 23.275 1.160 ;
        RECT 0.000 -0.450 23.520 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 3.210 0.575 4.250 ;
        RECT 3.125 4.020 4.855 4.250 ;
        RECT 3.125 3.440 3.355 4.020 ;
        RECT 4.625 3.210 4.855 4.020 ;
        RECT 8.970 3.710 9.200 4.250 ;
        RECT 5.545 3.480 9.200 3.710 ;
        RECT 5.545 3.210 5.775 3.480 ;
        RECT 8.970 3.440 9.200 3.480 ;
        RECT 0.345 2.980 2.775 3.210 ;
        RECT 4.625 2.980 5.775 3.210 ;
        RECT 2.545 1.600 2.775 2.980 ;
        RECT 6.155 2.965 7.590 3.195 ;
        RECT 7.360 2.735 7.590 2.965 ;
        RECT 8.250 2.735 8.535 3.250 ;
        RECT 9.990 2.915 10.220 4.250 ;
        RECT 11.010 3.210 11.240 4.250 ;
        RECT 13.050 3.210 13.280 4.250 ;
        RECT 14.790 3.250 15.020 4.250 ;
        RECT 11.010 2.980 13.280 3.210 ;
        RECT 14.250 3.020 15.020 3.250 ;
        RECT 15.810 4.020 20.000 4.250 ;
        RECT 9.990 2.735 10.535 2.915 ;
        RECT 4.650 1.600 4.990 2.735 ;
        RECT 7.360 2.505 7.955 2.735 ;
        RECT 8.250 2.520 9.695 2.735 ;
        RECT 9.990 2.685 13.955 2.735 ;
        RECT 8.450 2.505 9.695 2.520 ;
        RECT 10.310 2.505 13.955 2.685 ;
        RECT 7.360 2.100 7.590 2.505 ;
        RECT 0.245 1.370 4.990 1.600 ;
        RECT 6.210 1.870 7.590 2.100 ;
        RECT 0.245 0.800 0.475 1.370 ;
        RECT 6.210 1.270 6.440 1.870 ;
        RECT 6.670 1.410 8.220 1.640 ;
        RECT 3.270 1.065 3.610 1.085 ;
        RECT 3.270 1.040 6.105 1.065 ;
        RECT 6.670 1.040 6.900 1.410 ;
        RECT 3.270 0.835 6.900 1.040 ;
        RECT 6.000 0.810 6.900 0.835 ;
        RECT 7.990 0.985 8.220 1.410 ;
        RECT 8.450 1.215 8.680 2.505 ;
        RECT 9.190 0.985 9.420 1.325 ;
        RECT 10.310 0.985 10.540 2.505 ;
        RECT 14.250 2.275 14.480 3.020 ;
        RECT 11.535 2.045 14.480 2.275 ;
        RECT 10.835 1.815 11.175 1.960 ;
        RECT 10.835 1.585 14.020 1.815 ;
        RECT 13.790 0.985 14.020 1.585 ;
        RECT 14.250 1.215 14.480 2.045 ;
        RECT 14.790 0.985 15.020 2.790 ;
        RECT 15.810 1.555 16.040 4.020 ;
        RECT 15.390 1.215 16.040 1.555 ;
        RECT 16.270 0.985 16.500 2.790 ;
        RECT 16.730 1.215 17.060 3.780 ;
        RECT 17.410 3.550 19.540 3.780 ;
        RECT 17.410 2.450 17.640 3.550 ;
        RECT 19.310 2.215 19.540 3.550 ;
        RECT 19.770 2.525 20.000 4.020 ;
        RECT 19.310 1.985 20.585 2.215 ;
        RECT 7.990 0.755 9.420 0.985 ;
        RECT 13.790 0.755 16.500 0.985 ;
        RECT 19.990 0.800 20.220 1.985 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffrnq_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffrnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffrnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.320 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 2.330 4.490 2.735 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.144000 ;
    PORT
      LAYER Metal1 ;
        RECT 18.630 1.770 18.890 2.790 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 1.175 2.735 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.530 2.735 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.870 1.770 7.400 2.735 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.642000 ;
    PORT
      LAYER Metal1 ;
        RECT 22.425 1.620 22.655 4.250 ;
        RECT 24.230 1.620 24.895 4.250 ;
        RECT 22.425 1.390 24.895 1.620 ;
        RECT 22.425 0.840 22.655 1.390 ;
        RECT 24.230 1.210 24.895 1.390 ;
        RECT 24.665 0.840 24.895 1.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 26.320 5.490 ;
        RECT 1.510 3.440 1.740 4.590 ;
        RECT 5.525 3.440 5.755 4.590 ;
        RECT 7.640 3.940 7.980 4.590 ;
        RECT 12.825 3.450 13.055 4.590 ;
        RECT 14.585 3.440 14.815 4.590 ;
        RECT 18.885 4.350 19.115 4.590 ;
        RECT 20.925 3.440 21.155 4.590 ;
        RECT 23.495 3.440 23.725 4.590 ;
        RECT 25.645 3.440 25.875 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 26.750 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 26.750 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.585 0.450 1.815 1.080 ;
        RECT 5.945 0.450 6.175 0.645 ;
        RECT 7.965 0.450 8.195 0.620 ;
        RECT 13.945 0.450 14.175 1.380 ;
        RECT 18.445 0.450 18.675 1.380 ;
        RECT 21.305 0.450 21.535 1.160 ;
        RECT 23.545 0.450 23.775 1.160 ;
        RECT 25.785 0.450 26.015 1.160 ;
        RECT 0.000 -0.450 26.320 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.490 3.195 0.720 4.250 ;
        RECT 3.765 3.210 3.995 4.250 ;
        RECT 9.765 3.710 9.995 4.250 ;
        RECT 5.985 3.480 9.995 3.710 ;
        RECT 5.985 3.210 6.215 3.480 ;
        RECT 9.765 3.440 9.995 3.480 ;
        RECT 0.490 2.965 3.215 3.195 ;
        RECT 3.765 2.980 6.215 3.210 ;
        RECT 6.620 2.965 7.860 3.195 ;
        RECT 2.985 2.100 3.215 2.965 ;
        RECT 5.145 2.100 5.375 2.750 ;
        RECT 7.630 2.735 7.860 2.965 ;
        RECT 8.715 2.735 8.945 3.250 ;
        RECT 10.785 2.940 11.015 4.250 ;
        RECT 11.805 3.220 12.035 4.250 ;
        RECT 13.845 3.220 14.075 4.250 ;
        RECT 15.605 3.250 15.835 4.250 ;
        RECT 11.805 2.990 14.075 3.220 ;
        RECT 15.065 3.020 15.835 3.250 ;
        RECT 16.625 4.245 18.450 4.250 ;
        RECT 16.625 4.120 18.680 4.245 ;
        RECT 19.245 4.120 20.595 4.160 ;
        RECT 16.625 4.020 20.595 4.120 ;
        RECT 16.625 3.115 16.855 4.020 ;
        RECT 18.400 3.930 20.595 4.020 ;
        RECT 18.400 3.890 19.375 3.930 ;
        RECT 10.785 2.760 11.370 2.940 ;
        RECT 7.630 2.505 8.420 2.735 ;
        RECT 8.715 2.505 10.490 2.735 ;
        RECT 10.785 2.710 14.770 2.760 ;
        RECT 11.145 2.530 14.770 2.710 ;
        RECT 2.985 1.870 5.375 2.100 ;
        RECT 2.985 1.540 3.215 1.870 ;
        RECT 8.190 1.540 8.420 2.505 ;
        RECT 0.245 1.310 3.215 1.540 ;
        RECT 0.245 1.005 0.475 1.310 ;
        RECT 3.765 1.105 3.995 1.345 ;
        RECT 6.570 1.310 8.420 1.540 ;
        RECT 9.305 1.195 9.535 2.505 ;
        RECT 3.765 1.080 6.465 1.105 ;
        RECT 3.765 0.965 9.080 1.080 ;
        RECT 10.025 0.965 10.255 1.380 ;
        RECT 11.145 1.070 11.375 2.530 ;
        RECT 15.065 2.300 15.295 3.020 ;
        RECT 16.185 2.885 16.855 3.115 ;
        RECT 17.525 3.440 17.875 3.780 ;
        RECT 12.370 2.070 15.295 2.300 ;
        RECT 11.670 1.840 12.010 2.015 ;
        RECT 11.670 1.610 14.835 1.840 ;
        RECT 3.765 0.875 10.255 0.965 ;
        RECT 6.360 0.850 10.255 0.875 ;
        RECT 8.855 0.735 10.255 0.850 ;
        RECT 14.605 1.040 14.835 1.610 ;
        RECT 15.065 1.270 15.295 2.070 ;
        RECT 15.605 1.040 15.835 2.790 ;
        RECT 16.185 1.270 16.415 2.885 ;
        RECT 17.065 2.070 17.295 2.790 ;
        RECT 16.865 1.840 17.295 2.070 ;
        RECT 16.865 1.040 17.095 1.840 ;
        RECT 17.525 1.610 17.755 3.440 ;
        RECT 19.905 3.250 20.135 3.700 ;
        RECT 18.005 3.155 20.135 3.250 ;
        RECT 18.005 3.020 20.115 3.155 ;
        RECT 18.005 2.450 18.235 3.020 ;
        RECT 19.885 2.215 20.115 3.020 ;
        RECT 20.365 2.855 20.595 3.930 ;
        RECT 20.345 2.515 20.595 2.855 ;
        RECT 19.885 1.985 21.085 2.215 ;
        RECT 17.325 1.270 17.755 1.610 ;
        RECT 14.605 0.810 17.095 1.040 ;
        RECT 20.585 0.800 20.815 1.985 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffrnq_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.760 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 2.430 3.210 2.710 ;
        RECT 2.950 2.200 4.075 2.430 ;
        RECT 2.950 1.770 3.210 2.200 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.898000 ;
    PORT
      LAYER Metal1 ;
        RECT 21.430 1.770 21.795 2.710 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.145 0.940 2.710 ;
        RECT 0.150 1.770 0.410 2.145 ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.745 1.770 20.010 2.710 ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.090 2.710 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.310 2.330 7.130 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 24.775 2.560 25.050 4.075 ;
        RECT 24.775 2.330 25.515 2.560 ;
        RECT 25.285 0.845 25.515 2.330 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 25.760 5.490 ;
        RECT 1.340 3.435 1.570 4.590 ;
        RECT 5.110 3.905 5.340 4.590 ;
        RECT 7.030 4.005 7.370 4.590 ;
        RECT 12.125 4.330 12.355 4.590 ;
        RECT 15.245 4.505 15.475 4.590 ;
        RECT 19.275 4.070 19.505 4.590 ;
        RECT 21.480 4.265 21.820 4.590 ;
        RECT 23.575 3.740 23.805 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 26.190 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 26.190 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.335 0.450 1.675 1.080 ;
        RECT 5.530 0.450 5.760 0.535 ;
        RECT 7.385 0.450 7.615 1.135 ;
        RECT 13.425 0.450 13.655 1.425 ;
        RECT 20.970 0.450 21.310 1.080 ;
        RECT 24.165 0.450 24.395 1.600 ;
        RECT 0.000 -0.450 25.760 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.320 3.170 0.550 4.075 ;
        RECT 3.350 3.665 3.580 4.245 ;
        RECT 10.390 4.100 10.730 4.350 ;
        RECT 15.650 4.275 17.210 4.355 ;
        RECT 15.420 4.125 17.210 4.275 ;
        RECT 19.735 4.215 20.695 4.230 ;
        RECT 15.420 4.100 15.825 4.125 ;
        RECT 5.530 3.665 9.075 3.775 ;
        RECT 3.350 3.545 9.075 3.665 ;
        RECT 3.350 3.435 5.730 3.545 ;
        RECT 0.320 2.940 4.960 3.170 ;
        RECT 6.065 2.940 7.755 3.280 ;
        RECT 2.490 1.540 2.720 2.940 ;
        RECT 4.730 2.145 4.960 2.940 ;
        RECT 7.525 2.055 7.755 2.940 ;
        RECT 8.105 2.485 8.335 3.270 ;
        RECT 8.845 2.965 9.075 3.545 ;
        RECT 9.865 3.125 10.095 3.945 ;
        RECT 10.390 3.870 15.825 4.100 ;
        RECT 19.735 4.000 21.255 4.215 ;
        RECT 10.885 3.265 13.555 3.605 ;
        RECT 14.045 3.265 15.175 3.605 ;
        RECT 9.865 2.945 10.570 3.125 ;
        RECT 9.865 2.895 14.715 2.945 ;
        RECT 10.345 2.715 14.715 2.895 ;
        RECT 8.105 2.255 9.515 2.485 ;
        RECT 0.270 1.310 2.720 1.540 ;
        RECT 6.265 1.825 7.755 2.055 ;
        RECT 8.505 2.145 9.515 2.255 ;
        RECT 0.270 0.795 0.500 1.310 ;
        RECT 6.265 1.225 6.495 1.825 ;
        RECT 6.725 1.365 8.275 1.595 ;
        RECT 3.350 0.995 3.580 1.135 ;
        RECT 6.725 0.995 6.955 1.365 ;
        RECT 3.350 0.765 6.955 0.995 ;
        RECT 8.045 0.995 8.275 1.365 ;
        RECT 8.505 1.225 8.735 2.145 ;
        RECT 9.225 0.995 9.455 1.425 ;
        RECT 10.345 1.085 10.575 2.715 ;
        RECT 14.485 2.605 14.715 2.715 ;
        RECT 10.925 1.885 11.155 2.485 ;
        RECT 11.865 2.375 12.095 2.485 ;
        RECT 14.945 2.375 15.175 3.265 ;
        RECT 11.865 2.145 16.135 2.375 ;
        RECT 10.925 1.655 15.675 1.885 ;
        RECT 8.045 0.765 9.455 0.995 ;
        RECT 15.445 0.910 15.675 1.655 ;
        RECT 15.905 1.545 16.135 2.145 ;
        RECT 16.485 1.545 16.715 3.895 ;
        RECT 17.505 3.840 17.735 3.950 ;
        RECT 19.735 3.840 19.965 4.000 ;
        RECT 20.610 3.990 21.255 4.000 ;
        RECT 20.610 3.985 23.245 3.990 ;
        RECT 17.505 3.610 19.965 3.840 ;
        RECT 17.505 1.655 17.735 3.610 ;
        RECT 18.525 2.945 18.755 3.310 ;
        RECT 15.905 1.315 16.715 1.545 ;
        RECT 17.025 1.315 17.735 1.655 ;
        RECT 18.145 2.715 19.295 2.945 ;
        RECT 18.145 1.315 18.375 2.715 ;
        RECT 18.605 0.910 18.835 2.485 ;
        RECT 15.445 0.680 18.835 0.910 ;
        RECT 19.065 1.540 19.295 2.715 ;
        RECT 20.295 1.540 20.525 3.770 ;
        RECT 21.025 3.760 23.245 3.985 ;
        RECT 19.065 1.310 20.525 1.540 ;
        RECT 20.820 1.540 21.160 2.430 ;
        RECT 22.555 1.540 22.785 3.530 ;
        RECT 23.015 2.145 23.245 3.760 ;
        RECT 24.195 2.060 24.425 2.485 ;
        RECT 23.460 1.830 24.425 2.060 ;
        RECT 23.460 1.540 23.690 1.830 ;
        RECT 20.820 1.310 23.690 1.540 ;
        RECT 19.065 0.795 19.295 1.310 ;
        RECT 23.445 0.795 23.690 1.310 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.880 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 1.770 4.330 2.290 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.123000 ;
    PORT
      LAYER Metal1 ;
        RECT 21.430 2.355 21.690 2.710 ;
        RECT 21.430 2.015 21.935 2.355 ;
        RECT 21.430 1.770 21.690 2.015 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 1.770 0.970 2.300 ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.750 1.770 20.040 2.710 ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 1.770 2.090 2.345 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.310 2.330 7.130 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 25.145 2.710 25.375 4.080 ;
        RECT 25.145 0.790 25.610 2.710 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 26.880 5.490 ;
        RECT 1.415 3.270 1.645 4.590 ;
        RECT 5.085 3.440 5.315 4.590 ;
        RECT 7.190 4.125 7.530 4.590 ;
        RECT 12.210 4.565 12.550 4.590 ;
        RECT 15.350 4.565 15.690 4.590 ;
        RECT 19.395 3.910 19.625 4.590 ;
        RECT 21.665 4.300 21.895 4.590 ;
        RECT 23.725 3.270 23.955 4.590 ;
        RECT 26.165 3.270 26.395 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.320 27.310 5.470 ;
        RECT -0.430 2.265 0.430 2.320 ;
        RECT 21.385 2.265 27.310 2.320 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 9.180 2.280 18.695 2.320 ;
        RECT 8.440 2.265 18.695 2.280 ;
        RECT -0.430 -0.430 27.310 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.450 1.650 1.075 ;
        RECT 5.505 0.450 5.735 1.080 ;
        RECT 7.545 0.450 7.775 1.080 ;
        RECT 13.545 0.450 13.775 1.480 ;
        RECT 20.970 0.450 21.310 1.080 ;
        RECT 24.165 0.450 24.395 1.600 ;
        RECT 26.405 0.450 26.635 1.600 ;
        RECT 0.000 -0.450 26.880 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 10.530 4.105 17.310 4.335 ;
        RECT 0.395 2.805 0.625 4.080 ;
        RECT 3.325 3.210 3.555 4.080 ;
        RECT 5.545 3.665 9.215 3.895 ;
        RECT 5.545 3.210 5.775 3.665 ;
        RECT 3.325 2.980 5.775 3.210 ;
        RECT 6.225 3.095 7.590 3.435 ;
        RECT 0.395 2.750 2.745 2.805 ;
        RECT 0.395 2.575 4.835 2.750 ;
        RECT 2.595 2.520 4.835 2.575 ;
        RECT 2.595 1.540 2.825 2.520 ;
        RECT 4.605 2.015 4.835 2.520 ;
        RECT 7.360 2.110 7.590 3.095 ;
        RECT 8.265 2.565 8.495 3.435 ;
        RECT 8.985 3.085 9.215 3.665 ;
        RECT 10.005 2.970 10.235 3.930 ;
        RECT 14.165 3.645 16.815 3.875 ;
        RECT 19.855 3.840 23.375 4.070 ;
        RECT 11.025 3.270 13.675 3.610 ;
        RECT 14.165 3.535 16.135 3.645 ;
        RECT 14.305 2.970 14.535 3.080 ;
        RECT 10.005 2.740 14.535 2.970 ;
        RECT 8.265 2.335 9.655 2.565 ;
        RECT 8.665 2.225 9.655 2.335 ;
        RECT 7.360 2.000 8.215 2.110 ;
        RECT 6.425 1.770 8.215 2.000 ;
        RECT 0.245 1.310 2.825 1.540 ;
        RECT 3.325 1.310 6.195 1.540 ;
        RECT 0.245 0.790 0.475 1.310 ;
        RECT 3.325 0.790 3.555 1.310 ;
        RECT 5.965 0.940 6.195 1.310 ;
        RECT 6.425 1.170 6.655 1.770 ;
        RECT 6.885 1.310 8.435 1.540 ;
        RECT 6.885 0.940 7.115 1.310 ;
        RECT 5.965 0.710 7.115 0.940 ;
        RECT 8.205 0.940 8.435 1.310 ;
        RECT 8.665 1.170 8.895 2.225 ;
        RECT 9.465 0.940 9.695 1.480 ;
        RECT 10.585 1.370 10.815 2.740 ;
        RECT 15.905 2.510 16.135 3.535 ;
        RECT 16.585 3.065 16.815 3.645 ;
        RECT 17.605 3.680 19.215 3.765 ;
        RECT 19.855 3.680 20.085 3.840 ;
        RECT 17.605 3.535 20.085 3.680 ;
        RECT 17.605 2.970 17.835 3.535 ;
        RECT 19.035 3.450 20.085 3.535 ;
        RECT 11.165 1.940 11.395 2.355 ;
        RECT 12.005 2.170 16.135 2.510 ;
        RECT 11.165 1.710 15.675 1.940 ;
        RECT 8.205 0.710 9.695 0.940 ;
        RECT 15.445 1.020 15.675 1.710 ;
        RECT 15.905 1.370 16.135 2.170 ;
        RECT 17.025 2.740 17.835 2.970 ;
        RECT 18.625 2.815 18.855 3.305 ;
        RECT 20.400 3.270 20.645 3.610 ;
        RECT 17.025 1.370 17.255 2.740 ;
        RECT 18.145 2.585 19.295 2.815 ;
        RECT 18.145 1.370 18.375 2.585 ;
        RECT 18.605 1.020 18.835 2.355 ;
        RECT 19.065 1.540 19.295 2.585 ;
        RECT 20.400 1.540 20.630 3.270 ;
        RECT 19.065 1.310 20.630 1.540 ;
        RECT 20.860 1.540 21.200 2.300 ;
        RECT 22.685 1.540 22.915 3.610 ;
        RECT 23.145 2.415 23.375 3.840 ;
        RECT 24.605 2.195 24.835 2.355 ;
        RECT 23.445 1.965 24.835 2.195 ;
        RECT 23.445 1.540 23.675 1.965 ;
        RECT 20.860 1.310 23.675 1.540 ;
        RECT 19.065 1.025 19.295 1.310 ;
        RECT 15.445 0.680 18.835 1.020 ;
        RECT 23.445 0.845 23.675 1.310 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 29.120 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 1.770 3.770 2.710 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.123000 ;
    PORT
      LAYER Metal1 ;
        RECT 21.430 2.215 21.690 3.270 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.270 0.970 2.710 ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.130 2.950 20.010 3.270 ;
        RECT 19.655 2.740 20.010 2.950 ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 2.270 2.090 2.710 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 2.890 6.570 3.270 ;
        RECT 6.280 2.530 6.570 2.890 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 24.850 3.120 25.080 4.250 ;
        RECT 26.470 3.440 27.120 4.250 ;
        RECT 26.470 3.120 26.730 3.440 ;
        RECT 24.850 2.890 27.720 3.120 ;
        RECT 25.250 0.845 25.480 2.890 ;
        RECT 27.490 0.845 27.720 2.890 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 29.120 5.490 ;
        RECT 1.265 3.440 1.495 4.590 ;
        RECT 4.950 4.560 5.290 4.590 ;
        RECT 6.885 4.560 7.225 4.590 ;
        RECT 12.120 4.510 12.350 4.590 ;
        RECT 15.320 4.510 15.550 4.590 ;
        RECT 19.390 3.985 19.620 4.590 ;
        RECT 21.595 4.375 21.935 4.590 ;
        RECT 23.710 3.440 23.940 4.590 ;
        RECT 25.870 3.440 26.100 4.590 ;
        RECT 27.910 3.440 28.140 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 29.550 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 29.550 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.535 ;
        RECT 5.445 0.450 5.675 0.530 ;
        RECT 7.460 0.450 7.690 1.380 ;
        RECT 13.460 0.450 13.690 1.535 ;
        RECT 20.990 0.450 21.220 1.255 ;
        RECT 24.130 0.450 24.360 1.525 ;
        RECT 26.370 0.450 26.600 1.650 ;
        RECT 28.610 0.450 28.840 1.650 ;
        RECT 0.000 -0.450 29.120 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.170 0.475 4.250 ;
        RECT 3.025 4.100 9.130 4.330 ;
        RECT 3.025 3.440 3.255 4.100 ;
        RECT 5.700 3.500 7.830 3.840 ;
        RECT 0.245 2.940 4.835 3.170 ;
        RECT 2.445 2.040 2.675 2.940 ;
        RECT 4.605 2.215 4.835 2.940 ;
        RECT 7.600 2.300 7.830 3.500 ;
        RECT 8.180 2.555 8.410 3.870 ;
        RECT 8.900 3.065 9.130 4.100 ;
        RECT 10.445 4.050 17.355 4.280 ;
        RECT 19.850 3.915 23.360 4.145 ;
        RECT 9.920 3.215 10.150 3.875 ;
        RECT 10.940 3.440 13.590 3.780 ;
        RECT 14.080 3.550 16.860 3.780 ;
        RECT 19.850 3.755 20.080 3.915 ;
        RECT 14.080 3.440 14.310 3.550 ;
        RECT 15.640 3.440 16.860 3.550 ;
        RECT 17.650 3.525 20.080 3.755 ;
        RECT 9.920 3.210 10.550 3.215 ;
        RECT 14.520 3.210 14.750 3.320 ;
        RECT 9.920 2.985 14.750 3.210 ;
        RECT 10.500 2.980 14.750 2.985 ;
        RECT 8.180 2.325 9.570 2.555 ;
        RECT 0.245 1.810 2.675 2.040 ;
        RECT 6.340 2.070 7.830 2.300 ;
        RECT 8.580 2.215 9.570 2.325 ;
        RECT 0.245 1.195 0.475 1.810 ;
        RECT 3.325 0.990 3.555 1.535 ;
        RECT 6.340 1.220 6.570 2.070 ;
        RECT 6.800 1.610 8.350 1.840 ;
        RECT 6.800 0.990 7.030 1.610 ;
        RECT 3.325 0.760 7.030 0.990 ;
        RECT 8.120 0.990 8.350 1.610 ;
        RECT 8.580 1.220 8.810 2.215 ;
        RECT 9.380 0.990 9.610 1.535 ;
        RECT 10.500 1.195 10.730 2.980 ;
        RECT 15.640 2.565 15.870 3.440 ;
        RECT 17.650 3.175 17.880 3.525 ;
        RECT 11.920 2.225 15.870 2.565 ;
        RECT 11.080 1.995 11.310 2.115 ;
        RECT 11.080 1.765 15.410 1.995 ;
        RECT 8.120 0.760 9.610 0.990 ;
        RECT 15.180 0.910 15.410 1.765 ;
        RECT 15.640 1.195 15.870 2.225 ;
        RECT 16.760 2.945 17.880 3.175 ;
        RECT 16.760 1.195 16.990 2.945 ;
        RECT 18.670 2.680 18.900 3.295 ;
        RECT 17.880 2.510 19.255 2.680 ;
        RECT 20.410 2.510 20.640 3.685 ;
        RECT 17.880 2.450 20.640 2.510 ;
        RECT 17.880 1.195 18.110 2.450 ;
        RECT 19.030 2.280 20.640 2.450 ;
        RECT 18.340 0.910 18.680 2.220 ;
        RECT 19.030 1.145 19.260 2.280 ;
        RECT 20.795 1.985 21.135 2.110 ;
        RECT 22.670 1.985 22.900 3.685 ;
        RECT 23.130 2.215 23.360 3.915 ;
        RECT 24.570 1.985 24.800 2.555 ;
        RECT 20.795 1.755 24.800 1.985 ;
        RECT 15.180 0.680 18.680 0.910 ;
        RECT 23.410 0.845 23.640 1.755 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffsnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 24.640 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 1.770 3.995 2.710 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.275 0.970 2.710 ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 18.630 1.770 19.425 2.710 ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 2.275 2.090 2.710 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.310 2.275 7.130 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 23.670 0.845 24.285 4.060 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 24.640 5.490 ;
        RECT 1.315 3.400 1.545 4.590 ;
        RECT 5.145 3.250 5.375 4.590 ;
        RECT 7.450 3.970 7.790 4.590 ;
        RECT 12.595 3.835 12.825 4.590 ;
        RECT 14.955 3.090 15.185 4.590 ;
        RECT 18.955 3.400 19.185 4.590 ;
        RECT 21.195 4.310 21.425 4.590 ;
        RECT 22.985 3.250 23.215 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 25.070 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 25.070 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.450 ;
        RECT 5.455 0.450 5.685 0.630 ;
        RECT 7.555 0.450 7.785 1.140 ;
        RECT 12.640 0.450 12.980 0.625 ;
        RECT 20.875 0.450 21.105 0.610 ;
        RECT 22.935 0.450 23.165 1.165 ;
        RECT 0.000 -0.450 24.640 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.295 3.170 0.525 4.060 ;
        RECT 3.325 3.630 3.555 4.210 ;
        RECT 3.325 3.400 4.915 3.630 ;
        RECT 0.295 2.940 4.455 3.170 ;
        RECT 2.545 2.045 2.775 2.940 ;
        RECT 0.245 1.815 2.775 2.045 ;
        RECT 4.225 2.070 4.455 2.940 ;
        RECT 4.685 3.020 4.915 3.400 ;
        RECT 5.605 3.510 9.675 3.740 ;
        RECT 5.605 3.020 5.835 3.510 ;
        RECT 4.685 2.790 5.835 3.020 ;
        RECT 6.485 2.940 7.675 3.280 ;
        RECT 7.445 2.505 7.675 2.940 ;
        RECT 8.575 2.505 8.805 3.235 ;
        RECT 9.445 2.930 9.675 3.510 ;
        RECT 7.445 2.275 8.280 2.505 ;
        RECT 8.575 2.275 10.170 2.505 ;
        RECT 10.515 2.285 10.745 3.730 ;
        RECT 11.095 3.605 11.325 4.360 ;
        RECT 15.735 4.020 16.865 4.360 ;
        RECT 13.025 3.605 14.725 3.720 ;
        RECT 11.095 3.490 14.725 3.605 ;
        RECT 11.095 3.375 13.225 3.490 ;
        RECT 13.935 2.745 14.165 3.260 ;
        RECT 11.880 2.515 14.165 2.745 ;
        RECT 14.495 2.860 14.725 3.490 ;
        RECT 15.735 2.860 15.965 4.020 ;
        RECT 14.495 2.630 15.965 2.860 ;
        RECT 0.245 1.110 0.475 1.815 ;
        RECT 4.225 1.730 4.835 2.070 ;
        RECT 7.445 2.060 7.675 2.275 ;
        RECT 7.215 2.045 7.675 2.060 ;
        RECT 6.435 1.830 7.675 2.045 ;
        RECT 6.435 1.815 7.300 1.830 ;
        RECT 3.325 1.090 3.555 1.450 ;
        RECT 6.435 1.140 6.665 1.815 ;
        RECT 7.385 1.585 8.245 1.600 ;
        RECT 6.895 1.370 8.245 1.585 ;
        RECT 6.895 1.355 7.470 1.370 ;
        RECT 3.325 0.910 6.210 1.090 ;
        RECT 6.895 0.910 7.125 1.355 ;
        RECT 3.325 0.860 7.125 0.910 ;
        RECT 5.985 0.680 7.125 0.860 ;
        RECT 8.015 0.910 8.245 1.370 ;
        RECT 8.575 1.140 8.905 2.275 ;
        RECT 10.515 2.055 13.640 2.285 ;
        RECT 9.395 0.910 9.625 1.135 ;
        RECT 10.515 1.025 10.745 2.055 ;
        RECT 11.195 1.085 11.425 1.825 ;
        RECT 13.935 1.545 14.165 2.515 ;
        RECT 16.195 1.910 16.425 3.730 ;
        RECT 17.215 1.940 17.445 3.900 ;
        RECT 15.055 1.680 16.425 1.910 ;
        RECT 16.835 1.710 17.445 1.940 ;
        RECT 18.170 3.170 18.465 3.900 ;
        RECT 19.975 3.170 20.205 3.950 ;
        RECT 18.170 2.940 20.205 3.170 ;
        RECT 22.215 3.020 22.445 4.100 ;
        RECT 15.055 1.545 15.285 1.680 ;
        RECT 13.935 1.315 15.285 1.545 ;
        RECT 8.015 0.680 9.625 0.910 ;
        RECT 11.195 0.855 15.780 1.085 ;
        RECT 15.440 0.680 15.780 0.855 ;
        RECT 16.175 0.910 16.405 1.450 ;
        RECT 16.835 0.910 17.065 1.710 ;
        RECT 18.170 1.480 18.400 2.940 ;
        RECT 20.555 2.790 22.445 3.020 ;
        RECT 20.555 2.220 20.785 2.790 ;
        RECT 22.215 2.560 22.445 2.790 ;
        RECT 17.295 1.140 18.985 1.480 ;
        RECT 21.635 1.070 21.865 2.560 ;
        RECT 22.215 2.220 23.440 2.560 ;
        RECT 22.215 1.110 22.445 2.220 ;
        RECT 19.205 0.910 21.865 1.070 ;
        RECT 16.175 0.840 21.865 0.910 ;
        RECT 16.175 0.680 19.425 0.840 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffsnq_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffsnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.200 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 1.770 4.070 2.710 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.320 1.530 2.710 ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 18.630 2.265 19.110 2.605 ;
        RECT 18.630 1.210 18.890 2.265 ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 2.320 2.650 2.710 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.865 2.320 7.690 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 23.605 0.845 23.930 4.050 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 25.200 5.490 ;
        RECT 1.440 3.400 1.670 4.590 ;
        RECT 5.160 3.760 5.390 4.590 ;
        RECT 7.360 3.860 7.590 4.590 ;
        RECT 12.280 3.560 12.510 4.590 ;
        RECT 14.540 3.560 14.770 4.590 ;
        RECT 18.440 3.295 18.670 4.590 ;
        RECT 20.480 3.240 20.710 4.590 ;
        RECT 22.585 3.240 22.815 4.590 ;
        RECT 24.625 3.240 24.855 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 25.630 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 25.630 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.440 0.450 1.670 1.480 ;
        RECT 5.545 0.450 5.775 0.575 ;
        RECT 7.360 0.450 7.590 1.170 ;
        RECT 12.280 0.450 12.510 1.220 ;
        RECT 20.380 0.450 20.610 1.480 ;
        RECT 22.485 0.450 22.715 1.165 ;
        RECT 24.725 0.450 24.955 1.165 ;
        RECT 0.000 -0.450 25.200 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.420 3.170 0.650 4.050 ;
        RECT 3.400 3.630 3.630 4.210 ;
        RECT 7.820 3.915 9.480 4.145 ;
        RECT 5.605 3.630 7.220 3.675 ;
        RECT 7.820 3.630 8.050 3.915 ;
        RECT 3.400 3.530 4.970 3.630 ;
        RECT 5.605 3.530 8.050 3.630 ;
        RECT 3.400 3.445 8.050 3.530 ;
        RECT 3.400 3.400 5.820 3.445 ;
        RECT 7.080 3.400 8.050 3.445 ;
        RECT 4.780 3.300 5.820 3.400 ;
        RECT 6.340 3.170 6.570 3.215 ;
        RECT 0.420 3.070 4.590 3.170 ;
        RECT 0.420 2.940 4.910 3.070 ;
        RECT 2.880 2.090 3.110 2.940 ;
        RECT 4.400 2.840 4.910 2.940 ;
        RECT 6.340 2.940 8.150 3.170 ;
        RECT 6.340 2.875 6.570 2.940 ;
        RECT 4.680 2.265 4.910 2.840 ;
        RECT 7.920 2.090 8.150 2.940 ;
        RECT 0.320 1.860 3.110 2.090 ;
        RECT 6.240 1.860 8.150 2.090 ;
        RECT 8.380 2.550 8.610 3.685 ;
        RECT 9.250 3.090 9.480 3.915 ;
        RECT 8.380 2.320 9.975 2.550 ;
        RECT 0.320 1.140 0.550 1.860 ;
        RECT 3.400 1.035 3.630 1.480 ;
        RECT 6.240 1.260 6.470 1.860 ;
        RECT 6.700 1.400 8.050 1.630 ;
        RECT 3.400 1.030 6.190 1.035 ;
        RECT 6.700 1.030 6.930 1.400 ;
        RECT 3.400 0.805 6.930 1.030 ;
        RECT 6.140 0.800 6.930 0.805 ;
        RECT 7.820 0.910 8.050 1.400 ;
        RECT 8.380 1.140 8.710 2.320 ;
        RECT 10.320 2.315 10.550 3.730 ;
        RECT 10.900 3.330 11.130 4.360 ;
        RECT 12.740 3.960 14.310 4.190 ;
        RECT 12.740 3.330 12.970 3.960 ;
        RECT 10.900 3.100 12.970 3.330 ;
        RECT 13.520 2.745 13.750 3.730 ;
        RECT 14.080 3.330 14.310 3.960 ;
        RECT 15.200 3.975 16.330 4.315 ;
        RECT 15.200 3.330 15.430 3.975 ;
        RECT 14.080 3.100 15.430 3.330 ;
        RECT 15.660 2.745 15.890 3.685 ;
        RECT 11.785 2.515 15.890 2.745 ;
        RECT 10.320 2.285 11.670 2.315 ;
        RECT 10.320 2.085 13.225 2.285 ;
        RECT 9.200 0.910 9.430 1.220 ;
        RECT 10.320 1.110 10.550 2.085 ;
        RECT 11.555 2.055 13.225 2.085 ;
        RECT 10.845 1.825 11.185 1.855 ;
        RECT 10.845 1.595 12.970 1.825 ;
        RECT 7.820 0.680 9.430 0.910 ;
        RECT 12.740 0.910 12.970 1.595 ;
        RECT 14.540 1.140 14.770 2.515 ;
        RECT 16.680 2.115 16.910 3.845 ;
        RECT 17.720 3.065 17.950 3.845 ;
        RECT 19.460 3.065 19.690 4.050 ;
        RECT 17.720 2.835 19.690 3.065 ;
        RECT 21.680 3.010 21.910 4.050 ;
        RECT 16.320 1.885 16.910 2.115 ;
        RECT 16.320 1.480 16.550 1.885 ;
        RECT 18.170 1.655 18.400 2.835 ;
        RECT 20.040 2.780 23.255 3.010 ;
        RECT 20.040 2.265 20.270 2.780 ;
        RECT 20.500 2.320 21.385 2.550 ;
        RECT 20.500 1.940 20.730 2.320 ;
        RECT 15.660 1.140 16.550 1.480 ;
        RECT 16.780 1.315 18.400 1.655 ;
        RECT 19.120 1.710 20.730 1.940 ;
        RECT 16.320 0.980 16.550 1.140 ;
        RECT 19.120 0.980 19.350 1.710 ;
        RECT 12.740 0.680 15.265 0.910 ;
        RECT 16.320 0.750 19.350 0.980 ;
        RECT 21.680 0.845 21.910 2.780 ;
        RECT 23.025 2.265 23.255 2.780 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffsnq_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffsnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.440 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 1.770 4.330 2.215 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 1.770 0.970 2.215 ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 18.070 1.770 18.890 2.215 ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 1.770 2.090 2.215 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 2.330 6.910 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.559650 ;
    PORT
      LAYER Metal1 ;
        RECT 23.590 3.110 23.870 3.690 ;
        RECT 25.690 3.110 25.920 3.690 ;
        RECT 23.590 2.880 25.920 3.110 ;
        RECT 23.590 1.655 23.930 2.880 ;
        RECT 23.590 1.210 26.060 1.655 ;
        RECT 23.590 0.845 23.820 1.210 ;
        RECT 25.830 0.845 26.060 1.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 27.440 5.490 ;
        RECT 1.315 3.230 1.545 4.590 ;
        RECT 5.085 3.400 5.315 4.590 ;
        RECT 7.200 4.125 7.540 4.590 ;
        RECT 12.045 4.510 12.275 4.590 ;
        RECT 14.305 4.070 14.535 4.590 ;
        RECT 18.305 3.075 18.535 4.590 ;
        RECT 20.565 3.880 20.795 4.590 ;
        RECT 22.605 3.880 22.835 4.590 ;
        RECT 24.660 3.880 24.890 4.590 ;
        RECT 26.850 3.880 27.080 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 27.870 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 27.870 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.450 1.650 1.075 ;
        RECT 5.505 0.450 5.735 0.530 ;
        RECT 7.305 0.450 7.535 1.180 ;
        RECT 12.225 0.450 12.455 1.120 ;
        RECT 20.230 0.450 20.460 1.265 ;
        RECT 22.470 0.450 22.700 1.655 ;
        RECT 24.710 0.450 24.940 0.980 ;
        RECT 26.950 0.450 27.180 1.655 ;
        RECT 0.000 -0.450 27.440 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 10.590 4.050 13.975 4.280 ;
        RECT 0.295 2.685 0.525 4.040 ;
        RECT 3.325 3.170 3.555 4.040 ;
        RECT 5.545 3.665 9.275 3.895 ;
        RECT 5.545 3.170 5.775 3.665 ;
        RECT 3.325 2.940 5.775 3.170 ;
        RECT 6.235 3.095 7.370 3.435 ;
        RECT 8.275 3.095 8.655 3.435 ;
        RECT 0.295 2.455 4.835 2.685 ;
        RECT 2.545 1.540 2.775 2.455 ;
        RECT 4.605 1.930 4.835 2.455 ;
        RECT 7.140 2.215 7.370 3.095 ;
        RECT 8.425 2.215 8.655 3.095 ;
        RECT 9.045 3.065 9.275 3.665 ;
        RECT 10.065 2.215 10.295 3.875 ;
        RECT 13.745 3.840 13.975 4.050 ;
        RECT 16.005 3.840 16.235 4.360 ;
        RECT 13.285 2.675 13.515 3.770 ;
        RECT 13.745 3.610 16.235 3.840 ;
        RECT 13.745 3.095 13.975 3.610 ;
        RECT 15.545 2.675 15.775 3.380 ;
        RECT 16.005 3.095 16.235 3.610 ;
        RECT 11.330 2.445 15.775 2.675 ;
        RECT 7.140 2.100 7.980 2.215 ;
        RECT 0.245 1.310 2.775 1.540 ;
        RECT 6.185 1.870 7.980 2.100 ;
        RECT 8.425 1.985 9.720 2.215 ;
        RECT 10.065 1.985 13.170 2.215 ;
        RECT 0.245 0.925 0.475 1.310 ;
        RECT 6.185 1.270 6.415 1.870 ;
        RECT 6.645 1.410 8.195 1.640 ;
        RECT 3.325 0.990 3.555 1.130 ;
        RECT 6.645 0.990 6.875 1.410 ;
        RECT 3.325 0.760 6.875 0.990 ;
        RECT 7.965 0.990 8.195 1.410 ;
        RECT 8.425 1.220 8.655 1.985 ;
        RECT 9.145 0.990 9.375 1.120 ;
        RECT 7.965 0.760 9.375 0.990 ;
        RECT 10.065 0.925 10.495 1.985 ;
        RECT 10.790 1.525 12.915 1.755 ;
        RECT 12.685 0.910 12.915 1.525 ;
        RECT 14.405 1.315 14.635 2.445 ;
        RECT 16.565 1.960 16.795 3.900 ;
        RECT 16.185 1.730 16.795 1.960 ;
        RECT 17.585 2.845 17.815 3.900 ;
        RECT 19.325 2.845 19.555 3.715 ;
        RECT 17.585 2.615 19.555 2.845 ;
        RECT 21.585 2.785 21.815 3.690 ;
        RECT 19.905 2.760 21.815 2.785 ;
        RECT 16.185 1.425 16.415 1.730 ;
        RECT 17.585 1.500 17.815 2.615 ;
        RECT 19.905 2.445 23.275 2.760 ;
        RECT 21.350 2.420 23.275 2.445 ;
        RECT 19.120 1.985 21.055 2.215 ;
        RECT 15.525 1.085 16.415 1.425 ;
        RECT 16.645 1.160 18.320 1.500 ;
        RECT 16.185 0.930 16.415 1.085 ;
        RECT 19.120 0.930 19.350 1.985 ;
        RECT 12.685 0.680 15.130 0.910 ;
        RECT 16.185 0.700 19.350 0.930 ;
        RECT 21.350 0.845 21.580 2.420 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffsnq_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__tieh
  CLASS core TIEHIGH ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__tieh ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.240 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 2.890 1.530 3.700 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 2.240 5.490 ;
        RECT 0.250 2.945 0.480 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 2.670 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 2.670 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 0.450 0.480 1.355 ;
        RECT 0.000 -0.450 2.240 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.875 1.830 1.600 2.060 ;
        RECT 1.370 1.315 1.600 1.830 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__tieh

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__tiel
  CLASS core TIELOW ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__tiel ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.240 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.290400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.215 1.210 1.595 1.590 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 2.240 5.490 ;
        RECT 0.345 2.945 0.575 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 2.670 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 2.670 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.355 ;
        RECT 0.000 -0.450 2.240 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 2.700 1.595 3.685 ;
        RECT 0.870 2.470 1.595 2.700 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__tiel

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__xnor2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xnor2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.720 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.560500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.885 2.580 3.770 2.810 ;
        RECT 1.885 2.065 2.115 2.580 ;
        RECT 3.510 2.350 3.770 2.580 ;
        RECT 3.510 2.120 4.400 2.350 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.560500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.205 3.040 4.890 3.270 ;
        RECT 1.205 2.350 1.435 3.040 ;
        RECT 4.430 2.890 4.890 3.040 ;
        RECT 0.810 2.120 1.435 2.350 ;
        RECT 4.660 2.350 4.890 2.890 ;
        RECT 4.660 2.120 5.470 2.350 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.821000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.675 3.730 3.905 4.310 ;
        RECT 3.675 3.500 5.535 3.730 ;
        RECT 5.305 2.810 5.535 3.500 ;
        RECT 5.305 2.580 6.010 2.810 ;
        RECT 5.750 1.370 6.010 2.580 ;
        RECT 4.690 1.140 6.010 1.370 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 6.720 5.490 ;
        RECT 0.285 3.500 0.515 4.590 ;
        RECT 2.325 3.500 2.555 4.590 ;
        RECT 5.765 3.500 5.995 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 7.150 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.150 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.325 0.450 2.555 1.355 ;
        RECT 0.000 -0.450 6.720 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.305 3.730 1.535 4.310 ;
        RECT 0.745 3.500 1.535 3.730 ;
        RECT 0.745 2.810 0.975 3.500 ;
        RECT 0.285 2.580 0.975 2.810 ;
        RECT 0.285 1.835 0.515 2.580 ;
        RECT 2.345 2.120 3.280 2.350 ;
        RECT 2.345 1.835 2.575 2.120 ;
        RECT 0.285 1.605 2.575 1.835 ;
        RECT 0.285 1.015 0.515 1.605 ;
        RECT 3.625 0.910 3.855 1.655 ;
        RECT 3.625 0.680 6.150 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xnor2_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__xnor2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xnor2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.560500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.995 2.515 4.455 2.745 ;
        RECT 1.995 2.000 2.225 2.515 ;
        RECT 4.070 1.210 4.455 2.515 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.560500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.535 2.975 5.475 3.205 ;
        RECT 1.535 2.285 1.765 2.975 ;
        RECT 0.870 2.055 1.765 2.285 ;
        RECT 5.190 2.135 5.475 2.975 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.821000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.665 1.590 7.895 3.775 ;
        RECT 7.430 1.210 7.895 1.590 ;
        RECT 7.665 0.680 7.895 1.210 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 9.520 5.490 ;
        RECT 2.435 3.435 2.665 4.590 ;
        RECT 6.545 3.875 6.775 4.590 ;
        RECT 8.685 2.965 8.915 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 9.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 0.965 ;
        RECT 2.485 0.450 2.715 0.965 ;
        RECT 5.825 0.450 6.055 1.310 ;
        RECT 6.545 0.450 6.775 1.310 ;
        RECT 8.785 0.450 9.015 1.435 ;
        RECT 0.000 -0.450 9.520 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.785 4.015 6.110 4.245 ;
        RECT 0.345 1.770 0.575 3.775 ;
        RECT 3.785 3.435 4.015 4.015 ;
        RECT 4.750 3.435 5.935 3.665 ;
        RECT 2.455 2.055 3.490 2.285 ;
        RECT 5.705 2.115 5.935 3.435 ;
        RECT 2.455 1.770 2.685 2.055 ;
        RECT 5.705 1.905 7.215 2.115 ;
        RECT 0.345 1.540 2.685 1.770 ;
        RECT 4.685 1.675 7.215 1.905 ;
        RECT 1.310 0.680 1.650 1.540 ;
        RECT 4.685 0.910 4.915 1.675 ;
        RECT 3.730 0.680 4.915 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xnor2_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__xnor2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xnor2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.760 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.170500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 2.630 3.850 2.860 ;
        RECT 1.830 1.770 2.090 2.630 ;
        RECT 3.620 2.400 3.850 2.630 ;
        RECT 3.620 2.170 4.510 2.400 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.170500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.755 3.090 4.855 3.320 ;
        RECT 0.755 2.455 0.985 3.090 ;
        RECT 4.625 2.830 4.855 3.090 ;
        RECT 4.625 2.600 5.475 2.830 ;
        RECT 0.710 1.770 0.985 2.455 ;
        RECT 5.245 2.115 5.475 2.600 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.459000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.665 3.270 7.895 3.685 ;
        RECT 7.430 2.890 7.895 3.270 ;
        RECT 7.665 1.950 7.895 2.890 ;
        RECT 9.855 1.950 10.135 3.685 ;
        RECT 7.665 1.720 10.135 1.950 ;
        RECT 7.665 0.680 7.895 1.720 ;
        RECT 9.905 0.680 10.135 1.720 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 11.760 5.490 ;
        RECT 2.665 3.875 2.895 4.590 ;
        RECT 6.645 3.875 6.875 4.590 ;
        RECT 8.735 3.875 8.965 4.590 ;
        RECT 10.925 2.875 11.155 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 12.190 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.190 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.020 ;
        RECT 2.485 0.450 2.715 1.020 ;
        RECT 5.825 0.450 6.055 1.425 ;
        RECT 6.545 0.450 6.775 1.425 ;
        RECT 8.785 0.450 9.015 1.490 ;
        RECT 11.025 0.450 11.255 1.490 ;
        RECT 0.000 -0.450 11.760 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.785 4.130 6.110 4.360 ;
        RECT 3.785 3.550 4.015 4.130 ;
        RECT 4.750 3.550 5.935 3.780 ;
        RECT 0.250 2.875 0.525 3.215 ;
        RECT 0.250 1.540 0.480 2.875 ;
        RECT 2.320 2.170 3.390 2.400 ;
        RECT 2.320 1.540 2.550 2.170 ;
        RECT 5.705 1.885 5.935 3.550 ;
        RECT 7.085 1.885 7.315 2.455 ;
        RECT 0.250 1.310 2.550 1.540 ;
        RECT 3.785 1.655 7.315 1.885 ;
        RECT 1.365 0.680 1.595 1.310 ;
        RECT 3.785 0.680 4.015 1.655 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xnor2_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__xnor3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xnor3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.880 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.995 2.330 3.900 2.710 ;
        RECT 1.995 1.815 2.225 2.330 ;
        RECT 3.670 2.100 3.900 2.330 ;
        RECT 3.670 1.870 4.510 2.100 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.300 2.940 5.475 3.170 ;
        RECT 1.300 2.150 1.530 2.940 ;
        RECT 0.870 1.770 1.530 2.150 ;
        RECT 5.245 1.815 5.475 2.940 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.560500 ;
    PORT
      LAYER Metal1 ;
        RECT 8.740 2.330 10.000 2.710 ;
        RECT 8.740 2.100 8.970 2.330 ;
        RECT 8.090 1.870 8.970 2.100 ;
        RECT 9.770 2.100 10.000 2.330 ;
        RECT 9.770 1.870 10.710 2.100 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.912500 ;
    PORT
      LAYER Metal1 ;
        RECT 9.985 3.720 10.215 4.360 ;
        RECT 9.985 3.645 11.855 3.720 ;
        RECT 9.985 3.490 12.190 3.645 ;
        RECT 11.685 3.415 12.190 3.490 ;
        RECT 11.960 1.590 12.190 3.415 ;
        RECT 10.950 1.210 12.190 1.590 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 12.880 5.490 ;
        RECT 2.435 3.550 2.665 4.590 ;
        RECT 6.545 3.855 6.775 4.590 ;
        RECT 8.815 3.875 9.045 4.590 ;
        RECT 12.025 3.875 12.255 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 13.310 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 13.310 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.080 ;
        RECT 2.485 0.450 2.715 1.080 ;
        RECT 5.825 0.450 6.055 1.080 ;
        RECT 8.585 0.450 8.815 1.080 ;
        RECT 0.000 -0.450 12.880 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.785 4.130 6.055 4.360 ;
        RECT 0.345 1.540 0.575 3.890 ;
        RECT 3.785 3.550 4.015 4.130 ;
        RECT 4.805 3.630 5.035 3.890 ;
        RECT 5.825 3.855 6.055 4.130 ;
        RECT 7.005 3.870 8.585 4.100 ;
        RECT 4.805 3.625 5.775 3.630 ;
        RECT 7.005 3.625 7.235 3.870 ;
        RECT 4.805 3.400 7.235 3.625 ;
        RECT 5.725 3.395 7.235 3.400 ;
        RECT 5.725 2.100 5.955 3.395 ;
        RECT 2.455 1.870 3.440 2.100 ;
        RECT 5.725 1.870 7.270 2.100 ;
        RECT 2.455 1.540 2.685 1.870 ;
        RECT 5.725 1.540 5.955 1.870 ;
        RECT 7.565 1.640 7.795 3.640 ;
        RECT 8.355 3.260 8.585 3.870 ;
        RECT 8.355 3.030 11.515 3.260 ;
        RECT 11.285 2.100 11.515 3.030 ;
        RECT 9.200 1.640 9.540 2.100 ;
        RECT 11.285 1.870 11.730 2.100 ;
        RECT 0.345 1.310 2.685 1.540 ;
        RECT 3.785 1.310 5.955 1.540 ;
        RECT 6.545 1.410 9.540 1.640 ;
        RECT 1.365 0.740 1.595 1.310 ;
        RECT 3.785 0.740 4.015 1.310 ;
        RECT 6.545 1.040 6.775 1.410 ;
        RECT 9.885 0.970 10.115 1.550 ;
        RECT 9.885 0.740 12.410 0.970 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xnor3_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__xnor3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xnor3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.680 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.165 1.950 2.395 2.520 ;
        RECT 4.070 2.180 4.575 2.520 ;
        RECT 4.070 1.950 4.330 2.180 ;
        RECT 2.165 1.720 4.330 1.950 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.025 3.210 5.595 3.440 ;
        RECT 1.025 2.180 1.255 3.210 ;
        RECT 5.190 2.180 5.595 3.210 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.560500 ;
    PORT
      LAYER Metal1 ;
        RECT 8.310 2.770 10.490 3.000 ;
        RECT 10.230 2.540 10.490 2.770 ;
        RECT 10.230 2.310 10.930 2.540 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.772000 ;
    PORT
      LAYER Metal1 ;
        RECT 13.015 3.385 13.245 4.360 ;
        RECT 15.155 3.385 15.385 4.360 ;
        RECT 13.015 3.155 15.385 3.385 ;
        RECT 13.915 1.945 14.145 3.155 ;
        RECT 12.965 1.715 15.435 1.945 ;
        RECT 12.965 0.845 13.290 1.715 ;
        RECT 15.205 0.845 15.435 1.715 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 15.680 5.490 ;
        RECT 2.605 3.670 2.835 4.590 ;
        RECT 8.805 3.615 9.035 4.590 ;
        RECT 14.035 3.615 14.265 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 16.110 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 16.110 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.365 0.450 0.595 1.185 ;
        RECT 2.605 0.450 2.835 1.185 ;
        RECT 5.945 0.450 6.175 1.185 ;
        RECT 6.665 0.450 6.895 1.185 ;
        RECT 9.085 0.450 9.315 1.180 ;
        RECT 12.245 0.450 12.475 1.160 ;
        RECT 14.085 0.450 14.315 1.485 ;
        RECT 0.000 -0.450 15.680 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.905 4.130 6.230 4.360 ;
        RECT 0.465 1.950 0.695 3.955 ;
        RECT 3.905 3.670 4.135 4.130 ;
        RECT 4.870 3.670 6.055 3.900 ;
        RECT 1.485 2.750 3.555 2.980 ;
        RECT 1.485 1.950 1.715 2.750 ;
        RECT 3.325 2.180 3.555 2.750 ;
        RECT 5.825 2.520 6.055 3.670 ;
        RECT 6.765 2.980 6.995 4.360 ;
        RECT 12.245 3.900 12.475 4.360 ;
        RECT 10.150 3.550 12.475 3.900 ;
        RECT 6.765 2.750 8.015 2.980 ;
        RECT 11.170 2.930 12.355 3.160 ;
        RECT 7.785 2.540 8.015 2.750 ;
        RECT 5.825 2.290 7.435 2.520 ;
        RECT 0.465 1.720 1.715 1.950 ;
        RECT 1.485 0.845 1.715 1.720 ;
        RECT 7.205 1.645 7.435 2.290 ;
        RECT 4.550 1.415 7.435 1.645 ;
        RECT 4.550 1.130 4.780 1.415 ;
        RECT 3.850 0.900 4.780 1.130 ;
        RECT 7.205 0.915 7.435 1.415 ;
        RECT 7.785 2.310 9.860 2.540 ;
        RECT 12.125 2.520 12.355 2.930 ;
        RECT 7.785 1.145 8.015 2.310 ;
        RECT 11.665 2.080 11.895 2.520 ;
        RECT 8.245 1.850 11.895 2.080 ;
        RECT 12.125 2.180 13.685 2.520 ;
        RECT 8.245 0.915 8.475 1.850 ;
        RECT 12.125 1.620 12.355 2.180 ;
        RECT 7.205 0.685 8.475 0.915 ;
        RECT 10.205 1.390 12.355 1.620 ;
        RECT 10.205 0.845 10.435 1.390 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xnor3_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__xnor3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xnor3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.920 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.859500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.990 2.000 2.330 2.360 ;
        RECT 3.990 2.000 4.330 2.395 ;
        RECT 1.990 1.770 4.330 2.000 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.859500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.960 3.050 3.970 3.280 ;
        RECT 0.960 2.110 1.190 3.050 ;
        RECT 3.510 2.890 3.970 3.050 ;
        RECT 3.740 2.855 3.970 2.890 ;
        RECT 3.740 2.625 5.350 2.855 ;
        RECT 5.010 2.165 5.350 2.625 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.170500 ;
    PORT
      LAYER Metal1 ;
        RECT 8.145 2.775 10.490 3.005 ;
        RECT 10.230 2.560 10.490 2.775 ;
        RECT 10.230 2.330 10.805 2.560 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.593000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.940 3.645 13.170 4.345 ;
        RECT 12.940 3.415 14.125 3.645 ;
        RECT 13.895 2.150 14.125 3.415 ;
        RECT 15.030 2.150 15.260 4.345 ;
        RECT 13.895 2.115 15.260 2.150 ;
        RECT 17.220 2.115 17.550 4.345 ;
        RECT 13.895 2.000 17.550 2.115 ;
        RECT 12.840 1.885 17.550 2.000 ;
        RECT 12.840 1.770 15.310 1.885 ;
        RECT 12.840 0.845 13.070 1.770 ;
        RECT 15.080 0.845 15.310 1.770 ;
        RECT 17.320 0.845 17.550 1.885 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.920 5.490 ;
        RECT 2.385 3.535 2.615 4.590 ;
        RECT 8.640 3.535 8.870 4.590 ;
        RECT 13.960 3.875 14.190 4.590 ;
        RECT 16.150 3.875 16.380 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 18.350 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 18.350 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 6.500 1.185 6.730 1.480 ;
        RECT 0.245 0.450 0.475 1.185 ;
        RECT 2.485 0.450 2.715 1.185 ;
        RECT 5.415 0.845 6.730 1.185 ;
        RECT 5.415 0.450 5.645 0.845 ;
        RECT 8.960 0.450 9.190 1.165 ;
        RECT 12.120 0.450 12.350 1.165 ;
        RECT 13.960 0.450 14.190 1.165 ;
        RECT 16.200 0.450 16.430 1.655 ;
        RECT 0.000 -0.450 17.920 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.605 4.105 6.110 4.335 ;
        RECT 0.345 1.880 0.575 3.875 ;
        RECT 3.605 3.535 3.835 4.105 ;
        RECT 4.625 3.315 4.855 3.875 ;
        RECT 5.880 3.535 6.110 4.105 ;
        RECT 10.080 4.130 12.350 4.360 ;
        RECT 4.625 3.085 5.810 3.315 ;
        RECT 1.420 2.590 3.290 2.820 ;
        RECT 1.420 1.880 1.650 2.590 ;
        RECT 5.580 1.940 5.810 3.085 ;
        RECT 6.600 2.910 6.830 3.875 ;
        RECT 10.080 3.550 10.310 4.130 ;
        RECT 6.600 2.680 7.850 2.910 ;
        RECT 7.620 2.545 7.850 2.680 ;
        RECT 11.100 2.545 11.330 3.900 ;
        RECT 12.120 3.550 12.350 4.130 ;
        RECT 7.040 1.940 7.270 2.450 ;
        RECT 5.580 1.935 7.270 1.940 ;
        RECT 0.345 1.650 1.650 1.880 ;
        RECT 1.365 0.845 1.650 1.650 ;
        RECT 4.560 1.710 7.270 1.935 ;
        RECT 4.560 1.705 5.630 1.710 ;
        RECT 4.560 1.130 4.790 1.705 ;
        RECT 3.550 0.900 4.790 1.130 ;
        RECT 7.040 0.910 7.270 1.710 ;
        RECT 7.620 2.315 9.785 2.545 ;
        RECT 11.100 2.315 13.665 2.545 ;
        RECT 7.620 1.140 7.850 2.315 ;
        RECT 12.055 2.230 13.665 2.315 ;
        RECT 8.080 1.855 11.825 2.085 ;
        RECT 8.080 0.910 8.310 1.855 ;
        RECT 12.055 1.625 12.285 2.230 ;
        RECT 7.040 0.680 8.310 0.910 ;
        RECT 10.080 1.395 12.285 1.625 ;
        RECT 10.080 0.815 10.310 1.395 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xnor3_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__xor2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xor2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.720 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.560500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.640 2.330 4.115 2.710 ;
        RECT 2.640 2.135 2.870 2.330 ;
        RECT 1.940 1.905 2.870 2.135 ;
        RECT 3.885 2.190 4.115 2.330 ;
        RECT 3.885 1.850 4.455 2.190 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.560500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.940 4.575 3.170 ;
        RECT 0.710 1.850 1.015 2.940 ;
        RECT 4.345 2.700 4.575 2.940 ;
        RECT 4.345 2.470 5.060 2.700 ;
        RECT 4.830 2.135 5.060 2.470 ;
        RECT 4.830 1.905 5.530 2.135 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.805 3.270 5.035 3.900 ;
        RECT 4.805 3.120 5.450 3.270 ;
        RECT 4.805 3.040 5.990 3.120 ;
        RECT 5.190 2.890 5.990 3.040 ;
        RECT 5.760 1.620 5.990 2.890 ;
        RECT 3.785 1.390 5.990 1.620 ;
        RECT 3.785 0.810 4.015 1.390 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 6.720 5.490 ;
        RECT 2.435 3.400 2.665 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 7.150 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.150 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.150 ;
        RECT 2.485 0.450 2.715 1.150 ;
        RECT 5.825 0.450 6.055 1.160 ;
        RECT 0.000 -0.450 6.720 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.785 4.130 6.055 4.360 ;
        RECT 0.250 3.400 0.575 3.740 ;
        RECT 3.785 3.400 4.015 4.130 ;
        RECT 5.825 3.400 6.055 4.130 ;
        RECT 0.250 1.620 0.480 3.400 ;
        RECT 3.100 1.620 3.440 2.100 ;
        RECT 0.250 1.390 3.440 1.620 ;
        RECT 1.365 0.810 1.595 1.390 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xor2_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__xor2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xor2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.560500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.320 2.500 4.355 2.730 ;
        RECT 2.320 2.100 2.550 2.500 ;
        RECT 1.790 1.870 2.550 2.100 ;
        RECT 4.070 1.770 4.355 2.500 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.560500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.860 2.960 5.375 3.190 ;
        RECT 1.860 2.710 2.090 2.960 ;
        RECT 1.270 2.465 2.090 2.710 ;
        RECT 0.770 2.330 2.090 2.465 ;
        RECT 0.770 2.235 1.460 2.330 ;
        RECT 5.145 2.180 5.375 2.960 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.665 1.590 7.895 4.230 ;
        RECT 7.430 1.210 7.895 1.590 ;
        RECT 7.665 0.840 7.895 1.210 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 9.520 5.490 ;
        RECT 0.245 3.585 0.475 4.590 ;
        RECT 2.285 3.585 2.515 4.590 ;
        RECT 5.725 3.880 5.955 4.590 ;
        RECT 6.645 3.585 6.875 4.590 ;
        RECT 8.685 3.585 8.915 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 9.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.285 0.450 2.515 1.180 ;
        RECT 6.545 0.450 6.775 1.445 ;
        RECT 8.785 0.450 9.015 1.650 ;
        RECT 0.000 -0.450 9.520 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.265 3.170 1.495 4.310 ;
        RECT 3.685 3.650 3.915 4.230 ;
        RECT 3.685 3.420 5.835 3.650 ;
        RECT 0.245 2.940 1.495 3.170 ;
        RECT 0.245 1.640 0.475 2.940 ;
        RECT 2.955 1.640 3.185 2.270 ;
        RECT 5.605 2.110 5.835 3.420 ;
        RECT 5.605 1.950 7.370 2.110 ;
        RECT 4.705 1.880 7.370 1.950 ;
        RECT 4.705 1.720 5.825 1.880 ;
        RECT 0.245 1.410 3.185 1.640 ;
        RECT 0.245 0.840 0.475 1.410 ;
        RECT 3.585 0.910 3.815 1.650 ;
        RECT 4.705 1.140 4.935 1.720 ;
        RECT 5.825 0.910 6.055 1.490 ;
        RECT 3.585 0.680 6.055 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xor2_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__xor2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xor2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.760 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.170500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.790 2.330 4.360 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.170500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.770 2.940 4.860 3.170 ;
        RECT 0.770 2.330 1.110 2.940 ;
        RECT 4.630 2.710 4.860 2.940 ;
        RECT 4.630 2.330 5.430 2.710 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.459000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.430 3.450 7.895 4.360 ;
        RECT 7.665 2.115 7.895 3.450 ;
        RECT 9.855 2.115 10.135 4.360 ;
        RECT 7.665 1.885 10.135 2.115 ;
        RECT 7.665 0.845 7.895 1.885 ;
        RECT 9.905 0.845 10.135 1.885 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 11.760 5.490 ;
        RECT 0.245 3.860 0.475 4.590 ;
        RECT 2.285 3.860 2.515 4.590 ;
        RECT 5.725 3.860 5.955 4.590 ;
        RECT 6.645 3.860 6.875 4.590 ;
        RECT 8.735 3.860 8.965 4.590 ;
        RECT 10.925 3.860 11.155 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 12.190 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.190 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.230 0.450 2.570 1.595 ;
        RECT 6.545 0.450 6.775 1.165 ;
        RECT 8.785 0.450 9.015 1.655 ;
        RECT 11.025 0.450 11.255 1.655 ;
        RECT 0.000 -0.450 11.760 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.265 3.630 1.495 4.065 ;
        RECT 0.190 3.400 1.495 3.630 ;
        RECT 3.635 3.630 3.865 4.360 ;
        RECT 3.635 3.400 5.890 3.630 ;
        RECT 0.190 2.100 0.420 3.400 ;
        RECT 5.660 2.210 5.890 3.400 ;
        RECT 5.660 2.100 7.315 2.210 ;
        RECT 0.190 1.870 3.290 2.100 ;
        RECT 4.705 1.870 7.315 2.100 ;
        RECT 0.190 1.365 0.530 1.870 ;
        RECT 3.585 1.060 3.815 1.650 ;
        RECT 4.705 1.310 4.935 1.870 ;
        RECT 5.825 1.060 6.055 1.640 ;
        RECT 3.585 0.830 6.055 1.060 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xor2_4

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__xor3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xor3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.880 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.890 1.770 2.650 2.155 ;
        RECT 2.420 1.640 2.650 1.770 ;
        RECT 4.225 1.640 4.455 2.210 ;
        RECT 2.420 1.410 4.455 1.640 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.925 3.075 1.530 3.270 ;
        RECT 0.925 2.845 5.475 3.075 ;
        RECT 0.925 1.870 1.155 2.845 ;
        RECT 5.245 1.870 5.475 2.845 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.560500 ;
    PORT
      LAYER Metal1 ;
        RECT 7.990 2.480 10.755 2.710 ;
        RECT 7.990 2.330 8.335 2.480 ;
        RECT 10.525 1.870 10.755 2.480 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 11.105 3.270 11.335 3.700 ;
        RECT 11.105 2.890 12.235 3.270 ;
        RECT 12.005 1.155 12.235 2.890 ;
        RECT 10.030 0.925 12.235 1.155 ;
        RECT 10.030 0.895 10.370 0.925 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 12.880 5.490 ;
        RECT 2.385 3.305 2.615 4.590 ;
        RECT 8.685 2.965 8.915 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 13.310 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 13.310 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.180 ;
        RECT 2.485 0.450 2.715 1.180 ;
        RECT 5.825 0.450 6.055 1.180 ;
        RECT 6.545 0.450 6.775 1.180 ;
        RECT 8.785 0.450 9.015 1.180 ;
        RECT 12.125 0.450 12.355 0.695 ;
        RECT 0.000 -0.450 12.880 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.785 3.830 6.110 4.115 ;
        RECT 10.085 4.005 12.635 4.235 ;
        RECT 0.345 1.640 0.575 3.645 ;
        RECT 3.785 3.305 4.015 3.830 ;
        RECT 4.750 3.360 5.935 3.590 ;
        RECT 1.385 2.385 3.335 2.615 ;
        RECT 1.385 1.640 1.615 2.385 ;
        RECT 3.105 1.870 3.335 2.385 ;
        RECT 5.705 1.640 5.935 3.360 ;
        RECT 6.630 2.670 6.860 3.775 ;
        RECT 10.085 3.305 10.315 4.005 ;
        RECT 12.405 3.425 12.635 4.005 ;
        RECT 6.630 2.440 7.760 2.670 ;
        RECT 7.070 1.640 7.300 2.210 ;
        RECT 7.530 2.100 7.760 2.440 ;
        RECT 9.400 2.100 9.740 2.155 ;
        RECT 7.530 1.890 9.740 2.100 ;
        RECT 0.345 1.410 1.615 1.640 ;
        RECT 1.365 0.840 1.615 1.410 ;
        RECT 4.685 1.620 7.300 1.640 ;
        RECT 7.665 1.870 9.740 1.890 ;
        RECT 4.685 1.410 7.435 1.620 ;
        RECT 4.685 1.125 4.915 1.410 ;
        RECT 3.730 0.895 4.915 1.125 ;
        RECT 7.205 0.910 7.435 1.410 ;
        RECT 7.665 1.140 7.895 1.870 ;
        RECT 11.545 1.640 11.775 2.210 ;
        RECT 8.325 1.410 11.775 1.640 ;
        RECT 8.325 0.910 8.555 1.410 ;
        RECT 7.205 0.680 8.555 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xor3_1

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__xor3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xor3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.680 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.740 2.170 2.200 ;
        RECT 4.225 1.740 4.455 2.025 ;
        RECT 1.830 1.510 4.455 1.740 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.910 2.890 3.900 3.270 ;
        RECT 0.910 1.915 1.140 2.890 ;
        RECT 3.670 2.485 3.900 2.890 ;
        RECT 3.670 2.255 5.530 2.485 ;
        RECT 5.190 1.970 5.530 2.255 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.560500 ;
    PORT
      LAYER Metal1 ;
        RECT 8.090 2.370 10.710 2.710 ;
        RECT 9.670 2.330 10.710 2.370 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.772000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.845 3.645 13.075 4.320 ;
        RECT 12.845 3.415 14.030 3.645 ;
        RECT 13.800 1.670 14.030 3.415 ;
        RECT 14.985 1.670 15.315 3.685 ;
        RECT 12.845 1.440 15.315 1.670 ;
        RECT 12.845 0.845 13.290 1.440 ;
        RECT 15.085 0.845 15.315 1.440 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 15.680 5.490 ;
        RECT 2.435 3.510 2.665 4.590 ;
        RECT 6.545 3.450 6.775 4.590 ;
        RECT 8.815 4.350 9.045 4.590 ;
        RECT 12.025 4.350 12.255 4.590 ;
        RECT 13.865 3.875 14.095 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 16.110 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 16.110 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.185 ;
        RECT 2.485 0.450 2.715 1.185 ;
        RECT 5.825 0.450 6.055 1.185 ;
        RECT 8.585 0.450 8.815 1.185 ;
        RECT 13.965 0.450 14.195 1.165 ;
        RECT 0.000 -0.450 15.680 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.785 4.130 6.055 4.360 ;
        RECT 0.345 1.685 0.575 3.850 ;
        RECT 3.785 3.510 4.015 4.130 ;
        RECT 4.805 2.945 5.035 3.900 ;
        RECT 5.825 3.175 6.055 4.130 ;
        RECT 9.930 4.135 11.360 4.155 ;
        RECT 9.930 3.925 11.940 4.135 ;
        RECT 11.265 3.905 11.940 3.925 ;
        RECT 7.005 3.465 11.170 3.695 ;
        RECT 7.005 2.945 7.235 3.465 ;
        RECT 4.805 2.715 7.235 2.945 ;
        RECT 1.370 2.430 3.440 2.660 ;
        RECT 1.370 1.685 1.600 2.430 ;
        RECT 3.100 1.970 3.440 2.430 ;
        RECT 0.345 1.455 1.600 1.685 ;
        RECT 7.005 1.645 7.235 2.715 ;
        RECT 1.365 0.845 1.600 1.455 ;
        RECT 4.685 1.415 7.235 1.645 ;
        RECT 7.565 2.140 7.795 3.235 ;
        RECT 10.940 2.410 11.170 3.465 ;
        RECT 11.710 2.870 11.940 3.905 ;
        RECT 11.710 2.640 12.190 2.870 ;
        RECT 10.940 2.180 11.730 2.410 ;
        RECT 7.565 1.910 9.540 2.140 ;
        RECT 11.960 2.130 12.190 2.640 ;
        RECT 11.960 1.950 13.570 2.130 ;
        RECT 4.685 1.130 4.915 1.415 ;
        RECT 7.565 1.130 7.795 1.910 ;
        RECT 11.005 1.900 13.570 1.950 ;
        RECT 11.005 1.720 12.185 1.900 ;
        RECT 3.730 0.900 4.915 1.130 ;
        RECT 6.490 0.900 7.795 1.130 ;
        RECT 9.885 0.910 10.115 1.655 ;
        RECT 11.005 1.140 11.235 1.720 ;
        RECT 12.125 0.910 12.355 1.490 ;
        RECT 9.885 0.680 12.355 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xor3_2

#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__xor3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xor3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.920 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.859500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 2.005 2.170 2.135 ;
        RECT 4.045 2.005 4.275 2.520 ;
        RECT 1.830 1.775 4.275 2.005 ;
        RECT 1.830 1.210 2.090 1.775 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.859500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.905 3.005 2.880 3.055 ;
        RECT 0.905 2.825 4.860 3.005 ;
        RECT 0.905 2.180 1.135 2.825 ;
        RECT 2.735 2.775 4.860 2.825 ;
        RECT 4.630 2.710 4.860 2.775 ;
        RECT 4.630 2.180 5.295 2.710 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.170500 ;
    PORT
      LAYER Metal1 ;
        RECT 7.910 2.475 10.480 2.710 ;
        RECT 9.670 2.330 10.480 2.475 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.593000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.765 3.465 12.995 4.360 ;
        RECT 12.765 3.235 13.950 3.465 ;
        RECT 13.720 2.030 13.950 3.235 ;
        RECT 14.955 2.115 15.185 4.360 ;
        RECT 17.045 2.115 17.375 4.360 ;
        RECT 14.955 2.030 17.375 2.115 ;
        RECT 13.720 1.885 17.375 2.030 ;
        RECT 13.720 1.720 15.135 1.885 ;
        RECT 13.590 1.490 15.135 1.720 ;
        RECT 12.665 1.210 15.135 1.490 ;
        RECT 12.665 0.680 12.895 1.210 ;
        RECT 14.905 0.845 15.135 1.210 ;
        RECT 17.145 0.845 17.375 1.885 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.920 5.490 ;
        RECT 2.385 3.695 2.615 4.590 ;
        RECT 6.365 3.015 6.595 4.590 ;
        RECT 8.685 3.865 8.915 4.590 ;
        RECT 11.845 4.350 12.075 4.590 ;
        RECT 13.785 3.695 14.015 4.590 ;
        RECT 15.975 3.695 16.205 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 18.350 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 18.350 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.185 ;
        RECT 2.485 0.450 2.715 1.185 ;
        RECT 5.645 0.450 5.875 1.185 ;
        RECT 8.405 0.450 8.635 1.185 ;
        RECT 13.785 0.450 14.015 0.695 ;
        RECT 16.025 0.450 16.255 1.655 ;
        RECT 0.000 -0.450 17.920 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.605 4.130 5.875 4.360 ;
        RECT 0.345 1.950 0.575 4.035 ;
        RECT 3.605 3.695 3.835 4.130 ;
        RECT 4.625 3.465 4.855 3.900 ;
        RECT 5.645 3.695 5.875 4.130 ;
        RECT 9.700 3.865 11.955 4.095 ;
        RECT 6.825 3.635 8.545 3.680 ;
        RECT 4.625 3.235 5.755 3.465 ;
        RECT 1.365 2.465 2.590 2.595 ;
        RECT 1.365 2.365 3.310 2.465 ;
        RECT 1.365 1.950 1.595 2.365 ;
        RECT 2.380 2.235 3.310 2.365 ;
        RECT 5.525 2.410 5.755 3.235 ;
        RECT 6.825 3.450 11.495 3.635 ;
        RECT 6.825 2.410 7.055 3.450 ;
        RECT 8.405 3.405 11.495 3.450 ;
        RECT 0.345 1.720 1.595 1.950 ;
        RECT 1.365 0.845 1.595 1.720 ;
        RECT 5.525 2.180 7.055 2.410 ;
        RECT 7.385 2.245 7.615 3.220 ;
        RECT 5.525 1.645 5.755 2.180 ;
        RECT 7.385 2.015 9.410 2.245 ;
        RECT 11.265 2.180 11.495 3.405 ;
        RECT 11.725 2.160 11.955 3.865 ;
        RECT 7.385 1.950 7.615 2.015 ;
        RECT 11.725 1.950 13.490 2.160 ;
        RECT 4.465 1.415 5.755 1.645 ;
        RECT 6.365 1.720 7.615 1.950 ;
        RECT 10.825 1.930 13.490 1.950 ;
        RECT 10.825 1.720 11.955 1.930 ;
        RECT 4.465 1.130 4.695 1.415 ;
        RECT 3.550 0.900 4.695 1.130 ;
        RECT 6.365 0.845 6.595 1.720 ;
        RECT 9.705 0.910 9.935 1.655 ;
        RECT 10.825 1.315 11.055 1.720 ;
        RECT 11.945 0.910 12.175 1.490 ;
        RECT 9.705 0.680 12.175 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xor3_4

#--------EOF---------


END LIBRARY
