magic
tech gf180mcuA
timestamp 1698431365
<< properties >>
string GDS_END 1001750
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 1000418
<< end >>
