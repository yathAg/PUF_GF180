magic
tech gf180mcuB
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -3832 3921 164 17697
<< pwell >>
rect 2092 11351 4268 16351
rect 4528 11351 6704 16351
rect 6964 11351 9140 16351
rect 9400 11351 11576 16351
rect 2092 5339 4268 10339
rect 4528 5339 6704 10339
rect 6964 5339 9140 10339
rect 9400 5339 11576 10339
<< mvndiff >>
rect 2092 16314 2180 16351
rect 2092 11388 2105 16314
rect 2151 11388 2180 16314
rect 2092 11351 2180 11388
rect 4180 16314 4268 16351
rect 4180 11388 4209 16314
rect 4255 11388 4268 16314
rect 4180 11351 4268 11388
rect 4528 16314 4616 16351
rect 4528 11388 4541 16314
rect 4587 11388 4616 16314
rect 4528 11351 4616 11388
rect 6616 16314 6704 16351
rect 6616 11388 6645 16314
rect 6691 11388 6704 16314
rect 6616 11351 6704 11388
rect 6964 16314 7052 16351
rect 6964 11388 6977 16314
rect 7023 11388 7052 16314
rect 6964 11351 7052 11388
rect 9052 16314 9140 16351
rect 9052 11388 9081 16314
rect 9127 11388 9140 16314
rect 9052 11351 9140 11388
rect 9400 16314 9488 16351
rect 9400 11388 9413 16314
rect 9459 11388 9488 16314
rect 9400 11351 9488 11388
rect 11488 16314 11576 16351
rect 11488 11388 11517 16314
rect 11563 11388 11576 16314
rect 11488 11351 11576 11388
rect 2092 10302 2180 10339
rect 2092 5376 2105 10302
rect 2151 5376 2180 10302
rect 2092 5339 2180 5376
rect 4180 10302 4268 10339
rect 4180 5376 4209 10302
rect 4255 5376 4268 10302
rect 4180 5339 4268 5376
rect 4528 10302 4616 10339
rect 4528 5376 4541 10302
rect 4587 5376 4616 10302
rect 4528 5339 4616 5376
rect 6616 10302 6704 10339
rect 6616 5376 6645 10302
rect 6691 5376 6704 10302
rect 6616 5339 6704 5376
rect 6964 10302 7052 10339
rect 6964 5376 6977 10302
rect 7023 5376 7052 10302
rect 6964 5339 7052 5376
rect 9052 10302 9140 10339
rect 9052 5376 9081 10302
rect 9127 5376 9140 10302
rect 9052 5339 9140 5376
rect 9400 10302 9488 10339
rect 9400 5376 9413 10302
rect 9459 5376 9488 10302
rect 9400 5339 9488 5376
rect 11488 10302 11576 10339
rect 11488 5376 11517 10302
rect 11563 5376 11576 10302
rect 11488 5339 11576 5376
<< mvndiffc >>
rect 2105 11388 2151 16314
rect 4209 11388 4255 16314
rect 4541 11388 4587 16314
rect 6645 11388 6691 16314
rect 6977 11388 7023 16314
rect 9081 11388 9127 16314
rect 9413 11388 9459 16314
rect 11517 11388 11563 16314
rect 2105 5376 2151 10302
rect 4209 5376 4255 10302
rect 4541 5376 4587 10302
rect 6645 5376 6691 10302
rect 6977 5376 7023 10302
rect 9081 5376 9127 10302
rect 9413 5376 9459 10302
rect 11517 5376 11563 10302
<< psubdiff >>
rect 1565 17016 12109 17038
rect 1565 16970 1587 17016
rect 1633 16970 1701 17016
rect 1747 16970 1855 17016
rect 1901 16970 1969 17016
rect 2015 16970 2083 17016
rect 2129 16970 2197 17016
rect 2243 16970 2311 17016
rect 2357 16970 2425 17016
rect 2471 16970 2539 17016
rect 2585 16970 2653 17016
rect 2699 16970 2767 17016
rect 2813 16970 2881 17016
rect 2927 16970 2995 17016
rect 3041 16970 3109 17016
rect 3155 16970 3223 17016
rect 3269 16970 3337 17016
rect 3383 16970 3451 17016
rect 3497 16970 3565 17016
rect 3611 16970 3679 17016
rect 3725 16970 3793 17016
rect 3839 16970 3907 17016
rect 3953 16970 4021 17016
rect 4067 16970 4135 17016
rect 4181 16970 4249 17016
rect 4295 16970 4363 17016
rect 4409 16970 4477 17016
rect 4523 16970 4591 17016
rect 4637 16970 4705 17016
rect 4751 16970 4819 17016
rect 4865 16970 4933 17016
rect 4979 16970 5047 17016
rect 5093 16970 5161 17016
rect 5207 16970 5275 17016
rect 5321 16970 5389 17016
rect 5435 16970 5503 17016
rect 5549 16970 5617 17016
rect 5663 16970 5731 17016
rect 5777 16970 5845 17016
rect 5891 16970 5959 17016
rect 6005 16970 6073 17016
rect 6119 16970 6187 17016
rect 6233 16970 6301 17016
rect 6347 16970 6415 17016
rect 6461 16970 6529 17016
rect 6575 16970 6643 17016
rect 6689 16970 6757 17016
rect 6803 16970 6871 17016
rect 6917 16970 6985 17016
rect 7031 16970 7099 17016
rect 7145 16970 7213 17016
rect 7259 16970 7327 17016
rect 7373 16970 7441 17016
rect 7487 16970 7555 17016
rect 7601 16970 7669 17016
rect 7715 16970 7783 17016
rect 7829 16970 7897 17016
rect 7943 16970 8011 17016
rect 8057 16970 8125 17016
rect 8171 16970 8239 17016
rect 8285 16970 8353 17016
rect 8399 16970 8467 17016
rect 8513 16970 8581 17016
rect 8627 16970 8695 17016
rect 8741 16970 8809 17016
rect 8855 16970 8923 17016
rect 8969 16970 9037 17016
rect 9083 16970 9151 17016
rect 9197 16970 9265 17016
rect 9311 16970 9379 17016
rect 9425 16970 9493 17016
rect 9539 16970 9607 17016
rect 9653 16970 9721 17016
rect 9767 16970 9835 17016
rect 9881 16970 9949 17016
rect 9995 16970 10063 17016
rect 10109 16970 10177 17016
rect 10223 16970 10291 17016
rect 10337 16970 10405 17016
rect 10451 16970 10519 17016
rect 10565 16970 10633 17016
rect 10679 16970 10747 17016
rect 10793 16970 10861 17016
rect 10907 16970 10975 17016
rect 11021 16970 11089 17016
rect 11135 16970 11203 17016
rect 11249 16970 11317 17016
rect 11363 16970 11431 17016
rect 11477 16970 11545 17016
rect 11591 16970 11659 17016
rect 11705 16970 11773 17016
rect 11819 16970 11927 17016
rect 11973 16970 12041 17016
rect 12087 16970 12109 17016
rect 1565 16902 12109 16970
rect 1565 16856 1587 16902
rect 1633 16856 1701 16902
rect 1747 16856 1855 16902
rect 1901 16856 1969 16902
rect 2015 16856 2083 16902
rect 2129 16856 2197 16902
rect 2243 16856 2311 16902
rect 2357 16856 2425 16902
rect 2471 16856 2539 16902
rect 2585 16856 2653 16902
rect 2699 16856 2767 16902
rect 2813 16856 2881 16902
rect 2927 16856 2995 16902
rect 3041 16856 3109 16902
rect 3155 16856 3223 16902
rect 3269 16856 3337 16902
rect 3383 16856 3451 16902
rect 3497 16856 3565 16902
rect 3611 16856 3679 16902
rect 3725 16856 3793 16902
rect 3839 16856 3907 16902
rect 3953 16856 4021 16902
rect 4067 16856 4135 16902
rect 4181 16856 4249 16902
rect 4295 16856 4363 16902
rect 4409 16856 4477 16902
rect 4523 16856 4591 16902
rect 4637 16856 4705 16902
rect 4751 16856 4819 16902
rect 4865 16856 4933 16902
rect 4979 16856 5047 16902
rect 5093 16856 5161 16902
rect 5207 16856 5275 16902
rect 5321 16856 5389 16902
rect 5435 16856 5503 16902
rect 5549 16856 5617 16902
rect 5663 16856 5731 16902
rect 5777 16856 5845 16902
rect 5891 16856 5959 16902
rect 6005 16856 6073 16902
rect 6119 16856 6187 16902
rect 6233 16856 6301 16902
rect 6347 16856 6415 16902
rect 6461 16856 6529 16902
rect 6575 16856 6643 16902
rect 6689 16856 6757 16902
rect 6803 16856 6871 16902
rect 6917 16856 6985 16902
rect 7031 16856 7099 16902
rect 7145 16856 7213 16902
rect 7259 16856 7327 16902
rect 7373 16856 7441 16902
rect 7487 16856 7555 16902
rect 7601 16856 7669 16902
rect 7715 16856 7783 16902
rect 7829 16856 7897 16902
rect 7943 16856 8011 16902
rect 8057 16856 8125 16902
rect 8171 16856 8239 16902
rect 8285 16856 8353 16902
rect 8399 16856 8467 16902
rect 8513 16856 8581 16902
rect 8627 16856 8695 16902
rect 8741 16856 8809 16902
rect 8855 16856 8923 16902
rect 8969 16856 9037 16902
rect 9083 16856 9151 16902
rect 9197 16856 9265 16902
rect 9311 16856 9379 16902
rect 9425 16856 9493 16902
rect 9539 16856 9607 16902
rect 9653 16856 9721 16902
rect 9767 16856 9835 16902
rect 9881 16856 9949 16902
rect 9995 16856 10063 16902
rect 10109 16856 10177 16902
rect 10223 16856 10291 16902
rect 10337 16856 10405 16902
rect 10451 16856 10519 16902
rect 10565 16856 10633 16902
rect 10679 16856 10747 16902
rect 10793 16856 10861 16902
rect 10907 16856 10975 16902
rect 11021 16856 11089 16902
rect 11135 16856 11203 16902
rect 11249 16856 11317 16902
rect 11363 16856 11431 16902
rect 11477 16856 11545 16902
rect 11591 16856 11659 16902
rect 11705 16856 11773 16902
rect 11819 16856 11927 16902
rect 11973 16856 12041 16902
rect 12087 16856 12109 16902
rect 1565 16834 12109 16856
rect 1565 16788 1769 16834
rect 1565 16742 1587 16788
rect 1633 16742 1701 16788
rect 1747 16742 1769 16788
rect 1565 16218 1769 16742
rect 11905 16788 12109 16834
rect 11905 16742 11927 16788
rect 11973 16742 12041 16788
rect 12087 16742 12109 16788
rect 11905 16674 12109 16742
rect 11905 16628 11927 16674
rect 11973 16628 12041 16674
rect 12087 16628 12109 16674
rect 11905 16560 12109 16628
rect 11905 16514 11927 16560
rect 11973 16514 12041 16560
rect 12087 16514 12109 16560
rect 11905 16446 12109 16514
rect 11905 16400 11927 16446
rect 11973 16400 12041 16446
rect 12087 16400 12109 16446
rect 1565 16172 1587 16218
rect 1633 16172 1701 16218
rect 1747 16172 1769 16218
rect 1565 16104 1769 16172
rect 1565 16058 1587 16104
rect 1633 16058 1701 16104
rect 1747 16058 1769 16104
rect 1565 15990 1769 16058
rect 1565 15944 1587 15990
rect 1633 15944 1701 15990
rect 1747 15944 1769 15990
rect 1565 15876 1769 15944
rect 1565 15830 1587 15876
rect 1633 15830 1701 15876
rect 1747 15830 1769 15876
rect 1565 15762 1769 15830
rect 1565 15716 1587 15762
rect 1633 15716 1701 15762
rect 1747 15716 1769 15762
rect 1565 15648 1769 15716
rect 1565 15602 1587 15648
rect 1633 15602 1701 15648
rect 1747 15602 1769 15648
rect 1565 15534 1769 15602
rect 1565 15488 1587 15534
rect 1633 15488 1701 15534
rect 1747 15488 1769 15534
rect 1565 15420 1769 15488
rect 1565 15374 1587 15420
rect 1633 15374 1701 15420
rect 1747 15374 1769 15420
rect 1565 15306 1769 15374
rect 1565 15260 1587 15306
rect 1633 15260 1701 15306
rect 1747 15260 1769 15306
rect 1565 15192 1769 15260
rect 1565 15146 1587 15192
rect 1633 15146 1701 15192
rect 1747 15146 1769 15192
rect 1565 15078 1769 15146
rect 1565 15032 1587 15078
rect 1633 15032 1701 15078
rect 1747 15032 1769 15078
rect 1565 14964 1769 15032
rect 1565 14918 1587 14964
rect 1633 14918 1701 14964
rect 1747 14918 1769 14964
rect 1565 14850 1769 14918
rect 1565 14804 1587 14850
rect 1633 14804 1701 14850
rect 1747 14804 1769 14850
rect 1565 14736 1769 14804
rect 1565 14690 1587 14736
rect 1633 14690 1701 14736
rect 1747 14690 1769 14736
rect 1565 14622 1769 14690
rect 1565 14576 1587 14622
rect 1633 14576 1701 14622
rect 1747 14576 1769 14622
rect 1565 14508 1769 14576
rect 1565 14462 1587 14508
rect 1633 14462 1701 14508
rect 1747 14462 1769 14508
rect 1565 14394 1769 14462
rect 1565 14348 1587 14394
rect 1633 14348 1701 14394
rect 1747 14348 1769 14394
rect 1565 14280 1769 14348
rect 1565 14234 1587 14280
rect 1633 14234 1701 14280
rect 1747 14234 1769 14280
rect 1565 14166 1769 14234
rect 1565 14120 1587 14166
rect 1633 14120 1701 14166
rect 1747 14120 1769 14166
rect 1565 14052 1769 14120
rect 1565 14006 1587 14052
rect 1633 14006 1701 14052
rect 1747 14006 1769 14052
rect 1565 13938 1769 14006
rect 1565 13892 1587 13938
rect 1633 13892 1701 13938
rect 1747 13892 1769 13938
rect 1565 13824 1769 13892
rect 1565 13778 1587 13824
rect 1633 13778 1701 13824
rect 1747 13778 1769 13824
rect 1565 13710 1769 13778
rect 1565 13664 1587 13710
rect 1633 13664 1701 13710
rect 1747 13664 1769 13710
rect 1565 13596 1769 13664
rect 1565 13550 1587 13596
rect 1633 13550 1701 13596
rect 1747 13550 1769 13596
rect 1565 13482 1769 13550
rect 1565 13436 1587 13482
rect 1633 13436 1701 13482
rect 1747 13436 1769 13482
rect 1565 13368 1769 13436
rect 1565 13322 1587 13368
rect 1633 13322 1701 13368
rect 1747 13322 1769 13368
rect 1565 13254 1769 13322
rect 1565 13208 1587 13254
rect 1633 13208 1701 13254
rect 1747 13208 1769 13254
rect 1565 13140 1769 13208
rect 1565 13094 1587 13140
rect 1633 13094 1701 13140
rect 1747 13094 1769 13140
rect 1565 13026 1769 13094
rect 1565 12980 1587 13026
rect 1633 12980 1701 13026
rect 1747 12980 1769 13026
rect 1565 12912 1769 12980
rect 1565 12866 1587 12912
rect 1633 12866 1701 12912
rect 1747 12866 1769 12912
rect 1565 12798 1769 12866
rect 1565 12752 1587 12798
rect 1633 12752 1701 12798
rect 1747 12752 1769 12798
rect 1565 12684 1769 12752
rect 1565 12638 1587 12684
rect 1633 12638 1701 12684
rect 1747 12638 1769 12684
rect 1565 12570 1769 12638
rect 1565 12524 1587 12570
rect 1633 12524 1701 12570
rect 1747 12524 1769 12570
rect 1565 12456 1769 12524
rect 1565 12410 1587 12456
rect 1633 12410 1701 12456
rect 1747 12410 1769 12456
rect 1565 12342 1769 12410
rect 1565 12296 1587 12342
rect 1633 12296 1701 12342
rect 1747 12296 1769 12342
rect 1565 12228 1769 12296
rect 1565 12182 1587 12228
rect 1633 12182 1701 12228
rect 1747 12182 1769 12228
rect 1565 12114 1769 12182
rect 1565 12068 1587 12114
rect 1633 12068 1701 12114
rect 1747 12068 1769 12114
rect 1565 12000 1769 12068
rect 1565 11954 1587 12000
rect 1633 11954 1701 12000
rect 1747 11954 1769 12000
rect 1565 11886 1769 11954
rect 1565 11840 1587 11886
rect 1633 11840 1701 11886
rect 1747 11840 1769 11886
rect 1565 11772 1769 11840
rect 1565 11726 1587 11772
rect 1633 11726 1701 11772
rect 1747 11726 1769 11772
rect 1565 11658 1769 11726
rect 1565 11612 1587 11658
rect 1633 11612 1701 11658
rect 1747 11612 1769 11658
rect 1565 11544 1769 11612
rect 1565 11498 1587 11544
rect 1633 11498 1701 11544
rect 1747 11498 1769 11544
rect 1565 11430 1769 11498
rect 1565 11384 1587 11430
rect 1633 11384 1701 11430
rect 1747 11384 1769 11430
rect 1565 11316 1769 11384
rect 11905 16332 12109 16400
rect 11905 16286 11927 16332
rect 11973 16286 12041 16332
rect 12087 16286 12109 16332
rect 11905 16218 12109 16286
rect 11905 16172 11927 16218
rect 11973 16172 12041 16218
rect 12087 16172 12109 16218
rect 11905 16104 12109 16172
rect 11905 16058 11927 16104
rect 11973 16058 12041 16104
rect 12087 16058 12109 16104
rect 11905 15990 12109 16058
rect 11905 15944 11927 15990
rect 11973 15944 12041 15990
rect 12087 15944 12109 15990
rect 11905 15876 12109 15944
rect 11905 15830 11927 15876
rect 11973 15830 12041 15876
rect 12087 15830 12109 15876
rect 11905 15762 12109 15830
rect 11905 15716 11927 15762
rect 11973 15716 12041 15762
rect 12087 15716 12109 15762
rect 11905 15648 12109 15716
rect 11905 15602 11927 15648
rect 11973 15602 12041 15648
rect 12087 15602 12109 15648
rect 11905 15534 12109 15602
rect 11905 15488 11927 15534
rect 11973 15488 12041 15534
rect 12087 15488 12109 15534
rect 11905 15420 12109 15488
rect 11905 15374 11927 15420
rect 11973 15374 12041 15420
rect 12087 15374 12109 15420
rect 11905 15306 12109 15374
rect 11905 15260 11927 15306
rect 11973 15260 12041 15306
rect 12087 15260 12109 15306
rect 11905 15192 12109 15260
rect 11905 15146 11927 15192
rect 11973 15146 12041 15192
rect 12087 15146 12109 15192
rect 11905 15078 12109 15146
rect 11905 15032 11927 15078
rect 11973 15032 12041 15078
rect 12087 15032 12109 15078
rect 11905 14964 12109 15032
rect 11905 14918 11927 14964
rect 11973 14918 12041 14964
rect 12087 14918 12109 14964
rect 11905 14850 12109 14918
rect 11905 14804 11927 14850
rect 11973 14804 12041 14850
rect 12087 14804 12109 14850
rect 11905 14736 12109 14804
rect 11905 14690 11927 14736
rect 11973 14690 12041 14736
rect 12087 14690 12109 14736
rect 11905 14622 12109 14690
rect 11905 14576 11927 14622
rect 11973 14576 12041 14622
rect 12087 14576 12109 14622
rect 11905 14508 12109 14576
rect 11905 14462 11927 14508
rect 11973 14462 12041 14508
rect 12087 14462 12109 14508
rect 11905 14394 12109 14462
rect 11905 14348 11927 14394
rect 11973 14348 12041 14394
rect 12087 14348 12109 14394
rect 11905 14280 12109 14348
rect 11905 14234 11927 14280
rect 11973 14234 12041 14280
rect 12087 14234 12109 14280
rect 11905 14166 12109 14234
rect 11905 14120 11927 14166
rect 11973 14120 12041 14166
rect 12087 14120 12109 14166
rect 11905 14052 12109 14120
rect 11905 14006 11927 14052
rect 11973 14006 12041 14052
rect 12087 14006 12109 14052
rect 11905 13938 12109 14006
rect 11905 13892 11927 13938
rect 11973 13892 12041 13938
rect 12087 13892 12109 13938
rect 11905 13824 12109 13892
rect 11905 13778 11927 13824
rect 11973 13778 12041 13824
rect 12087 13778 12109 13824
rect 11905 13710 12109 13778
rect 11905 13664 11927 13710
rect 11973 13664 12041 13710
rect 12087 13664 12109 13710
rect 11905 13596 12109 13664
rect 11905 13550 11927 13596
rect 11973 13550 12041 13596
rect 12087 13550 12109 13596
rect 11905 13482 12109 13550
rect 11905 13436 11927 13482
rect 11973 13436 12041 13482
rect 12087 13436 12109 13482
rect 11905 13368 12109 13436
rect 11905 13322 11927 13368
rect 11973 13322 12041 13368
rect 12087 13322 12109 13368
rect 11905 13254 12109 13322
rect 11905 13208 11927 13254
rect 11973 13208 12041 13254
rect 12087 13208 12109 13254
rect 11905 13140 12109 13208
rect 11905 13094 11927 13140
rect 11973 13094 12041 13140
rect 12087 13094 12109 13140
rect 11905 13026 12109 13094
rect 11905 12980 11927 13026
rect 11973 12980 12041 13026
rect 12087 12980 12109 13026
rect 11905 12912 12109 12980
rect 11905 12866 11927 12912
rect 11973 12866 12041 12912
rect 12087 12866 12109 12912
rect 11905 12798 12109 12866
rect 11905 12752 11927 12798
rect 11973 12752 12041 12798
rect 12087 12752 12109 12798
rect 11905 12684 12109 12752
rect 11905 12638 11927 12684
rect 11973 12638 12041 12684
rect 12087 12638 12109 12684
rect 11905 12570 12109 12638
rect 11905 12524 11927 12570
rect 11973 12524 12041 12570
rect 12087 12524 12109 12570
rect 11905 12456 12109 12524
rect 11905 12410 11927 12456
rect 11973 12410 12041 12456
rect 12087 12410 12109 12456
rect 11905 12342 12109 12410
rect 11905 12296 11927 12342
rect 11973 12296 12041 12342
rect 12087 12296 12109 12342
rect 11905 12228 12109 12296
rect 11905 12182 11927 12228
rect 11973 12182 12041 12228
rect 12087 12182 12109 12228
rect 11905 12114 12109 12182
rect 11905 12068 11927 12114
rect 11973 12068 12041 12114
rect 12087 12068 12109 12114
rect 11905 12000 12109 12068
rect 11905 11954 11927 12000
rect 11973 11954 12041 12000
rect 12087 11954 12109 12000
rect 11905 11886 12109 11954
rect 11905 11840 11927 11886
rect 11973 11840 12041 11886
rect 12087 11840 12109 11886
rect 11905 11772 12109 11840
rect 11905 11726 11927 11772
rect 11973 11726 12041 11772
rect 12087 11726 12109 11772
rect 11905 11658 12109 11726
rect 11905 11612 11927 11658
rect 11973 11612 12041 11658
rect 12087 11612 12109 11658
rect 11905 11544 12109 11612
rect 11905 11498 11927 11544
rect 11973 11498 12041 11544
rect 12087 11498 12109 11544
rect 11905 11430 12109 11498
rect 11905 11384 11927 11430
rect 11973 11384 12041 11430
rect 12087 11384 12109 11430
rect 1565 11270 1587 11316
rect 1633 11270 1701 11316
rect 1747 11270 1769 11316
rect 1565 11202 1769 11270
rect 11905 11316 12109 11384
rect 11905 11270 11927 11316
rect 11973 11270 12041 11316
rect 12087 11270 12109 11316
rect 1565 11156 1587 11202
rect 1633 11156 1701 11202
rect 1747 11156 1769 11202
rect 1565 11088 1769 11156
rect 1565 11042 1587 11088
rect 1633 11042 1701 11088
rect 1747 11042 1769 11088
rect 1565 10974 1769 11042
rect 1565 10928 1587 10974
rect 1633 10928 1701 10974
rect 1747 10947 1769 10974
rect 11905 11202 12109 11270
rect 11905 11156 11927 11202
rect 11973 11156 12041 11202
rect 12087 11156 12109 11202
rect 11905 11088 12109 11156
rect 11905 11042 11927 11088
rect 11973 11042 12041 11088
rect 12087 11042 12109 11088
rect 11905 10974 12109 11042
rect 11905 10947 11927 10974
rect 1747 10928 11927 10947
rect 11973 10928 12041 10974
rect 12087 10928 12109 10974
rect 1565 10925 12109 10928
rect 1565 10879 1855 10925
rect 1901 10879 1969 10925
rect 2015 10879 2083 10925
rect 2129 10879 2197 10925
rect 2243 10879 2311 10925
rect 2357 10879 2425 10925
rect 2471 10879 2539 10925
rect 2585 10879 2653 10925
rect 2699 10879 2767 10925
rect 2813 10879 2881 10925
rect 2927 10879 2995 10925
rect 3041 10879 3109 10925
rect 3155 10879 3223 10925
rect 3269 10879 3337 10925
rect 3383 10879 3451 10925
rect 3497 10879 3565 10925
rect 3611 10879 3679 10925
rect 3725 10879 3793 10925
rect 3839 10879 3907 10925
rect 3953 10879 4021 10925
rect 4067 10879 4135 10925
rect 4181 10879 4249 10925
rect 4295 10879 4363 10925
rect 4409 10879 4477 10925
rect 4523 10879 4591 10925
rect 4637 10879 4705 10925
rect 4751 10879 4819 10925
rect 4865 10879 4933 10925
rect 4979 10879 5047 10925
rect 5093 10879 5161 10925
rect 5207 10879 5275 10925
rect 5321 10879 5389 10925
rect 5435 10879 5503 10925
rect 5549 10879 5617 10925
rect 5663 10879 5731 10925
rect 5777 10879 5845 10925
rect 5891 10879 5959 10925
rect 6005 10879 6073 10925
rect 6119 10879 6187 10925
rect 6233 10879 6301 10925
rect 6347 10879 6415 10925
rect 6461 10879 6529 10925
rect 6575 10879 6643 10925
rect 6689 10879 6757 10925
rect 6803 10879 6871 10925
rect 6917 10879 6985 10925
rect 7031 10879 7099 10925
rect 7145 10879 7213 10925
rect 7259 10879 7327 10925
rect 7373 10879 7441 10925
rect 7487 10879 7555 10925
rect 7601 10879 7669 10925
rect 7715 10879 7783 10925
rect 7829 10879 7897 10925
rect 7943 10879 8011 10925
rect 8057 10879 8125 10925
rect 8171 10879 8239 10925
rect 8285 10879 8353 10925
rect 8399 10879 8467 10925
rect 8513 10879 8581 10925
rect 8627 10879 8695 10925
rect 8741 10879 8809 10925
rect 8855 10879 8923 10925
rect 8969 10879 9037 10925
rect 9083 10879 9151 10925
rect 9197 10879 9265 10925
rect 9311 10879 9379 10925
rect 9425 10879 9493 10925
rect 9539 10879 9607 10925
rect 9653 10879 9721 10925
rect 9767 10879 9835 10925
rect 9881 10879 9949 10925
rect 9995 10879 10063 10925
rect 10109 10879 10177 10925
rect 10223 10879 10291 10925
rect 10337 10879 10405 10925
rect 10451 10879 10519 10925
rect 10565 10879 10633 10925
rect 10679 10879 10747 10925
rect 10793 10879 10861 10925
rect 10907 10879 10975 10925
rect 11021 10879 11089 10925
rect 11135 10879 11203 10925
rect 11249 10879 11317 10925
rect 11363 10879 11431 10925
rect 11477 10879 11545 10925
rect 11591 10879 11659 10925
rect 11705 10879 11773 10925
rect 11819 10879 12109 10925
rect 1565 10860 12109 10879
rect 1565 10814 1587 10860
rect 1633 10814 1701 10860
rect 1747 10814 11927 10860
rect 11973 10814 12041 10860
rect 12087 10814 12109 10860
rect 1565 10811 12109 10814
rect 1565 10765 1855 10811
rect 1901 10765 1969 10811
rect 2015 10765 2083 10811
rect 2129 10765 2197 10811
rect 2243 10765 2311 10811
rect 2357 10765 2425 10811
rect 2471 10765 2539 10811
rect 2585 10765 2653 10811
rect 2699 10765 2767 10811
rect 2813 10765 2881 10811
rect 2927 10765 2995 10811
rect 3041 10765 3109 10811
rect 3155 10765 3223 10811
rect 3269 10765 3337 10811
rect 3383 10765 3451 10811
rect 3497 10765 3565 10811
rect 3611 10765 3679 10811
rect 3725 10765 3793 10811
rect 3839 10765 3907 10811
rect 3953 10765 4021 10811
rect 4067 10765 4135 10811
rect 4181 10765 4249 10811
rect 4295 10765 4363 10811
rect 4409 10765 4477 10811
rect 4523 10765 4591 10811
rect 4637 10765 4705 10811
rect 4751 10765 4819 10811
rect 4865 10765 4933 10811
rect 4979 10765 5047 10811
rect 5093 10765 5161 10811
rect 5207 10765 5275 10811
rect 5321 10765 5389 10811
rect 5435 10765 5503 10811
rect 5549 10765 5617 10811
rect 5663 10765 5731 10811
rect 5777 10765 5845 10811
rect 5891 10765 5959 10811
rect 6005 10765 6073 10811
rect 6119 10765 6187 10811
rect 6233 10765 6301 10811
rect 6347 10765 6415 10811
rect 6461 10765 6529 10811
rect 6575 10765 6643 10811
rect 6689 10765 6757 10811
rect 6803 10765 6871 10811
rect 6917 10765 6985 10811
rect 7031 10765 7099 10811
rect 7145 10765 7213 10811
rect 7259 10765 7327 10811
rect 7373 10765 7441 10811
rect 7487 10765 7555 10811
rect 7601 10765 7669 10811
rect 7715 10765 7783 10811
rect 7829 10765 7897 10811
rect 7943 10765 8011 10811
rect 8057 10765 8125 10811
rect 8171 10765 8239 10811
rect 8285 10765 8353 10811
rect 8399 10765 8467 10811
rect 8513 10765 8581 10811
rect 8627 10765 8695 10811
rect 8741 10765 8809 10811
rect 8855 10765 8923 10811
rect 8969 10765 9037 10811
rect 9083 10765 9151 10811
rect 9197 10765 9265 10811
rect 9311 10765 9379 10811
rect 9425 10765 9493 10811
rect 9539 10765 9607 10811
rect 9653 10765 9721 10811
rect 9767 10765 9835 10811
rect 9881 10765 9949 10811
rect 9995 10765 10063 10811
rect 10109 10765 10177 10811
rect 10223 10765 10291 10811
rect 10337 10765 10405 10811
rect 10451 10765 10519 10811
rect 10565 10765 10633 10811
rect 10679 10765 10747 10811
rect 10793 10765 10861 10811
rect 10907 10765 10975 10811
rect 11021 10765 11089 10811
rect 11135 10765 11203 10811
rect 11249 10765 11317 10811
rect 11363 10765 11431 10811
rect 11477 10765 11545 10811
rect 11591 10765 11659 10811
rect 11705 10765 11773 10811
rect 11819 10765 12109 10811
rect 1565 10746 12109 10765
rect 1565 10700 1587 10746
rect 1633 10700 1701 10746
rect 1747 10743 11927 10746
rect 1747 10700 1769 10743
rect 1565 10632 1769 10700
rect 1565 10586 1587 10632
rect 1633 10586 1701 10632
rect 1747 10586 1769 10632
rect 1565 10518 1769 10586
rect 1565 10472 1587 10518
rect 1633 10472 1701 10518
rect 1747 10472 1769 10518
rect 1565 10404 1769 10472
rect 11905 10700 11927 10743
rect 11973 10700 12041 10746
rect 12087 10700 12109 10746
rect 11905 10632 12109 10700
rect 11905 10586 11927 10632
rect 11973 10586 12041 10632
rect 12087 10586 12109 10632
rect 11905 10518 12109 10586
rect 11905 10472 11927 10518
rect 11973 10472 12041 10518
rect 12087 10472 12109 10518
rect 1565 10358 1587 10404
rect 1633 10358 1701 10404
rect 1747 10358 1769 10404
rect 1565 10290 1769 10358
rect 11905 10404 12109 10472
rect 11905 10358 11927 10404
rect 11973 10358 12041 10404
rect 12087 10358 12109 10404
rect 1565 10244 1587 10290
rect 1633 10244 1701 10290
rect 1747 10244 1769 10290
rect 1565 10176 1769 10244
rect 1565 10130 1587 10176
rect 1633 10130 1701 10176
rect 1747 10130 1769 10176
rect 1565 10062 1769 10130
rect 1565 10016 1587 10062
rect 1633 10016 1701 10062
rect 1747 10016 1769 10062
rect 1565 9948 1769 10016
rect 1565 9902 1587 9948
rect 1633 9902 1701 9948
rect 1747 9902 1769 9948
rect 1565 9834 1769 9902
rect 1565 9788 1587 9834
rect 1633 9788 1701 9834
rect 1747 9788 1769 9834
rect 1565 9720 1769 9788
rect 1565 9674 1587 9720
rect 1633 9674 1701 9720
rect 1747 9674 1769 9720
rect 1565 9606 1769 9674
rect 1565 9560 1587 9606
rect 1633 9560 1701 9606
rect 1747 9560 1769 9606
rect 1565 9492 1769 9560
rect 1565 9446 1587 9492
rect 1633 9446 1701 9492
rect 1747 9446 1769 9492
rect 1565 9378 1769 9446
rect 1565 9332 1587 9378
rect 1633 9332 1701 9378
rect 1747 9332 1769 9378
rect 1565 9264 1769 9332
rect 1565 9218 1587 9264
rect 1633 9218 1701 9264
rect 1747 9218 1769 9264
rect 1565 9150 1769 9218
rect 1565 9104 1587 9150
rect 1633 9104 1701 9150
rect 1747 9104 1769 9150
rect 1565 9036 1769 9104
rect 1565 8990 1587 9036
rect 1633 8990 1701 9036
rect 1747 8990 1769 9036
rect 1565 8922 1769 8990
rect 1565 8876 1587 8922
rect 1633 8876 1701 8922
rect 1747 8876 1769 8922
rect 1565 8808 1769 8876
rect 1565 8762 1587 8808
rect 1633 8762 1701 8808
rect 1747 8762 1769 8808
rect 1565 8694 1769 8762
rect 1565 8648 1587 8694
rect 1633 8648 1701 8694
rect 1747 8648 1769 8694
rect 1565 8580 1769 8648
rect 1565 8534 1587 8580
rect 1633 8534 1701 8580
rect 1747 8534 1769 8580
rect 1565 8466 1769 8534
rect 1565 8420 1587 8466
rect 1633 8420 1701 8466
rect 1747 8420 1769 8466
rect 1565 8352 1769 8420
rect 1565 8306 1587 8352
rect 1633 8306 1701 8352
rect 1747 8306 1769 8352
rect 1565 8238 1769 8306
rect 1565 8192 1587 8238
rect 1633 8192 1701 8238
rect 1747 8192 1769 8238
rect 1565 8124 1769 8192
rect 1565 8078 1587 8124
rect 1633 8078 1701 8124
rect 1747 8078 1769 8124
rect 1565 8010 1769 8078
rect 1565 7964 1587 8010
rect 1633 7964 1701 8010
rect 1747 7964 1769 8010
rect 1565 7896 1769 7964
rect 1565 7850 1587 7896
rect 1633 7850 1701 7896
rect 1747 7850 1769 7896
rect 1565 7782 1769 7850
rect 1565 7736 1587 7782
rect 1633 7736 1701 7782
rect 1747 7736 1769 7782
rect 1565 7668 1769 7736
rect 1565 7622 1587 7668
rect 1633 7622 1701 7668
rect 1747 7622 1769 7668
rect 1565 7554 1769 7622
rect 1565 7508 1587 7554
rect 1633 7508 1701 7554
rect 1747 7508 1769 7554
rect 1565 7440 1769 7508
rect 1565 7394 1587 7440
rect 1633 7394 1701 7440
rect 1747 7394 1769 7440
rect 1565 7326 1769 7394
rect 1565 7280 1587 7326
rect 1633 7280 1701 7326
rect 1747 7280 1769 7326
rect 1565 7212 1769 7280
rect 1565 7166 1587 7212
rect 1633 7166 1701 7212
rect 1747 7166 1769 7212
rect 1565 7098 1769 7166
rect 1565 7052 1587 7098
rect 1633 7052 1701 7098
rect 1747 7052 1769 7098
rect 1565 6984 1769 7052
rect 1565 6938 1587 6984
rect 1633 6938 1701 6984
rect 1747 6938 1769 6984
rect 1565 6870 1769 6938
rect 1565 6824 1587 6870
rect 1633 6824 1701 6870
rect 1747 6824 1769 6870
rect 1565 6756 1769 6824
rect 1565 6710 1587 6756
rect 1633 6710 1701 6756
rect 1747 6710 1769 6756
rect 1565 6642 1769 6710
rect 1565 6596 1587 6642
rect 1633 6596 1701 6642
rect 1747 6596 1769 6642
rect 1565 6528 1769 6596
rect 1565 6482 1587 6528
rect 1633 6482 1701 6528
rect 1747 6482 1769 6528
rect 1565 6414 1769 6482
rect 1565 6368 1587 6414
rect 1633 6368 1701 6414
rect 1747 6368 1769 6414
rect 1565 6300 1769 6368
rect 1565 6254 1587 6300
rect 1633 6254 1701 6300
rect 1747 6254 1769 6300
rect 1565 6186 1769 6254
rect 1565 6140 1587 6186
rect 1633 6140 1701 6186
rect 1747 6140 1769 6186
rect 1565 6072 1769 6140
rect 1565 6026 1587 6072
rect 1633 6026 1701 6072
rect 1747 6026 1769 6072
rect 1565 5958 1769 6026
rect 1565 5912 1587 5958
rect 1633 5912 1701 5958
rect 1747 5912 1769 5958
rect 1565 5844 1769 5912
rect 1565 5798 1587 5844
rect 1633 5798 1701 5844
rect 1747 5798 1769 5844
rect 1565 5730 1769 5798
rect 1565 5684 1587 5730
rect 1633 5684 1701 5730
rect 1747 5684 1769 5730
rect 1565 5616 1769 5684
rect 1565 5570 1587 5616
rect 1633 5570 1701 5616
rect 1747 5570 1769 5616
rect 1565 5502 1769 5570
rect 1565 5456 1587 5502
rect 1633 5456 1701 5502
rect 1747 5456 1769 5502
rect 1565 5046 1769 5456
rect 11905 10290 12109 10358
rect 11905 10244 11927 10290
rect 11973 10244 12041 10290
rect 12087 10244 12109 10290
rect 11905 10176 12109 10244
rect 11905 10130 11927 10176
rect 11973 10130 12041 10176
rect 12087 10130 12109 10176
rect 11905 10062 12109 10130
rect 11905 10016 11927 10062
rect 11973 10016 12041 10062
rect 12087 10016 12109 10062
rect 11905 9948 12109 10016
rect 11905 9902 11927 9948
rect 11973 9902 12041 9948
rect 12087 9902 12109 9948
rect 11905 9834 12109 9902
rect 11905 9788 11927 9834
rect 11973 9788 12041 9834
rect 12087 9788 12109 9834
rect 11905 9720 12109 9788
rect 11905 9674 11927 9720
rect 11973 9674 12041 9720
rect 12087 9674 12109 9720
rect 11905 9606 12109 9674
rect 11905 9560 11927 9606
rect 11973 9560 12041 9606
rect 12087 9560 12109 9606
rect 11905 9492 12109 9560
rect 11905 9446 11927 9492
rect 11973 9446 12041 9492
rect 12087 9446 12109 9492
rect 11905 9378 12109 9446
rect 11905 9332 11927 9378
rect 11973 9332 12041 9378
rect 12087 9332 12109 9378
rect 11905 9264 12109 9332
rect 11905 9218 11927 9264
rect 11973 9218 12041 9264
rect 12087 9218 12109 9264
rect 11905 9150 12109 9218
rect 11905 9104 11927 9150
rect 11973 9104 12041 9150
rect 12087 9104 12109 9150
rect 11905 9036 12109 9104
rect 11905 8990 11927 9036
rect 11973 8990 12041 9036
rect 12087 8990 12109 9036
rect 11905 8922 12109 8990
rect 11905 8876 11927 8922
rect 11973 8876 12041 8922
rect 12087 8876 12109 8922
rect 11905 8808 12109 8876
rect 11905 8762 11927 8808
rect 11973 8762 12041 8808
rect 12087 8762 12109 8808
rect 11905 8694 12109 8762
rect 11905 8648 11927 8694
rect 11973 8648 12041 8694
rect 12087 8648 12109 8694
rect 11905 8580 12109 8648
rect 11905 8534 11927 8580
rect 11973 8534 12041 8580
rect 12087 8534 12109 8580
rect 11905 8466 12109 8534
rect 11905 8420 11927 8466
rect 11973 8420 12041 8466
rect 12087 8420 12109 8466
rect 11905 8352 12109 8420
rect 11905 8306 11927 8352
rect 11973 8306 12041 8352
rect 12087 8306 12109 8352
rect 11905 8238 12109 8306
rect 11905 8192 11927 8238
rect 11973 8192 12041 8238
rect 12087 8192 12109 8238
rect 11905 8124 12109 8192
rect 11905 8078 11927 8124
rect 11973 8078 12041 8124
rect 12087 8078 12109 8124
rect 11905 8010 12109 8078
rect 11905 7964 11927 8010
rect 11973 7964 12041 8010
rect 12087 7964 12109 8010
rect 11905 7896 12109 7964
rect 11905 7850 11927 7896
rect 11973 7850 12041 7896
rect 12087 7850 12109 7896
rect 11905 7782 12109 7850
rect 11905 7736 11927 7782
rect 11973 7736 12041 7782
rect 12087 7736 12109 7782
rect 11905 7668 12109 7736
rect 11905 7622 11927 7668
rect 11973 7622 12041 7668
rect 12087 7622 12109 7668
rect 11905 7554 12109 7622
rect 11905 7508 11927 7554
rect 11973 7508 12041 7554
rect 12087 7508 12109 7554
rect 11905 7440 12109 7508
rect 11905 7394 11927 7440
rect 11973 7394 12041 7440
rect 12087 7394 12109 7440
rect 11905 7326 12109 7394
rect 11905 7280 11927 7326
rect 11973 7280 12041 7326
rect 12087 7280 12109 7326
rect 11905 7212 12109 7280
rect 11905 7166 11927 7212
rect 11973 7166 12041 7212
rect 12087 7166 12109 7212
rect 11905 7098 12109 7166
rect 11905 7052 11927 7098
rect 11973 7052 12041 7098
rect 12087 7052 12109 7098
rect 11905 6984 12109 7052
rect 11905 6938 11927 6984
rect 11973 6938 12041 6984
rect 12087 6938 12109 6984
rect 11905 6870 12109 6938
rect 11905 6824 11927 6870
rect 11973 6824 12041 6870
rect 12087 6824 12109 6870
rect 11905 6756 12109 6824
rect 11905 6710 11927 6756
rect 11973 6710 12041 6756
rect 12087 6710 12109 6756
rect 11905 6642 12109 6710
rect 11905 6596 11927 6642
rect 11973 6596 12041 6642
rect 12087 6596 12109 6642
rect 11905 6528 12109 6596
rect 11905 6482 11927 6528
rect 11973 6482 12041 6528
rect 12087 6482 12109 6528
rect 11905 6414 12109 6482
rect 11905 6368 11927 6414
rect 11973 6368 12041 6414
rect 12087 6368 12109 6414
rect 11905 6300 12109 6368
rect 11905 6254 11927 6300
rect 11973 6254 12041 6300
rect 12087 6254 12109 6300
rect 11905 6186 12109 6254
rect 11905 6140 11927 6186
rect 11973 6140 12041 6186
rect 12087 6140 12109 6186
rect 11905 6072 12109 6140
rect 11905 6026 11927 6072
rect 11973 6026 12041 6072
rect 12087 6026 12109 6072
rect 11905 5958 12109 6026
rect 11905 5912 11927 5958
rect 11973 5912 12041 5958
rect 12087 5912 12109 5958
rect 11905 5844 12109 5912
rect 11905 5798 11927 5844
rect 11973 5798 12041 5844
rect 12087 5798 12109 5844
rect 11905 5730 12109 5798
rect 11905 5684 11927 5730
rect 11973 5684 12041 5730
rect 12087 5684 12109 5730
rect 11905 5616 12109 5684
rect 11905 5570 11927 5616
rect 11973 5570 12041 5616
rect 12087 5570 12109 5616
rect 11905 5502 12109 5570
rect 11905 5456 11927 5502
rect 11973 5456 12041 5502
rect 12087 5456 12109 5502
rect 11905 5388 12109 5456
rect 11905 5342 11927 5388
rect 11973 5342 12041 5388
rect 12087 5342 12109 5388
rect 11905 5274 12109 5342
rect 1565 5000 1587 5046
rect 1633 5000 1701 5046
rect 1747 5000 1769 5046
rect 1565 4954 1769 5000
rect 11905 5228 11927 5274
rect 11973 5228 12041 5274
rect 12087 5228 12109 5274
rect 11905 5160 12109 5228
rect 11905 5114 11927 5160
rect 11973 5114 12041 5160
rect 12087 5114 12109 5160
rect 11905 5046 12109 5114
rect 11905 5000 11927 5046
rect 11973 5000 12041 5046
rect 12087 5000 12109 5046
rect 11905 4954 12109 5000
rect 1565 4932 12109 4954
rect 1565 4886 1587 4932
rect 1633 4886 1701 4932
rect 1747 4886 1855 4932
rect 1901 4886 1969 4932
rect 2015 4886 2083 4932
rect 2129 4886 2197 4932
rect 2243 4886 2311 4932
rect 2357 4886 2425 4932
rect 2471 4886 2539 4932
rect 2585 4886 2653 4932
rect 2699 4886 2767 4932
rect 2813 4886 2881 4932
rect 2927 4886 2995 4932
rect 3041 4886 3109 4932
rect 3155 4886 3223 4932
rect 3269 4886 3337 4932
rect 3383 4886 3451 4932
rect 3497 4886 3565 4932
rect 3611 4886 3679 4932
rect 3725 4886 3793 4932
rect 3839 4886 3907 4932
rect 3953 4886 4021 4932
rect 4067 4886 4135 4932
rect 4181 4886 4249 4932
rect 4295 4886 4363 4932
rect 4409 4886 4477 4932
rect 4523 4886 4591 4932
rect 4637 4886 4705 4932
rect 4751 4886 4819 4932
rect 4865 4886 4933 4932
rect 4979 4886 5047 4932
rect 5093 4886 5161 4932
rect 5207 4886 5275 4932
rect 5321 4886 5389 4932
rect 5435 4886 5503 4932
rect 5549 4886 5617 4932
rect 5663 4886 5731 4932
rect 5777 4886 5845 4932
rect 5891 4886 5959 4932
rect 6005 4886 6073 4932
rect 6119 4886 6187 4932
rect 6233 4886 6301 4932
rect 6347 4886 6415 4932
rect 6461 4886 6529 4932
rect 6575 4886 6643 4932
rect 6689 4886 6757 4932
rect 6803 4886 6871 4932
rect 6917 4886 6985 4932
rect 7031 4886 7099 4932
rect 7145 4886 7213 4932
rect 7259 4886 7327 4932
rect 7373 4886 7441 4932
rect 7487 4886 7555 4932
rect 7601 4886 7669 4932
rect 7715 4886 7783 4932
rect 7829 4886 7897 4932
rect 7943 4886 8011 4932
rect 8057 4886 8125 4932
rect 8171 4886 8239 4932
rect 8285 4886 8353 4932
rect 8399 4886 8467 4932
rect 8513 4886 8581 4932
rect 8627 4886 8695 4932
rect 8741 4886 8809 4932
rect 8855 4886 8923 4932
rect 8969 4886 9037 4932
rect 9083 4886 9151 4932
rect 9197 4886 9265 4932
rect 9311 4886 9379 4932
rect 9425 4886 9493 4932
rect 9539 4886 9607 4932
rect 9653 4886 9721 4932
rect 9767 4886 9835 4932
rect 9881 4886 9949 4932
rect 9995 4886 10063 4932
rect 10109 4886 10177 4932
rect 10223 4886 10291 4932
rect 10337 4886 10405 4932
rect 10451 4886 10519 4932
rect 10565 4886 10633 4932
rect 10679 4886 10747 4932
rect 10793 4886 10861 4932
rect 10907 4886 10975 4932
rect 11021 4886 11089 4932
rect 11135 4886 11203 4932
rect 11249 4886 11317 4932
rect 11363 4886 11431 4932
rect 11477 4886 11545 4932
rect 11591 4886 11659 4932
rect 11705 4886 11773 4932
rect 11819 4886 11927 4932
rect 11973 4886 12041 4932
rect 12087 4886 12109 4932
rect 1565 4818 12109 4886
rect 1565 4772 1587 4818
rect 1633 4772 1701 4818
rect 1747 4772 1855 4818
rect 1901 4772 1969 4818
rect 2015 4772 2083 4818
rect 2129 4772 2197 4818
rect 2243 4772 2311 4818
rect 2357 4772 2425 4818
rect 2471 4772 2539 4818
rect 2585 4772 2653 4818
rect 2699 4772 2767 4818
rect 2813 4772 2881 4818
rect 2927 4772 2995 4818
rect 3041 4772 3109 4818
rect 3155 4772 3223 4818
rect 3269 4772 3337 4818
rect 3383 4772 3451 4818
rect 3497 4772 3565 4818
rect 3611 4772 3679 4818
rect 3725 4772 3793 4818
rect 3839 4772 3907 4818
rect 3953 4772 4021 4818
rect 4067 4772 4135 4818
rect 4181 4772 4249 4818
rect 4295 4772 4363 4818
rect 4409 4772 4477 4818
rect 4523 4772 4591 4818
rect 4637 4772 4705 4818
rect 4751 4772 4819 4818
rect 4865 4772 4933 4818
rect 4979 4772 5047 4818
rect 5093 4772 5161 4818
rect 5207 4772 5275 4818
rect 5321 4772 5389 4818
rect 5435 4772 5503 4818
rect 5549 4772 5617 4818
rect 5663 4772 5731 4818
rect 5777 4772 5845 4818
rect 5891 4772 5959 4818
rect 6005 4772 6073 4818
rect 6119 4772 6187 4818
rect 6233 4772 6301 4818
rect 6347 4772 6415 4818
rect 6461 4772 6529 4818
rect 6575 4772 6643 4818
rect 6689 4772 6757 4818
rect 6803 4772 6871 4818
rect 6917 4772 6985 4818
rect 7031 4772 7099 4818
rect 7145 4772 7213 4818
rect 7259 4772 7327 4818
rect 7373 4772 7441 4818
rect 7487 4772 7555 4818
rect 7601 4772 7669 4818
rect 7715 4772 7783 4818
rect 7829 4772 7897 4818
rect 7943 4772 8011 4818
rect 8057 4772 8125 4818
rect 8171 4772 8239 4818
rect 8285 4772 8353 4818
rect 8399 4772 8467 4818
rect 8513 4772 8581 4818
rect 8627 4772 8695 4818
rect 8741 4772 8809 4818
rect 8855 4772 8923 4818
rect 8969 4772 9037 4818
rect 9083 4772 9151 4818
rect 9197 4772 9265 4818
rect 9311 4772 9379 4818
rect 9425 4772 9493 4818
rect 9539 4772 9607 4818
rect 9653 4772 9721 4818
rect 9767 4772 9835 4818
rect 9881 4772 9949 4818
rect 9995 4772 10063 4818
rect 10109 4772 10177 4818
rect 10223 4772 10291 4818
rect 10337 4772 10405 4818
rect 10451 4772 10519 4818
rect 10565 4772 10633 4818
rect 10679 4772 10747 4818
rect 10793 4772 10861 4818
rect 10907 4772 10975 4818
rect 11021 4772 11089 4818
rect 11135 4772 11203 4818
rect 11249 4772 11317 4818
rect 11363 4772 11431 4818
rect 11477 4772 11545 4818
rect 11591 4772 11659 4818
rect 11705 4772 11773 4818
rect 11819 4772 11927 4818
rect 11973 4772 12041 4818
rect 12087 4772 12109 4818
rect 1565 4750 12109 4772
<< nsubdiff >>
rect -3749 17592 81 17614
rect -3749 17546 -3727 17592
rect -3681 17546 -3573 17592
rect -3527 17546 -3469 17592
rect -3423 17546 -3365 17592
rect -3319 17546 -3261 17592
rect -3215 17546 -3157 17592
rect -3111 17546 -3053 17592
rect -3007 17546 -2949 17592
rect -2903 17546 -2845 17592
rect -2799 17546 -2741 17592
rect -2695 17546 -2637 17592
rect -2591 17546 -2533 17592
rect -2487 17546 -2429 17592
rect -2383 17546 -2325 17592
rect -2279 17546 -2221 17592
rect -2175 17546 -2117 17592
rect -2071 17546 -2013 17592
rect -1967 17546 -1909 17592
rect -1863 17546 -1805 17592
rect -1759 17546 -1701 17592
rect -1655 17546 -1597 17592
rect -1551 17546 -1493 17592
rect -1447 17546 -1389 17592
rect -1343 17546 -1285 17592
rect -1239 17546 -1181 17592
rect -1135 17546 -1077 17592
rect -1031 17546 -973 17592
rect -927 17546 -869 17592
rect -823 17546 -765 17592
rect -719 17546 -661 17592
rect -615 17546 -557 17592
rect -511 17546 -453 17592
rect -407 17546 -349 17592
rect -303 17546 -245 17592
rect -199 17546 -141 17592
rect -95 17546 13 17592
rect 59 17546 81 17592
rect -3749 17524 81 17546
rect -3749 17488 -3659 17524
rect -3749 17442 -3727 17488
rect -3681 17442 -3659 17488
rect -3749 17384 -3659 17442
rect -3749 17338 -3727 17384
rect -3681 17338 -3659 17384
rect -3749 17280 -3659 17338
rect -9 17488 81 17524
rect -9 17442 13 17488
rect 59 17442 81 17488
rect -9 17384 81 17442
rect -9 17338 13 17384
rect 59 17338 81 17384
rect -3749 17234 -3727 17280
rect -3681 17234 -3659 17280
rect -3749 17176 -3659 17234
rect -3749 17130 -3727 17176
rect -3681 17130 -3659 17176
rect -3749 17072 -3659 17130
rect -3749 17026 -3727 17072
rect -3681 17026 -3659 17072
rect -3749 16968 -3659 17026
rect -3749 16922 -3727 16968
rect -3681 16922 -3659 16968
rect -3749 16864 -3659 16922
rect -3749 16818 -3727 16864
rect -3681 16818 -3659 16864
rect -3749 16760 -3659 16818
rect -3749 16714 -3727 16760
rect -3681 16714 -3659 16760
rect -3749 16656 -3659 16714
rect -3749 16610 -3727 16656
rect -3681 16610 -3659 16656
rect -3749 16552 -3659 16610
rect -3749 16506 -3727 16552
rect -3681 16506 -3659 16552
rect -3749 16448 -3659 16506
rect -3749 16402 -3727 16448
rect -3681 16402 -3659 16448
rect -3749 16344 -3659 16402
rect -3749 16298 -3727 16344
rect -3681 16298 -3659 16344
rect -3749 16240 -3659 16298
rect -3749 16194 -3727 16240
rect -3681 16194 -3659 16240
rect -3749 16136 -3659 16194
rect -3749 16090 -3727 16136
rect -3681 16090 -3659 16136
rect -3749 16032 -3659 16090
rect -3749 15986 -3727 16032
rect -3681 15986 -3659 16032
rect -3749 15928 -3659 15986
rect -3749 15882 -3727 15928
rect -3681 15882 -3659 15928
rect -3749 15824 -3659 15882
rect -3749 15778 -3727 15824
rect -3681 15778 -3659 15824
rect -3749 15720 -3659 15778
rect -3749 15674 -3727 15720
rect -3681 15674 -3659 15720
rect -3749 15616 -3659 15674
rect -3749 15570 -3727 15616
rect -3681 15570 -3659 15616
rect -3749 15512 -3659 15570
rect -3749 15466 -3727 15512
rect -3681 15466 -3659 15512
rect -3749 15408 -3659 15466
rect -3749 15362 -3727 15408
rect -3681 15362 -3659 15408
rect -3749 15304 -3659 15362
rect -3749 15258 -3727 15304
rect -3681 15258 -3659 15304
rect -3749 15200 -3659 15258
rect -3749 15154 -3727 15200
rect -3681 15154 -3659 15200
rect -3749 15096 -3659 15154
rect -3749 15050 -3727 15096
rect -3681 15050 -3659 15096
rect -3749 14992 -3659 15050
rect -3749 14946 -3727 14992
rect -3681 14946 -3659 14992
rect -3749 14888 -3659 14946
rect -3749 14842 -3727 14888
rect -3681 14842 -3659 14888
rect -3749 14784 -3659 14842
rect -3749 14738 -3727 14784
rect -3681 14738 -3659 14784
rect -3749 14680 -3659 14738
rect -3749 14634 -3727 14680
rect -3681 14634 -3659 14680
rect -3749 14576 -3659 14634
rect -3749 14530 -3727 14576
rect -3681 14530 -3659 14576
rect -3749 14472 -3659 14530
rect -3749 14426 -3727 14472
rect -3681 14426 -3659 14472
rect -3749 14368 -3659 14426
rect -3749 14322 -3727 14368
rect -3681 14322 -3659 14368
rect -3749 14264 -3659 14322
rect -3749 14218 -3727 14264
rect -3681 14218 -3659 14264
rect -3749 14160 -3659 14218
rect -3749 14114 -3727 14160
rect -3681 14114 -3659 14160
rect -3749 14056 -3659 14114
rect -3749 14010 -3727 14056
rect -3681 14010 -3659 14056
rect -3749 13952 -3659 14010
rect -3749 13906 -3727 13952
rect -3681 13906 -3659 13952
rect -3749 13848 -3659 13906
rect -3749 13802 -3727 13848
rect -3681 13802 -3659 13848
rect -3749 13744 -3659 13802
rect -3749 13698 -3727 13744
rect -3681 13698 -3659 13744
rect -3749 13640 -3659 13698
rect -3749 13594 -3727 13640
rect -3681 13594 -3659 13640
rect -3749 13536 -3659 13594
rect -3749 13490 -3727 13536
rect -3681 13490 -3659 13536
rect -3749 13432 -3659 13490
rect -3749 13386 -3727 13432
rect -3681 13386 -3659 13432
rect -3749 13328 -3659 13386
rect -3749 13282 -3727 13328
rect -3681 13282 -3659 13328
rect -3749 13224 -3659 13282
rect -3749 13178 -3727 13224
rect -3681 13178 -3659 13224
rect -3749 13120 -3659 13178
rect -3749 13074 -3727 13120
rect -3681 13074 -3659 13120
rect -3749 13016 -3659 13074
rect -3749 12970 -3727 13016
rect -3681 12970 -3659 13016
rect -3749 12912 -3659 12970
rect -3749 12866 -3727 12912
rect -3681 12866 -3659 12912
rect -3749 12808 -3659 12866
rect -3749 12762 -3727 12808
rect -3681 12762 -3659 12808
rect -3749 12704 -3659 12762
rect -3749 12658 -3727 12704
rect -3681 12658 -3659 12704
rect -3749 12600 -3659 12658
rect -3749 12554 -3727 12600
rect -3681 12554 -3659 12600
rect -3749 12496 -3659 12554
rect -3749 12450 -3727 12496
rect -3681 12450 -3659 12496
rect -3749 12392 -3659 12450
rect -3749 12346 -3727 12392
rect -3681 12346 -3659 12392
rect -3749 12288 -3659 12346
rect -3749 12242 -3727 12288
rect -3681 12242 -3659 12288
rect -3749 12184 -3659 12242
rect -3749 12138 -3727 12184
rect -3681 12138 -3659 12184
rect -3749 12080 -3659 12138
rect -3749 12034 -3727 12080
rect -3681 12034 -3659 12080
rect -3749 11976 -3659 12034
rect -3749 11930 -3727 11976
rect -3681 11930 -3659 11976
rect -3749 11872 -3659 11930
rect -3749 11826 -3727 11872
rect -3681 11826 -3659 11872
rect -3749 11768 -3659 11826
rect -3749 11722 -3727 11768
rect -3681 11722 -3659 11768
rect -3749 11664 -3659 11722
rect -3749 11618 -3727 11664
rect -3681 11618 -3659 11664
rect -3749 11560 -3659 11618
rect -3749 11514 -3727 11560
rect -3681 11514 -3659 11560
rect -3749 11456 -3659 11514
rect -3749 11410 -3727 11456
rect -3681 11410 -3659 11456
rect -3749 11352 -3659 11410
rect -3749 11306 -3727 11352
rect -3681 11306 -3659 11352
rect -3749 11248 -3659 11306
rect -3749 11202 -3727 11248
rect -3681 11202 -3659 11248
rect -3749 11144 -3659 11202
rect -3749 11098 -3727 11144
rect -3681 11098 -3659 11144
rect -3749 11040 -3659 11098
rect -3749 10994 -3727 11040
rect -3681 10994 -3659 11040
rect -3749 10936 -3659 10994
rect -3749 10890 -3727 10936
rect -3681 10890 -3659 10936
rect -3749 10832 -3659 10890
rect -3749 10786 -3727 10832
rect -3681 10786 -3659 10832
rect -3749 10728 -3659 10786
rect -3749 10682 -3727 10728
rect -3681 10682 -3659 10728
rect -3749 10624 -3659 10682
rect -3749 10578 -3727 10624
rect -3681 10578 -3659 10624
rect -3749 10520 -3659 10578
rect -3749 10474 -3727 10520
rect -3681 10474 -3659 10520
rect -3749 10416 -3659 10474
rect -3749 10370 -3727 10416
rect -3681 10370 -3659 10416
rect -3749 10312 -3659 10370
rect -3749 10266 -3727 10312
rect -3681 10266 -3659 10312
rect -3749 10208 -3659 10266
rect -3749 10162 -3727 10208
rect -3681 10162 -3659 10208
rect -3749 10104 -3659 10162
rect -3749 10058 -3727 10104
rect -3681 10058 -3659 10104
rect -3749 10000 -3659 10058
rect -3749 9954 -3727 10000
rect -3681 9954 -3659 10000
rect -3749 9896 -3659 9954
rect -3749 9850 -3727 9896
rect -3681 9850 -3659 9896
rect -3749 9792 -3659 9850
rect -3749 9746 -3727 9792
rect -3681 9746 -3659 9792
rect -3749 9688 -3659 9746
rect -3749 9642 -3727 9688
rect -3681 9642 -3659 9688
rect -3749 9584 -3659 9642
rect -3749 9538 -3727 9584
rect -3681 9538 -3659 9584
rect -3749 9480 -3659 9538
rect -3749 9434 -3727 9480
rect -3681 9434 -3659 9480
rect -3749 9376 -3659 9434
rect -3749 9330 -3727 9376
rect -3681 9330 -3659 9376
rect -3749 9272 -3659 9330
rect -3749 9226 -3727 9272
rect -3681 9226 -3659 9272
rect -3749 9168 -3659 9226
rect -3749 9122 -3727 9168
rect -3681 9122 -3659 9168
rect -3749 9064 -3659 9122
rect -3749 9018 -3727 9064
rect -3681 9018 -3659 9064
rect -3749 8960 -3659 9018
rect -3749 8914 -3727 8960
rect -3681 8914 -3659 8960
rect -3749 8856 -3659 8914
rect -3749 8810 -3727 8856
rect -3681 8810 -3659 8856
rect -3749 8752 -3659 8810
rect -3749 8706 -3727 8752
rect -3681 8706 -3659 8752
rect -3749 8648 -3659 8706
rect -3749 8602 -3727 8648
rect -3681 8602 -3659 8648
rect -3749 8544 -3659 8602
rect -3749 8498 -3727 8544
rect -3681 8498 -3659 8544
rect -3749 8440 -3659 8498
rect -3749 8394 -3727 8440
rect -3681 8394 -3659 8440
rect -3749 8336 -3659 8394
rect -3749 8290 -3727 8336
rect -3681 8290 -3659 8336
rect -3749 8232 -3659 8290
rect -3749 8186 -3727 8232
rect -3681 8186 -3659 8232
rect -3749 8128 -3659 8186
rect -3749 8082 -3727 8128
rect -3681 8082 -3659 8128
rect -3749 8024 -3659 8082
rect -3749 7978 -3727 8024
rect -3681 7978 -3659 8024
rect -3749 7920 -3659 7978
rect -3749 7874 -3727 7920
rect -3681 7874 -3659 7920
rect -3749 7816 -3659 7874
rect -3749 7770 -3727 7816
rect -3681 7770 -3659 7816
rect -3749 7712 -3659 7770
rect -3749 7666 -3727 7712
rect -3681 7666 -3659 7712
rect -3749 7608 -3659 7666
rect -3749 7562 -3727 7608
rect -3681 7562 -3659 7608
rect -3749 7504 -3659 7562
rect -3749 7458 -3727 7504
rect -3681 7458 -3659 7504
rect -3749 7400 -3659 7458
rect -3749 7354 -3727 7400
rect -3681 7354 -3659 7400
rect -3749 7296 -3659 7354
rect -3749 7250 -3727 7296
rect -3681 7250 -3659 7296
rect -3749 7192 -3659 7250
rect -3749 7146 -3727 7192
rect -3681 7146 -3659 7192
rect -3749 7088 -3659 7146
rect -3749 7042 -3727 7088
rect -3681 7042 -3659 7088
rect -3749 6984 -3659 7042
rect -3749 6938 -3727 6984
rect -3681 6938 -3659 6984
rect -3749 6880 -3659 6938
rect -3749 6834 -3727 6880
rect -3681 6834 -3659 6880
rect -3749 6776 -3659 6834
rect -3749 6730 -3727 6776
rect -3681 6730 -3659 6776
rect -3749 6672 -3659 6730
rect -3749 6626 -3727 6672
rect -3681 6626 -3659 6672
rect -3749 6568 -3659 6626
rect -3749 6522 -3727 6568
rect -3681 6522 -3659 6568
rect -3749 6464 -3659 6522
rect -3749 6418 -3727 6464
rect -3681 6418 -3659 6464
rect -3749 6360 -3659 6418
rect -3749 6314 -3727 6360
rect -3681 6314 -3659 6360
rect -3749 6256 -3659 6314
rect -3749 6210 -3727 6256
rect -3681 6210 -3659 6256
rect -3749 6152 -3659 6210
rect -3749 6106 -3727 6152
rect -3681 6106 -3659 6152
rect -3749 6048 -3659 6106
rect -3749 6002 -3727 6048
rect -3681 6002 -3659 6048
rect -3749 5944 -3659 6002
rect -3749 5898 -3727 5944
rect -3681 5898 -3659 5944
rect -3749 5840 -3659 5898
rect -3749 5794 -3727 5840
rect -3681 5794 -3659 5840
rect -3749 5736 -3659 5794
rect -3749 5690 -3727 5736
rect -3681 5690 -3659 5736
rect -3749 5632 -3659 5690
rect -3749 5586 -3727 5632
rect -3681 5586 -3659 5632
rect -3749 5528 -3659 5586
rect -3749 5482 -3727 5528
rect -3681 5482 -3659 5528
rect -3749 5424 -3659 5482
rect -3749 5378 -3727 5424
rect -3681 5378 -3659 5424
rect -3749 5320 -3659 5378
rect -3749 5274 -3727 5320
rect -3681 5274 -3659 5320
rect -3749 5216 -3659 5274
rect -3749 5170 -3727 5216
rect -3681 5170 -3659 5216
rect -3749 5112 -3659 5170
rect -3749 5066 -3727 5112
rect -3681 5066 -3659 5112
rect -3749 5008 -3659 5066
rect -3749 4962 -3727 5008
rect -3681 4962 -3659 5008
rect -3749 4904 -3659 4962
rect -3749 4858 -3727 4904
rect -3681 4858 -3659 4904
rect -3749 4800 -3659 4858
rect -3749 4754 -3727 4800
rect -3681 4754 -3659 4800
rect -3749 4696 -3659 4754
rect -3749 4650 -3727 4696
rect -3681 4650 -3659 4696
rect -3749 4592 -3659 4650
rect -3749 4546 -3727 4592
rect -3681 4546 -3659 4592
rect -3749 4488 -3659 4546
rect -3749 4442 -3727 4488
rect -3681 4442 -3659 4488
rect -3749 4384 -3659 4442
rect -3749 4338 -3727 4384
rect -3681 4338 -3659 4384
rect -3749 4280 -3659 4338
rect -9 17280 81 17338
rect -9 17234 13 17280
rect 59 17234 81 17280
rect -9 17176 81 17234
rect -9 17130 13 17176
rect 59 17130 81 17176
rect -9 17072 81 17130
rect -9 17026 13 17072
rect 59 17026 81 17072
rect -9 16968 81 17026
rect -9 16922 13 16968
rect 59 16922 81 16968
rect -9 16864 81 16922
rect -9 16818 13 16864
rect 59 16818 81 16864
rect -9 16760 81 16818
rect -9 16714 13 16760
rect 59 16714 81 16760
rect -9 16656 81 16714
rect -9 16610 13 16656
rect 59 16610 81 16656
rect -9 16552 81 16610
rect -9 16506 13 16552
rect 59 16506 81 16552
rect -9 16448 81 16506
rect -9 16402 13 16448
rect 59 16402 81 16448
rect -9 16344 81 16402
rect -9 16298 13 16344
rect 59 16298 81 16344
rect -9 16240 81 16298
rect -9 16194 13 16240
rect 59 16194 81 16240
rect -9 16136 81 16194
rect -9 16090 13 16136
rect 59 16090 81 16136
rect -9 16032 81 16090
rect -9 15986 13 16032
rect 59 15986 81 16032
rect -9 15928 81 15986
rect -9 15882 13 15928
rect 59 15882 81 15928
rect -9 15824 81 15882
rect -9 15778 13 15824
rect 59 15778 81 15824
rect -9 15720 81 15778
rect -9 15674 13 15720
rect 59 15674 81 15720
rect -9 15616 81 15674
rect -9 15570 13 15616
rect 59 15570 81 15616
rect -9 15512 81 15570
rect -9 15466 13 15512
rect 59 15466 81 15512
rect -9 15408 81 15466
rect -9 15362 13 15408
rect 59 15362 81 15408
rect -9 15304 81 15362
rect -9 15258 13 15304
rect 59 15258 81 15304
rect -9 15200 81 15258
rect -9 15154 13 15200
rect 59 15154 81 15200
rect -9 15096 81 15154
rect -9 15050 13 15096
rect 59 15050 81 15096
rect -9 14992 81 15050
rect -9 14946 13 14992
rect 59 14946 81 14992
rect -9 14888 81 14946
rect -9 14842 13 14888
rect 59 14842 81 14888
rect -9 14784 81 14842
rect -9 14738 13 14784
rect 59 14738 81 14784
rect -9 14680 81 14738
rect -9 14634 13 14680
rect 59 14634 81 14680
rect -9 14576 81 14634
rect -9 14530 13 14576
rect 59 14530 81 14576
rect -9 14472 81 14530
rect -9 14426 13 14472
rect 59 14426 81 14472
rect -9 14368 81 14426
rect -9 14322 13 14368
rect 59 14322 81 14368
rect -9 14264 81 14322
rect -9 14218 13 14264
rect 59 14218 81 14264
rect -9 14160 81 14218
rect -9 14114 13 14160
rect 59 14114 81 14160
rect -9 14056 81 14114
rect -9 14010 13 14056
rect 59 14010 81 14056
rect -9 13952 81 14010
rect -9 13906 13 13952
rect 59 13906 81 13952
rect -9 13848 81 13906
rect -9 13802 13 13848
rect 59 13802 81 13848
rect -9 13744 81 13802
rect -9 13698 13 13744
rect 59 13698 81 13744
rect -9 13640 81 13698
rect -9 13594 13 13640
rect 59 13594 81 13640
rect -9 13536 81 13594
rect -9 13490 13 13536
rect 59 13490 81 13536
rect -9 13432 81 13490
rect -9 13386 13 13432
rect 59 13386 81 13432
rect -9 13328 81 13386
rect -9 13282 13 13328
rect 59 13282 81 13328
rect -9 13224 81 13282
rect -9 13178 13 13224
rect 59 13178 81 13224
rect -9 13120 81 13178
rect -9 13074 13 13120
rect 59 13074 81 13120
rect -9 13016 81 13074
rect -9 12970 13 13016
rect 59 12970 81 13016
rect -9 12912 81 12970
rect -9 12866 13 12912
rect 59 12866 81 12912
rect -9 12808 81 12866
rect -9 12762 13 12808
rect 59 12762 81 12808
rect -9 12704 81 12762
rect -9 12658 13 12704
rect 59 12658 81 12704
rect -9 12600 81 12658
rect -9 12554 13 12600
rect 59 12554 81 12600
rect -9 12496 81 12554
rect -9 12450 13 12496
rect 59 12450 81 12496
rect -9 12392 81 12450
rect -9 12346 13 12392
rect 59 12346 81 12392
rect -9 12288 81 12346
rect -9 12242 13 12288
rect 59 12242 81 12288
rect -9 12184 81 12242
rect -9 12138 13 12184
rect 59 12138 81 12184
rect -9 12080 81 12138
rect -9 12034 13 12080
rect 59 12034 81 12080
rect -9 11976 81 12034
rect -9 11930 13 11976
rect 59 11930 81 11976
rect -9 11872 81 11930
rect -9 11826 13 11872
rect 59 11826 81 11872
rect -9 11768 81 11826
rect -9 11722 13 11768
rect 59 11722 81 11768
rect -9 11664 81 11722
rect -9 11618 13 11664
rect 59 11618 81 11664
rect -9 11560 81 11618
rect -9 11514 13 11560
rect 59 11514 81 11560
rect -9 11456 81 11514
rect -9 11410 13 11456
rect 59 11410 81 11456
rect -9 11352 81 11410
rect -9 11306 13 11352
rect 59 11306 81 11352
rect -9 11248 81 11306
rect -9 11202 13 11248
rect 59 11202 81 11248
rect -9 11144 81 11202
rect -9 11098 13 11144
rect 59 11098 81 11144
rect -9 11040 81 11098
rect -9 10994 13 11040
rect 59 10994 81 11040
rect -9 10936 81 10994
rect -9 10890 13 10936
rect 59 10890 81 10936
rect -9 10832 81 10890
rect -9 10786 13 10832
rect 59 10786 81 10832
rect -9 10728 81 10786
rect -9 10682 13 10728
rect 59 10682 81 10728
rect -9 10624 81 10682
rect -9 10578 13 10624
rect 59 10578 81 10624
rect -9 10520 81 10578
rect -9 10474 13 10520
rect 59 10474 81 10520
rect -9 10416 81 10474
rect -9 10370 13 10416
rect 59 10370 81 10416
rect -9 10312 81 10370
rect -9 10266 13 10312
rect 59 10266 81 10312
rect -9 10208 81 10266
rect -9 10162 13 10208
rect 59 10162 81 10208
rect -9 10104 81 10162
rect -9 10058 13 10104
rect 59 10058 81 10104
rect -9 10000 81 10058
rect -9 9954 13 10000
rect 59 9954 81 10000
rect -9 9896 81 9954
rect -9 9850 13 9896
rect 59 9850 81 9896
rect -9 9792 81 9850
rect -9 9746 13 9792
rect 59 9746 81 9792
rect -9 9688 81 9746
rect -9 9642 13 9688
rect 59 9642 81 9688
rect -9 9584 81 9642
rect -9 9538 13 9584
rect 59 9538 81 9584
rect -9 9480 81 9538
rect -9 9434 13 9480
rect 59 9434 81 9480
rect -9 9376 81 9434
rect -9 9330 13 9376
rect 59 9330 81 9376
rect -9 9272 81 9330
rect -9 9226 13 9272
rect 59 9226 81 9272
rect -9 9168 81 9226
rect -9 9122 13 9168
rect 59 9122 81 9168
rect -9 9064 81 9122
rect -9 9018 13 9064
rect 59 9018 81 9064
rect -9 8960 81 9018
rect -9 8914 13 8960
rect 59 8914 81 8960
rect -9 8856 81 8914
rect -9 8810 13 8856
rect 59 8810 81 8856
rect -9 8752 81 8810
rect -9 8706 13 8752
rect 59 8706 81 8752
rect -9 8648 81 8706
rect -9 8602 13 8648
rect 59 8602 81 8648
rect -9 8544 81 8602
rect -9 8498 13 8544
rect 59 8498 81 8544
rect -9 8440 81 8498
rect -9 8394 13 8440
rect 59 8394 81 8440
rect -9 8336 81 8394
rect -9 8290 13 8336
rect 59 8290 81 8336
rect -9 8232 81 8290
rect -9 8186 13 8232
rect 59 8186 81 8232
rect -9 8128 81 8186
rect -9 8082 13 8128
rect 59 8082 81 8128
rect -9 8024 81 8082
rect -9 7978 13 8024
rect 59 7978 81 8024
rect -9 7920 81 7978
rect -9 7874 13 7920
rect 59 7874 81 7920
rect -9 7816 81 7874
rect -9 7770 13 7816
rect 59 7770 81 7816
rect -9 7712 81 7770
rect -9 7666 13 7712
rect 59 7666 81 7712
rect -9 7608 81 7666
rect -9 7562 13 7608
rect 59 7562 81 7608
rect -9 7504 81 7562
rect -9 7458 13 7504
rect 59 7458 81 7504
rect -9 7400 81 7458
rect -9 7354 13 7400
rect 59 7354 81 7400
rect -9 7296 81 7354
rect -9 7250 13 7296
rect 59 7250 81 7296
rect -9 7192 81 7250
rect -9 7146 13 7192
rect 59 7146 81 7192
rect -9 7088 81 7146
rect -9 7042 13 7088
rect 59 7042 81 7088
rect -9 6984 81 7042
rect -9 6938 13 6984
rect 59 6938 81 6984
rect -9 6880 81 6938
rect -9 6834 13 6880
rect 59 6834 81 6880
rect -9 6776 81 6834
rect -9 6730 13 6776
rect 59 6730 81 6776
rect -9 6672 81 6730
rect -9 6626 13 6672
rect 59 6626 81 6672
rect -9 6568 81 6626
rect -9 6522 13 6568
rect 59 6522 81 6568
rect -9 6464 81 6522
rect -9 6418 13 6464
rect 59 6418 81 6464
rect -9 6360 81 6418
rect -9 6314 13 6360
rect 59 6314 81 6360
rect -9 6256 81 6314
rect -9 6210 13 6256
rect 59 6210 81 6256
rect -9 6152 81 6210
rect -9 6106 13 6152
rect 59 6106 81 6152
rect -9 6048 81 6106
rect -9 6002 13 6048
rect 59 6002 81 6048
rect -9 5944 81 6002
rect -9 5898 13 5944
rect 59 5898 81 5944
rect -9 5840 81 5898
rect -9 5794 13 5840
rect 59 5794 81 5840
rect -9 5736 81 5794
rect -9 5690 13 5736
rect 59 5690 81 5736
rect -9 5632 81 5690
rect -9 5586 13 5632
rect 59 5586 81 5632
rect -9 5528 81 5586
rect -9 5482 13 5528
rect 59 5482 81 5528
rect -9 5424 81 5482
rect -9 5378 13 5424
rect 59 5378 81 5424
rect -9 5320 81 5378
rect -9 5274 13 5320
rect 59 5274 81 5320
rect -9 5216 81 5274
rect -9 5170 13 5216
rect 59 5170 81 5216
rect -9 5112 81 5170
rect -9 5066 13 5112
rect 59 5066 81 5112
rect -9 5008 81 5066
rect -9 4962 13 5008
rect 59 4962 81 5008
rect -9 4904 81 4962
rect -9 4858 13 4904
rect 59 4858 81 4904
rect -9 4800 81 4858
rect -9 4754 13 4800
rect 59 4754 81 4800
rect -9 4696 81 4754
rect -9 4650 13 4696
rect 59 4650 81 4696
rect -9 4592 81 4650
rect -9 4546 13 4592
rect 59 4546 81 4592
rect -3749 4234 -3727 4280
rect -3681 4234 -3659 4280
rect -3749 4176 -3659 4234
rect -3749 4130 -3727 4176
rect -3681 4130 -3659 4176
rect -3749 4094 -3659 4130
rect -9 4176 81 4546
rect -9 4130 13 4176
rect 59 4130 81 4176
rect -9 4094 81 4130
rect -3749 4072 81 4094
rect -3749 4026 -3727 4072
rect -3681 4026 -3573 4072
rect -3527 4026 -3469 4072
rect -3423 4026 -3365 4072
rect -3319 4026 -3261 4072
rect -3215 4026 -3157 4072
rect -3111 4026 -3053 4072
rect -3007 4026 -2949 4072
rect -2903 4026 -2845 4072
rect -2799 4026 -2741 4072
rect -2695 4026 -2637 4072
rect -2591 4026 -2533 4072
rect -2487 4026 -2429 4072
rect -2383 4026 -2325 4072
rect -2279 4026 -2221 4072
rect -2175 4026 -2117 4072
rect -2071 4026 -2013 4072
rect -1967 4026 -1909 4072
rect -1863 4026 -1805 4072
rect -1759 4026 -1701 4072
rect -1655 4026 -1597 4072
rect -1551 4026 -1493 4072
rect -1447 4026 -1389 4072
rect -1343 4026 -1285 4072
rect -1239 4026 -1181 4072
rect -1135 4026 -1077 4072
rect -1031 4026 -973 4072
rect -927 4026 -869 4072
rect -823 4026 -765 4072
rect -719 4026 -661 4072
rect -615 4026 -557 4072
rect -511 4026 -453 4072
rect -407 4026 -349 4072
rect -303 4026 -245 4072
rect -199 4026 -141 4072
rect -95 4026 13 4072
rect 59 4026 81 4072
rect -3749 4004 81 4026
<< psubdiffcont >>
rect 1587 16970 1633 17016
rect 1701 16970 1747 17016
rect 1855 16970 1901 17016
rect 1969 16970 2015 17016
rect 2083 16970 2129 17016
rect 2197 16970 2243 17016
rect 2311 16970 2357 17016
rect 2425 16970 2471 17016
rect 2539 16970 2585 17016
rect 2653 16970 2699 17016
rect 2767 16970 2813 17016
rect 2881 16970 2927 17016
rect 2995 16970 3041 17016
rect 3109 16970 3155 17016
rect 3223 16970 3269 17016
rect 3337 16970 3383 17016
rect 3451 16970 3497 17016
rect 3565 16970 3611 17016
rect 3679 16970 3725 17016
rect 3793 16970 3839 17016
rect 3907 16970 3953 17016
rect 4021 16970 4067 17016
rect 4135 16970 4181 17016
rect 4249 16970 4295 17016
rect 4363 16970 4409 17016
rect 4477 16970 4523 17016
rect 4591 16970 4637 17016
rect 4705 16970 4751 17016
rect 4819 16970 4865 17016
rect 4933 16970 4979 17016
rect 5047 16970 5093 17016
rect 5161 16970 5207 17016
rect 5275 16970 5321 17016
rect 5389 16970 5435 17016
rect 5503 16970 5549 17016
rect 5617 16970 5663 17016
rect 5731 16970 5777 17016
rect 5845 16970 5891 17016
rect 5959 16970 6005 17016
rect 6073 16970 6119 17016
rect 6187 16970 6233 17016
rect 6301 16970 6347 17016
rect 6415 16970 6461 17016
rect 6529 16970 6575 17016
rect 6643 16970 6689 17016
rect 6757 16970 6803 17016
rect 6871 16970 6917 17016
rect 6985 16970 7031 17016
rect 7099 16970 7145 17016
rect 7213 16970 7259 17016
rect 7327 16970 7373 17016
rect 7441 16970 7487 17016
rect 7555 16970 7601 17016
rect 7669 16970 7715 17016
rect 7783 16970 7829 17016
rect 7897 16970 7943 17016
rect 8011 16970 8057 17016
rect 8125 16970 8171 17016
rect 8239 16970 8285 17016
rect 8353 16970 8399 17016
rect 8467 16970 8513 17016
rect 8581 16970 8627 17016
rect 8695 16970 8741 17016
rect 8809 16970 8855 17016
rect 8923 16970 8969 17016
rect 9037 16970 9083 17016
rect 9151 16970 9197 17016
rect 9265 16970 9311 17016
rect 9379 16970 9425 17016
rect 9493 16970 9539 17016
rect 9607 16970 9653 17016
rect 9721 16970 9767 17016
rect 9835 16970 9881 17016
rect 9949 16970 9995 17016
rect 10063 16970 10109 17016
rect 10177 16970 10223 17016
rect 10291 16970 10337 17016
rect 10405 16970 10451 17016
rect 10519 16970 10565 17016
rect 10633 16970 10679 17016
rect 10747 16970 10793 17016
rect 10861 16970 10907 17016
rect 10975 16970 11021 17016
rect 11089 16970 11135 17016
rect 11203 16970 11249 17016
rect 11317 16970 11363 17016
rect 11431 16970 11477 17016
rect 11545 16970 11591 17016
rect 11659 16970 11705 17016
rect 11773 16970 11819 17016
rect 11927 16970 11973 17016
rect 12041 16970 12087 17016
rect 1587 16856 1633 16902
rect 1701 16856 1747 16902
rect 1855 16856 1901 16902
rect 1969 16856 2015 16902
rect 2083 16856 2129 16902
rect 2197 16856 2243 16902
rect 2311 16856 2357 16902
rect 2425 16856 2471 16902
rect 2539 16856 2585 16902
rect 2653 16856 2699 16902
rect 2767 16856 2813 16902
rect 2881 16856 2927 16902
rect 2995 16856 3041 16902
rect 3109 16856 3155 16902
rect 3223 16856 3269 16902
rect 3337 16856 3383 16902
rect 3451 16856 3497 16902
rect 3565 16856 3611 16902
rect 3679 16856 3725 16902
rect 3793 16856 3839 16902
rect 3907 16856 3953 16902
rect 4021 16856 4067 16902
rect 4135 16856 4181 16902
rect 4249 16856 4295 16902
rect 4363 16856 4409 16902
rect 4477 16856 4523 16902
rect 4591 16856 4637 16902
rect 4705 16856 4751 16902
rect 4819 16856 4865 16902
rect 4933 16856 4979 16902
rect 5047 16856 5093 16902
rect 5161 16856 5207 16902
rect 5275 16856 5321 16902
rect 5389 16856 5435 16902
rect 5503 16856 5549 16902
rect 5617 16856 5663 16902
rect 5731 16856 5777 16902
rect 5845 16856 5891 16902
rect 5959 16856 6005 16902
rect 6073 16856 6119 16902
rect 6187 16856 6233 16902
rect 6301 16856 6347 16902
rect 6415 16856 6461 16902
rect 6529 16856 6575 16902
rect 6643 16856 6689 16902
rect 6757 16856 6803 16902
rect 6871 16856 6917 16902
rect 6985 16856 7031 16902
rect 7099 16856 7145 16902
rect 7213 16856 7259 16902
rect 7327 16856 7373 16902
rect 7441 16856 7487 16902
rect 7555 16856 7601 16902
rect 7669 16856 7715 16902
rect 7783 16856 7829 16902
rect 7897 16856 7943 16902
rect 8011 16856 8057 16902
rect 8125 16856 8171 16902
rect 8239 16856 8285 16902
rect 8353 16856 8399 16902
rect 8467 16856 8513 16902
rect 8581 16856 8627 16902
rect 8695 16856 8741 16902
rect 8809 16856 8855 16902
rect 8923 16856 8969 16902
rect 9037 16856 9083 16902
rect 9151 16856 9197 16902
rect 9265 16856 9311 16902
rect 9379 16856 9425 16902
rect 9493 16856 9539 16902
rect 9607 16856 9653 16902
rect 9721 16856 9767 16902
rect 9835 16856 9881 16902
rect 9949 16856 9995 16902
rect 10063 16856 10109 16902
rect 10177 16856 10223 16902
rect 10291 16856 10337 16902
rect 10405 16856 10451 16902
rect 10519 16856 10565 16902
rect 10633 16856 10679 16902
rect 10747 16856 10793 16902
rect 10861 16856 10907 16902
rect 10975 16856 11021 16902
rect 11089 16856 11135 16902
rect 11203 16856 11249 16902
rect 11317 16856 11363 16902
rect 11431 16856 11477 16902
rect 11545 16856 11591 16902
rect 11659 16856 11705 16902
rect 11773 16856 11819 16902
rect 11927 16856 11973 16902
rect 12041 16856 12087 16902
rect 1587 16742 1633 16788
rect 1701 16742 1747 16788
rect 11927 16742 11973 16788
rect 12041 16742 12087 16788
rect 11927 16628 11973 16674
rect 12041 16628 12087 16674
rect 11927 16514 11973 16560
rect 12041 16514 12087 16560
rect 11927 16400 11973 16446
rect 12041 16400 12087 16446
rect 1587 16172 1633 16218
rect 1701 16172 1747 16218
rect 1587 16058 1633 16104
rect 1701 16058 1747 16104
rect 1587 15944 1633 15990
rect 1701 15944 1747 15990
rect 1587 15830 1633 15876
rect 1701 15830 1747 15876
rect 1587 15716 1633 15762
rect 1701 15716 1747 15762
rect 1587 15602 1633 15648
rect 1701 15602 1747 15648
rect 1587 15488 1633 15534
rect 1701 15488 1747 15534
rect 1587 15374 1633 15420
rect 1701 15374 1747 15420
rect 1587 15260 1633 15306
rect 1701 15260 1747 15306
rect 1587 15146 1633 15192
rect 1701 15146 1747 15192
rect 1587 15032 1633 15078
rect 1701 15032 1747 15078
rect 1587 14918 1633 14964
rect 1701 14918 1747 14964
rect 1587 14804 1633 14850
rect 1701 14804 1747 14850
rect 1587 14690 1633 14736
rect 1701 14690 1747 14736
rect 1587 14576 1633 14622
rect 1701 14576 1747 14622
rect 1587 14462 1633 14508
rect 1701 14462 1747 14508
rect 1587 14348 1633 14394
rect 1701 14348 1747 14394
rect 1587 14234 1633 14280
rect 1701 14234 1747 14280
rect 1587 14120 1633 14166
rect 1701 14120 1747 14166
rect 1587 14006 1633 14052
rect 1701 14006 1747 14052
rect 1587 13892 1633 13938
rect 1701 13892 1747 13938
rect 1587 13778 1633 13824
rect 1701 13778 1747 13824
rect 1587 13664 1633 13710
rect 1701 13664 1747 13710
rect 1587 13550 1633 13596
rect 1701 13550 1747 13596
rect 1587 13436 1633 13482
rect 1701 13436 1747 13482
rect 1587 13322 1633 13368
rect 1701 13322 1747 13368
rect 1587 13208 1633 13254
rect 1701 13208 1747 13254
rect 1587 13094 1633 13140
rect 1701 13094 1747 13140
rect 1587 12980 1633 13026
rect 1701 12980 1747 13026
rect 1587 12866 1633 12912
rect 1701 12866 1747 12912
rect 1587 12752 1633 12798
rect 1701 12752 1747 12798
rect 1587 12638 1633 12684
rect 1701 12638 1747 12684
rect 1587 12524 1633 12570
rect 1701 12524 1747 12570
rect 1587 12410 1633 12456
rect 1701 12410 1747 12456
rect 1587 12296 1633 12342
rect 1701 12296 1747 12342
rect 1587 12182 1633 12228
rect 1701 12182 1747 12228
rect 1587 12068 1633 12114
rect 1701 12068 1747 12114
rect 1587 11954 1633 12000
rect 1701 11954 1747 12000
rect 1587 11840 1633 11886
rect 1701 11840 1747 11886
rect 1587 11726 1633 11772
rect 1701 11726 1747 11772
rect 1587 11612 1633 11658
rect 1701 11612 1747 11658
rect 1587 11498 1633 11544
rect 1701 11498 1747 11544
rect 1587 11384 1633 11430
rect 1701 11384 1747 11430
rect 11927 16286 11973 16332
rect 12041 16286 12087 16332
rect 11927 16172 11973 16218
rect 12041 16172 12087 16218
rect 11927 16058 11973 16104
rect 12041 16058 12087 16104
rect 11927 15944 11973 15990
rect 12041 15944 12087 15990
rect 11927 15830 11973 15876
rect 12041 15830 12087 15876
rect 11927 15716 11973 15762
rect 12041 15716 12087 15762
rect 11927 15602 11973 15648
rect 12041 15602 12087 15648
rect 11927 15488 11973 15534
rect 12041 15488 12087 15534
rect 11927 15374 11973 15420
rect 12041 15374 12087 15420
rect 11927 15260 11973 15306
rect 12041 15260 12087 15306
rect 11927 15146 11973 15192
rect 12041 15146 12087 15192
rect 11927 15032 11973 15078
rect 12041 15032 12087 15078
rect 11927 14918 11973 14964
rect 12041 14918 12087 14964
rect 11927 14804 11973 14850
rect 12041 14804 12087 14850
rect 11927 14690 11973 14736
rect 12041 14690 12087 14736
rect 11927 14576 11973 14622
rect 12041 14576 12087 14622
rect 11927 14462 11973 14508
rect 12041 14462 12087 14508
rect 11927 14348 11973 14394
rect 12041 14348 12087 14394
rect 11927 14234 11973 14280
rect 12041 14234 12087 14280
rect 11927 14120 11973 14166
rect 12041 14120 12087 14166
rect 11927 14006 11973 14052
rect 12041 14006 12087 14052
rect 11927 13892 11973 13938
rect 12041 13892 12087 13938
rect 11927 13778 11973 13824
rect 12041 13778 12087 13824
rect 11927 13664 11973 13710
rect 12041 13664 12087 13710
rect 11927 13550 11973 13596
rect 12041 13550 12087 13596
rect 11927 13436 11973 13482
rect 12041 13436 12087 13482
rect 11927 13322 11973 13368
rect 12041 13322 12087 13368
rect 11927 13208 11973 13254
rect 12041 13208 12087 13254
rect 11927 13094 11973 13140
rect 12041 13094 12087 13140
rect 11927 12980 11973 13026
rect 12041 12980 12087 13026
rect 11927 12866 11973 12912
rect 12041 12866 12087 12912
rect 11927 12752 11973 12798
rect 12041 12752 12087 12798
rect 11927 12638 11973 12684
rect 12041 12638 12087 12684
rect 11927 12524 11973 12570
rect 12041 12524 12087 12570
rect 11927 12410 11973 12456
rect 12041 12410 12087 12456
rect 11927 12296 11973 12342
rect 12041 12296 12087 12342
rect 11927 12182 11973 12228
rect 12041 12182 12087 12228
rect 11927 12068 11973 12114
rect 12041 12068 12087 12114
rect 11927 11954 11973 12000
rect 12041 11954 12087 12000
rect 11927 11840 11973 11886
rect 12041 11840 12087 11886
rect 11927 11726 11973 11772
rect 12041 11726 12087 11772
rect 11927 11612 11973 11658
rect 12041 11612 12087 11658
rect 11927 11498 11973 11544
rect 12041 11498 12087 11544
rect 11927 11384 11973 11430
rect 12041 11384 12087 11430
rect 1587 11270 1633 11316
rect 1701 11270 1747 11316
rect 11927 11270 11973 11316
rect 12041 11270 12087 11316
rect 1587 11156 1633 11202
rect 1701 11156 1747 11202
rect 1587 11042 1633 11088
rect 1701 11042 1747 11088
rect 1587 10928 1633 10974
rect 1701 10928 1747 10974
rect 11927 11156 11973 11202
rect 12041 11156 12087 11202
rect 11927 11042 11973 11088
rect 12041 11042 12087 11088
rect 11927 10928 11973 10974
rect 12041 10928 12087 10974
rect 1855 10879 1901 10925
rect 1969 10879 2015 10925
rect 2083 10879 2129 10925
rect 2197 10879 2243 10925
rect 2311 10879 2357 10925
rect 2425 10879 2471 10925
rect 2539 10879 2585 10925
rect 2653 10879 2699 10925
rect 2767 10879 2813 10925
rect 2881 10879 2927 10925
rect 2995 10879 3041 10925
rect 3109 10879 3155 10925
rect 3223 10879 3269 10925
rect 3337 10879 3383 10925
rect 3451 10879 3497 10925
rect 3565 10879 3611 10925
rect 3679 10879 3725 10925
rect 3793 10879 3839 10925
rect 3907 10879 3953 10925
rect 4021 10879 4067 10925
rect 4135 10879 4181 10925
rect 4249 10879 4295 10925
rect 4363 10879 4409 10925
rect 4477 10879 4523 10925
rect 4591 10879 4637 10925
rect 4705 10879 4751 10925
rect 4819 10879 4865 10925
rect 4933 10879 4979 10925
rect 5047 10879 5093 10925
rect 5161 10879 5207 10925
rect 5275 10879 5321 10925
rect 5389 10879 5435 10925
rect 5503 10879 5549 10925
rect 5617 10879 5663 10925
rect 5731 10879 5777 10925
rect 5845 10879 5891 10925
rect 5959 10879 6005 10925
rect 6073 10879 6119 10925
rect 6187 10879 6233 10925
rect 6301 10879 6347 10925
rect 6415 10879 6461 10925
rect 6529 10879 6575 10925
rect 6643 10879 6689 10925
rect 6757 10879 6803 10925
rect 6871 10879 6917 10925
rect 6985 10879 7031 10925
rect 7099 10879 7145 10925
rect 7213 10879 7259 10925
rect 7327 10879 7373 10925
rect 7441 10879 7487 10925
rect 7555 10879 7601 10925
rect 7669 10879 7715 10925
rect 7783 10879 7829 10925
rect 7897 10879 7943 10925
rect 8011 10879 8057 10925
rect 8125 10879 8171 10925
rect 8239 10879 8285 10925
rect 8353 10879 8399 10925
rect 8467 10879 8513 10925
rect 8581 10879 8627 10925
rect 8695 10879 8741 10925
rect 8809 10879 8855 10925
rect 8923 10879 8969 10925
rect 9037 10879 9083 10925
rect 9151 10879 9197 10925
rect 9265 10879 9311 10925
rect 9379 10879 9425 10925
rect 9493 10879 9539 10925
rect 9607 10879 9653 10925
rect 9721 10879 9767 10925
rect 9835 10879 9881 10925
rect 9949 10879 9995 10925
rect 10063 10879 10109 10925
rect 10177 10879 10223 10925
rect 10291 10879 10337 10925
rect 10405 10879 10451 10925
rect 10519 10879 10565 10925
rect 10633 10879 10679 10925
rect 10747 10879 10793 10925
rect 10861 10879 10907 10925
rect 10975 10879 11021 10925
rect 11089 10879 11135 10925
rect 11203 10879 11249 10925
rect 11317 10879 11363 10925
rect 11431 10879 11477 10925
rect 11545 10879 11591 10925
rect 11659 10879 11705 10925
rect 11773 10879 11819 10925
rect 1587 10814 1633 10860
rect 1701 10814 1747 10860
rect 11927 10814 11973 10860
rect 12041 10814 12087 10860
rect 1855 10765 1901 10811
rect 1969 10765 2015 10811
rect 2083 10765 2129 10811
rect 2197 10765 2243 10811
rect 2311 10765 2357 10811
rect 2425 10765 2471 10811
rect 2539 10765 2585 10811
rect 2653 10765 2699 10811
rect 2767 10765 2813 10811
rect 2881 10765 2927 10811
rect 2995 10765 3041 10811
rect 3109 10765 3155 10811
rect 3223 10765 3269 10811
rect 3337 10765 3383 10811
rect 3451 10765 3497 10811
rect 3565 10765 3611 10811
rect 3679 10765 3725 10811
rect 3793 10765 3839 10811
rect 3907 10765 3953 10811
rect 4021 10765 4067 10811
rect 4135 10765 4181 10811
rect 4249 10765 4295 10811
rect 4363 10765 4409 10811
rect 4477 10765 4523 10811
rect 4591 10765 4637 10811
rect 4705 10765 4751 10811
rect 4819 10765 4865 10811
rect 4933 10765 4979 10811
rect 5047 10765 5093 10811
rect 5161 10765 5207 10811
rect 5275 10765 5321 10811
rect 5389 10765 5435 10811
rect 5503 10765 5549 10811
rect 5617 10765 5663 10811
rect 5731 10765 5777 10811
rect 5845 10765 5891 10811
rect 5959 10765 6005 10811
rect 6073 10765 6119 10811
rect 6187 10765 6233 10811
rect 6301 10765 6347 10811
rect 6415 10765 6461 10811
rect 6529 10765 6575 10811
rect 6643 10765 6689 10811
rect 6757 10765 6803 10811
rect 6871 10765 6917 10811
rect 6985 10765 7031 10811
rect 7099 10765 7145 10811
rect 7213 10765 7259 10811
rect 7327 10765 7373 10811
rect 7441 10765 7487 10811
rect 7555 10765 7601 10811
rect 7669 10765 7715 10811
rect 7783 10765 7829 10811
rect 7897 10765 7943 10811
rect 8011 10765 8057 10811
rect 8125 10765 8171 10811
rect 8239 10765 8285 10811
rect 8353 10765 8399 10811
rect 8467 10765 8513 10811
rect 8581 10765 8627 10811
rect 8695 10765 8741 10811
rect 8809 10765 8855 10811
rect 8923 10765 8969 10811
rect 9037 10765 9083 10811
rect 9151 10765 9197 10811
rect 9265 10765 9311 10811
rect 9379 10765 9425 10811
rect 9493 10765 9539 10811
rect 9607 10765 9653 10811
rect 9721 10765 9767 10811
rect 9835 10765 9881 10811
rect 9949 10765 9995 10811
rect 10063 10765 10109 10811
rect 10177 10765 10223 10811
rect 10291 10765 10337 10811
rect 10405 10765 10451 10811
rect 10519 10765 10565 10811
rect 10633 10765 10679 10811
rect 10747 10765 10793 10811
rect 10861 10765 10907 10811
rect 10975 10765 11021 10811
rect 11089 10765 11135 10811
rect 11203 10765 11249 10811
rect 11317 10765 11363 10811
rect 11431 10765 11477 10811
rect 11545 10765 11591 10811
rect 11659 10765 11705 10811
rect 11773 10765 11819 10811
rect 1587 10700 1633 10746
rect 1701 10700 1747 10746
rect 1587 10586 1633 10632
rect 1701 10586 1747 10632
rect 1587 10472 1633 10518
rect 1701 10472 1747 10518
rect 11927 10700 11973 10746
rect 12041 10700 12087 10746
rect 11927 10586 11973 10632
rect 12041 10586 12087 10632
rect 11927 10472 11973 10518
rect 12041 10472 12087 10518
rect 1587 10358 1633 10404
rect 1701 10358 1747 10404
rect 11927 10358 11973 10404
rect 12041 10358 12087 10404
rect 1587 10244 1633 10290
rect 1701 10244 1747 10290
rect 1587 10130 1633 10176
rect 1701 10130 1747 10176
rect 1587 10016 1633 10062
rect 1701 10016 1747 10062
rect 1587 9902 1633 9948
rect 1701 9902 1747 9948
rect 1587 9788 1633 9834
rect 1701 9788 1747 9834
rect 1587 9674 1633 9720
rect 1701 9674 1747 9720
rect 1587 9560 1633 9606
rect 1701 9560 1747 9606
rect 1587 9446 1633 9492
rect 1701 9446 1747 9492
rect 1587 9332 1633 9378
rect 1701 9332 1747 9378
rect 1587 9218 1633 9264
rect 1701 9218 1747 9264
rect 1587 9104 1633 9150
rect 1701 9104 1747 9150
rect 1587 8990 1633 9036
rect 1701 8990 1747 9036
rect 1587 8876 1633 8922
rect 1701 8876 1747 8922
rect 1587 8762 1633 8808
rect 1701 8762 1747 8808
rect 1587 8648 1633 8694
rect 1701 8648 1747 8694
rect 1587 8534 1633 8580
rect 1701 8534 1747 8580
rect 1587 8420 1633 8466
rect 1701 8420 1747 8466
rect 1587 8306 1633 8352
rect 1701 8306 1747 8352
rect 1587 8192 1633 8238
rect 1701 8192 1747 8238
rect 1587 8078 1633 8124
rect 1701 8078 1747 8124
rect 1587 7964 1633 8010
rect 1701 7964 1747 8010
rect 1587 7850 1633 7896
rect 1701 7850 1747 7896
rect 1587 7736 1633 7782
rect 1701 7736 1747 7782
rect 1587 7622 1633 7668
rect 1701 7622 1747 7668
rect 1587 7508 1633 7554
rect 1701 7508 1747 7554
rect 1587 7394 1633 7440
rect 1701 7394 1747 7440
rect 1587 7280 1633 7326
rect 1701 7280 1747 7326
rect 1587 7166 1633 7212
rect 1701 7166 1747 7212
rect 1587 7052 1633 7098
rect 1701 7052 1747 7098
rect 1587 6938 1633 6984
rect 1701 6938 1747 6984
rect 1587 6824 1633 6870
rect 1701 6824 1747 6870
rect 1587 6710 1633 6756
rect 1701 6710 1747 6756
rect 1587 6596 1633 6642
rect 1701 6596 1747 6642
rect 1587 6482 1633 6528
rect 1701 6482 1747 6528
rect 1587 6368 1633 6414
rect 1701 6368 1747 6414
rect 1587 6254 1633 6300
rect 1701 6254 1747 6300
rect 1587 6140 1633 6186
rect 1701 6140 1747 6186
rect 1587 6026 1633 6072
rect 1701 6026 1747 6072
rect 1587 5912 1633 5958
rect 1701 5912 1747 5958
rect 1587 5798 1633 5844
rect 1701 5798 1747 5844
rect 1587 5684 1633 5730
rect 1701 5684 1747 5730
rect 1587 5570 1633 5616
rect 1701 5570 1747 5616
rect 1587 5456 1633 5502
rect 1701 5456 1747 5502
rect 11927 10244 11973 10290
rect 12041 10244 12087 10290
rect 11927 10130 11973 10176
rect 12041 10130 12087 10176
rect 11927 10016 11973 10062
rect 12041 10016 12087 10062
rect 11927 9902 11973 9948
rect 12041 9902 12087 9948
rect 11927 9788 11973 9834
rect 12041 9788 12087 9834
rect 11927 9674 11973 9720
rect 12041 9674 12087 9720
rect 11927 9560 11973 9606
rect 12041 9560 12087 9606
rect 11927 9446 11973 9492
rect 12041 9446 12087 9492
rect 11927 9332 11973 9378
rect 12041 9332 12087 9378
rect 11927 9218 11973 9264
rect 12041 9218 12087 9264
rect 11927 9104 11973 9150
rect 12041 9104 12087 9150
rect 11927 8990 11973 9036
rect 12041 8990 12087 9036
rect 11927 8876 11973 8922
rect 12041 8876 12087 8922
rect 11927 8762 11973 8808
rect 12041 8762 12087 8808
rect 11927 8648 11973 8694
rect 12041 8648 12087 8694
rect 11927 8534 11973 8580
rect 12041 8534 12087 8580
rect 11927 8420 11973 8466
rect 12041 8420 12087 8466
rect 11927 8306 11973 8352
rect 12041 8306 12087 8352
rect 11927 8192 11973 8238
rect 12041 8192 12087 8238
rect 11927 8078 11973 8124
rect 12041 8078 12087 8124
rect 11927 7964 11973 8010
rect 12041 7964 12087 8010
rect 11927 7850 11973 7896
rect 12041 7850 12087 7896
rect 11927 7736 11973 7782
rect 12041 7736 12087 7782
rect 11927 7622 11973 7668
rect 12041 7622 12087 7668
rect 11927 7508 11973 7554
rect 12041 7508 12087 7554
rect 11927 7394 11973 7440
rect 12041 7394 12087 7440
rect 11927 7280 11973 7326
rect 12041 7280 12087 7326
rect 11927 7166 11973 7212
rect 12041 7166 12087 7212
rect 11927 7052 11973 7098
rect 12041 7052 12087 7098
rect 11927 6938 11973 6984
rect 12041 6938 12087 6984
rect 11927 6824 11973 6870
rect 12041 6824 12087 6870
rect 11927 6710 11973 6756
rect 12041 6710 12087 6756
rect 11927 6596 11973 6642
rect 12041 6596 12087 6642
rect 11927 6482 11973 6528
rect 12041 6482 12087 6528
rect 11927 6368 11973 6414
rect 12041 6368 12087 6414
rect 11927 6254 11973 6300
rect 12041 6254 12087 6300
rect 11927 6140 11973 6186
rect 12041 6140 12087 6186
rect 11927 6026 11973 6072
rect 12041 6026 12087 6072
rect 11927 5912 11973 5958
rect 12041 5912 12087 5958
rect 11927 5798 11973 5844
rect 12041 5798 12087 5844
rect 11927 5684 11973 5730
rect 12041 5684 12087 5730
rect 11927 5570 11973 5616
rect 12041 5570 12087 5616
rect 11927 5456 11973 5502
rect 12041 5456 12087 5502
rect 11927 5342 11973 5388
rect 12041 5342 12087 5388
rect 1587 5000 1633 5046
rect 1701 5000 1747 5046
rect 11927 5228 11973 5274
rect 12041 5228 12087 5274
rect 11927 5114 11973 5160
rect 12041 5114 12087 5160
rect 11927 5000 11973 5046
rect 12041 5000 12087 5046
rect 1587 4886 1633 4932
rect 1701 4886 1747 4932
rect 1855 4886 1901 4932
rect 1969 4886 2015 4932
rect 2083 4886 2129 4932
rect 2197 4886 2243 4932
rect 2311 4886 2357 4932
rect 2425 4886 2471 4932
rect 2539 4886 2585 4932
rect 2653 4886 2699 4932
rect 2767 4886 2813 4932
rect 2881 4886 2927 4932
rect 2995 4886 3041 4932
rect 3109 4886 3155 4932
rect 3223 4886 3269 4932
rect 3337 4886 3383 4932
rect 3451 4886 3497 4932
rect 3565 4886 3611 4932
rect 3679 4886 3725 4932
rect 3793 4886 3839 4932
rect 3907 4886 3953 4932
rect 4021 4886 4067 4932
rect 4135 4886 4181 4932
rect 4249 4886 4295 4932
rect 4363 4886 4409 4932
rect 4477 4886 4523 4932
rect 4591 4886 4637 4932
rect 4705 4886 4751 4932
rect 4819 4886 4865 4932
rect 4933 4886 4979 4932
rect 5047 4886 5093 4932
rect 5161 4886 5207 4932
rect 5275 4886 5321 4932
rect 5389 4886 5435 4932
rect 5503 4886 5549 4932
rect 5617 4886 5663 4932
rect 5731 4886 5777 4932
rect 5845 4886 5891 4932
rect 5959 4886 6005 4932
rect 6073 4886 6119 4932
rect 6187 4886 6233 4932
rect 6301 4886 6347 4932
rect 6415 4886 6461 4932
rect 6529 4886 6575 4932
rect 6643 4886 6689 4932
rect 6757 4886 6803 4932
rect 6871 4886 6917 4932
rect 6985 4886 7031 4932
rect 7099 4886 7145 4932
rect 7213 4886 7259 4932
rect 7327 4886 7373 4932
rect 7441 4886 7487 4932
rect 7555 4886 7601 4932
rect 7669 4886 7715 4932
rect 7783 4886 7829 4932
rect 7897 4886 7943 4932
rect 8011 4886 8057 4932
rect 8125 4886 8171 4932
rect 8239 4886 8285 4932
rect 8353 4886 8399 4932
rect 8467 4886 8513 4932
rect 8581 4886 8627 4932
rect 8695 4886 8741 4932
rect 8809 4886 8855 4932
rect 8923 4886 8969 4932
rect 9037 4886 9083 4932
rect 9151 4886 9197 4932
rect 9265 4886 9311 4932
rect 9379 4886 9425 4932
rect 9493 4886 9539 4932
rect 9607 4886 9653 4932
rect 9721 4886 9767 4932
rect 9835 4886 9881 4932
rect 9949 4886 9995 4932
rect 10063 4886 10109 4932
rect 10177 4886 10223 4932
rect 10291 4886 10337 4932
rect 10405 4886 10451 4932
rect 10519 4886 10565 4932
rect 10633 4886 10679 4932
rect 10747 4886 10793 4932
rect 10861 4886 10907 4932
rect 10975 4886 11021 4932
rect 11089 4886 11135 4932
rect 11203 4886 11249 4932
rect 11317 4886 11363 4932
rect 11431 4886 11477 4932
rect 11545 4886 11591 4932
rect 11659 4886 11705 4932
rect 11773 4886 11819 4932
rect 11927 4886 11973 4932
rect 12041 4886 12087 4932
rect 1587 4772 1633 4818
rect 1701 4772 1747 4818
rect 1855 4772 1901 4818
rect 1969 4772 2015 4818
rect 2083 4772 2129 4818
rect 2197 4772 2243 4818
rect 2311 4772 2357 4818
rect 2425 4772 2471 4818
rect 2539 4772 2585 4818
rect 2653 4772 2699 4818
rect 2767 4772 2813 4818
rect 2881 4772 2927 4818
rect 2995 4772 3041 4818
rect 3109 4772 3155 4818
rect 3223 4772 3269 4818
rect 3337 4772 3383 4818
rect 3451 4772 3497 4818
rect 3565 4772 3611 4818
rect 3679 4772 3725 4818
rect 3793 4772 3839 4818
rect 3907 4772 3953 4818
rect 4021 4772 4067 4818
rect 4135 4772 4181 4818
rect 4249 4772 4295 4818
rect 4363 4772 4409 4818
rect 4477 4772 4523 4818
rect 4591 4772 4637 4818
rect 4705 4772 4751 4818
rect 4819 4772 4865 4818
rect 4933 4772 4979 4818
rect 5047 4772 5093 4818
rect 5161 4772 5207 4818
rect 5275 4772 5321 4818
rect 5389 4772 5435 4818
rect 5503 4772 5549 4818
rect 5617 4772 5663 4818
rect 5731 4772 5777 4818
rect 5845 4772 5891 4818
rect 5959 4772 6005 4818
rect 6073 4772 6119 4818
rect 6187 4772 6233 4818
rect 6301 4772 6347 4818
rect 6415 4772 6461 4818
rect 6529 4772 6575 4818
rect 6643 4772 6689 4818
rect 6757 4772 6803 4818
rect 6871 4772 6917 4818
rect 6985 4772 7031 4818
rect 7099 4772 7145 4818
rect 7213 4772 7259 4818
rect 7327 4772 7373 4818
rect 7441 4772 7487 4818
rect 7555 4772 7601 4818
rect 7669 4772 7715 4818
rect 7783 4772 7829 4818
rect 7897 4772 7943 4818
rect 8011 4772 8057 4818
rect 8125 4772 8171 4818
rect 8239 4772 8285 4818
rect 8353 4772 8399 4818
rect 8467 4772 8513 4818
rect 8581 4772 8627 4818
rect 8695 4772 8741 4818
rect 8809 4772 8855 4818
rect 8923 4772 8969 4818
rect 9037 4772 9083 4818
rect 9151 4772 9197 4818
rect 9265 4772 9311 4818
rect 9379 4772 9425 4818
rect 9493 4772 9539 4818
rect 9607 4772 9653 4818
rect 9721 4772 9767 4818
rect 9835 4772 9881 4818
rect 9949 4772 9995 4818
rect 10063 4772 10109 4818
rect 10177 4772 10223 4818
rect 10291 4772 10337 4818
rect 10405 4772 10451 4818
rect 10519 4772 10565 4818
rect 10633 4772 10679 4818
rect 10747 4772 10793 4818
rect 10861 4772 10907 4818
rect 10975 4772 11021 4818
rect 11089 4772 11135 4818
rect 11203 4772 11249 4818
rect 11317 4772 11363 4818
rect 11431 4772 11477 4818
rect 11545 4772 11591 4818
rect 11659 4772 11705 4818
rect 11773 4772 11819 4818
rect 11927 4772 11973 4818
rect 12041 4772 12087 4818
<< nsubdiffcont >>
rect -3727 17546 -3681 17592
rect -3573 17546 -3527 17592
rect -3469 17546 -3423 17592
rect -3365 17546 -3319 17592
rect -3261 17546 -3215 17592
rect -3157 17546 -3111 17592
rect -3053 17546 -3007 17592
rect -2949 17546 -2903 17592
rect -2845 17546 -2799 17592
rect -2741 17546 -2695 17592
rect -2637 17546 -2591 17592
rect -2533 17546 -2487 17592
rect -2429 17546 -2383 17592
rect -2325 17546 -2279 17592
rect -2221 17546 -2175 17592
rect -2117 17546 -2071 17592
rect -2013 17546 -1967 17592
rect -1909 17546 -1863 17592
rect -1805 17546 -1759 17592
rect -1701 17546 -1655 17592
rect -1597 17546 -1551 17592
rect -1493 17546 -1447 17592
rect -1389 17546 -1343 17592
rect -1285 17546 -1239 17592
rect -1181 17546 -1135 17592
rect -1077 17546 -1031 17592
rect -973 17546 -927 17592
rect -869 17546 -823 17592
rect -765 17546 -719 17592
rect -661 17546 -615 17592
rect -557 17546 -511 17592
rect -453 17546 -407 17592
rect -349 17546 -303 17592
rect -245 17546 -199 17592
rect -141 17546 -95 17592
rect 13 17546 59 17592
rect -3727 17442 -3681 17488
rect -3727 17338 -3681 17384
rect 13 17442 59 17488
rect 13 17338 59 17384
rect -3727 17234 -3681 17280
rect -3727 17130 -3681 17176
rect -3727 17026 -3681 17072
rect -3727 16922 -3681 16968
rect -3727 16818 -3681 16864
rect -3727 16714 -3681 16760
rect -3727 16610 -3681 16656
rect -3727 16506 -3681 16552
rect -3727 16402 -3681 16448
rect -3727 16298 -3681 16344
rect -3727 16194 -3681 16240
rect -3727 16090 -3681 16136
rect -3727 15986 -3681 16032
rect -3727 15882 -3681 15928
rect -3727 15778 -3681 15824
rect -3727 15674 -3681 15720
rect -3727 15570 -3681 15616
rect -3727 15466 -3681 15512
rect -3727 15362 -3681 15408
rect -3727 15258 -3681 15304
rect -3727 15154 -3681 15200
rect -3727 15050 -3681 15096
rect -3727 14946 -3681 14992
rect -3727 14842 -3681 14888
rect -3727 14738 -3681 14784
rect -3727 14634 -3681 14680
rect -3727 14530 -3681 14576
rect -3727 14426 -3681 14472
rect -3727 14322 -3681 14368
rect -3727 14218 -3681 14264
rect -3727 14114 -3681 14160
rect -3727 14010 -3681 14056
rect -3727 13906 -3681 13952
rect -3727 13802 -3681 13848
rect -3727 13698 -3681 13744
rect -3727 13594 -3681 13640
rect -3727 13490 -3681 13536
rect -3727 13386 -3681 13432
rect -3727 13282 -3681 13328
rect -3727 13178 -3681 13224
rect -3727 13074 -3681 13120
rect -3727 12970 -3681 13016
rect -3727 12866 -3681 12912
rect -3727 12762 -3681 12808
rect -3727 12658 -3681 12704
rect -3727 12554 -3681 12600
rect -3727 12450 -3681 12496
rect -3727 12346 -3681 12392
rect -3727 12242 -3681 12288
rect -3727 12138 -3681 12184
rect -3727 12034 -3681 12080
rect -3727 11930 -3681 11976
rect -3727 11826 -3681 11872
rect -3727 11722 -3681 11768
rect -3727 11618 -3681 11664
rect -3727 11514 -3681 11560
rect -3727 11410 -3681 11456
rect -3727 11306 -3681 11352
rect -3727 11202 -3681 11248
rect -3727 11098 -3681 11144
rect -3727 10994 -3681 11040
rect -3727 10890 -3681 10936
rect -3727 10786 -3681 10832
rect -3727 10682 -3681 10728
rect -3727 10578 -3681 10624
rect -3727 10474 -3681 10520
rect -3727 10370 -3681 10416
rect -3727 10266 -3681 10312
rect -3727 10162 -3681 10208
rect -3727 10058 -3681 10104
rect -3727 9954 -3681 10000
rect -3727 9850 -3681 9896
rect -3727 9746 -3681 9792
rect -3727 9642 -3681 9688
rect -3727 9538 -3681 9584
rect -3727 9434 -3681 9480
rect -3727 9330 -3681 9376
rect -3727 9226 -3681 9272
rect -3727 9122 -3681 9168
rect -3727 9018 -3681 9064
rect -3727 8914 -3681 8960
rect -3727 8810 -3681 8856
rect -3727 8706 -3681 8752
rect -3727 8602 -3681 8648
rect -3727 8498 -3681 8544
rect -3727 8394 -3681 8440
rect -3727 8290 -3681 8336
rect -3727 8186 -3681 8232
rect -3727 8082 -3681 8128
rect -3727 7978 -3681 8024
rect -3727 7874 -3681 7920
rect -3727 7770 -3681 7816
rect -3727 7666 -3681 7712
rect -3727 7562 -3681 7608
rect -3727 7458 -3681 7504
rect -3727 7354 -3681 7400
rect -3727 7250 -3681 7296
rect -3727 7146 -3681 7192
rect -3727 7042 -3681 7088
rect -3727 6938 -3681 6984
rect -3727 6834 -3681 6880
rect -3727 6730 -3681 6776
rect -3727 6626 -3681 6672
rect -3727 6522 -3681 6568
rect -3727 6418 -3681 6464
rect -3727 6314 -3681 6360
rect -3727 6210 -3681 6256
rect -3727 6106 -3681 6152
rect -3727 6002 -3681 6048
rect -3727 5898 -3681 5944
rect -3727 5794 -3681 5840
rect -3727 5690 -3681 5736
rect -3727 5586 -3681 5632
rect -3727 5482 -3681 5528
rect -3727 5378 -3681 5424
rect -3727 5274 -3681 5320
rect -3727 5170 -3681 5216
rect -3727 5066 -3681 5112
rect -3727 4962 -3681 5008
rect -3727 4858 -3681 4904
rect -3727 4754 -3681 4800
rect -3727 4650 -3681 4696
rect -3727 4546 -3681 4592
rect -3727 4442 -3681 4488
rect -3727 4338 -3681 4384
rect 13 17234 59 17280
rect 13 17130 59 17176
rect 13 17026 59 17072
rect 13 16922 59 16968
rect 13 16818 59 16864
rect 13 16714 59 16760
rect 13 16610 59 16656
rect 13 16506 59 16552
rect 13 16402 59 16448
rect 13 16298 59 16344
rect 13 16194 59 16240
rect 13 16090 59 16136
rect 13 15986 59 16032
rect 13 15882 59 15928
rect 13 15778 59 15824
rect 13 15674 59 15720
rect 13 15570 59 15616
rect 13 15466 59 15512
rect 13 15362 59 15408
rect 13 15258 59 15304
rect 13 15154 59 15200
rect 13 15050 59 15096
rect 13 14946 59 14992
rect 13 14842 59 14888
rect 13 14738 59 14784
rect 13 14634 59 14680
rect 13 14530 59 14576
rect 13 14426 59 14472
rect 13 14322 59 14368
rect 13 14218 59 14264
rect 13 14114 59 14160
rect 13 14010 59 14056
rect 13 13906 59 13952
rect 13 13802 59 13848
rect 13 13698 59 13744
rect 13 13594 59 13640
rect 13 13490 59 13536
rect 13 13386 59 13432
rect 13 13282 59 13328
rect 13 13178 59 13224
rect 13 13074 59 13120
rect 13 12970 59 13016
rect 13 12866 59 12912
rect 13 12762 59 12808
rect 13 12658 59 12704
rect 13 12554 59 12600
rect 13 12450 59 12496
rect 13 12346 59 12392
rect 13 12242 59 12288
rect 13 12138 59 12184
rect 13 12034 59 12080
rect 13 11930 59 11976
rect 13 11826 59 11872
rect 13 11722 59 11768
rect 13 11618 59 11664
rect 13 11514 59 11560
rect 13 11410 59 11456
rect 13 11306 59 11352
rect 13 11202 59 11248
rect 13 11098 59 11144
rect 13 10994 59 11040
rect 13 10890 59 10936
rect 13 10786 59 10832
rect 13 10682 59 10728
rect 13 10578 59 10624
rect 13 10474 59 10520
rect 13 10370 59 10416
rect 13 10266 59 10312
rect 13 10162 59 10208
rect 13 10058 59 10104
rect 13 9954 59 10000
rect 13 9850 59 9896
rect 13 9746 59 9792
rect 13 9642 59 9688
rect 13 9538 59 9584
rect 13 9434 59 9480
rect 13 9330 59 9376
rect 13 9226 59 9272
rect 13 9122 59 9168
rect 13 9018 59 9064
rect 13 8914 59 8960
rect 13 8810 59 8856
rect 13 8706 59 8752
rect 13 8602 59 8648
rect 13 8498 59 8544
rect 13 8394 59 8440
rect 13 8290 59 8336
rect 13 8186 59 8232
rect 13 8082 59 8128
rect 13 7978 59 8024
rect 13 7874 59 7920
rect 13 7770 59 7816
rect 13 7666 59 7712
rect 13 7562 59 7608
rect 13 7458 59 7504
rect 13 7354 59 7400
rect 13 7250 59 7296
rect 13 7146 59 7192
rect 13 7042 59 7088
rect 13 6938 59 6984
rect 13 6834 59 6880
rect 13 6730 59 6776
rect 13 6626 59 6672
rect 13 6522 59 6568
rect 13 6418 59 6464
rect 13 6314 59 6360
rect 13 6210 59 6256
rect 13 6106 59 6152
rect 13 6002 59 6048
rect 13 5898 59 5944
rect 13 5794 59 5840
rect 13 5690 59 5736
rect 13 5586 59 5632
rect 13 5482 59 5528
rect 13 5378 59 5424
rect 13 5274 59 5320
rect 13 5170 59 5216
rect 13 5066 59 5112
rect 13 4962 59 5008
rect 13 4858 59 4904
rect 13 4754 59 4800
rect 13 4650 59 4696
rect 13 4546 59 4592
rect -3727 4234 -3681 4280
rect -3727 4130 -3681 4176
rect 13 4130 59 4176
rect -3727 4026 -3681 4072
rect -3573 4026 -3527 4072
rect -3469 4026 -3423 4072
rect -3365 4026 -3319 4072
rect -3261 4026 -3215 4072
rect -3157 4026 -3111 4072
rect -3053 4026 -3007 4072
rect -2949 4026 -2903 4072
rect -2845 4026 -2799 4072
rect -2741 4026 -2695 4072
rect -2637 4026 -2591 4072
rect -2533 4026 -2487 4072
rect -2429 4026 -2383 4072
rect -2325 4026 -2279 4072
rect -2221 4026 -2175 4072
rect -2117 4026 -2071 4072
rect -2013 4026 -1967 4072
rect -1909 4026 -1863 4072
rect -1805 4026 -1759 4072
rect -1701 4026 -1655 4072
rect -1597 4026 -1551 4072
rect -1493 4026 -1447 4072
rect -1389 4026 -1343 4072
rect -1285 4026 -1239 4072
rect -1181 4026 -1135 4072
rect -1077 4026 -1031 4072
rect -973 4026 -927 4072
rect -869 4026 -823 4072
rect -765 4026 -719 4072
rect -661 4026 -615 4072
rect -557 4026 -511 4072
rect -453 4026 -407 4072
rect -349 4026 -303 4072
rect -245 4026 -199 4072
rect -141 4026 -95 4072
rect 13 4026 59 4072
<< mvnmoscap >>
rect 2180 11351 4180 16351
rect 4616 11351 6616 16351
rect 7052 11351 9052 16351
rect 9488 11351 11488 16351
rect 2180 5339 4180 10339
rect 4616 5339 6616 10339
rect 7052 5339 9052 10339
rect 9488 5339 11488 10339
<< polysilicon >>
rect -3454 17287 -3294 17300
rect -3454 17241 -3397 17287
rect -3351 17241 -3294 17287
rect -3454 17198 -3294 17241
rect -3454 4384 -3294 4427
rect -3454 4338 -3397 4384
rect -3351 4338 -3294 4384
rect -3454 4325 -3294 4338
rect -3174 17287 -3014 17300
rect -3174 17241 -3117 17287
rect -3071 17241 -3014 17287
rect -3174 17198 -3014 17241
rect -3174 4384 -3014 4427
rect -3174 4338 -3117 4384
rect -3071 4338 -3014 4384
rect -3174 4325 -3014 4338
rect -2894 17287 -2734 17300
rect -2894 17241 -2837 17287
rect -2791 17241 -2734 17287
rect -2894 17198 -2734 17241
rect -2894 4384 -2734 4427
rect -2894 4338 -2837 4384
rect -2791 4338 -2734 4384
rect -2894 4325 -2734 4338
rect -2614 17287 -2454 17300
rect -2614 17241 -2557 17287
rect -2511 17241 -2454 17287
rect -2614 17198 -2454 17241
rect -2614 4384 -2454 4427
rect -2614 4338 -2557 4384
rect -2511 4338 -2454 4384
rect -2614 4325 -2454 4338
rect -2334 17287 -2174 17300
rect -2334 17241 -2277 17287
rect -2231 17241 -2174 17287
rect -2334 17198 -2174 17241
rect -2334 4384 -2174 4427
rect -2334 4338 -2277 4384
rect -2231 4338 -2174 4384
rect -2334 4325 -2174 4338
rect -2054 17287 -1894 17300
rect -2054 17241 -1997 17287
rect -1951 17241 -1894 17287
rect -2054 17198 -1894 17241
rect -2054 4384 -1894 4427
rect -2054 4338 -1997 4384
rect -1951 4338 -1894 4384
rect -2054 4325 -1894 4338
rect -1774 17287 -1614 17300
rect -1774 17241 -1717 17287
rect -1671 17241 -1614 17287
rect -1774 17198 -1614 17241
rect -1774 4384 -1614 4427
rect -1774 4338 -1717 4384
rect -1671 4338 -1614 4384
rect -1774 4325 -1614 4338
rect -1494 17287 -1334 17300
rect -1494 17241 -1437 17287
rect -1391 17241 -1334 17287
rect -1494 17198 -1334 17241
rect -1494 4384 -1334 4427
rect -1494 4338 -1437 4384
rect -1391 4338 -1334 4384
rect -1494 4325 -1334 4338
rect -1214 17287 -1054 17300
rect -1214 17241 -1157 17287
rect -1111 17241 -1054 17287
rect -1214 17198 -1054 17241
rect -1214 4384 -1054 4427
rect -1214 4338 -1157 4384
rect -1111 4338 -1054 4384
rect -1214 4325 -1054 4338
rect -934 17287 -774 17300
rect -934 17241 -877 17287
rect -831 17241 -774 17287
rect -934 17198 -774 17241
rect -934 4384 -774 4427
rect -934 4338 -877 4384
rect -831 4338 -774 4384
rect -934 4325 -774 4338
rect -654 17287 -494 17300
rect -654 17241 -597 17287
rect -551 17241 -494 17287
rect -654 17198 -494 17241
rect -654 4384 -494 4427
rect -654 4338 -597 4384
rect -551 4338 -494 4384
rect -654 4325 -494 4338
rect -374 17287 -214 17300
rect -374 17241 -317 17287
rect -271 17241 -214 17287
rect -374 17198 -214 17241
rect -374 4384 -214 4427
rect -374 4338 -317 4384
rect -271 4338 -214 4384
rect -374 4325 -214 4338
rect 2180 16430 4180 16443
rect 2180 16384 2233 16430
rect 4127 16384 4180 16430
rect 2180 16351 4180 16384
rect 4616 16430 6616 16443
rect 4616 16384 4669 16430
rect 6563 16384 6616 16430
rect 4616 16351 6616 16384
rect 7052 16430 9052 16443
rect 7052 16384 7105 16430
rect 8999 16384 9052 16430
rect 7052 16351 9052 16384
rect 9488 16430 11488 16443
rect 9488 16384 9541 16430
rect 11435 16384 11488 16430
rect 9488 16351 11488 16384
rect 2180 11318 4180 11351
rect 2180 11272 2233 11318
rect 4127 11272 4180 11318
rect 2180 11259 4180 11272
rect 4616 11318 6616 11351
rect 4616 11272 4669 11318
rect 6563 11272 6616 11318
rect 4616 11259 6616 11272
rect 7052 11318 9052 11351
rect 7052 11272 7105 11318
rect 8999 11272 9052 11318
rect 7052 11259 9052 11272
rect 9488 11318 11488 11351
rect 9488 11272 9541 11318
rect 11435 11272 11488 11318
rect 9488 11259 11488 11272
rect 2180 10418 4180 10431
rect 2180 10372 2233 10418
rect 4127 10372 4180 10418
rect 2180 10339 4180 10372
rect 4616 10418 6616 10431
rect 4616 10372 4669 10418
rect 6563 10372 6616 10418
rect 4616 10339 6616 10372
rect 7052 10418 9052 10431
rect 7052 10372 7105 10418
rect 8999 10372 9052 10418
rect 7052 10339 9052 10372
rect 9488 10418 11488 10431
rect 9488 10372 9541 10418
rect 11435 10372 11488 10418
rect 9488 10339 11488 10372
rect 2180 5306 4180 5339
rect 2180 5260 2233 5306
rect 4127 5260 4180 5306
rect 2180 5247 4180 5260
rect 4616 5306 6616 5339
rect 4616 5260 4669 5306
rect 6563 5260 6616 5306
rect 4616 5247 6616 5260
rect 7052 5306 9052 5339
rect 7052 5260 7105 5306
rect 8999 5260 9052 5306
rect 7052 5247 9052 5260
rect 9488 5306 11488 5339
rect 9488 5260 9541 5306
rect 11435 5260 11488 5306
rect 9488 5247 11488 5260
<< polycontact >>
rect -3397 17241 -3351 17287
rect -3397 4338 -3351 4384
rect -3117 17241 -3071 17287
rect -3117 4338 -3071 4384
rect -2837 17241 -2791 17287
rect -2837 4338 -2791 4384
rect -2557 17241 -2511 17287
rect -2557 4338 -2511 4384
rect -2277 17241 -2231 17287
rect -2277 4338 -2231 4384
rect -1997 17241 -1951 17287
rect -1997 4338 -1951 4384
rect -1717 17241 -1671 17287
rect -1717 4338 -1671 4384
rect -1437 17241 -1391 17287
rect -1437 4338 -1391 4384
rect -1157 17241 -1111 17287
rect -1157 4338 -1111 4384
rect -877 17241 -831 17287
rect -877 4338 -831 4384
rect -597 17241 -551 17287
rect -597 4338 -551 4384
rect -317 17241 -271 17287
rect -317 4338 -271 4384
rect 2233 16384 4127 16430
rect 4669 16384 6563 16430
rect 7105 16384 8999 16430
rect 9541 16384 11435 16430
rect 2233 11272 4127 11318
rect 4669 11272 6563 11318
rect 7105 11272 8999 11318
rect 9541 11272 11435 11318
rect 2233 10372 4127 10418
rect 4669 10372 6563 10418
rect 7105 10372 8999 10418
rect 9541 10372 11435 10418
rect 2233 5260 4127 5306
rect 4669 5260 6563 5306
rect 7105 5260 8999 5306
rect 9541 5260 11435 5306
<< ppolyres >>
rect -3454 4427 -3294 17198
rect -3174 4427 -3014 17198
rect -2894 4427 -2734 17198
rect -2614 4427 -2454 17198
rect -2334 4427 -2174 17198
rect -2054 4427 -1894 17198
rect -1774 4427 -1614 17198
rect -1494 4427 -1334 17198
rect -1214 4427 -1054 17198
rect -934 4427 -774 17198
rect -654 4427 -494 17198
rect -374 4427 -214 17198
<< metal1 >>
rect -3742 17592 74 17603
rect -3742 17546 -3727 17592
rect -3681 17546 -3573 17592
rect -3527 17546 -3469 17592
rect -3423 17546 -3365 17592
rect -3319 17546 -3261 17592
rect -3215 17546 -3157 17592
rect -3111 17546 -3053 17592
rect -3007 17546 -2949 17592
rect -2903 17546 -2845 17592
rect -2799 17546 -2741 17592
rect -2695 17546 -2637 17592
rect -2591 17546 -2533 17592
rect -2487 17546 -2429 17592
rect -2383 17546 -2325 17592
rect -2279 17546 -2221 17592
rect -2175 17546 -2117 17592
rect -2071 17546 -2013 17592
rect -1967 17546 -1909 17592
rect -1863 17546 -1805 17592
rect -1759 17546 -1701 17592
rect -1655 17546 -1597 17592
rect -1551 17546 -1493 17592
rect -1447 17546 -1389 17592
rect -1343 17546 -1285 17592
rect -1239 17546 -1181 17592
rect -1135 17546 -1077 17592
rect -1031 17546 -973 17592
rect -927 17546 -869 17592
rect -823 17546 -765 17592
rect -719 17546 -661 17592
rect -615 17546 -557 17592
rect -511 17546 -453 17592
rect -407 17546 -349 17592
rect -303 17546 -245 17592
rect -199 17546 -141 17592
rect -95 17546 13 17592
rect 59 17546 74 17592
rect -3742 17535 74 17546
rect -3742 17488 -3666 17535
rect -3742 17442 -3727 17488
rect -3681 17442 -3666 17488
rect -3742 17384 -3666 17442
rect -3742 17338 -3727 17384
rect -3681 17338 -3666 17384
rect -3742 17280 -3666 17338
rect -2 17488 74 17535
rect -2 17442 13 17488
rect 59 17442 74 17488
rect -2 17384 74 17442
rect -2 17338 13 17384
rect 59 17338 74 17384
rect -3742 17234 -3727 17280
rect -3681 17234 -3666 17280
rect -3742 17176 -3666 17234
rect -3452 17287 -3016 17298
rect -3452 17241 -3397 17287
rect -3351 17241 -3117 17287
rect -3071 17241 -3016 17287
rect -3452 17230 -3016 17241
rect -2892 17287 -2456 17298
rect -2892 17241 -2837 17287
rect -2791 17241 -2557 17287
rect -2511 17241 -2456 17287
rect -2892 17230 -2456 17241
rect -2332 17287 -1896 17298
rect -2332 17241 -2277 17287
rect -2231 17241 -1997 17287
rect -1951 17241 -1896 17287
rect -2332 17230 -1896 17241
rect -1772 17287 -1336 17298
rect -1772 17241 -1717 17287
rect -1671 17241 -1437 17287
rect -1391 17241 -1336 17287
rect -1772 17230 -1336 17241
rect -1212 17287 -776 17298
rect -1212 17241 -1157 17287
rect -1111 17241 -877 17287
rect -831 17241 -776 17287
rect -1212 17230 -776 17241
rect -652 17287 -216 17298
rect -652 17241 -597 17287
rect -551 17241 -317 17287
rect -271 17241 -216 17287
rect -652 17230 -216 17241
rect -2 17280 74 17338
rect -2 17234 13 17280
rect 59 17234 74 17280
rect -3742 17130 -3727 17176
rect -3681 17130 -3666 17176
rect -3742 17072 -3666 17130
rect -3742 17026 -3727 17072
rect -3681 17026 -3666 17072
rect -3742 16968 -3666 17026
rect -3742 16922 -3727 16968
rect -3681 16922 -3666 16968
rect -3742 16864 -3666 16922
rect -3742 16818 -3727 16864
rect -3681 16818 -3666 16864
rect -3742 16760 -3666 16818
rect -3742 16714 -3727 16760
rect -3681 16714 -3666 16760
rect -3742 16656 -3666 16714
rect -3742 16610 -3727 16656
rect -3681 16610 -3666 16656
rect -3742 16552 -3666 16610
rect -3742 16506 -3727 16552
rect -3681 16506 -3666 16552
rect -3742 16448 -3666 16506
rect -3742 16402 -3727 16448
rect -3681 16402 -3666 16448
rect -3742 16344 -3666 16402
rect -3742 16298 -3727 16344
rect -3681 16298 -3666 16344
rect -3742 16240 -3666 16298
rect -3742 16194 -3727 16240
rect -3681 16194 -3666 16240
rect -3742 16136 -3666 16194
rect -3742 16090 -3727 16136
rect -3681 16090 -3666 16136
rect -3742 16032 -3666 16090
rect -3742 15986 -3727 16032
rect -3681 15986 -3666 16032
rect -3742 15928 -3666 15986
rect -3742 15882 -3727 15928
rect -3681 15882 -3666 15928
rect -3742 15824 -3666 15882
rect -3742 15778 -3727 15824
rect -3681 15778 -3666 15824
rect -3742 15720 -3666 15778
rect -3742 15674 -3727 15720
rect -3681 15674 -3666 15720
rect -3742 15616 -3666 15674
rect -3742 15570 -3727 15616
rect -3681 15570 -3666 15616
rect -3742 15512 -3666 15570
rect -3742 15466 -3727 15512
rect -3681 15466 -3666 15512
rect -3742 15408 -3666 15466
rect -3742 15362 -3727 15408
rect -3681 15362 -3666 15408
rect -3742 15304 -3666 15362
rect -3742 15258 -3727 15304
rect -3681 15258 -3666 15304
rect -3742 15200 -3666 15258
rect -3742 15154 -3727 15200
rect -3681 15154 -3666 15200
rect -3742 15096 -3666 15154
rect -3742 15050 -3727 15096
rect -3681 15050 -3666 15096
rect -3742 14992 -3666 15050
rect -3742 14946 -3727 14992
rect -3681 14946 -3666 14992
rect -3742 14888 -3666 14946
rect -3742 14842 -3727 14888
rect -3681 14842 -3666 14888
rect -3742 14784 -3666 14842
rect -3742 14738 -3727 14784
rect -3681 14738 -3666 14784
rect -3742 14680 -3666 14738
rect -3742 14634 -3727 14680
rect -3681 14634 -3666 14680
rect -3742 14576 -3666 14634
rect -3742 14530 -3727 14576
rect -3681 14530 -3666 14576
rect -3742 14472 -3666 14530
rect -3742 14426 -3727 14472
rect -3681 14426 -3666 14472
rect -3742 14368 -3666 14426
rect -3742 14322 -3727 14368
rect -3681 14322 -3666 14368
rect -3742 14264 -3666 14322
rect -3742 14218 -3727 14264
rect -3681 14218 -3666 14264
rect -3742 14160 -3666 14218
rect -3742 14114 -3727 14160
rect -3681 14114 -3666 14160
rect -3742 14056 -3666 14114
rect -3742 14010 -3727 14056
rect -3681 14010 -3666 14056
rect -3742 13952 -3666 14010
rect -3742 13906 -3727 13952
rect -3681 13906 -3666 13952
rect -3742 13848 -3666 13906
rect -3742 13802 -3727 13848
rect -3681 13802 -3666 13848
rect -3742 13744 -3666 13802
rect -3742 13698 -3727 13744
rect -3681 13698 -3666 13744
rect -3742 13640 -3666 13698
rect -3742 13594 -3727 13640
rect -3681 13594 -3666 13640
rect -3742 13536 -3666 13594
rect -3742 13490 -3727 13536
rect -3681 13490 -3666 13536
rect -3742 13432 -3666 13490
rect -3742 13386 -3727 13432
rect -3681 13386 -3666 13432
rect -3742 13328 -3666 13386
rect -3742 13282 -3727 13328
rect -3681 13282 -3666 13328
rect -3742 13224 -3666 13282
rect -3742 13178 -3727 13224
rect -3681 13178 -3666 13224
rect -3742 13120 -3666 13178
rect -3742 13074 -3727 13120
rect -3681 13074 -3666 13120
rect -3742 13016 -3666 13074
rect -3742 12970 -3727 13016
rect -3681 12970 -3666 13016
rect -3742 12912 -3666 12970
rect -3742 12866 -3727 12912
rect -3681 12866 -3666 12912
rect -3742 12808 -3666 12866
rect -3742 12762 -3727 12808
rect -3681 12762 -3666 12808
rect -3742 12704 -3666 12762
rect -3742 12658 -3727 12704
rect -3681 12658 -3666 12704
rect -3742 12600 -3666 12658
rect -3742 12554 -3727 12600
rect -3681 12554 -3666 12600
rect -3742 12496 -3666 12554
rect -3742 12450 -3727 12496
rect -3681 12450 -3666 12496
rect -3742 12392 -3666 12450
rect -3742 12346 -3727 12392
rect -3681 12346 -3666 12392
rect -3742 12288 -3666 12346
rect -3742 12242 -3727 12288
rect -3681 12242 -3666 12288
rect -3742 12184 -3666 12242
rect -3742 12138 -3727 12184
rect -3681 12138 -3666 12184
rect -3742 12080 -3666 12138
rect -3742 12034 -3727 12080
rect -3681 12034 -3666 12080
rect -3742 11976 -3666 12034
rect -3742 11930 -3727 11976
rect -3681 11930 -3666 11976
rect -3742 11872 -3666 11930
rect -3742 11826 -3727 11872
rect -3681 11826 -3666 11872
rect -3742 11768 -3666 11826
rect -3742 11722 -3727 11768
rect -3681 11722 -3666 11768
rect -3742 11664 -3666 11722
rect -3742 11618 -3727 11664
rect -3681 11618 -3666 11664
rect -3742 11560 -3666 11618
rect -3742 11514 -3727 11560
rect -3681 11514 -3666 11560
rect -3742 11456 -3666 11514
rect -3742 11410 -3727 11456
rect -3681 11410 -3666 11456
rect -3742 11352 -3666 11410
rect -3742 11306 -3727 11352
rect -3681 11306 -3666 11352
rect -3742 11248 -3666 11306
rect -3742 11202 -3727 11248
rect -3681 11202 -3666 11248
rect -3742 11144 -3666 11202
rect -3742 11098 -3727 11144
rect -3681 11098 -3666 11144
rect -3742 11040 -3666 11098
rect -3742 10994 -3727 11040
rect -3681 10994 -3666 11040
rect -3742 10936 -3666 10994
rect -3742 10890 -3727 10936
rect -3681 10890 -3666 10936
rect -3742 10832 -3666 10890
rect -3742 10786 -3727 10832
rect -3681 10786 -3666 10832
rect -3742 10728 -3666 10786
rect -3742 10682 -3727 10728
rect -3681 10682 -3666 10728
rect -3742 10624 -3666 10682
rect -3742 10578 -3727 10624
rect -3681 10578 -3666 10624
rect -3742 10520 -3666 10578
rect -3742 10474 -3727 10520
rect -3681 10474 -3666 10520
rect -3742 10416 -3666 10474
rect -3742 10370 -3727 10416
rect -3681 10370 -3666 10416
rect -3742 10312 -3666 10370
rect -3742 10266 -3727 10312
rect -3681 10266 -3666 10312
rect -3742 10208 -3666 10266
rect -3742 10162 -3727 10208
rect -3681 10162 -3666 10208
rect -3742 10104 -3666 10162
rect -3742 10058 -3727 10104
rect -3681 10058 -3666 10104
rect -3742 10000 -3666 10058
rect -3742 9954 -3727 10000
rect -3681 9954 -3666 10000
rect -3742 9896 -3666 9954
rect -3742 9850 -3727 9896
rect -3681 9850 -3666 9896
rect -3742 9792 -3666 9850
rect -3742 9746 -3727 9792
rect -3681 9746 -3666 9792
rect -3742 9688 -3666 9746
rect -3742 9642 -3727 9688
rect -3681 9642 -3666 9688
rect -3742 9584 -3666 9642
rect -3742 9538 -3727 9584
rect -3681 9538 -3666 9584
rect -3742 9480 -3666 9538
rect -3742 9434 -3727 9480
rect -3681 9434 -3666 9480
rect -3742 9376 -3666 9434
rect -3742 9330 -3727 9376
rect -3681 9330 -3666 9376
rect -3742 9272 -3666 9330
rect -3742 9226 -3727 9272
rect -3681 9226 -3666 9272
rect -3742 9168 -3666 9226
rect -3742 9122 -3727 9168
rect -3681 9122 -3666 9168
rect -3742 9064 -3666 9122
rect -3742 9018 -3727 9064
rect -3681 9018 -3666 9064
rect -3742 8960 -3666 9018
rect -3742 8914 -3727 8960
rect -3681 8914 -3666 8960
rect -3742 8856 -3666 8914
rect -3742 8810 -3727 8856
rect -3681 8810 -3666 8856
rect -3742 8752 -3666 8810
rect -3742 8706 -3727 8752
rect -3681 8706 -3666 8752
rect -3742 8648 -3666 8706
rect -3742 8602 -3727 8648
rect -3681 8602 -3666 8648
rect -3742 8544 -3666 8602
rect -3742 8498 -3727 8544
rect -3681 8498 -3666 8544
rect -3742 8440 -3666 8498
rect -3742 8394 -3727 8440
rect -3681 8394 -3666 8440
rect -3742 8336 -3666 8394
rect -3742 8290 -3727 8336
rect -3681 8290 -3666 8336
rect -3742 8232 -3666 8290
rect -3742 8186 -3727 8232
rect -3681 8186 -3666 8232
rect -3742 8128 -3666 8186
rect -3742 8082 -3727 8128
rect -3681 8082 -3666 8128
rect -3742 8024 -3666 8082
rect -3742 7978 -3727 8024
rect -3681 7978 -3666 8024
rect -3742 7920 -3666 7978
rect -3742 7874 -3727 7920
rect -3681 7874 -3666 7920
rect -3742 7816 -3666 7874
rect -3742 7770 -3727 7816
rect -3681 7770 -3666 7816
rect -3742 7712 -3666 7770
rect -3742 7666 -3727 7712
rect -3681 7666 -3666 7712
rect -3742 7608 -3666 7666
rect -3742 7562 -3727 7608
rect -3681 7562 -3666 7608
rect -3742 7504 -3666 7562
rect -3742 7458 -3727 7504
rect -3681 7458 -3666 7504
rect -3742 7400 -3666 7458
rect -3742 7354 -3727 7400
rect -3681 7354 -3666 7400
rect -3742 7296 -3666 7354
rect -3742 7250 -3727 7296
rect -3681 7250 -3666 7296
rect -3742 7192 -3666 7250
rect -3742 7146 -3727 7192
rect -3681 7146 -3666 7192
rect -3742 7088 -3666 7146
rect -3742 7042 -3727 7088
rect -3681 7042 -3666 7088
rect -3742 6984 -3666 7042
rect -3742 6938 -3727 6984
rect -3681 6938 -3666 6984
rect -3742 6880 -3666 6938
rect -3742 6834 -3727 6880
rect -3681 6834 -3666 6880
rect -3742 6776 -3666 6834
rect -3742 6730 -3727 6776
rect -3681 6730 -3666 6776
rect -3742 6672 -3666 6730
rect -3742 6626 -3727 6672
rect -3681 6626 -3666 6672
rect -3742 6568 -3666 6626
rect -3742 6522 -3727 6568
rect -3681 6522 -3666 6568
rect -3742 6464 -3666 6522
rect -3742 6418 -3727 6464
rect -3681 6418 -3666 6464
rect -3742 6360 -3666 6418
rect -3742 6314 -3727 6360
rect -3681 6314 -3666 6360
rect -3742 6256 -3666 6314
rect -3742 6210 -3727 6256
rect -3681 6210 -3666 6256
rect -3742 6152 -3666 6210
rect -3742 6106 -3727 6152
rect -3681 6106 -3666 6152
rect -3742 6048 -3666 6106
rect -3742 6002 -3727 6048
rect -3681 6002 -3666 6048
rect -3742 5944 -3666 6002
rect -3742 5898 -3727 5944
rect -3681 5898 -3666 5944
rect -3742 5840 -3666 5898
rect -3742 5794 -3727 5840
rect -3681 5794 -3666 5840
rect -3742 5736 -3666 5794
rect -3742 5690 -3727 5736
rect -3681 5690 -3666 5736
rect -3742 5632 -3666 5690
rect -3742 5586 -3727 5632
rect -3681 5586 -3666 5632
rect -3742 5528 -3666 5586
rect -3742 5482 -3727 5528
rect -3681 5482 -3666 5528
rect -3742 5424 -3666 5482
rect -3742 5378 -3727 5424
rect -3681 5378 -3666 5424
rect -3742 5320 -3666 5378
rect -3742 5274 -3727 5320
rect -3681 5274 -3666 5320
rect -3742 5216 -3666 5274
rect -3742 5170 -3727 5216
rect -3681 5170 -3666 5216
rect -3742 5112 -3666 5170
rect -3742 5066 -3727 5112
rect -3681 5066 -3666 5112
rect -3742 5008 -3666 5066
rect -3742 4962 -3727 5008
rect -3681 4962 -3666 5008
rect -3742 4904 -3666 4962
rect -3742 4858 -3727 4904
rect -3681 4858 -3666 4904
rect -3742 4800 -3666 4858
rect -3742 4754 -3727 4800
rect -3681 4754 -3666 4800
rect -3742 4696 -3666 4754
rect -3742 4650 -3727 4696
rect -3681 4650 -3666 4696
rect -3742 4592 -3666 4650
rect -3742 4546 -3727 4592
rect -3681 4546 -3666 4592
rect -3742 4488 -3666 4546
rect -3742 4442 -3727 4488
rect -3681 4442 -3666 4488
rect -2 17176 74 17234
rect -2 17130 13 17176
rect 59 17130 74 17176
rect -2 17072 74 17130
rect -2 17026 13 17072
rect 59 17026 74 17072
rect -2 16968 74 17026
rect -2 16922 13 16968
rect 59 16922 74 16968
rect -2 16864 74 16922
rect -2 16818 13 16864
rect 59 16818 74 16864
rect -2 16760 74 16818
rect -2 16714 13 16760
rect 59 16714 74 16760
rect -2 16656 74 16714
rect 1576 17016 12098 17028
rect 1576 16970 1587 17016
rect 1633 16970 1701 17016
rect 1747 16970 1855 17016
rect 1901 16970 1969 17016
rect 2015 16970 2083 17016
rect 2129 16970 2197 17016
rect 2243 16970 2311 17016
rect 2357 16970 2425 17016
rect 2471 16970 2539 17016
rect 2585 16970 2653 17016
rect 2699 16970 2767 17016
rect 2813 16970 2881 17016
rect 2927 16970 2995 17016
rect 3041 16970 3109 17016
rect 3155 16970 3223 17016
rect 3269 16970 3337 17016
rect 3383 16970 3451 17016
rect 3497 16970 3565 17016
rect 3611 16970 3679 17016
rect 3725 16970 3793 17016
rect 3839 16970 3907 17016
rect 3953 16970 4021 17016
rect 4067 16970 4135 17016
rect 4181 16970 4249 17016
rect 4295 16970 4363 17016
rect 4409 16970 4477 17016
rect 4523 16970 4591 17016
rect 4637 16970 4705 17016
rect 4751 16970 4819 17016
rect 4865 16970 4933 17016
rect 4979 16970 5047 17016
rect 5093 16970 5161 17016
rect 5207 16970 5275 17016
rect 5321 16970 5389 17016
rect 5435 16970 5503 17016
rect 5549 16970 5617 17016
rect 5663 16970 5731 17016
rect 5777 16970 5845 17016
rect 5891 16970 5959 17016
rect 6005 16970 6073 17016
rect 6119 16970 6187 17016
rect 6233 16970 6301 17016
rect 6347 16970 6415 17016
rect 6461 16970 6529 17016
rect 6575 16970 6643 17016
rect 6689 16970 6757 17016
rect 6803 16970 6871 17016
rect 6917 16970 6985 17016
rect 7031 16970 7099 17016
rect 7145 16970 7213 17016
rect 7259 16970 7327 17016
rect 7373 16970 7441 17016
rect 7487 16970 7555 17016
rect 7601 16970 7669 17016
rect 7715 16970 7783 17016
rect 7829 16970 7897 17016
rect 7943 16970 8011 17016
rect 8057 16970 8125 17016
rect 8171 16970 8239 17016
rect 8285 16970 8353 17016
rect 8399 16970 8467 17016
rect 8513 16970 8581 17016
rect 8627 16970 8695 17016
rect 8741 16970 8809 17016
rect 8855 16970 8923 17016
rect 8969 16970 9037 17016
rect 9083 16970 9151 17016
rect 9197 16970 9265 17016
rect 9311 16970 9379 17016
rect 9425 16970 9493 17016
rect 9539 16970 9607 17016
rect 9653 16970 9721 17016
rect 9767 16970 9835 17016
rect 9881 16970 9949 17016
rect 9995 16970 10063 17016
rect 10109 16970 10177 17016
rect 10223 16970 10291 17016
rect 10337 16970 10405 17016
rect 10451 16970 10519 17016
rect 10565 16970 10633 17016
rect 10679 16970 10747 17016
rect 10793 16970 10861 17016
rect 10907 16970 10975 17016
rect 11021 16970 11089 17016
rect 11135 16970 11203 17016
rect 11249 16970 11317 17016
rect 11363 16970 11431 17016
rect 11477 16970 11545 17016
rect 11591 16970 11659 17016
rect 11705 16970 11773 17016
rect 11819 16970 11927 17016
rect 11973 16970 12041 17016
rect 12087 16970 12098 17016
rect 1576 16902 12098 16970
rect 1576 16856 1587 16902
rect 1633 16856 1701 16902
rect 1747 16856 1855 16902
rect 1901 16856 1969 16902
rect 2015 16856 2083 16902
rect 2129 16856 2197 16902
rect 2243 16856 2311 16902
rect 2357 16856 2425 16902
rect 2471 16856 2539 16902
rect 2585 16856 2653 16902
rect 2699 16856 2767 16902
rect 2813 16856 2881 16902
rect 2927 16856 2995 16902
rect 3041 16856 3109 16902
rect 3155 16856 3223 16902
rect 3269 16856 3337 16902
rect 3383 16856 3451 16902
rect 3497 16856 3565 16902
rect 3611 16856 3679 16902
rect 3725 16856 3793 16902
rect 3839 16856 3907 16902
rect 3953 16856 4021 16902
rect 4067 16856 4135 16902
rect 4181 16856 4249 16902
rect 4295 16856 4363 16902
rect 4409 16856 4477 16902
rect 4523 16856 4591 16902
rect 4637 16856 4705 16902
rect 4751 16856 4819 16902
rect 4865 16856 4933 16902
rect 4979 16856 5047 16902
rect 5093 16856 5161 16902
rect 5207 16856 5275 16902
rect 5321 16856 5389 16902
rect 5435 16856 5503 16902
rect 5549 16856 5617 16902
rect 5663 16856 5731 16902
rect 5777 16856 5845 16902
rect 5891 16856 5959 16902
rect 6005 16856 6073 16902
rect 6119 16856 6187 16902
rect 6233 16856 6301 16902
rect 6347 16856 6415 16902
rect 6461 16856 6529 16902
rect 6575 16856 6643 16902
rect 6689 16856 6757 16902
rect 6803 16856 6871 16902
rect 6917 16856 6985 16902
rect 7031 16856 7099 16902
rect 7145 16856 7213 16902
rect 7259 16856 7327 16902
rect 7373 16856 7441 16902
rect 7487 16856 7555 16902
rect 7601 16856 7669 16902
rect 7715 16856 7783 16902
rect 7829 16856 7897 16902
rect 7943 16856 8011 16902
rect 8057 16856 8125 16902
rect 8171 16856 8239 16902
rect 8285 16856 8353 16902
rect 8399 16856 8467 16902
rect 8513 16856 8581 16902
rect 8627 16856 8695 16902
rect 8741 16856 8809 16902
rect 8855 16856 8923 16902
rect 8969 16856 9037 16902
rect 9083 16856 9151 16902
rect 9197 16856 9265 16902
rect 9311 16856 9379 16902
rect 9425 16856 9493 16902
rect 9539 16856 9607 16902
rect 9653 16856 9721 16902
rect 9767 16856 9835 16902
rect 9881 16856 9949 16902
rect 9995 16856 10063 16902
rect 10109 16856 10177 16902
rect 10223 16856 10291 16902
rect 10337 16856 10405 16902
rect 10451 16856 10519 16902
rect 10565 16856 10633 16902
rect 10679 16856 10747 16902
rect 10793 16856 10861 16902
rect 10907 16856 10975 16902
rect 11021 16856 11089 16902
rect 11135 16856 11203 16902
rect 11249 16856 11317 16902
rect 11363 16856 11431 16902
rect 11477 16856 11545 16902
rect 11591 16856 11659 16902
rect 11705 16856 11773 16902
rect 11819 16856 11927 16902
rect 11973 16856 12041 16902
rect 12087 16856 12098 16902
rect 1576 16844 12098 16856
rect 1576 16788 1758 16844
rect 1576 16742 1587 16788
rect 1633 16742 1701 16788
rect 1747 16742 1758 16788
rect 1576 16681 1758 16742
rect 11916 16788 12098 16844
rect 11916 16742 11927 16788
rect 11973 16742 12041 16788
rect 12087 16742 12098 16788
rect -2 16610 13 16656
rect 59 16610 74 16656
rect -2 16552 74 16610
rect 11916 16674 12098 16742
rect 11916 16628 11927 16674
rect 11973 16628 12041 16674
rect 12087 16628 12098 16674
rect -2 16506 13 16552
rect 59 16506 74 16552
rect -2 16448 74 16506
rect -2 16402 13 16448
rect 59 16402 74 16448
rect -2 16344 74 16402
rect -2 16298 13 16344
rect 59 16298 74 16344
rect -2 16240 74 16298
rect -2 16194 13 16240
rect 59 16194 74 16240
rect -2 16136 74 16194
rect -2 16090 13 16136
rect 59 16090 74 16136
rect -2 16032 74 16090
rect -2 15986 13 16032
rect 59 15986 74 16032
rect -2 15928 74 15986
rect -2 15882 13 15928
rect 59 15882 74 15928
rect -2 15824 74 15882
rect -2 15778 13 15824
rect 59 15778 74 15824
rect -2 15720 74 15778
rect -2 15674 13 15720
rect 59 15674 74 15720
rect -2 15616 74 15674
rect -2 15570 13 15616
rect 59 15570 74 15616
rect -2 15512 74 15570
rect -2 15466 13 15512
rect 59 15466 74 15512
rect -2 15408 74 15466
rect -2 15362 13 15408
rect 59 15362 74 15408
rect -2 15304 74 15362
rect -2 15258 13 15304
rect 59 15258 74 15304
rect -2 15200 74 15258
rect -2 15154 13 15200
rect 59 15154 74 15200
rect -2 15096 74 15154
rect -2 15050 13 15096
rect 59 15050 74 15096
rect -2 14992 74 15050
rect -2 14946 13 14992
rect 59 14946 74 14992
rect -2 14888 74 14946
rect -2 14842 13 14888
rect 59 14842 74 14888
rect -2 14784 74 14842
rect -2 14738 13 14784
rect 59 14738 74 14784
rect -2 14680 74 14738
rect -2 14634 13 14680
rect 59 14634 74 14680
rect -2 14576 74 14634
rect -2 14530 13 14576
rect 59 14530 74 14576
rect -2 14472 74 14530
rect -2 14426 13 14472
rect 59 14426 74 14472
rect -2 14368 74 14426
rect -2 14322 13 14368
rect 59 14322 74 14368
rect -2 14264 74 14322
rect -2 14218 13 14264
rect 59 14218 74 14264
rect -2 14160 74 14218
rect -2 14114 13 14160
rect 59 14114 74 14160
rect -2 14056 74 14114
rect -2 14010 13 14056
rect 59 14010 74 14056
rect -2 13952 74 14010
rect -2 13906 13 13952
rect 59 13906 74 13952
rect -2 13848 74 13906
rect -2 13802 13 13848
rect 59 13802 74 13848
rect -2 13744 74 13802
rect -2 13698 13 13744
rect 59 13698 74 13744
rect -2 13640 74 13698
rect -2 13594 13 13640
rect 59 13594 74 13640
rect -2 13536 74 13594
rect -2 13490 13 13536
rect 59 13490 74 13536
rect -2 13432 74 13490
rect -2 13386 13 13432
rect 59 13386 74 13432
rect -2 13328 74 13386
rect -2 13282 13 13328
rect 59 13282 74 13328
rect -2 13224 74 13282
rect -2 13178 13 13224
rect 59 13178 74 13224
rect -2 13120 74 13178
rect -2 13074 13 13120
rect 59 13074 74 13120
rect -2 13016 74 13074
rect -2 12970 13 13016
rect 59 12970 74 13016
rect -2 12912 74 12970
rect -2 12866 13 12912
rect 59 12866 74 12912
rect -2 12808 74 12866
rect -2 12762 13 12808
rect 59 12762 74 12808
rect -2 12704 74 12762
rect -2 12658 13 12704
rect 59 12658 74 12704
rect -2 12600 74 12658
rect -2 12554 13 12600
rect 59 12554 74 12600
rect -2 12496 74 12554
rect -2 12450 13 12496
rect 59 12450 74 12496
rect -2 12392 74 12450
rect -2 12346 13 12392
rect 59 12346 74 12392
rect -2 12288 74 12346
rect -2 12242 13 12288
rect 59 12242 74 12288
rect -2 12184 74 12242
rect -2 12138 13 12184
rect 59 12138 74 12184
rect -2 12080 74 12138
rect -2 12034 13 12080
rect 59 12034 74 12080
rect -2 11976 74 12034
rect -2 11930 13 11976
rect 59 11930 74 11976
rect -2 11872 74 11930
rect -2 11826 13 11872
rect 59 11826 74 11872
rect -2 11768 74 11826
rect -2 11722 13 11768
rect 59 11722 74 11768
rect -2 11664 74 11722
rect -2 11618 13 11664
rect 59 11618 74 11664
rect -2 11560 74 11618
rect -2 11514 13 11560
rect 59 11514 74 11560
rect -2 11456 74 11514
rect -2 11410 13 11456
rect 59 11410 74 11456
rect -2 11352 74 11410
rect -2 11306 13 11352
rect 59 11306 74 11352
rect -2 11248 74 11306
rect -2 11202 13 11248
rect 59 11202 74 11248
rect -2 11144 74 11202
rect -2 11098 13 11144
rect 59 11098 74 11144
rect -2 11040 74 11098
rect -2 10994 13 11040
rect 59 10994 74 11040
rect -2 10936 74 10994
rect -2 10890 13 10936
rect 59 10890 74 10936
rect -2 10832 74 10890
rect -2 10786 13 10832
rect 59 10786 74 10832
rect -2 10728 74 10786
rect -2 10682 13 10728
rect 59 10682 74 10728
rect -2 10624 74 10682
rect -2 10578 13 10624
rect 59 10578 74 10624
rect -2 10520 74 10578
rect -2 10474 13 10520
rect 59 10474 74 10520
rect -2 10416 74 10474
rect -2 10370 13 10416
rect 59 10370 74 10416
rect -2 10312 74 10370
rect -2 10266 13 10312
rect 59 10266 74 10312
rect -2 10208 74 10266
rect -2 10162 13 10208
rect 59 10162 74 10208
rect -2 10104 74 10162
rect -2 10058 13 10104
rect 59 10058 74 10104
rect -2 10000 74 10058
rect -2 9954 13 10000
rect 59 9954 74 10000
rect -2 9896 74 9954
rect -2 9850 13 9896
rect 59 9850 74 9896
rect -2 9792 74 9850
rect -2 9746 13 9792
rect 59 9746 74 9792
rect -2 9688 74 9746
rect -2 9642 13 9688
rect 59 9642 74 9688
rect -2 9584 74 9642
rect -2 9538 13 9584
rect 59 9538 74 9584
rect -2 9480 74 9538
rect -2 9434 13 9480
rect 59 9434 74 9480
rect -2 9376 74 9434
rect -2 9330 13 9376
rect 59 9330 74 9376
rect -2 9272 74 9330
rect -2 9226 13 9272
rect 59 9226 74 9272
rect -2 9168 74 9226
rect -2 9122 13 9168
rect 59 9122 74 9168
rect -2 9064 74 9122
rect -2 9018 13 9064
rect 59 9018 74 9064
rect -2 8960 74 9018
rect -2 8914 13 8960
rect 59 8914 74 8960
rect -2 8856 74 8914
rect -2 8810 13 8856
rect 59 8810 74 8856
rect -2 8752 74 8810
rect -2 8706 13 8752
rect 59 8706 74 8752
rect -2 8648 74 8706
rect -2 8602 13 8648
rect 59 8602 74 8648
rect -2 8544 74 8602
rect -2 8498 13 8544
rect 59 8498 74 8544
rect -2 8440 74 8498
rect -2 8394 13 8440
rect 59 8394 74 8440
rect -2 8336 74 8394
rect -2 8290 13 8336
rect 59 8290 74 8336
rect -2 8232 74 8290
rect -2 8186 13 8232
rect 59 8186 74 8232
rect -2 8128 74 8186
rect -2 8082 13 8128
rect 59 8082 74 8128
rect -2 8024 74 8082
rect -2 7978 13 8024
rect 59 7978 74 8024
rect -2 7920 74 7978
rect -2 7874 13 7920
rect 59 7874 74 7920
rect -2 7816 74 7874
rect -2 7770 13 7816
rect 59 7770 74 7816
rect -2 7712 74 7770
rect -2 7666 13 7712
rect 59 7666 74 7712
rect -2 7608 74 7666
rect -2 7562 13 7608
rect 59 7562 74 7608
rect -2 7504 74 7562
rect -2 7458 13 7504
rect 59 7458 74 7504
rect -2 7400 74 7458
rect -2 7354 13 7400
rect 59 7354 74 7400
rect -2 7296 74 7354
rect -2 7250 13 7296
rect 59 7250 74 7296
rect -2 7192 74 7250
rect -2 7146 13 7192
rect 59 7146 74 7192
rect -2 7088 74 7146
rect -2 7042 13 7088
rect 59 7042 74 7088
rect -2 6984 74 7042
rect -2 6938 13 6984
rect 59 6938 74 6984
rect -2 6880 74 6938
rect -2 6834 13 6880
rect 59 6834 74 6880
rect -2 6776 74 6834
rect -2 6730 13 6776
rect 59 6730 74 6776
rect -2 6672 74 6730
rect -2 6626 13 6672
rect 59 6626 74 6672
rect -2 6568 74 6626
rect -2 6522 13 6568
rect 59 6522 74 6568
rect -2 6464 74 6522
rect -2 6418 13 6464
rect 59 6418 74 6464
rect -2 6360 74 6418
rect -2 6314 13 6360
rect 59 6314 74 6360
rect -2 6256 74 6314
rect -2 6210 13 6256
rect 59 6210 74 6256
rect -2 6152 74 6210
rect -2 6106 13 6152
rect 59 6106 74 6152
rect -2 6048 74 6106
rect -2 6002 13 6048
rect 59 6002 74 6048
rect -2 5944 74 6002
rect -2 5898 13 5944
rect 59 5898 74 5944
rect -2 5840 74 5898
rect -2 5794 13 5840
rect 59 5794 74 5840
rect -2 5736 74 5794
rect -2 5690 13 5736
rect 59 5690 74 5736
rect -2 5632 74 5690
rect -2 5586 13 5632
rect 59 5586 74 5632
rect -2 5528 74 5586
rect -2 5482 13 5528
rect 59 5482 74 5528
rect -2 5424 74 5482
rect -2 5378 13 5424
rect 59 5378 74 5424
rect -2 5320 74 5378
rect -2 5274 13 5320
rect 59 5274 74 5320
rect -2 5216 74 5274
rect -2 5170 13 5216
rect 59 5170 74 5216
rect -2 5112 74 5170
rect -2 5066 13 5112
rect 59 5066 74 5112
rect -2 5008 74 5066
rect -2 4962 13 5008
rect 59 4962 74 5008
rect -2 4904 74 4962
rect -2 4858 13 4904
rect 59 4858 74 4904
rect -2 4800 74 4858
rect -2 4754 13 4800
rect 59 4754 74 4800
rect -2 4696 74 4754
rect -2 4650 13 4696
rect 59 4650 74 4696
rect -2 4592 74 4650
rect -2 4546 13 4592
rect 59 4546 74 4592
rect -2 4455 74 4546
rect 355 16441 11446 16573
rect 355 16430 4138 16441
rect 355 16411 2233 16430
rect 355 5279 423 16411
rect 2222 16384 2233 16411
rect 4127 16384 4138 16430
rect 2222 16373 4138 16384
rect 4658 16430 6574 16441
rect 4658 16384 4669 16430
rect 6563 16384 6574 16430
rect 4658 16373 6574 16384
rect 7094 16430 9010 16441
rect 7094 16384 7105 16430
rect 8999 16384 9010 16430
rect 7094 16373 9010 16384
rect 9530 16430 11446 16441
rect 9530 16384 9541 16430
rect 11435 16384 11446 16430
rect 9530 16373 11446 16384
rect 11916 16560 12098 16628
rect 11916 16514 11927 16560
rect 11973 16514 12041 16560
rect 12087 16514 12098 16560
rect 11916 16446 12098 16514
rect 11916 16400 11927 16446
rect 11973 16400 12041 16446
rect 12087 16400 12098 16446
rect 1576 16314 2162 16351
rect 1576 16218 2105 16314
rect 1576 16172 1587 16218
rect 1633 16172 1701 16218
rect 1747 16172 2105 16218
rect 1576 16104 2105 16172
rect 1576 16058 1587 16104
rect 1633 16058 1701 16104
rect 1747 16058 2105 16104
rect 1576 15990 2105 16058
rect 1576 15944 1587 15990
rect 1633 15944 1701 15990
rect 1747 15944 2105 15990
rect 1576 15876 2105 15944
rect 1576 15830 1587 15876
rect 1633 15830 1701 15876
rect 1747 15830 2105 15876
rect 1576 15762 2105 15830
rect 1576 15716 1587 15762
rect 1633 15716 1701 15762
rect 1747 15716 2105 15762
rect 1576 15648 2105 15716
rect 1576 15602 1587 15648
rect 1633 15602 1701 15648
rect 1747 15602 2105 15648
rect 1576 15534 2105 15602
rect 1576 15488 1587 15534
rect 1633 15488 1701 15534
rect 1747 15488 2105 15534
rect 1576 15420 2105 15488
rect 1576 15374 1587 15420
rect 1633 15374 1701 15420
rect 1747 15374 2105 15420
rect 1576 15306 2105 15374
rect 1576 15260 1587 15306
rect 1633 15260 1701 15306
rect 1747 15260 2105 15306
rect 1576 15192 2105 15260
rect 1576 15146 1587 15192
rect 1633 15146 1701 15192
rect 1747 15146 2105 15192
rect 1576 15078 2105 15146
rect 1576 15032 1587 15078
rect 1633 15032 1701 15078
rect 1747 15032 2105 15078
rect 1576 14964 2105 15032
rect 1576 14918 1587 14964
rect 1633 14918 1701 14964
rect 1747 14918 2105 14964
rect 1576 14850 2105 14918
rect 1576 14804 1587 14850
rect 1633 14804 1701 14850
rect 1747 14804 2105 14850
rect 1576 14736 2105 14804
rect 1576 14690 1587 14736
rect 1633 14690 1701 14736
rect 1747 14690 2105 14736
rect 1576 14622 2105 14690
rect 1576 14576 1587 14622
rect 1633 14576 1701 14622
rect 1747 14576 2105 14622
rect 1576 14508 2105 14576
rect 1576 14462 1587 14508
rect 1633 14462 1701 14508
rect 1747 14462 2105 14508
rect 1576 14394 2105 14462
rect 1576 14348 1587 14394
rect 1633 14348 1701 14394
rect 1747 14348 2105 14394
rect 1576 14280 2105 14348
rect 1576 14234 1587 14280
rect 1633 14234 1701 14280
rect 1747 14234 2105 14280
rect 1576 14166 2105 14234
rect 1576 14120 1587 14166
rect 1633 14120 1701 14166
rect 1747 14120 2105 14166
rect 1576 14052 2105 14120
rect 1576 14006 1587 14052
rect 1633 14006 1701 14052
rect 1747 14006 2105 14052
rect 1576 13938 2105 14006
rect 1576 13892 1587 13938
rect 1633 13892 1701 13938
rect 1747 13892 2105 13938
rect 1576 13824 2105 13892
rect 1576 13778 1587 13824
rect 1633 13778 1701 13824
rect 1747 13778 2105 13824
rect 1576 13710 2105 13778
rect 1576 13664 1587 13710
rect 1633 13664 1701 13710
rect 1747 13664 2105 13710
rect 1576 13596 2105 13664
rect 1576 13550 1587 13596
rect 1633 13550 1701 13596
rect 1747 13550 2105 13596
rect 1576 13482 2105 13550
rect 1576 13436 1587 13482
rect 1633 13436 1701 13482
rect 1747 13436 2105 13482
rect 1576 13368 2105 13436
rect 1576 13322 1587 13368
rect 1633 13322 1701 13368
rect 1747 13322 2105 13368
rect 1576 13254 2105 13322
rect 1576 13208 1587 13254
rect 1633 13208 1701 13254
rect 1747 13208 2105 13254
rect 1576 13140 2105 13208
rect 1576 13094 1587 13140
rect 1633 13094 1701 13140
rect 1747 13094 2105 13140
rect 1576 13026 2105 13094
rect 1576 12980 1587 13026
rect 1633 12980 1701 13026
rect 1747 12980 2105 13026
rect 1576 12912 2105 12980
rect 1576 12866 1587 12912
rect 1633 12866 1701 12912
rect 1747 12866 2105 12912
rect 1576 12798 2105 12866
rect 1576 12752 1587 12798
rect 1633 12752 1701 12798
rect 1747 12752 2105 12798
rect 1576 12684 2105 12752
rect 1576 12638 1587 12684
rect 1633 12638 1701 12684
rect 1747 12638 2105 12684
rect 1576 12570 2105 12638
rect 1576 12524 1587 12570
rect 1633 12524 1701 12570
rect 1747 12524 2105 12570
rect 1576 12456 2105 12524
rect 1576 12410 1587 12456
rect 1633 12410 1701 12456
rect 1747 12410 2105 12456
rect 1576 12342 2105 12410
rect 1576 12296 1587 12342
rect 1633 12296 1701 12342
rect 1747 12296 2105 12342
rect 1576 12228 2105 12296
rect 1576 12182 1587 12228
rect 1633 12182 1701 12228
rect 1747 12182 2105 12228
rect 1576 12114 2105 12182
rect 1576 12068 1587 12114
rect 1633 12068 1701 12114
rect 1747 12068 2105 12114
rect 1576 12000 2105 12068
rect 1576 11954 1587 12000
rect 1633 11954 1701 12000
rect 1747 11954 2105 12000
rect 1576 11886 2105 11954
rect 1576 11840 1587 11886
rect 1633 11840 1701 11886
rect 1747 11840 2105 11886
rect 1576 11772 2105 11840
rect 1576 11726 1587 11772
rect 1633 11726 1701 11772
rect 1747 11726 2105 11772
rect 1576 11658 2105 11726
rect 1576 11612 1587 11658
rect 1633 11612 1701 11658
rect 1747 11612 2105 11658
rect 1576 11544 2105 11612
rect 1576 11498 1587 11544
rect 1633 11498 1701 11544
rect 1747 11498 2105 11544
rect 1576 11430 2105 11498
rect 1576 11384 1587 11430
rect 1633 11384 1701 11430
rect 1747 11388 2105 11430
rect 2151 11388 2162 16314
rect 1747 11384 2162 11388
rect 1576 11316 2162 11384
rect 2680 11329 3680 16373
rect 4198 16314 4598 16351
rect 4198 11388 4209 16314
rect 4255 11388 4541 16314
rect 4587 11388 4598 16314
rect 1576 11270 1587 11316
rect 1633 11270 1701 11316
rect 1747 11270 2162 11316
rect 1576 11202 2162 11270
rect 2222 11318 4138 11329
rect 2222 11272 2233 11318
rect 4127 11272 4138 11318
rect 2222 11261 4138 11272
rect 1576 11156 1587 11202
rect 1633 11156 1701 11202
rect 1747 11201 2162 11202
rect 4198 11201 4598 11388
rect 5116 11329 6116 16373
rect 6634 16314 7034 16351
rect 6634 11388 6645 16314
rect 6691 11388 6977 16314
rect 7023 11388 7034 16314
rect 4658 11318 6574 11329
rect 4658 11272 4669 11318
rect 6563 11272 6574 11318
rect 4658 11261 6574 11272
rect 6634 11201 7034 11388
rect 7552 11329 8552 16373
rect 9070 16314 9470 16351
rect 9070 11388 9081 16314
rect 9127 11388 9413 16314
rect 9459 11388 9470 16314
rect 7094 11318 9010 11329
rect 7094 11272 7105 11318
rect 8999 11272 9010 11318
rect 7094 11261 9010 11272
rect 9070 11201 9470 11388
rect 9988 11329 10988 16373
rect 11916 16351 12098 16400
rect 11506 16332 12098 16351
rect 11506 16314 11927 16332
rect 11506 11388 11517 16314
rect 11563 16286 11927 16314
rect 11973 16286 12041 16332
rect 12087 16286 12098 16332
rect 11563 16218 12098 16286
rect 11563 16172 11927 16218
rect 11973 16172 12041 16218
rect 12087 16172 12098 16218
rect 11563 16104 12098 16172
rect 11563 16058 11927 16104
rect 11973 16058 12041 16104
rect 12087 16058 12098 16104
rect 11563 15990 12098 16058
rect 11563 15944 11927 15990
rect 11973 15944 12041 15990
rect 12087 15944 12098 15990
rect 11563 15876 12098 15944
rect 11563 15830 11927 15876
rect 11973 15830 12041 15876
rect 12087 15830 12098 15876
rect 11563 15762 12098 15830
rect 11563 15716 11927 15762
rect 11973 15716 12041 15762
rect 12087 15716 12098 15762
rect 11563 15648 12098 15716
rect 11563 15602 11927 15648
rect 11973 15602 12041 15648
rect 12087 15602 12098 15648
rect 11563 15534 12098 15602
rect 11563 15488 11927 15534
rect 11973 15488 12041 15534
rect 12087 15488 12098 15534
rect 11563 15420 12098 15488
rect 11563 15374 11927 15420
rect 11973 15374 12041 15420
rect 12087 15374 12098 15420
rect 11563 15306 12098 15374
rect 11563 15260 11927 15306
rect 11973 15260 12041 15306
rect 12087 15260 12098 15306
rect 11563 15192 12098 15260
rect 11563 15146 11927 15192
rect 11973 15146 12041 15192
rect 12087 15146 12098 15192
rect 11563 15078 12098 15146
rect 11563 15032 11927 15078
rect 11973 15032 12041 15078
rect 12087 15032 12098 15078
rect 11563 14964 12098 15032
rect 11563 14918 11927 14964
rect 11973 14918 12041 14964
rect 12087 14918 12098 14964
rect 11563 14850 12098 14918
rect 11563 14804 11927 14850
rect 11973 14804 12041 14850
rect 12087 14804 12098 14850
rect 11563 14736 12098 14804
rect 11563 14690 11927 14736
rect 11973 14690 12041 14736
rect 12087 14690 12098 14736
rect 11563 14622 12098 14690
rect 11563 14576 11927 14622
rect 11973 14576 12041 14622
rect 12087 14576 12098 14622
rect 11563 14508 12098 14576
rect 11563 14462 11927 14508
rect 11973 14462 12041 14508
rect 12087 14462 12098 14508
rect 11563 14394 12098 14462
rect 11563 14348 11927 14394
rect 11973 14348 12041 14394
rect 12087 14348 12098 14394
rect 11563 14280 12098 14348
rect 11563 14234 11927 14280
rect 11973 14234 12041 14280
rect 12087 14234 12098 14280
rect 11563 14166 12098 14234
rect 11563 14120 11927 14166
rect 11973 14120 12041 14166
rect 12087 14120 12098 14166
rect 11563 14052 12098 14120
rect 11563 14006 11927 14052
rect 11973 14006 12041 14052
rect 12087 14006 12098 14052
rect 11563 13938 12098 14006
rect 11563 13892 11927 13938
rect 11973 13892 12041 13938
rect 12087 13892 12098 13938
rect 11563 13824 12098 13892
rect 11563 13778 11927 13824
rect 11973 13778 12041 13824
rect 12087 13778 12098 13824
rect 11563 13710 12098 13778
rect 11563 13664 11927 13710
rect 11973 13664 12041 13710
rect 12087 13664 12098 13710
rect 11563 13596 12098 13664
rect 11563 13550 11927 13596
rect 11973 13550 12041 13596
rect 12087 13550 12098 13596
rect 11563 13482 12098 13550
rect 11563 13436 11927 13482
rect 11973 13436 12041 13482
rect 12087 13436 12098 13482
rect 11563 13368 12098 13436
rect 11563 13322 11927 13368
rect 11973 13322 12041 13368
rect 12087 13322 12098 13368
rect 11563 13254 12098 13322
rect 11563 13208 11927 13254
rect 11973 13208 12041 13254
rect 12087 13208 12098 13254
rect 11563 13140 12098 13208
rect 11563 13094 11927 13140
rect 11973 13094 12041 13140
rect 12087 13094 12098 13140
rect 11563 13026 12098 13094
rect 11563 12980 11927 13026
rect 11973 12980 12041 13026
rect 12087 12980 12098 13026
rect 11563 12912 12098 12980
rect 11563 12866 11927 12912
rect 11973 12866 12041 12912
rect 12087 12866 12098 12912
rect 11563 12798 12098 12866
rect 11563 12752 11927 12798
rect 11973 12752 12041 12798
rect 12087 12752 12098 12798
rect 11563 12684 12098 12752
rect 11563 12638 11927 12684
rect 11973 12638 12041 12684
rect 12087 12638 12098 12684
rect 11563 12570 12098 12638
rect 11563 12524 11927 12570
rect 11973 12524 12041 12570
rect 12087 12524 12098 12570
rect 11563 12456 12098 12524
rect 11563 12410 11927 12456
rect 11973 12410 12041 12456
rect 12087 12410 12098 12456
rect 11563 12342 12098 12410
rect 11563 12296 11927 12342
rect 11973 12296 12041 12342
rect 12087 12296 12098 12342
rect 11563 12228 12098 12296
rect 11563 12182 11927 12228
rect 11973 12182 12041 12228
rect 12087 12182 12098 12228
rect 11563 12114 12098 12182
rect 11563 12068 11927 12114
rect 11973 12068 12041 12114
rect 12087 12068 12098 12114
rect 11563 12000 12098 12068
rect 11563 11954 11927 12000
rect 11973 11954 12041 12000
rect 12087 11954 12098 12000
rect 11563 11886 12098 11954
rect 11563 11840 11927 11886
rect 11973 11840 12041 11886
rect 12087 11840 12098 11886
rect 11563 11772 12098 11840
rect 11563 11726 11927 11772
rect 11973 11726 12041 11772
rect 12087 11726 12098 11772
rect 11563 11658 12098 11726
rect 11563 11612 11927 11658
rect 11973 11612 12041 11658
rect 12087 11612 12098 11658
rect 11563 11544 12098 11612
rect 11563 11498 11927 11544
rect 11973 11498 12041 11544
rect 12087 11498 12098 11544
rect 11563 11430 12098 11498
rect 11563 11388 11927 11430
rect 11506 11384 11927 11388
rect 11973 11384 12041 11430
rect 12087 11384 12098 11430
rect 9530 11318 11446 11329
rect 9530 11272 9541 11318
rect 11435 11272 11446 11318
rect 9530 11261 11446 11272
rect 11506 11316 12098 11384
rect 11506 11270 11927 11316
rect 11973 11270 12041 11316
rect 12087 11270 12098 11316
rect 11506 11202 12098 11270
rect 11506 11201 11927 11202
rect 1747 11156 11927 11201
rect 11973 11156 12041 11202
rect 12087 11156 12098 11202
rect 1576 11088 12098 11156
rect 1576 11042 1587 11088
rect 1633 11042 1701 11088
rect 1747 11042 11927 11088
rect 11973 11042 12041 11088
rect 12087 11042 12098 11088
rect 1576 10974 12098 11042
rect 1576 10928 1587 10974
rect 1633 10928 1701 10974
rect 1747 10928 11927 10974
rect 11973 10928 12041 10974
rect 12087 10928 12098 10974
rect 1576 10925 12098 10928
rect 1576 10879 1855 10925
rect 1901 10879 1969 10925
rect 2015 10879 2083 10925
rect 2129 10879 2197 10925
rect 2243 10879 2311 10925
rect 2357 10879 2425 10925
rect 2471 10879 2539 10925
rect 2585 10879 2653 10925
rect 2699 10879 2767 10925
rect 2813 10879 2881 10925
rect 2927 10879 2995 10925
rect 3041 10879 3109 10925
rect 3155 10879 3223 10925
rect 3269 10879 3337 10925
rect 3383 10879 3451 10925
rect 3497 10879 3565 10925
rect 3611 10879 3679 10925
rect 3725 10879 3793 10925
rect 3839 10879 3907 10925
rect 3953 10879 4021 10925
rect 4067 10879 4135 10925
rect 4181 10879 4249 10925
rect 4295 10879 4363 10925
rect 4409 10879 4477 10925
rect 4523 10879 4591 10925
rect 4637 10879 4705 10925
rect 4751 10879 4819 10925
rect 4865 10879 4933 10925
rect 4979 10879 5047 10925
rect 5093 10879 5161 10925
rect 5207 10879 5275 10925
rect 5321 10879 5389 10925
rect 5435 10879 5503 10925
rect 5549 10879 5617 10925
rect 5663 10879 5731 10925
rect 5777 10879 5845 10925
rect 5891 10879 5959 10925
rect 6005 10879 6073 10925
rect 6119 10879 6187 10925
rect 6233 10879 6301 10925
rect 6347 10879 6415 10925
rect 6461 10879 6529 10925
rect 6575 10879 6643 10925
rect 6689 10879 6757 10925
rect 6803 10879 6871 10925
rect 6917 10879 6985 10925
rect 7031 10879 7099 10925
rect 7145 10879 7213 10925
rect 7259 10879 7327 10925
rect 7373 10879 7441 10925
rect 7487 10879 7555 10925
rect 7601 10879 7669 10925
rect 7715 10879 7783 10925
rect 7829 10879 7897 10925
rect 7943 10879 8011 10925
rect 8057 10879 8125 10925
rect 8171 10879 8239 10925
rect 8285 10879 8353 10925
rect 8399 10879 8467 10925
rect 8513 10879 8581 10925
rect 8627 10879 8695 10925
rect 8741 10879 8809 10925
rect 8855 10879 8923 10925
rect 8969 10879 9037 10925
rect 9083 10879 9151 10925
rect 9197 10879 9265 10925
rect 9311 10879 9379 10925
rect 9425 10879 9493 10925
rect 9539 10879 9607 10925
rect 9653 10879 9721 10925
rect 9767 10879 9835 10925
rect 9881 10879 9949 10925
rect 9995 10879 10063 10925
rect 10109 10879 10177 10925
rect 10223 10879 10291 10925
rect 10337 10879 10405 10925
rect 10451 10879 10519 10925
rect 10565 10879 10633 10925
rect 10679 10879 10747 10925
rect 10793 10879 10861 10925
rect 10907 10879 10975 10925
rect 11021 10879 11089 10925
rect 11135 10879 11203 10925
rect 11249 10879 11317 10925
rect 11363 10879 11431 10925
rect 11477 10879 11545 10925
rect 11591 10879 11659 10925
rect 11705 10879 11773 10925
rect 11819 10879 12098 10925
rect 1576 10860 12098 10879
rect 1576 10814 1587 10860
rect 1633 10814 1701 10860
rect 1747 10814 11927 10860
rect 11973 10814 12041 10860
rect 12087 10814 12098 10860
rect 1576 10811 12098 10814
rect 1576 10765 1855 10811
rect 1901 10765 1969 10811
rect 2015 10765 2083 10811
rect 2129 10765 2197 10811
rect 2243 10765 2311 10811
rect 2357 10765 2425 10811
rect 2471 10765 2539 10811
rect 2585 10765 2653 10811
rect 2699 10765 2767 10811
rect 2813 10765 2881 10811
rect 2927 10765 2995 10811
rect 3041 10765 3109 10811
rect 3155 10765 3223 10811
rect 3269 10765 3337 10811
rect 3383 10765 3451 10811
rect 3497 10765 3565 10811
rect 3611 10765 3679 10811
rect 3725 10765 3793 10811
rect 3839 10765 3907 10811
rect 3953 10765 4021 10811
rect 4067 10765 4135 10811
rect 4181 10765 4249 10811
rect 4295 10765 4363 10811
rect 4409 10765 4477 10811
rect 4523 10765 4591 10811
rect 4637 10765 4705 10811
rect 4751 10765 4819 10811
rect 4865 10765 4933 10811
rect 4979 10765 5047 10811
rect 5093 10765 5161 10811
rect 5207 10765 5275 10811
rect 5321 10765 5389 10811
rect 5435 10765 5503 10811
rect 5549 10765 5617 10811
rect 5663 10765 5731 10811
rect 5777 10765 5845 10811
rect 5891 10765 5959 10811
rect 6005 10765 6073 10811
rect 6119 10765 6187 10811
rect 6233 10765 6301 10811
rect 6347 10765 6415 10811
rect 6461 10765 6529 10811
rect 6575 10765 6643 10811
rect 6689 10765 6757 10811
rect 6803 10765 6871 10811
rect 6917 10765 6985 10811
rect 7031 10765 7099 10811
rect 7145 10765 7213 10811
rect 7259 10765 7327 10811
rect 7373 10765 7441 10811
rect 7487 10765 7555 10811
rect 7601 10765 7669 10811
rect 7715 10765 7783 10811
rect 7829 10765 7897 10811
rect 7943 10765 8011 10811
rect 8057 10765 8125 10811
rect 8171 10765 8239 10811
rect 8285 10765 8353 10811
rect 8399 10765 8467 10811
rect 8513 10765 8581 10811
rect 8627 10765 8695 10811
rect 8741 10765 8809 10811
rect 8855 10765 8923 10811
rect 8969 10765 9037 10811
rect 9083 10765 9151 10811
rect 9197 10765 9265 10811
rect 9311 10765 9379 10811
rect 9425 10765 9493 10811
rect 9539 10765 9607 10811
rect 9653 10765 9721 10811
rect 9767 10765 9835 10811
rect 9881 10765 9949 10811
rect 9995 10765 10063 10811
rect 10109 10765 10177 10811
rect 10223 10765 10291 10811
rect 10337 10765 10405 10811
rect 10451 10765 10519 10811
rect 10565 10765 10633 10811
rect 10679 10765 10747 10811
rect 10793 10765 10861 10811
rect 10907 10765 10975 10811
rect 11021 10765 11089 10811
rect 11135 10765 11203 10811
rect 11249 10765 11317 10811
rect 11363 10765 11431 10811
rect 11477 10765 11545 10811
rect 11591 10765 11659 10811
rect 11705 10765 11773 10811
rect 11819 10765 12098 10811
rect 1576 10746 12098 10765
rect 1576 10700 1587 10746
rect 1633 10700 1701 10746
rect 1747 10700 11927 10746
rect 11973 10700 12041 10746
rect 12087 10700 12098 10746
rect 1576 10632 12098 10700
rect 1576 10586 1587 10632
rect 1633 10586 1701 10632
rect 1747 10586 11927 10632
rect 11973 10586 12041 10632
rect 12087 10586 12098 10632
rect 1576 10518 12098 10586
rect 1576 10472 1587 10518
rect 1633 10472 1701 10518
rect 1747 10489 11927 10518
rect 1747 10472 2162 10489
rect 1576 10404 2162 10472
rect 1576 10358 1587 10404
rect 1633 10358 1701 10404
rect 1747 10358 2162 10404
rect 2222 10418 4138 10429
rect 2222 10372 2233 10418
rect 4127 10372 4138 10418
rect 2222 10361 4138 10372
rect 1576 10302 2162 10358
rect 1576 10290 2105 10302
rect 1576 10244 1587 10290
rect 1633 10244 1701 10290
rect 1747 10244 2105 10290
rect 1576 10176 2105 10244
rect 1576 10130 1587 10176
rect 1633 10130 1701 10176
rect 1747 10130 2105 10176
rect 1576 10062 2105 10130
rect 1576 10016 1587 10062
rect 1633 10016 1701 10062
rect 1747 10016 2105 10062
rect 1576 9948 2105 10016
rect 1576 9902 1587 9948
rect 1633 9902 1701 9948
rect 1747 9902 2105 9948
rect 1576 9834 2105 9902
rect 1576 9788 1587 9834
rect 1633 9788 1701 9834
rect 1747 9788 2105 9834
rect 1576 9720 2105 9788
rect 1576 9674 1587 9720
rect 1633 9674 1701 9720
rect 1747 9674 2105 9720
rect 1576 9606 2105 9674
rect 1576 9560 1587 9606
rect 1633 9560 1701 9606
rect 1747 9560 2105 9606
rect 1576 9492 2105 9560
rect 1576 9446 1587 9492
rect 1633 9446 1701 9492
rect 1747 9446 2105 9492
rect 1576 9378 2105 9446
rect 1576 9332 1587 9378
rect 1633 9332 1701 9378
rect 1747 9332 2105 9378
rect 1576 9264 2105 9332
rect 1576 9218 1587 9264
rect 1633 9218 1701 9264
rect 1747 9218 2105 9264
rect 1576 9150 2105 9218
rect 1576 9104 1587 9150
rect 1633 9104 1701 9150
rect 1747 9104 2105 9150
rect 1576 9036 2105 9104
rect 1576 8990 1587 9036
rect 1633 8990 1701 9036
rect 1747 8990 2105 9036
rect 1576 8922 2105 8990
rect 1576 8876 1587 8922
rect 1633 8876 1701 8922
rect 1747 8876 2105 8922
rect 1576 8808 2105 8876
rect 1576 8762 1587 8808
rect 1633 8762 1701 8808
rect 1747 8762 2105 8808
rect 1576 8694 2105 8762
rect 1576 8648 1587 8694
rect 1633 8648 1701 8694
rect 1747 8648 2105 8694
rect 1576 8580 2105 8648
rect 1576 8534 1587 8580
rect 1633 8534 1701 8580
rect 1747 8534 2105 8580
rect 1576 8466 2105 8534
rect 1576 8420 1587 8466
rect 1633 8420 1701 8466
rect 1747 8420 2105 8466
rect 1576 8352 2105 8420
rect 1576 8306 1587 8352
rect 1633 8306 1701 8352
rect 1747 8306 2105 8352
rect 1576 8238 2105 8306
rect 1576 8192 1587 8238
rect 1633 8192 1701 8238
rect 1747 8192 2105 8238
rect 1576 8124 2105 8192
rect 1576 8078 1587 8124
rect 1633 8078 1701 8124
rect 1747 8078 2105 8124
rect 1576 8010 2105 8078
rect 1576 7964 1587 8010
rect 1633 7964 1701 8010
rect 1747 7964 2105 8010
rect 1576 7896 2105 7964
rect 1576 7850 1587 7896
rect 1633 7850 1701 7896
rect 1747 7850 2105 7896
rect 1576 7782 2105 7850
rect 1576 7736 1587 7782
rect 1633 7736 1701 7782
rect 1747 7736 2105 7782
rect 1576 7668 2105 7736
rect 1576 7622 1587 7668
rect 1633 7622 1701 7668
rect 1747 7622 2105 7668
rect 1576 7554 2105 7622
rect 1576 7508 1587 7554
rect 1633 7508 1701 7554
rect 1747 7508 2105 7554
rect 1576 7440 2105 7508
rect 1576 7394 1587 7440
rect 1633 7394 1701 7440
rect 1747 7394 2105 7440
rect 1576 7326 2105 7394
rect 1576 7280 1587 7326
rect 1633 7280 1701 7326
rect 1747 7280 2105 7326
rect 1576 7212 2105 7280
rect 1576 7166 1587 7212
rect 1633 7166 1701 7212
rect 1747 7166 2105 7212
rect 1576 7098 2105 7166
rect 1576 7052 1587 7098
rect 1633 7052 1701 7098
rect 1747 7052 2105 7098
rect 1576 6984 2105 7052
rect 1576 6938 1587 6984
rect 1633 6938 1701 6984
rect 1747 6938 2105 6984
rect 1576 6870 2105 6938
rect 1576 6824 1587 6870
rect 1633 6824 1701 6870
rect 1747 6824 2105 6870
rect 1576 6756 2105 6824
rect 1576 6710 1587 6756
rect 1633 6710 1701 6756
rect 1747 6710 2105 6756
rect 1576 6642 2105 6710
rect 1576 6596 1587 6642
rect 1633 6596 1701 6642
rect 1747 6596 2105 6642
rect 1576 6528 2105 6596
rect 1576 6482 1587 6528
rect 1633 6482 1701 6528
rect 1747 6482 2105 6528
rect 1576 6414 2105 6482
rect 1576 6368 1587 6414
rect 1633 6368 1701 6414
rect 1747 6368 2105 6414
rect 1576 6300 2105 6368
rect 1576 6254 1587 6300
rect 1633 6254 1701 6300
rect 1747 6254 2105 6300
rect 1576 6186 2105 6254
rect 1576 6140 1587 6186
rect 1633 6140 1701 6186
rect 1747 6140 2105 6186
rect 1576 6072 2105 6140
rect 1576 6026 1587 6072
rect 1633 6026 1701 6072
rect 1747 6026 2105 6072
rect 1576 5958 2105 6026
rect 1576 5912 1587 5958
rect 1633 5912 1701 5958
rect 1747 5912 2105 5958
rect 1576 5844 2105 5912
rect 1576 5798 1587 5844
rect 1633 5798 1701 5844
rect 1747 5798 2105 5844
rect 1576 5730 2105 5798
rect 1576 5684 1587 5730
rect 1633 5684 1701 5730
rect 1747 5684 2105 5730
rect 1576 5616 2105 5684
rect 1576 5570 1587 5616
rect 1633 5570 1701 5616
rect 1747 5570 2105 5616
rect 1576 5502 2105 5570
rect 1576 5456 1587 5502
rect 1633 5456 1701 5502
rect 1747 5456 2105 5502
rect 1576 5376 2105 5456
rect 2151 5376 2162 10302
rect 1576 5339 2162 5376
rect 2680 5317 3680 10361
rect 4198 10302 4598 10489
rect 4658 10418 6574 10429
rect 4658 10372 4669 10418
rect 6563 10372 6574 10418
rect 4658 10361 6574 10372
rect 4198 5376 4209 10302
rect 4255 5376 4541 10302
rect 4587 5376 4598 10302
rect 4198 5339 4598 5376
rect 5116 5317 6116 10361
rect 6634 10302 7034 10489
rect 7094 10418 9010 10429
rect 7094 10372 7105 10418
rect 8999 10372 9010 10418
rect 7094 10361 9010 10372
rect 6634 5376 6645 10302
rect 6691 5376 6977 10302
rect 7023 5376 7034 10302
rect 6634 5339 7034 5376
rect 7552 5317 8552 10361
rect 9070 10302 9470 10489
rect 11506 10472 11927 10489
rect 11973 10472 12041 10518
rect 12087 10472 12098 10518
rect 9530 10418 11446 10429
rect 9530 10372 9541 10418
rect 11435 10372 11446 10418
rect 9530 10361 11446 10372
rect 11506 10404 12098 10472
rect 9070 5376 9081 10302
rect 9127 5376 9413 10302
rect 9459 5376 9470 10302
rect 9070 5339 9470 5376
rect 9988 5317 10988 10361
rect 11506 10358 11927 10404
rect 11973 10358 12041 10404
rect 12087 10358 12098 10404
rect 11506 10302 12098 10358
rect 11506 5376 11517 10302
rect 11563 10290 12098 10302
rect 11563 10244 11927 10290
rect 11973 10244 12041 10290
rect 12087 10244 12098 10290
rect 11563 10176 12098 10244
rect 11563 10130 11927 10176
rect 11973 10130 12041 10176
rect 12087 10130 12098 10176
rect 11563 10062 12098 10130
rect 11563 10016 11927 10062
rect 11973 10016 12041 10062
rect 12087 10016 12098 10062
rect 11563 9948 12098 10016
rect 11563 9902 11927 9948
rect 11973 9902 12041 9948
rect 12087 9902 12098 9948
rect 11563 9834 12098 9902
rect 11563 9788 11927 9834
rect 11973 9788 12041 9834
rect 12087 9788 12098 9834
rect 11563 9720 12098 9788
rect 11563 9674 11927 9720
rect 11973 9674 12041 9720
rect 12087 9674 12098 9720
rect 11563 9606 12098 9674
rect 11563 9560 11927 9606
rect 11973 9560 12041 9606
rect 12087 9560 12098 9606
rect 11563 9492 12098 9560
rect 11563 9446 11927 9492
rect 11973 9446 12041 9492
rect 12087 9446 12098 9492
rect 11563 9378 12098 9446
rect 11563 9332 11927 9378
rect 11973 9332 12041 9378
rect 12087 9332 12098 9378
rect 11563 9264 12098 9332
rect 11563 9218 11927 9264
rect 11973 9218 12041 9264
rect 12087 9218 12098 9264
rect 11563 9150 12098 9218
rect 11563 9104 11927 9150
rect 11973 9104 12041 9150
rect 12087 9104 12098 9150
rect 11563 9036 12098 9104
rect 11563 8990 11927 9036
rect 11973 8990 12041 9036
rect 12087 8990 12098 9036
rect 11563 8922 12098 8990
rect 11563 8876 11927 8922
rect 11973 8876 12041 8922
rect 12087 8876 12098 8922
rect 11563 8808 12098 8876
rect 11563 8762 11927 8808
rect 11973 8762 12041 8808
rect 12087 8762 12098 8808
rect 11563 8694 12098 8762
rect 11563 8648 11927 8694
rect 11973 8648 12041 8694
rect 12087 8648 12098 8694
rect 11563 8580 12098 8648
rect 11563 8534 11927 8580
rect 11973 8534 12041 8580
rect 12087 8534 12098 8580
rect 11563 8466 12098 8534
rect 11563 8420 11927 8466
rect 11973 8420 12041 8466
rect 12087 8420 12098 8466
rect 11563 8352 12098 8420
rect 11563 8306 11927 8352
rect 11973 8306 12041 8352
rect 12087 8306 12098 8352
rect 11563 8238 12098 8306
rect 11563 8192 11927 8238
rect 11973 8192 12041 8238
rect 12087 8192 12098 8238
rect 11563 8124 12098 8192
rect 11563 8078 11927 8124
rect 11973 8078 12041 8124
rect 12087 8078 12098 8124
rect 11563 8010 12098 8078
rect 11563 7964 11927 8010
rect 11973 7964 12041 8010
rect 12087 7964 12098 8010
rect 11563 7896 12098 7964
rect 11563 7850 11927 7896
rect 11973 7850 12041 7896
rect 12087 7850 12098 7896
rect 11563 7782 12098 7850
rect 11563 7736 11927 7782
rect 11973 7736 12041 7782
rect 12087 7736 12098 7782
rect 11563 7668 12098 7736
rect 11563 7622 11927 7668
rect 11973 7622 12041 7668
rect 12087 7622 12098 7668
rect 11563 7554 12098 7622
rect 11563 7508 11927 7554
rect 11973 7508 12041 7554
rect 12087 7508 12098 7554
rect 11563 7440 12098 7508
rect 11563 7394 11927 7440
rect 11973 7394 12041 7440
rect 12087 7394 12098 7440
rect 11563 7326 12098 7394
rect 11563 7280 11927 7326
rect 11973 7280 12041 7326
rect 12087 7280 12098 7326
rect 11563 7212 12098 7280
rect 11563 7166 11927 7212
rect 11973 7166 12041 7212
rect 12087 7166 12098 7212
rect 11563 7098 12098 7166
rect 11563 7052 11927 7098
rect 11973 7052 12041 7098
rect 12087 7052 12098 7098
rect 11563 6984 12098 7052
rect 11563 6938 11927 6984
rect 11973 6938 12041 6984
rect 12087 6938 12098 6984
rect 11563 6870 12098 6938
rect 11563 6824 11927 6870
rect 11973 6824 12041 6870
rect 12087 6824 12098 6870
rect 11563 6756 12098 6824
rect 11563 6710 11927 6756
rect 11973 6710 12041 6756
rect 12087 6710 12098 6756
rect 11563 6642 12098 6710
rect 11563 6596 11927 6642
rect 11973 6596 12041 6642
rect 12087 6596 12098 6642
rect 11563 6528 12098 6596
rect 11563 6482 11927 6528
rect 11973 6482 12041 6528
rect 12087 6482 12098 6528
rect 11563 6414 12098 6482
rect 11563 6368 11927 6414
rect 11973 6368 12041 6414
rect 12087 6368 12098 6414
rect 11563 6300 12098 6368
rect 11563 6254 11927 6300
rect 11973 6254 12041 6300
rect 12087 6254 12098 6300
rect 11563 6186 12098 6254
rect 11563 6140 11927 6186
rect 11973 6140 12041 6186
rect 12087 6140 12098 6186
rect 11563 6072 12098 6140
rect 11563 6026 11927 6072
rect 11973 6026 12041 6072
rect 12087 6026 12098 6072
rect 11563 5958 12098 6026
rect 11563 5912 11927 5958
rect 11973 5912 12041 5958
rect 12087 5912 12098 5958
rect 11563 5844 12098 5912
rect 11563 5798 11927 5844
rect 11973 5798 12041 5844
rect 12087 5798 12098 5844
rect 11563 5730 12098 5798
rect 11563 5684 11927 5730
rect 11973 5684 12041 5730
rect 12087 5684 12098 5730
rect 11563 5616 12098 5684
rect 11563 5570 11927 5616
rect 11973 5570 12041 5616
rect 12087 5570 12098 5616
rect 11563 5502 12098 5570
rect 11563 5456 11927 5502
rect 11973 5456 12041 5502
rect 12087 5456 12098 5502
rect 11563 5388 12098 5456
rect 11563 5376 11927 5388
rect 11506 5342 11927 5376
rect 11973 5342 12041 5388
rect 12087 5342 12098 5388
rect 11506 5339 12098 5342
rect 2222 5306 4138 5317
rect 2222 5279 2233 5306
rect 355 5260 2233 5279
rect 4127 5260 4138 5306
rect 355 5249 4138 5260
rect 4658 5306 6574 5317
rect 4658 5260 4669 5306
rect 6563 5260 6574 5306
rect 4658 5249 6574 5260
rect 7094 5306 9010 5317
rect 7094 5260 7105 5306
rect 8999 5260 9010 5306
rect 7094 5249 9010 5260
rect 9530 5306 11446 5317
rect 9530 5260 9541 5306
rect 11435 5260 11446 5306
rect 9530 5249 11446 5260
rect 355 5117 11446 5249
rect 11916 5274 12098 5339
rect 11916 5228 11927 5274
rect 11973 5228 12041 5274
rect 12087 5228 12098 5274
rect 11916 5160 12098 5228
rect -3742 4395 -3666 4442
rect 355 4395 423 5117
rect 11916 5114 11927 5160
rect 11973 5114 12041 5160
rect 12087 5114 12098 5160
rect 1576 5046 1758 5067
rect 1576 5000 1587 5046
rect 1633 5000 1701 5046
rect 1747 5000 1758 5046
rect 1576 4944 1758 5000
rect 11916 5046 12098 5114
rect 11916 5000 11927 5046
rect 11973 5000 12041 5046
rect 12087 5000 12098 5046
rect 11916 4944 12098 5000
rect 1576 4932 12098 4944
rect 1576 4886 1587 4932
rect 1633 4886 1701 4932
rect 1747 4886 1855 4932
rect 1901 4886 1969 4932
rect 2015 4886 2083 4932
rect 2129 4886 2197 4932
rect 2243 4886 2311 4932
rect 2357 4886 2425 4932
rect 2471 4886 2539 4932
rect 2585 4886 2653 4932
rect 2699 4886 2767 4932
rect 2813 4886 2881 4932
rect 2927 4886 2995 4932
rect 3041 4886 3109 4932
rect 3155 4886 3223 4932
rect 3269 4886 3337 4932
rect 3383 4886 3451 4932
rect 3497 4886 3565 4932
rect 3611 4886 3679 4932
rect 3725 4886 3793 4932
rect 3839 4886 3907 4932
rect 3953 4886 4021 4932
rect 4067 4886 4135 4932
rect 4181 4886 4249 4932
rect 4295 4886 4363 4932
rect 4409 4886 4477 4932
rect 4523 4886 4591 4932
rect 4637 4886 4705 4932
rect 4751 4886 4819 4932
rect 4865 4886 4933 4932
rect 4979 4886 5047 4932
rect 5093 4886 5161 4932
rect 5207 4886 5275 4932
rect 5321 4886 5389 4932
rect 5435 4886 5503 4932
rect 5549 4886 5617 4932
rect 5663 4886 5731 4932
rect 5777 4886 5845 4932
rect 5891 4886 5959 4932
rect 6005 4886 6073 4932
rect 6119 4886 6187 4932
rect 6233 4886 6301 4932
rect 6347 4886 6415 4932
rect 6461 4886 6529 4932
rect 6575 4886 6643 4932
rect 6689 4886 6757 4932
rect 6803 4886 6871 4932
rect 6917 4886 6985 4932
rect 7031 4886 7099 4932
rect 7145 4886 7213 4932
rect 7259 4886 7327 4932
rect 7373 4886 7441 4932
rect 7487 4886 7555 4932
rect 7601 4886 7669 4932
rect 7715 4886 7783 4932
rect 7829 4886 7897 4932
rect 7943 4886 8011 4932
rect 8057 4886 8125 4932
rect 8171 4886 8239 4932
rect 8285 4886 8353 4932
rect 8399 4886 8467 4932
rect 8513 4886 8581 4932
rect 8627 4886 8695 4932
rect 8741 4886 8809 4932
rect 8855 4886 8923 4932
rect 8969 4886 9037 4932
rect 9083 4886 9151 4932
rect 9197 4886 9265 4932
rect 9311 4886 9379 4932
rect 9425 4886 9493 4932
rect 9539 4886 9607 4932
rect 9653 4886 9721 4932
rect 9767 4886 9835 4932
rect 9881 4886 9949 4932
rect 9995 4886 10063 4932
rect 10109 4886 10177 4932
rect 10223 4886 10291 4932
rect 10337 4886 10405 4932
rect 10451 4886 10519 4932
rect 10565 4886 10633 4932
rect 10679 4886 10747 4932
rect 10793 4886 10861 4932
rect 10907 4886 10975 4932
rect 11021 4886 11089 4932
rect 11135 4886 11203 4932
rect 11249 4886 11317 4932
rect 11363 4886 11431 4932
rect 11477 4886 11545 4932
rect 11591 4886 11659 4932
rect 11705 4886 11773 4932
rect 11819 4886 11927 4932
rect 11973 4886 12041 4932
rect 12087 4886 12098 4932
rect 1576 4818 12098 4886
rect 1576 4772 1587 4818
rect 1633 4772 1701 4818
rect 1747 4772 1855 4818
rect 1901 4772 1969 4818
rect 2015 4772 2083 4818
rect 2129 4772 2197 4818
rect 2243 4772 2311 4818
rect 2357 4772 2425 4818
rect 2471 4772 2539 4818
rect 2585 4772 2653 4818
rect 2699 4772 2767 4818
rect 2813 4772 2881 4818
rect 2927 4772 2995 4818
rect 3041 4772 3109 4818
rect 3155 4772 3223 4818
rect 3269 4772 3337 4818
rect 3383 4772 3451 4818
rect 3497 4772 3565 4818
rect 3611 4772 3679 4818
rect 3725 4772 3793 4818
rect 3839 4772 3907 4818
rect 3953 4772 4021 4818
rect 4067 4772 4135 4818
rect 4181 4772 4249 4818
rect 4295 4772 4363 4818
rect 4409 4772 4477 4818
rect 4523 4772 4591 4818
rect 4637 4772 4705 4818
rect 4751 4772 4819 4818
rect 4865 4772 4933 4818
rect 4979 4772 5047 4818
rect 5093 4772 5161 4818
rect 5207 4772 5275 4818
rect 5321 4772 5389 4818
rect 5435 4772 5503 4818
rect 5549 4772 5617 4818
rect 5663 4772 5731 4818
rect 5777 4772 5845 4818
rect 5891 4772 5959 4818
rect 6005 4772 6073 4818
rect 6119 4772 6187 4818
rect 6233 4772 6301 4818
rect 6347 4772 6415 4818
rect 6461 4772 6529 4818
rect 6575 4772 6643 4818
rect 6689 4772 6757 4818
rect 6803 4772 6871 4818
rect 6917 4772 6985 4818
rect 7031 4772 7099 4818
rect 7145 4772 7213 4818
rect 7259 4772 7327 4818
rect 7373 4772 7441 4818
rect 7487 4772 7555 4818
rect 7601 4772 7669 4818
rect 7715 4772 7783 4818
rect 7829 4772 7897 4818
rect 7943 4772 8011 4818
rect 8057 4772 8125 4818
rect 8171 4772 8239 4818
rect 8285 4772 8353 4818
rect 8399 4772 8467 4818
rect 8513 4772 8581 4818
rect 8627 4772 8695 4818
rect 8741 4772 8809 4818
rect 8855 4772 8923 4818
rect 8969 4772 9037 4818
rect 9083 4772 9151 4818
rect 9197 4772 9265 4818
rect 9311 4772 9379 4818
rect 9425 4772 9493 4818
rect 9539 4772 9607 4818
rect 9653 4772 9721 4818
rect 9767 4772 9835 4818
rect 9881 4772 9949 4818
rect 9995 4772 10063 4818
rect 10109 4772 10177 4818
rect 10223 4772 10291 4818
rect 10337 4772 10405 4818
rect 10451 4772 10519 4818
rect 10565 4772 10633 4818
rect 10679 4772 10747 4818
rect 10793 4772 10861 4818
rect 10907 4772 10975 4818
rect 11021 4772 11089 4818
rect 11135 4772 11203 4818
rect 11249 4772 11317 4818
rect 11363 4772 11431 4818
rect 11477 4772 11545 4818
rect 11591 4772 11659 4818
rect 11705 4772 11773 4818
rect 11819 4772 11927 4818
rect 11973 4772 12041 4818
rect 12087 4772 12098 4818
rect 1576 4760 12098 4772
rect -3742 4384 -3296 4395
rect -3742 4338 -3727 4384
rect -3681 4338 -3397 4384
rect -3351 4338 -3296 4384
rect -3742 4327 -3296 4338
rect -3172 4384 -2736 4395
rect -3172 4338 -3117 4384
rect -3071 4338 -2837 4384
rect -2791 4338 -2736 4384
rect -3172 4327 -2736 4338
rect -2612 4384 -2176 4395
rect -2612 4338 -2557 4384
rect -2511 4338 -2277 4384
rect -2231 4338 -2176 4384
rect -2612 4327 -2176 4338
rect -2052 4384 -1616 4395
rect -2052 4338 -1997 4384
rect -1951 4338 -1717 4384
rect -1671 4338 -1616 4384
rect -2052 4327 -1616 4338
rect -1492 4384 -1056 4395
rect -1492 4338 -1437 4384
rect -1391 4338 -1157 4384
rect -1111 4338 -1056 4384
rect -1492 4327 -1056 4338
rect -932 4384 -496 4395
rect -932 4338 -877 4384
rect -831 4338 -597 4384
rect -551 4338 -496 4384
rect -932 4327 -496 4338
rect -372 4384 423 4395
rect -372 4338 -317 4384
rect -271 4338 423 4384
rect -372 4327 423 4338
rect -3742 4280 -3666 4327
rect -3742 4234 -3727 4280
rect -3681 4234 -3666 4280
rect -3742 4176 -3666 4234
rect -3742 4130 -3727 4176
rect -3681 4130 -3666 4176
rect -3742 4083 -3666 4130
rect 2 4176 70 4267
rect 2 4130 13 4176
rect 59 4130 70 4176
rect 2 4083 70 4130
rect -3742 4072 70 4083
rect -3742 4026 -3727 4072
rect -3681 4026 -3573 4072
rect -3527 4026 -3469 4072
rect -3423 4026 -3365 4072
rect -3319 4026 -3261 4072
rect -3215 4026 -3157 4072
rect -3111 4026 -3053 4072
rect -3007 4026 -2949 4072
rect -2903 4026 -2845 4072
rect -2799 4026 -2741 4072
rect -2695 4026 -2637 4072
rect -2591 4026 -2533 4072
rect -2487 4026 -2429 4072
rect -2383 4026 -2325 4072
rect -2279 4026 -2221 4072
rect -2175 4026 -2117 4072
rect -2071 4026 -2013 4072
rect -1967 4026 -1909 4072
rect -1863 4026 -1805 4072
rect -1759 4026 -1701 4072
rect -1655 4026 -1597 4072
rect -1551 4026 -1493 4072
rect -1447 4026 -1389 4072
rect -1343 4026 -1285 4072
rect -1239 4026 -1181 4072
rect -1135 4026 -1077 4072
rect -1031 4026 -973 4072
rect -927 4026 -869 4072
rect -823 4026 -765 4072
rect -719 4026 -661 4072
rect -615 4026 -557 4072
rect -511 4026 -453 4072
rect -407 4026 -349 4072
rect -303 4026 -245 4072
rect -199 4026 -141 4072
rect -95 4026 13 4072
rect 59 4026 70 4072
rect -3742 4015 70 4026
use M1_NWELL_CDNS_40661954729280  M1_NWELL_CDNS_40661954729280_0
timestamp 1698431365
transform -1 0 -3704 0 -1 10809
box 0 0 1 1
use M1_NWELL_CDNS_40661954729281  M1_NWELL_CDNS_40661954729281_0
timestamp 1698431365
transform 0 -1 -1834 1 0 17569
box 0 0 1 1
use M1_NWELL_CDNS_40661954729281  M1_NWELL_CDNS_40661954729281_1
timestamp 1698431365
transform 0 -1 -1834 1 0 4049
box 0 0 1 1
use M1_PSUB_CDNS_40661954729136  M1_PSUB_CDNS_40661954729136_0
timestamp 1698431365
transform 1 0 12007 0 1 10894
box 0 0 1 1
use M1_PSUB_CDNS_40661954729138  M1_PSUB_CDNS_40661954729138_0
timestamp 1698431365
transform 0 -1 6837 1 0 10845
box 0 0 1 1
use M1_PSUB_CDNS_40661954729138  M1_PSUB_CDNS_40661954729138_1
timestamp 1698431365
transform 0 -1 6837 1 0 4852
box 0 0 1 1
use M1_PSUB_CDNS_40661954729138  M1_PSUB_CDNS_40661954729138_2
timestamp 1698431365
transform 0 -1 6837 1 0 16936
box 0 0 1 1
use nmoscap_6p0_CDNS_406619547290  nmoscap_6p0_CDNS_406619547290_0
timestamp 1698431365
transform 1 0 2180 0 -1 10339
box 0 0 1 1
use nmoscap_6p0_CDNS_406619547290  nmoscap_6p0_CDNS_406619547290_1
timestamp 1698431365
transform 1 0 4616 0 -1 10339
box 0 0 1 1
use nmoscap_6p0_CDNS_406619547290  nmoscap_6p0_CDNS_406619547290_2
timestamp 1698431365
transform 1 0 7052 0 -1 10339
box 0 0 1 1
use nmoscap_6p0_CDNS_406619547290  nmoscap_6p0_CDNS_406619547290_3
timestamp 1698431365
transform 1 0 9488 0 -1 10339
box 0 0 1 1
use nmoscap_6p0_CDNS_406619547290  nmoscap_6p0_CDNS_406619547290_4
timestamp 1698431365
transform 1 0 9488 0 1 11351
box 0 0 1 1
use nmoscap_6p0_CDNS_406619547290  nmoscap_6p0_CDNS_406619547290_5
timestamp 1698431365
transform 1 0 7052 0 1 11351
box 0 0 1 1
use nmoscap_6p0_CDNS_406619547290  nmoscap_6p0_CDNS_406619547290_6
timestamp 1698431365
transform 1 0 4616 0 1 11351
box 0 0 1 1
use nmoscap_6p0_CDNS_406619547290  nmoscap_6p0_CDNS_406619547290_7
timestamp 1698431365
transform 1 0 2180 0 1 11351
box 0 0 1 1
use ppolyf_u_CDNS_406619547295  ppolyf_u_CDNS_406619547295_0
timestamp 1698431365
transform 0 1 -1774 1 0 4325
box 0 0 1 1
use ppolyf_u_CDNS_406619547295  ppolyf_u_CDNS_406619547295_1
timestamp 1698431365
transform 0 1 -654 1 0 4325
box 0 0 1 1
use ppolyf_u_CDNS_406619547295  ppolyf_u_CDNS_406619547295_2
timestamp 1698431365
transform 0 1 -2334 1 0 4325
box 0 0 1 1
use ppolyf_u_CDNS_406619547295  ppolyf_u_CDNS_406619547295_3
timestamp 1698431365
transform 0 1 -1214 1 0 4325
box 0 0 1 1
use ppolyf_u_CDNS_406619547295  ppolyf_u_CDNS_406619547295_4
timestamp 1698431365
transform 0 1 -2894 1 0 4325
box 0 0 1 1
use ppolyf_u_CDNS_406619547295  ppolyf_u_CDNS_406619547295_5
timestamp 1698431365
transform 0 1 -374 -1 0 17300
box 0 0 1 1
use ppolyf_u_CDNS_406619547295  ppolyf_u_CDNS_406619547295_6
timestamp 1698431365
transform 0 1 -934 -1 0 17300
box 0 0 1 1
use ppolyf_u_CDNS_406619547295  ppolyf_u_CDNS_406619547295_7
timestamp 1698431365
transform 0 1 -3174 -1 0 17300
box 0 0 1 1
use ppolyf_u_CDNS_406619547295  ppolyf_u_CDNS_406619547295_8
timestamp 1698431365
transform 0 1 -1494 -1 0 17300
box 0 0 1 1
use ppolyf_u_CDNS_406619547295  ppolyf_u_CDNS_406619547295_9
timestamp 1698431365
transform 0 1 -2614 -1 0 17300
box 0 0 1 1
use ppolyf_u_CDNS_406619547295  ppolyf_u_CDNS_406619547295_10
timestamp 1698431365
transform 0 1 -2054 -1 0 17300
box 0 0 1 1
use ppolyf_u_CDNS_406619547295  ppolyf_u_CDNS_406619547295_11
timestamp 1698431365
transform 0 -1 -3294 1 0 4325
box 0 0 1 1
<< labels >>
rlabel metal1 s 984 16493 984 16493 4 VRC
port 1 nsew
rlabel metal1 s -3704 4447 -3704 4447 4 VPLUS
port 2 nsew
rlabel metal1 s 6835 10844 6835 10844 4 VMINUS
port 3 nsew
<< properties >>
string GDS_END 6644804
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 6618804
<< end >>
