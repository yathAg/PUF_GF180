magic
tech gf180mcuD
timestamp 1698431365
<< properties >>
string GDS_END 17158894
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 17089066
<< end >>
