magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
use M1_NACTIVE$$203393068_256x8m81  M1_NACTIVE$$203393068_256x8m81_0
timestamp 1698431365
transform 1 0 14063 0 1 29759
box 0 0 1 1
use M1_NWELL$$204218412_256x8m81  M1_NWELL$$204218412_256x8m81_0
timestamp 1698431365
transform -1 0 25568 0 1 29686
box 0 0 1 1
use M1_NWELL$$204218412_256x8m81  M1_NWELL$$204218412_256x8m81_1
timestamp 1698431365
transform 1 0 2200 0 1 29686
box 0 0 1 1
use M1_PACTIVE$$204148780_256x8m81  M1_PACTIVE$$204148780_256x8m81_0
timestamp 1698431365
transform 1 0 11463 0 1 29759
box 0 0 1 1
use M1_PACTIVE$$204148780_256x8m81  M1_PACTIVE$$204148780_256x8m81_1
timestamp 1698431365
transform 1 0 21475 0 1 29759
box 0 0 1 1
use M1_PACTIVE$$204148780_256x8m81  M1_PACTIVE$$204148780_256x8m81_2
timestamp 1698431365
transform 1 0 4390 0 1 29759
box 0 0 1 1
use M1_PACTIVE$$204149804_256x8m81  M1_PACTIVE$$204149804_256x8m81_0
timestamp 1698431365
transform 1 0 15860 0 1 29759
box 0 0 1 1
use M1_POLY2$$204150828_256x8m81  M1_POLY2$$204150828_256x8m81_0
timestamp 1698431365
transform 1 0 9381 0 1 29448
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_0
timestamp 1698431365
transform 1 0 15413 0 1 29741
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_0
timestamp 1698431365
transform 0 -1 13712 1 0 29693
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_1
timestamp 1698431365
transform 1 0 15625 0 1 29401
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_2
timestamp 1698431365
transform 1 0 18313 0 1 29436
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_3
timestamp 1698431365
transform 1 0 12040 0 1 29361
box 0 0 1 1
use M2_M1$$201262124_256x8m81  M2_M1$$201262124_256x8m81_0
timestamp 1698431365
transform 1 0 13701 0 1 29691
box 0 0 1 1
use M2_M1$$204138540_256x8m81  M2_M1$$204138540_256x8m81_0
timestamp 1698431365
transform 1 0 10402 0 1 29448
box 0 0 1 1
use M2_M1$$204138540_256x8m81  M2_M1$$204138540_256x8m81_1
timestamp 1698431365
transform 1 0 14059 0 1 29752
box 0 0 1 1
use M2_M1$$204139564_256x8m81  M2_M1$$204139564_256x8m81_0
timestamp 1698431365
transform 1 0 11601 0 1 29705
box 0 0 1 1
use M2_M1$$204140588_256x8m81  M2_M1$$204140588_256x8m81_0
timestamp 1698431365
transform 1 0 12359 0 1 29217
box 0 0 1 1
use M2_M1$$204141612_256x8m81  M2_M1$$204141612_256x8m81_0
timestamp 1698431365
transform 1 0 15126 0 1 29752
box 0 0 1 1
use M2_M1$$204141612_256x8m81  M2_M1$$204141612_256x8m81_1
timestamp 1698431365
transform 1 0 20177 0 1 29680
box 0 0 1 1
use M2_M1$$204141612_256x8m81  M2_M1$$204141612_256x8m81_2
timestamp 1698431365
transform 1 0 20177 0 1 29217
box 0 0 1 1
use M2_M1$$204220460_256x8m81  M2_M1$$204220460_256x8m81_0
timestamp 1698431365
transform 1 0 6792 0 1 29217
box 0 0 1 1
use M2_M1$$204220460_256x8m81  M2_M1$$204220460_256x8m81_1
timestamp 1698431365
transform 1 0 22430 0 1 29217
box 0 0 1 1
use M2_M1$$204220460_256x8m81  M2_M1$$204220460_256x8m81_2
timestamp 1698431365
transform 1 0 4399 0 1 29219
box 0 0 1 1
use M2_M1$$204220460_256x8m81  M2_M1$$204220460_256x8m81_3
timestamp 1698431365
transform 1 0 6792 0 1 29680
box 0 0 1 1
use M2_M1$$204221484_256x8m81  M2_M1$$204221484_256x8m81_0
timestamp 1698431365
transform -1 0 25612 0 1 29700
box 0 0 1 1
use M2_M1$$204221484_256x8m81  M2_M1$$204221484_256x8m81_1
timestamp 1698431365
transform 1 0 2156 0 1 29700
box 0 0 1 1
use M2_M1$$204222508_256x8m81  M2_M1$$204222508_256x8m81_0
timestamp 1698431365
transform 1 0 21486 0 1 29700
box 0 0 1 1
use M2_M1$$204222508_256x8m81  M2_M1$$204222508_256x8m81_1
timestamp 1698431365
transform 1 0 5639 0 1 29700
box 0 0 1 1
use M3_M2$$204142636_256x8m81  M3_M2$$204142636_256x8m81_0
timestamp 1698431365
transform 1 0 5639 0 1 29700
box 0 0 1 1
use M3_M2$$204142636_256x8m81  M3_M2$$204142636_256x8m81_1
timestamp 1698431365
transform 1 0 8250 0 1 29217
box 0 0 1 1
use M3_M2$$204142636_256x8m81  M3_M2$$204142636_256x8m81_2
timestamp 1698431365
transform 1 0 21486 0 1 29700
box 0 0 1 1
use M3_M2$$204143660_256x8m81  M3_M2$$204143660_256x8m81_0
timestamp 1698431365
transform 1 0 11601 0 1 29700
box 0 0 1 1
use M3_M2$$204144684_256x8m81  M3_M2$$204144684_256x8m81_0
timestamp 1698431365
transform 1 0 22430 0 1 29217
box 0 0 1 1
use M3_M2$$204144684_256x8m81  M3_M2$$204144684_256x8m81_1
timestamp 1698431365
transform 1 0 4399 0 1 29219
box 0 0 1 1
use M3_M2$$204145708_256x8m81  M3_M2$$204145708_256x8m81_0
timestamp 1698431365
transform 1 0 12359 0 1 29217
box 0 0 1 1
use M3_M2$$204146732_256x8m81  M3_M2$$204146732_256x8m81_0
timestamp 1698431365
transform 1 0 14059 0 1 29210
box 0 0 1 1
use M3_M2$$204147756_256x8m81  M3_M2$$204147756_256x8m81_0
timestamp 1698431365
transform 1 0 12339 0 1 28800
box 0 0 1 1
use nmos_1p2$$204213292_R90_256x8m81  nmos_1p2$$204213292_R90_256x8m81_0
timestamp 1698431365
transform 0 -1 6346 1 0 29303
box -31 0 -30 1
use nmos_1p2$$204215340_256x8m81  nmos_1p2$$204215340_256x8m81_0
timestamp 1698431365
transform 0 -1 13604 -1 0 29362
box -31 0 -30 1
use nmos_5p04310590878199_256x8m81  nmos_5p04310590878199_256x8m81_0
timestamp 1698431365
transform 0 -1 23346 1 0 29272
box 0 0 1 1
use nmos_5p043105908781111_256x8m81  nmos_5p043105908781111_256x8m81_0
timestamp 1698431365
transform 0 -1 16283 1 0 29272
box 0 0 1 1
use nmos_5p043105908781111_256x8m81  nmos_5p043105908781111_256x8m81_1
timestamp 1698431365
transform 0 -1 11913 1 0 29272
box 0 0 1 1
use pmos_1p2$$204216364_256x8m81  pmos_1p2$$204216364_256x8m81_0
timestamp 1698431365
transform 0 -1 20950 1 0 29303
box -31 0 -30 1
use pmos_1p2$$204216364_256x8m81  pmos_1p2$$204216364_256x8m81_1
timestamp 1698431365
transform 0 -1 9245 1 0 29303
box -31 0 -30 1
use pmos_1p2$$204217388_256x8m81  pmos_1p2$$204217388_256x8m81_0
timestamp 1698431365
transform 0 -1 11004 1 0 29303
box -31 0 -30 1
use pmos_5p043105908781101_256x8m81  pmos_5p043105908781101_256x8m81_0
timestamp 1698431365
transform 0 -1 15304 1 0 29272
box 0 0 1 1
use pmos_5p043105908781101_256x8m81  pmos_5p043105908781101_256x8m81_1
timestamp 1698431365
transform 0 -1 17974 1 0 29272
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_0
timestamp 1698431365
transform 0 -1 2203 -1 0 28950
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_1
timestamp 1698431365
transform 0 -1 2203 -1 0 27150
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_2
timestamp 1698431365
transform 0 -1 2203 -1 0 25350
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_3
timestamp 1698431365
transform 0 -1 2203 -1 0 23550
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_4
timestamp 1698431365
transform 0 -1 2203 -1 0 21750
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_5
timestamp 1698431365
transform 0 -1 2203 -1 0 19950
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_6
timestamp 1698431365
transform 0 -1 2203 -1 0 18150
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_7
timestamp 1698431365
transform 0 -1 2203 -1 0 16350
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_8
timestamp 1698431365
transform 0 -1 2203 -1 0 14550
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_9
timestamp 1698431365
transform 0 -1 2203 -1 0 12750
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_10
timestamp 1698431365
transform 0 -1 2203 -1 0 10950
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_11
timestamp 1698431365
transform 0 -1 2203 -1 0 9150
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_12
timestamp 1698431365
transform 0 -1 2203 -1 0 7350
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_13
timestamp 1698431365
transform 0 -1 2203 -1 0 5550
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_14
timestamp 1698431365
transform 0 -1 2203 -1 0 3750
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_15
timestamp 1698431365
transform 0 -1 2203 -1 0 1950
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_16
timestamp 1698431365
transform 0 1 25566 -1 0 28950
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_17
timestamp 1698431365
transform 0 1 25566 -1 0 27150
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_18
timestamp 1698431365
transform 0 1 25566 -1 0 25350
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_19
timestamp 1698431365
transform 0 1 25566 -1 0 23550
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_20
timestamp 1698431365
transform 0 1 25566 -1 0 21750
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_21
timestamp 1698431365
transform 0 1 25566 -1 0 19950
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_22
timestamp 1698431365
transform 0 1 25566 -1 0 18150
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_23
timestamp 1698431365
transform 0 1 25566 -1 0 16350
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_24
timestamp 1698431365
transform 0 1 25566 -1 0 14550
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_25
timestamp 1698431365
transform 0 1 25566 -1 0 12750
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_26
timestamp 1698431365
transform 0 1 25566 -1 0 10950
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_27
timestamp 1698431365
transform 0 1 25566 -1 0 9150
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_28
timestamp 1698431365
transform 0 1 25566 -1 0 7350
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_29
timestamp 1698431365
transform 0 1 25566 -1 0 5550
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_30
timestamp 1698431365
transform 0 1 25566 -1 0 3750
box 0 0 1 1
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_31
timestamp 1698431365
transform 0 1 25566 -1 0 1950
box 0 0 1 1
use pmoscap_W2_5_R270_256x8m81  pmoscap_W2_5_R270_256x8m81_0
timestamp 1698431365
transform 0 -1 2203 -1 0 29850
box 150 220 1051 2048
use pmoscap_W2_5_R270_256x8m81  pmoscap_W2_5_R270_256x8m81_1
timestamp 1698431365
transform 0 1 25566 -1 0 29850
box 150 220 1051 2048
use xdec32_256x8m81  xdec32_256x8m81_0
timestamp 1698431365
transform 1 0 1726 0 1 0
box 1426 -1 22889 28801
<< properties >>
string GDS_END 2364970
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 2346198
<< end >>
