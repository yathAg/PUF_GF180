magic
tech gf180mcuD
magscale 1 10
timestamp 1698431365
use M1_NACTIVE$$204211244_128x8m81  M1_NACTIVE$$204211244_128x8m81_0
timestamp 1698431365
transform 1 0 605 0 1 220
box 0 0 1 1
use M1_PACTIVE$$20421_R270_128x8m81  M1_PACTIVE$$20421_R270_128x8m81_0
timestamp 1698431365
transform 1 0 605 0 1 2047
box 0 0 1 1
use M1_POLY2$$204395564_128x8m81  M1_POLY2$$204395564_128x8m81_0
timestamp 1698431365
transform 1 0 601 0 1 1741
box 0 0 1 1
use M2_M1$$204396588_R270_128x8m81  M2_M1$$204396588_R270_128x8m81_0
timestamp 1698431365
transform 1 0 150 0 1 955
box 0 0 1 1
use M2_M1$$204396588_R270_128x8m81  M2_M1$$204396588_R270_128x8m81_1
timestamp 1698431365
transform 1 0 1050 0 1 955
box 0 0 1 1
use M3_M2$$204397612_R270_128x8m81  M3_M2$$204397612_R270_128x8m81_0
timestamp 1698431365
transform 1 0 1050 0 1 955
box 0 0 1 1
<< properties >>
string GDS_END 1686232
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 1683472
<< end >>
