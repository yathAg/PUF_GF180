magic
tech gf180mcuB
magscale 1 10
timestamp 1698431365
use npn_10p00x10p00_0  npn_10p00x10p00_0_0
timestamp 1698431365
transform 1 0 1320 0 1 1320
box -1264 -1264 3264 3264
<< labels >>
flabel metal1 s 1325 1325 1325 1325 0 FreeSans 200 0 0 0 I1_default_E
port 3 nsew
flabel metal1 s 61 4505 61 4505 0 FreeSans 200 0 0 0 I1_default_S
port 4 nsew
flabel metal1 s 4505 61 4505 61 0 FreeSans 200 0 0 0 I1_default_S
port 4 nsew
flabel metal1 s 4005 61 4005 61 0 FreeSans 200 0 0 0 I1_default_S
port 4 nsew
flabel metal1 s 61 61 61 61 0 FreeSans 200 0 0 0 I1_default_S
port 4 nsew
flabel metal1 s 61 61 61 61 0 FreeSans 200 0 0 0 I1_default_S
port 4 nsew
flabel metal1 s 1029 1029 1029 1029 0 FreeSans 200 0 0 0 I1_default_C
port 1 nsew
flabel metal1 s 3537 1029 3537 1029 0 FreeSans 200 0 0 0 I1_default_C
port 1 nsew
flabel metal1 s 1029 3537 1029 3537 0 FreeSans 200 0 0 0 I1_default_C
port 1 nsew
flabel metal1 s 1177 1177 1177 1177 0 FreeSans 200 0 0 0 I1_default_B
port 2 nsew
flabel metal1 s 3389 1177 3389 1177 0 FreeSans 200 0 0 0 I1_default_B
port 2 nsew
flabel metal1 s 1177 3389 1177 3389 0 FreeSans 200 0 0 0 I1_default_B
port 2 nsew
<< properties >>
string GDS_END 38826
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_pr/gds/npn_10p00x10p00.gds
string GDS_START 37916
string device primitive
<< end >>
