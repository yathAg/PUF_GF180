magic
tech gf180mcuB
magscale 1 10
timestamp 1698431365
<< isosubstrate >>
rect -496 -83 693 2575
<< nwell >>
rect -247 1551 693 2575
rect 1033 1281 4434 2575
<< mvnmos >>
rect -92 263 48 1063
rect 152 263 292 1063
rect 1655 270 1795 520
rect 1899 270 2039 520
rect 2559 270 2699 570
rect 2803 270 2943 570
rect 3047 270 3187 570
rect 3291 270 3431 570
rect 3535 270 3675 570
rect 3779 270 3919 570
<< mvpmos >>
rect 152 1811 292 2211
rect 1411 1522 1551 2022
rect 1655 1522 1795 2022
rect 1899 1522 2039 2022
rect 2143 1522 2283 2022
rect 2559 1522 2699 2222
rect 2803 1522 2943 2222
rect 3047 1522 3187 2222
rect 3291 1522 3431 2222
rect 3535 1522 3675 2222
rect 3779 1522 3919 2222
<< mvndiff >>
rect -180 1050 -92 1063
rect -180 1004 -167 1050
rect -121 1004 -92 1050
rect -180 946 -92 1004
rect -180 900 -167 946
rect -121 900 -92 946
rect -180 842 -92 900
rect -180 796 -167 842
rect -121 796 -92 842
rect -180 738 -92 796
rect -180 692 -167 738
rect -121 692 -92 738
rect -180 634 -92 692
rect -180 588 -167 634
rect -121 588 -92 634
rect -180 530 -92 588
rect -180 484 -167 530
rect -121 484 -92 530
rect -180 426 -92 484
rect -180 380 -167 426
rect -121 380 -92 426
rect -180 322 -92 380
rect -180 276 -167 322
rect -121 276 -92 322
rect -180 263 -92 276
rect 48 1050 152 1063
rect 48 1004 77 1050
rect 123 1004 152 1050
rect 48 946 152 1004
rect 48 900 77 946
rect 123 900 152 946
rect 48 842 152 900
rect 48 796 77 842
rect 123 796 152 842
rect 48 738 152 796
rect 48 692 77 738
rect 123 692 152 738
rect 48 634 152 692
rect 48 588 77 634
rect 123 588 152 634
rect 48 530 152 588
rect 48 484 77 530
rect 123 484 152 530
rect 48 426 152 484
rect 48 380 77 426
rect 123 380 152 426
rect 48 322 152 380
rect 48 276 77 322
rect 123 276 152 322
rect 48 263 152 276
rect 292 1050 380 1063
rect 292 1004 321 1050
rect 367 1004 380 1050
rect 292 946 380 1004
rect 292 900 321 946
rect 367 900 380 946
rect 292 842 380 900
rect 292 796 321 842
rect 367 796 380 842
rect 292 738 380 796
rect 292 692 321 738
rect 367 692 380 738
rect 292 634 380 692
rect 292 588 321 634
rect 367 588 380 634
rect 292 530 380 588
rect 292 484 321 530
rect 367 484 380 530
rect 292 426 380 484
rect 292 380 321 426
rect 367 380 380 426
rect 292 322 380 380
rect 292 276 321 322
rect 367 276 380 322
rect 292 263 380 276
rect 2471 557 2559 570
rect 1567 507 1655 520
rect 1567 461 1580 507
rect 1626 461 1655 507
rect 1567 329 1655 461
rect 1567 283 1580 329
rect 1626 283 1655 329
rect 1567 270 1655 283
rect 1795 507 1899 520
rect 1795 461 1824 507
rect 1870 461 1899 507
rect 1795 329 1899 461
rect 1795 283 1824 329
rect 1870 283 1899 329
rect 1795 270 1899 283
rect 2039 507 2127 520
rect 2039 461 2068 507
rect 2114 461 2127 507
rect 2039 329 2127 461
rect 2039 283 2068 329
rect 2114 283 2127 329
rect 2039 270 2127 283
rect 2471 511 2484 557
rect 2530 511 2559 557
rect 2471 443 2559 511
rect 2471 397 2484 443
rect 2530 397 2559 443
rect 2471 329 2559 397
rect 2471 283 2484 329
rect 2530 283 2559 329
rect 2471 270 2559 283
rect 2699 557 2803 570
rect 2699 511 2728 557
rect 2774 511 2803 557
rect 2699 443 2803 511
rect 2699 397 2728 443
rect 2774 397 2803 443
rect 2699 329 2803 397
rect 2699 283 2728 329
rect 2774 283 2803 329
rect 2699 270 2803 283
rect 2943 557 3047 570
rect 2943 511 2972 557
rect 3018 511 3047 557
rect 2943 443 3047 511
rect 2943 397 2972 443
rect 3018 397 3047 443
rect 2943 329 3047 397
rect 2943 283 2972 329
rect 3018 283 3047 329
rect 2943 270 3047 283
rect 3187 557 3291 570
rect 3187 511 3216 557
rect 3262 511 3291 557
rect 3187 443 3291 511
rect 3187 397 3216 443
rect 3262 397 3291 443
rect 3187 329 3291 397
rect 3187 283 3216 329
rect 3262 283 3291 329
rect 3187 270 3291 283
rect 3431 557 3535 570
rect 3431 511 3460 557
rect 3506 511 3535 557
rect 3431 443 3535 511
rect 3431 397 3460 443
rect 3506 397 3535 443
rect 3431 329 3535 397
rect 3431 283 3460 329
rect 3506 283 3535 329
rect 3431 270 3535 283
rect 3675 557 3779 570
rect 3675 511 3704 557
rect 3750 511 3779 557
rect 3675 443 3779 511
rect 3675 397 3704 443
rect 3750 397 3779 443
rect 3675 329 3779 397
rect 3675 283 3704 329
rect 3750 283 3779 329
rect 3675 270 3779 283
rect 3919 557 4007 570
rect 3919 511 3948 557
rect 3994 511 4007 557
rect 3919 443 4007 511
rect 3919 397 3948 443
rect 3994 397 4007 443
rect 3919 329 4007 397
rect 3919 283 3948 329
rect 3994 283 4007 329
rect 3919 270 4007 283
<< mvpdiff >>
rect 64 2198 152 2211
rect 64 2152 77 2198
rect 123 2152 152 2198
rect 64 2089 152 2152
rect 64 2043 77 2089
rect 123 2043 152 2089
rect 64 1980 152 2043
rect 64 1934 77 1980
rect 123 1934 152 1980
rect 64 1870 152 1934
rect 64 1824 77 1870
rect 123 1824 152 1870
rect 64 1811 152 1824
rect 292 2198 380 2211
rect 292 2152 321 2198
rect 367 2152 380 2198
rect 292 2089 380 2152
rect 292 2043 321 2089
rect 367 2043 380 2089
rect 292 1980 380 2043
rect 292 1934 321 1980
rect 367 1934 380 1980
rect 292 1870 380 1934
rect 292 1824 321 1870
rect 367 1824 380 1870
rect 292 1811 380 1824
rect 2471 2209 2559 2222
rect 2471 2163 2484 2209
rect 2530 2163 2559 2209
rect 2471 2105 2559 2163
rect 2471 2059 2484 2105
rect 2530 2059 2559 2105
rect 1323 2009 1411 2022
rect 1323 1963 1336 2009
rect 1382 1963 1411 2009
rect 1323 1902 1411 1963
rect 1323 1856 1336 1902
rect 1382 1856 1411 1902
rect 1323 1795 1411 1856
rect 1323 1749 1336 1795
rect 1382 1749 1411 1795
rect 1323 1688 1411 1749
rect 1323 1642 1336 1688
rect 1382 1642 1411 1688
rect 1323 1581 1411 1642
rect 1323 1535 1336 1581
rect 1382 1535 1411 1581
rect 1323 1522 1411 1535
rect 1551 2009 1655 2022
rect 1551 1963 1580 2009
rect 1626 1963 1655 2009
rect 1551 1902 1655 1963
rect 1551 1856 1580 1902
rect 1626 1856 1655 1902
rect 1551 1795 1655 1856
rect 1551 1749 1580 1795
rect 1626 1749 1655 1795
rect 1551 1688 1655 1749
rect 1551 1642 1580 1688
rect 1626 1642 1655 1688
rect 1551 1581 1655 1642
rect 1551 1535 1580 1581
rect 1626 1535 1655 1581
rect 1551 1522 1655 1535
rect 1795 2009 1899 2022
rect 1795 1963 1824 2009
rect 1870 1963 1899 2009
rect 1795 1902 1899 1963
rect 1795 1856 1824 1902
rect 1870 1856 1899 1902
rect 1795 1795 1899 1856
rect 1795 1749 1824 1795
rect 1870 1749 1899 1795
rect 1795 1688 1899 1749
rect 1795 1642 1824 1688
rect 1870 1642 1899 1688
rect 1795 1581 1899 1642
rect 1795 1535 1824 1581
rect 1870 1535 1899 1581
rect 1795 1522 1899 1535
rect 2039 2009 2143 2022
rect 2039 1963 2068 2009
rect 2114 1963 2143 2009
rect 2039 1902 2143 1963
rect 2039 1856 2068 1902
rect 2114 1856 2143 1902
rect 2039 1795 2143 1856
rect 2039 1749 2068 1795
rect 2114 1749 2143 1795
rect 2039 1688 2143 1749
rect 2039 1642 2068 1688
rect 2114 1642 2143 1688
rect 2039 1581 2143 1642
rect 2039 1535 2068 1581
rect 2114 1535 2143 1581
rect 2039 1522 2143 1535
rect 2283 2009 2371 2022
rect 2283 1963 2312 2009
rect 2358 1963 2371 2009
rect 2283 1902 2371 1963
rect 2283 1856 2312 1902
rect 2358 1856 2371 1902
rect 2283 1795 2371 1856
rect 2283 1749 2312 1795
rect 2358 1749 2371 1795
rect 2283 1688 2371 1749
rect 2283 1642 2312 1688
rect 2358 1642 2371 1688
rect 2283 1581 2371 1642
rect 2283 1535 2312 1581
rect 2358 1535 2371 1581
rect 2283 1522 2371 1535
rect 2471 2001 2559 2059
rect 2471 1955 2484 2001
rect 2530 1955 2559 2001
rect 2471 1896 2559 1955
rect 2471 1850 2484 1896
rect 2530 1850 2559 1896
rect 2471 1791 2559 1850
rect 2471 1745 2484 1791
rect 2530 1745 2559 1791
rect 2471 1686 2559 1745
rect 2471 1640 2484 1686
rect 2530 1640 2559 1686
rect 2471 1581 2559 1640
rect 2471 1535 2484 1581
rect 2530 1535 2559 1581
rect 2471 1522 2559 1535
rect 2699 2209 2803 2222
rect 2699 2163 2728 2209
rect 2774 2163 2803 2209
rect 2699 2105 2803 2163
rect 2699 2059 2728 2105
rect 2774 2059 2803 2105
rect 2699 2001 2803 2059
rect 2699 1955 2728 2001
rect 2774 1955 2803 2001
rect 2699 1896 2803 1955
rect 2699 1850 2728 1896
rect 2774 1850 2803 1896
rect 2699 1791 2803 1850
rect 2699 1745 2728 1791
rect 2774 1745 2803 1791
rect 2699 1686 2803 1745
rect 2699 1640 2728 1686
rect 2774 1640 2803 1686
rect 2699 1581 2803 1640
rect 2699 1535 2728 1581
rect 2774 1535 2803 1581
rect 2699 1522 2803 1535
rect 2943 2209 3047 2222
rect 2943 2163 2972 2209
rect 3018 2163 3047 2209
rect 2943 2105 3047 2163
rect 2943 2059 2972 2105
rect 3018 2059 3047 2105
rect 2943 2001 3047 2059
rect 2943 1955 2972 2001
rect 3018 1955 3047 2001
rect 2943 1896 3047 1955
rect 2943 1850 2972 1896
rect 3018 1850 3047 1896
rect 2943 1791 3047 1850
rect 2943 1745 2972 1791
rect 3018 1745 3047 1791
rect 2943 1686 3047 1745
rect 2943 1640 2972 1686
rect 3018 1640 3047 1686
rect 2943 1581 3047 1640
rect 2943 1535 2972 1581
rect 3018 1535 3047 1581
rect 2943 1522 3047 1535
rect 3187 2209 3291 2222
rect 3187 2163 3216 2209
rect 3262 2163 3291 2209
rect 3187 2105 3291 2163
rect 3187 2059 3216 2105
rect 3262 2059 3291 2105
rect 3187 2001 3291 2059
rect 3187 1955 3216 2001
rect 3262 1955 3291 2001
rect 3187 1896 3291 1955
rect 3187 1850 3216 1896
rect 3262 1850 3291 1896
rect 3187 1791 3291 1850
rect 3187 1745 3216 1791
rect 3262 1745 3291 1791
rect 3187 1686 3291 1745
rect 3187 1640 3216 1686
rect 3262 1640 3291 1686
rect 3187 1581 3291 1640
rect 3187 1535 3216 1581
rect 3262 1535 3291 1581
rect 3187 1522 3291 1535
rect 3431 2209 3535 2222
rect 3431 2163 3460 2209
rect 3506 2163 3535 2209
rect 3431 2105 3535 2163
rect 3431 2059 3460 2105
rect 3506 2059 3535 2105
rect 3431 2001 3535 2059
rect 3431 1955 3460 2001
rect 3506 1955 3535 2001
rect 3431 1896 3535 1955
rect 3431 1850 3460 1896
rect 3506 1850 3535 1896
rect 3431 1791 3535 1850
rect 3431 1745 3460 1791
rect 3506 1745 3535 1791
rect 3431 1686 3535 1745
rect 3431 1640 3460 1686
rect 3506 1640 3535 1686
rect 3431 1581 3535 1640
rect 3431 1535 3460 1581
rect 3506 1535 3535 1581
rect 3431 1522 3535 1535
rect 3675 2209 3779 2222
rect 3675 2163 3704 2209
rect 3750 2163 3779 2209
rect 3675 2105 3779 2163
rect 3675 2059 3704 2105
rect 3750 2059 3779 2105
rect 3675 2001 3779 2059
rect 3675 1955 3704 2001
rect 3750 1955 3779 2001
rect 3675 1896 3779 1955
rect 3675 1850 3704 1896
rect 3750 1850 3779 1896
rect 3675 1791 3779 1850
rect 3675 1745 3704 1791
rect 3750 1745 3779 1791
rect 3675 1686 3779 1745
rect 3675 1640 3704 1686
rect 3750 1640 3779 1686
rect 3675 1581 3779 1640
rect 3675 1535 3704 1581
rect 3750 1535 3779 1581
rect 3675 1522 3779 1535
rect 3919 2209 4007 2222
rect 3919 2163 3948 2209
rect 3994 2163 4007 2209
rect 3919 2105 4007 2163
rect 3919 2059 3948 2105
rect 3994 2059 4007 2105
rect 3919 2001 4007 2059
rect 3919 1955 3948 2001
rect 3994 1955 4007 2001
rect 3919 1896 4007 1955
rect 3919 1850 3948 1896
rect 3994 1850 4007 1896
rect 3919 1791 4007 1850
rect 3919 1745 3948 1791
rect 3994 1745 4007 1791
rect 3919 1686 4007 1745
rect 3919 1640 3948 1686
rect 3994 1640 4007 1686
rect 3919 1581 4007 1640
rect 3919 1535 3948 1581
rect 3994 1535 4007 1581
rect 3919 1522 4007 1535
<< mvndiffc >>
rect -167 1004 -121 1050
rect -167 900 -121 946
rect -167 796 -121 842
rect -167 692 -121 738
rect -167 588 -121 634
rect -167 484 -121 530
rect -167 380 -121 426
rect -167 276 -121 322
rect 77 1004 123 1050
rect 77 900 123 946
rect 77 796 123 842
rect 77 692 123 738
rect 77 588 123 634
rect 77 484 123 530
rect 77 380 123 426
rect 77 276 123 322
rect 321 1004 367 1050
rect 321 900 367 946
rect 321 796 367 842
rect 321 692 367 738
rect 321 588 367 634
rect 321 484 367 530
rect 321 380 367 426
rect 321 276 367 322
rect 1580 461 1626 507
rect 1580 283 1626 329
rect 1824 461 1870 507
rect 1824 283 1870 329
rect 2068 461 2114 507
rect 2068 283 2114 329
rect 2484 511 2530 557
rect 2484 397 2530 443
rect 2484 283 2530 329
rect 2728 511 2774 557
rect 2728 397 2774 443
rect 2728 283 2774 329
rect 2972 511 3018 557
rect 2972 397 3018 443
rect 2972 283 3018 329
rect 3216 511 3262 557
rect 3216 397 3262 443
rect 3216 283 3262 329
rect 3460 511 3506 557
rect 3460 397 3506 443
rect 3460 283 3506 329
rect 3704 511 3750 557
rect 3704 397 3750 443
rect 3704 283 3750 329
rect 3948 511 3994 557
rect 3948 397 3994 443
rect 3948 283 3994 329
<< mvpdiffc >>
rect 77 2152 123 2198
rect 77 2043 123 2089
rect 77 1934 123 1980
rect 77 1824 123 1870
rect 321 2152 367 2198
rect 321 2043 367 2089
rect 321 1934 367 1980
rect 321 1824 367 1870
rect 2484 2163 2530 2209
rect 2484 2059 2530 2105
rect 1336 1963 1382 2009
rect 1336 1856 1382 1902
rect 1336 1749 1382 1795
rect 1336 1642 1382 1688
rect 1336 1535 1382 1581
rect 1580 1963 1626 2009
rect 1580 1856 1626 1902
rect 1580 1749 1626 1795
rect 1580 1642 1626 1688
rect 1580 1535 1626 1581
rect 1824 1963 1870 2009
rect 1824 1856 1870 1902
rect 1824 1749 1870 1795
rect 1824 1642 1870 1688
rect 1824 1535 1870 1581
rect 2068 1963 2114 2009
rect 2068 1856 2114 1902
rect 2068 1749 2114 1795
rect 2068 1642 2114 1688
rect 2068 1535 2114 1581
rect 2312 1963 2358 2009
rect 2312 1856 2358 1902
rect 2312 1749 2358 1795
rect 2312 1642 2358 1688
rect 2312 1535 2358 1581
rect 2484 1955 2530 2001
rect 2484 1850 2530 1896
rect 2484 1745 2530 1791
rect 2484 1640 2530 1686
rect 2484 1535 2530 1581
rect 2728 2163 2774 2209
rect 2728 2059 2774 2105
rect 2728 1955 2774 2001
rect 2728 1850 2774 1896
rect 2728 1745 2774 1791
rect 2728 1640 2774 1686
rect 2728 1535 2774 1581
rect 2972 2163 3018 2209
rect 2972 2059 3018 2105
rect 2972 1955 3018 2001
rect 2972 1850 3018 1896
rect 2972 1745 3018 1791
rect 2972 1640 3018 1686
rect 2972 1535 3018 1581
rect 3216 2163 3262 2209
rect 3216 2059 3262 2105
rect 3216 1955 3262 2001
rect 3216 1850 3262 1896
rect 3216 1745 3262 1791
rect 3216 1640 3262 1686
rect 3216 1535 3262 1581
rect 3460 2163 3506 2209
rect 3460 2059 3506 2105
rect 3460 1955 3506 2001
rect 3460 1850 3506 1896
rect 3460 1745 3506 1791
rect 3460 1640 3506 1686
rect 3460 1535 3506 1581
rect 3704 2163 3750 2209
rect 3704 2059 3750 2105
rect 3704 1955 3750 2001
rect 3704 1850 3750 1896
rect 3704 1745 3750 1791
rect 3704 1640 3750 1686
rect 3704 1535 3750 1581
rect 3948 2163 3994 2209
rect 3948 2059 3994 2105
rect 3948 1955 3994 2001
rect 3948 1850 3994 1896
rect 3948 1745 3994 1791
rect 3948 1640 3994 1686
rect 3948 1535 3994 1581
<< psubdiff >>
rect -443 1196 -353 1218
rect -443 22 -421 1196
rect -375 90 -353 1196
rect 520 1196 610 1218
rect 520 90 542 1196
rect -375 68 542 90
rect 471 22 542 68
rect 588 22 610 1196
rect -443 0 610 22
rect 1116 1008 1206 1030
rect 1116 22 1138 1008
rect 1184 90 1206 1008
rect 4244 1008 4334 1030
rect 4244 90 4266 1008
rect 1184 68 4266 90
rect 1184 22 1292 68
rect 4158 22 4266 68
rect 4312 22 4334 1008
rect 1116 0 4334 22
<< nsubdiff >>
rect -164 2470 610 2492
rect -164 1766 -142 2470
rect -96 2424 12 2470
rect 434 2424 542 2470
rect -96 2402 542 2424
rect -96 1766 -74 2402
rect -164 1744 -74 1766
rect 520 1766 542 2402
rect 588 1766 610 2470
rect 520 1744 610 1766
rect 1116 2470 4300 2492
rect 1116 1484 1138 2470
rect 1184 2424 1260 2470
rect 4126 2424 4232 2470
rect 1184 2402 4232 2424
rect 1184 1484 1206 2402
rect 1116 1462 1206 1484
rect 4210 1484 4232 2402
rect 4278 1484 4300 2470
rect 4210 1462 4300 1484
<< psubdiffcont >>
rect -421 68 -375 1196
rect -421 22 471 68
rect 542 22 588 1196
rect 1138 22 1184 1008
rect 1292 22 4158 68
rect 4266 22 4312 1008
<< nsubdiffcont >>
rect -142 1766 -96 2470
rect 12 2424 434 2470
rect 542 1766 588 2470
rect 1138 1484 1184 2470
rect 1260 2424 4126 2470
rect 4232 1484 4278 2470
<< polysilicon >>
rect 152 2211 292 2255
rect -92 1412 48 1431
rect -92 1272 -47 1412
rect -1 1272 48 1412
rect -92 1063 48 1272
rect 152 1412 292 1811
rect 2559 2222 2699 2266
rect 2803 2222 2943 2266
rect 3047 2222 3187 2266
rect 3291 2222 3431 2266
rect 3535 2222 3675 2266
rect 3779 2222 3919 2266
rect 1411 2022 1551 2066
rect 1655 2022 1795 2066
rect 1899 2022 2039 2066
rect 2143 2022 2283 2066
rect 152 1272 199 1412
rect 245 1272 292 1412
rect 152 1063 292 1272
rect 1411 1265 1551 1522
rect -92 219 48 263
rect 152 219 292 263
rect 1411 1125 1458 1265
rect 1504 1125 1551 1265
rect 1411 1106 1551 1125
rect 1655 1265 1795 1522
rect 1655 1125 1702 1265
rect 1748 1125 1795 1265
rect 1655 520 1795 1125
rect 1899 1265 2039 1522
rect 1899 1125 1946 1265
rect 1992 1125 2039 1265
rect 1899 520 2039 1125
rect 2143 1265 2283 1522
rect 2143 1125 2190 1265
rect 2236 1125 2283 1265
rect 2143 1106 2283 1125
rect 2559 1265 2699 1522
rect 2559 1125 2606 1265
rect 2652 1125 2699 1265
rect 2559 570 2699 1125
rect 2803 1265 2943 1522
rect 2803 1125 2850 1265
rect 2896 1125 2943 1265
rect 2803 570 2943 1125
rect 3047 1265 3187 1522
rect 3047 1125 3094 1265
rect 3140 1125 3187 1265
rect 3047 570 3187 1125
rect 3291 1265 3431 1522
rect 3291 1125 3338 1265
rect 3384 1125 3431 1265
rect 3291 570 3431 1125
rect 3535 1265 3675 1522
rect 3535 1125 3582 1265
rect 3628 1125 3675 1265
rect 3535 570 3675 1125
rect 3779 1265 3919 1522
rect 3779 1125 3826 1265
rect 3872 1125 3919 1265
rect 3779 570 3919 1125
rect 1655 226 1795 270
rect 1899 226 2039 270
rect 2559 226 2699 270
rect 2803 226 2943 270
rect 3047 226 3187 270
rect 3291 226 3431 270
rect 3535 226 3675 270
rect 3779 226 3919 270
<< polycontact >>
rect -47 1272 -1 1412
rect 199 1272 245 1412
rect 1458 1125 1504 1265
rect 1702 1125 1748 1265
rect 1946 1125 1992 1265
rect 2190 1125 2236 1265
rect 2606 1125 2652 1265
rect 2850 1125 2896 1265
rect 3094 1125 3140 1265
rect 3338 1125 3384 1265
rect 3582 1125 3628 1265
rect 3826 1125 3872 1265
<< metal1 >>
rect -153 2470 599 2481
rect -153 1766 -142 2470
rect -96 2424 12 2470
rect 434 2424 542 2470
rect -96 2413 542 2424
rect -96 1766 -85 2413
rect 62 2198 138 2413
rect 62 2152 77 2198
rect 123 2152 138 2198
rect 62 2089 138 2152
rect 62 2043 77 2089
rect 123 2043 138 2089
rect 62 1980 138 2043
rect 62 1934 77 1980
rect 123 1934 138 1980
rect 62 1870 138 1934
rect 62 1824 77 1870
rect 123 1824 138 1870
rect 62 1811 138 1824
rect 306 2198 382 2211
rect 306 2152 321 2198
rect 367 2152 382 2198
rect 306 2089 382 2152
rect 306 2043 321 2089
rect 367 2043 382 2089
rect 306 1980 382 2043
rect 306 1934 321 1980
rect 367 1934 382 1980
rect 306 1870 382 1934
rect 306 1824 321 1870
rect 367 1824 382 1870
rect -153 1755 -85 1766
rect 306 1441 382 1824
rect 531 1766 542 2413
rect 588 1766 599 2470
rect 531 1755 599 1766
rect 1127 2470 4289 2481
rect 1127 1484 1138 2470
rect 1184 2424 1260 2470
rect 4126 2424 4232 2470
rect 1184 2413 4232 2424
rect 1184 1484 1195 2413
rect 1321 2009 1397 2413
rect 1321 1963 1336 2009
rect 1382 1963 1397 2009
rect 1321 1902 1397 1963
rect 1580 2009 1626 2022
rect 1580 1958 1626 1963
rect 1809 2009 1885 2413
rect 1809 1963 1824 2009
rect 1870 1963 1885 2009
rect 1321 1856 1336 1902
rect 1382 1856 1397 1902
rect 1321 1795 1397 1856
rect 1321 1749 1336 1795
rect 1382 1749 1397 1795
rect 1321 1688 1397 1749
rect 1321 1642 1336 1688
rect 1382 1642 1397 1688
rect 1321 1581 1397 1642
rect 1321 1535 1336 1581
rect 1382 1535 1397 1581
rect 1321 1522 1397 1535
rect 1565 1902 1641 1958
rect 1565 1856 1580 1902
rect 1626 1856 1641 1902
rect 1565 1795 1641 1856
rect 1565 1749 1580 1795
rect 1626 1749 1641 1795
rect 1565 1688 1641 1749
rect 1565 1642 1580 1688
rect 1626 1642 1641 1688
rect 1565 1581 1641 1642
rect 1565 1535 1580 1581
rect 1626 1535 1641 1581
rect 1127 1473 1195 1484
rect 1565 1442 1641 1535
rect 1809 1902 1885 1963
rect 2068 2009 2114 2022
rect 2068 1958 2114 1963
rect 2297 2009 2373 2413
rect 2297 1963 2312 2009
rect 2358 1963 2373 2009
rect 1809 1856 1824 1902
rect 1870 1856 1885 1902
rect 1809 1795 1885 1856
rect 1809 1749 1824 1795
rect 1870 1749 1885 1795
rect 1809 1688 1885 1749
rect 1809 1642 1824 1688
rect 1870 1642 1885 1688
rect 1809 1581 1885 1642
rect 1809 1535 1824 1581
rect 1870 1535 1885 1581
rect 1809 1522 1885 1535
rect 2053 1902 2129 1958
rect 2053 1856 2068 1902
rect 2114 1856 2129 1902
rect 2053 1795 2129 1856
rect 2053 1749 2068 1795
rect 2114 1749 2129 1795
rect 2053 1688 2129 1749
rect 2053 1642 2068 1688
rect 2114 1642 2129 1688
rect 2053 1581 2129 1642
rect 2053 1535 2068 1581
rect 2114 1535 2129 1581
rect 2053 1442 2129 1535
rect 2297 1902 2373 1963
rect 2297 1856 2312 1902
rect 2358 1856 2373 1902
rect 2297 1795 2373 1856
rect 2297 1749 2312 1795
rect 2358 1749 2373 1795
rect 2297 1688 2373 1749
rect 2297 1642 2312 1688
rect 2358 1642 2373 1688
rect 2297 1581 2373 1642
rect 2297 1535 2312 1581
rect 2358 1535 2373 1581
rect 2297 1522 2373 1535
rect 2469 2209 2545 2413
rect 2469 2163 2484 2209
rect 2530 2163 2545 2209
rect 2469 2105 2545 2163
rect 2469 2059 2484 2105
rect 2530 2059 2545 2105
rect 2469 2001 2545 2059
rect 2469 1955 2484 2001
rect 2530 1955 2545 2001
rect 2469 1896 2545 1955
rect 2469 1850 2484 1896
rect 2530 1850 2545 1896
rect 2469 1791 2545 1850
rect 2469 1745 2484 1791
rect 2530 1745 2545 1791
rect 2469 1686 2545 1745
rect 2469 1640 2484 1686
rect 2530 1640 2545 1686
rect 2469 1581 2545 1640
rect 2469 1535 2484 1581
rect 2530 1535 2545 1581
rect 2469 1522 2545 1535
rect 2713 2209 2789 2222
rect 2713 2163 2728 2209
rect 2774 2163 2789 2209
rect 2713 2105 2789 2163
rect 2713 2059 2728 2105
rect 2774 2059 2789 2105
rect 2713 2001 2789 2059
rect 2713 1955 2728 2001
rect 2774 1955 2789 2001
rect 2713 1896 2789 1955
rect 2713 1850 2728 1896
rect 2774 1850 2789 1896
rect 2713 1791 2789 1850
rect 2713 1745 2728 1791
rect 2774 1745 2789 1791
rect 2713 1686 2789 1745
rect 2713 1640 2728 1686
rect 2774 1640 2789 1686
rect 2713 1581 2789 1640
rect 2713 1535 2728 1581
rect 2774 1535 2789 1581
rect 2713 1442 2789 1535
rect 2957 2209 3033 2413
rect 2957 2163 2972 2209
rect 3018 2163 3033 2209
rect 2957 2105 3033 2163
rect 2957 2059 2972 2105
rect 3018 2059 3033 2105
rect 2957 2001 3033 2059
rect 2957 1955 2972 2001
rect 3018 1955 3033 2001
rect 2957 1896 3033 1955
rect 2957 1850 2972 1896
rect 3018 1850 3033 1896
rect 2957 1791 3033 1850
rect 2957 1745 2972 1791
rect 3018 1745 3033 1791
rect 2957 1686 3033 1745
rect 2957 1640 2972 1686
rect 3018 1640 3033 1686
rect 2957 1581 3033 1640
rect 2957 1535 2972 1581
rect 3018 1535 3033 1581
rect 2957 1522 3033 1535
rect 3201 2209 3277 2222
rect 3201 2163 3216 2209
rect 3262 2163 3277 2209
rect 3201 2105 3277 2163
rect 3201 2059 3216 2105
rect 3262 2059 3277 2105
rect 3201 2001 3277 2059
rect 3201 1955 3216 2001
rect 3262 1955 3277 2001
rect 3201 1896 3277 1955
rect 3201 1850 3216 1896
rect 3262 1850 3277 1896
rect 3201 1791 3277 1850
rect 3201 1745 3216 1791
rect 3262 1745 3277 1791
rect 3201 1686 3277 1745
rect 3201 1640 3216 1686
rect 3262 1640 3277 1686
rect 3201 1581 3277 1640
rect 3201 1535 3216 1581
rect 3262 1535 3277 1581
rect 3201 1442 3277 1535
rect 3445 2209 3521 2413
rect 3445 2163 3460 2209
rect 3506 2163 3521 2209
rect 3445 2105 3521 2163
rect 3445 2059 3460 2105
rect 3506 2059 3521 2105
rect 3445 2001 3521 2059
rect 3445 1955 3460 2001
rect 3506 1955 3521 2001
rect 3445 1896 3521 1955
rect 3445 1850 3460 1896
rect 3506 1850 3521 1896
rect 3445 1791 3521 1850
rect 3445 1745 3460 1791
rect 3506 1745 3521 1791
rect 3445 1686 3521 1745
rect 3445 1640 3460 1686
rect 3506 1640 3521 1686
rect 3445 1581 3521 1640
rect 3445 1535 3460 1581
rect 3506 1535 3521 1581
rect 3445 1522 3521 1535
rect 3689 2209 3765 2222
rect 3689 2163 3704 2209
rect 3750 2163 3765 2209
rect 3689 2105 3765 2163
rect 3689 2059 3704 2105
rect 3750 2059 3765 2105
rect 3689 2001 3765 2059
rect 3689 1955 3704 2001
rect 3750 1955 3765 2001
rect 3689 1896 3765 1955
rect 3689 1850 3704 1896
rect 3750 1850 3765 1896
rect 3689 1791 3765 1850
rect 3689 1745 3704 1791
rect 3750 1745 3765 1791
rect 3689 1686 3765 1745
rect 3689 1640 3704 1686
rect 3750 1640 3765 1686
rect 3689 1581 3765 1640
rect 3689 1535 3704 1581
rect 3750 1535 3765 1581
rect 3689 1442 3765 1535
rect 3933 2209 4009 2413
rect 3933 2163 3948 2209
rect 3994 2163 4009 2209
rect 3933 2105 4009 2163
rect 3933 2059 3948 2105
rect 3994 2059 4009 2105
rect 3933 2001 4009 2059
rect 3933 1955 3948 2001
rect 3994 1955 4009 2001
rect 3933 1896 4009 1955
rect 3933 1850 3948 1896
rect 3994 1850 4009 1896
rect 3933 1791 4009 1850
rect 3933 1745 3948 1791
rect 3994 1745 4009 1791
rect 3933 1686 4009 1745
rect 3933 1640 3948 1686
rect 3994 1640 4009 1686
rect 3933 1581 4009 1640
rect 3933 1535 3948 1581
rect 3994 1535 4009 1581
rect 3933 1522 4009 1535
rect 4221 1484 4232 2413
rect 4278 1484 4289 2470
rect 4221 1473 4289 1484
rect -58 1412 10 1423
rect -58 1272 -47 1412
rect -1 1272 10 1412
rect -58 1261 10 1272
rect 188 1412 256 1423
rect 188 1272 199 1412
rect 245 1272 256 1412
rect 188 1261 256 1272
rect 306 1341 937 1441
rect 1565 1366 2667 1442
rect 2713 1366 4066 1442
rect -432 1196 -364 1207
rect -432 22 -421 1196
rect -375 79 -364 1196
rect -167 1050 -121 1063
rect -167 946 -121 1004
rect 77 1050 123 1063
rect 77 990 123 1004
rect 306 1050 382 1341
rect 837 1276 937 1341
rect 2591 1276 2667 1366
rect 837 1265 2247 1276
rect 306 1004 321 1050
rect 367 1004 382 1050
rect -167 842 -121 900
rect -167 738 -121 796
rect -182 696 -167 708
rect 62 946 138 990
rect 62 900 77 946
rect 123 900 138 946
rect 62 842 138 900
rect 62 796 77 842
rect 123 796 138 842
rect 62 738 138 796
rect -121 696 -106 708
rect -182 332 -170 696
rect -118 332 -106 696
rect -182 322 -106 332
rect -182 320 -167 322
rect -121 320 -106 322
rect 62 692 77 738
rect 123 692 138 738
rect 62 634 138 692
rect 62 588 77 634
rect 123 588 138 634
rect 62 530 138 588
rect 62 484 77 530
rect 123 484 138 530
rect 62 426 138 484
rect 62 380 77 426
rect 123 380 138 426
rect 62 322 138 380
rect -167 263 -121 276
rect 62 276 77 322
rect 123 276 138 322
rect 62 79 138 276
rect 306 946 382 1004
rect 306 900 321 946
rect 367 900 382 946
rect 306 842 382 900
rect 306 796 321 842
rect 367 796 382 842
rect 306 738 382 796
rect 306 696 321 738
rect 367 696 382 738
rect 306 332 318 696
rect 370 332 382 696
rect 306 322 382 332
rect 306 276 321 322
rect 367 276 382 322
rect 306 263 382 276
rect 531 1196 599 1207
rect 531 79 542 1196
rect -375 68 542 79
rect 471 22 542 68
rect 588 22 599 1196
rect 837 1125 1458 1265
rect 1504 1125 1702 1265
rect 1748 1125 1946 1265
rect 1992 1125 2190 1265
rect 2236 1125 2247 1265
rect 837 1114 2247 1125
rect 2591 1265 3883 1276
rect 2591 1125 2606 1265
rect 2652 1125 2850 1265
rect 2896 1125 3094 1265
rect 3140 1125 3338 1265
rect 3384 1125 3582 1265
rect 3628 1125 3826 1265
rect 3872 1125 3883 1265
rect 2591 1114 3883 1125
rect -432 11 599 22
rect 1127 1008 1195 1019
rect 1127 22 1138 1008
rect 1184 79 1195 1008
rect 2591 819 2667 1114
rect 3990 819 4066 1366
rect 1809 743 2667 819
rect 2713 743 4066 819
rect 4255 1008 4323 1019
rect 1580 507 1626 520
rect 1565 461 1580 470
rect 1809 507 1885 743
rect 2469 557 2545 570
rect 1626 461 1641 470
rect 1565 329 1641 461
rect 1565 283 1580 329
rect 1626 283 1641 329
rect 1565 79 1641 283
rect 1809 461 1824 507
rect 1870 461 1885 507
rect 2068 507 2114 520
rect 1809 329 1885 461
rect 1809 283 1824 329
rect 1870 283 1885 329
rect 1809 270 1885 283
rect 2053 461 2068 470
rect 2469 511 2484 557
rect 2530 511 2545 557
rect 2114 461 2129 470
rect 2053 329 2129 461
rect 2053 283 2068 329
rect 2114 283 2129 329
rect 2053 79 2129 283
rect 2469 443 2545 511
rect 2469 397 2484 443
rect 2530 397 2545 443
rect 2469 329 2545 397
rect 2469 283 2484 329
rect 2530 283 2545 329
rect 2469 79 2545 283
rect 2713 557 2789 743
rect 2713 511 2728 557
rect 2774 511 2789 557
rect 2713 443 2789 511
rect 2713 397 2728 443
rect 2774 397 2789 443
rect 2713 329 2789 397
rect 2713 283 2728 329
rect 2774 283 2789 329
rect 2713 270 2789 283
rect 2957 557 3033 570
rect 2957 511 2972 557
rect 3018 511 3033 557
rect 2957 443 3033 511
rect 2957 397 2972 443
rect 3018 397 3033 443
rect 2957 329 3033 397
rect 2957 283 2972 329
rect 3018 283 3033 329
rect 2957 79 3033 283
rect 3201 557 3277 743
rect 3201 511 3216 557
rect 3262 511 3277 557
rect 3201 443 3277 511
rect 3201 397 3216 443
rect 3262 397 3277 443
rect 3201 329 3277 397
rect 3201 283 3216 329
rect 3262 283 3277 329
rect 3201 270 3277 283
rect 3445 557 3521 570
rect 3445 511 3460 557
rect 3506 511 3521 557
rect 3445 443 3521 511
rect 3445 397 3460 443
rect 3506 397 3521 443
rect 3445 329 3521 397
rect 3445 283 3460 329
rect 3506 283 3521 329
rect 3445 79 3521 283
rect 3689 557 3765 743
rect 3689 511 3704 557
rect 3750 511 3765 557
rect 3689 443 3765 511
rect 3689 397 3704 443
rect 3750 397 3765 443
rect 3689 329 3765 397
rect 3689 283 3704 329
rect 3750 283 3765 329
rect 3689 270 3765 283
rect 3931 557 4007 570
rect 3931 511 3948 557
rect 3994 511 4007 557
rect 3931 443 4007 511
rect 3931 397 3948 443
rect 3994 397 4007 443
rect 3931 329 4007 397
rect 3931 283 3948 329
rect 3994 283 4007 329
rect 3931 79 4007 283
rect 4255 79 4266 1008
rect 1184 68 4266 79
rect 1184 22 1292 68
rect 4158 22 4266 68
rect 4312 22 4323 1008
rect 1127 11 4323 22
<< via1 >>
rect -170 692 -167 696
rect -167 692 -121 696
rect -121 692 -118 696
rect -170 634 -118 692
rect -170 588 -167 634
rect -167 588 -121 634
rect -121 588 -118 634
rect -170 530 -118 588
rect -170 484 -167 530
rect -167 484 -121 530
rect -121 484 -118 530
rect -170 426 -118 484
rect -170 380 -167 426
rect -167 380 -121 426
rect -121 380 -118 426
rect -170 332 -118 380
rect 318 692 321 696
rect 321 692 367 696
rect 367 692 370 696
rect 318 634 370 692
rect 318 588 321 634
rect 321 588 367 634
rect 367 588 370 634
rect 318 530 370 588
rect 318 484 321 530
rect 321 484 367 530
rect 367 484 370 530
rect 318 426 370 484
rect 318 380 321 426
rect 321 380 367 426
rect 367 380 370 426
rect 318 332 370 380
<< metal2 >>
rect -182 696 -106 708
rect -182 332 -170 696
rect -118 573 -106 696
rect 306 696 382 708
rect 306 573 318 696
rect -118 435 318 573
rect -118 332 -106 435
rect -182 320 -106 332
rect 306 332 318 435
rect 370 332 382 696
rect 306 320 382 332
use M1_NWELL_CDNS_40661954729411  M1_NWELL_CDNS_40661954729411_0
timestamp 1698431365
transform 1 0 223 0 1 2447
box 0 0 1 1
use M1_NWELL_CDNS_40661954729412  M1_NWELL_CDNS_40661954729412_0
timestamp 1698431365
transform 1 0 4255 0 1 1977
box 0 0 1 1
use M1_NWELL_CDNS_40661954729412  M1_NWELL_CDNS_40661954729412_1
timestamp 1698431365
transform 1 0 1161 0 1 1977
box 0 0 1 1
use M1_NWELL_CDNS_40661954729429  M1_NWELL_CDNS_40661954729429_0
timestamp 1698431365
transform 1 0 2693 0 1 2447
box 0 0 1 1
use M1_NWELL_CDNS_40661954729432  M1_NWELL_CDNS_40661954729432_0
timestamp 1698431365
transform 1 0 565 0 1 2118
box 0 0 1 1
use M1_NWELL_CDNS_40661954729432  M1_NWELL_CDNS_40661954729432_1
timestamp 1698431365
transform 1 0 -119 0 1 2118
box 0 0 1 1
use M1_POLY2_CDNS_40661954729415  M1_POLY2_CDNS_40661954729415_0
timestamp 1698431365
transform 1 0 3849 0 1 1195
box 0 0 1 1
use M1_POLY2_CDNS_40661954729415  M1_POLY2_CDNS_40661954729415_1
timestamp 1698431365
transform 1 0 3605 0 1 1195
box 0 0 1 1
use M1_POLY2_CDNS_40661954729415  M1_POLY2_CDNS_40661954729415_2
timestamp 1698431365
transform 1 0 -24 0 1 1342
box 0 0 1 1
use M1_POLY2_CDNS_40661954729415  M1_POLY2_CDNS_40661954729415_3
timestamp 1698431365
transform 1 0 222 0 1 1342
box 0 0 1 1
use M1_POLY2_CDNS_40661954729415  M1_POLY2_CDNS_40661954729415_4
timestamp 1698431365
transform 1 0 1725 0 1 1195
box 0 0 1 1
use M1_POLY2_CDNS_40661954729415  M1_POLY2_CDNS_40661954729415_5
timestamp 1698431365
transform 1 0 1481 0 1 1195
box 0 0 1 1
use M1_POLY2_CDNS_40661954729415  M1_POLY2_CDNS_40661954729415_6
timestamp 1698431365
transform 1 0 2629 0 1 1195
box 0 0 1 1
use M1_POLY2_CDNS_40661954729415  M1_POLY2_CDNS_40661954729415_7
timestamp 1698431365
transform 1 0 2873 0 1 1195
box 0 0 1 1
use M1_POLY2_CDNS_40661954729415  M1_POLY2_CDNS_40661954729415_8
timestamp 1698431365
transform 1 0 2213 0 1 1195
box 0 0 1 1
use M1_POLY2_CDNS_40661954729415  M1_POLY2_CDNS_40661954729415_9
timestamp 1698431365
transform 1 0 3361 0 1 1195
box 0 0 1 1
use M1_POLY2_CDNS_40661954729415  M1_POLY2_CDNS_40661954729415_10
timestamp 1698431365
transform 1 0 3117 0 1 1195
box 0 0 1 1
use M1_POLY2_CDNS_40661954729415  M1_POLY2_CDNS_40661954729415_11
timestamp 1698431365
transform 1 0 1969 0 1 1195
box 0 0 1 1
use M1_PSUB_CDNS_40661954729413  M1_PSUB_CDNS_40661954729413_0
timestamp 1698431365
transform 1 0 1161 0 -1 515
box 0 0 1 1
use M1_PSUB_CDNS_40661954729413  M1_PSUB_CDNS_40661954729413_1
timestamp 1698431365
transform 1 0 4289 0 -1 515
box 0 0 1 1
use M1_PSUB_CDNS_40661954729428  M1_PSUB_CDNS_40661954729428_0
timestamp 1698431365
transform 1 0 72 0 -1 45
box 0 0 1 1
use M1_PSUB_CDNS_40661954729430  M1_PSUB_CDNS_40661954729430_0
timestamp 1698431365
transform 1 0 565 0 -1 609
box 0 0 1 1
use M1_PSUB_CDNS_40661954729430  M1_PSUB_CDNS_40661954729430_1
timestamp 1698431365
transform 1 0 -398 0 -1 609
box 0 0 1 1
use M1_PSUB_CDNS_40661954729431  M1_PSUB_CDNS_40661954729431_0
timestamp 1698431365
transform 1 0 2725 0 -1 45
box 0 0 1 1
use M2_M1_CDNS_40661954729404  M2_M1_CDNS_40661954729404_0
timestamp 1698431365
transform 1 0 344 0 1 514
box 0 0 1 1
use M2_M1_CDNS_40661954729404  M2_M1_CDNS_40661954729404_1
timestamp 1698431365
transform 1 0 -144 0 1 514
box 0 0 1 1
use nmos_6p0_CDNS_4066195472929  nmos_6p0_CDNS_4066195472929_0
timestamp 1698431365
transform 1 0 -92 0 1 263
box 0 0 1 1
use nmos_6p0_CDNS_4066195472931  nmos_6p0_CDNS_4066195472931_0
timestamp 1698431365
transform 1 0 2559 0 1 270
box 0 0 1 1
use nmos_6p0_CDNS_4066195472932  nmos_6p0_CDNS_4066195472932_0
timestamp 1698431365
transform 1 0 1655 0 1 270
box 0 0 1 1
use pmos_6p0_CDNS_4066195472917  pmos_6p0_CDNS_4066195472917_0
timestamp 1698431365
transform 1 0 152 0 1 1811
box 0 0 1 1
use pmos_6p0_CDNS_4066195472928  pmos_6p0_CDNS_4066195472928_0
timestamp 1698431365
transform 1 0 1411 0 1 1522
box 0 0 1 1
use pmos_6p0_CDNS_4066195472930  pmos_6p0_CDNS_4066195472930_0
timestamp 1698431365
transform 1 0 2559 0 1 1522
box 0 0 1 1
<< labels >>
rlabel metal1 s 2 2452 2 2452 4 DVDD
port 1 nsew
rlabel metal1 s 225 1326 225 1326 4 A
port 2 nsew
rlabel metal1 s 80 45 80 45 4 DVSS
port 3 nsew
rlabel metal1 s 1852 2452 1852 2452 4 VDD
port 4 nsew
rlabel metal1 s 1482 45 1482 45 4 VSS
port 5 nsew
rlabel metal1 s 3512 1200 3512 1200 4 Z
port 6 nsew
rlabel metal1 s -21 1326 -21 1326 4 A
port 2 nsew
<< properties >>
string GDS_END 1465840
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 1459986
string path 80.975 20.475 80.975 6.750 
<< end >>
