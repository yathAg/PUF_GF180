magic
tech gf180mcuB
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 352 758 870
<< pwell >>
rect -86 -86 758 352
<< metal1 >>
rect 0 724 672 844
rect 49 506 95 724
rect 141 424 207 575
rect 253 547 299 676
rect 466 593 534 724
rect 253 472 542 547
rect 141 347 394 424
rect 141 238 207 347
rect 466 301 542 472
rect 273 254 542 301
rect 49 60 95 208
rect 273 136 319 254
rect 497 60 543 208
rect 0 -60 672 60
<< labels >>
rlabel metal1 s 141 238 207 347 6 I
port 1 nsew default input
rlabel metal1 s 141 347 394 424 6 I
port 1 nsew default input
rlabel metal1 s 141 424 207 575 6 I
port 1 nsew default input
rlabel metal1 s 273 136 319 254 6 ZN
port 2 nsew default output
rlabel metal1 s 273 254 542 301 6 ZN
port 2 nsew default output
rlabel metal1 s 466 301 542 472 6 ZN
port 2 nsew default output
rlabel metal1 s 253 472 542 547 6 ZN
port 2 nsew default output
rlabel metal1 s 253 547 299 676 6 ZN
port 2 nsew default output
rlabel metal1 s 466 593 534 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 506 95 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 724 672 844 6 VDD
port 3 nsew power bidirectional abutment
rlabel nwell s -86 352 758 870 6 VNW
port 4 nsew power bidirectional
rlabel pwell s -86 -86 758 352 6 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 0 -60 672 60 8 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 497 60 543 208 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 208 6 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 672 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 820038
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 817426
<< end >>
