magic
tech gf180mcuA
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 407 2550 870
rect -86 352 575 407
rect 943 352 2550 407
<< pwell >>
rect 575 352 943 407
rect -86 -86 2550 352
<< mvnmos >>
rect 124 68 244 232
rect 348 68 468 232
rect 572 68 692 232
rect 1064 68 1184 232
rect 1288 68 1408 232
rect 1512 68 1632 232
rect 1736 68 1856 232
rect 1960 68 2080 232
rect 2184 68 2304 232
<< mvpmos >>
rect 172 527 272 716
rect 376 527 476 716
rect 660 527 760 716
rect 1144 481 1244 716
rect 1348 481 1448 716
rect 1552 481 1652 716
rect 1756 481 1856 716
rect 1960 481 2060 716
rect 2164 481 2264 716
<< mvndiff >>
rect 752 274 824 287
rect 752 232 765 274
rect 36 219 124 232
rect 36 173 49 219
rect 95 173 124 219
rect 36 68 124 173
rect 244 128 348 232
rect 244 82 273 128
rect 319 82 348 128
rect 244 68 348 82
rect 468 169 572 232
rect 468 123 497 169
rect 543 123 572 169
rect 468 68 572 123
rect 692 228 765 232
rect 811 228 824 274
rect 692 68 824 228
rect 932 95 1064 232
rect 932 49 945 95
rect 991 68 1064 95
rect 1184 219 1288 232
rect 1184 173 1213 219
rect 1259 173 1288 219
rect 1184 68 1288 173
rect 1408 127 1512 232
rect 1408 81 1437 127
rect 1483 81 1512 127
rect 1408 68 1512 81
rect 1632 219 1736 232
rect 1632 173 1661 219
rect 1707 173 1736 219
rect 1632 68 1736 173
rect 1856 127 1960 232
rect 1856 81 1885 127
rect 1931 81 1960 127
rect 1856 68 1960 81
rect 2080 219 2184 232
rect 2080 173 2109 219
rect 2155 173 2184 219
rect 2080 68 2184 173
rect 2304 127 2392 232
rect 2304 81 2333 127
rect 2379 81 2392 127
rect 2304 68 2392 81
rect 991 49 1004 68
rect 932 36 1004 49
<< mvpdiff >>
rect 84 602 172 716
rect 84 556 97 602
rect 143 556 172 602
rect 84 527 172 556
rect 272 698 376 716
rect 272 652 301 698
rect 347 652 376 698
rect 272 527 376 652
rect 476 678 660 716
rect 476 632 585 678
rect 631 632 660 678
rect 476 527 660 632
rect 760 586 848 716
rect 760 540 789 586
rect 835 540 848 586
rect 760 527 848 540
rect 1056 703 1144 716
rect 1056 657 1069 703
rect 1115 657 1144 703
rect 1056 481 1144 657
rect 1244 665 1348 716
rect 1244 525 1273 665
rect 1319 525 1348 665
rect 1244 481 1348 525
rect 1448 703 1552 716
rect 1448 657 1477 703
rect 1523 657 1552 703
rect 1448 481 1552 657
rect 1652 665 1756 716
rect 1652 525 1681 665
rect 1727 525 1756 665
rect 1652 481 1756 525
rect 1856 703 1960 716
rect 1856 657 1885 703
rect 1931 657 1960 703
rect 1856 481 1960 657
rect 2060 665 2164 716
rect 2060 525 2089 665
rect 2135 525 2164 665
rect 2060 481 2164 525
rect 2264 703 2352 716
rect 2264 657 2293 703
rect 2339 657 2352 703
rect 2264 481 2352 657
<< mvndiffc >>
rect 49 173 95 219
rect 273 82 319 128
rect 497 123 543 169
rect 765 228 811 274
rect 945 49 991 95
rect 1213 173 1259 219
rect 1437 81 1483 127
rect 1661 173 1707 219
rect 1885 81 1931 127
rect 2109 173 2155 219
rect 2333 81 2379 127
<< mvpdiffc >>
rect 97 556 143 602
rect 301 652 347 698
rect 585 632 631 678
rect 789 540 835 586
rect 1069 657 1115 703
rect 1273 525 1319 665
rect 1477 657 1523 703
rect 1681 525 1727 665
rect 1885 657 1931 703
rect 2089 525 2135 665
rect 2293 657 2339 703
<< polysilicon >>
rect 172 716 272 760
rect 376 716 476 760
rect 660 716 760 760
rect 1144 716 1244 760
rect 1348 716 1448 760
rect 1552 716 1652 760
rect 1756 716 1856 760
rect 1960 716 2060 760
rect 2164 716 2264 760
rect 172 413 272 527
rect 376 413 476 527
rect 660 493 760 527
rect 660 447 673 493
rect 719 447 760 493
rect 660 434 760 447
rect 1144 420 1244 481
rect 1348 420 1448 481
rect 124 412 612 413
rect 124 366 185 412
rect 231 373 612 412
rect 231 366 244 373
rect 124 232 244 366
rect 348 311 468 324
rect 348 265 385 311
rect 431 265 468 311
rect 348 232 468 265
rect 572 288 612 373
rect 1064 407 1448 420
rect 1064 361 1119 407
rect 1353 387 1448 407
rect 1552 439 1652 481
rect 1552 393 1593 439
rect 1639 420 1652 439
rect 1756 439 1856 481
rect 1756 420 1769 439
rect 1639 393 1769 420
rect 1815 420 1856 439
rect 1960 439 2060 481
rect 1960 420 1973 439
rect 1815 393 1973 420
rect 2019 420 2060 439
rect 2164 420 2264 481
rect 2019 393 2264 420
rect 1353 361 1408 387
rect 1552 380 2264 393
rect 1064 348 1408 361
rect 572 232 692 288
rect 1064 232 1184 348
rect 1288 232 1408 348
rect 1512 319 2304 332
rect 1512 273 1547 319
rect 1593 292 1749 319
rect 1593 273 1632 292
rect 1512 232 1632 273
rect 1736 273 1749 292
rect 1795 292 1973 319
rect 1795 273 1856 292
rect 1736 232 1856 273
rect 1960 273 1973 292
rect 2019 292 2304 319
rect 2019 273 2080 292
rect 1960 232 2080 273
rect 2184 232 2304 292
rect 124 24 244 68
rect 348 24 468 68
rect 572 24 692 68
rect 1064 24 1184 68
rect 1288 24 1408 68
rect 1512 24 1632 68
rect 1736 24 1856 68
rect 1960 24 2080 68
rect 2184 24 2304 68
<< polycontact >>
rect 673 447 719 493
rect 185 366 231 412
rect 385 265 431 311
rect 1119 361 1353 407
rect 1593 393 1639 439
rect 1769 393 1815 439
rect 1973 393 2019 439
rect 1547 273 1593 319
rect 1749 273 1795 319
rect 1973 273 2019 319
<< metal1 >>
rect 0 724 2464 844
rect 290 698 358 724
rect 290 652 301 698
rect 347 652 358 698
rect 1058 703 1126 724
rect 574 632 585 678
rect 631 632 965 678
rect 1058 657 1069 703
rect 1115 657 1126 703
rect 1466 703 1534 724
rect 1262 665 1330 676
rect 84 556 97 602
rect 143 556 431 602
rect 385 504 431 556
rect 778 540 789 586
rect 835 540 846 586
rect 385 493 730 504
rect 385 447 673 493
rect 719 447 730 493
rect 130 412 318 430
rect 130 366 185 412
rect 231 366 318 412
rect 130 354 318 366
rect 385 311 431 447
rect 778 401 846 540
rect 38 219 431 265
rect 497 355 846 401
rect 919 552 965 632
rect 1262 552 1273 665
rect 919 525 1273 552
rect 1319 552 1330 665
rect 1466 657 1477 703
rect 1523 657 1534 703
rect 1874 703 1942 724
rect 1670 665 1738 676
rect 1319 525 1549 552
rect 919 506 1549 525
rect 38 173 49 219
rect 95 173 106 219
rect 38 170 106 173
rect 497 169 543 355
rect 919 309 965 506
rect 1503 439 1549 506
rect 1670 525 1681 665
rect 1727 560 1738 665
rect 1874 657 1885 703
rect 1931 657 1942 703
rect 2282 703 2350 724
rect 2078 665 2146 676
rect 2078 560 2089 665
rect 1727 525 2089 560
rect 2135 552 2146 665
rect 2282 657 2293 703
rect 2339 657 2350 703
rect 2135 525 2222 552
rect 1670 504 2222 525
rect 1026 407 1438 430
rect 1026 361 1119 407
rect 1353 361 1438 407
rect 1503 393 1593 439
rect 1639 393 1769 439
rect 1815 393 1973 439
rect 2019 393 2030 439
rect 1026 354 1438 361
rect 754 274 965 309
rect 754 228 765 274
rect 811 263 965 274
rect 1503 273 1547 319
rect 1593 273 1749 319
rect 1795 273 1973 319
rect 2019 273 2030 319
rect 811 228 822 263
rect 1503 219 1549 273
rect 2146 227 2222 504
rect 1139 187 1213 219
rect 262 128 330 131
rect 262 82 273 128
rect 319 82 330 128
rect 843 173 1213 187
rect 1259 173 1549 219
rect 1632 219 2222 227
rect 1632 173 1661 219
rect 1707 173 2109 219
rect 2155 173 2222 219
rect 843 152 1189 173
rect 543 141 1189 152
rect 543 123 888 141
rect 497 106 888 123
rect 262 60 330 82
rect 934 60 945 95
rect 0 49 945 60
rect 991 60 1002 95
rect 1426 81 1437 127
rect 1483 81 1494 127
rect 1426 60 1494 81
rect 1874 81 1885 127
rect 1931 81 1942 127
rect 1874 60 1942 81
rect 2322 81 2333 127
rect 2379 81 2390 127
rect 2322 60 2390 81
rect 991 49 2464 60
rect 0 -60 2464 49
<< labels >>
flabel metal1 s 2078 560 2146 676 0 FreeSans 400 0 0 0 Z
port 3 nsew default output
flabel metal1 s 130 354 318 430 0 FreeSans 600 0 0 0 EN
port 1 nsew default input
flabel metal1 s 1026 354 1438 430 0 FreeSans 400 0 0 0 I
port 2 nsew default input
flabel metal1 s 262 127 330 131 0 FreeSans 400 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel metal1 s 0 724 2464 844 0 FreeSans 400 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 5 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 6 nsew ground bidirectional
rlabel metal1 s 1670 560 1738 676 1 Z
port 3 nsew default output
rlabel metal1 s 1670 552 2146 560 1 Z
port 3 nsew default output
rlabel metal1 s 1670 504 2222 552 1 Z
port 3 nsew default output
rlabel metal1 s 2146 227 2222 504 1 Z
port 3 nsew default output
rlabel metal1 s 1632 173 2222 227 1 Z
port 3 nsew default output
rlabel metal1 s 2282 657 2350 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1874 657 1942 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1466 657 1534 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1058 657 1126 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 290 657 358 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 290 652 358 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2322 95 2390 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1874 95 1942 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1426 95 1494 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 95 330 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2322 60 2390 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1874 60 1942 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1426 60 1494 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 934 60 1002 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 60 330 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 2464 60 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2464 784
string GDS_END 1408856
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1402790
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
