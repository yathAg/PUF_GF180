magic
tech gf180mcuC
timestamp 1698431365
<< properties >>
string GDS_END 912700
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 856034
<< end >>
