magic
tech gf180mcuD
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 453 3222 1094
<< pwell >>
rect -86 -86 3222 453
<< mvnmos >>
rect 125 134 245 292
rect 385 134 505 274
rect 753 69 873 209
rect 921 69 1041 209
rect 1145 69 1265 209
rect 1405 69 1525 227
rect 1629 69 1749 227
rect 1853 69 1973 227
rect 2113 69 2233 333
rect 2337 69 2457 333
rect 2561 69 2681 333
rect 2785 69 2905 333
<< mvpmos >>
rect 145 615 245 891
rect 385 615 485 815
rect 833 649 933 849
rect 981 649 1081 849
rect 1185 649 1285 849
rect 1425 573 1525 849
rect 1629 573 1729 849
rect 1833 573 1933 849
rect 2073 573 2173 939
rect 2277 573 2377 939
rect 2481 573 2581 939
rect 2685 573 2785 939
<< mvndiff >>
rect 37 193 125 292
rect 37 147 50 193
rect 96 147 125 193
rect 37 134 125 147
rect 245 274 325 292
rect 245 193 385 274
rect 245 147 274 193
rect 320 147 385 193
rect 245 134 385 147
rect 505 193 593 274
rect 2033 227 2113 333
rect 1325 209 1405 227
rect 505 147 534 193
rect 580 147 593 193
rect 505 134 593 147
rect 665 193 753 209
rect 665 147 678 193
rect 724 147 753 193
rect 665 69 753 147
rect 873 69 921 209
rect 1041 193 1145 209
rect 1041 147 1070 193
rect 1116 147 1145 193
rect 1041 69 1145 147
rect 1265 69 1405 209
rect 1525 193 1629 227
rect 1525 147 1554 193
rect 1600 147 1629 193
rect 1525 69 1629 147
rect 1749 193 1853 227
rect 1749 147 1778 193
rect 1824 147 1853 193
rect 1749 69 1853 147
rect 1973 193 2113 227
rect 1973 147 2002 193
rect 2048 147 2113 193
rect 1973 69 2113 147
rect 2233 287 2337 333
rect 2233 147 2262 287
rect 2308 147 2337 287
rect 2233 69 2337 147
rect 2457 185 2561 333
rect 2457 139 2486 185
rect 2532 139 2561 185
rect 2457 69 2561 139
rect 2681 287 2785 333
rect 2681 147 2710 287
rect 2756 147 2785 287
rect 2681 69 2785 147
rect 2905 287 2993 333
rect 2905 147 2934 287
rect 2980 147 2993 287
rect 2905 69 2993 147
<< mvpdiff >>
rect 57 802 145 891
rect 57 662 70 802
rect 116 662 145 802
rect 57 615 145 662
rect 245 815 325 891
rect 1993 849 2073 939
rect 245 802 385 815
rect 245 662 274 802
rect 320 662 385 802
rect 245 615 385 662
rect 485 802 573 815
rect 485 662 514 802
rect 560 662 573 802
rect 485 615 573 662
rect 745 802 833 849
rect 745 662 758 802
rect 804 662 833 802
rect 745 649 833 662
rect 933 649 981 849
rect 1081 802 1185 849
rect 1081 662 1110 802
rect 1156 662 1185 802
rect 1081 649 1185 662
rect 1285 649 1425 849
rect 1345 573 1425 649
rect 1525 802 1629 849
rect 1525 662 1554 802
rect 1600 662 1629 802
rect 1525 573 1629 662
rect 1729 802 1833 849
rect 1729 662 1758 802
rect 1804 662 1833 802
rect 1729 573 1833 662
rect 1933 802 2073 849
rect 1933 662 1962 802
rect 2008 662 2073 802
rect 1933 573 2073 662
rect 2173 802 2277 939
rect 2173 662 2202 802
rect 2248 662 2277 802
rect 2173 573 2277 662
rect 2377 802 2481 939
rect 2377 662 2406 802
rect 2452 662 2481 802
rect 2377 573 2481 662
rect 2581 802 2685 939
rect 2581 662 2610 802
rect 2656 662 2685 802
rect 2581 573 2685 662
rect 2785 802 2873 939
rect 2785 662 2814 802
rect 2860 662 2873 802
rect 2785 573 2873 662
<< mvndiffc >>
rect 50 147 96 193
rect 274 147 320 193
rect 534 147 580 193
rect 678 147 724 193
rect 1070 147 1116 193
rect 1554 147 1600 193
rect 1778 147 1824 193
rect 2002 147 2048 193
rect 2262 147 2308 287
rect 2486 139 2532 185
rect 2710 147 2756 287
rect 2934 147 2980 287
<< mvpdiffc >>
rect 70 662 116 802
rect 274 662 320 802
rect 514 662 560 802
rect 758 662 804 802
rect 1110 662 1156 802
rect 1554 662 1600 802
rect 1758 662 1804 802
rect 1962 662 2008 802
rect 2202 662 2248 802
rect 2406 662 2452 802
rect 2610 662 2656 802
rect 2814 662 2860 802
<< polysilicon >>
rect 385 941 1081 981
rect 145 891 245 935
rect 385 815 485 941
rect 833 849 933 893
rect 981 849 1081 941
rect 2073 939 2173 983
rect 2277 939 2377 983
rect 2481 939 2581 983
rect 2685 939 2785 983
rect 1185 849 1285 893
rect 1425 849 1525 893
rect 1629 849 1729 893
rect 1833 849 1933 893
rect 145 419 245 615
rect 145 373 158 419
rect 204 373 245 419
rect 145 336 245 373
rect 125 292 245 336
rect 385 419 485 615
rect 833 605 933 649
rect 981 605 1081 649
rect 833 432 873 605
rect 385 373 398 419
rect 444 373 485 419
rect 385 318 485 373
rect 753 419 873 432
rect 753 373 814 419
rect 860 373 873 419
rect 385 274 505 318
rect 753 209 873 373
rect 921 419 993 432
rect 921 373 934 419
rect 980 373 993 419
rect 1041 426 1081 605
rect 1185 605 1285 649
rect 1185 546 1284 605
rect 1153 533 1284 546
rect 1153 487 1166 533
rect 1212 487 1284 533
rect 1153 474 1284 487
rect 1041 386 1265 426
rect 921 253 993 373
rect 921 209 1041 253
rect 1145 209 1265 386
rect 1425 419 1525 573
rect 1425 373 1466 419
rect 1512 373 1525 419
rect 1425 271 1525 373
rect 1405 227 1525 271
rect 1629 513 1729 573
rect 1833 513 1933 573
rect 2073 513 2173 573
rect 2277 513 2377 573
rect 2481 513 2581 573
rect 2685 513 2785 573
rect 1629 441 2905 513
rect 1629 419 1749 441
rect 1629 373 1642 419
rect 1688 373 1749 419
rect 1629 227 1749 373
rect 1853 227 1973 441
rect 2113 333 2233 441
rect 2337 333 2457 441
rect 2561 333 2681 441
rect 2785 333 2905 441
rect 125 90 245 134
rect 385 90 505 134
rect 753 25 873 69
rect 921 25 1041 69
rect 1145 25 1265 69
rect 1405 25 1525 69
rect 1629 25 1749 69
rect 1853 25 1973 69
rect 2113 25 2233 69
rect 2337 25 2457 69
rect 2561 25 2681 69
rect 2785 25 2905 69
<< polycontact >>
rect 158 373 204 419
rect 398 373 444 419
rect 814 373 860 419
rect 934 373 980 419
rect 1166 487 1212 533
rect 1466 373 1512 419
rect 1642 373 1688 419
<< metal1 >>
rect 0 918 3136 1098
rect 50 802 116 813
rect 50 662 70 802
rect 50 651 116 662
rect 274 802 320 918
rect 274 651 320 662
rect 514 802 560 813
rect 50 308 96 651
rect 514 544 560 662
rect 758 802 804 918
rect 758 651 804 662
rect 1110 802 1156 813
rect 1110 636 1156 662
rect 1554 802 1600 918
rect 1554 651 1600 662
rect 1758 802 1824 813
rect 1804 662 1824 802
rect 1110 590 1304 636
rect 142 419 204 542
rect 514 533 1212 544
rect 514 487 1166 533
rect 514 476 1212 487
rect 142 373 158 419
rect 142 354 204 373
rect 398 419 444 430
rect 398 308 444 373
rect 50 262 444 308
rect 50 193 96 262
rect 50 136 96 147
rect 274 193 320 204
rect 274 90 320 147
rect 514 193 580 476
rect 814 419 866 430
rect 860 373 866 419
rect 814 242 866 373
rect 934 419 980 476
rect 934 362 980 373
rect 1258 204 1304 590
rect 1758 522 1824 662
rect 1962 802 2008 918
rect 1962 651 2008 662
rect 2202 802 2248 813
rect 1466 476 1824 522
rect 1466 419 1512 476
rect 1466 362 1512 373
rect 1642 419 1688 430
rect 1642 296 1688 373
rect 514 147 534 193
rect 514 136 580 147
rect 678 193 724 204
rect 678 90 724 147
rect 1070 193 1304 204
rect 1116 182 1304 193
rect 1462 250 1688 296
rect 1462 182 1508 250
rect 1116 147 1508 182
rect 1070 136 1508 147
rect 1554 193 1600 204
rect 1554 90 1600 147
rect 1778 193 1824 476
rect 2202 430 2248 662
rect 2406 802 2452 918
rect 2406 651 2452 662
rect 2610 802 2656 813
rect 2202 384 2322 430
rect 2262 288 2322 384
rect 2610 298 2656 662
rect 2814 802 2860 918
rect 2814 651 2860 662
rect 2610 288 2756 298
rect 2262 287 2756 288
rect 1778 136 1824 147
rect 2002 193 2048 204
rect 2002 90 2048 147
rect 2308 242 2710 287
rect 2262 136 2308 147
rect 2486 185 2532 196
rect 2486 90 2532 139
rect 2710 136 2756 147
rect 2934 287 2980 298
rect 2934 90 2980 147
rect 0 -90 3136 90
<< labels >>
flabel metal1 s 814 242 866 430 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 142 354 204 542 0 FreeSans 200 0 0 0 E
port 2 nsew clock input
flabel metal1 s 2610 430 2656 813 0 FreeSans 200 0 0 0 Q
port 3 nsew default output
flabel metal1 s 0 918 3136 1098 0 FreeSans 200 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 2934 204 2980 298 0 FreeSans 200 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 5 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 6 nsew ground bidirectional
rlabel metal1 s 2202 430 2248 813 1 Q
port 3 nsew default output
rlabel metal1 s 2610 384 2656 430 1 Q
port 3 nsew default output
rlabel metal1 s 2202 384 2322 430 1 Q
port 3 nsew default output
rlabel metal1 s 2610 298 2656 384 1 Q
port 3 nsew default output
rlabel metal1 s 2262 298 2322 384 1 Q
port 3 nsew default output
rlabel metal1 s 2610 288 2756 298 1 Q
port 3 nsew default output
rlabel metal1 s 2262 288 2322 298 1 Q
port 3 nsew default output
rlabel metal1 s 2262 242 2756 288 1 Q
port 3 nsew default output
rlabel metal1 s 2710 136 2756 242 1 Q
port 3 nsew default output
rlabel metal1 s 2262 136 2308 242 1 Q
port 3 nsew default output
rlabel metal1 s 2814 651 2860 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2406 651 2452 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1962 651 2008 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1554 651 1600 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 758 651 804 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 274 651 320 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2934 196 2980 204 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2002 196 2048 204 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1554 196 1600 204 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 678 196 724 204 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 274 196 320 204 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2934 90 2980 196 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2486 90 2532 196 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2002 90 2048 196 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1554 90 1600 196 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 678 90 724 196 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 274 90 320 196 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 3136 90 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3136 1008
string GDS_END 1001938
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 995070
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
