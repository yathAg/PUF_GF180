magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 377 5126 870
rect -86 352 1121 377
rect 4085 352 5126 377
<< pwell >>
rect 1121 352 4085 377
rect -86 -86 5126 352
<< mvnmos >>
rect 124 156 244 228
rect 348 156 468 228
rect 516 156 636 228
rect 740 156 860 228
rect 908 156 1028 228
rect 1185 135 1305 228
rect 1648 139 1768 232
rect 2060 124 2180 196
rect 2284 124 2404 196
rect 2452 124 2572 196
rect 2692 124 2812 196
rect 3004 185 3124 257
rect 3228 185 3348 257
rect 3452 185 3572 257
rect 3690 185 3810 257
rect 4002 124 4122 232
rect 4186 124 4306 232
rect 4554 70 4674 232
rect 4778 70 4898 232
<< mvpmos >>
rect 124 502 224 628
rect 348 502 448 628
rect 496 502 596 628
rect 740 502 840 628
rect 888 502 988 628
rect 1185 502 1285 687
rect 1648 497 1748 660
rect 2054 502 2154 628
rect 2258 502 2358 628
rect 2462 502 2562 628
rect 2754 502 2854 628
rect 3102 502 3202 628
rect 3306 502 3406 628
rect 3539 502 3639 628
rect 3743 502 3843 628
rect 4002 502 4102 686
rect 4206 502 4306 686
rect 4564 472 4664 715
rect 4778 472 4878 715
<< mvndiff >>
rect 1365 244 1437 257
rect 1365 228 1378 244
rect 36 215 124 228
rect 36 169 49 215
rect 95 169 124 215
rect 36 156 124 169
rect 244 215 348 228
rect 244 169 273 215
rect 319 169 348 215
rect 244 156 348 169
rect 468 156 516 228
rect 636 215 740 228
rect 636 169 665 215
rect 711 169 740 215
rect 636 156 740 169
rect 860 156 908 228
rect 1028 194 1185 228
rect 1028 156 1110 194
rect 1097 148 1110 156
rect 1156 148 1185 194
rect 1097 135 1185 148
rect 1305 198 1378 228
rect 1424 198 1437 244
rect 1828 244 1900 257
rect 1828 232 1841 244
rect 1305 135 1437 198
rect 1560 198 1648 232
rect 1560 152 1573 198
rect 1619 152 1648 198
rect 1560 139 1648 152
rect 1768 198 1841 232
rect 1887 198 1900 244
rect 1768 139 1900 198
rect 2872 196 3004 257
rect 1972 183 2060 196
rect 1972 137 1985 183
rect 2031 137 2060 183
rect 1972 124 2060 137
rect 2180 183 2284 196
rect 2180 137 2209 183
rect 2255 137 2284 183
rect 2180 124 2284 137
rect 2404 124 2452 196
rect 2572 124 2692 196
rect 2812 185 3004 196
rect 3124 244 3228 257
rect 3124 198 3153 244
rect 3199 198 3228 244
rect 3124 185 3228 198
rect 3348 244 3452 257
rect 3348 198 3377 244
rect 3423 198 3452 244
rect 3348 185 3452 198
rect 3572 244 3690 257
rect 3572 198 3615 244
rect 3661 198 3690 244
rect 3572 185 3690 198
rect 3810 232 3942 257
rect 3810 185 4002 232
rect 2812 183 2944 185
rect 2812 137 2885 183
rect 2931 137 2944 183
rect 3870 183 4002 185
rect 2812 124 2944 137
rect 3870 137 3883 183
rect 3929 137 4002 183
rect 3870 124 4002 137
rect 4122 124 4186 232
rect 4306 219 4394 232
rect 4306 173 4335 219
rect 4381 173 4394 219
rect 4306 124 4394 173
rect 4466 168 4554 232
rect 4466 122 4479 168
rect 4525 122 4554 168
rect 4466 70 4554 122
rect 4674 202 4778 232
rect 4674 156 4703 202
rect 4749 156 4778 202
rect 4674 70 4778 156
rect 4898 168 4986 232
rect 4898 122 4927 168
rect 4973 122 4986 168
rect 4898 70 4986 122
<< mvpdiff >>
rect 1516 716 1588 729
rect 1048 634 1185 687
rect 1048 628 1075 634
rect 36 585 124 628
rect 36 539 49 585
rect 95 539 124 585
rect 36 502 124 539
rect 224 615 348 628
rect 224 569 263 615
rect 309 569 348 615
rect 224 502 348 569
rect 448 502 496 628
rect 596 595 740 628
rect 596 549 665 595
rect 711 549 740 595
rect 596 502 740 549
rect 840 502 888 628
rect 988 588 1075 628
rect 1121 588 1185 634
rect 988 502 1185 588
rect 1285 561 1393 687
rect 1285 515 1322 561
rect 1368 515 1393 561
rect 1285 502 1393 515
rect 1516 670 1529 716
rect 1575 670 1588 716
rect 1516 660 1588 670
rect 1516 497 1648 660
rect 1748 558 1836 660
rect 2622 647 2694 660
rect 2622 628 2635 647
rect 1748 512 1777 558
rect 1823 512 1836 558
rect 1748 497 1836 512
rect 1966 589 2054 628
rect 1966 543 1979 589
rect 2025 543 2054 589
rect 1966 502 2054 543
rect 2154 585 2258 628
rect 2154 539 2183 585
rect 2229 539 2258 585
rect 2154 502 2258 539
rect 2358 584 2462 628
rect 2358 538 2387 584
rect 2433 538 2462 584
rect 2358 502 2462 538
rect 2562 601 2635 628
rect 2681 628 2694 647
rect 3903 628 4002 686
rect 2681 601 2754 628
rect 2562 502 2754 601
rect 2854 584 2942 628
rect 2854 538 2883 584
rect 2929 538 2942 584
rect 2854 502 2942 538
rect 3014 590 3102 628
rect 3014 544 3027 590
rect 3073 544 3102 590
rect 3014 502 3102 544
rect 3202 582 3306 628
rect 3202 536 3231 582
rect 3277 536 3306 582
rect 3202 502 3306 536
rect 3406 595 3539 628
rect 3406 549 3435 595
rect 3481 549 3539 595
rect 3406 502 3539 549
rect 3639 561 3743 628
rect 3639 515 3668 561
rect 3714 515 3743 561
rect 3639 502 3743 515
rect 3843 615 4002 628
rect 3843 569 3907 615
rect 3953 569 4002 615
rect 3843 502 4002 569
rect 4102 561 4206 686
rect 4102 515 4131 561
rect 4177 515 4206 561
rect 4102 502 4206 515
rect 4306 669 4394 686
rect 4306 529 4335 669
rect 4381 529 4394 669
rect 4306 502 4394 529
rect 4476 680 4564 715
rect 4476 634 4489 680
rect 4535 634 4564 680
rect 4476 575 4564 634
rect 4476 529 4489 575
rect 4535 529 4564 575
rect 4476 472 4564 529
rect 4664 660 4778 715
rect 4664 614 4703 660
rect 4749 614 4778 660
rect 4664 546 4778 614
rect 4664 500 4703 546
rect 4749 500 4778 546
rect 4664 472 4778 500
rect 4878 680 4966 715
rect 4878 634 4907 680
rect 4953 634 4966 680
rect 4878 575 4966 634
rect 4878 529 4907 575
rect 4953 529 4966 575
rect 4878 472 4966 529
<< mvndiffc >>
rect 49 169 95 215
rect 273 169 319 215
rect 665 169 711 215
rect 1110 148 1156 194
rect 1378 198 1424 244
rect 1573 152 1619 198
rect 1841 198 1887 244
rect 1985 137 2031 183
rect 2209 137 2255 183
rect 3153 198 3199 244
rect 3377 198 3423 244
rect 3615 198 3661 244
rect 2885 137 2931 183
rect 3883 137 3929 183
rect 4335 173 4381 219
rect 4479 122 4525 168
rect 4703 156 4749 202
rect 4927 122 4973 168
<< mvpdiffc >>
rect 49 539 95 585
rect 263 569 309 615
rect 665 549 711 595
rect 1075 588 1121 634
rect 1322 515 1368 561
rect 1529 670 1575 716
rect 1777 512 1823 558
rect 1979 543 2025 589
rect 2183 539 2229 585
rect 2387 538 2433 584
rect 2635 601 2681 647
rect 2883 538 2929 584
rect 3027 544 3073 590
rect 3231 536 3277 582
rect 3435 549 3481 595
rect 3668 515 3714 561
rect 3907 569 3953 615
rect 4131 515 4177 561
rect 4335 529 4381 669
rect 4489 634 4535 680
rect 4489 529 4535 575
rect 4703 614 4749 660
rect 4703 500 4749 546
rect 4907 634 4953 680
rect 4907 529 4953 575
<< polysilicon >>
rect 124 720 988 760
rect 124 628 224 720
rect 348 628 448 672
rect 496 628 596 672
rect 740 628 840 672
rect 888 628 988 720
rect 1185 687 1285 731
rect 1648 720 3406 760
rect 1648 660 1748 720
rect 124 432 224 502
rect 124 351 244 432
rect 124 305 150 351
rect 196 305 244 351
rect 124 228 244 305
rect 348 351 448 502
rect 496 469 596 502
rect 496 423 525 469
rect 571 423 596 469
rect 496 410 596 423
rect 348 305 374 351
rect 420 305 448 351
rect 348 272 448 305
rect 740 407 840 502
rect 888 458 988 502
rect 740 361 753 407
rect 799 361 840 407
rect 1185 415 1285 502
rect 2054 628 2154 672
rect 2258 628 2358 720
rect 2462 628 2562 672
rect 2754 628 2854 672
rect 3102 628 3202 672
rect 3306 628 3406 720
rect 4002 686 4102 731
rect 4206 686 4306 731
rect 4564 715 4664 759
rect 4778 715 4878 759
rect 3539 628 3639 673
rect 3743 628 3843 673
rect 1185 369 1213 415
rect 1259 413 1285 415
rect 1648 448 1748 497
rect 1259 369 1305 413
rect 740 272 840 361
rect 908 335 1028 361
rect 908 289 926 335
rect 972 289 1028 335
rect 348 228 468 272
rect 516 228 636 272
rect 740 228 860 272
rect 908 228 1028 289
rect 1185 228 1305 369
rect 1648 402 1661 448
rect 1707 402 1748 448
rect 1648 277 1748 402
rect 2054 407 2154 502
rect 2258 458 2358 502
rect 2462 460 2562 502
rect 2054 361 2067 407
rect 2113 372 2154 407
rect 2462 414 2503 460
rect 2549 414 2562 460
rect 2754 427 2854 502
rect 3102 442 3202 502
rect 2462 406 2562 414
rect 2113 361 2404 372
rect 2054 326 2404 361
rect 2284 325 2404 326
rect 2284 279 2301 325
rect 2347 279 2404 325
rect 124 64 244 156
rect 348 112 468 156
rect 516 64 636 156
rect 740 112 860 156
rect 908 112 1028 156
rect 1648 232 1768 277
rect 2060 196 2180 240
rect 2284 196 2404 279
rect 2462 240 2572 406
rect 2452 196 2572 240
rect 2692 346 2854 427
rect 3004 402 3202 442
rect 3306 442 3406 502
rect 3539 469 3639 502
rect 3306 402 3469 442
rect 3539 423 3552 469
rect 3598 423 3639 469
rect 3743 442 3843 502
rect 3539 410 3639 423
rect 3004 368 3124 402
rect 2692 196 2812 346
rect 3004 322 3017 368
rect 3063 322 3124 368
rect 3429 372 3469 402
rect 3710 407 3843 442
rect 3004 257 3124 322
rect 3228 336 3348 349
rect 3228 290 3274 336
rect 3320 290 3348 336
rect 3429 332 3492 372
rect 3228 257 3348 290
rect 3452 301 3492 332
rect 3710 361 3736 407
rect 3782 361 3843 407
rect 3710 317 3843 361
rect 3710 301 3810 317
rect 3452 257 3572 301
rect 3690 257 3810 301
rect 4002 311 4102 502
rect 4002 265 4023 311
rect 4069 276 4102 311
rect 4206 469 4306 502
rect 4206 423 4223 469
rect 4269 423 4306 469
rect 4206 276 4306 423
rect 4564 439 4664 472
rect 4564 299 4583 439
rect 4629 388 4664 439
rect 4778 388 4878 472
rect 4629 320 4878 388
rect 4629 299 4674 320
rect 4564 277 4674 299
rect 4069 265 4122 276
rect 1185 91 1305 135
rect 124 24 636 64
rect 1648 64 1768 139
rect 4002 232 4122 265
rect 4186 232 4306 276
rect 4554 232 4674 277
rect 4778 277 4878 320
rect 4778 232 4898 277
rect 3004 141 3124 185
rect 3228 141 3348 185
rect 3452 141 3572 185
rect 3690 141 3810 185
rect 2060 64 2180 124
rect 2284 80 2404 124
rect 2452 80 2572 124
rect 1648 24 2180 64
rect 2692 64 2812 124
rect 4002 64 4122 124
rect 4186 80 4306 124
rect 2692 24 4122 64
rect 4554 26 4674 70
rect 4778 26 4898 70
<< polycontact >>
rect 150 305 196 351
rect 525 423 571 469
rect 374 305 420 351
rect 753 361 799 407
rect 1213 369 1259 415
rect 926 289 972 335
rect 1661 402 1707 448
rect 2067 361 2113 407
rect 2503 414 2549 460
rect 2301 279 2347 325
rect 3552 423 3598 469
rect 3017 322 3063 368
rect 3274 290 3320 336
rect 3736 361 3782 407
rect 4023 265 4069 311
rect 4223 423 4269 469
rect 4583 299 4629 439
<< metal1 >>
rect 0 724 5040 844
rect 252 615 320 724
rect 49 585 95 608
rect 252 569 263 615
rect 309 569 320 615
rect 1075 634 1121 724
rect 1518 716 1586 724
rect 654 549 665 595
rect 711 549 1015 595
rect 1075 577 1121 588
rect 1217 632 1472 678
rect 1518 670 1529 716
rect 1575 670 1586 716
rect 49 523 95 539
rect 969 531 1015 549
rect 1217 531 1263 632
rect 1426 624 1472 632
rect 1641 632 2025 678
rect 1641 624 1687 632
rect 1426 578 1687 624
rect 1979 589 2025 632
rect 2624 647 2692 724
rect 49 477 571 523
rect 969 484 1263 531
rect 1322 561 1368 578
rect 1777 558 1823 569
rect 1368 515 1707 524
rect 1322 477 1707 515
rect 49 215 95 477
rect 525 469 571 477
rect 49 156 95 169
rect 141 351 206 430
rect 141 305 150 351
rect 196 305 206 351
rect 141 119 206 305
rect 365 351 430 430
rect 365 305 374 351
rect 420 305 430 351
rect 273 215 319 228
rect 273 60 319 169
rect 365 119 430 305
rect 525 307 571 423
rect 619 407 878 438
rect 619 361 753 407
rect 799 361 878 407
rect 619 353 878 361
rect 1026 415 1326 431
rect 1026 369 1213 415
rect 1259 369 1326 415
rect 1026 353 1326 369
rect 926 335 972 350
rect 525 289 926 307
rect 525 261 972 289
rect 1018 252 1321 298
rect 1389 255 1435 477
rect 1661 448 1707 477
rect 1661 382 1707 402
rect 1979 529 2025 543
rect 2183 585 2229 625
rect 2624 601 2635 647
rect 2681 601 2692 647
rect 1777 407 1823 512
rect 2183 459 2229 539
rect 2387 584 2433 601
rect 2624 600 2692 601
rect 2883 584 2929 601
rect 2433 538 2883 552
rect 2387 506 2929 538
rect 3027 590 3073 724
rect 3431 632 3815 678
rect 3027 533 3073 544
rect 3231 582 3277 607
rect 3231 460 3277 536
rect 2183 413 2439 459
rect 2492 414 2503 460
rect 2549 414 3277 460
rect 3431 595 3492 632
rect 3431 549 3435 595
rect 3481 549 3492 595
rect 3431 538 3492 549
rect 3644 561 3714 586
rect 1777 361 2067 407
rect 2113 361 2124 407
rect 1777 360 2124 361
rect 1018 215 1064 252
rect 650 169 665 215
rect 711 169 1064 215
rect 1110 194 1156 205
rect 1110 60 1156 148
rect 1275 152 1321 252
rect 1367 244 1435 255
rect 1367 198 1378 244
rect 1424 198 1435 244
rect 1481 259 1736 306
rect 1481 152 1527 259
rect 1275 106 1527 152
rect 1573 198 1619 209
rect 1573 60 1619 152
rect 1690 152 1736 259
rect 1830 244 1898 360
rect 1830 198 1841 244
rect 1887 198 1898 244
rect 1985 183 2031 194
rect 1690 137 1985 152
rect 1690 106 2031 137
rect 2209 183 2255 413
rect 2393 368 2439 413
rect 2301 325 2347 344
rect 2393 322 3017 368
rect 3063 322 3074 368
rect 2301 275 2347 279
rect 2301 229 3042 275
rect 2209 126 2255 137
rect 2874 137 2885 183
rect 2931 137 2942 183
rect 2874 60 2942 137
rect 2996 152 3042 229
rect 3142 244 3210 414
rect 3142 198 3153 244
rect 3199 198 3210 244
rect 3274 336 3320 347
rect 3274 152 3320 290
rect 3431 244 3477 538
rect 3644 515 3668 561
rect 3644 484 3714 515
rect 3769 523 3815 632
rect 3896 615 3964 724
rect 3896 569 3907 615
rect 3953 569 3964 615
rect 4039 631 4269 678
rect 4039 523 4085 631
rect 3366 198 3377 244
rect 3423 198 3477 244
rect 3523 469 3598 480
rect 3523 423 3552 469
rect 3523 412 3598 423
rect 3523 152 3569 412
rect 3644 349 3690 484
rect 3769 477 4085 523
rect 4131 561 4177 572
rect 4131 431 4177 515
rect 3615 302 3690 349
rect 3736 407 4177 431
rect 3782 385 4177 407
rect 4223 469 4269 631
rect 4335 669 4381 724
rect 4335 514 4381 529
rect 4489 680 4535 724
rect 4907 680 4953 724
rect 4489 575 4535 634
rect 4489 512 4535 529
rect 4692 660 4796 672
rect 4692 614 4703 660
rect 4749 614 4796 660
rect 4692 546 4796 614
rect 4692 500 4703 546
rect 4749 500 4796 546
rect 4907 575 4953 634
rect 4907 512 4953 529
rect 4223 406 4269 423
rect 4583 439 4629 450
rect 3736 336 3782 361
rect 4131 327 4177 385
rect 3831 311 4082 327
rect 3615 244 3661 302
rect 3831 265 4023 311
rect 4069 265 4082 311
rect 4131 299 4583 327
rect 4131 281 4629 299
rect 3831 242 4082 265
rect 3615 158 3661 198
rect 4007 204 4082 242
rect 4335 219 4381 281
rect 2996 106 3569 152
rect 3872 137 3883 183
rect 3929 137 3940 183
rect 3872 60 3940 137
rect 4007 133 4140 204
rect 4692 202 4796 500
rect 4335 162 4381 173
rect 4479 168 4525 185
rect 4479 60 4525 122
rect 4692 156 4703 202
rect 4749 156 4796 202
rect 4692 120 4796 156
rect 4927 168 4973 185
rect 4927 60 4973 122
rect 0 -60 5040 60
<< labels >>
flabel metal1 s 4692 120 4796 672 0 FreeSans 400 0 0 0 Q
port 6 nsew default output
flabel metal1 s 3831 242 4082 327 0 FreeSans 400 0 0 0 RN
port 2 nsew default input
flabel metal1 s 141 119 206 430 0 FreeSans 400 0 0 0 SE
port 3 nsew default input
flabel metal1 s 365 119 430 430 0 FreeSans 400 0 0 0 SI
port 4 nsew default input
flabel metal1 s 0 724 5040 844 0 FreeSans 400 0 0 0 VDD
port 7 nsew power bidirectional abutment
flabel metal1 s 273 209 319 228 0 FreeSans 400 0 0 0 VSS
port 10 nsew ground bidirectional abutment
flabel metal1 s 1026 353 1326 431 0 FreeSans 400 0 0 0 CLK
port 5 nsew clock input
flabel metal1 s 619 353 878 438 0 FreeSans 400 0 0 0 D
port 1 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 8 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 9 nsew ground bidirectional
rlabel metal1 s 4007 204 4082 242 1 RN
port 2 nsew default input
rlabel metal1 s 4007 133 4140 204 1 RN
port 2 nsew default input
rlabel metal1 s 4907 670 4953 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4489 670 4535 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4335 670 4381 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3896 670 3964 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3027 670 3073 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2624 670 2692 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1518 670 1586 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1075 670 1121 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 252 670 320 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4907 600 4953 670 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4489 600 4535 670 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4335 600 4381 670 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3896 600 3964 670 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3027 600 3073 670 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2624 600 2692 670 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1075 600 1121 670 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 252 600 320 670 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4907 577 4953 600 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4489 577 4535 600 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4335 577 4381 600 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3896 577 3964 600 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3027 577 3073 600 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1075 577 1121 600 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 252 577 320 600 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4907 569 4953 577 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4489 569 4535 577 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4335 569 4381 577 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3896 569 3964 577 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3027 569 3073 577 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 252 569 320 577 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4907 533 4953 569 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4489 533 4535 569 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4335 533 4381 569 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3027 533 3073 569 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4907 514 4953 533 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4489 514 4535 533 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4335 514 4381 533 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4907 512 4953 514 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4489 512 4535 514 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1573 205 1619 209 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 273 205 319 209 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 1573 185 1619 205 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 1110 185 1156 205 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 273 185 319 205 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 4927 183 4973 185 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 4479 183 4525 185 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 1573 183 1619 185 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 1110 183 1156 185 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 273 183 319 185 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 4927 60 4973 183 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 4479 60 4525 183 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 3872 60 3940 183 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 2874 60 2942 183 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 1573 60 1619 183 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 1110 60 1156 183 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 273 60 319 183 1 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 5040 60 1 VSS
port 10 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 5040 784
string GDS_END 232690
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 221860
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
