magic
tech gf180mcuD
timestamp 1698431365
<< properties >>
string GDS_END 13421480
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 13231460
<< end >>
