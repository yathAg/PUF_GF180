magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< polysilicon >>
rect 794 8377 972 8396
rect 794 8331 813 8377
rect 953 8331 972 8377
rect 794 8312 972 8331
rect 2598 8377 2776 8396
rect 2598 8331 2617 8377
rect 2757 8331 2776 8377
rect 2598 8312 2776 8331
rect 3002 8377 3180 8396
rect 3002 8331 3021 8377
rect 3161 8331 3180 8377
rect 3002 8312 3180 8331
rect 4806 8377 4984 8396
rect 4806 8331 4825 8377
rect 4965 8331 4984 8377
rect 4806 8312 4984 8331
rect 5210 8377 5388 8396
rect 5210 8331 5229 8377
rect 5369 8331 5388 8377
rect 5210 8312 5388 8331
rect 7014 8377 7192 8396
rect 7014 8331 7033 8377
rect 7173 8331 7192 8377
rect 7014 8312 7192 8331
rect 7418 8377 7596 8396
rect 7418 8331 7437 8377
rect 7577 8331 7596 8377
rect 7418 8312 7596 8331
rect 9222 8377 9400 8396
rect 9222 8331 9241 8377
rect 9381 8331 9400 8377
rect 9222 8312 9400 8331
rect 803 8300 963 8312
rect 2607 8300 2767 8312
rect 3011 8300 3171 8312
rect 4815 8300 4975 8312
rect 5219 8300 5379 8312
rect 7023 8300 7183 8312
rect 7427 8300 7587 8312
rect 9231 8300 9391 8312
rect 794 706 972 725
rect 794 660 813 706
rect 953 660 972 706
rect 794 641 972 660
rect 2598 706 2776 725
rect 2598 660 2617 706
rect 2757 660 2776 706
rect 2598 641 2776 660
rect 3002 706 3180 725
rect 3002 660 3021 706
rect 3161 660 3180 706
rect 3002 641 3180 660
rect 4806 706 4984 725
rect 4806 660 4825 706
rect 4965 660 4984 706
rect 4806 641 4984 660
rect 5211 706 5389 725
rect 5211 660 5230 706
rect 5370 660 5389 706
rect 5211 641 5389 660
rect 7014 706 7192 725
rect 7014 660 7033 706
rect 7173 660 7192 706
rect 7014 641 7192 660
rect 7417 706 7595 725
rect 7417 660 7436 706
rect 7576 660 7595 706
rect 7417 641 7595 660
rect 9222 706 9400 725
rect 9222 660 9241 706
rect 9381 660 9400 706
rect 9222 641 9400 660
<< polycontact >>
rect 813 8331 953 8377
rect 2617 8331 2757 8377
rect 3021 8331 3161 8377
rect 4825 8331 4965 8377
rect 5229 8331 5369 8377
rect 7033 8331 7173 8377
rect 7437 8331 7577 8377
rect 9241 8331 9381 8377
rect 813 660 953 706
rect 2617 660 2757 706
rect 3021 660 3161 706
rect 4825 660 4965 706
rect 5230 660 5370 706
rect 7033 660 7173 706
rect 7436 660 7576 706
rect 9241 660 9381 706
<< metal1 >>
rect -251 9400 4976 9508
rect -251 9240 3172 9340
rect -251 9080 2768 9180
rect -251 8920 964 9020
rect 802 8377 964 8920
rect 802 8331 813 8377
rect 953 8331 964 8377
rect 802 8320 964 8331
rect 2606 8377 2768 9080
rect 2606 8331 2617 8377
rect 2757 8331 2768 8377
rect 2606 8320 2768 8331
rect 3010 8377 3172 9240
rect 3010 8331 3021 8377
rect 3161 8331 3172 8377
rect 3010 8320 3172 8331
rect 4814 8377 4976 9400
rect 4814 8331 4825 8377
rect 4965 8331 4976 8377
rect 4814 8320 4976 8331
rect 5218 9400 10510 9508
rect 5218 8377 5380 9400
rect 5218 8331 5229 8377
rect 5369 8331 5380 8377
rect 5218 8320 5380 8331
rect 7022 9240 10510 9340
rect 7022 8377 7184 9240
rect 7022 8331 7033 8377
rect 7173 8331 7184 8377
rect 7022 8320 7184 8331
rect 7426 9080 10510 9180
rect 7426 8377 7588 9080
rect 7426 8331 7437 8377
rect 7577 8331 7588 8377
rect 7426 8320 7588 8331
rect 9230 8920 10510 9020
rect 9230 8377 9392 8920
rect 9230 8331 9241 8377
rect 9381 8331 9392 8377
rect 9230 8320 9392 8331
rect 302 363 559 8212
rect 849 717 895 8320
rect 2675 717 2721 8320
rect 3057 717 3103 8320
rect 4883 717 4929 8320
rect 5265 717 5311 8320
rect 7091 717 7137 8320
rect 7473 717 7519 8320
rect 9299 717 9345 8320
rect 9391 812 9967 8212
rect 802 706 964 717
rect 802 660 813 706
rect 953 660 964 706
rect 802 649 964 660
rect 2606 706 2768 717
rect 2606 660 2617 706
rect 2757 660 2768 706
rect 2606 649 2768 660
rect 3010 706 3172 717
rect 3010 660 3021 706
rect 3161 660 3172 706
rect 3010 649 3172 660
rect 4814 706 4976 717
rect 4814 660 4825 706
rect 4965 660 4976 706
rect 4814 649 4976 660
rect 5219 706 5381 717
rect 5219 660 5230 706
rect 5370 660 5381 706
rect 5219 649 5381 660
rect 7022 706 7184 717
rect 7022 660 7033 706
rect 7173 660 7184 706
rect 7022 649 7184 660
rect 7425 706 7587 717
rect 7425 660 7436 706
rect 7576 660 7587 706
rect 7425 649 7587 660
rect 9230 706 9392 717
rect 9230 660 9241 706
rect 9381 660 9392 706
rect 9230 649 9392 660
rect 9730 363 9967 812
use comp018green_out_drv_nleg_6T  comp018green_out_drv_nleg_6T_0
timestamp 1698431365
transform 1 0 7221 0 1 680
box 48 44 2328 7632
use comp018green_out_drv_nleg_6T  comp018green_out_drv_nleg_6T_1
timestamp 1698431365
transform 1 0 5013 0 1 680
box 48 44 2328 7632
use comp018green_out_drv_nleg_6T  comp018green_out_drv_nleg_6T_2
timestamp 1698431365
transform 1 0 2805 0 1 680
box 48 44 2328 7632
use comp018green_out_drv_nleg_6T  comp018green_out_drv_nleg_6T_3
timestamp 1698431365
transform 1 0 597 0 1 680
box 48 44 2328 7632
use GR_NMOS  GR_NMOS_0
timestamp 1698431365
transform 1 0 363 0 1 436
box -1789 -834 11222 10481
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_0
timestamp 1698431365
transform 0 1 9311 1 0 8354
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_1
timestamp 1698431365
transform 0 1 5299 1 0 8354
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_2
timestamp 1698431365
transform 0 1 7103 1 0 8354
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_3
timestamp 1698431365
transform 0 1 7507 1 0 8354
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_4
timestamp 1698431365
transform 0 -1 4895 1 0 683
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_5
timestamp 1698431365
transform 0 -1 9311 1 0 683
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_6
timestamp 1698431365
transform 0 -1 7506 1 0 683
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_7
timestamp 1698431365
transform 0 -1 7103 1 0 683
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_8
timestamp 1698431365
transform 0 -1 5300 1 0 683
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_9
timestamp 1698431365
transform 0 -1 3091 1 0 8354
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_10
timestamp 1698431365
transform 0 -1 2687 1 0 8354
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_11
timestamp 1698431365
transform 0 -1 4895 1 0 8354
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_12
timestamp 1698431365
transform 0 -1 883 1 0 8354
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_13
timestamp 1698431365
transform 0 -1 3091 1 0 683
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_14
timestamp 1698431365
transform 0 -1 883 1 0 683
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_15
timestamp 1698431365
transform 0 -1 2687 1 0 683
box 0 0 1 1
use nmos_metal_stack  nmos_metal_stack_0
timestamp 1698431365
transform -1 0 9591 0 1 812
box -44 0 2004 7400
use nmos_metal_stack  nmos_metal_stack_1
timestamp 1698431365
transform 1 0 7227 0 1 812
box -44 0 2004 7400
use nmos_metal_stack  nmos_metal_stack_2
timestamp 1698431365
transform 1 0 5019 0 1 812
box -44 0 2004 7400
use nmos_metal_stack  nmos_metal_stack_3
timestamp 1698431365
transform 1 0 2811 0 1 812
box -44 0 2004 7400
use nmos_metal_stack  nmos_metal_stack_4
timestamp 1698431365
transform 1 0 603 0 1 812
box -44 0 2004 7400
<< properties >>
string GDS_END 2348664
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 2343818
string path 233.050 208.025 233.050 17.675 
<< end >>
