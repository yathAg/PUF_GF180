magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 352 3894 870
<< pwell >>
rect -86 -86 3894 352
<< mvnmos >>
rect 124 68 244 232
rect 348 68 468 232
rect 572 68 692 232
rect 796 68 916 232
rect 1020 68 1140 232
rect 1244 68 1364 232
rect 1468 68 1588 232
rect 1692 68 1812 232
rect 1916 68 2036 232
rect 2140 68 2260 232
rect 2364 68 2484 232
rect 2588 68 2708 232
rect 2812 68 2932 232
rect 3036 68 3156 232
rect 3260 68 3380 232
rect 3484 68 3604 232
<< mvpmos >>
rect 124 472 224 716
rect 348 472 448 716
rect 572 472 672 716
rect 796 472 896 716
rect 1020 472 1120 716
rect 1244 472 1344 716
rect 1468 472 1568 716
rect 1692 472 1792 716
rect 1916 472 2016 716
rect 2140 472 2240 716
rect 2364 472 2464 716
rect 2588 472 2688 716
rect 2812 472 2912 716
rect 3036 472 3136 716
rect 3260 472 3360 716
rect 3484 472 3584 716
<< mvndiff >>
rect 36 192 124 232
rect 36 146 49 192
rect 95 146 124 192
rect 36 68 124 146
rect 244 192 348 232
rect 244 146 273 192
rect 319 146 348 192
rect 244 68 348 146
rect 468 127 572 232
rect 468 81 497 127
rect 543 81 572 127
rect 468 68 572 81
rect 692 192 796 232
rect 692 146 721 192
rect 767 146 796 192
rect 692 68 796 146
rect 916 127 1020 232
rect 916 81 945 127
rect 991 81 1020 127
rect 916 68 1020 81
rect 1140 192 1244 232
rect 1140 146 1169 192
rect 1215 146 1244 192
rect 1140 68 1244 146
rect 1364 127 1468 232
rect 1364 81 1393 127
rect 1439 81 1468 127
rect 1364 68 1468 81
rect 1588 192 1692 232
rect 1588 146 1617 192
rect 1663 146 1692 192
rect 1588 68 1692 146
rect 1812 127 1916 232
rect 1812 81 1841 127
rect 1887 81 1916 127
rect 1812 68 1916 81
rect 2036 192 2140 232
rect 2036 146 2065 192
rect 2111 146 2140 192
rect 2036 68 2140 146
rect 2260 127 2364 232
rect 2260 81 2289 127
rect 2335 81 2364 127
rect 2260 68 2364 81
rect 2484 192 2588 232
rect 2484 146 2513 192
rect 2559 146 2588 192
rect 2484 68 2588 146
rect 2708 127 2812 232
rect 2708 81 2737 127
rect 2783 81 2812 127
rect 2708 68 2812 81
rect 2932 192 3036 232
rect 2932 146 2961 192
rect 3007 146 3036 192
rect 2932 68 3036 146
rect 3156 127 3260 232
rect 3156 81 3185 127
rect 3231 81 3260 127
rect 3156 68 3260 81
rect 3380 192 3484 232
rect 3380 146 3409 192
rect 3455 146 3484 192
rect 3380 68 3484 146
rect 3604 192 3692 232
rect 3604 146 3633 192
rect 3679 146 3692 192
rect 3604 68 3692 146
<< mvpdiff >>
rect 36 687 124 716
rect 36 547 49 687
rect 95 547 124 687
rect 36 472 124 547
rect 224 665 348 716
rect 224 525 273 665
rect 319 525 348 665
rect 224 472 348 525
rect 448 703 572 716
rect 448 657 477 703
rect 523 657 572 703
rect 448 472 572 657
rect 672 665 796 716
rect 672 525 701 665
rect 747 525 796 665
rect 672 472 796 525
rect 896 703 1020 716
rect 896 657 925 703
rect 971 657 1020 703
rect 896 472 1020 657
rect 1120 665 1244 716
rect 1120 525 1149 665
rect 1195 525 1244 665
rect 1120 472 1244 525
rect 1344 703 1468 716
rect 1344 657 1373 703
rect 1419 657 1468 703
rect 1344 472 1468 657
rect 1568 665 1692 716
rect 1568 525 1616 665
rect 1662 525 1692 665
rect 1568 472 1692 525
rect 1792 703 1916 716
rect 1792 657 1821 703
rect 1867 657 1916 703
rect 1792 472 1916 657
rect 2016 665 2140 716
rect 2016 525 2045 665
rect 2091 525 2140 665
rect 2016 472 2140 525
rect 2240 703 2364 716
rect 2240 657 2269 703
rect 2315 657 2364 703
rect 2240 472 2364 657
rect 2464 665 2588 716
rect 2464 525 2493 665
rect 2539 525 2588 665
rect 2464 472 2588 525
rect 2688 703 2812 716
rect 2688 657 2717 703
rect 2763 657 2812 703
rect 2688 472 2812 657
rect 2912 665 3036 716
rect 2912 525 2941 665
rect 2987 525 3036 665
rect 2912 472 3036 525
rect 3136 703 3260 716
rect 3136 657 3165 703
rect 3211 657 3260 703
rect 3136 472 3260 657
rect 3360 665 3484 716
rect 3360 525 3389 665
rect 3435 525 3484 665
rect 3360 472 3484 525
rect 3584 687 3672 716
rect 3584 547 3613 687
rect 3659 547 3672 687
rect 3584 472 3672 547
<< mvndiffc >>
rect 49 146 95 192
rect 273 146 319 192
rect 497 81 543 127
rect 721 146 767 192
rect 945 81 991 127
rect 1169 146 1215 192
rect 1393 81 1439 127
rect 1617 146 1663 192
rect 1841 81 1887 127
rect 2065 146 2111 192
rect 2289 81 2335 127
rect 2513 146 2559 192
rect 2737 81 2783 127
rect 2961 146 3007 192
rect 3185 81 3231 127
rect 3409 146 3455 192
rect 3633 146 3679 192
<< mvpdiffc >>
rect 49 547 95 687
rect 273 525 319 665
rect 477 657 523 703
rect 701 525 747 665
rect 925 657 971 703
rect 1149 525 1195 665
rect 1373 657 1419 703
rect 1616 525 1662 665
rect 1821 657 1867 703
rect 2045 525 2091 665
rect 2269 657 2315 703
rect 2493 525 2539 665
rect 2717 657 2763 703
rect 2941 525 2987 665
rect 3165 657 3211 703
rect 3389 525 3435 665
rect 3613 547 3659 687
<< polysilicon >>
rect 124 716 224 760
rect 348 716 448 760
rect 572 716 672 760
rect 796 716 896 760
rect 1020 716 1120 760
rect 1244 716 1344 760
rect 1468 716 1568 760
rect 1692 716 1792 760
rect 1916 716 2016 760
rect 2140 716 2240 760
rect 2364 716 2464 760
rect 2588 716 2688 760
rect 2812 716 2912 760
rect 3036 716 3136 760
rect 3260 716 3360 760
rect 3484 716 3584 760
rect 124 412 224 472
rect 348 412 448 472
rect 572 412 672 472
rect 796 412 896 472
rect 1020 412 1120 472
rect 1244 412 1344 472
rect 1468 412 1568 472
rect 1692 412 1792 472
rect 1916 412 2016 472
rect 2140 412 2240 472
rect 2364 412 2464 472
rect 2588 412 2688 472
rect 2812 412 2912 472
rect 3036 412 3136 472
rect 3260 412 3360 472
rect 3484 412 3584 472
rect 124 399 3584 412
rect 124 353 137 399
rect 1687 353 2016 399
rect 3566 353 3584 399
rect 124 340 3584 353
rect 124 232 244 340
rect 348 232 468 340
rect 572 232 692 340
rect 796 232 916 340
rect 1020 232 1140 340
rect 1244 232 1364 340
rect 1468 232 1588 340
rect 1692 232 1812 340
rect 1916 232 2036 340
rect 2140 232 2260 340
rect 2364 232 2484 340
rect 2588 232 2708 340
rect 2812 232 2932 340
rect 3036 232 3156 340
rect 3260 232 3380 340
rect 3484 288 3584 340
rect 3484 232 3604 288
rect 124 24 244 68
rect 348 24 468 68
rect 572 24 692 68
rect 796 24 916 68
rect 1020 24 1140 68
rect 1244 24 1364 68
rect 1468 24 1588 68
rect 1692 24 1812 68
rect 1916 24 2036 68
rect 2140 24 2260 68
rect 2364 24 2484 68
rect 2588 24 2708 68
rect 2812 24 2932 68
rect 3036 24 3156 68
rect 3260 24 3380 68
rect 3484 24 3604 68
<< polycontact >>
rect 137 353 1687 399
rect 2016 353 3566 399
<< metal1 >>
rect 0 724 3808 844
rect 49 687 95 724
rect 477 703 523 724
rect 49 536 95 547
rect 273 665 319 678
rect 925 703 971 724
rect 477 646 523 657
rect 701 665 747 678
rect 319 525 701 600
rect 1373 703 1419 724
rect 925 646 971 657
rect 1149 665 1195 678
rect 747 525 1149 600
rect 1821 703 1867 724
rect 1373 646 1419 657
rect 1616 665 1662 678
rect 1195 525 1616 600
rect 2269 703 2315 724
rect 1821 646 1867 657
rect 2045 665 2091 678
rect 1662 525 2045 600
rect 2717 703 2763 724
rect 2269 646 2315 657
rect 2493 665 2539 678
rect 2091 525 2493 600
rect 3165 703 3211 724
rect 2717 646 2763 657
rect 2941 665 2987 678
rect 2539 525 2941 600
rect 3613 687 3659 724
rect 3165 646 3211 657
rect 3389 665 3435 678
rect 2987 525 3389 600
rect 3613 536 3659 547
rect 273 484 3435 525
rect 124 399 1702 438
rect 124 353 137 399
rect 1687 353 1702 399
rect 1758 289 1938 484
rect 2003 399 3584 438
rect 2003 353 2016 399
rect 3566 353 3584 399
rect 49 192 95 203
rect 49 60 95 146
rect 273 192 3455 289
rect 319 173 721 192
rect 319 146 325 173
rect 273 135 325 146
rect 767 173 1169 192
rect 721 135 767 146
rect 1215 173 1617 192
rect 1169 135 1215 146
rect 1663 173 2065 192
rect 1617 135 1663 146
rect 2111 173 2513 192
rect 2065 135 2111 146
rect 2559 173 2961 192
rect 2513 135 2559 146
rect 3007 173 3409 192
rect 2961 135 3007 146
rect 3409 135 3455 146
rect 3633 192 3679 203
rect 486 81 497 127
rect 543 81 554 127
rect 486 60 554 81
rect 934 81 945 127
rect 991 81 1002 127
rect 934 60 1002 81
rect 1382 81 1393 127
rect 1439 81 1450 127
rect 1382 60 1450 81
rect 1830 81 1841 127
rect 1887 81 1898 127
rect 1830 60 1898 81
rect 2278 81 2289 127
rect 2335 81 2346 127
rect 2278 60 2346 81
rect 2726 81 2737 127
rect 2783 81 2794 127
rect 2726 60 2794 81
rect 3174 81 3185 127
rect 3231 81 3242 127
rect 3174 60 3242 81
rect 3633 60 3679 146
rect 0 -60 3808 60
<< labels >>
flabel metal1 s 3633 127 3679 203 0 FreeSans 400 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel metal1 s 3389 600 3435 678 0 FreeSans 400 0 0 0 ZN
port 2 nsew default output
flabel metal1 s 124 353 1702 438 0 FreeSans 400 0 0 0 I
port 1 nsew default input
flabel metal1 s 0 724 3808 844 0 FreeSans 400 0 0 0 VDD
port 3 nsew power bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 4 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 2003 353 3584 438 1 I
port 1 nsew default input
rlabel metal1 s 2941 600 2987 678 1 ZN
port 2 nsew default output
rlabel metal1 s 2493 600 2539 678 1 ZN
port 2 nsew default output
rlabel metal1 s 2045 600 2091 678 1 ZN
port 2 nsew default output
rlabel metal1 s 1616 600 1662 678 1 ZN
port 2 nsew default output
rlabel metal1 s 1149 600 1195 678 1 ZN
port 2 nsew default output
rlabel metal1 s 701 600 747 678 1 ZN
port 2 nsew default output
rlabel metal1 s 273 600 319 678 1 ZN
port 2 nsew default output
rlabel metal1 s 273 484 3435 600 1 ZN
port 2 nsew default output
rlabel metal1 s 1758 289 1938 484 1 ZN
port 2 nsew default output
rlabel metal1 s 273 173 3455 289 1 ZN
port 2 nsew default output
rlabel metal1 s 3409 135 3455 173 1 ZN
port 2 nsew default output
rlabel metal1 s 2961 135 3007 173 1 ZN
port 2 nsew default output
rlabel metal1 s 2513 135 2559 173 1 ZN
port 2 nsew default output
rlabel metal1 s 2065 135 2111 173 1 ZN
port 2 nsew default output
rlabel metal1 s 1617 135 1663 173 1 ZN
port 2 nsew default output
rlabel metal1 s 1169 135 1215 173 1 ZN
port 2 nsew default output
rlabel metal1 s 721 135 767 173 1 ZN
port 2 nsew default output
rlabel metal1 s 273 135 325 173 1 ZN
port 2 nsew default output
rlabel metal1 s 3613 646 3659 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3165 646 3211 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2717 646 2763 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2269 646 2315 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1821 646 1867 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1373 646 1419 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 925 646 971 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 477 646 523 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 646 95 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3613 536 3659 646 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 536 95 646 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 127 95 203 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3633 60 3679 127 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3174 60 3242 127 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2726 60 2794 127 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2278 60 2346 127 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1830 60 1898 127 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1382 60 1450 127 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 934 60 1002 127 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 486 60 554 127 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 127 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3808 60 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3808 784
string GDS_END 506636
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 497912
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
