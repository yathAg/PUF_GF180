magic
tech gf180mcuB
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 453 3670 1094
<< pwell >>
rect -86 -86 3670 453
<< metal1 >>
rect 0 918 3584 1098
rect 0 -90 3584 90
<< labels >>
rlabel metal1 s 0 918 3584 1098 6 VDD
port 1 nsew power bidirectional abutment
rlabel nwell s -86 453 3670 1094 6 VNW
port 2 nsew power bidirectional
rlabel pwell s -86 -86 3670 453 6 VPW
port 3 nsew ground bidirectional
rlabel metal1 s 0 -90 3584 90 8 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3584 1008
string LEFclass core SPACER
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 772408
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 771246
<< end >>
