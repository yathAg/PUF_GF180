magic
tech gf180mcuD
magscale 1 10
timestamp 1698431365
<< psubdiff >>
rect 0 69842 200 69968
rect 0 13186 77 69842
rect 123 13186 200 69842
rect 0 13097 200 13186
<< psubdiffcont >>
rect 77 13186 123 69842
<< metal1 >>
rect -32 69842 232 69957
rect -32 64942 77 69842
rect 123 64942 232 69842
rect -32 64890 75 64942
rect 127 64890 232 64942
rect -32 64830 77 64890
rect 123 64830 232 64890
rect -32 64778 75 64830
rect 127 64778 232 64830
rect -32 64718 77 64778
rect 123 64718 232 64778
rect -32 64666 75 64718
rect 127 64666 232 64718
rect -32 64606 77 64666
rect 123 64606 232 64666
rect -32 64554 75 64606
rect 127 64554 232 64606
rect -32 64494 77 64554
rect 123 64494 232 64554
rect -32 64442 75 64494
rect 127 64442 232 64494
rect -32 64382 77 64442
rect 123 64382 232 64442
rect -32 64330 75 64382
rect 127 64330 232 64382
rect -32 64270 77 64330
rect 123 64270 232 64330
rect -32 64218 75 64270
rect 127 64218 232 64270
rect -32 64158 77 64218
rect 123 64158 232 64218
rect -32 64106 75 64158
rect 127 64106 232 64158
rect -32 64046 77 64106
rect 123 64046 232 64106
rect -32 63994 75 64046
rect 127 63994 232 64046
rect -32 63934 77 63994
rect 123 63934 232 63994
rect -32 63882 75 63934
rect 127 63882 232 63934
rect -32 63822 77 63882
rect 123 63822 232 63882
rect -32 63770 75 63822
rect 127 63770 232 63822
rect -32 63710 77 63770
rect 123 63710 232 63770
rect -32 63658 75 63710
rect 127 63658 232 63710
rect -32 50536 77 63658
rect 123 50536 232 63658
rect -32 50484 76 50536
rect 128 50484 232 50536
rect -32 50424 77 50484
rect 123 50424 232 50484
rect -32 50372 76 50424
rect 128 50372 232 50424
rect -32 50312 77 50372
rect 123 50312 232 50372
rect -32 50260 76 50312
rect 128 50260 232 50312
rect -32 50200 77 50260
rect 123 50200 232 50260
rect -32 50148 76 50200
rect 128 50148 232 50200
rect -32 50088 77 50148
rect 123 50088 232 50148
rect -32 50036 76 50088
rect 128 50036 232 50088
rect -32 49976 77 50036
rect 123 49976 232 50036
rect -32 49924 76 49976
rect 128 49924 232 49976
rect -32 49864 77 49924
rect 123 49864 232 49924
rect -32 49812 76 49864
rect 128 49812 232 49864
rect -32 49752 77 49812
rect 123 49752 232 49812
rect -32 49700 76 49752
rect 128 49700 232 49752
rect -32 49640 77 49700
rect 123 49640 232 49700
rect -32 49588 76 49640
rect 128 49588 232 49640
rect -32 49528 77 49588
rect 123 49528 232 49588
rect -32 49476 76 49528
rect 128 49476 232 49528
rect -32 49416 77 49476
rect 123 49416 232 49476
rect -32 49364 76 49416
rect 128 49364 232 49416
rect -32 49304 77 49364
rect 123 49304 232 49364
rect -32 49252 76 49304
rect 128 49252 232 49304
rect -32 13186 77 49252
rect 123 13186 232 49252
rect -32 13097 232 13186
<< via1 >>
rect 75 64890 77 64942
rect 77 64890 123 64942
rect 123 64890 127 64942
rect 75 64778 77 64830
rect 77 64778 123 64830
rect 123 64778 127 64830
rect 75 64666 77 64718
rect 77 64666 123 64718
rect 123 64666 127 64718
rect 75 64554 77 64606
rect 77 64554 123 64606
rect 123 64554 127 64606
rect 75 64442 77 64494
rect 77 64442 123 64494
rect 123 64442 127 64494
rect 75 64330 77 64382
rect 77 64330 123 64382
rect 123 64330 127 64382
rect 75 64218 77 64270
rect 77 64218 123 64270
rect 123 64218 127 64270
rect 75 64106 77 64158
rect 77 64106 123 64158
rect 123 64106 127 64158
rect 75 63994 77 64046
rect 77 63994 123 64046
rect 123 63994 127 64046
rect 75 63882 77 63934
rect 77 63882 123 63934
rect 123 63882 127 63934
rect 75 63770 77 63822
rect 77 63770 123 63822
rect 123 63770 127 63822
rect 75 63658 77 63710
rect 77 63658 123 63710
rect 123 63658 127 63710
rect 76 50484 77 50536
rect 77 50484 123 50536
rect 123 50484 128 50536
rect 76 50372 77 50424
rect 77 50372 123 50424
rect 123 50372 128 50424
rect 76 50260 77 50312
rect 77 50260 123 50312
rect 123 50260 128 50312
rect 76 50148 77 50200
rect 77 50148 123 50200
rect 123 50148 128 50200
rect 76 50036 77 50088
rect 77 50036 123 50088
rect 123 50036 128 50088
rect 76 49924 77 49976
rect 77 49924 123 49976
rect 123 49924 128 49976
rect 76 49812 77 49864
rect 77 49812 123 49864
rect 123 49812 128 49864
rect 76 49700 77 49752
rect 77 49700 123 49752
rect 123 49700 128 49752
rect 76 49588 77 49640
rect 77 49588 123 49640
rect 123 49588 128 49640
rect 76 49476 77 49528
rect 77 49476 123 49528
rect 123 49476 128 49528
rect 76 49364 77 49416
rect 77 49364 123 49416
rect 123 49364 128 49416
rect 76 49252 77 49304
rect 77 49252 123 49304
rect 123 49252 128 49304
<< metal2 >>
rect 0 64944 200 65000
rect 0 64888 73 64944
rect 129 64888 200 64944
rect 0 64832 200 64888
rect 0 64776 73 64832
rect 129 64776 200 64832
rect 0 64720 200 64776
rect 0 64664 73 64720
rect 129 64664 200 64720
rect 0 64608 200 64664
rect 0 64552 73 64608
rect 129 64552 200 64608
rect 0 64496 200 64552
rect 0 64440 73 64496
rect 129 64440 200 64496
rect 0 64384 200 64440
rect 0 64328 73 64384
rect 129 64328 200 64384
rect 0 64272 200 64328
rect 0 64216 73 64272
rect 129 64216 200 64272
rect 0 64160 200 64216
rect 0 64104 73 64160
rect 129 64104 200 64160
rect 0 64048 200 64104
rect 0 63992 73 64048
rect 129 63992 200 64048
rect 0 63936 200 63992
rect 0 63880 73 63936
rect 129 63880 200 63936
rect 0 63824 200 63880
rect 0 63768 73 63824
rect 129 63768 200 63824
rect 0 63712 200 63768
rect 0 63656 73 63712
rect 129 63656 200 63712
rect 0 63600 200 63656
rect 0 50538 200 50600
rect 0 50482 74 50538
rect 130 50482 200 50538
rect 0 50426 200 50482
rect 0 50370 74 50426
rect 130 50370 200 50426
rect 0 50314 200 50370
rect 0 50258 74 50314
rect 130 50258 200 50314
rect 0 50202 200 50258
rect 0 50146 74 50202
rect 130 50146 200 50202
rect 0 50090 200 50146
rect 0 50034 74 50090
rect 130 50034 200 50090
rect 0 49978 200 50034
rect 0 49922 74 49978
rect 130 49922 200 49978
rect 0 49866 200 49922
rect 0 49810 74 49866
rect 130 49810 200 49866
rect 0 49754 200 49810
rect 0 49698 74 49754
rect 130 49698 200 49754
rect 0 49642 200 49698
rect 0 49586 74 49642
rect 130 49586 200 49642
rect 0 49530 200 49586
rect 0 49474 74 49530
rect 130 49474 200 49530
rect 0 49418 200 49474
rect 0 49362 74 49418
rect 130 49362 200 49418
rect 0 49306 200 49362
rect 0 49250 74 49306
rect 130 49250 200 49306
rect 0 49200 200 49250
<< via2 >>
rect 73 64942 129 64944
rect 73 64890 75 64942
rect 75 64890 127 64942
rect 127 64890 129 64942
rect 73 64888 129 64890
rect 73 64830 129 64832
rect 73 64778 75 64830
rect 75 64778 127 64830
rect 127 64778 129 64830
rect 73 64776 129 64778
rect 73 64718 129 64720
rect 73 64666 75 64718
rect 75 64666 127 64718
rect 127 64666 129 64718
rect 73 64664 129 64666
rect 73 64606 129 64608
rect 73 64554 75 64606
rect 75 64554 127 64606
rect 127 64554 129 64606
rect 73 64552 129 64554
rect 73 64494 129 64496
rect 73 64442 75 64494
rect 75 64442 127 64494
rect 127 64442 129 64494
rect 73 64440 129 64442
rect 73 64382 129 64384
rect 73 64330 75 64382
rect 75 64330 127 64382
rect 127 64330 129 64382
rect 73 64328 129 64330
rect 73 64270 129 64272
rect 73 64218 75 64270
rect 75 64218 127 64270
rect 127 64218 129 64270
rect 73 64216 129 64218
rect 73 64158 129 64160
rect 73 64106 75 64158
rect 75 64106 127 64158
rect 127 64106 129 64158
rect 73 64104 129 64106
rect 73 64046 129 64048
rect 73 63994 75 64046
rect 75 63994 127 64046
rect 127 63994 129 64046
rect 73 63992 129 63994
rect 73 63934 129 63936
rect 73 63882 75 63934
rect 75 63882 127 63934
rect 127 63882 129 63934
rect 73 63880 129 63882
rect 73 63822 129 63824
rect 73 63770 75 63822
rect 75 63770 127 63822
rect 127 63770 129 63822
rect 73 63768 129 63770
rect 73 63710 129 63712
rect 73 63658 75 63710
rect 75 63658 127 63710
rect 127 63658 129 63710
rect 73 63656 129 63658
rect 74 50536 130 50538
rect 74 50484 76 50536
rect 76 50484 128 50536
rect 128 50484 130 50536
rect 74 50482 130 50484
rect 74 50424 130 50426
rect 74 50372 76 50424
rect 76 50372 128 50424
rect 128 50372 130 50424
rect 74 50370 130 50372
rect 74 50312 130 50314
rect 74 50260 76 50312
rect 76 50260 128 50312
rect 128 50260 130 50312
rect 74 50258 130 50260
rect 74 50200 130 50202
rect 74 50148 76 50200
rect 76 50148 128 50200
rect 128 50148 130 50200
rect 74 50146 130 50148
rect 74 50088 130 50090
rect 74 50036 76 50088
rect 76 50036 128 50088
rect 128 50036 130 50088
rect 74 50034 130 50036
rect 74 49976 130 49978
rect 74 49924 76 49976
rect 76 49924 128 49976
rect 128 49924 130 49976
rect 74 49922 130 49924
rect 74 49864 130 49866
rect 74 49812 76 49864
rect 76 49812 128 49864
rect 128 49812 130 49864
rect 74 49810 130 49812
rect 74 49752 130 49754
rect 74 49700 76 49752
rect 76 49700 128 49752
rect 128 49700 130 49752
rect 74 49698 130 49700
rect 74 49640 130 49642
rect 74 49588 76 49640
rect 76 49588 128 49640
rect 128 49588 130 49640
rect 74 49586 130 49588
rect 74 49528 130 49530
rect 74 49476 76 49528
rect 76 49476 128 49528
rect 128 49476 130 49528
rect 74 49474 130 49476
rect 74 49416 130 49418
rect 74 49364 76 49416
rect 76 49364 128 49416
rect 128 49364 130 49416
rect 74 49362 130 49364
rect 74 49304 130 49306
rect 74 49252 76 49304
rect 76 49252 128 49304
rect 128 49252 130 49304
rect 74 49250 130 49252
<< metal3 >>
rect 0 68400 200 69678
rect 0 66800 200 68200
rect 0 65200 200 66600
rect 0 64944 200 65000
rect 0 64888 73 64944
rect 129 64888 200 64944
rect 0 64832 200 64888
rect 0 64776 73 64832
rect 129 64776 200 64832
rect 0 64720 200 64776
rect 0 64664 73 64720
rect 129 64664 200 64720
rect 0 64608 200 64664
rect 0 64552 73 64608
rect 129 64552 200 64608
rect 0 64496 200 64552
rect 0 64440 73 64496
rect 129 64440 200 64496
rect 0 64384 200 64440
rect 0 64328 73 64384
rect 129 64328 200 64384
rect 0 64272 200 64328
rect 0 64216 73 64272
rect 129 64216 200 64272
rect 0 64160 200 64216
rect 0 64104 73 64160
rect 129 64104 200 64160
rect 0 64048 200 64104
rect 0 63992 73 64048
rect 129 63992 200 64048
rect 0 63936 200 63992
rect 0 63880 73 63936
rect 129 63880 200 63936
rect 0 63824 200 63880
rect 0 63768 73 63824
rect 129 63768 200 63824
rect 0 63712 200 63768
rect 0 63656 73 63712
rect 129 63656 200 63712
rect 0 63600 200 63656
rect 0 62000 200 63400
rect 0 60400 200 61800
rect 0 58800 200 60200
rect 0 57200 200 58600
rect 0 55600 200 57000
rect 0 54000 200 55400
rect 0 52400 200 53800
rect 0 50800 200 52200
rect 0 50538 200 50600
rect 0 50482 74 50538
rect 130 50482 200 50538
rect 0 50426 200 50482
rect 0 50370 74 50426
rect 130 50370 200 50426
rect 0 50314 200 50370
rect 0 50258 74 50314
rect 130 50258 200 50314
rect 0 50202 200 50258
rect 0 50146 74 50202
rect 130 50146 200 50202
rect 0 50090 200 50146
rect 0 50034 74 50090
rect 130 50034 200 50090
rect 0 49978 200 50034
rect 0 49922 74 49978
rect 130 49922 200 49978
rect 0 49866 200 49922
rect 0 49810 74 49866
rect 130 49810 200 49866
rect 0 49754 200 49810
rect 0 49698 74 49754
rect 130 49698 200 49754
rect 0 49642 200 49698
rect 0 49586 74 49642
rect 130 49586 200 49642
rect 0 49530 200 49586
rect 0 49474 74 49530
rect 130 49474 200 49530
rect 0 49418 200 49474
rect 0 49362 74 49418
rect 130 49362 200 49418
rect 0 49306 200 49362
rect 0 49250 74 49306
rect 130 49250 200 49306
rect 0 49200 200 49250
rect 0 46000 200 49000
rect 0 42800 200 45800
rect 0 41200 200 42600
rect 0 39600 200 41000
rect 0 36400 200 39400
rect 0 33200 200 36200
rect 0 30000 200 33000
rect 0 26800 200 29800
rect 0 25200 200 26600
rect 0 23600 200 25000
rect 0 20400 200 23400
rect 0 17200 200 20200
rect 0 14000 200 17000
use M1_PSUB_CDNS_4066195314525  M1_PSUB_CDNS_4066195314525_0
timestamp 1698431365
transform 1 0 100 0 1 41514
box 0 0 1 1
use M2_M1_CDNS_4066195314526  M2_M1_CDNS_4066195314526_0
timestamp 1698431365
transform 1 0 102 0 1 49894
box 0 0 1 1
use M2_M1_CDNS_4066195314527  M2_M1_CDNS_4066195314527_0
timestamp 1698431365
transform 1 0 101 0 1 64300
box 0 0 1 1
use M3_M2_CDNS_4066195314528  M3_M2_CDNS_4066195314528_0
timestamp 1698431365
transform 1 0 102 0 1 49894
box 0 0 1 1
use M3_M2_CDNS_4066195314529  M3_M2_CDNS_4066195314529_0
timestamp 1698431365
transform 1 0 101 0 1 64300
box 0 0 1 1
<< labels >>
rlabel metal3 s 94 64258 94 64258 4 VSS
port 1 nsew
rlabel metal3 s 94 50023 94 50023 4 VSS
port 1 nsew
rlabel metal3 s 94 51458 94 51458 4 VDD
port 2 nsew
rlabel metal3 s 94 62823 94 62823 4 VDD
port 2 nsew
rlabel metal3 s 94 18921 94 18921 4 DVSS
port 3 nsew
rlabel metal3 s 94 15750 94 15750 4 DVSS
port 3 nsew
rlabel metal3 s 94 21907 94 21907 4 DVSS
port 3 nsew
rlabel metal3 s 94 26100 94 26100 4 DVSS
port 3 nsew
rlabel metal3 s 94 40342 94 40342 4 DVSS
port 3 nsew
rlabel metal3 s 94 47595 94 47595 4 DVSS
port 3 nsew
rlabel metal3 s 94 57858 94 57858 4 DVSS
port 3 nsew
rlabel metal3 s 94 61058 94 61058 4 DVSS
port 3 nsew
rlabel metal3 s 94 66023 94 66023 4 DVSS
port 3 nsew
rlabel metal3 s 94 69049 94 69049 4 DVSS
port 3 nsew
rlabel metal3 s 94 67458 94 67458 4 DVDD
port 4 nsew
rlabel metal3 s 94 59623 94 59623 4 DVDD
port 4 nsew
rlabel metal3 s 94 56423 94 56423 4 DVDD
port 4 nsew
rlabel metal3 s 94 54658 94 54658 4 DVDD
port 4 nsew
rlabel metal3 s 94 53223 94 53223 4 DVDD
port 4 nsew
rlabel metal3 s 94 44368 94 44368 4 DVDD
port 4 nsew
rlabel metal3 s 94 41977 94 41977 4 DVDD
port 4 nsew
rlabel metal3 s 94 37959 94 37959 4 DVDD
port 4 nsew
rlabel metal3 s 94 34723 94 34723 4 DVDD
port 4 nsew
rlabel metal3 s 94 31609 94 31609 4 DVDD
port 4 nsew
rlabel metal3 s 94 28394 94 28394 4 DVDD
port 4 nsew
rlabel metal3 s 94 24284 94 24284 4 DVDD
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 200 70000
string GDS_END 5032048
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 5028714
<< end >>
