magic
tech gf180mcuB
magscale 1 5
timestamp 1698431365
<< nwell >>
rect -43 176 155 435
<< pwell >>
rect -43 -43 155 176
<< metal1 >>
rect 0 362 112 422
rect 0 -30 112 30
<< labels >>
rlabel metal1 s 0 362 112 422 6 VDD
port 1 nsew power bidirectional abutment
rlabel nwell s -43 176 155 435 6 VNW
port 2 nsew power bidirectional
rlabel pwell s -43 -43 155 176 6 VPW
port 3 nsew ground bidirectional
rlabel metal1 s 0 -30 112 30 8 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 112 392
string LEFclass core SPACER
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1148476
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1147316
<< end >>
