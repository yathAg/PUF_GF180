magic
tech gf180mcuD
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 352 3222 870
<< pwell >>
rect -86 -86 3222 352
<< mvnmos >>
rect 124 93 244 165
rect 348 93 468 165
rect 608 93 728 165
rect 832 93 952 165
rect 1016 93 1136 165
rect 1400 93 1520 165
rect 1624 93 1744 165
rect 1884 68 2004 232
rect 2108 68 2228 232
rect 2292 68 2412 232
rect 2668 68 2788 232
rect 2892 68 3012 232
<< mvpmos >>
rect 144 561 244 638
rect 368 561 468 638
rect 628 526 728 638
rect 832 526 932 638
rect 1036 526 1136 638
rect 1435 526 1535 638
rect 1644 526 1744 638
rect 1904 472 2004 716
rect 2123 472 2223 716
rect 2327 472 2427 716
rect 2678 472 2778 716
rect 2902 472 3002 716
<< mvndiff >>
rect 1804 165 1884 232
rect 36 152 124 165
rect 36 106 49 152
rect 95 106 124 152
rect 36 93 124 106
rect 244 152 348 165
rect 244 106 273 152
rect 319 106 348 152
rect 244 93 348 106
rect 468 152 608 165
rect 468 106 514 152
rect 560 106 608 152
rect 468 93 608 106
rect 728 152 832 165
rect 728 106 757 152
rect 803 106 832 152
rect 728 93 832 106
rect 952 93 1016 165
rect 1136 152 1224 165
rect 1136 106 1165 152
rect 1211 106 1224 152
rect 1136 93 1224 106
rect 1312 152 1400 165
rect 1312 106 1325 152
rect 1371 106 1400 152
rect 1312 93 1400 106
rect 1520 152 1624 165
rect 1520 106 1549 152
rect 1595 106 1624 152
rect 1520 93 1624 106
rect 1744 152 1884 165
rect 1744 106 1809 152
rect 1855 106 1884 152
rect 1744 93 1884 106
rect 1804 68 1884 93
rect 2004 152 2108 232
rect 2004 106 2033 152
rect 2079 106 2108 152
rect 2004 68 2108 106
rect 2228 68 2292 232
rect 2412 127 2500 232
rect 2412 81 2441 127
rect 2487 81 2500 127
rect 2412 68 2500 81
rect 2580 192 2668 232
rect 2580 146 2593 192
rect 2639 146 2668 192
rect 2580 68 2668 146
rect 2788 184 2892 232
rect 2788 138 2817 184
rect 2863 138 2892 184
rect 2788 68 2892 138
rect 3012 193 3100 232
rect 3012 147 3041 193
rect 3087 147 3100 193
rect 3012 68 3100 147
<< mvpdiff >>
rect 1816 698 1904 716
rect 1816 638 1829 698
rect 56 622 144 638
rect 56 576 69 622
rect 115 576 144 622
rect 56 561 144 576
rect 244 561 368 638
rect 468 625 628 638
rect 468 579 497 625
rect 543 579 628 625
rect 468 561 628 579
rect 548 526 628 561
rect 728 625 832 638
rect 728 579 757 625
rect 803 579 832 625
rect 728 526 832 579
rect 932 585 1036 638
rect 932 539 961 585
rect 1007 539 1036 585
rect 932 526 1036 539
rect 1136 625 1224 638
rect 1136 579 1165 625
rect 1211 579 1224 625
rect 1136 526 1224 579
rect 1347 585 1435 638
rect 1347 539 1360 585
rect 1406 539 1435 585
rect 1347 526 1435 539
rect 1535 526 1644 638
rect 1744 558 1829 638
rect 1875 558 1904 698
rect 1744 526 1904 558
rect 1816 472 1904 526
rect 2004 678 2123 716
rect 2004 632 2048 678
rect 2094 632 2123 678
rect 2004 472 2123 632
rect 2223 586 2327 716
rect 2223 540 2252 586
rect 2298 540 2327 586
rect 2223 472 2327 540
rect 2427 678 2515 716
rect 2427 632 2456 678
rect 2502 632 2515 678
rect 2427 472 2515 632
rect 2590 665 2678 716
rect 2590 525 2603 665
rect 2649 525 2678 665
rect 2590 472 2678 525
rect 2778 665 2902 716
rect 2778 619 2807 665
rect 2853 619 2902 665
rect 2778 472 2902 619
rect 3002 665 3090 716
rect 3002 525 3031 665
rect 3077 525 3090 665
rect 3002 472 3090 525
<< mvndiffc >>
rect 49 106 95 152
rect 273 106 319 152
rect 514 106 560 152
rect 757 106 803 152
rect 1165 106 1211 152
rect 1325 106 1371 152
rect 1549 106 1595 152
rect 1809 106 1855 152
rect 2033 106 2079 152
rect 2441 81 2487 127
rect 2593 146 2639 192
rect 2817 138 2863 184
rect 3041 147 3087 193
<< mvpdiffc >>
rect 69 576 115 622
rect 497 579 543 625
rect 757 579 803 625
rect 961 539 1007 585
rect 1165 579 1211 625
rect 1360 539 1406 585
rect 1829 558 1875 698
rect 2048 632 2094 678
rect 2252 540 2298 586
rect 2456 632 2502 678
rect 2603 525 2649 665
rect 2807 619 2853 665
rect 3031 525 3077 665
<< polysilicon >>
rect 144 638 244 682
rect 368 638 468 682
rect 628 638 728 682
rect 832 638 932 682
rect 1036 638 1136 682
rect 1435 638 1535 719
rect 1644 638 1744 719
rect 1904 716 2004 760
rect 2123 716 2223 760
rect 2327 716 2427 760
rect 2678 716 2778 760
rect 2902 716 3002 760
rect 144 528 244 561
rect 144 482 181 528
rect 227 482 244 528
rect 144 215 244 482
rect 368 303 468 561
rect 368 257 409 303
rect 455 257 468 303
rect 368 215 468 257
rect 628 399 728 526
rect 628 353 653 399
rect 699 353 728 399
rect 628 215 728 353
rect 124 165 244 215
rect 348 165 468 215
rect 608 165 728 215
rect 832 304 932 526
rect 832 258 861 304
rect 907 258 932 304
rect 832 215 932 258
rect 1036 413 1136 526
rect 1036 367 1062 413
rect 1108 367 1136 413
rect 1036 215 1136 367
rect 1435 482 1535 526
rect 1435 260 1520 482
rect 832 165 952 215
rect 1016 165 1136 215
rect 1400 245 1520 260
rect 1400 199 1426 245
rect 1472 199 1520 245
rect 1644 411 1744 526
rect 1644 365 1680 411
rect 1726 365 1744 411
rect 1644 215 1744 365
rect 1904 311 2004 472
rect 1904 276 1922 311
rect 1884 265 1922 276
rect 1968 265 2004 311
rect 2123 311 2223 472
rect 2123 276 2148 311
rect 1884 232 2004 265
rect 2108 265 2148 276
rect 2194 276 2223 311
rect 2327 428 2427 472
rect 2327 416 2412 428
rect 2327 370 2353 416
rect 2399 370 2412 416
rect 2327 276 2412 370
rect 2678 409 2778 472
rect 2678 363 2703 409
rect 2749 363 2778 409
rect 2678 357 2778 363
rect 2902 409 3002 472
rect 2902 363 2923 409
rect 2969 363 3002 409
rect 2902 357 3002 363
rect 2678 311 3002 357
rect 2678 288 2788 311
rect 2194 265 2228 276
rect 2108 232 2228 265
rect 2292 232 2412 276
rect 2668 232 2788 288
rect 2892 288 3002 311
rect 2892 232 3012 288
rect 1400 165 1520 199
rect 1624 165 1744 215
rect 124 49 244 93
rect 348 49 468 93
rect 608 49 728 93
rect 832 49 952 93
rect 1016 49 1136 93
rect 1400 49 1520 93
rect 1624 49 1744 93
rect 1884 24 2004 68
rect 2108 24 2228 68
rect 2292 24 2412 68
rect 2668 24 2788 68
rect 2892 24 3012 68
<< polycontact >>
rect 181 482 227 528
rect 409 257 455 303
rect 653 353 699 399
rect 861 258 907 304
rect 1062 367 1108 413
rect 1426 199 1472 245
rect 1680 365 1726 411
rect 1922 265 1968 311
rect 2148 265 2194 311
rect 2353 370 2399 416
rect 2703 363 2749 409
rect 2923 363 2969 409
<< metal1 >>
rect 0 724 3136 844
rect 69 622 115 638
rect 484 625 556 724
rect 1818 698 1886 724
rect 484 579 497 625
rect 543 579 556 625
rect 744 631 1211 678
rect 744 625 816 631
rect 744 579 757 625
rect 803 579 816 625
rect 1152 625 1211 631
rect 69 245 115 576
rect 950 539 961 585
rect 1007 539 1018 585
rect 1152 579 1165 625
rect 1152 568 1211 579
rect 1257 631 1613 678
rect 165 528 848 531
rect 165 482 181 528
rect 227 482 848 528
rect 165 477 848 482
rect 787 420 848 477
rect 950 513 1018 539
rect 1257 513 1303 631
rect 950 467 1303 513
rect 787 413 1143 420
rect 273 353 653 399
rect 699 353 714 399
rect 787 367 1062 413
rect 1108 367 1143 413
rect 787 363 1143 367
rect 273 245 330 353
rect 387 304 981 307
rect 387 303 861 304
rect 387 257 409 303
rect 455 258 861 303
rect 907 258 981 304
rect 455 257 981 258
rect 387 253 981 257
rect 69 198 330 245
rect 1257 245 1303 467
rect 1349 539 1360 585
rect 1406 539 1417 585
rect 1349 419 1417 539
rect 1567 511 1613 631
rect 1818 558 1829 698
rect 1875 558 1886 698
rect 2009 632 2048 678
rect 2094 632 2456 678
rect 2502 632 2515 678
rect 2603 665 2659 678
rect 1818 557 1886 558
rect 2223 540 2252 586
rect 2298 540 2515 586
rect 1567 494 2177 511
rect 1567 465 2399 494
rect 2131 448 2399 465
rect 1349 372 1606 419
rect 1538 276 1606 372
rect 1660 411 2085 419
rect 1660 365 1680 411
rect 1726 365 2085 411
rect 1660 363 2085 365
rect 2034 322 2085 363
rect 2353 416 2399 448
rect 2353 343 2399 370
rect 2469 409 2515 540
rect 2649 536 2659 665
rect 2807 665 2853 724
rect 2807 590 2853 619
rect 3031 665 3107 678
rect 2649 525 3031 536
rect 3077 525 3107 665
rect 2603 472 3107 525
rect 2469 363 2703 409
rect 2749 363 2923 409
rect 2969 363 2983 409
rect 2034 311 2215 322
rect 1903 276 1922 311
rect 1538 265 1922 276
rect 1968 265 1981 311
rect 1257 244 1426 245
rect 262 152 330 198
rect 1046 199 1426 244
rect 1472 199 1487 245
rect 1046 198 1487 199
rect 1538 230 1981 265
rect 2034 265 2148 311
rect 2194 265 2215 311
rect 2034 242 2215 265
rect 1046 152 1092 198
rect 1538 152 1606 230
rect 2469 219 2515 363
rect 3031 312 3107 472
rect 38 106 49 152
rect 95 106 106 152
rect 262 106 273 152
rect 319 106 330 152
rect 503 106 514 152
rect 560 106 571 152
rect 746 106 757 152
rect 803 106 1092 152
rect 1154 106 1165 152
rect 1211 106 1222 152
rect 38 60 106 106
rect 503 60 571 106
rect 1154 60 1222 106
rect 1314 106 1325 152
rect 1371 106 1382 152
rect 1538 106 1549 152
rect 1595 106 1606 152
rect 1809 152 1855 178
rect 2281 173 2515 219
rect 2593 248 3107 312
rect 2593 192 2662 248
rect 2281 153 2342 173
rect 2007 152 2342 153
rect 2007 106 2033 152
rect 2079 106 2342 152
rect 2639 146 2662 192
rect 1314 60 1382 106
rect 1809 60 1855 106
rect 2430 81 2441 127
rect 2487 81 2498 127
rect 2593 120 2662 146
rect 2817 184 2863 195
rect 2430 60 2498 81
rect 2817 60 2863 138
rect 3031 193 3107 248
rect 3031 147 3041 193
rect 3087 147 3107 193
rect 3031 120 3107 147
rect 0 -60 3136 60
<< labels >>
flabel metal1 s 1660 363 2085 419 0 FreeSans 400 0 0 0 A3
port 3 nsew default input
flabel metal1 s 0 724 3136 844 0 FreeSans 400 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 2817 178 2863 195 0 FreeSans 400 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel metal1 s 3031 536 3107 678 0 FreeSans 400 0 0 0 ZN
port 4 nsew default output
flabel metal1 s 387 253 981 307 0 FreeSans 400 0 0 0 A1
port 1 nsew default input
flabel metal1 s 165 477 848 531 0 FreeSans 400 0 0 0 A2
port 2 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 6 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 787 420 848 477 1 A2
port 2 nsew default input
rlabel metal1 s 787 363 1143 420 1 A2
port 2 nsew default input
rlabel metal1 s 2034 322 2085 363 1 A3
port 3 nsew default input
rlabel metal1 s 2034 242 2215 322 1 A3
port 3 nsew default input
rlabel metal1 s 2603 536 2659 678 1 ZN
port 4 nsew default output
rlabel metal1 s 2603 472 3107 536 1 ZN
port 4 nsew default output
rlabel metal1 s 3031 312 3107 472 1 ZN
port 4 nsew default output
rlabel metal1 s 2593 248 3107 312 1 ZN
port 4 nsew default output
rlabel metal1 s 3031 120 3107 248 1 ZN
port 4 nsew default output
rlabel metal1 s 2593 120 2662 248 1 ZN
port 4 nsew default output
rlabel metal1 s 2807 590 2853 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1818 590 1886 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 484 590 556 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1818 579 1886 590 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 484 579 556 590 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1818 557 1886 579 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2817 152 2863 178 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1809 152 1855 178 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2817 127 2863 152 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1809 127 1855 152 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1314 127 1382 152 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1154 127 1222 152 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 503 127 571 152 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 38 127 106 152 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2817 60 2863 127 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2430 60 2498 127 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1809 60 1855 127 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1314 60 1382 127 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1154 60 1222 127 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 503 60 571 127 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 38 60 106 127 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3136 60 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3136 784
string GDS_END 348236
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 341132
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
