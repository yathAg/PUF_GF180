magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 352 3558 870
<< pwell >>
rect -86 -86 3558 352
<< metal1 >>
rect 0 724 3472 844
rect 297 657 365 724
rect 1293 657 1361 724
rect 2349 635 2417 724
rect 186 240 681 320
rect 2679 532 2747 639
rect 2893 635 2961 724
rect 3108 532 3230 651
rect 3311 541 3379 724
rect 2679 485 3230 532
rect 3108 231 3230 485
rect 2679 185 3230 231
rect 317 60 385 127
rect 1333 60 1401 127
rect 2385 60 2431 139
rect 2679 135 2726 185
rect 3108 146 3230 185
rect 2904 60 2950 139
rect 3352 60 3398 139
rect 0 -60 3472 60
<< obsm1 >>
rect 49 481 117 621
rect 49 413 653 481
rect 49 180 95 413
rect 744 361 790 632
rect 877 575 1252 621
rect 744 293 1160 361
rect 1206 350 1252 575
rect 1780 564 1857 632
rect 1780 375 1826 564
rect 1944 493 1990 632
rect 1944 447 2338 493
rect 1206 304 1623 350
rect 1780 307 2216 375
rect 2274 352 2338 447
rect 49 134 117 180
rect 744 154 821 293
rect 1206 200 1252 304
rect 897 154 1252 200
rect 1780 143 1826 307
rect 2274 306 2938 352
rect 2274 211 2338 306
rect 1944 143 2338 211
<< labels >>
rlabel metal1 s 186 240 681 320 6 I
port 1 nsew default input
rlabel metal1 s 3108 146 3230 185 6 Z
port 2 nsew default output
rlabel metal1 s 2679 135 2726 185 6 Z
port 2 nsew default output
rlabel metal1 s 2679 185 3230 231 6 Z
port 2 nsew default output
rlabel metal1 s 3108 231 3230 485 6 Z
port 2 nsew default output
rlabel metal1 s 2679 485 3230 532 6 Z
port 2 nsew default output
rlabel metal1 s 3108 532 3230 651 6 Z
port 2 nsew default output
rlabel metal1 s 2679 532 2747 639 6 Z
port 2 nsew default output
rlabel metal1 s 3311 541 3379 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2893 635 2961 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2349 635 2417 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1293 657 1361 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 297 657 365 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 724 3472 844 6 VDD
port 3 nsew power bidirectional abutment
rlabel nwell s -86 352 3558 870 6 VNW
port 4 nsew power bidirectional
rlabel pwell s -86 -86 3558 352 6 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 0 -60 3472 60 8 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3352 60 3398 139 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2904 60 2950 139 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2385 60 2431 139 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1333 60 1401 127 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 317 60 385 127 6 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3472 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1122016
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1115372
<< end >>
