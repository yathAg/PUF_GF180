magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 377 3782 870
rect -86 352 227 377
rect 1799 352 3782 377
<< pwell >>
rect -86 -86 3782 352
<< mvnmos >>
rect 124 68 244 232
rect 392 93 512 257
rect 616 93 736 257
rect 840 93 960 257
rect 1064 93 1184 257
rect 1288 93 1408 257
rect 1512 93 1632 257
rect 1780 68 1900 232
rect 2004 68 2124 232
rect 2208 68 2328 232
rect 2432 68 2552 232
rect 2616 68 2736 232
rect 2840 68 2960 232
rect 3024 68 3144 232
rect 3248 68 3368 232
rect 3432 68 3552 232
<< mvpmos >>
rect 144 497 244 716
rect 412 497 512 716
rect 616 497 716 716
rect 860 497 960 716
rect 1064 497 1164 716
rect 1308 497 1408 716
rect 1512 497 1612 716
rect 1780 497 1880 716
rect 2024 519 2124 716
rect 2228 519 2328 716
rect 2432 519 2532 716
rect 2636 519 2736 716
rect 2840 519 2940 716
rect 3044 519 3144 716
rect 3248 519 3348 716
rect 3452 519 3552 716
<< mvndiff >>
rect 304 244 392 257
rect 304 232 317 244
rect 36 152 124 232
rect 36 106 49 152
rect 95 106 124 152
rect 36 68 124 106
rect 244 198 317 232
rect 363 198 392 244
rect 244 93 392 198
rect 512 152 616 257
rect 512 106 541 152
rect 587 106 616 152
rect 512 93 616 106
rect 736 244 840 257
rect 736 198 765 244
rect 811 198 840 244
rect 736 93 840 198
rect 960 152 1064 257
rect 960 106 989 152
rect 1035 106 1064 152
rect 960 93 1064 106
rect 1184 244 1288 257
rect 1184 198 1213 244
rect 1259 198 1288 244
rect 1184 93 1288 198
rect 1408 152 1512 257
rect 1408 106 1437 152
rect 1483 106 1512 152
rect 1408 93 1512 106
rect 1632 244 1720 257
rect 1632 198 1661 244
rect 1707 232 1720 244
rect 1707 198 1780 232
rect 1632 93 1780 198
rect 244 68 324 93
rect 1700 68 1780 93
rect 1900 152 2004 232
rect 1900 106 1929 152
rect 1975 106 2004 152
rect 1900 68 2004 106
rect 2124 68 2208 232
rect 2328 127 2432 232
rect 2328 81 2357 127
rect 2403 81 2432 127
rect 2328 68 2432 81
rect 2552 68 2616 232
rect 2736 152 2840 232
rect 2736 106 2765 152
rect 2811 106 2840 152
rect 2736 68 2840 106
rect 2960 68 3024 232
rect 3144 127 3248 232
rect 3144 81 3173 127
rect 3219 81 3248 127
rect 3144 68 3248 81
rect 3368 68 3432 232
rect 3552 219 3640 232
rect 3552 173 3581 219
rect 3627 173 3640 219
rect 3552 68 3640 173
<< mvpdiff >>
rect 56 665 144 716
rect 56 525 69 665
rect 115 525 144 665
rect 56 497 144 525
rect 244 497 412 716
rect 512 665 616 716
rect 512 525 541 665
rect 587 525 616 665
rect 512 497 616 525
rect 716 497 860 716
rect 960 703 1064 716
rect 960 657 989 703
rect 1035 657 1064 703
rect 960 497 1064 657
rect 1164 497 1308 716
rect 1408 639 1512 716
rect 1408 593 1437 639
rect 1483 593 1512 639
rect 1408 497 1512 593
rect 1612 497 1780 716
rect 1880 703 2024 716
rect 1880 657 1929 703
rect 1975 657 2024 703
rect 1880 519 2024 657
rect 2124 639 2228 716
rect 2124 593 2153 639
rect 2199 593 2228 639
rect 2124 519 2228 593
rect 2328 703 2432 716
rect 2328 657 2357 703
rect 2403 657 2432 703
rect 2328 519 2432 657
rect 2532 639 2636 716
rect 2532 593 2561 639
rect 2607 593 2636 639
rect 2532 519 2636 593
rect 2736 703 2840 716
rect 2736 657 2765 703
rect 2811 657 2840 703
rect 2736 519 2840 657
rect 2940 639 3044 716
rect 2940 593 2969 639
rect 3015 593 3044 639
rect 2940 519 3044 593
rect 3144 703 3248 716
rect 3144 657 3173 703
rect 3219 657 3248 703
rect 3144 519 3248 657
rect 3348 639 3452 716
rect 3348 593 3377 639
rect 3423 593 3452 639
rect 3348 519 3452 593
rect 3552 672 3640 716
rect 3552 532 3581 672
rect 3627 532 3640 672
rect 3552 519 3640 532
rect 1880 497 1960 519
<< mvndiffc >>
rect 49 106 95 152
rect 317 198 363 244
rect 541 106 587 152
rect 765 198 811 244
rect 989 106 1035 152
rect 1213 198 1259 244
rect 1437 106 1483 152
rect 1661 198 1707 244
rect 1929 106 1975 152
rect 2357 81 2403 127
rect 2765 106 2811 152
rect 3173 81 3219 127
rect 3581 173 3627 219
<< mvpdiffc >>
rect 69 525 115 665
rect 541 525 587 665
rect 989 657 1035 703
rect 1437 593 1483 639
rect 1929 657 1975 703
rect 2153 593 2199 639
rect 2357 657 2403 703
rect 2561 593 2607 639
rect 2765 657 2811 703
rect 2969 593 3015 639
rect 3173 657 3219 703
rect 3377 593 3423 639
rect 3581 532 3627 672
<< polysilicon >>
rect 144 716 244 760
rect 412 716 512 760
rect 616 716 716 760
rect 860 716 960 760
rect 1064 716 1164 760
rect 1308 716 1408 760
rect 1512 716 1612 760
rect 1780 716 1880 760
rect 2024 716 2124 760
rect 2228 716 2328 760
rect 2432 716 2532 760
rect 2636 716 2736 760
rect 2840 716 2940 760
rect 3044 716 3144 760
rect 3248 716 3348 760
rect 3452 716 3552 760
rect 144 428 244 497
rect 144 401 171 428
rect 124 382 171 401
rect 217 382 244 428
rect 412 401 512 497
rect 616 401 716 497
rect 860 428 960 497
rect 860 401 887 428
rect 124 232 244 382
rect 392 344 736 401
rect 392 336 512 344
rect 392 290 429 336
rect 475 290 512 336
rect 392 257 512 290
rect 616 336 736 344
rect 616 290 653 336
rect 699 290 736 336
rect 616 257 736 290
rect 840 382 887 401
rect 933 401 960 428
rect 1064 428 1164 497
rect 1064 401 1091 428
rect 933 382 1091 401
rect 1137 401 1164 428
rect 1308 413 1408 497
rect 1308 401 1335 413
rect 1137 382 1184 401
rect 840 344 1184 382
rect 840 257 960 344
rect 1064 257 1184 344
rect 1288 367 1335 401
rect 1381 401 1408 413
rect 1512 413 1612 497
rect 1512 401 1539 413
rect 1381 367 1539 401
rect 1585 401 1612 413
rect 1780 413 1880 497
rect 1585 367 1632 401
rect 1288 344 1632 367
rect 1288 257 1408 344
rect 1512 257 1632 344
rect 1780 367 1809 413
rect 1855 401 1880 413
rect 2024 413 2124 519
rect 2024 401 2050 413
rect 1855 367 1900 401
rect 1780 232 1900 367
rect 2004 367 2050 401
rect 2096 367 2124 413
rect 2228 413 2328 519
rect 2228 401 2255 413
rect 2004 232 2124 367
rect 2208 367 2255 401
rect 2301 401 2328 413
rect 2432 413 2532 519
rect 2432 401 2459 413
rect 2301 367 2459 401
rect 2505 401 2532 413
rect 2636 401 2736 519
rect 2840 401 2940 519
rect 3044 413 3144 519
rect 3044 401 3071 413
rect 2505 367 2552 401
rect 2208 344 2552 367
rect 2208 232 2328 344
rect 2432 232 2552 344
rect 2616 344 2960 401
rect 2616 311 2736 344
rect 2616 265 2653 311
rect 2699 265 2736 311
rect 2616 232 2736 265
rect 2840 311 2960 344
rect 2840 265 2877 311
rect 2923 265 2960 311
rect 2840 232 2960 265
rect 3024 367 3071 401
rect 3117 401 3144 413
rect 3248 413 3348 519
rect 3248 401 3275 413
rect 3117 367 3275 401
rect 3321 401 3348 413
rect 3452 401 3552 519
rect 3321 367 3368 401
rect 3024 344 3368 367
rect 3024 232 3144 344
rect 3248 232 3368 344
rect 3432 311 3552 401
rect 3432 265 3465 311
rect 3511 265 3552 311
rect 3432 232 3552 265
rect 124 24 244 68
rect 392 24 512 93
rect 616 24 736 93
rect 840 24 960 93
rect 1064 24 1184 93
rect 1288 24 1408 93
rect 1512 24 1632 93
rect 1780 24 1900 68
rect 2004 24 2124 68
rect 2208 24 2328 68
rect 2432 24 2552 68
rect 2616 24 2736 68
rect 2840 24 2960 68
rect 3024 24 3144 68
rect 3248 24 3368 68
rect 3432 24 3552 68
<< polycontact >>
rect 171 382 217 428
rect 429 290 475 336
rect 653 290 699 336
rect 887 382 933 428
rect 1091 382 1137 428
rect 1335 367 1381 413
rect 1539 367 1585 413
rect 1809 367 1855 413
rect 2050 367 2096 413
rect 2255 367 2301 413
rect 2459 367 2505 413
rect 2653 265 2699 311
rect 2877 265 2923 311
rect 3071 367 3117 413
rect 3275 367 3321 413
rect 3465 265 3511 311
<< metal1 >>
rect 0 724 3696 844
rect 69 665 115 724
rect 978 703 1046 724
rect 69 506 115 525
rect 530 525 541 665
rect 587 648 598 665
rect 978 657 989 703
rect 1035 657 1046 703
rect 1918 703 1986 724
rect 1918 657 1929 703
rect 1975 657 1986 703
rect 2346 703 2414 724
rect 2346 657 2357 703
rect 2403 657 2414 703
rect 2754 703 2822 724
rect 2754 657 2765 703
rect 2811 657 2822 703
rect 3162 703 3230 724
rect 3162 657 3173 703
rect 3219 657 3230 703
rect 3581 672 3627 724
rect 587 605 928 648
rect 1095 639 1868 648
rect 1095 605 1437 639
rect 587 593 1437 605
rect 1483 605 1868 639
rect 2035 639 2296 648
rect 2035 605 2153 639
rect 1483 593 2153 605
rect 2199 611 2296 639
rect 2464 639 2704 648
rect 2464 611 2561 639
rect 2199 593 2561 611
rect 2607 611 2704 639
rect 2872 639 3112 648
rect 2872 611 2969 639
rect 2607 593 2969 611
rect 3015 611 3112 639
rect 3280 639 3490 648
rect 3280 611 3377 639
rect 3015 593 3377 611
rect 3423 593 3490 639
rect 587 584 3490 593
rect 587 525 598 584
rect 878 559 1145 584
rect 1818 559 3490 584
rect 530 495 598 525
rect 1191 472 1776 536
rect 1191 428 1241 472
rect 124 382 171 428
rect 217 382 887 428
rect 933 382 1091 428
rect 1137 382 1241 428
rect 1708 424 1776 472
rect 1308 413 1662 424
rect 1308 367 1335 413
rect 1381 367 1539 413
rect 1585 367 1662 413
rect 1308 354 1662 367
rect 1708 413 1882 424
rect 1708 367 1809 413
rect 1855 367 1882 413
rect 1708 354 1882 367
rect 1308 336 1358 354
rect 392 290 429 336
rect 475 290 653 336
rect 699 290 1358 336
rect 1928 244 1992 559
rect 3581 519 3627 532
rect 2040 413 2104 485
rect 2040 367 2050 413
rect 2096 367 2104 413
rect 2040 311 2104 367
rect 2150 413 3368 424
rect 2150 367 2255 413
rect 2301 367 2459 413
rect 2505 367 3071 413
rect 3117 367 3275 413
rect 3321 367 3368 413
rect 2150 360 3368 367
rect 2040 265 2653 311
rect 2699 265 2877 311
rect 2923 265 3465 311
rect 3511 265 3552 311
rect 2586 244 3016 265
rect 304 198 317 244
rect 363 198 765 244
rect 811 198 1213 244
rect 1259 198 1661 244
rect 1707 198 1992 244
rect 2131 173 2510 219
rect 2131 152 2177 173
rect 36 106 49 152
rect 95 106 541 152
rect 587 106 989 152
rect 1035 106 1437 152
rect 1483 106 1929 152
rect 1975 106 2177 152
rect 2464 152 2510 173
rect 3066 173 3581 219
rect 3627 173 3640 219
rect 3066 152 3112 173
rect 2346 81 2357 127
rect 2403 81 2414 127
rect 2464 106 2765 152
rect 2811 106 3112 152
rect 2346 60 2414 81
rect 3162 81 3173 127
rect 3219 81 3230 127
rect 3162 60 3230 81
rect 0 -60 3696 60
<< labels >>
flabel metal1 s 2040 311 2104 485 0 FreeSans 400 0 0 0 B
port 3 nsew default input
flabel metal1 s 2150 360 3368 424 0 FreeSans 400 0 0 0 C
port 4 nsew default input
flabel metal1 s 0 724 3696 844 0 FreeSans 400 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 3162 60 3230 127 0 FreeSans 400 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel metal1 s 530 648 598 665 0 FreeSans 400 0 0 0 ZN
port 5 nsew default output
flabel metal1 s 1308 354 1662 424 0 FreeSans 400 0 0 0 A1
port 1 nsew default input
flabel metal1 s 1191 472 1776 536 0 FreeSans 400 0 0 0 A2
port 2 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 7 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 8 nsew ground bidirectional
rlabel metal1 s 1308 336 1358 354 1 A1
port 1 nsew default input
rlabel metal1 s 392 290 1358 336 1 A1
port 1 nsew default input
rlabel metal1 s 1708 428 1776 472 1 A2
port 2 nsew default input
rlabel metal1 s 1191 428 1241 472 1 A2
port 2 nsew default input
rlabel metal1 s 1708 424 1776 428 1 A2
port 2 nsew default input
rlabel metal1 s 124 424 1241 428 1 A2
port 2 nsew default input
rlabel metal1 s 1708 382 1882 424 1 A2
port 2 nsew default input
rlabel metal1 s 124 382 1241 424 1 A2
port 2 nsew default input
rlabel metal1 s 1708 354 1882 382 1 A2
port 2 nsew default input
rlabel metal1 s 2040 265 3552 311 1 B
port 3 nsew default input
rlabel metal1 s 2586 244 3016 265 1 B
port 3 nsew default input
rlabel metal1 s 3280 611 3490 648 1 ZN
port 5 nsew default output
rlabel metal1 s 2872 611 3112 648 1 ZN
port 5 nsew default output
rlabel metal1 s 2464 611 2704 648 1 ZN
port 5 nsew default output
rlabel metal1 s 2035 611 2296 648 1 ZN
port 5 nsew default output
rlabel metal1 s 1095 611 1868 648 1 ZN
port 5 nsew default output
rlabel metal1 s 530 611 928 648 1 ZN
port 5 nsew default output
rlabel metal1 s 2035 605 3490 611 1 ZN
port 5 nsew default output
rlabel metal1 s 1095 605 1868 611 1 ZN
port 5 nsew default output
rlabel metal1 s 530 605 928 611 1 ZN
port 5 nsew default output
rlabel metal1 s 530 584 3490 605 1 ZN
port 5 nsew default output
rlabel metal1 s 1818 559 3490 584 1 ZN
port 5 nsew default output
rlabel metal1 s 878 559 1145 584 1 ZN
port 5 nsew default output
rlabel metal1 s 530 559 598 584 1 ZN
port 5 nsew default output
rlabel metal1 s 1928 495 1992 559 1 ZN
port 5 nsew default output
rlabel metal1 s 530 495 598 559 1 ZN
port 5 nsew default output
rlabel metal1 s 1928 244 1992 495 1 ZN
port 5 nsew default output
rlabel metal1 s 304 198 1992 244 1 ZN
port 5 nsew default output
rlabel metal1 s 3581 657 3627 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3162 657 3230 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2754 657 2822 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2346 657 2414 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1918 657 1986 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 978 657 1046 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 69 657 115 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3581 519 3627 657 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 69 519 115 657 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 69 506 115 519 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2346 60 2414 127 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3696 60 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3696 784
string GDS_END 104678
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 97608
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
