magic
tech gf180mcuB
timestamp 1698431365
<< properties >>
string GDS_END 10712178
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 10710510
<< end >>
