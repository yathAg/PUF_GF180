magic
tech gf180mcuD
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 352 2550 870
<< pwell >>
rect -86 -86 2550 352
<< mvnmos >>
rect 179 68 299 140
rect 403 68 523 140
rect 571 68 691 140
rect 1027 68 1147 141
rect 1195 68 1315 141
rect 1525 68 1645 232
rect 1749 68 1869 232
rect 1973 68 2093 232
rect 2197 68 2317 232
<< mvpmos >>
rect 179 644 279 716
rect 403 644 503 716
rect 571 644 671 716
rect 1027 622 1127 694
rect 1195 622 1295 694
rect 1555 472 1655 716
rect 1759 472 1859 716
rect 1963 472 2063 716
rect 2197 472 2297 716
<< mvndiff >>
rect 47 180 119 193
rect 47 134 60 180
rect 106 140 119 180
rect 751 200 823 213
rect 751 154 764 200
rect 810 154 823 200
rect 751 140 823 154
rect 106 134 179 140
rect 47 68 179 134
rect 299 127 403 140
rect 299 81 328 127
rect 374 81 403 127
rect 299 68 403 81
rect 523 68 571 140
rect 691 68 823 140
rect 895 200 967 213
rect 895 154 908 200
rect 954 154 967 200
rect 895 141 967 154
rect 1445 141 1525 232
rect 895 68 1027 141
rect 1147 68 1195 141
rect 1315 127 1525 141
rect 1315 81 1344 127
rect 1390 81 1525 127
rect 1315 68 1525 81
rect 1645 192 1749 232
rect 1645 146 1674 192
rect 1720 146 1749 192
rect 1645 68 1749 146
rect 1869 127 1973 232
rect 1869 81 1898 127
rect 1944 81 1973 127
rect 1869 68 1973 81
rect 2093 192 2197 232
rect 2093 146 2122 192
rect 2168 146 2197 192
rect 2093 68 2197 146
rect 2317 184 2405 232
rect 2317 138 2346 184
rect 2392 138 2405 184
rect 2317 68 2405 138
<< mvpdiff >>
rect 47 644 179 716
rect 279 703 403 716
rect 279 657 308 703
rect 354 657 403 703
rect 279 644 403 657
rect 503 644 571 716
rect 671 644 803 716
rect 1445 694 1555 716
rect 47 621 119 644
rect 47 575 60 621
rect 106 575 119 621
rect 47 562 119 575
rect 731 621 803 644
rect 731 575 744 621
rect 790 575 803 621
rect 731 562 803 575
rect 895 622 1027 694
rect 1127 622 1195 694
rect 1295 681 1555 694
rect 1295 635 1324 681
rect 1370 665 1555 681
rect 1370 635 1480 665
rect 1295 622 1480 635
rect 895 621 967 622
rect 895 575 908 621
rect 954 575 967 621
rect 895 562 967 575
rect 1445 525 1480 622
rect 1526 525 1555 665
rect 1445 472 1555 525
rect 1655 665 1759 716
rect 1655 525 1684 665
rect 1730 525 1759 665
rect 1655 472 1759 525
rect 1859 665 1963 716
rect 1859 525 1888 665
rect 1934 525 1963 665
rect 1859 472 1963 525
rect 2063 665 2197 716
rect 2063 525 2122 665
rect 2168 525 2197 665
rect 2063 472 2197 525
rect 2297 665 2385 716
rect 2297 525 2326 665
rect 2372 525 2385 665
rect 2297 472 2385 525
<< mvndiffc >>
rect 60 134 106 180
rect 764 154 810 200
rect 328 81 374 127
rect 908 154 954 200
rect 1344 81 1390 127
rect 1674 146 1720 192
rect 1898 81 1944 127
rect 2122 146 2168 192
rect 2346 138 2392 184
<< mvpdiffc >>
rect 308 657 354 703
rect 60 575 106 621
rect 744 575 790 621
rect 1324 635 1370 681
rect 908 575 954 621
rect 1480 525 1526 665
rect 1684 525 1730 665
rect 1888 525 1934 665
rect 2122 525 2168 665
rect 2326 525 2372 665
<< polysilicon >>
rect 179 716 279 760
rect 403 716 503 760
rect 571 716 671 760
rect 1027 694 1127 738
rect 1195 694 1295 738
rect 1555 716 1655 760
rect 1759 716 1859 760
rect 1963 716 2063 760
rect 2197 716 2297 760
rect 179 303 279 644
rect 179 257 192 303
rect 238 257 279 303
rect 179 184 279 257
rect 403 483 503 644
rect 571 483 671 644
rect 403 470 671 483
rect 403 424 416 470
rect 462 424 596 470
rect 642 424 671 470
rect 403 411 671 424
rect 403 184 503 411
rect 571 184 671 411
rect 1027 399 1127 622
rect 1195 399 1295 622
rect 1027 382 1295 399
rect 1555 384 1655 472
rect 1759 384 1859 472
rect 1963 384 2063 472
rect 2197 384 2297 472
rect 1027 336 1040 382
rect 1086 344 1295 382
rect 1086 336 1127 344
rect 1027 251 1127 336
rect 1195 251 1295 344
rect 1525 371 2317 384
rect 1525 325 1538 371
rect 2054 325 2317 371
rect 1525 312 2317 325
rect 179 140 299 184
rect 403 140 523 184
rect 571 140 691 184
rect 1027 141 1147 251
rect 1195 141 1315 251
rect 1525 232 1645 312
rect 1749 232 1869 312
rect 1973 232 2093 312
rect 2197 232 2317 312
rect 179 24 299 68
rect 403 24 523 68
rect 571 24 691 68
rect 1027 24 1147 68
rect 1195 24 1315 68
rect 1525 24 1645 68
rect 1749 24 1869 68
rect 1973 24 2093 68
rect 2197 24 2317 68
<< polycontact >>
rect 192 257 238 303
rect 416 424 462 470
rect 596 424 642 470
rect 1040 336 1086 382
rect 1538 325 2054 371
<< metal1 >>
rect 0 724 2464 844
rect 297 703 365 724
rect 297 657 308 703
rect 354 657 365 703
rect 1313 681 1537 724
rect 1313 635 1324 681
rect 1370 665 1537 681
rect 1370 635 1480 665
rect 744 621 790 632
rect 49 575 60 621
rect 106 575 117 621
rect 49 481 117 575
rect 49 470 653 481
rect 49 424 416 470
rect 462 424 596 470
rect 642 424 653 470
rect 49 413 653 424
rect 49 180 95 413
rect 744 382 790 575
rect 908 621 954 632
rect 908 493 954 575
rect 1471 525 1480 635
rect 1526 525 1537 665
rect 1471 506 1537 525
rect 1684 665 1730 676
rect 908 447 1231 493
rect 744 336 1040 382
rect 1086 336 1097 382
rect 1167 371 1231 447
rect 1684 468 1730 525
rect 1888 665 1934 724
rect 1888 514 1934 525
rect 2122 665 2236 676
rect 2168 525 2236 665
rect 2122 468 2236 525
rect 2326 665 2372 724
rect 2326 506 2372 525
rect 1684 421 2236 468
rect 186 303 672 320
rect 186 257 192 303
rect 238 257 672 303
rect 186 240 672 257
rect 744 200 821 336
rect 1167 325 1538 371
rect 2054 325 2072 371
rect 1167 211 1231 325
rect 2122 243 2236 421
rect 49 134 60 180
rect 106 134 117 180
rect 744 154 764 200
rect 810 154 821 200
rect 908 200 1231 211
rect 954 154 1231 200
rect 908 143 1231 154
rect 1674 192 2236 243
rect 1344 127 1390 138
rect 317 81 328 127
rect 374 81 385 127
rect 317 60 385 81
rect 1674 106 1720 146
rect 2168 146 2236 192
rect 1344 60 1390 81
rect 1887 81 1898 127
rect 1944 81 1955 127
rect 2122 110 2236 146
rect 2346 184 2392 223
rect 1887 60 1955 81
rect 2346 60 2392 138
rect 0 -60 2464 60
<< labels >>
flabel metal1 s 2346 138 2392 223 0 FreeSans 400 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel metal1 s 2122 468 2236 676 0 FreeSans 400 0 0 0 Z
port 2 nsew default output
flabel metal1 s 186 240 672 320 0 FreeSans 400 0 0 0 I
port 1 nsew default input
flabel metal1 s 0 724 2464 844 0 FreeSans 400 0 0 0 VDD
port 3 nsew power bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 4 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 1684 468 1730 676 1 Z
port 2 nsew default output
rlabel metal1 s 1684 421 2236 468 1 Z
port 2 nsew default output
rlabel metal1 s 2122 243 2236 421 1 Z
port 2 nsew default output
rlabel metal1 s 1674 192 2236 243 1 Z
port 2 nsew default output
rlabel metal1 s 2122 110 2236 192 1 Z
port 2 nsew default output
rlabel metal1 s 1674 110 1720 192 1 Z
port 2 nsew default output
rlabel metal1 s 1674 106 1720 110 1 Z
port 2 nsew default output
rlabel metal1 s 2326 657 2372 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1888 657 1934 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1313 657 1537 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 297 657 365 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2326 635 2372 657 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1888 635 1934 657 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1313 635 1537 657 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2326 514 2372 635 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1888 514 1934 635 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1471 514 1537 635 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2326 506 2372 514 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1471 506 1537 514 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2346 127 2392 138 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1344 127 1390 138 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2346 60 2392 127 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1887 60 1955 127 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1344 60 1390 127 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 317 60 385 127 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 2464 60 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2464 784
string GDS_END 1104100
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1098704
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
