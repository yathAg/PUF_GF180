magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< metal1 >>
rect 742 2136 1686 2148
rect 742 2084 754 2136
rect 806 2084 878 2136
rect 930 2084 1002 2136
rect 1054 2084 1126 2136
rect 1178 2084 1250 2136
rect 1302 2084 1374 2136
rect 1426 2084 1498 2136
rect 1550 2084 1622 2136
rect 1674 2084 1686 2136
rect 742 2012 1686 2084
rect 742 1960 754 2012
rect 806 1960 878 2012
rect 930 1960 1002 2012
rect 1054 1960 1126 2012
rect 1178 1960 1250 2012
rect 1302 1960 1374 2012
rect 1426 1960 1498 2012
rect 1550 1960 1622 2012
rect 1674 1960 1686 2012
rect 742 1888 1686 1960
rect 742 1836 754 1888
rect 806 1836 878 1888
rect 930 1836 1002 1888
rect 1054 1836 1126 1888
rect 1178 1836 1250 1888
rect 1302 1836 1374 1888
rect 1426 1836 1498 1888
rect 1550 1836 1622 1888
rect 1674 1836 1686 1888
rect 742 1824 1686 1836
<< via1 >>
rect 754 2084 806 2136
rect 878 2084 930 2136
rect 1002 2084 1054 2136
rect 1126 2084 1178 2136
rect 1250 2084 1302 2136
rect 1374 2084 1426 2136
rect 1498 2084 1550 2136
rect 1622 2084 1674 2136
rect 754 1960 806 2012
rect 878 1960 930 2012
rect 1002 1960 1054 2012
rect 1126 1960 1178 2012
rect 1250 1960 1302 2012
rect 1374 1960 1426 2012
rect 1498 1960 1550 2012
rect 1622 1960 1674 2012
rect 754 1836 806 1888
rect 878 1836 930 1888
rect 1002 1836 1054 1888
rect 1126 1836 1178 1888
rect 1250 1836 1302 1888
rect 1374 1836 1426 1888
rect 1498 1836 1550 1888
rect 1622 1836 1674 1888
<< metal2 >>
rect 742 2138 1686 2148
rect 742 2082 752 2138
rect 808 2082 876 2138
rect 932 2082 1000 2138
rect 1056 2082 1124 2138
rect 1180 2082 1248 2138
rect 1304 2082 1372 2138
rect 1428 2082 1496 2138
rect 1552 2082 1620 2138
rect 1676 2082 1686 2138
rect 742 2014 1686 2082
rect 742 1958 752 2014
rect 808 1958 876 2014
rect 932 1958 1000 2014
rect 1056 1958 1124 2014
rect 1180 1958 1248 2014
rect 1304 1958 1372 2014
rect 1428 1958 1496 2014
rect 1552 1958 1620 2014
rect 1676 1958 1686 2014
rect 742 1890 1686 1958
rect 742 1834 752 1890
rect 808 1834 876 1890
rect 932 1834 1000 1890
rect 1056 1834 1124 1890
rect 1180 1834 1248 1890
rect 1304 1834 1372 1890
rect 1428 1834 1496 1890
rect 1552 1834 1620 1890
rect 1676 1834 1686 1890
rect 742 1824 1686 1834
<< via2 >>
rect 752 2136 808 2138
rect 752 2084 754 2136
rect 754 2084 806 2136
rect 806 2084 808 2136
rect 752 2082 808 2084
rect 876 2136 932 2138
rect 876 2084 878 2136
rect 878 2084 930 2136
rect 930 2084 932 2136
rect 876 2082 932 2084
rect 1000 2136 1056 2138
rect 1000 2084 1002 2136
rect 1002 2084 1054 2136
rect 1054 2084 1056 2136
rect 1000 2082 1056 2084
rect 1124 2136 1180 2138
rect 1124 2084 1126 2136
rect 1126 2084 1178 2136
rect 1178 2084 1180 2136
rect 1124 2082 1180 2084
rect 1248 2136 1304 2138
rect 1248 2084 1250 2136
rect 1250 2084 1302 2136
rect 1302 2084 1304 2136
rect 1248 2082 1304 2084
rect 1372 2136 1428 2138
rect 1372 2084 1374 2136
rect 1374 2084 1426 2136
rect 1426 2084 1428 2136
rect 1372 2082 1428 2084
rect 1496 2136 1552 2138
rect 1496 2084 1498 2136
rect 1498 2084 1550 2136
rect 1550 2084 1552 2136
rect 1496 2082 1552 2084
rect 1620 2136 1676 2138
rect 1620 2084 1622 2136
rect 1622 2084 1674 2136
rect 1674 2084 1676 2136
rect 1620 2082 1676 2084
rect 752 2012 808 2014
rect 752 1960 754 2012
rect 754 1960 806 2012
rect 806 1960 808 2012
rect 752 1958 808 1960
rect 876 2012 932 2014
rect 876 1960 878 2012
rect 878 1960 930 2012
rect 930 1960 932 2012
rect 876 1958 932 1960
rect 1000 2012 1056 2014
rect 1000 1960 1002 2012
rect 1002 1960 1054 2012
rect 1054 1960 1056 2012
rect 1000 1958 1056 1960
rect 1124 2012 1180 2014
rect 1124 1960 1126 2012
rect 1126 1960 1178 2012
rect 1178 1960 1180 2012
rect 1124 1958 1180 1960
rect 1248 2012 1304 2014
rect 1248 1960 1250 2012
rect 1250 1960 1302 2012
rect 1302 1960 1304 2012
rect 1248 1958 1304 1960
rect 1372 2012 1428 2014
rect 1372 1960 1374 2012
rect 1374 1960 1426 2012
rect 1426 1960 1428 2012
rect 1372 1958 1428 1960
rect 1496 2012 1552 2014
rect 1496 1960 1498 2012
rect 1498 1960 1550 2012
rect 1550 1960 1552 2012
rect 1496 1958 1552 1960
rect 1620 2012 1676 2014
rect 1620 1960 1622 2012
rect 1622 1960 1674 2012
rect 1674 1960 1676 2012
rect 1620 1958 1676 1960
rect 752 1888 808 1890
rect 752 1836 754 1888
rect 754 1836 806 1888
rect 806 1836 808 1888
rect 752 1834 808 1836
rect 876 1888 932 1890
rect 876 1836 878 1888
rect 878 1836 930 1888
rect 930 1836 932 1888
rect 876 1834 932 1836
rect 1000 1888 1056 1890
rect 1000 1836 1002 1888
rect 1002 1836 1054 1888
rect 1054 1836 1056 1888
rect 1000 1834 1056 1836
rect 1124 1888 1180 1890
rect 1124 1836 1126 1888
rect 1126 1836 1178 1888
rect 1178 1836 1180 1888
rect 1124 1834 1180 1836
rect 1248 1888 1304 1890
rect 1248 1836 1250 1888
rect 1250 1836 1302 1888
rect 1302 1836 1304 1888
rect 1248 1834 1304 1836
rect 1372 1888 1428 1890
rect 1372 1836 1374 1888
rect 1374 1836 1426 1888
rect 1426 1836 1428 1888
rect 1372 1834 1428 1836
rect 1496 1888 1552 1890
rect 1496 1836 1498 1888
rect 1498 1836 1550 1888
rect 1550 1836 1552 1888
rect 1496 1834 1552 1836
rect 1620 1888 1676 1890
rect 1620 1836 1622 1888
rect 1622 1836 1674 1888
rect 1674 1836 1676 1888
rect 1620 1834 1676 1836
<< metal3 >>
rect 714 2138 1714 2430
rect 714 2082 752 2138
rect 808 2082 876 2138
rect 932 2082 1000 2138
rect 1056 2082 1124 2138
rect 1180 2082 1248 2138
rect 1304 2082 1372 2138
rect 1428 2082 1496 2138
rect 1552 2082 1620 2138
rect 1676 2082 1714 2138
rect 714 2014 1714 2082
rect 714 1958 752 2014
rect 808 1958 876 2014
rect 932 1958 1000 2014
rect 1056 1958 1124 2014
rect 1180 1958 1248 2014
rect 1304 1958 1372 2014
rect 1428 1958 1496 2014
rect 1552 1958 1620 2014
rect 1676 1958 1714 2014
rect 714 1890 1714 1958
rect 714 1834 752 1890
rect 808 1834 876 1890
rect 932 1834 1000 1890
rect 1056 1834 1124 1890
rect 1180 1834 1248 1890
rect 1304 1834 1372 1890
rect 1428 1834 1496 1890
rect 1552 1834 1620 1890
rect 1676 1834 1714 1890
rect 714 1822 1714 1834
use M2_M14310590878179_256x8m81  M2_M14310590878179_256x8m81_0
timestamp 1698431365
transform 1 0 1214 0 1 1986
box 0 0 1 1
use M3_M24310590878178_256x8m81  M3_M24310590878178_256x8m81_0
timestamp 1698431365
transform 1 0 1214 0 1 1986
box 0 0 1 1
<< properties >>
string GDS_END 2396058
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 2395886
<< end >>
