magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 377 2662 870
rect -86 352 689 377
rect 1084 352 2662 377
<< pwell >>
rect 689 352 1084 377
rect -86 -86 2662 352
<< mvnmos >>
rect 135 68 255 232
rect 359 68 479 232
rect 583 68 703 232
rect 1070 68 1190 232
rect 1330 68 1450 176
rect 1554 68 1674 176
rect 1856 68 1976 232
rect 2080 68 2200 232
rect 2304 68 2424 232
<< mvpmos >>
rect 184 497 284 716
rect 388 497 488 716
rect 592 497 692 716
rect 1080 497 1180 716
rect 1320 515 1420 716
rect 1524 515 1624 716
rect 1764 480 1864 716
rect 1968 480 2068 716
rect 2172 480 2272 716
<< mvndiff >>
rect 763 244 835 257
rect 763 232 776 244
rect 47 192 135 232
rect 47 146 60 192
rect 106 146 135 192
rect 47 68 135 146
rect 255 139 359 232
rect 255 93 284 139
rect 330 93 359 139
rect 255 68 359 93
rect 479 166 583 232
rect 479 120 508 166
rect 554 120 583 166
rect 479 68 583 120
rect 703 198 776 232
rect 822 198 835 244
rect 703 68 835 198
rect 938 244 1010 257
rect 938 198 951 244
rect 997 232 1010 244
rect 997 198 1070 232
rect 938 68 1070 198
rect 1190 176 1270 232
rect 1776 176 1856 232
rect 1190 127 1330 176
rect 1190 81 1237 127
rect 1283 81 1330 127
rect 1190 68 1330 81
rect 1450 163 1554 176
rect 1450 117 1479 163
rect 1525 117 1554 163
rect 1450 68 1554 117
rect 1674 141 1856 176
rect 1674 95 1745 141
rect 1791 95 1856 141
rect 1674 68 1856 95
rect 1976 200 2080 232
rect 1976 154 2005 200
rect 2051 154 2080 200
rect 1976 68 2080 154
rect 2200 127 2304 232
rect 2200 81 2229 127
rect 2275 81 2304 127
rect 2200 68 2304 81
rect 2424 200 2512 232
rect 2424 154 2453 200
rect 2499 154 2512 200
rect 2424 68 2512 154
<< mvpdiff >>
rect 96 650 184 716
rect 96 510 109 650
rect 155 510 184 650
rect 96 497 184 510
rect 284 670 388 716
rect 284 624 313 670
rect 359 624 388 670
rect 284 497 388 624
rect 488 677 592 716
rect 488 631 517 677
rect 563 631 592 677
rect 488 497 592 631
rect 692 567 780 716
rect 692 521 721 567
rect 767 521 780 567
rect 692 497 780 521
rect 992 556 1080 716
rect 992 510 1005 556
rect 1051 510 1080 556
rect 992 497 1080 510
rect 1180 703 1320 716
rect 1180 657 1228 703
rect 1274 657 1320 703
rect 1180 515 1320 657
rect 1420 611 1524 716
rect 1420 565 1449 611
rect 1495 565 1524 611
rect 1420 515 1524 565
rect 1624 703 1764 716
rect 1624 563 1667 703
rect 1713 563 1764 703
rect 1624 515 1764 563
rect 1180 497 1260 515
rect 1684 480 1764 515
rect 1864 633 1968 716
rect 1864 493 1893 633
rect 1939 493 1968 633
rect 1864 480 1968 493
rect 2068 690 2172 716
rect 2068 644 2097 690
rect 2143 644 2172 690
rect 2068 480 2172 644
rect 2272 633 2360 716
rect 2272 493 2301 633
rect 2347 493 2360 633
rect 2272 480 2360 493
<< mvndiffc >>
rect 60 146 106 192
rect 284 93 330 139
rect 508 120 554 166
rect 776 198 822 244
rect 951 198 997 244
rect 1237 81 1283 127
rect 1479 117 1525 163
rect 1745 95 1791 141
rect 2005 154 2051 200
rect 2229 81 2275 127
rect 2453 154 2499 200
<< mvpdiffc >>
rect 109 510 155 650
rect 313 624 359 670
rect 517 631 563 677
rect 721 521 767 567
rect 1005 510 1051 556
rect 1228 657 1274 703
rect 1449 565 1495 611
rect 1667 563 1713 703
rect 1893 493 1939 633
rect 2097 644 2143 690
rect 2301 493 2347 633
<< polysilicon >>
rect 184 716 284 760
rect 388 716 488 760
rect 592 716 692 760
rect 1080 716 1180 760
rect 1320 716 1420 760
rect 1524 716 1624 760
rect 1764 716 1864 760
rect 1968 716 2068 760
rect 2172 716 2272 760
rect 184 412 284 497
rect 388 412 488 497
rect 592 464 692 497
rect 592 418 605 464
rect 651 418 692 464
rect 135 377 544 412
rect 592 405 692 418
rect 1080 410 1180 497
rect 135 331 183 377
rect 229 372 544 377
rect 229 331 255 372
rect 135 232 255 331
rect 504 357 544 372
rect 1080 364 1107 410
rect 1153 364 1180 410
rect 359 311 431 324
rect 504 317 623 357
rect 1080 326 1180 364
rect 359 265 372 311
rect 418 276 431 311
rect 583 288 623 317
rect 418 265 479 276
rect 359 232 479 265
rect 583 232 703 288
rect 1070 287 1180 326
rect 1320 459 1420 515
rect 1320 319 1349 459
rect 1395 324 1420 459
rect 1524 324 1624 515
rect 1764 439 1864 480
rect 1764 393 1791 439
rect 1837 420 1864 439
rect 1968 439 2068 480
rect 1968 420 1996 439
rect 1837 393 1996 420
rect 2042 420 2068 439
rect 2172 439 2272 480
rect 2172 420 2202 439
rect 2042 393 2202 420
rect 2248 393 2272 439
rect 1764 380 2272 393
rect 1395 319 1624 324
rect 1320 311 1624 319
rect 1070 232 1190 287
rect 1320 280 1443 311
rect 1330 265 1443 280
rect 1583 288 1624 311
rect 1856 319 2424 332
rect 1583 265 1674 288
rect 1330 252 1674 265
rect 1330 176 1450 252
rect 1554 176 1674 252
rect 1856 273 1889 319
rect 1935 292 2119 319
rect 1935 273 1976 292
rect 1856 232 1976 273
rect 2080 273 2119 292
rect 2165 292 2317 319
rect 2165 273 2200 292
rect 2080 232 2200 273
rect 2304 273 2317 292
rect 2363 273 2424 319
rect 2304 232 2424 273
rect 135 24 255 68
rect 359 24 479 68
rect 583 24 703 68
rect 1070 24 1190 68
rect 1330 24 1450 68
rect 1554 24 1674 68
rect 1856 24 1976 68
rect 2080 24 2200 68
rect 2304 24 2424 68
<< polycontact >>
rect 605 418 651 464
rect 183 331 229 377
rect 1107 364 1153 410
rect 372 265 418 311
rect 1349 319 1395 459
rect 1791 393 1837 439
rect 1996 393 2042 439
rect 2202 393 2248 439
rect 1443 265 1583 311
rect 1889 273 1935 319
rect 2119 273 2165 319
rect 2317 273 2363 319
<< metal1 >>
rect 0 724 2576 844
rect 313 670 359 724
rect 1217 703 1285 724
rect 109 650 155 661
rect 506 677 1143 678
rect 506 631 517 677
rect 563 631 1143 677
rect 1217 657 1228 703
rect 1274 657 1285 703
rect 1667 703 1713 724
rect 313 613 359 624
rect 720 567 767 578
rect 155 510 651 558
rect 109 499 651 510
rect 372 464 651 499
rect 132 377 320 430
rect 132 331 183 377
rect 229 331 320 377
rect 132 330 320 331
rect 372 418 605 464
rect 372 407 651 418
rect 720 521 721 567
rect 372 311 418 407
rect 720 361 767 521
rect 372 245 418 265
rect 60 198 418 245
rect 606 315 767 361
rect 60 192 106 198
rect 606 177 652 315
rect 813 269 859 631
rect 1097 611 1143 631
rect 1005 556 1051 574
rect 1097 565 1449 611
rect 1495 565 1621 611
rect 1051 510 1395 518
rect 1005 471 1395 510
rect 1349 459 1395 471
rect 906 410 1222 425
rect 906 364 1107 410
rect 1153 364 1222 410
rect 906 358 1222 364
rect 1575 439 1621 565
rect 2097 690 2143 724
rect 2097 633 2143 644
rect 1667 552 1713 563
rect 1882 493 1893 633
rect 1939 532 1950 633
rect 2290 532 2301 633
rect 1939 493 2301 532
rect 2347 550 2358 633
rect 2347 493 2552 550
rect 1882 485 2552 493
rect 1575 393 1791 439
rect 1837 393 1996 439
rect 2042 393 2202 439
rect 2248 393 2273 439
rect 1575 392 2273 393
rect 1349 312 1395 319
rect 763 244 859 269
rect 1024 311 1395 312
rect 1024 265 1443 311
rect 1583 265 1594 311
rect 1640 273 1889 319
rect 1935 273 2119 319
rect 2165 273 2317 319
rect 2363 273 2374 319
rect 1024 244 1070 265
rect 763 198 776 244
rect 822 198 859 244
rect 940 198 951 244
rect 997 198 1070 244
rect 1640 219 1686 273
rect 2453 220 2552 485
rect 508 166 652 177
rect 60 135 106 146
rect 284 139 330 152
rect 554 152 652 166
rect 1116 173 1686 219
rect 2005 200 2552 220
rect 1116 152 1162 173
rect 554 120 1162 152
rect 1479 163 1525 173
rect 508 106 1162 120
rect 284 60 330 93
rect 1226 81 1237 127
rect 1283 81 1294 127
rect 1479 106 1525 117
rect 1745 141 1791 180
rect 1226 60 1294 81
rect 2051 173 2453 200
rect 2005 123 2051 154
rect 2499 154 2552 200
rect 1745 60 1791 95
rect 2218 81 2229 127
rect 2275 81 2286 127
rect 2453 122 2552 154
rect 2218 60 2286 81
rect 0 -60 2576 60
<< labels >>
flabel metal1 s 0 724 2576 844 0 FreeSans 400 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 1745 152 1791 180 0 FreeSans 400 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel metal1 s 2290 550 2358 633 0 FreeSans 400 0 0 0 ZN
port 3 nsew default output
flabel metal1 s 132 330 320 430 0 FreeSans 400 0 0 0 EN
port 1 nsew default input
flabel metal1 s 906 358 1222 425 0 FreeSans 400 0 0 0 I
port 2 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 5 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 6 nsew ground bidirectional
rlabel metal1 s 1882 550 1950 633 1 ZN
port 3 nsew default output
rlabel metal1 s 2290 532 2552 550 1 ZN
port 3 nsew default output
rlabel metal1 s 1882 532 1950 550 1 ZN
port 3 nsew default output
rlabel metal1 s 1882 485 2552 532 1 ZN
port 3 nsew default output
rlabel metal1 s 2453 220 2552 485 1 ZN
port 3 nsew default output
rlabel metal1 s 2005 173 2552 220 1 ZN
port 3 nsew default output
rlabel metal1 s 2453 123 2552 173 1 ZN
port 3 nsew default output
rlabel metal1 s 2005 123 2051 173 1 ZN
port 3 nsew default output
rlabel metal1 s 2453 122 2552 123 1 ZN
port 3 nsew default output
rlabel metal1 s 2097 657 2143 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1667 657 1713 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1217 657 1285 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 313 657 359 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2097 633 2143 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1667 633 1713 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 313 633 359 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1667 613 1713 633 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 313 613 359 633 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1667 552 1713 613 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1745 127 1791 152 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 284 127 330 152 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2218 60 2286 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1745 60 1791 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1226 60 1294 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 284 60 330 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 2576 60 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2576 784
string GDS_END 534198
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 527684
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
