magic
tech gf180mcuA
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 352 1654 870
<< pwell >>
rect -86 -86 1654 352
<< mvnmos >>
rect 124 72 244 165
rect 348 72 468 165
rect 572 72 692 165
rect 796 72 916 165
rect 1056 68 1176 232
rect 1280 68 1400 232
<< mvpmos >>
rect 144 472 244 716
rect 368 472 468 716
rect 592 472 692 716
rect 816 472 916 716
rect 1066 472 1166 716
rect 1280 472 1380 716
<< mvndiff >>
rect 976 165 1056 232
rect 36 131 124 165
rect 36 85 49 131
rect 95 85 124 131
rect 36 72 124 85
rect 244 152 348 165
rect 244 106 273 152
rect 319 106 348 152
rect 244 72 348 106
rect 468 131 572 165
rect 468 85 497 131
rect 543 85 572 131
rect 468 72 572 85
rect 692 152 796 165
rect 692 106 721 152
rect 767 106 796 152
rect 692 72 796 106
rect 916 131 1056 165
rect 916 85 945 131
rect 991 85 1056 131
rect 916 72 1056 85
rect 976 68 1056 72
rect 1176 192 1280 232
rect 1176 146 1205 192
rect 1251 146 1280 192
rect 1176 68 1280 146
rect 1400 157 1488 232
rect 1400 111 1429 157
rect 1475 111 1488 157
rect 1400 68 1488 111
<< mvpdiff >>
rect 56 665 144 716
rect 56 525 69 665
rect 115 525 144 665
rect 56 472 144 525
rect 244 472 368 716
rect 468 472 592 716
rect 692 472 816 716
rect 916 665 1066 716
rect 916 525 964 665
rect 1010 525 1066 665
rect 916 472 1066 525
rect 1166 665 1280 716
rect 1166 525 1195 665
rect 1241 525 1280 665
rect 1166 472 1280 525
rect 1380 664 1468 716
rect 1380 618 1409 664
rect 1455 618 1468 664
rect 1380 472 1468 618
<< mvndiffc >>
rect 49 85 95 131
rect 273 106 319 152
rect 497 85 543 131
rect 721 106 767 152
rect 945 85 991 131
rect 1205 146 1251 192
rect 1429 111 1475 157
<< mvpdiffc >>
rect 69 525 115 665
rect 964 525 1010 665
rect 1195 525 1241 665
rect 1409 618 1455 664
<< polysilicon >>
rect 144 716 244 760
rect 368 716 468 760
rect 592 716 692 760
rect 816 716 916 760
rect 1066 716 1166 760
rect 1280 716 1380 760
rect 144 408 244 472
rect 368 408 468 472
rect 592 408 692 472
rect 816 408 916 472
rect 124 389 244 408
rect 124 343 147 389
rect 193 343 244 389
rect 124 165 244 343
rect 348 389 468 408
rect 348 343 371 389
rect 417 343 468 389
rect 348 165 468 343
rect 572 389 692 408
rect 572 343 595 389
rect 641 343 692 389
rect 572 165 692 343
rect 796 389 916 408
rect 796 343 819 389
rect 865 343 916 389
rect 796 165 916 343
rect 1066 415 1166 472
rect 1066 369 1094 415
rect 1140 394 1166 415
rect 1280 415 1380 472
rect 1280 394 1293 415
rect 1140 369 1293 394
rect 1339 369 1380 415
rect 1066 348 1380 369
rect 1066 277 1176 348
rect 1056 232 1176 277
rect 1280 277 1380 348
rect 1280 232 1400 277
rect 124 28 244 72
rect 348 28 468 72
rect 572 28 692 72
rect 796 28 916 72
rect 1056 24 1176 68
rect 1280 24 1400 68
<< polycontact >>
rect 147 343 193 389
rect 371 343 417 389
rect 595 343 641 389
rect 819 343 865 389
rect 1094 369 1140 415
rect 1293 369 1339 415
<< metal1 >>
rect 0 724 1568 844
rect 69 665 115 678
rect 115 525 308 552
rect 69 506 308 525
rect 132 389 204 458
rect 132 343 147 389
rect 193 343 204 389
rect 132 203 204 343
rect 262 236 308 506
rect 356 389 428 678
rect 356 343 371 389
rect 417 343 428 389
rect 356 296 428 343
rect 580 389 652 678
rect 580 343 595 389
rect 641 343 652 389
rect 580 296 652 343
rect 804 389 876 678
rect 964 665 1010 724
rect 964 506 1010 525
rect 1194 665 1317 678
rect 1194 525 1195 665
rect 1241 536 1317 665
rect 1409 664 1455 724
rect 1409 598 1455 618
rect 1241 525 1456 536
rect 1194 472 1456 525
rect 804 343 819 389
rect 865 343 876 389
rect 804 296 876 343
rect 1006 369 1094 415
rect 1140 369 1293 415
rect 1339 369 1350 415
rect 1006 236 1052 369
rect 1402 312 1456 472
rect 262 189 1052 236
rect 1205 248 1456 312
rect 1205 192 1317 248
rect 262 152 330 189
rect 38 85 49 131
rect 95 85 106 131
rect 262 106 273 152
rect 319 106 330 152
rect 710 152 778 189
rect 38 60 106 85
rect 486 85 497 131
rect 543 85 554 131
rect 710 106 721 152
rect 767 106 778 152
rect 1251 146 1317 192
rect 486 60 554 85
rect 934 85 945 131
rect 991 85 1002 131
rect 1205 106 1317 146
rect 1429 157 1475 180
rect 934 60 1002 85
rect 1429 60 1475 111
rect 0 -60 1568 60
<< labels >>
flabel metal1 s 132 203 204 458 0 FreeSans 400 0 0 0 A1
port 1 nsew default input
flabel metal1 s 580 296 652 678 0 FreeSans 400 0 0 0 A3
port 3 nsew default input
flabel metal1 s 804 296 876 678 0 FreeSans 400 0 0 0 A4
port 4 nsew default input
flabel metal1 s 0 724 1568 844 0 FreeSans 400 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 1429 131 1475 180 0 FreeSans 400 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel metal1 s 1194 536 1317 678 0 FreeSans 400 0 0 0 Z
port 5 nsew default output
flabel metal1 s 356 296 428 678 0 FreeSans 400 0 0 0 A2
port 2 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 7 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 8 nsew ground bidirectional
rlabel metal1 s 1194 472 1456 536 1 Z
port 5 nsew default output
rlabel metal1 s 1402 312 1456 472 1 Z
port 5 nsew default output
rlabel metal1 s 1205 248 1456 312 1 Z
port 5 nsew default output
rlabel metal1 s 1205 106 1317 248 1 Z
port 5 nsew default output
rlabel metal1 s 1409 598 1455 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 964 598 1010 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 964 506 1010 598 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1429 60 1475 131 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 934 60 1002 131 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 486 60 554 131 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 38 60 106 131 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 1568 60 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1568 784
string GDS_END 175942
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 171784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
