magic
tech gf180mcuA
magscale 1 10
timestamp 1698431365
<< isosubstrate >>
rect -1470 -83 6872 2575
<< nwell >>
rect -1402 1487 6872 2575
rect 0 1281 6872 1487
rect 251 1215 1051 1281
<< mvnmos >>
rect 459 280 599 680
rect 703 280 843 680
rect 1170 620 1310 920
rect 1747 280 1887 920
rect 1991 280 2131 920
rect 2235 280 2375 920
rect 2479 280 2619 920
rect 2723 280 2863 920
rect 3203 338 3343 868
rect 3447 338 3587 868
rect 3691 338 3831 868
rect 3935 338 4075 868
rect 4323 268 4463 868
rect 4567 268 4707 868
rect 4811 268 4951 868
rect 5055 268 5195 868
rect 5443 608 5583 868
rect 5831 731 5971 1031
rect 6219 731 6359 1031
<< mvpmos >>
rect 459 1335 599 2135
rect 703 1335 843 2135
rect 1669 1797 1809 2097
rect 1913 1797 2053 2097
rect 2365 1797 2505 2197
rect 2609 1797 2749 2197
rect 2853 1797 2993 2197
rect 3315 1730 3455 2110
rect 3559 1730 3699 2110
rect 4183 1730 4323 2160
rect 4427 1730 4567 2160
rect 4815 1730 4955 2110
rect 5059 1730 5199 2110
rect 5831 1637 5971 2037
rect 6219 1637 6359 2037
<< mvndiff >>
rect 1082 907 1170 920
rect 1082 861 1095 907
rect 1141 861 1170 907
rect 1082 793 1170 861
rect 1082 747 1095 793
rect 1141 747 1170 793
rect 371 667 459 680
rect 371 621 384 667
rect 430 621 459 667
rect 371 558 459 621
rect 371 512 384 558
rect 430 512 459 558
rect 371 449 459 512
rect 371 403 384 449
rect 430 403 459 449
rect 371 339 459 403
rect 371 293 384 339
rect 430 293 459 339
rect 371 280 459 293
rect 599 667 703 680
rect 599 621 628 667
rect 674 621 703 667
rect 599 558 703 621
rect 599 512 628 558
rect 674 512 703 558
rect 599 449 703 512
rect 599 403 628 449
rect 674 403 703 449
rect 599 339 703 403
rect 599 293 628 339
rect 674 293 703 339
rect 599 280 703 293
rect 843 667 931 680
rect 843 621 872 667
rect 918 621 931 667
rect 843 558 931 621
rect 1082 679 1170 747
rect 1082 633 1095 679
rect 1141 633 1170 679
rect 1082 620 1170 633
rect 1310 907 1398 920
rect 1310 861 1339 907
rect 1385 861 1398 907
rect 1310 793 1398 861
rect 1310 747 1339 793
rect 1385 747 1398 793
rect 1310 679 1398 747
rect 1310 633 1339 679
rect 1385 633 1398 679
rect 1310 620 1398 633
rect 1659 907 1747 920
rect 1659 861 1672 907
rect 1718 861 1747 907
rect 1659 794 1747 861
rect 1659 748 1672 794
rect 1718 748 1747 794
rect 1659 681 1747 748
rect 1659 635 1672 681
rect 1718 635 1747 681
rect 843 512 872 558
rect 918 512 931 558
rect 843 449 931 512
rect 843 403 872 449
rect 918 403 931 449
rect 843 339 931 403
rect 843 293 872 339
rect 918 293 931 339
rect 843 280 931 293
rect 1659 567 1747 635
rect 1659 521 1672 567
rect 1718 521 1747 567
rect 1659 453 1747 521
rect 1659 407 1672 453
rect 1718 407 1747 453
rect 1659 339 1747 407
rect 1659 293 1672 339
rect 1718 293 1747 339
rect 1659 280 1747 293
rect 1887 907 1991 920
rect 1887 861 1916 907
rect 1962 861 1991 907
rect 1887 794 1991 861
rect 1887 748 1916 794
rect 1962 748 1991 794
rect 1887 681 1991 748
rect 1887 635 1916 681
rect 1962 635 1991 681
rect 1887 567 1991 635
rect 1887 521 1916 567
rect 1962 521 1991 567
rect 1887 453 1991 521
rect 1887 407 1916 453
rect 1962 407 1991 453
rect 1887 339 1991 407
rect 1887 293 1916 339
rect 1962 293 1991 339
rect 1887 280 1991 293
rect 2131 907 2235 920
rect 2131 861 2160 907
rect 2206 861 2235 907
rect 2131 794 2235 861
rect 2131 748 2160 794
rect 2206 748 2235 794
rect 2131 681 2235 748
rect 2131 635 2160 681
rect 2206 635 2235 681
rect 2131 567 2235 635
rect 2131 521 2160 567
rect 2206 521 2235 567
rect 2131 453 2235 521
rect 2131 407 2160 453
rect 2206 407 2235 453
rect 2131 339 2235 407
rect 2131 293 2160 339
rect 2206 293 2235 339
rect 2131 280 2235 293
rect 2375 907 2479 920
rect 2375 861 2404 907
rect 2450 861 2479 907
rect 2375 794 2479 861
rect 2375 748 2404 794
rect 2450 748 2479 794
rect 2375 681 2479 748
rect 2375 635 2404 681
rect 2450 635 2479 681
rect 2375 567 2479 635
rect 2375 521 2404 567
rect 2450 521 2479 567
rect 2375 453 2479 521
rect 2375 407 2404 453
rect 2450 407 2479 453
rect 2375 339 2479 407
rect 2375 293 2404 339
rect 2450 293 2479 339
rect 2375 280 2479 293
rect 2619 907 2723 920
rect 2619 861 2648 907
rect 2694 861 2723 907
rect 2619 794 2723 861
rect 2619 748 2648 794
rect 2694 748 2723 794
rect 2619 681 2723 748
rect 2619 635 2648 681
rect 2694 635 2723 681
rect 2619 567 2723 635
rect 2619 521 2648 567
rect 2694 521 2723 567
rect 2619 453 2723 521
rect 2619 407 2648 453
rect 2694 407 2723 453
rect 2619 339 2723 407
rect 2619 293 2648 339
rect 2694 293 2723 339
rect 2619 280 2723 293
rect 2863 907 2951 920
rect 2863 861 2892 907
rect 2938 861 2951 907
rect 5743 1018 5831 1031
rect 5743 972 5756 1018
rect 5802 972 5831 1018
rect 5743 904 5831 972
rect 2863 794 2951 861
rect 2863 748 2892 794
rect 2938 748 2951 794
rect 2863 681 2951 748
rect 2863 635 2892 681
rect 2938 635 2951 681
rect 2863 567 2951 635
rect 2863 521 2892 567
rect 2938 521 2951 567
rect 2863 453 2951 521
rect 2863 407 2892 453
rect 2938 407 2951 453
rect 2863 339 2951 407
rect 2863 293 2892 339
rect 2938 293 2951 339
rect 3115 855 3203 868
rect 3115 809 3128 855
rect 3174 809 3203 855
rect 3115 741 3203 809
rect 3115 695 3128 741
rect 3174 695 3203 741
rect 3115 627 3203 695
rect 3115 581 3128 627
rect 3174 581 3203 627
rect 3115 512 3203 581
rect 3115 466 3128 512
rect 3174 466 3203 512
rect 3115 397 3203 466
rect 3115 351 3128 397
rect 3174 351 3203 397
rect 3115 338 3203 351
rect 3343 855 3447 868
rect 3343 809 3372 855
rect 3418 809 3447 855
rect 3343 741 3447 809
rect 3343 695 3372 741
rect 3418 695 3447 741
rect 3343 627 3447 695
rect 3343 581 3372 627
rect 3418 581 3447 627
rect 3343 512 3447 581
rect 3343 466 3372 512
rect 3418 466 3447 512
rect 3343 397 3447 466
rect 3343 351 3372 397
rect 3418 351 3447 397
rect 3343 338 3447 351
rect 3587 855 3691 868
rect 3587 809 3616 855
rect 3662 809 3691 855
rect 3587 741 3691 809
rect 3587 695 3616 741
rect 3662 695 3691 741
rect 3587 627 3691 695
rect 3587 581 3616 627
rect 3662 581 3691 627
rect 3587 512 3691 581
rect 3587 466 3616 512
rect 3662 466 3691 512
rect 3587 397 3691 466
rect 3587 351 3616 397
rect 3662 351 3691 397
rect 3587 338 3691 351
rect 3831 855 3935 868
rect 3831 809 3860 855
rect 3906 809 3935 855
rect 3831 741 3935 809
rect 3831 695 3860 741
rect 3906 695 3935 741
rect 3831 627 3935 695
rect 3831 581 3860 627
rect 3906 581 3935 627
rect 3831 512 3935 581
rect 3831 466 3860 512
rect 3906 466 3935 512
rect 3831 397 3935 466
rect 3831 351 3860 397
rect 3906 351 3935 397
rect 3831 338 3935 351
rect 4075 855 4163 868
rect 4075 809 4104 855
rect 4150 809 4163 855
rect 4075 741 4163 809
rect 4075 695 4104 741
rect 4150 695 4163 741
rect 4075 627 4163 695
rect 4075 581 4104 627
rect 4150 581 4163 627
rect 4075 512 4163 581
rect 4075 466 4104 512
rect 4150 466 4163 512
rect 4075 397 4163 466
rect 4075 351 4104 397
rect 4150 351 4163 397
rect 4075 338 4163 351
rect 4235 855 4323 868
rect 4235 809 4248 855
rect 4294 809 4323 855
rect 4235 750 4323 809
rect 4235 704 4248 750
rect 4294 704 4323 750
rect 4235 645 4323 704
rect 4235 599 4248 645
rect 4294 599 4323 645
rect 4235 539 4323 599
rect 4235 493 4248 539
rect 4294 493 4323 539
rect 4235 433 4323 493
rect 4235 387 4248 433
rect 4294 387 4323 433
rect 4235 327 4323 387
rect 2863 280 2951 293
rect 4235 281 4248 327
rect 4294 281 4323 327
rect 4235 268 4323 281
rect 4463 855 4567 868
rect 4463 809 4492 855
rect 4538 809 4567 855
rect 4463 750 4567 809
rect 4463 704 4492 750
rect 4538 704 4567 750
rect 4463 645 4567 704
rect 4463 599 4492 645
rect 4538 599 4567 645
rect 4463 539 4567 599
rect 4463 493 4492 539
rect 4538 493 4567 539
rect 4463 433 4567 493
rect 4463 387 4492 433
rect 4538 387 4567 433
rect 4463 327 4567 387
rect 4463 281 4492 327
rect 4538 281 4567 327
rect 4463 268 4567 281
rect 4707 855 4811 868
rect 4707 809 4736 855
rect 4782 809 4811 855
rect 4707 750 4811 809
rect 4707 704 4736 750
rect 4782 704 4811 750
rect 4707 645 4811 704
rect 4707 599 4736 645
rect 4782 599 4811 645
rect 4707 539 4811 599
rect 4707 493 4736 539
rect 4782 493 4811 539
rect 4707 433 4811 493
rect 4707 387 4736 433
rect 4782 387 4811 433
rect 4707 327 4811 387
rect 4707 281 4736 327
rect 4782 281 4811 327
rect 4707 268 4811 281
rect 4951 855 5055 868
rect 4951 809 4980 855
rect 5026 809 5055 855
rect 4951 750 5055 809
rect 4951 704 4980 750
rect 5026 704 5055 750
rect 4951 645 5055 704
rect 4951 599 4980 645
rect 5026 599 5055 645
rect 4951 539 5055 599
rect 4951 493 4980 539
rect 5026 493 5055 539
rect 4951 433 5055 493
rect 4951 387 4980 433
rect 5026 387 5055 433
rect 4951 327 5055 387
rect 4951 281 4980 327
rect 5026 281 5055 327
rect 4951 268 5055 281
rect 5195 855 5283 868
rect 5195 809 5224 855
rect 5270 809 5283 855
rect 5195 750 5283 809
rect 5195 704 5224 750
rect 5270 704 5283 750
rect 5195 645 5283 704
rect 5195 599 5224 645
rect 5270 599 5283 645
rect 5355 855 5443 868
rect 5355 809 5368 855
rect 5414 809 5443 855
rect 5355 667 5443 809
rect 5355 621 5368 667
rect 5414 621 5443 667
rect 5355 608 5443 621
rect 5583 855 5671 868
rect 5583 809 5612 855
rect 5658 809 5671 855
rect 5583 667 5671 809
rect 5743 858 5756 904
rect 5802 858 5831 904
rect 5743 790 5831 858
rect 5743 744 5756 790
rect 5802 744 5831 790
rect 5743 731 5831 744
rect 5971 1018 6059 1031
rect 5971 972 6000 1018
rect 6046 972 6059 1018
rect 5971 904 6059 972
rect 5971 858 6000 904
rect 6046 858 6059 904
rect 5971 790 6059 858
rect 5971 744 6000 790
rect 6046 744 6059 790
rect 5971 731 6059 744
rect 6131 1018 6219 1031
rect 6131 972 6144 1018
rect 6190 972 6219 1018
rect 6131 904 6219 972
rect 6131 858 6144 904
rect 6190 858 6219 904
rect 6131 790 6219 858
rect 6131 744 6144 790
rect 6190 744 6219 790
rect 6131 731 6219 744
rect 6359 1018 6447 1031
rect 6359 972 6388 1018
rect 6434 972 6447 1018
rect 6359 904 6447 972
rect 6359 858 6388 904
rect 6434 858 6447 904
rect 6359 790 6447 858
rect 6359 744 6388 790
rect 6434 744 6447 790
rect 6359 731 6447 744
rect 5583 621 5612 667
rect 5658 621 5671 667
rect 5583 608 5671 621
rect 5195 539 5283 599
rect 5195 493 5224 539
rect 5270 493 5283 539
rect 5195 433 5283 493
rect 5195 387 5224 433
rect 5270 387 5283 433
rect 5195 327 5283 387
rect 5195 281 5224 327
rect 5270 281 5283 327
rect 5195 268 5283 281
<< mvpdiff >>
rect 2277 2184 2365 2197
rect 371 2122 459 2135
rect 371 2076 384 2122
rect 430 2076 459 2122
rect 371 2018 459 2076
rect 371 1972 384 2018
rect 430 1972 459 2018
rect 371 1914 459 1972
rect 371 1868 384 1914
rect 430 1868 459 1914
rect 371 1810 459 1868
rect 371 1764 384 1810
rect 430 1764 459 1810
rect 371 1706 459 1764
rect 371 1660 384 1706
rect 430 1660 459 1706
rect 371 1602 459 1660
rect 371 1556 384 1602
rect 430 1556 459 1602
rect 371 1498 459 1556
rect 371 1452 384 1498
rect 430 1452 459 1498
rect 371 1394 459 1452
rect 371 1348 384 1394
rect 430 1348 459 1394
rect 371 1335 459 1348
rect 599 2122 703 2135
rect 599 2076 628 2122
rect 674 2076 703 2122
rect 599 2018 703 2076
rect 599 1972 628 2018
rect 674 1972 703 2018
rect 599 1914 703 1972
rect 599 1868 628 1914
rect 674 1868 703 1914
rect 599 1810 703 1868
rect 599 1764 628 1810
rect 674 1764 703 1810
rect 599 1706 703 1764
rect 599 1660 628 1706
rect 674 1660 703 1706
rect 599 1602 703 1660
rect 599 1556 628 1602
rect 674 1556 703 1602
rect 599 1498 703 1556
rect 599 1452 628 1498
rect 674 1452 703 1498
rect 599 1394 703 1452
rect 599 1348 628 1394
rect 674 1348 703 1394
rect 599 1335 703 1348
rect 843 2122 931 2135
rect 843 2076 872 2122
rect 918 2076 931 2122
rect 2277 2138 2290 2184
rect 2336 2138 2365 2184
rect 843 2018 931 2076
rect 843 1972 872 2018
rect 918 1972 931 2018
rect 843 1914 931 1972
rect 843 1868 872 1914
rect 918 1868 931 1914
rect 843 1810 931 1868
rect 843 1764 872 1810
rect 918 1764 931 1810
rect 1581 2084 1669 2097
rect 1581 2038 1594 2084
rect 1640 2038 1669 2084
rect 1581 1970 1669 2038
rect 1581 1924 1594 1970
rect 1640 1924 1669 1970
rect 1581 1856 1669 1924
rect 1581 1810 1594 1856
rect 1640 1810 1669 1856
rect 1581 1797 1669 1810
rect 1809 2084 1913 2097
rect 1809 2038 1838 2084
rect 1884 2038 1913 2084
rect 1809 1970 1913 2038
rect 1809 1924 1838 1970
rect 1884 1924 1913 1970
rect 1809 1856 1913 1924
rect 1809 1810 1838 1856
rect 1884 1810 1913 1856
rect 1809 1797 1913 1810
rect 2053 2084 2141 2097
rect 2053 2038 2082 2084
rect 2128 2038 2141 2084
rect 2053 1970 2141 2038
rect 2053 1924 2082 1970
rect 2128 1924 2141 1970
rect 2053 1856 2141 1924
rect 2053 1810 2082 1856
rect 2128 1810 2141 1856
rect 2053 1797 2141 1810
rect 2277 2074 2365 2138
rect 2277 2028 2290 2074
rect 2336 2028 2365 2074
rect 2277 1965 2365 2028
rect 2277 1919 2290 1965
rect 2336 1919 2365 1965
rect 2277 1856 2365 1919
rect 2277 1810 2290 1856
rect 2336 1810 2365 1856
rect 2277 1797 2365 1810
rect 2505 2184 2609 2197
rect 2505 2138 2534 2184
rect 2580 2138 2609 2184
rect 2505 2074 2609 2138
rect 2505 2028 2534 2074
rect 2580 2028 2609 2074
rect 2505 1965 2609 2028
rect 2505 1919 2534 1965
rect 2580 1919 2609 1965
rect 2505 1856 2609 1919
rect 2505 1810 2534 1856
rect 2580 1810 2609 1856
rect 2505 1797 2609 1810
rect 2749 2184 2853 2197
rect 2749 2138 2778 2184
rect 2824 2138 2853 2184
rect 2749 2074 2853 2138
rect 2749 2028 2778 2074
rect 2824 2028 2853 2074
rect 2749 1965 2853 2028
rect 2749 1919 2778 1965
rect 2824 1919 2853 1965
rect 2749 1856 2853 1919
rect 2749 1810 2778 1856
rect 2824 1810 2853 1856
rect 2749 1797 2853 1810
rect 2993 2184 3081 2197
rect 2993 2138 3022 2184
rect 3068 2138 3081 2184
rect 2993 2074 3081 2138
rect 4095 2147 4183 2160
rect 2993 2028 3022 2074
rect 3068 2028 3081 2074
rect 2993 1965 3081 2028
rect 2993 1919 3022 1965
rect 3068 1919 3081 1965
rect 2993 1856 3081 1919
rect 2993 1810 3022 1856
rect 3068 1810 3081 1856
rect 2993 1797 3081 1810
rect 3227 2097 3315 2110
rect 3227 1949 3240 2097
rect 3286 1949 3315 2097
rect 3227 1892 3315 1949
rect 3227 1846 3240 1892
rect 3286 1846 3315 1892
rect 843 1706 931 1764
rect 843 1660 872 1706
rect 918 1660 931 1706
rect 843 1602 931 1660
rect 3227 1789 3315 1846
rect 3227 1743 3240 1789
rect 3286 1743 3315 1789
rect 3227 1730 3315 1743
rect 3455 2097 3559 2110
rect 3455 1949 3484 2097
rect 3530 1949 3559 2097
rect 3455 1892 3559 1949
rect 3455 1846 3484 1892
rect 3530 1846 3559 1892
rect 3455 1789 3559 1846
rect 3455 1743 3484 1789
rect 3530 1743 3559 1789
rect 3455 1730 3559 1743
rect 3699 2097 3787 2110
rect 3699 1949 3728 2097
rect 3774 1949 3787 2097
rect 3699 1892 3787 1949
rect 3699 1846 3728 1892
rect 3774 1846 3787 1892
rect 3699 1789 3787 1846
rect 3699 1743 3728 1789
rect 3774 1743 3787 1789
rect 3699 1730 3787 1743
rect 4095 2101 4108 2147
rect 4154 2101 4183 2147
rect 4095 2028 4183 2101
rect 4095 1982 4108 2028
rect 4154 1982 4183 2028
rect 4095 1909 4183 1982
rect 4095 1863 4108 1909
rect 4154 1863 4183 1909
rect 4095 1789 4183 1863
rect 4095 1743 4108 1789
rect 4154 1743 4183 1789
rect 4095 1730 4183 1743
rect 4323 2147 4427 2160
rect 4323 2101 4352 2147
rect 4398 2101 4427 2147
rect 4323 2028 4427 2101
rect 4323 1982 4352 2028
rect 4398 1982 4427 2028
rect 4323 1909 4427 1982
rect 4323 1863 4352 1909
rect 4398 1863 4427 1909
rect 4323 1789 4427 1863
rect 4323 1743 4352 1789
rect 4398 1743 4427 1789
rect 4323 1730 4427 1743
rect 4567 2147 4655 2160
rect 4567 2101 4596 2147
rect 4642 2101 4655 2147
rect 4567 2028 4655 2101
rect 4567 1982 4596 2028
rect 4642 1982 4655 2028
rect 4567 1909 4655 1982
rect 4567 1863 4596 1909
rect 4642 1863 4655 1909
rect 4567 1789 4655 1863
rect 4567 1743 4596 1789
rect 4642 1743 4655 1789
rect 4567 1730 4655 1743
rect 4727 2097 4815 2110
rect 4727 1949 4740 2097
rect 4786 1949 4815 2097
rect 4727 1892 4815 1949
rect 4727 1846 4740 1892
rect 4786 1846 4815 1892
rect 4727 1789 4815 1846
rect 4727 1743 4740 1789
rect 4786 1743 4815 1789
rect 4727 1730 4815 1743
rect 4955 2097 5059 2110
rect 4955 1949 4984 2097
rect 5030 1949 5059 2097
rect 4955 1892 5059 1949
rect 4955 1846 4984 1892
rect 5030 1846 5059 1892
rect 4955 1789 5059 1846
rect 4955 1743 4984 1789
rect 5030 1743 5059 1789
rect 4955 1730 5059 1743
rect 5199 2097 5287 2110
rect 5199 1949 5228 2097
rect 5274 1949 5287 2097
rect 5199 1892 5287 1949
rect 5199 1846 5228 1892
rect 5274 1846 5287 1892
rect 5199 1789 5287 1846
rect 5199 1743 5228 1789
rect 5274 1743 5287 1789
rect 5199 1730 5287 1743
rect 5743 2024 5831 2037
rect 5743 1978 5756 2024
rect 5802 1978 5831 2024
rect 5743 1914 5831 1978
rect 5743 1868 5756 1914
rect 5802 1868 5831 1914
rect 5743 1805 5831 1868
rect 5743 1759 5756 1805
rect 5802 1759 5831 1805
rect 5743 1696 5831 1759
rect 5743 1650 5756 1696
rect 5802 1650 5831 1696
rect 843 1556 872 1602
rect 918 1556 931 1602
rect 5743 1637 5831 1650
rect 5971 2024 6059 2037
rect 5971 1978 6000 2024
rect 6046 1978 6059 2024
rect 5971 1914 6059 1978
rect 5971 1868 6000 1914
rect 6046 1868 6059 1914
rect 5971 1805 6059 1868
rect 5971 1759 6000 1805
rect 6046 1759 6059 1805
rect 5971 1696 6059 1759
rect 5971 1650 6000 1696
rect 6046 1650 6059 1696
rect 5971 1637 6059 1650
rect 6131 2024 6219 2037
rect 6131 1978 6144 2024
rect 6190 1978 6219 2024
rect 6131 1914 6219 1978
rect 6131 1868 6144 1914
rect 6190 1868 6219 1914
rect 6131 1805 6219 1868
rect 6131 1759 6144 1805
rect 6190 1759 6219 1805
rect 6131 1696 6219 1759
rect 6131 1650 6144 1696
rect 6190 1650 6219 1696
rect 6131 1637 6219 1650
rect 6359 2024 6447 2037
rect 6359 1978 6388 2024
rect 6434 1978 6447 2024
rect 6359 1914 6447 1978
rect 6359 1868 6388 1914
rect 6434 1868 6447 1914
rect 6359 1805 6447 1868
rect 6359 1759 6388 1805
rect 6434 1759 6447 1805
rect 6359 1696 6447 1759
rect 6359 1650 6388 1696
rect 6434 1650 6447 1696
rect 6359 1637 6447 1650
rect 843 1498 931 1556
rect 843 1452 872 1498
rect 918 1452 931 1498
rect 843 1394 931 1452
rect 843 1348 872 1394
rect 918 1348 931 1394
rect 843 1335 931 1348
<< mvndiffc >>
rect 1095 861 1141 907
rect 1095 747 1141 793
rect 384 621 430 667
rect 384 512 430 558
rect 384 403 430 449
rect 384 293 430 339
rect 628 621 674 667
rect 628 512 674 558
rect 628 403 674 449
rect 628 293 674 339
rect 872 621 918 667
rect 1095 633 1141 679
rect 1339 861 1385 907
rect 1339 747 1385 793
rect 1339 633 1385 679
rect 1672 861 1718 907
rect 1672 748 1718 794
rect 1672 635 1718 681
rect 872 512 918 558
rect 872 403 918 449
rect 872 293 918 339
rect 1672 521 1718 567
rect 1672 407 1718 453
rect 1672 293 1718 339
rect 1916 861 1962 907
rect 1916 748 1962 794
rect 1916 635 1962 681
rect 1916 521 1962 567
rect 1916 407 1962 453
rect 1916 293 1962 339
rect 2160 861 2206 907
rect 2160 748 2206 794
rect 2160 635 2206 681
rect 2160 521 2206 567
rect 2160 407 2206 453
rect 2160 293 2206 339
rect 2404 861 2450 907
rect 2404 748 2450 794
rect 2404 635 2450 681
rect 2404 521 2450 567
rect 2404 407 2450 453
rect 2404 293 2450 339
rect 2648 861 2694 907
rect 2648 748 2694 794
rect 2648 635 2694 681
rect 2648 521 2694 567
rect 2648 407 2694 453
rect 2648 293 2694 339
rect 2892 861 2938 907
rect 5756 972 5802 1018
rect 2892 748 2938 794
rect 2892 635 2938 681
rect 2892 521 2938 567
rect 2892 407 2938 453
rect 2892 293 2938 339
rect 3128 809 3174 855
rect 3128 695 3174 741
rect 3128 581 3174 627
rect 3128 466 3174 512
rect 3128 351 3174 397
rect 3372 809 3418 855
rect 3372 695 3418 741
rect 3372 581 3418 627
rect 3372 466 3418 512
rect 3372 351 3418 397
rect 3616 809 3662 855
rect 3616 695 3662 741
rect 3616 581 3662 627
rect 3616 466 3662 512
rect 3616 351 3662 397
rect 3860 809 3906 855
rect 3860 695 3906 741
rect 3860 581 3906 627
rect 3860 466 3906 512
rect 3860 351 3906 397
rect 4104 809 4150 855
rect 4104 695 4150 741
rect 4104 581 4150 627
rect 4104 466 4150 512
rect 4104 351 4150 397
rect 4248 809 4294 855
rect 4248 704 4294 750
rect 4248 599 4294 645
rect 4248 493 4294 539
rect 4248 387 4294 433
rect 4248 281 4294 327
rect 4492 809 4538 855
rect 4492 704 4538 750
rect 4492 599 4538 645
rect 4492 493 4538 539
rect 4492 387 4538 433
rect 4492 281 4538 327
rect 4736 809 4782 855
rect 4736 704 4782 750
rect 4736 599 4782 645
rect 4736 493 4782 539
rect 4736 387 4782 433
rect 4736 281 4782 327
rect 4980 809 5026 855
rect 4980 704 5026 750
rect 4980 599 5026 645
rect 4980 493 5026 539
rect 4980 387 5026 433
rect 4980 281 5026 327
rect 5224 809 5270 855
rect 5224 704 5270 750
rect 5224 599 5270 645
rect 5368 809 5414 855
rect 5368 621 5414 667
rect 5612 809 5658 855
rect 5756 858 5802 904
rect 5756 744 5802 790
rect 6000 972 6046 1018
rect 6000 858 6046 904
rect 6000 744 6046 790
rect 6144 972 6190 1018
rect 6144 858 6190 904
rect 6144 744 6190 790
rect 6388 972 6434 1018
rect 6388 858 6434 904
rect 6388 744 6434 790
rect 5612 621 5658 667
rect 5224 493 5270 539
rect 5224 387 5270 433
rect 5224 281 5270 327
<< mvpdiffc >>
rect 384 2076 430 2122
rect 384 1972 430 2018
rect 384 1868 430 1914
rect 384 1764 430 1810
rect 384 1660 430 1706
rect 384 1556 430 1602
rect 384 1452 430 1498
rect 384 1348 430 1394
rect 628 2076 674 2122
rect 628 1972 674 2018
rect 628 1868 674 1914
rect 628 1764 674 1810
rect 628 1660 674 1706
rect 628 1556 674 1602
rect 628 1452 674 1498
rect 628 1348 674 1394
rect 872 2076 918 2122
rect 2290 2138 2336 2184
rect 872 1972 918 2018
rect 872 1868 918 1914
rect 872 1764 918 1810
rect 1594 2038 1640 2084
rect 1594 1924 1640 1970
rect 1594 1810 1640 1856
rect 1838 2038 1884 2084
rect 1838 1924 1884 1970
rect 1838 1810 1884 1856
rect 2082 2038 2128 2084
rect 2082 1924 2128 1970
rect 2082 1810 2128 1856
rect 2290 2028 2336 2074
rect 2290 1919 2336 1965
rect 2290 1810 2336 1856
rect 2534 2138 2580 2184
rect 2534 2028 2580 2074
rect 2534 1919 2580 1965
rect 2534 1810 2580 1856
rect 2778 2138 2824 2184
rect 2778 2028 2824 2074
rect 2778 1919 2824 1965
rect 2778 1810 2824 1856
rect 3022 2138 3068 2184
rect 3022 2028 3068 2074
rect 3022 1919 3068 1965
rect 3022 1810 3068 1856
rect 3240 1949 3286 2097
rect 3240 1846 3286 1892
rect 872 1660 918 1706
rect 3240 1743 3286 1789
rect 3484 1949 3530 2097
rect 3484 1846 3530 1892
rect 3484 1743 3530 1789
rect 3728 1949 3774 2097
rect 3728 1846 3774 1892
rect 3728 1743 3774 1789
rect 4108 2101 4154 2147
rect 4108 1982 4154 2028
rect 4108 1863 4154 1909
rect 4108 1743 4154 1789
rect 4352 2101 4398 2147
rect 4352 1982 4398 2028
rect 4352 1863 4398 1909
rect 4352 1743 4398 1789
rect 4596 2101 4642 2147
rect 4596 1982 4642 2028
rect 4596 1863 4642 1909
rect 4596 1743 4642 1789
rect 4740 1949 4786 2097
rect 4740 1846 4786 1892
rect 4740 1743 4786 1789
rect 4984 1949 5030 2097
rect 4984 1846 5030 1892
rect 4984 1743 5030 1789
rect 5228 1949 5274 2097
rect 5228 1846 5274 1892
rect 5228 1743 5274 1789
rect 5756 1978 5802 2024
rect 5756 1868 5802 1914
rect 5756 1759 5802 1805
rect 5756 1650 5802 1696
rect 872 1556 918 1602
rect 6000 1978 6046 2024
rect 6000 1868 6046 1914
rect 6000 1759 6046 1805
rect 6000 1650 6046 1696
rect 6144 1978 6190 2024
rect 6144 1868 6190 1914
rect 6144 1759 6190 1805
rect 6144 1650 6190 1696
rect 6388 1978 6434 2024
rect 6388 1868 6434 1914
rect 6388 1759 6434 1805
rect 6388 1650 6434 1696
rect 872 1452 918 1498
rect 872 1348 918 1394
<< psubdiff >>
rect -1319 1008 19 1030
rect -1319 962 -1297 1008
rect -1251 962 -1193 1008
rect -1147 962 -1089 1008
rect -1043 962 -985 1008
rect -939 962 -881 1008
rect -835 962 -777 1008
rect -731 962 -673 1008
rect -627 962 -569 1008
rect -523 962 -465 1008
rect -419 962 -361 1008
rect -315 962 -257 1008
rect -211 962 -153 1008
rect -107 962 -49 1008
rect -3 962 19 1008
rect -1319 904 19 962
rect -1319 858 -1297 904
rect -1251 858 -1193 904
rect -1147 858 -1089 904
rect -1043 858 -985 904
rect -939 858 -881 904
rect -835 858 -777 904
rect -731 858 -673 904
rect -627 858 -569 904
rect -523 858 -465 904
rect -419 858 -361 904
rect -315 858 -257 904
rect -211 858 -153 904
rect -107 858 -49 904
rect -3 858 19 904
rect -1319 800 19 858
rect -1319 754 -1297 800
rect -1251 754 -1193 800
rect -1147 754 -1089 800
rect -1043 754 -985 800
rect -939 754 -881 800
rect -835 754 -777 800
rect -731 754 -673 800
rect -627 754 -569 800
rect -523 754 -465 800
rect -419 754 -361 800
rect -315 754 -257 800
rect -211 754 -153 800
rect -107 754 -49 800
rect -3 754 19 800
rect -1319 696 19 754
rect -1319 650 -1297 696
rect -1251 650 -1193 696
rect -1147 650 -1089 696
rect -1043 650 -985 696
rect -939 650 -881 696
rect -835 650 -777 696
rect -731 650 -673 696
rect -627 650 -569 696
rect -523 650 -465 696
rect -419 650 -361 696
rect -315 650 -257 696
rect -211 650 -153 696
rect -107 650 -49 696
rect -3 650 19 696
rect -1319 592 19 650
rect -1319 546 -1297 592
rect -1251 546 -1193 592
rect -1147 546 -1089 592
rect -1043 546 -985 592
rect -939 546 -881 592
rect -835 546 -777 592
rect -731 546 -673 592
rect -627 546 -569 592
rect -523 546 -465 592
rect -419 546 -361 592
rect -315 546 -257 592
rect -211 546 -153 592
rect -107 546 -49 592
rect -3 546 19 592
rect -1319 488 19 546
rect -1319 442 -1297 488
rect -1251 442 -1193 488
rect -1147 442 -1089 488
rect -1043 442 -985 488
rect -939 442 -881 488
rect -835 442 -777 488
rect -731 442 -673 488
rect -627 442 -569 488
rect -523 442 -465 488
rect -419 442 -361 488
rect -315 442 -257 488
rect -211 442 -153 488
rect -107 442 -49 488
rect -3 442 19 488
rect -1319 384 19 442
rect -1319 338 -1297 384
rect -1251 338 -1193 384
rect -1147 338 -1089 384
rect -1043 338 -985 384
rect -939 338 -881 384
rect -835 338 -777 384
rect -731 338 -673 384
rect -627 338 -569 384
rect -523 338 -465 384
rect -419 338 -361 384
rect -315 338 -257 384
rect -211 338 -153 384
rect -107 338 -49 384
rect -3 338 19 384
rect -1319 280 19 338
rect -1319 234 -1297 280
rect -1251 234 -1193 280
rect -1147 234 -1089 280
rect -1043 234 -985 280
rect -939 234 -881 280
rect -835 234 -777 280
rect -731 234 -673 280
rect -627 234 -569 280
rect -523 234 -465 280
rect -419 234 -361 280
rect -315 234 -257 280
rect -211 234 -153 280
rect -107 234 -49 280
rect -3 234 19 280
rect -1319 176 19 234
rect -1319 130 -1297 176
rect -1251 130 -1193 176
rect -1147 130 -1089 176
rect -1043 130 -985 176
rect -939 130 -881 176
rect -835 130 -777 176
rect -731 130 -673 176
rect -627 130 -569 176
rect -523 130 -465 176
rect -419 130 -361 176
rect -315 130 -257 176
rect -211 130 -153 176
rect -107 130 -49 176
rect -3 130 19 176
rect -1319 108 19 130
rect 83 1008 173 1030
rect 83 22 105 1008
rect 151 90 173 1008
rect 6699 1008 6789 1030
rect 6699 90 6721 1008
rect 151 68 6721 90
rect 151 22 269 68
rect 6613 22 6721 68
rect 6767 22 6789 1008
rect 83 0 6789 22
<< nsubdiff >>
rect -1319 2470 19 2492
rect -1319 2424 -1297 2470
rect -1251 2424 -1193 2470
rect -1147 2424 -1089 2470
rect -1043 2424 -985 2470
rect -939 2424 -881 2470
rect -835 2424 -777 2470
rect -731 2424 -673 2470
rect -627 2424 -569 2470
rect -523 2424 -465 2470
rect -419 2424 -361 2470
rect -315 2424 -257 2470
rect -211 2424 -153 2470
rect -107 2424 -49 2470
rect -3 2424 19 2470
rect -1319 2366 19 2424
rect -1319 2320 -1297 2366
rect -1251 2320 -1193 2366
rect -1147 2320 -1089 2366
rect -1043 2320 -985 2366
rect -939 2320 -881 2366
rect -835 2320 -777 2366
rect -731 2320 -673 2366
rect -627 2320 -569 2366
rect -523 2320 -465 2366
rect -419 2320 -361 2366
rect -315 2320 -257 2366
rect -211 2320 -153 2366
rect -107 2320 -49 2366
rect -3 2320 19 2366
rect -1319 2262 19 2320
rect -1319 2216 -1297 2262
rect -1251 2216 -1193 2262
rect -1147 2216 -1089 2262
rect -1043 2216 -985 2262
rect -939 2216 -881 2262
rect -835 2216 -777 2262
rect -731 2216 -673 2262
rect -627 2216 -569 2262
rect -523 2216 -465 2262
rect -419 2216 -361 2262
rect -315 2216 -257 2262
rect -211 2216 -153 2262
rect -107 2216 -49 2262
rect -3 2216 19 2262
rect -1319 2158 19 2216
rect -1319 2112 -1297 2158
rect -1251 2112 -1193 2158
rect -1147 2112 -1089 2158
rect -1043 2112 -985 2158
rect -939 2112 -881 2158
rect -835 2112 -777 2158
rect -731 2112 -673 2158
rect -627 2112 -569 2158
rect -523 2112 -465 2158
rect -419 2112 -361 2158
rect -315 2112 -257 2158
rect -211 2112 -153 2158
rect -107 2112 -49 2158
rect -3 2112 19 2158
rect -1319 2054 19 2112
rect -1319 2008 -1297 2054
rect -1251 2008 -1193 2054
rect -1147 2008 -1089 2054
rect -1043 2008 -985 2054
rect -939 2008 -881 2054
rect -835 2008 -777 2054
rect -731 2008 -673 2054
rect -627 2008 -569 2054
rect -523 2008 -465 2054
rect -419 2008 -361 2054
rect -315 2008 -257 2054
rect -211 2008 -153 2054
rect -107 2008 -49 2054
rect -3 2008 19 2054
rect -1319 1950 19 2008
rect -1319 1904 -1297 1950
rect -1251 1904 -1193 1950
rect -1147 1904 -1089 1950
rect -1043 1904 -985 1950
rect -939 1904 -881 1950
rect -835 1904 -777 1950
rect -731 1904 -673 1950
rect -627 1904 -569 1950
rect -523 1904 -465 1950
rect -419 1904 -361 1950
rect -315 1904 -257 1950
rect -211 1904 -153 1950
rect -107 1904 -49 1950
rect -3 1904 19 1950
rect -1319 1846 19 1904
rect -1319 1800 -1297 1846
rect -1251 1800 -1193 1846
rect -1147 1800 -1089 1846
rect -1043 1800 -985 1846
rect -939 1800 -881 1846
rect -835 1800 -777 1846
rect -731 1800 -673 1846
rect -627 1800 -569 1846
rect -523 1800 -465 1846
rect -419 1800 -361 1846
rect -315 1800 -257 1846
rect -211 1800 -153 1846
rect -107 1800 -49 1846
rect -3 1800 19 1846
rect -1319 1742 19 1800
rect -1319 1696 -1297 1742
rect -1251 1696 -1193 1742
rect -1147 1696 -1089 1742
rect -1043 1696 -985 1742
rect -939 1696 -881 1742
rect -835 1696 -777 1742
rect -731 1696 -673 1742
rect -627 1696 -569 1742
rect -523 1696 -465 1742
rect -419 1696 -361 1742
rect -315 1696 -257 1742
rect -211 1696 -153 1742
rect -107 1696 -49 1742
rect -3 1696 19 1742
rect -1319 1638 19 1696
rect -1319 1592 -1297 1638
rect -1251 1592 -1193 1638
rect -1147 1592 -1089 1638
rect -1043 1592 -985 1638
rect -939 1592 -881 1638
rect -835 1592 -777 1638
rect -731 1592 -673 1638
rect -627 1592 -569 1638
rect -523 1592 -465 1638
rect -419 1592 -361 1638
rect -315 1592 -257 1638
rect -211 1592 -153 1638
rect -107 1592 -49 1638
rect -3 1592 19 1638
rect -1319 1570 19 1592
rect 83 2470 6789 2492
rect 83 1484 105 2470
rect 151 2424 269 2470
rect 6613 2424 6721 2470
rect 151 2402 6721 2424
rect 151 1484 173 2402
rect 83 1462 173 1484
rect 6699 1484 6721 2402
rect 6767 1484 6789 2470
rect 6699 1462 6789 1484
<< psubdiffcont >>
rect -1297 962 -1251 1008
rect -1193 962 -1147 1008
rect -1089 962 -1043 1008
rect -985 962 -939 1008
rect -881 962 -835 1008
rect -777 962 -731 1008
rect -673 962 -627 1008
rect -569 962 -523 1008
rect -465 962 -419 1008
rect -361 962 -315 1008
rect -257 962 -211 1008
rect -153 962 -107 1008
rect -49 962 -3 1008
rect -1297 858 -1251 904
rect -1193 858 -1147 904
rect -1089 858 -1043 904
rect -985 858 -939 904
rect -881 858 -835 904
rect -777 858 -731 904
rect -673 858 -627 904
rect -569 858 -523 904
rect -465 858 -419 904
rect -361 858 -315 904
rect -257 858 -211 904
rect -153 858 -107 904
rect -49 858 -3 904
rect -1297 754 -1251 800
rect -1193 754 -1147 800
rect -1089 754 -1043 800
rect -985 754 -939 800
rect -881 754 -835 800
rect -777 754 -731 800
rect -673 754 -627 800
rect -569 754 -523 800
rect -465 754 -419 800
rect -361 754 -315 800
rect -257 754 -211 800
rect -153 754 -107 800
rect -49 754 -3 800
rect -1297 650 -1251 696
rect -1193 650 -1147 696
rect -1089 650 -1043 696
rect -985 650 -939 696
rect -881 650 -835 696
rect -777 650 -731 696
rect -673 650 -627 696
rect -569 650 -523 696
rect -465 650 -419 696
rect -361 650 -315 696
rect -257 650 -211 696
rect -153 650 -107 696
rect -49 650 -3 696
rect -1297 546 -1251 592
rect -1193 546 -1147 592
rect -1089 546 -1043 592
rect -985 546 -939 592
rect -881 546 -835 592
rect -777 546 -731 592
rect -673 546 -627 592
rect -569 546 -523 592
rect -465 546 -419 592
rect -361 546 -315 592
rect -257 546 -211 592
rect -153 546 -107 592
rect -49 546 -3 592
rect -1297 442 -1251 488
rect -1193 442 -1147 488
rect -1089 442 -1043 488
rect -985 442 -939 488
rect -881 442 -835 488
rect -777 442 -731 488
rect -673 442 -627 488
rect -569 442 -523 488
rect -465 442 -419 488
rect -361 442 -315 488
rect -257 442 -211 488
rect -153 442 -107 488
rect -49 442 -3 488
rect -1297 338 -1251 384
rect -1193 338 -1147 384
rect -1089 338 -1043 384
rect -985 338 -939 384
rect -881 338 -835 384
rect -777 338 -731 384
rect -673 338 -627 384
rect -569 338 -523 384
rect -465 338 -419 384
rect -361 338 -315 384
rect -257 338 -211 384
rect -153 338 -107 384
rect -49 338 -3 384
rect -1297 234 -1251 280
rect -1193 234 -1147 280
rect -1089 234 -1043 280
rect -985 234 -939 280
rect -881 234 -835 280
rect -777 234 -731 280
rect -673 234 -627 280
rect -569 234 -523 280
rect -465 234 -419 280
rect -361 234 -315 280
rect -257 234 -211 280
rect -153 234 -107 280
rect -49 234 -3 280
rect -1297 130 -1251 176
rect -1193 130 -1147 176
rect -1089 130 -1043 176
rect -985 130 -939 176
rect -881 130 -835 176
rect -777 130 -731 176
rect -673 130 -627 176
rect -569 130 -523 176
rect -465 130 -419 176
rect -361 130 -315 176
rect -257 130 -211 176
rect -153 130 -107 176
rect -49 130 -3 176
rect 105 22 151 1008
rect 269 22 6613 68
rect 6721 22 6767 1008
<< nsubdiffcont >>
rect -1297 2424 -1251 2470
rect -1193 2424 -1147 2470
rect -1089 2424 -1043 2470
rect -985 2424 -939 2470
rect -881 2424 -835 2470
rect -777 2424 -731 2470
rect -673 2424 -627 2470
rect -569 2424 -523 2470
rect -465 2424 -419 2470
rect -361 2424 -315 2470
rect -257 2424 -211 2470
rect -153 2424 -107 2470
rect -49 2424 -3 2470
rect -1297 2320 -1251 2366
rect -1193 2320 -1147 2366
rect -1089 2320 -1043 2366
rect -985 2320 -939 2366
rect -881 2320 -835 2366
rect -777 2320 -731 2366
rect -673 2320 -627 2366
rect -569 2320 -523 2366
rect -465 2320 -419 2366
rect -361 2320 -315 2366
rect -257 2320 -211 2366
rect -153 2320 -107 2366
rect -49 2320 -3 2366
rect -1297 2216 -1251 2262
rect -1193 2216 -1147 2262
rect -1089 2216 -1043 2262
rect -985 2216 -939 2262
rect -881 2216 -835 2262
rect -777 2216 -731 2262
rect -673 2216 -627 2262
rect -569 2216 -523 2262
rect -465 2216 -419 2262
rect -361 2216 -315 2262
rect -257 2216 -211 2262
rect -153 2216 -107 2262
rect -49 2216 -3 2262
rect -1297 2112 -1251 2158
rect -1193 2112 -1147 2158
rect -1089 2112 -1043 2158
rect -985 2112 -939 2158
rect -881 2112 -835 2158
rect -777 2112 -731 2158
rect -673 2112 -627 2158
rect -569 2112 -523 2158
rect -465 2112 -419 2158
rect -361 2112 -315 2158
rect -257 2112 -211 2158
rect -153 2112 -107 2158
rect -49 2112 -3 2158
rect -1297 2008 -1251 2054
rect -1193 2008 -1147 2054
rect -1089 2008 -1043 2054
rect -985 2008 -939 2054
rect -881 2008 -835 2054
rect -777 2008 -731 2054
rect -673 2008 -627 2054
rect -569 2008 -523 2054
rect -465 2008 -419 2054
rect -361 2008 -315 2054
rect -257 2008 -211 2054
rect -153 2008 -107 2054
rect -49 2008 -3 2054
rect -1297 1904 -1251 1950
rect -1193 1904 -1147 1950
rect -1089 1904 -1043 1950
rect -985 1904 -939 1950
rect -881 1904 -835 1950
rect -777 1904 -731 1950
rect -673 1904 -627 1950
rect -569 1904 -523 1950
rect -465 1904 -419 1950
rect -361 1904 -315 1950
rect -257 1904 -211 1950
rect -153 1904 -107 1950
rect -49 1904 -3 1950
rect -1297 1800 -1251 1846
rect -1193 1800 -1147 1846
rect -1089 1800 -1043 1846
rect -985 1800 -939 1846
rect -881 1800 -835 1846
rect -777 1800 -731 1846
rect -673 1800 -627 1846
rect -569 1800 -523 1846
rect -465 1800 -419 1846
rect -361 1800 -315 1846
rect -257 1800 -211 1846
rect -153 1800 -107 1846
rect -49 1800 -3 1846
rect -1297 1696 -1251 1742
rect -1193 1696 -1147 1742
rect -1089 1696 -1043 1742
rect -985 1696 -939 1742
rect -881 1696 -835 1742
rect -777 1696 -731 1742
rect -673 1696 -627 1742
rect -569 1696 -523 1742
rect -465 1696 -419 1742
rect -361 1696 -315 1742
rect -257 1696 -211 1742
rect -153 1696 -107 1742
rect -49 1696 -3 1742
rect -1297 1592 -1251 1638
rect -1193 1592 -1147 1638
rect -1089 1592 -1043 1638
rect -985 1592 -939 1638
rect -881 1592 -835 1638
rect -777 1592 -731 1638
rect -673 1592 -627 1638
rect -569 1592 -523 1638
rect -465 1592 -419 1638
rect -361 1592 -315 1638
rect -257 1592 -211 1638
rect -153 1592 -107 1638
rect -49 1592 -3 1638
rect 105 1484 151 2470
rect 269 2424 6613 2470
rect 6721 1484 6767 2470
<< polysilicon >>
rect 2365 2197 2505 2241
rect 2609 2197 2749 2241
rect 2853 2197 2993 2241
rect 459 2135 599 2179
rect 703 2135 843 2179
rect 1669 2097 1809 2141
rect 1913 2097 2053 2141
rect 4183 2160 4323 2204
rect 4427 2160 4567 2204
rect 3315 2110 3455 2154
rect 3559 2110 3699 2154
rect 1669 1644 1809 1797
rect 1913 1644 2053 1797
rect 2365 1644 2505 1797
rect 2609 1644 2749 1797
rect 2853 1644 2993 1797
rect 4815 2110 4955 2154
rect 5059 2110 5199 2154
rect 5831 2037 5971 2081
rect 6219 2037 6359 2081
rect 3315 1644 3455 1730
rect 3559 1644 3699 1730
rect 4183 1644 4323 1730
rect 4427 1644 4567 1730
rect 4815 1644 4955 1730
rect 5059 1644 5199 1730
rect 1650 1625 1828 1644
rect 1650 1579 1669 1625
rect 1809 1579 1828 1625
rect 1650 1560 1828 1579
rect 1894 1625 2072 1644
rect 1894 1579 1913 1625
rect 2053 1579 2072 1625
rect 1894 1560 2072 1579
rect 2346 1625 2524 1644
rect 2346 1579 2365 1625
rect 2505 1579 2524 1625
rect 2346 1560 2524 1579
rect 2590 1625 2768 1644
rect 2590 1579 2609 1625
rect 2749 1579 2768 1625
rect 2590 1560 2768 1579
rect 2834 1625 3012 1644
rect 2834 1579 2853 1625
rect 2993 1579 3012 1625
rect 2834 1560 3012 1579
rect 3296 1625 3474 1644
rect 3296 1579 3315 1625
rect 3455 1579 3474 1625
rect 3296 1560 3474 1579
rect 3540 1625 3718 1644
rect 3540 1579 3559 1625
rect 3699 1579 3718 1625
rect 3540 1560 3718 1579
rect 4164 1625 4342 1644
rect 4164 1579 4183 1625
rect 4323 1579 4342 1625
rect 4164 1560 4342 1579
rect 4408 1625 4586 1644
rect 4408 1579 4427 1625
rect 4567 1579 4586 1625
rect 4408 1560 4586 1579
rect 4796 1625 4974 1644
rect 4796 1579 4815 1625
rect 4955 1579 4974 1625
rect 4796 1560 4974 1579
rect 5040 1625 5218 1644
rect 5040 1579 5059 1625
rect 5199 1579 5218 1625
rect 5040 1560 5218 1579
rect 5831 1528 5971 1637
rect 6219 1528 6359 1637
rect 5812 1509 5990 1528
rect 5812 1463 5831 1509
rect 5971 1463 5990 1509
rect 5812 1444 5990 1463
rect 6200 1509 6378 1528
rect 6200 1463 6219 1509
rect 6359 1463 6378 1509
rect 6200 1444 6378 1463
rect 459 1027 599 1335
rect 459 887 506 1027
rect 552 887 599 1027
rect 459 680 599 887
rect 703 1027 843 1335
rect 5812 1213 5990 1232
rect 5812 1167 5831 1213
rect 5971 1167 5990 1213
rect 5812 1148 5990 1167
rect 6200 1213 6378 1232
rect 6200 1167 6219 1213
rect 6359 1167 6378 1213
rect 6200 1148 6378 1167
rect 1151 1101 1329 1120
rect 1151 1055 1170 1101
rect 1310 1055 1329 1101
rect 1151 1036 1329 1055
rect 1728 1101 1906 1120
rect 1728 1055 1747 1101
rect 1887 1055 1906 1101
rect 1728 1036 1906 1055
rect 1972 1101 2150 1120
rect 1972 1055 1991 1101
rect 2131 1055 2150 1101
rect 1972 1036 2150 1055
rect 2216 1101 2394 1120
rect 2216 1055 2235 1101
rect 2375 1055 2394 1101
rect 2216 1036 2394 1055
rect 2460 1101 2638 1120
rect 2460 1055 2479 1101
rect 2619 1055 2638 1101
rect 2460 1036 2638 1055
rect 2704 1101 2882 1120
rect 2704 1055 2723 1101
rect 2863 1055 2882 1101
rect 2704 1036 2882 1055
rect 3184 1101 3362 1120
rect 3184 1055 3203 1101
rect 3343 1055 3362 1101
rect 3184 1036 3362 1055
rect 3428 1101 3606 1120
rect 3428 1055 3447 1101
rect 3587 1055 3606 1101
rect 3428 1036 3606 1055
rect 3672 1101 3850 1120
rect 3672 1055 3691 1101
rect 3831 1055 3850 1101
rect 3672 1036 3850 1055
rect 3916 1101 4094 1120
rect 3916 1055 3935 1101
rect 4075 1055 4094 1101
rect 3916 1036 4094 1055
rect 4304 1101 4482 1120
rect 4304 1055 4323 1101
rect 4463 1055 4482 1101
rect 4304 1036 4482 1055
rect 4548 1101 4726 1120
rect 4548 1055 4567 1101
rect 4707 1055 4726 1101
rect 4548 1036 4726 1055
rect 4792 1101 4970 1120
rect 4792 1055 4811 1101
rect 4951 1055 4970 1101
rect 4792 1036 4970 1055
rect 5036 1101 5214 1120
rect 5036 1055 5055 1101
rect 5195 1055 5214 1101
rect 5036 1036 5214 1055
rect 703 887 750 1027
rect 796 887 843 1027
rect 1170 920 1310 1036
rect 1747 920 1887 1036
rect 1991 920 2131 1036
rect 2235 920 2375 1036
rect 2479 920 2619 1036
rect 2723 920 2863 1036
rect 703 680 843 887
rect 1170 576 1310 620
rect 3203 868 3343 1036
rect 3447 868 3587 1036
rect 3691 868 3831 1036
rect 3935 868 4075 1036
rect 4323 868 4463 1036
rect 4567 868 4707 1036
rect 4811 868 4951 1036
rect 5055 868 5195 1036
rect 5831 1031 5971 1148
rect 6219 1031 6359 1148
rect 5443 868 5583 912
rect 3203 294 3343 338
rect 3447 294 3587 338
rect 3691 294 3831 338
rect 3935 294 4075 338
rect 459 236 599 280
rect 703 236 843 280
rect 1747 236 1887 280
rect 1991 236 2131 280
rect 2235 236 2375 280
rect 2479 236 2619 280
rect 2723 236 2863 280
rect 5831 687 5971 731
rect 6219 687 6359 731
rect 5443 513 5583 608
rect 5443 494 5621 513
rect 5443 448 5462 494
rect 5602 448 5621 494
rect 5443 429 5621 448
rect 4323 224 4463 268
rect 4567 224 4707 268
rect 4811 224 4951 268
rect 5055 224 5195 268
<< polycontact >>
rect 1669 1579 1809 1625
rect 1913 1579 2053 1625
rect 2365 1579 2505 1625
rect 2609 1579 2749 1625
rect 2853 1579 2993 1625
rect 3315 1579 3455 1625
rect 3559 1579 3699 1625
rect 4183 1579 4323 1625
rect 4427 1579 4567 1625
rect 4815 1579 4955 1625
rect 5059 1579 5199 1625
rect 5831 1463 5971 1509
rect 6219 1463 6359 1509
rect 506 887 552 1027
rect 5831 1167 5971 1213
rect 6219 1167 6359 1213
rect 1170 1055 1310 1101
rect 1747 1055 1887 1101
rect 1991 1055 2131 1101
rect 2235 1055 2375 1101
rect 2479 1055 2619 1101
rect 2723 1055 2863 1101
rect 3203 1055 3343 1101
rect 3447 1055 3587 1101
rect 3691 1055 3831 1101
rect 3935 1055 4075 1101
rect 4323 1055 4463 1101
rect 4567 1055 4707 1101
rect 4811 1055 4951 1101
rect 5055 1055 5195 1101
rect 750 887 796 1027
rect 5462 448 5602 494
<< metal1 >>
rect 8 2481 148 2489
rect -1308 2470 6778 2481
rect -1308 2424 -1297 2470
rect -1251 2424 -1193 2470
rect -1147 2424 -1089 2470
rect -1043 2424 -985 2470
rect -939 2424 -881 2470
rect -835 2424 -777 2470
rect -731 2424 -673 2470
rect -627 2424 -569 2470
rect -523 2424 -465 2470
rect -419 2424 -361 2470
rect -315 2424 -257 2470
rect -211 2424 -153 2470
rect -107 2424 -49 2470
rect -3 2424 105 2470
rect -1308 2366 105 2424
rect -1308 2320 -1297 2366
rect -1251 2320 -1193 2366
rect -1147 2320 -1089 2366
rect -1043 2320 -985 2366
rect -939 2320 -881 2366
rect -835 2320 -777 2366
rect -731 2320 -673 2366
rect -627 2320 -569 2366
rect -523 2320 -465 2366
rect -419 2320 -361 2366
rect -315 2320 -257 2366
rect -211 2320 -153 2366
rect -107 2320 -49 2366
rect -3 2320 105 2366
rect -1308 2262 105 2320
rect -1308 2216 -1297 2262
rect -1251 2216 -1193 2262
rect -1147 2216 -1089 2262
rect -1043 2216 -985 2262
rect -939 2216 -881 2262
rect -835 2216 -777 2262
rect -731 2216 -673 2262
rect -627 2216 -569 2262
rect -523 2216 -465 2262
rect -419 2216 -361 2262
rect -315 2216 -257 2262
rect -211 2216 -153 2262
rect -107 2216 -49 2262
rect -3 2216 105 2262
rect -1308 2158 105 2216
rect -1308 2112 -1297 2158
rect -1251 2112 -1193 2158
rect -1147 2112 -1089 2158
rect -1043 2112 -985 2158
rect -939 2112 -881 2158
rect -835 2112 -777 2158
rect -731 2112 -673 2158
rect -627 2112 -569 2158
rect -523 2112 -465 2158
rect -419 2112 -361 2158
rect -315 2112 -257 2158
rect -211 2112 -153 2158
rect -107 2112 -49 2158
rect -3 2112 105 2158
rect -1308 2054 105 2112
rect -1308 2008 -1297 2054
rect -1251 2008 -1193 2054
rect -1147 2008 -1089 2054
rect -1043 2008 -985 2054
rect -939 2008 -881 2054
rect -835 2008 -777 2054
rect -731 2008 -673 2054
rect -627 2008 -569 2054
rect -523 2008 -465 2054
rect -419 2008 -361 2054
rect -315 2008 -257 2054
rect -211 2008 -153 2054
rect -107 2008 -49 2054
rect -3 2008 105 2054
rect -1308 1950 105 2008
rect -1308 1904 -1297 1950
rect -1251 1904 -1193 1950
rect -1147 1904 -1089 1950
rect -1043 1904 -985 1950
rect -939 1904 -881 1950
rect -835 1904 -777 1950
rect -731 1904 -673 1950
rect -627 1904 -569 1950
rect -523 1904 -465 1950
rect -419 1904 -361 1950
rect -315 1904 -257 1950
rect -211 1904 -153 1950
rect -107 1904 -49 1950
rect -3 1904 105 1950
rect -1308 1846 105 1904
rect -1308 1800 -1297 1846
rect -1251 1800 -1193 1846
rect -1147 1800 -1089 1846
rect -1043 1800 -985 1846
rect -939 1800 -881 1846
rect -835 1800 -777 1846
rect -731 1800 -673 1846
rect -627 1800 -569 1846
rect -523 1800 -465 1846
rect -419 1800 -361 1846
rect -315 1800 -257 1846
rect -211 1800 -153 1846
rect -107 1800 -49 1846
rect -3 1800 105 1846
rect -1308 1742 105 1800
rect -1308 1696 -1297 1742
rect -1251 1696 -1193 1742
rect -1147 1696 -1089 1742
rect -1043 1696 -985 1742
rect -939 1696 -881 1742
rect -835 1696 -777 1742
rect -731 1696 -673 1742
rect -627 1696 -569 1742
rect -523 1696 -465 1742
rect -419 1696 -361 1742
rect -315 1696 -257 1742
rect -211 1696 -153 1742
rect -107 1696 -49 1742
rect -3 1696 105 1742
rect -1308 1638 105 1696
rect -1308 1592 -1297 1638
rect -1251 1592 -1193 1638
rect -1147 1592 -1089 1638
rect -1043 1592 -985 1638
rect -939 1592 -881 1638
rect -835 1592 -777 1638
rect -731 1592 -673 1638
rect -627 1592 -569 1638
rect -523 1592 -465 1638
rect -419 1592 -361 1638
rect -315 1592 -257 1638
rect -211 1592 -153 1638
rect -107 1592 -49 1638
rect -3 1592 105 1638
rect -1308 1581 105 1592
rect 94 1484 105 1581
rect 151 2424 269 2470
rect 6613 2424 6721 2470
rect 151 2413 6721 2424
rect 151 1484 162 2413
rect 94 1473 162 1484
rect 384 2122 430 2413
rect 384 2018 430 2076
rect 384 1914 430 1972
rect 384 1810 430 1868
rect 384 1706 430 1764
rect 384 1602 430 1660
rect 384 1498 430 1556
rect 384 1394 430 1452
rect 384 1335 430 1348
rect 613 2122 689 2135
rect 613 2076 628 2122
rect 674 2076 689 2122
rect 613 2018 689 2076
rect 613 1972 628 2018
rect 674 1972 689 2018
rect 613 1914 689 1972
rect 613 1868 628 1914
rect 674 1868 689 1914
rect 613 1810 689 1868
rect 613 1764 628 1810
rect 674 1764 689 1810
rect 613 1706 689 1764
rect 613 1660 628 1706
rect 674 1660 689 1706
rect 613 1602 689 1660
rect 613 1556 628 1602
rect 674 1556 689 1602
rect 613 1498 689 1556
rect 613 1452 628 1498
rect 674 1452 689 1498
rect 613 1394 689 1452
rect 613 1348 628 1394
rect 674 1348 689 1394
rect 613 1224 689 1348
rect 872 2122 918 2413
rect 872 2018 918 2076
rect 872 1914 918 1972
rect 872 1810 918 1868
rect 1594 2084 1640 2413
rect 1594 1970 1640 2038
rect 1838 2084 1884 2097
rect 1838 1977 1884 2038
rect 2082 2084 2128 2413
rect 1594 1856 1640 1924
rect 1594 1797 1640 1810
rect 1823 1970 1899 1977
rect 1823 1965 1838 1970
rect 1884 1965 1899 1970
rect 1823 1809 1835 1965
rect 1887 1809 1899 1965
rect 1823 1797 1899 1809
rect 2082 1970 2128 2038
rect 2082 1856 2128 1924
rect 2082 1797 2128 1810
rect 2290 2184 2346 2413
rect 2336 2138 2346 2184
rect 2290 2074 2346 2138
rect 2336 2028 2346 2074
rect 2290 1965 2346 2028
rect 2336 1919 2346 1965
rect 2290 1856 2346 1919
rect 2336 1810 2346 1856
rect 872 1706 918 1764
rect 2290 1745 2346 1810
rect 2528 2301 3072 2357
rect 2528 2184 2584 2301
rect 2528 2138 2534 2184
rect 2580 2138 2584 2184
rect 2528 2074 2584 2138
rect 2528 2028 2534 2074
rect 2580 2028 2584 2074
rect 2528 1965 2584 2028
rect 2528 1919 2534 1965
rect 2580 1919 2584 1965
rect 2528 1856 2584 1919
rect 2528 1810 2534 1856
rect 2580 1810 2584 1856
rect 2528 1797 2584 1810
rect 2773 2184 2829 2197
rect 2773 2138 2778 2184
rect 2824 2138 2829 2184
rect 2773 2074 2829 2138
rect 2773 2028 2778 2074
rect 2824 2028 2829 2074
rect 2773 1965 2829 2028
rect 2773 1919 2778 1965
rect 2824 1919 2829 1965
rect 2773 1856 2829 1919
rect 3016 2184 3072 2301
rect 3016 2138 3022 2184
rect 3068 2138 3072 2184
rect 3016 2074 3072 2138
rect 3016 2028 3022 2074
rect 3068 2028 3072 2074
rect 3016 1965 3072 2028
rect 3016 1919 3022 1965
rect 3068 1919 3072 1965
rect 3016 1910 3072 1919
rect 3227 2210 3303 2222
rect 3227 2054 3239 2210
rect 3291 2054 3303 2210
rect 3227 1949 3240 2054
rect 3286 1949 3303 2054
rect 2773 1810 2778 1856
rect 2824 1810 2829 1856
rect 2773 1745 2829 1810
rect 2290 1689 2829 1745
rect 3006 1898 3082 1910
rect 3006 1742 3018 1898
rect 3070 1742 3082 1898
rect 3006 1730 3082 1742
rect 3227 1892 3303 1949
rect 3227 1846 3240 1892
rect 3286 1846 3303 1892
rect 3227 1789 3303 1846
rect 3227 1743 3240 1789
rect 3286 1743 3303 1789
rect 3227 1730 3303 1743
rect 3469 2097 3545 2413
rect 4979 2285 6620 2341
rect 3601 2254 4171 2266
rect 3601 2202 3613 2254
rect 3769 2202 4171 2254
rect 3601 2190 4171 2202
rect 4095 2147 4171 2190
rect 4095 2110 4108 2147
rect 3469 1949 3484 2097
rect 3530 1949 3545 2097
rect 3469 1892 3545 1949
rect 3469 1846 3484 1892
rect 3530 1846 3545 1892
rect 3469 1789 3545 1846
rect 3469 1743 3484 1789
rect 3530 1743 3545 1789
rect 3469 1730 3545 1743
rect 3728 2106 4108 2110
rect 4154 2106 4171 2147
rect 3728 2097 4107 2106
rect 3774 1950 4107 2097
rect 4159 1950 4171 2106
rect 3774 1949 4171 1950
rect 3728 1909 4171 1949
rect 4352 2147 4398 2160
rect 4352 2028 4398 2101
rect 4352 1910 4398 1982
rect 4579 2147 4655 2206
rect 4579 2106 4596 2147
rect 4642 2110 4655 2147
rect 4642 2106 4786 2110
rect 4579 1950 4591 2106
rect 4643 2097 4786 2106
rect 4643 1950 4740 2097
rect 4579 1949 4740 1950
rect 3728 1892 4108 1909
rect 3774 1863 4108 1892
rect 4154 1863 4171 1909
rect 3774 1846 4171 1863
rect 3728 1789 4171 1846
rect 3774 1743 4108 1789
rect 4154 1743 4171 1789
rect 3728 1730 4171 1743
rect 4337 1909 4413 1910
rect 4337 1898 4352 1909
rect 4398 1898 4413 1909
rect 4337 1742 4349 1898
rect 4401 1742 4413 1898
rect 4337 1730 4413 1742
rect 4579 1909 4786 1949
rect 4579 1863 4596 1909
rect 4642 1892 4786 1909
rect 4642 1863 4740 1892
rect 4579 1846 4740 1863
rect 4579 1789 4786 1846
rect 4579 1743 4596 1789
rect 4642 1743 4740 1789
rect 4979 2097 5035 2285
rect 4979 1949 4984 2097
rect 5030 1949 5035 2097
rect 4979 1892 5035 1949
rect 4979 1846 4984 1892
rect 5030 1846 5035 1892
rect 4979 1789 5035 1846
rect 4979 1766 4984 1789
rect 4579 1730 4786 1743
rect 5030 1766 5035 1789
rect 5203 2106 5279 2118
rect 5203 1950 5215 2106
rect 5267 2097 5279 2106
rect 5203 1949 5228 1950
rect 5274 1949 5279 2097
rect 5203 1892 5279 1949
rect 5203 1846 5228 1892
rect 5274 1846 5279 1892
rect 5203 1789 5279 1846
rect 4984 1730 5030 1743
rect 5203 1743 5228 1789
rect 5274 1743 5279 1789
rect 5203 1730 5279 1743
rect 5741 2024 5817 2037
rect 5741 1978 5756 2024
rect 5802 1978 5817 2024
rect 5741 1914 5817 1978
rect 5741 1868 5756 1914
rect 5802 1868 5817 1914
rect 5741 1805 5817 1868
rect 5741 1804 5756 1805
rect 5802 1804 5817 1805
rect 872 1602 918 1660
rect 5741 1648 5753 1804
rect 5805 1648 5817 1804
rect 3876 1636 4056 1644
rect 5741 1636 5817 1648
rect 6000 2024 6190 2037
rect 6046 1978 6144 2024
rect 6000 1914 6190 1978
rect 6046 1868 6144 1914
rect 6000 1805 6190 1868
rect 6388 2024 6434 2037
rect 6388 1914 6434 1978
rect 6388 1817 6434 1868
rect 6000 1696 6017 1759
rect 6173 1696 6190 1759
rect 6000 1649 6017 1650
rect 6173 1649 6190 1650
rect 6000 1637 6190 1649
rect 6373 1805 6449 1817
rect 6373 1649 6385 1805
rect 6437 1649 6449 1805
rect 6564 1793 6620 2285
rect 6373 1637 6449 1649
rect 6554 1781 6630 1793
rect 872 1498 918 1556
rect 1492 1625 2064 1636
rect 1492 1579 1669 1625
rect 1809 1579 1913 1625
rect 2053 1579 2064 1625
rect 1492 1568 2064 1579
rect 2354 1625 3004 1636
rect 2354 1579 2365 1625
rect 2505 1579 2609 1625
rect 2749 1624 2853 1625
rect 2779 1579 2853 1624
rect 2993 1579 3004 1625
rect 2354 1572 2623 1579
rect 2779 1572 3004 1579
rect 2354 1568 3004 1572
rect 3304 1632 4578 1636
rect 3304 1625 3888 1632
rect 3304 1579 3315 1625
rect 3455 1579 3559 1625
rect 3699 1580 3888 1625
rect 4044 1625 4578 1632
rect 4044 1580 4183 1625
rect 3699 1579 4183 1580
rect 4323 1579 4427 1625
rect 4567 1579 4578 1625
rect 3304 1568 4578 1579
rect 4804 1625 5817 1636
rect 4804 1579 4815 1625
rect 4955 1579 5059 1625
rect 5199 1579 5817 1625
rect 6554 1625 6566 1781
rect 6618 1625 6630 1781
rect 6554 1613 6630 1625
rect 4804 1568 5817 1579
rect 872 1394 918 1452
rect 872 1335 918 1348
rect 1142 1506 1322 1518
rect 1142 1454 1154 1506
rect 1310 1454 1322 1506
rect 1142 1442 1322 1454
rect 1142 1224 1240 1442
rect 1492 1244 1560 1568
rect 2611 1560 2791 1568
rect 1640 1508 1820 1518
rect 5820 1509 6370 1520
rect 5820 1508 5831 1509
rect 1640 1506 5831 1508
rect 1640 1454 1652 1506
rect 1808 1463 5831 1506
rect 5971 1463 6219 1509
rect 6359 1508 6370 1509
rect 6359 1463 6472 1508
rect 6710 1484 6721 2413
rect 6767 1484 6778 2470
rect 6710 1473 6778 1484
rect 1808 1454 6472 1463
rect 1640 1452 6472 1454
rect 1640 1442 1820 1452
rect 2954 1364 6472 1396
rect 2954 1363 4361 1364
rect 2954 1311 2966 1363
rect 3122 1312 4361 1363
rect 4517 1312 4873 1364
rect 5029 1312 6017 1364
rect 6173 1312 6472 1364
rect 3122 1311 6472 1312
rect 2954 1280 6472 1311
rect 1492 1232 1672 1244
rect 613 1168 1321 1224
rect 1492 1180 1504 1232
rect 1660 1224 1672 1232
rect 1660 1213 6472 1224
rect 1660 1180 5831 1213
rect 1492 1168 5831 1180
rect 495 1027 811 1038
rect -1308 1008 162 1019
rect -1308 962 -1297 1008
rect -1251 962 -1193 1008
rect -1147 962 -1089 1008
rect -1043 962 -985 1008
rect -939 962 -881 1008
rect -835 962 -777 1008
rect -731 962 -673 1008
rect -627 962 -569 1008
rect -523 962 -465 1008
rect -419 962 -361 1008
rect -315 962 -257 1008
rect -211 962 -153 1008
rect -107 962 -49 1008
rect -3 962 105 1008
rect -1308 904 105 962
rect -1308 858 -1297 904
rect -1251 858 -1193 904
rect -1147 858 -1089 904
rect -1043 858 -985 904
rect -939 858 -881 904
rect -835 858 -777 904
rect -731 858 -673 904
rect -627 858 -569 904
rect -523 858 -465 904
rect -419 858 -361 904
rect -315 858 -257 904
rect -211 858 -153 904
rect -107 858 -49 904
rect -3 858 105 904
rect -1308 800 105 858
rect -1308 754 -1297 800
rect -1251 754 -1193 800
rect -1147 754 -1089 800
rect -1043 754 -985 800
rect -939 754 -881 800
rect -835 754 -777 800
rect -731 754 -673 800
rect -627 754 -569 800
rect -523 754 -465 800
rect -419 754 -361 800
rect -315 754 -257 800
rect -211 754 -153 800
rect -107 754 -49 800
rect -3 754 105 800
rect -1308 696 105 754
rect -1308 650 -1297 696
rect -1251 650 -1193 696
rect -1147 650 -1089 696
rect -1043 650 -985 696
rect -939 650 -881 696
rect -835 650 -777 696
rect -731 650 -673 696
rect -627 650 -569 696
rect -523 650 -465 696
rect -419 650 -361 696
rect -315 650 -257 696
rect -211 650 -153 696
rect -107 650 -49 696
rect -3 650 105 696
rect -1308 592 105 650
rect -1308 546 -1297 592
rect -1251 546 -1193 592
rect -1147 546 -1089 592
rect -1043 546 -985 592
rect -939 546 -881 592
rect -835 546 -777 592
rect -731 546 -673 592
rect -627 546 -569 592
rect -523 546 -465 592
rect -419 546 -361 592
rect -315 546 -257 592
rect -211 546 -153 592
rect -107 546 -49 592
rect -3 546 105 592
rect -1308 488 105 546
rect -1308 442 -1297 488
rect -1251 442 -1193 488
rect -1147 442 -1089 488
rect -1043 442 -985 488
rect -939 442 -881 488
rect -835 442 -777 488
rect -731 442 -673 488
rect -627 442 -569 488
rect -523 442 -465 488
rect -419 442 -361 488
rect -315 442 -257 488
rect -211 442 -153 488
rect -107 442 -49 488
rect -3 442 105 488
rect -1308 384 105 442
rect -1308 338 -1297 384
rect -1251 338 -1193 384
rect -1147 338 -1089 384
rect -1043 338 -985 384
rect -939 338 -881 384
rect -835 338 -777 384
rect -731 338 -673 384
rect -627 338 -569 384
rect -523 338 -465 384
rect -419 338 -361 384
rect -315 338 -257 384
rect -211 338 -153 384
rect -107 338 -49 384
rect -3 338 105 384
rect -1308 280 105 338
rect -1308 234 -1297 280
rect -1251 234 -1193 280
rect -1147 234 -1089 280
rect -1043 234 -985 280
rect -939 234 -881 280
rect -835 234 -777 280
rect -731 234 -673 280
rect -627 234 -569 280
rect -523 234 -465 280
rect -419 234 -361 280
rect -315 234 -257 280
rect -211 234 -153 280
rect -107 234 -49 280
rect -3 234 105 280
rect -1308 176 105 234
rect -1308 130 -1297 176
rect -1251 130 -1193 176
rect -1147 130 -1089 176
rect -1043 130 -985 176
rect -939 130 -881 176
rect -835 130 -777 176
rect -731 130 -673 176
rect -627 130 -569 176
rect -523 130 -465 176
rect -419 130 -361 176
rect -315 130 -257 176
rect -211 130 -153 176
rect -107 130 -49 176
rect -3 130 105 176
rect -1308 119 105 130
rect 8 22 105 119
rect 151 79 162 1008
rect 495 887 506 1027
rect 552 982 750 1027
rect 552 930 630 982
rect 552 887 750 930
rect 796 887 811 1027
rect 495 876 811 887
rect 905 826 981 1168
rect 1159 1101 1321 1168
rect 5820 1167 5831 1168
rect 5971 1167 6219 1213
rect 6359 1168 6472 1213
rect 6359 1167 6370 1168
rect 5820 1156 6370 1167
rect 4016 1112 4196 1120
rect 1159 1055 1170 1101
rect 1310 1055 1321 1101
rect 1159 1044 1321 1055
rect 1508 1101 2874 1112
rect 1508 1055 1747 1101
rect 1887 1055 1991 1101
rect 2131 1055 2235 1101
rect 2375 1055 2479 1101
rect 2619 1100 2723 1101
rect 2619 1055 2623 1100
rect 2863 1055 2874 1101
rect 1508 1048 2623 1055
rect 2779 1048 2874 1055
rect 1508 1044 2874 1048
rect 3192 1108 5206 1112
rect 3192 1101 4028 1108
rect 4184 1101 5206 1108
rect 3192 1055 3203 1101
rect 3343 1055 3447 1101
rect 3587 1055 3691 1101
rect 3831 1055 3935 1101
rect 4184 1056 4323 1101
rect 4075 1055 4323 1056
rect 4463 1055 4567 1101
rect 4707 1055 4811 1101
rect 4951 1055 5055 1101
rect 5195 1055 5206 1101
rect 3192 1044 5206 1055
rect 615 750 981 826
rect 1095 907 1141 920
rect 1095 793 1141 861
rect 384 667 430 680
rect 384 558 430 621
rect 384 449 430 512
rect 384 339 430 403
rect 384 79 430 293
rect 615 667 687 750
rect 615 621 628 667
rect 674 621 687 667
rect 615 558 687 621
rect 615 512 628 558
rect 674 512 687 558
rect 615 449 687 512
rect 615 403 628 449
rect 674 403 687 449
rect 615 339 687 403
rect 615 293 628 339
rect 674 293 687 339
rect 615 280 687 293
rect 872 667 918 680
rect 872 558 918 621
rect 872 449 918 512
rect 872 339 918 403
rect 1095 679 1141 747
rect 1095 349 1141 633
rect 1339 907 1385 920
rect 1339 793 1385 861
rect 1339 679 1385 747
rect 872 79 918 293
rect 1092 337 1272 349
rect 1092 285 1104 337
rect 1260 285 1272 337
rect 1092 273 1272 285
rect 1339 79 1385 633
rect 1508 135 1576 1044
rect 2611 1036 2791 1044
rect 5741 1019 5817 1031
rect 1672 907 1718 920
rect 1672 794 1718 861
rect 1657 748 1672 754
rect 1901 907 1977 920
rect 1901 861 1916 907
rect 1962 861 1977 907
rect 1901 794 1977 861
rect 1718 748 1733 754
rect 1657 742 1733 748
rect 1657 586 1669 742
rect 1721 586 1733 742
rect 1657 574 1733 586
rect 1901 748 1916 794
rect 1962 748 1977 794
rect 2160 907 2206 920
rect 2160 794 2206 861
rect 1901 681 1977 748
rect 1901 635 1916 681
rect 1962 635 1977 681
rect 1672 567 1718 574
rect 1672 453 1718 521
rect 1672 339 1718 407
rect 1672 79 1718 293
rect 1901 567 1977 635
rect 2145 748 2160 754
rect 2389 907 2465 920
rect 2389 861 2404 907
rect 2450 861 2465 907
rect 2389 794 2465 861
rect 2206 748 2221 754
rect 2145 742 2221 748
rect 2145 586 2157 742
rect 2209 586 2221 742
rect 2145 574 2221 586
rect 2389 748 2404 794
rect 2450 748 2465 794
rect 2648 907 2694 920
rect 2648 794 2694 861
rect 2389 681 2465 748
rect 2389 635 2404 681
rect 2450 635 2465 681
rect 1901 521 1916 567
rect 1962 521 1977 567
rect 1901 453 1977 521
rect 1901 407 1916 453
rect 1962 407 1977 453
rect 1901 339 1977 407
rect 1901 293 1916 339
rect 1962 293 1977 339
rect 1901 217 1977 293
rect 2160 567 2206 574
rect 2160 453 2206 521
rect 2160 339 2206 407
rect 2160 280 2206 293
rect 2389 567 2465 635
rect 2634 748 2648 754
rect 2877 918 3921 994
rect 2877 907 2953 918
rect 2877 861 2892 907
rect 2938 861 2953 907
rect 2877 794 2953 861
rect 2694 748 2710 754
rect 2634 742 2710 748
rect 2634 586 2646 742
rect 2698 586 2710 742
rect 2634 574 2710 586
rect 2877 748 2892 794
rect 2938 748 2953 794
rect 2877 681 2953 748
rect 2877 635 2892 681
rect 2938 635 2953 681
rect 2389 521 2404 567
rect 2450 521 2465 567
rect 2389 453 2465 521
rect 2389 407 2404 453
rect 2450 407 2465 453
rect 2389 339 2465 407
rect 2389 293 2404 339
rect 2450 293 2465 339
rect 2389 219 2465 293
rect 2648 567 2694 574
rect 2648 453 2694 521
rect 2648 339 2694 407
rect 2648 280 2694 293
rect 2877 567 2953 635
rect 2877 521 2892 567
rect 2938 521 2953 567
rect 2877 453 2953 521
rect 2877 407 2892 453
rect 2938 407 2953 453
rect 2877 339 2953 407
rect 2877 293 2892 339
rect 2938 293 2953 339
rect 2877 219 2953 293
rect 2389 217 2953 219
rect 1901 159 2953 217
rect 3113 855 3189 868
rect 3113 809 3128 855
rect 3174 809 3189 855
rect 3113 741 3189 809
rect 3113 695 3128 741
rect 3174 695 3189 741
rect 3113 627 3189 695
rect 3113 581 3128 627
rect 3174 581 3189 627
rect 3113 512 3189 581
rect 3113 466 3128 512
rect 3174 466 3189 512
rect 3113 397 3189 466
rect 3113 351 3128 397
rect 3174 351 3189 397
rect 3113 235 3189 351
rect 3357 855 3433 918
rect 3357 809 3372 855
rect 3418 809 3433 855
rect 3357 741 3433 809
rect 3357 695 3372 741
rect 3418 695 3433 741
rect 3357 627 3433 695
rect 3357 581 3372 627
rect 3418 581 3433 627
rect 3357 512 3433 581
rect 3357 466 3372 512
rect 3418 466 3433 512
rect 3357 397 3433 466
rect 3357 351 3372 397
rect 3418 351 3433 397
rect 3357 338 3433 351
rect 3601 855 3677 868
rect 3601 809 3616 855
rect 3662 809 3677 855
rect 3601 741 3677 809
rect 3601 695 3616 741
rect 3662 695 3677 741
rect 3601 627 3677 695
rect 3601 581 3616 627
rect 3662 581 3677 627
rect 3601 512 3677 581
rect 3601 466 3616 512
rect 3662 466 3677 512
rect 3601 397 3677 466
rect 3601 351 3616 397
rect 3662 351 3677 397
rect 3601 235 3677 351
rect 3845 855 3921 918
rect 4233 948 5658 994
rect 4233 918 5285 948
rect 4233 868 4309 918
rect 3845 809 3860 855
rect 3906 809 3921 855
rect 3845 741 3921 809
rect 3845 695 3860 741
rect 3906 695 3921 741
rect 3845 627 3921 695
rect 3845 581 3860 627
rect 3906 581 3921 627
rect 3845 512 3921 581
rect 3845 466 3860 512
rect 3906 466 3921 512
rect 3845 397 3921 466
rect 3845 351 3860 397
rect 3906 351 3921 397
rect 3845 338 3921 351
rect 4089 855 4311 868
rect 4089 809 4104 855
rect 4150 809 4248 855
rect 4294 809 4311 855
rect 4089 750 4311 809
rect 4089 741 4248 750
rect 4089 695 4104 741
rect 4150 704 4248 741
rect 4294 704 4311 750
rect 4150 695 4311 704
rect 4089 645 4311 695
rect 4477 856 4553 868
rect 4477 700 4489 856
rect 4541 700 4553 856
rect 4477 688 4553 700
rect 4721 855 4797 918
rect 4721 809 4736 855
rect 4782 809 4797 855
rect 4721 750 4797 809
rect 4721 704 4736 750
rect 4782 704 4797 750
rect 4089 627 4248 645
rect 4089 581 4104 627
rect 4150 599 4248 627
rect 4294 599 4311 645
rect 4150 581 4311 599
rect 4089 539 4311 581
rect 4089 512 4248 539
rect 4089 466 4104 512
rect 4150 493 4248 512
rect 4294 493 4311 539
rect 4150 466 4311 493
rect 4089 433 4311 466
rect 4089 397 4248 433
rect 4089 351 4104 397
rect 4150 387 4248 397
rect 4294 387 4311 433
rect 4150 351 4311 387
rect 4089 327 4311 351
rect 4089 281 4248 327
rect 4294 281 4311 327
rect 4089 235 4311 281
rect 4492 645 4538 688
rect 4492 539 4538 599
rect 4492 433 4538 493
rect 4492 327 4538 387
rect 4492 268 4538 281
rect 4721 645 4797 704
rect 4965 857 5041 869
rect 4965 701 4977 857
rect 5029 701 5041 857
rect 4965 689 5041 701
rect 5209 855 5285 918
rect 5209 809 5224 855
rect 5270 809 5285 855
rect 5209 750 5285 809
rect 5209 704 5224 750
rect 5270 704 5285 750
rect 4721 599 4736 645
rect 4782 599 4797 645
rect 4721 539 4797 599
rect 4721 493 4736 539
rect 4782 493 4797 539
rect 4721 433 4797 493
rect 4721 387 4736 433
rect 4782 387 4797 433
rect 4721 327 4797 387
rect 4721 281 4736 327
rect 4782 281 4797 327
rect 3113 233 4311 235
rect 4721 233 4797 281
rect 4980 645 5026 689
rect 4980 539 5026 599
rect 4980 433 5026 493
rect 4980 327 5026 387
rect 4980 268 5026 281
rect 5209 645 5285 704
rect 5353 856 5429 868
rect 5353 700 5365 856
rect 5417 700 5429 856
rect 5353 688 5429 700
rect 5612 855 5658 948
rect 5209 599 5224 645
rect 5270 599 5285 645
rect 5368 667 5414 688
rect 5368 608 5414 621
rect 5612 667 5658 809
rect 5741 863 5753 1019
rect 5805 863 5817 1019
rect 5741 858 5756 863
rect 5802 858 5817 863
rect 5741 790 5817 858
rect 5741 751 5756 790
rect 5802 751 5817 790
rect 6000 1019 6190 1031
rect 6000 1018 6017 1019
rect 6173 1018 6190 1019
rect 6000 904 6017 972
rect 6173 904 6190 972
rect 6046 858 6144 863
rect 6000 790 6190 858
rect 5756 731 5802 744
rect 6046 744 6144 790
rect 6000 731 6190 744
rect 6373 1019 6449 1031
rect 6373 863 6385 1019
rect 6437 863 6449 1019
rect 6373 858 6388 863
rect 6434 858 6449 863
rect 6373 790 6449 858
rect 6373 744 6388 790
rect 6434 744 6449 790
rect 5612 608 5658 621
rect 5209 539 5285 599
rect 5209 493 5224 539
rect 5270 493 5285 539
rect 6373 505 6449 744
rect 5209 433 5285 493
rect 5451 494 6449 505
rect 5451 448 5462 494
rect 5602 448 6449 494
rect 5451 437 6449 448
rect 6710 1008 6778 1019
rect 5209 387 5224 433
rect 5270 387 5285 433
rect 5209 327 5285 387
rect 5209 281 5224 327
rect 5270 281 5285 327
rect 5209 233 5285 281
rect 3113 159 4165 233
rect 6450 79 6630 87
rect 6710 79 6721 1008
rect 151 75 6721 79
rect 151 68 6462 75
rect 151 22 269 68
rect 6618 23 6721 75
rect 6613 22 6721 23
rect 6767 22 6778 1008
rect 8 11 6778 22
<< via1 >>
rect 1835 1924 1838 1965
rect 1838 1924 1884 1965
rect 1884 1924 1887 1965
rect 1835 1856 1887 1924
rect 1835 1810 1838 1856
rect 1838 1810 1884 1856
rect 1884 1810 1887 1856
rect 1835 1809 1887 1810
rect 3239 2097 3291 2210
rect 3239 2054 3240 2097
rect 3240 2054 3286 2097
rect 3286 2054 3291 2097
rect 3018 1856 3070 1898
rect 3018 1810 3022 1856
rect 3022 1810 3068 1856
rect 3068 1810 3070 1856
rect 3018 1742 3070 1810
rect 3613 2202 3769 2254
rect 4107 2101 4108 2106
rect 4108 2101 4154 2106
rect 4154 2101 4159 2106
rect 4107 2028 4159 2101
rect 4107 1982 4108 2028
rect 4108 1982 4154 2028
rect 4154 1982 4159 2028
rect 4107 1950 4159 1982
rect 4591 2101 4596 2106
rect 4596 2101 4642 2106
rect 4642 2101 4643 2106
rect 4591 2028 4643 2101
rect 4591 1982 4596 2028
rect 4596 1982 4642 2028
rect 4642 1982 4643 2028
rect 4591 1950 4643 1982
rect 4349 1863 4352 1898
rect 4352 1863 4398 1898
rect 4398 1863 4401 1898
rect 4349 1789 4401 1863
rect 4349 1743 4352 1789
rect 4352 1743 4398 1789
rect 4398 1743 4401 1789
rect 4349 1742 4401 1743
rect 5215 2097 5267 2106
rect 5215 1950 5228 2097
rect 5228 1950 5267 2097
rect 5753 1759 5756 1804
rect 5756 1759 5802 1804
rect 5802 1759 5805 1804
rect 5753 1696 5805 1759
rect 5753 1650 5756 1696
rect 5756 1650 5802 1696
rect 5802 1650 5805 1696
rect 5753 1648 5805 1650
rect 6017 1759 6046 1805
rect 6046 1759 6144 1805
rect 6144 1759 6173 1805
rect 6017 1696 6173 1759
rect 6017 1650 6046 1696
rect 6046 1650 6144 1696
rect 6144 1650 6173 1696
rect 6017 1649 6173 1650
rect 6385 1759 6388 1805
rect 6388 1759 6434 1805
rect 6434 1759 6437 1805
rect 6385 1696 6437 1759
rect 6385 1650 6388 1696
rect 6388 1650 6434 1696
rect 6434 1650 6437 1696
rect 6385 1649 6437 1650
rect 2623 1579 2749 1624
rect 2749 1579 2779 1624
rect 2623 1572 2779 1579
rect 3888 1580 4044 1632
rect 6566 1625 6618 1781
rect 1154 1454 1310 1506
rect 1652 1454 1808 1506
rect 2966 1311 3122 1363
rect 4361 1312 4517 1364
rect 4873 1312 5029 1364
rect 6017 1312 6173 1364
rect 1504 1180 1660 1232
rect 630 930 750 982
rect 750 930 786 982
rect 2623 1055 2723 1100
rect 2723 1055 2779 1100
rect 2623 1048 2779 1055
rect 4028 1101 4184 1108
rect 4028 1056 4075 1101
rect 4075 1056 4184 1101
rect 1104 285 1260 337
rect 1669 681 1721 742
rect 1669 635 1672 681
rect 1672 635 1718 681
rect 1718 635 1721 681
rect 1669 586 1721 635
rect 2157 681 2209 742
rect 2157 635 2160 681
rect 2160 635 2206 681
rect 2206 635 2209 681
rect 2157 586 2209 635
rect 2646 681 2698 742
rect 2646 635 2648 681
rect 2648 635 2694 681
rect 2694 635 2698 681
rect 2646 586 2698 635
rect 4489 855 4541 856
rect 4489 809 4492 855
rect 4492 809 4538 855
rect 4538 809 4541 855
rect 4489 750 4541 809
rect 4489 704 4492 750
rect 4492 704 4538 750
rect 4538 704 4541 750
rect 4489 700 4541 704
rect 4977 855 5029 857
rect 4977 809 4980 855
rect 4980 809 5026 855
rect 5026 809 5029 855
rect 4977 750 5029 809
rect 4977 704 4980 750
rect 4980 704 5026 750
rect 5026 704 5029 750
rect 4977 701 5029 704
rect 5365 855 5417 856
rect 5365 809 5368 855
rect 5368 809 5414 855
rect 5414 809 5417 855
rect 5365 700 5417 809
rect 5753 1018 5805 1019
rect 5753 972 5756 1018
rect 5756 972 5802 1018
rect 5802 972 5805 1018
rect 5753 904 5805 972
rect 5753 863 5756 904
rect 5756 863 5802 904
rect 5802 863 5805 904
rect 6017 1018 6173 1019
rect 6017 972 6046 1018
rect 6046 972 6144 1018
rect 6144 972 6173 1018
rect 6017 904 6173 972
rect 6017 863 6046 904
rect 6046 863 6144 904
rect 6144 863 6173 904
rect 6385 1018 6437 1019
rect 6385 972 6388 1018
rect 6388 972 6434 1018
rect 6434 972 6437 1018
rect 6385 904 6437 972
rect 6385 863 6388 904
rect 6388 863 6434 904
rect 6434 863 6437 904
rect 6462 68 6618 75
rect 6462 23 6613 68
rect 6613 23 6618 68
<< metal2 >>
rect 3227 2254 3781 2266
rect 3227 2210 3613 2254
rect 3227 2054 3239 2210
rect 3291 2202 3613 2210
rect 3769 2202 3781 2254
rect 3291 2190 3781 2202
rect 3291 2054 3303 2190
rect 3227 2042 3303 2054
rect 4095 2106 5279 2118
rect 1823 1965 1968 1977
rect 1823 1809 1835 1965
rect 1887 1809 1968 1965
rect 4095 1950 4107 2106
rect 4159 2042 4591 2106
rect 4159 1950 4171 2042
rect 4095 1938 4171 1950
rect 1823 1797 1968 1809
rect 1142 1506 1820 1518
rect 1142 1454 1154 1506
rect 1310 1454 1652 1506
rect 1808 1454 1820 1506
rect 1142 1442 1820 1454
rect 1150 1232 1672 1244
rect 1150 1180 1504 1232
rect 1660 1180 1672 1232
rect 1150 1168 1672 1180
rect 1150 994 1330 1168
rect 1896 1029 1968 1797
rect 3006 1898 3082 1910
rect 3006 1742 3018 1898
rect 3070 1742 3082 1898
rect 2611 1624 2791 1636
rect 2611 1572 2623 1624
rect 2779 1572 2791 1624
rect 2611 1100 2791 1572
rect 3006 1396 3082 1742
rect 4326 1898 4435 1967
rect 4579 1950 4591 2042
rect 4643 2042 5215 2106
rect 4643 1950 4655 2042
rect 4579 1938 4655 1950
rect 5203 1950 5215 2042
rect 5267 1950 5279 2106
rect 5203 1938 5279 1950
rect 4326 1742 4349 1898
rect 4401 1742 4435 1898
rect 3876 1632 4056 1644
rect 3876 1580 3888 1632
rect 4044 1580 4056 1632
rect 3876 1568 4056 1580
rect 2954 1363 3134 1396
rect 2954 1311 2966 1363
rect 3122 1311 3134 1363
rect 2954 1280 3134 1311
rect 2611 1048 2623 1100
rect 2779 1048 2791 1100
rect 2611 1036 2791 1048
rect 3915 1120 4019 1568
rect 4326 1376 4435 1742
rect 4326 1364 4553 1376
rect 4326 1312 4361 1364
rect 4517 1312 4553 1364
rect 4326 1300 4553 1312
rect 4861 1364 5041 1376
rect 4861 1312 4873 1364
rect 5029 1312 5041 1364
rect 4861 1300 5041 1312
rect 3915 1108 4196 1120
rect 3915 1056 4028 1108
rect 4184 1056 4196 1108
rect 3915 1044 4196 1056
rect 618 982 798 994
rect 618 930 630 982
rect 786 930 798 982
rect 618 918 798 930
rect 826 918 1330 994
rect 1480 953 1968 1029
rect 1480 485 1556 953
rect 4477 856 4553 1300
rect 1657 742 2710 754
rect 1657 586 1669 742
rect 1721 586 2157 742
rect 2209 586 2646 742
rect 2698 586 2710 742
rect 4477 700 4489 856
rect 4541 700 4553 856
rect 4477 688 4553 700
rect 4965 857 5041 1300
rect 5364 1052 5468 2252
rect 5555 926 5631 2481
rect 4965 701 4977 857
rect 5029 701 5041 857
rect 4965 689 5041 701
rect 5353 861 5631 926
rect 5741 1804 5817 1816
rect 5741 1648 5753 1804
rect 5805 1648 5817 1804
rect 5741 1019 5817 1648
rect 5741 863 5753 1019
rect 5805 863 5817 1019
rect 5353 856 5429 861
rect 5353 700 5365 856
rect 5417 700 5429 856
rect 5353 688 5429 700
rect 1657 574 2710 586
rect 5741 485 5817 863
rect 6005 1805 6185 1817
rect 6005 1649 6017 1805
rect 6173 1649 6185 1805
rect 6005 1364 6185 1649
rect 6005 1312 6017 1364
rect 6173 1312 6185 1364
rect 6005 1019 6185 1312
rect 6005 863 6017 1019
rect 6173 863 6185 1019
rect 6005 851 6185 863
rect 6373 1805 6449 1817
rect 6373 1649 6385 1805
rect 6437 1649 6449 1805
rect 6373 1019 6449 1649
rect 6373 863 6385 1019
rect 6437 863 6449 1019
rect 1480 409 5817 485
rect 6373 349 6449 863
rect 1092 337 6449 349
rect 1092 285 1104 337
rect 1260 285 6449 337
rect 1092 273 6449 285
rect 6554 1781 6630 1793
rect 6554 1625 6566 1781
rect 6618 1625 6630 1781
rect 6554 87 6630 1625
rect 6450 75 6630 87
rect 6450 23 6462 75
rect 6618 23 6630 75
rect 6450 11 6630 23
use M1_NWELL_CDNS_40661956134418  M1_NWELL_CDNS_40661956134418_0
timestamp 1698431365
transform 1 0 6744 0 1 1977
box 0 0 1 1
use M1_NWELL_CDNS_40661956134418  M1_NWELL_CDNS_40661956134418_1
timestamp 1698431365
transform 1 0 128 0 1 1977
box 0 0 1 1
use M1_NWELL_CDNS_40661956134421  M1_NWELL_CDNS_40661956134421_0
timestamp 1698431365
transform 1 0 3441 0 1 2447
box 0 0 1 1
use M1_NWELL_CDNS_40661956134423  M1_NWELL_CDNS_40661956134423_0
timestamp 1698431365
transform 1 0 -650 0 1 2031
box 0 0 1 1
use M1_POLY2_CDNS_40661956134128  M1_POLY2_CDNS_40661956134128_0
timestamp 1698431365
transform 1 0 2549 0 1 1078
box 0 0 1 1
use M1_POLY2_CDNS_40661956134128  M1_POLY2_CDNS_40661956134128_1
timestamp 1698431365
transform 1 0 2061 0 1 1078
box 0 0 1 1
use M1_POLY2_CDNS_40661956134128  M1_POLY2_CDNS_40661956134128_2
timestamp 1698431365
transform 1 0 5532 0 1 471
box 0 0 1 1
use M1_POLY2_CDNS_40661956134128  M1_POLY2_CDNS_40661956134128_3
timestamp 1698431365
transform 1 0 1240 0 1 1078
box 0 0 1 1
use M1_POLY2_CDNS_40661956134128  M1_POLY2_CDNS_40661956134128_4
timestamp 1698431365
transform 1 0 2305 0 1 1078
box 0 0 1 1
use M1_POLY2_CDNS_40661956134128  M1_POLY2_CDNS_40661956134128_5
timestamp 1698431365
transform 1 0 2793 0 1 1078
box 0 0 1 1
use M1_POLY2_CDNS_40661956134128  M1_POLY2_CDNS_40661956134128_6
timestamp 1698431365
transform 1 0 1817 0 1 1078
box 0 0 1 1
use M1_POLY2_CDNS_40661956134326  M1_POLY2_CDNS_40661956134326_0
timestamp 1698431365
transform 0 1 6289 1 0 1486
box 0 0 1 1
use M1_POLY2_CDNS_40661956134326  M1_POLY2_CDNS_40661956134326_1
timestamp 1698431365
transform 0 1 5901 1 0 1486
box 0 0 1 1
use M1_POLY2_CDNS_40661956134326  M1_POLY2_CDNS_40661956134326_2
timestamp 1698431365
transform 1 0 529 0 -1 957
box 0 0 1 1
use M1_POLY2_CDNS_40661956134326  M1_POLY2_CDNS_40661956134326_3
timestamp 1698431365
transform 1 0 773 0 -1 957
box 0 0 1 1
use M1_POLY2_CDNS_40661956134326  M1_POLY2_CDNS_40661956134326_4
timestamp 1698431365
transform 0 1 5901 -1 0 1190
box 0 0 1 1
use M1_POLY2_CDNS_40661956134326  M1_POLY2_CDNS_40661956134326_5
timestamp 1698431365
transform 0 1 6289 -1 0 1190
box 0 0 1 1
use M1_POLY2_CDNS_40661956134326  M1_POLY2_CDNS_40661956134326_6
timestamp 1698431365
transform 0 -1 3629 1 0 1602
box 0 0 1 1
use M1_POLY2_CDNS_40661956134326  M1_POLY2_CDNS_40661956134326_7
timestamp 1698431365
transform 0 -1 5129 1 0 1602
box 0 0 1 1
use M1_POLY2_CDNS_40661956134326  M1_POLY2_CDNS_40661956134326_8
timestamp 1698431365
transform 0 -1 3385 1 0 1602
box 0 0 1 1
use M1_POLY2_CDNS_40661956134326  M1_POLY2_CDNS_40661956134326_9
timestamp 1698431365
transform 0 -1 4253 1 0 1602
box 0 0 1 1
use M1_POLY2_CDNS_40661956134326  M1_POLY2_CDNS_40661956134326_10
timestamp 1698431365
transform 0 -1 4881 1 0 1078
box 0 0 1 1
use M1_POLY2_CDNS_40661956134326  M1_POLY2_CDNS_40661956134326_11
timestamp 1698431365
transform 0 -1 3761 1 0 1078
box 0 0 1 1
use M1_POLY2_CDNS_40661956134326  M1_POLY2_CDNS_40661956134326_12
timestamp 1698431365
transform 0 -1 3273 1 0 1078
box 0 0 1 1
use M1_POLY2_CDNS_40661956134326  M1_POLY2_CDNS_40661956134326_13
timestamp 1698431365
transform 0 -1 3517 1 0 1078
box 0 0 1 1
use M1_POLY2_CDNS_40661956134326  M1_POLY2_CDNS_40661956134326_14
timestamp 1698431365
transform 0 -1 5125 1 0 1078
box 0 0 1 1
use M1_POLY2_CDNS_40661956134326  M1_POLY2_CDNS_40661956134326_15
timestamp 1698431365
transform 0 -1 4637 1 0 1078
box 0 0 1 1
use M1_POLY2_CDNS_40661956134326  M1_POLY2_CDNS_40661956134326_16
timestamp 1698431365
transform 0 -1 4393 1 0 1078
box 0 0 1 1
use M1_POLY2_CDNS_40661956134326  M1_POLY2_CDNS_40661956134326_17
timestamp 1698431365
transform 0 -1 4885 1 0 1602
box 0 0 1 1
use M1_POLY2_CDNS_40661956134326  M1_POLY2_CDNS_40661956134326_18
timestamp 1698431365
transform 0 -1 4497 1 0 1602
box 0 0 1 1
use M1_POLY2_CDNS_40661956134326  M1_POLY2_CDNS_40661956134326_19
timestamp 1698431365
transform 0 -1 1983 1 0 1602
box 0 0 1 1
use M1_POLY2_CDNS_40661956134326  M1_POLY2_CDNS_40661956134326_20
timestamp 1698431365
transform 0 -1 1739 1 0 1602
box 0 0 1 1
use M1_POLY2_CDNS_40661956134326  M1_POLY2_CDNS_40661956134326_21
timestamp 1698431365
transform 0 -1 2923 1 0 1602
box 0 0 1 1
use M1_POLY2_CDNS_40661956134326  M1_POLY2_CDNS_40661956134326_22
timestamp 1698431365
transform 0 -1 2679 1 0 1602
box 0 0 1 1
use M1_POLY2_CDNS_40661956134326  M1_POLY2_CDNS_40661956134326_23
timestamp 1698431365
transform 0 -1 4005 1 0 1078
box 0 0 1 1
use M1_POLY2_CDNS_40661956134326  M1_POLY2_CDNS_40661956134326_24
timestamp 1698431365
transform 0 -1 2435 1 0 1602
box 0 0 1 1
use M1_PSUB_CDNS_40661956134330  M1_PSUB_CDNS_40661956134330_0
timestamp 1698431365
transform 1 0 6744 0 -1 515
box 0 0 1 1
use M1_PSUB_CDNS_40661956134330  M1_PSUB_CDNS_40661956134330_1
timestamp 1698431365
transform 1 0 128 0 -1 515
box 0 0 1 1
use M1_PSUB_CDNS_40661956134420  M1_PSUB_CDNS_40661956134420_0
timestamp 1698431365
transform 1 0 3441 0 -1 45
box 0 0 1 1
use M1_PSUB_CDNS_40661956134422  M1_PSUB_CDNS_40661956134422_0
timestamp 1698431365
transform 1 0 -650 0 1 569
box 0 0 1 1
use M2_M1_CDNS_40661956134235  M2_M1_CDNS_40661956134235_0
timestamp 1698431365
transform 1 0 6095 0 1 1727
box 0 0 1 1
use M2_M1_CDNS_40661956134235  M2_M1_CDNS_40661956134235_1
timestamp 1698431365
transform 1 0 6095 0 1 941
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_0
timestamp 1698431365
transform 1 0 6540 0 1 49
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_1
timestamp 1698431365
transform 1 0 3966 0 1 1606
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_2
timestamp 1698431365
transform 1 0 1730 0 1 1480
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_3
timestamp 1698431365
transform 1 0 4439 0 1 1338
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_4
timestamp 1698431365
transform 1 0 6095 0 1 1338
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_5
timestamp 1698431365
transform 1 0 3044 0 1 1337
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_6
timestamp 1698431365
transform 1 0 2701 0 1 1598
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_7
timestamp 1698431365
transform 1 0 2701 0 1 1074
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_8
timestamp 1698431365
transform 1 0 4951 0 1 1338
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_9
timestamp 1698431365
transform 1 0 3691 0 1 2228
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_10
timestamp 1698431365
transform 1 0 1582 0 1 1206
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_11
timestamp 1698431365
transform 1 0 1232 0 1 1480
box 0 0 1 1
use M2_M1_CDNS_40661956134237  M2_M1_CDNS_40661956134237_12
timestamp 1698431365
transform 1 0 4106 0 1 1082
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_0
timestamp 1698431365
transform 0 -1 708 1 0 956
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_1
timestamp 1698431365
transform 0 -1 1182 1 0 311
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_2
timestamp 1698431365
transform 1 0 4375 0 1 1820
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_3
timestamp 1698431365
transform 1 0 4133 0 1 2028
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_4
timestamp 1698431365
transform 1 0 3265 0 1 2132
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_5
timestamp 1698431365
transform 1 0 2672 0 1 664
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_6
timestamp 1698431365
transform 1 0 5003 0 1 779
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_7
timestamp 1698431365
transform 1 0 4515 0 1 778
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_8
timestamp 1698431365
transform 1 0 5391 0 1 778
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_9
timestamp 1698431365
transform 1 0 2183 0 1 664
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_10
timestamp 1698431365
transform 1 0 4617 0 1 2028
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_11
timestamp 1698431365
transform 1 0 1861 0 1 1887
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_12
timestamp 1698431365
transform 1 0 5779 0 1 1726
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_13
timestamp 1698431365
transform 1 0 6411 0 1 941
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_14
timestamp 1698431365
transform 1 0 5779 0 1 941
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_15
timestamp 1698431365
transform 1 0 6411 0 1 1727
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_16
timestamp 1698431365
transform 1 0 5241 0 1 2028
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_17
timestamp 1698431365
transform 1 0 1695 0 1 664
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_18
timestamp 1698431365
transform 1 0 3044 0 1 1820
box 0 0 1 1
use M2_M1_CDNS_40661956134270  M2_M1_CDNS_40661956134270_19
timestamp 1698431365
transform 1 0 6592 0 1 1703
box 0 0 1 1
use nmos_6p0_CDNS_4066195613430  nmos_6p0_CDNS_4066195613430_0
timestamp 1698431365
transform 1 0 6219 0 1 731
box 0 0 1 1
use nmos_6p0_CDNS_4066195613435  nmos_6p0_CDNS_4066195613435_0
timestamp 1698431365
transform 1 0 459 0 1 280
box 0 0 1 1
use nmos_6p0_CDNS_4066195613436  nmos_6p0_CDNS_4066195613436_0
timestamp 1698431365
transform -1 0 1310 0 -1 920
box 0 0 1 1
use nmos_6p0_CDNS_4066195613436  nmos_6p0_CDNS_4066195613436_1
timestamp 1698431365
transform 1 0 5831 0 1 731
box 0 0 1 1
use nmos_6p0_CDNS_4066195613437  nmos_6p0_CDNS_4066195613437_0
timestamp 1698431365
transform 1 0 1747 0 1 280
box 0 0 1 1
use nmos_6p0_CDNS_4066195613440  nmos_6p0_CDNS_4066195613440_0
timestamp 1698431365
transform 1 0 5443 0 1 608
box 0 0 1 1
use nmos_6p0_CDNS_4066195613441  nmos_6p0_CDNS_4066195613441_0
timestamp 1698431365
transform 1 0 3203 0 1 338
box 0 0 1 1
use nmos_6p0_CDNS_4066195613442  nmos_6p0_CDNS_4066195613442_0
timestamp 1698431365
transform 1 0 4323 0 1 268
box 0 0 1 1
use pmos_6p0_CDNS_4066195613434  pmos_6p0_CDNS_4066195613434_0
timestamp 1698431365
transform -1 0 2053 0 1 1797
box 0 0 1 1
use pmos_6p0_CDNS_4066195613438  pmos_6p0_CDNS_4066195613438_0
timestamp 1698431365
transform 1 0 4183 0 1 1730
box 0 0 1 1
use pmos_6p0_CDNS_4066195613439  pmos_6p0_CDNS_4066195613439_0
timestamp 1698431365
transform 1 0 6219 0 -1 2037
box 0 0 1 1
use pmos_6p0_CDNS_4066195613439  pmos_6p0_CDNS_4066195613439_1
timestamp 1698431365
transform -1 0 5971 0 -1 2037
box 0 0 1 1
use pmos_6p0_CDNS_4066195613443  pmos_6p0_CDNS_4066195613443_0
timestamp 1698431365
transform -1 0 2993 0 -1 2197
box 0 0 1 1
use pmos_6p0_CDNS_4066195613444  pmos_6p0_CDNS_4066195613444_0
timestamp 1698431365
transform 1 0 4815 0 1 1730
box 0 0 1 1
use pmos_6p0_CDNS_4066195613444  pmos_6p0_CDNS_4066195613444_1
timestamp 1698431365
transform 1 0 3315 0 1 1730
box 0 0 1 1
use pmos_6p0_CDNS_4066195613445  pmos_6p0_CDNS_4066195613445_0
timestamp 1698431365
transform -1 0 843 0 1 1335
box 0 0 1 1
<< labels >>
rlabel metal2 s 2695 1339 2695 1339 4 IE
port 1 nsew
rlabel metal2 s 855 960 855 960 4 CS
port 2 nsew
rlabel metal1 s 884 2452 884 2452 4 DVDD
port 3 nsew
rlabel metal1 s 4228 1072 4228 1072 4 A
port 4 nsew
rlabel metal1 s 320 39 320 39 4 DVSS
port 5 nsew
rlabel metal1 s 6269 1344 6269 1344 4 Z
port 6 nsew
<< properties >>
string GDS_END 1119770
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 1104652
string path 80.675 55.700 93.150 55.700 
<< end >>
