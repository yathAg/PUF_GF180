magic
tech gf180mcuB
magscale 1 10
timestamp 1698431365
<< obsm1 >>
rect 13108 13108 71000 71000
<< obsm2 >>
rect 13606 13594 70901 70890
<< metal3 >>
rect 14000 70800 17000 71000
rect 17200 70800 20200 71000
rect 20400 70800 23400 71000
rect 23600 70800 25000 71000
rect 25200 70800 26600 71000
rect 26800 70800 29800 71000
rect 30000 70800 33000 71000
rect 33200 70800 36200 71000
rect 36400 70800 39400 71000
rect 39600 70800 41000 71000
rect 41200 70800 42600 71000
rect 42800 70800 45800 71000
rect 46000 70800 49000 71000
rect 49200 70800 50600 71000
rect 50800 70800 52200 71000
rect 52400 70800 53800 71000
rect 54000 70800 55400 71000
rect 55600 70800 57000 71000
rect 57200 70800 58600 71000
rect 58800 70800 60200 71000
rect 60400 70800 61800 71000
rect 62000 70800 63400 71000
rect 63600 70800 65000 71000
rect 65200 70800 66600 71000
rect 66800 70800 68200 71000
rect 68400 70800 69678 71000
rect 70800 68400 71000 69678
rect 70800 66800 71000 68200
rect 70800 65200 71000 66600
rect 70800 63600 71000 65000
rect 70800 62000 71000 63400
rect 70800 60400 71000 61800
rect 70800 58800 71000 60200
rect 70800 57200 71000 58600
rect 70800 55600 71000 57000
rect 70800 54000 71000 55400
rect 70800 52400 71000 53800
rect 70800 50800 71000 52200
rect 70800 49200 71000 50600
rect 70800 46000 71000 49000
rect 70800 42800 71000 45800
rect 70800 41200 71000 42600
rect 70800 39600 71000 41000
rect 70800 36400 71000 39400
rect 70800 33200 71000 36200
rect 70800 30000 71000 33000
rect 70800 26800 71000 29800
rect 70800 25200 71000 26600
rect 70800 23600 71000 25000
rect 70800 20400 71000 23400
rect 70800 17200 71000 20200
rect 70800 14000 71000 17000
<< obsm3 >>
rect 17060 70740 17140 70890
rect 20260 70740 20340 70890
rect 23460 70740 23540 70890
rect 25060 70740 25140 70890
rect 26660 70740 26740 70890
rect 29860 70740 29940 70890
rect 33060 70740 33140 70890
rect 36260 70740 36340 70890
rect 39460 70740 39540 70890
rect 41060 70740 41140 70890
rect 42660 70740 42740 70890
rect 45860 70740 45940 70890
rect 49060 70740 49140 70890
rect 50660 70740 50740 70890
rect 52260 70740 52340 70890
rect 53860 70740 53940 70890
rect 55460 70740 55540 70890
rect 57060 70740 57140 70890
rect 58660 70740 58740 70890
rect 60260 70740 60340 70890
rect 61860 70740 61940 70890
rect 63460 70740 63540 70890
rect 65060 70740 65140 70890
rect 66660 70740 66740 70890
rect 68260 70740 68340 70890
rect 69738 70740 70800 70890
rect 14000 69738 70800 70740
rect 14000 68340 70740 69738
rect 14000 68260 70800 68340
rect 14000 66740 70740 68260
rect 14000 66660 70800 66740
rect 14000 65140 70740 66660
rect 14000 65060 70800 65140
rect 14000 63540 70740 65060
rect 14000 63460 70800 63540
rect 14000 61940 70740 63460
rect 14000 61860 70800 61940
rect 14000 60340 70740 61860
rect 14000 60260 70800 60340
rect 14000 58740 70740 60260
rect 14000 58660 70800 58740
rect 14000 57140 70740 58660
rect 14000 57060 70800 57140
rect 14000 55540 70740 57060
rect 14000 55460 70800 55540
rect 14000 53940 70740 55460
rect 14000 53860 70800 53940
rect 14000 52340 70740 53860
rect 14000 52260 70800 52340
rect 14000 50740 70740 52260
rect 14000 50660 70800 50740
rect 14000 49140 70740 50660
rect 14000 49060 70800 49140
rect 14000 45940 70740 49060
rect 14000 45860 70800 45940
rect 14000 42740 70740 45860
rect 14000 42660 70800 42740
rect 14000 41140 70740 42660
rect 14000 41060 70800 41140
rect 14000 39540 70740 41060
rect 14000 39460 70800 39540
rect 14000 36340 70740 39460
rect 14000 36260 70800 36340
rect 14000 33140 70740 36260
rect 14000 33060 70800 33140
rect 14000 29940 70740 33060
rect 14000 29860 70800 29940
rect 14000 26740 70740 29860
rect 14000 26660 70800 26740
rect 14000 25140 70740 26660
rect 14000 25060 70800 25140
rect 14000 23540 70740 25060
rect 14000 23460 70800 23540
rect 14000 20340 70740 23460
rect 14000 20260 70800 20340
rect 14000 17140 70740 20260
rect 14000 17060 70800 17140
rect 14000 14000 70740 17060
<< metal4 >>
rect 14000 70800 17000 71000
rect 17200 70800 20200 71000
rect 20400 70800 23400 71000
rect 23600 70800 25000 71000
rect 25200 70800 26600 71000
rect 26800 70800 29800 71000
rect 30000 70800 33000 71000
rect 33200 70800 36200 71000
rect 36400 70800 39400 71000
rect 39600 70800 41000 71000
rect 41200 70800 42600 71000
rect 42800 70800 45800 71000
rect 46000 70800 49000 71000
rect 49200 70800 50600 71000
rect 50800 70800 52200 71000
rect 52400 70800 53800 71000
rect 54000 70800 55400 71000
rect 55600 70800 57000 71000
rect 57200 70800 58600 71000
rect 58800 70800 60200 71000
rect 60400 70800 61800 71000
rect 62000 70800 63400 71000
rect 63600 70800 65000 71000
rect 65200 70800 66600 71000
rect 66800 70800 68200 71000
rect 68400 70800 69678 71000
rect 70800 68400 71000 69678
rect 70800 66800 71000 68200
rect 70800 65200 71000 66600
rect 70800 63600 71000 65000
rect 70800 62000 71000 63400
rect 70800 60400 71000 61800
rect 70800 58800 71000 60200
rect 70800 57200 71000 58600
rect 70800 55600 71000 57000
rect 70800 54000 71000 55400
rect 70800 52400 71000 53800
rect 70800 50800 71000 52200
rect 70800 49200 71000 50600
rect 70800 46000 71000 49000
rect 70800 42800 71000 45800
rect 70800 41200 71000 42600
rect 70800 39600 71000 41000
rect 70800 36400 71000 39400
rect 70800 33200 71000 36200
rect 70800 30000 71000 33000
rect 70800 26800 71000 29800
rect 70800 25200 71000 26600
rect 70800 23600 71000 25000
rect 70800 20400 71000 23400
rect 70800 17200 71000 20200
rect 70800 14000 71000 17000
<< obsm4 >>
rect 69778 70700 70800 70800
rect 14000 69778 70800 70700
rect 14000 14000 70700 69778
<< labels >>
rlabel metal3 s 66800 70800 68200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 66800 71000 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 58800 70800 60200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 58800 71000 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 55600 70800 57000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 55600 71000 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 54000 70800 55400 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 54000 71000 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 52400 70800 53800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 52400 71000 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 42800 70800 45800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 42800 71000 45800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 41200 70800 42600 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 41200 71000 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 36400 70800 39400 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 36400 71000 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 33200 70800 36200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 33200 71000 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 30000 70800 33000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 30000 71000 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 26800 70800 29800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 26800 71000 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 23600 70800 25000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 66800 70800 68200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 66800 71000 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 58800 70800 60200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 58800 71000 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 55600 70800 57000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 55600 71000 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 54000 70800 55400 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 54000 71000 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 52400 70800 53800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 52400 71000 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 42800 70800 45800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 42800 71000 45800 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 41200 70800 42600 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 41200 71000 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 36400 70800 39400 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 36400 71000 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 33200 70800 36200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 33200 71000 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 30000 70800 33000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 30000 71000 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 26800 70800 29800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 26800 71000 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 23600 70800 25000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 23600 71000 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 23600 71000 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 68400 70800 69678 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 68400 71000 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 65200 70800 66600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 65200 71000 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 60400 70800 61800 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 60400 71000 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 57200 70800 58600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 57200 71000 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 46000 70800 49000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 46000 71000 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 39600 70800 41000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 39600 71000 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 25200 70800 26600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 25200 71000 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 20400 70800 23400 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 20400 71000 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 17200 70800 20200 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 17200 71000 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 14000 70800 17000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 68400 70800 69678 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 68400 71000 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 65200 70800 66600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 65200 71000 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 60400 70800 61800 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 60400 71000 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 57200 70800 58600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 57200 71000 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 46000 70800 49000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 46000 71000 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 39600 70800 41000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 39600 71000 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 25200 70800 26600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 25200 71000 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 20400 70800 23400 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 20400 71000 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 17200 70800 20200 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 17200 71000 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 14000 70800 17000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 14000 71000 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 14000 71000 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 62000 70800 63400 71000 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 70800 62000 71000 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 50800 70800 52200 71000 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 62000 70800 63400 71000 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 70800 62000 71000 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 50800 70800 52200 71000 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 70800 50800 71000 52200 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 70800 50800 71000 52200 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 63600 70800 65000 71000 6 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 70800 63600 71000 65000 6 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 49200 70800 50600 71000 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 63600 70800 65000 71000 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 70800 63600 71000 65000 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 49200 70800 50600 71000 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 70800 49200 71000 50600 6 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 70800 49200 71000 50600 6 VSS
port 4 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 71000 71000
string LEFclass ENDCAP BOTTOMLEFT
string LEFsite GF_COR_Site
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 12063666
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 12059128
<< end >>
