magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< obsm1 >>
rect -32 13108 1032 69957
<< obsm2 >>
rect 0 13470 1000 69660
<< metal3 >>
rect 0 68400 200 69678
rect 800 68400 1000 69678
rect 0 66800 200 68200
rect 800 66800 1000 68200
rect 0 65200 200 66600
rect 800 65200 1000 66600
rect 0 63600 200 65000
rect 800 63600 1000 65000
rect 0 62000 200 63400
rect 800 62000 1000 63400
rect 0 60400 200 61800
rect 800 60400 1000 61800
rect 0 58800 200 60200
rect 800 58800 1000 60200
rect 0 57200 200 58600
rect 800 57200 1000 58600
rect 0 55600 200 57000
rect 800 55600 1000 57000
rect 0 54000 200 55400
rect 800 54000 1000 55400
rect 0 52400 200 53800
rect 800 52400 1000 53800
rect 0 50800 200 52200
rect 800 50800 1000 52200
rect 0 49200 200 50600
rect 800 49200 1000 50600
rect 0 46000 200 49000
rect 800 46000 1000 49000
rect 0 42800 200 45800
rect 800 42800 1000 45800
rect 0 41200 200 42600
rect 800 41200 1000 42600
rect 0 39600 200 41000
rect 800 39600 1000 41000
rect 0 36400 200 39400
rect 800 36400 1000 39400
rect 0 33200 200 36200
rect 800 33200 1000 36200
rect 0 30000 200 33000
rect 800 30000 1000 33000
rect 0 26800 200 29800
rect 800 26800 1000 29800
rect 0 25200 200 26600
rect 800 25200 1000 26600
rect 0 23600 200 25000
rect 800 23600 1000 25000
rect 0 20400 200 23400
rect 800 20400 1000 23400
rect 0 17200 200 20200
rect 800 17200 1000 20200
rect 0 14000 200 17000
rect 800 14000 1000 17000
<< obsm3 >>
rect 260 68340 740 69678
rect 200 68260 800 68340
rect 260 66740 740 68260
rect 200 66660 800 66740
rect 260 65140 740 66660
rect 200 65060 800 65140
rect 260 63540 740 65060
rect 200 63460 800 63540
rect 260 61940 740 63460
rect 200 61860 800 61940
rect 260 60340 740 61860
rect 200 60260 800 60340
rect 260 58740 740 60260
rect 200 58660 800 58740
rect 260 57140 740 58660
rect 200 57060 800 57140
rect 260 55540 740 57060
rect 200 55460 800 55540
rect 260 53940 740 55460
rect 200 53860 800 53940
rect 260 52340 740 53860
rect 200 52260 800 52340
rect 260 50740 740 52260
rect 200 50660 800 50740
rect 260 49140 740 50660
rect 200 49060 800 49140
rect 260 45940 740 49060
rect 200 45860 800 45940
rect 260 42740 740 45860
rect 200 42660 800 42740
rect 260 41140 740 42660
rect 200 41060 800 41140
rect 260 39540 740 41060
rect 200 39460 800 39540
rect 260 36340 740 39460
rect 200 36260 800 36340
rect 260 33140 740 36260
rect 200 33060 800 33140
rect 260 29940 740 33060
rect 200 29860 800 29940
rect 260 26740 740 29860
rect 200 26660 800 26740
rect 260 25140 740 26660
rect 200 25060 800 25140
rect 260 23540 740 25060
rect 200 23460 800 23540
rect 260 20340 740 23460
rect 200 20260 800 20340
rect 260 17140 740 20260
rect 200 17060 800 17140
rect 260 14000 740 17060
<< metal4 >>
rect 0 68400 200 69678
rect 800 68400 1000 69678
rect 0 66800 200 68200
rect 800 66800 1000 68200
rect 0 65200 200 66600
rect 800 65200 1000 66600
rect 0 63600 200 65000
rect 800 63600 1000 65000
rect 0 62000 200 63400
rect 800 62000 1000 63400
rect 0 60400 200 61800
rect 800 60400 1000 61800
rect 0 58800 200 60200
rect 800 58800 1000 60200
rect 0 57200 200 58600
rect 800 57200 1000 58600
rect 0 55600 200 57000
rect 800 55600 1000 57000
rect 0 54000 200 55400
rect 800 54000 1000 55400
rect 0 52400 200 53800
rect 800 52400 1000 53800
rect 0 50800 200 52200
rect 800 50800 1000 52200
rect 0 49200 200 50600
rect 800 49200 1000 50600
rect 0 46000 200 49000
rect 800 46000 1000 49000
rect 0 42800 200 45800
rect 800 42800 1000 45800
rect 0 41200 200 42600
rect 800 41200 1000 42600
rect 0 39600 200 41000
rect 800 39600 1000 41000
rect 0 36400 200 39400
rect 800 36400 1000 39400
rect 0 33200 200 36200
rect 800 33200 1000 36200
rect 0 30000 200 33000
rect 800 30000 1000 33000
rect 0 26800 200 29800
rect 800 26800 1000 29800
rect 0 25200 200 26600
rect 800 25200 1000 26600
rect 0 23600 200 25000
rect 800 23600 1000 25000
rect 0 20400 200 23400
rect 800 20400 1000 23400
rect 0 17200 200 20200
rect 800 17200 1000 20200
rect 0 14000 200 17000
rect 800 14000 1000 17000
<< obsm4 >>
rect 260 68340 740 69678
rect 200 68260 800 68340
rect 260 66740 740 68260
rect 200 66660 800 66740
rect 260 65140 740 66660
rect 200 65060 800 65140
rect 260 63540 740 65060
rect 200 63460 800 63540
rect 260 61940 740 63460
rect 200 61860 800 61940
rect 260 60340 740 61860
rect 200 60260 800 60340
rect 260 58740 740 60260
rect 200 58660 800 58740
rect 260 57140 740 58660
rect 200 57060 800 57140
rect 260 55540 740 57060
rect 200 55460 800 55540
rect 260 53940 740 55460
rect 200 53860 800 53940
rect 260 52340 740 53860
rect 200 52260 800 52340
rect 260 50740 740 52260
rect 200 50660 800 50740
rect 260 49140 740 50660
rect 200 49060 800 49140
rect 260 45940 740 49060
rect 200 45860 800 45940
rect 260 42740 740 45860
rect 200 42660 800 42740
rect 260 41140 740 42660
rect 200 41060 800 41140
rect 260 39540 740 41060
rect 200 39460 800 39540
rect 260 36340 740 39460
rect 200 36260 800 36340
rect 260 33140 740 36260
rect 200 33060 800 33140
rect 260 29940 740 33060
rect 200 29860 800 29940
rect 260 26740 740 29860
rect 200 26660 800 26740
rect 260 25140 740 26660
rect 200 25060 800 25140
rect 260 23540 740 25060
rect 200 23460 800 23540
rect 260 20340 740 23460
rect 200 20260 800 20340
rect 260 17140 740 20260
rect 200 17060 800 17140
rect 260 14000 740 17060
<< metal5 >>
rect 0 68400 200 69678
rect 0 66800 200 68200
rect 0 65200 200 66600
rect 0 63600 200 65000
rect 0 62000 200 63400
rect 0 60400 200 61800
rect 0 58800 200 60200
rect 0 57200 200 58600
rect 0 55600 200 57000
rect 0 54000 200 55400
rect 0 52400 200 53800
rect 0 50800 200 52200
rect 0 49200 200 50600
rect 0 46000 200 49000
rect 0 42800 200 45800
rect 0 41200 200 42600
rect 0 39600 200 41000
rect 0 36400 200 39400
rect 0 33200 200 36200
rect 0 30000 200 33000
rect 0 26800 200 29800
rect 0 25200 200 26600
rect 0 23600 200 25000
rect 0 20400 200 23400
rect 0 17200 200 20200
rect 0 14000 200 17000
rect 800 68400 1000 69678
rect 800 66800 1000 68200
rect 800 65200 1000 66600
rect 800 63600 1000 65000
rect 800 62000 1000 63400
rect 800 60400 1000 61800
rect 800 58800 1000 60200
rect 800 57200 1000 58600
rect 800 55600 1000 57000
rect 800 54000 1000 55400
rect 800 52400 1000 53800
rect 800 50800 1000 52200
rect 800 49200 1000 50600
rect 800 46000 1000 49000
rect 800 42800 1000 45800
rect 800 41200 1000 42600
rect 800 39600 1000 41000
rect 800 36400 1000 39400
rect 800 33200 1000 36200
rect 800 30000 1000 33000
rect 800 26800 1000 29800
rect 800 25200 1000 26600
rect 800 23600 1000 25000
rect 800 20400 1000 23400
rect 800 17200 1000 20200
rect 800 14000 1000 17000
<< obsm5 >>
rect 320 14000 680 69678
<< labels >>
rlabel metal5 s 800 26800 1000 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 800 30000 1000 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 800 33200 1000 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 800 36400 1000 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 800 42800 1000 45800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 800 23600 1000 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 800 41200 1000 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 800 52400 1000 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 800 54000 1000 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 800 55600 1000 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 800 58800 1000 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 800 66800 1000 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 800 26800 1000 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 800 30000 1000 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 800 33200 1000 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 800 36400 1000 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 800 42800 1000 45800 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 800 23600 1000 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 800 41200 1000 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 800 52400 1000 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 800 54000 1000 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 800 55600 1000 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 800 58800 1000 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 800 66800 1000 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 26800 1000 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 30000 1000 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 33200 1000 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 36400 1000 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 42800 1000 45800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 23600 1000 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 41200 1000 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 52400 1000 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 54000 1000 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 55600 1000 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 58800 1000 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 66800 1000 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 66800 200 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 58800 200 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 55600 200 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 54000 200 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 52400 200 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 42800 200 45800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 41200 200 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 36400 200 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 33200 200 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 30000 200 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 26800 200 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 66800 200 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 58800 200 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 55600 200 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 54000 200 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 52400 200 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 42800 200 45800 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 41200 200 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 36400 200 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 33200 200 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 30000 200 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 26800 200 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 66800 200 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 58800 200 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 55600 200 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 54000 200 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 52400 200 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 42800 200 45800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 41200 200 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 36400 200 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 33200 200 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 30000 200 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 26800 200 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 23600 200 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 23600 200 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 23600 200 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 800 14000 1000 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 800 17200 1000 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 800 20400 1000 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 800 46000 1000 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 800 25200 1000 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 800 39600 1000 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 800 57200 1000 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 800 60400 1000 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 800 65200 1000 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 800 68400 1000 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 800 14000 1000 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 800 17200 1000 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 800 20400 1000 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 800 46000 1000 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 800 25200 1000 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 800 39600 1000 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 800 57200 1000 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 800 60400 1000 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 800 65200 1000 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 800 68400 1000 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 14000 1000 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 17200 1000 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 20400 1000 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 46000 1000 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 25200 1000 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 39600 1000 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 57200 1000 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 60400 1000 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 65200 1000 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 68400 1000 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 68400 200 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 65200 200 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 60400 200 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 57200 200 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 46000 200 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 39600 200 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 25200 200 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 20400 200 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 17200 200 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 68400 200 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 65200 200 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 60400 200 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 57200 200 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 46000 200 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 39600 200 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 25200 200 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 20400 200 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 17200 200 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 68400 200 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 65200 200 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 60400 200 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 57200 200 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 46000 200 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 39600 200 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 25200 200 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 20400 200 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 17200 200 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 14000 200 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 14000 200 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 14000 200 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 800 50800 1000 52200 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 800 62000 1000 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 800 50800 1000 52200 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 800 62000 1000 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 800 50800 1000 52200 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 800 62000 1000 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 0 62000 200 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 0 62000 200 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 0 62000 200 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 0 50800 200 52200 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 0 50800 200 52200 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 0 50800 200 52200 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 800 49200 1000 50600 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 800 63600 1000 65000 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 800 49200 1000 50600 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 800 63600 1000 65000 6 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 800 49200 1000 50600 6 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 800 63600 1000 65000 6 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 0 63600 200 65000 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 0 63600 200 65000 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 0 63600 200 65000 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 0 49200 200 50600 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 0 49200 200 50600 6 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 0 49200 200 50600 6 VSS
port 4 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 1000 70000
string LEFclass PAD SPACER
string LEFsite GF_IO_Site
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 5105772
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 5096184
<< end >>
