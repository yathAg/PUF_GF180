magic
tech gf180mcuD
timestamp 1698431365
<< properties >>
string GDS_END 12325440
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 12323324
<< end >>
