magic
tech gf180mcuB
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 453 2662 1094
<< pwell >>
rect -86 -86 2662 453
<< mvnmos >>
rect 124 146 244 218
rect 348 146 468 218
rect 608 146 728 278
rect 832 146 952 278
rect 1016 146 1136 278
rect 1384 146 1504 278
rect 1568 146 1688 278
rect 1828 69 1948 333
rect 2052 69 2172 333
rect 2276 69 2396 333
<< mvpmos >>
rect 144 691 244 790
rect 358 691 458 790
rect 618 691 718 874
rect 832 691 932 874
rect 1036 691 1136 874
rect 1384 658 1484 841
rect 1588 658 1688 841
rect 1838 573 1938 939
rect 2072 573 2172 939
rect 2276 573 2376 939
<< mvndiff >>
rect 1748 278 1828 333
rect 528 218 608 278
rect 36 205 124 218
rect 36 159 49 205
rect 95 159 124 205
rect 36 146 124 159
rect 244 205 348 218
rect 244 159 273 205
rect 319 159 348 205
rect 244 146 348 159
rect 468 205 608 218
rect 468 159 497 205
rect 543 159 608 205
rect 468 146 608 159
rect 728 205 832 278
rect 728 159 757 205
rect 803 159 832 205
rect 728 146 832 159
rect 952 146 1016 278
rect 1136 205 1224 278
rect 1136 159 1165 205
rect 1211 159 1224 205
rect 1136 146 1224 159
rect 1296 265 1384 278
rect 1296 219 1309 265
rect 1355 219 1384 265
rect 1296 146 1384 219
rect 1504 146 1568 278
rect 1688 205 1828 278
rect 1688 159 1717 205
rect 1763 159 1828 205
rect 1688 146 1828 159
rect 1748 69 1828 146
rect 1948 299 2052 333
rect 1948 159 1977 299
rect 2023 159 2052 299
rect 1948 69 2052 159
rect 2172 318 2276 333
rect 2172 272 2201 318
rect 2247 272 2276 318
rect 2172 69 2276 272
rect 2396 194 2484 333
rect 2396 148 2425 194
rect 2471 148 2484 194
rect 2396 69 2484 148
<< mvpdiff >>
rect 1750 926 1838 939
rect 538 790 618 874
rect 56 767 144 790
rect 56 721 69 767
rect 115 721 144 767
rect 56 691 144 721
rect 244 691 358 790
rect 458 767 618 790
rect 458 721 487 767
rect 533 721 618 767
rect 458 691 618 721
rect 718 861 832 874
rect 718 721 757 861
rect 803 721 832 861
rect 718 691 832 721
rect 932 767 1036 874
rect 932 721 961 767
rect 1007 721 1036 767
rect 932 691 1036 721
rect 1136 828 1224 874
rect 1750 841 1763 926
rect 1136 782 1165 828
rect 1211 782 1224 828
rect 1136 691 1224 782
rect 1296 828 1384 841
rect 1296 782 1309 828
rect 1355 782 1384 828
rect 1296 658 1384 782
rect 1484 717 1588 841
rect 1484 671 1513 717
rect 1559 671 1588 717
rect 1484 658 1588 671
rect 1688 786 1763 841
rect 1809 786 1838 926
rect 1688 658 1838 786
rect 1758 573 1838 658
rect 1938 861 2072 939
rect 1938 721 1997 861
rect 2043 721 2072 861
rect 1938 573 2072 721
rect 2172 573 2276 939
rect 2376 926 2464 939
rect 2376 786 2405 926
rect 2451 786 2464 926
rect 2376 573 2464 786
<< mvndiffc >>
rect 49 159 95 205
rect 273 159 319 205
rect 497 159 543 205
rect 757 159 803 205
rect 1165 159 1211 205
rect 1309 219 1355 265
rect 1717 159 1763 205
rect 1977 159 2023 299
rect 2201 272 2247 318
rect 2425 148 2471 194
<< mvpdiffc >>
rect 69 721 115 767
rect 487 721 533 767
rect 757 721 803 861
rect 961 721 1007 767
rect 1165 782 1211 828
rect 1309 782 1355 828
rect 1513 671 1559 717
rect 1763 786 1809 926
rect 1997 721 2043 861
rect 2405 786 2451 926
<< polysilicon >>
rect 1838 939 1938 983
rect 2072 939 2172 983
rect 2276 939 2376 983
rect 618 874 718 918
rect 832 874 932 918
rect 1036 874 1136 918
rect 144 790 244 834
rect 358 790 458 834
rect 1384 841 1484 885
rect 1588 841 1688 885
rect 144 420 244 691
rect 144 374 185 420
rect 231 374 244 420
rect 144 262 244 374
rect 358 420 458 691
rect 358 374 399 420
rect 445 374 458 420
rect 358 262 458 374
rect 618 420 718 691
rect 618 374 631 420
rect 677 374 718 420
rect 618 322 718 374
rect 832 420 932 691
rect 832 374 845 420
rect 891 374 932 420
rect 832 322 932 374
rect 1036 420 1136 691
rect 1036 374 1049 420
rect 1095 374 1136 420
rect 1036 322 1136 374
rect 608 278 728 322
rect 832 278 952 322
rect 1016 278 1136 322
rect 1384 420 1484 658
rect 1384 374 1397 420
rect 1443 374 1484 420
rect 1384 322 1484 374
rect 1588 420 1688 658
rect 1588 374 1629 420
rect 1675 374 1688 420
rect 1838 420 1938 573
rect 1838 377 1851 420
rect 1588 322 1688 374
rect 1828 374 1851 377
rect 1897 377 1938 420
rect 2072 420 2172 573
rect 2072 377 2085 420
rect 1897 374 1948 377
rect 1828 333 1948 374
rect 2052 374 2085 377
rect 2131 374 2172 420
rect 2052 333 2172 374
rect 2276 420 2376 573
rect 2276 374 2289 420
rect 2335 377 2376 420
rect 2335 374 2396 377
rect 2276 333 2396 374
rect 1384 278 1504 322
rect 1568 278 1688 322
rect 124 218 244 262
rect 348 218 468 262
rect 124 102 244 146
rect 348 102 468 146
rect 608 102 728 146
rect 832 102 952 146
rect 1016 102 1136 146
rect 1384 102 1504 146
rect 1568 102 1688 146
rect 1828 25 1948 69
rect 2052 25 2172 69
rect 2276 25 2396 69
<< polycontact >>
rect 185 374 231 420
rect 399 374 445 420
rect 631 374 677 420
rect 845 374 891 420
rect 1049 374 1095 420
rect 1397 374 1443 420
rect 1629 374 1675 420
rect 1851 374 1897 420
rect 2085 374 2131 420
rect 2289 374 2335 420
<< metal1 >>
rect 0 926 2576 1098
rect 0 918 1763 926
rect 69 767 115 778
rect 69 308 115 721
rect 487 767 533 918
rect 487 710 533 721
rect 757 861 1211 872
rect 803 828 1211 861
rect 803 826 1165 828
rect 757 710 803 721
rect 961 767 1007 778
rect 1165 771 1211 782
rect 1309 828 1355 918
rect 1309 771 1355 782
rect 1401 774 1717 820
rect 1809 918 2405 926
rect 1763 775 1809 786
rect 1997 861 2043 872
rect 1007 725 1155 726
rect 1401 725 1447 774
rect 1007 721 1447 725
rect 961 680 1447 721
rect 1145 679 1447 680
rect 1513 717 1559 728
rect 260 588 1095 634
rect 260 430 306 588
rect 174 420 306 430
rect 174 374 185 420
rect 231 374 306 420
rect 174 354 306 374
rect 399 466 780 542
rect 399 420 445 466
rect 734 420 780 466
rect 1049 420 1095 588
rect 399 363 445 374
rect 491 374 631 420
rect 677 374 688 420
rect 734 374 845 420
rect 891 374 902 420
rect 491 308 537 374
rect 1049 363 1095 374
rect 1145 420 1191 679
rect 1145 374 1397 420
rect 1443 374 1454 420
rect 1145 308 1191 374
rect 1513 328 1559 671
rect 1671 652 1717 774
rect 2451 918 2576 926
rect 2405 775 2451 786
rect 2043 729 2371 744
rect 2043 721 2438 729
rect 1997 698 2438 721
rect 2337 683 2438 698
rect 1671 606 2303 652
rect 1748 466 2000 542
rect 1748 420 1794 466
rect 1954 420 2000 466
rect 2257 420 2303 606
rect 1618 374 1629 420
rect 1675 374 1794 420
rect 1840 374 1851 420
rect 1897 374 1908 420
rect 1954 374 2085 420
rect 2131 374 2142 420
rect 2257 374 2289 420
rect 2335 374 2346 420
rect 1840 328 1908 374
rect 69 262 537 308
rect 757 262 1191 308
rect 1309 282 1908 328
rect 2392 318 2438 683
rect 1977 299 2023 310
rect 1309 265 1355 282
rect 49 205 95 216
rect 49 90 95 159
rect 273 205 319 262
rect 273 148 319 159
rect 497 205 543 216
rect 497 90 543 159
rect 757 205 803 262
rect 757 148 803 159
rect 1165 205 1211 216
rect 1309 208 1355 219
rect 1165 90 1211 159
rect 1717 205 1763 216
rect 1717 90 1763 159
rect 2190 272 2201 318
rect 2247 272 2438 318
rect 2190 242 2438 272
rect 2023 159 2425 194
rect 1977 148 2425 159
rect 2471 148 2482 194
rect 0 -90 2576 90
<< labels >>
flabel metal1 s 399 466 780 542 0 FreeSans 200 0 0 0 A1
port 1 nsew default input
flabel metal1 s 260 588 1095 634 0 FreeSans 200 0 0 0 A2
port 2 nsew default input
flabel metal1 s 1748 466 2000 542 0 FreeSans 200 0 0 0 A3
port 3 nsew default input
flabel metal1 s 0 918 2576 1098 0 FreeSans 200 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 1717 90 1763 216 0 FreeSans 200 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel metal1 s 1997 744 2043 872 0 FreeSans 200 0 0 0 ZN
port 4 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 6 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 734 420 780 466 1 A1
port 1 nsew default input
rlabel metal1 s 399 420 445 466 1 A1
port 1 nsew default input
rlabel metal1 s 734 374 902 420 1 A1
port 1 nsew default input
rlabel metal1 s 399 374 445 420 1 A1
port 1 nsew default input
rlabel metal1 s 399 363 445 374 1 A1
port 1 nsew default input
rlabel metal1 s 1049 430 1095 588 1 A2
port 2 nsew default input
rlabel metal1 s 260 430 306 588 1 A2
port 2 nsew default input
rlabel metal1 s 1049 363 1095 430 1 A2
port 2 nsew default input
rlabel metal1 s 174 363 306 430 1 A2
port 2 nsew default input
rlabel metal1 s 174 354 306 363 1 A2
port 2 nsew default input
rlabel metal1 s 1954 420 2000 466 1 A3
port 3 nsew default input
rlabel metal1 s 1748 420 1794 466 1 A3
port 3 nsew default input
rlabel metal1 s 1954 374 2142 420 1 A3
port 3 nsew default input
rlabel metal1 s 1618 374 1794 420 1 A3
port 3 nsew default input
rlabel metal1 s 1997 729 2371 744 1 ZN
port 4 nsew default output
rlabel metal1 s 1997 698 2438 729 1 ZN
port 4 nsew default output
rlabel metal1 s 2337 683 2438 698 1 ZN
port 4 nsew default output
rlabel metal1 s 2392 318 2438 683 1 ZN
port 4 nsew default output
rlabel metal1 s 2190 242 2438 318 1 ZN
port 4 nsew default output
rlabel metal1 s 2405 775 2451 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1763 775 1809 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1309 775 1355 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 487 775 533 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1309 771 1355 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 487 771 533 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 487 710 533 771 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1165 90 1211 216 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 497 90 543 216 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 49 90 95 216 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 2576 90 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2576 1008
string GDS_END 467310
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 460972
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
