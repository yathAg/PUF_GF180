magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< isosubstrate >>
rect -51 -51 12313 14512
<< nwell >>
rect -51 13856 12313 14512
rect -51 8012 605 13856
rect 11657 8012 12313 13856
rect -51 7356 12313 8012
rect 601 591 11661 6463
<< psubdiff >>
rect 684 13765 11578 13787
rect 684 13719 750 13765
rect 11512 13719 11578 13765
rect 684 13611 11578 13719
rect 684 13589 1032 13611
rect 684 8279 706 13589
rect 752 13580 1032 13589
rect 752 12500 860 13580
rect 906 13565 1032 13580
rect 11230 13589 11578 13611
rect 11230 13580 11510 13589
rect 11230 13565 11356 13580
rect 906 13543 11356 13565
rect 906 12537 928 13543
rect 11334 12537 11356 13543
rect 906 12515 11356 12537
rect 906 12500 1032 12515
rect 752 12469 1032 12500
rect 11230 12500 11356 12515
rect 11402 12500 11510 13580
rect 11230 12469 11510 12500
rect 752 12361 11510 12469
rect 752 12315 891 12361
rect 11371 12315 11510 12361
rect 752 12207 11510 12315
rect 752 12176 1032 12207
rect 752 11096 860 12176
rect 906 12161 1032 12176
rect 11230 12176 11510 12207
rect 11230 12161 11356 12176
rect 906 12139 11356 12161
rect 906 11133 928 12139
rect 11334 11133 11356 12139
rect 906 11111 11356 11133
rect 906 11096 1032 11111
rect 752 11065 1032 11096
rect 11230 11096 11356 11111
rect 11402 11096 11510 12176
rect 11230 11065 11510 11096
rect 752 10957 11510 11065
rect 752 10911 891 10957
rect 11371 10911 11510 10957
rect 752 10803 11510 10911
rect 752 10772 1032 10803
rect 752 9692 860 10772
rect 906 10757 1032 10772
rect 11230 10772 11510 10803
rect 11230 10757 11356 10772
rect 906 10735 11356 10757
rect 906 9729 928 10735
rect 11334 9729 11356 10735
rect 906 9707 11356 9729
rect 906 9692 1032 9707
rect 752 9661 1032 9692
rect 11230 9692 11356 9707
rect 11402 9692 11510 10772
rect 11230 9661 11510 9692
rect 752 9553 11510 9661
rect 752 9507 891 9553
rect 11371 9507 11510 9553
rect 752 9399 11510 9507
rect 752 9368 1032 9399
rect 752 8288 860 9368
rect 906 9353 1032 9368
rect 11230 9368 11510 9399
rect 11230 9353 11356 9368
rect 906 9331 11356 9353
rect 906 8325 928 9331
rect 11334 8325 11356 9331
rect 906 8303 11356 8325
rect 906 8288 1032 8303
rect 752 8279 1032 8288
rect 684 8257 1032 8279
rect 11230 8288 11356 8303
rect 11402 8288 11510 9368
rect 11230 8279 11510 8288
rect 11556 8279 11578 13589
rect 11230 8257 11578 8279
rect 684 8149 11578 8257
rect 684 8103 750 8149
rect 11512 8103 11578 8149
rect 684 8081 11578 8103
rect 32 7000 12230 7022
rect 32 54 54 7000
rect 500 6554 608 7000
rect 11654 6554 11762 7000
rect 500 6532 11762 6554
rect 500 522 522 6532
rect 11740 522 11762 6532
rect 500 500 11762 522
rect 500 54 608 500
rect 11654 54 11762 500
rect 12208 54 12230 7000
rect 32 32 12230 54
<< nsubdiff >>
rect 32 14407 12230 14429
rect 32 7461 54 14407
rect 500 13961 608 14407
rect 11654 13961 11762 14407
rect 500 13939 11762 13961
rect 500 7929 522 13939
rect 11740 7929 11762 13939
rect 500 7907 11762 7929
rect 500 7461 608 7907
rect 11654 7461 11762 7907
rect 12208 7461 12230 14407
rect 32 7439 12230 7461
rect 684 6358 11578 6380
rect 684 6312 750 6358
rect 11512 6312 11578 6358
rect 684 6204 11578 6312
rect 684 6182 1032 6204
rect 684 872 706 6182
rect 752 6173 1032 6182
rect 752 5093 860 6173
rect 906 6158 1032 6173
rect 11230 6182 11578 6204
rect 11230 6173 11510 6182
rect 11230 6158 11356 6173
rect 906 6136 11356 6158
rect 906 5130 928 6136
rect 11334 5130 11356 6136
rect 906 5108 11356 5130
rect 906 5093 1032 5108
rect 752 5062 1032 5093
rect 11230 5093 11356 5108
rect 11402 5093 11510 6173
rect 11230 5062 11510 5093
rect 752 4954 11510 5062
rect 752 4908 891 4954
rect 11371 4908 11510 4954
rect 752 4800 11510 4908
rect 752 4769 1032 4800
rect 752 3689 860 4769
rect 906 4754 1032 4769
rect 11230 4769 11510 4800
rect 11230 4754 11356 4769
rect 906 4732 11356 4754
rect 906 3726 928 4732
rect 11334 3726 11356 4732
rect 906 3704 11356 3726
rect 906 3689 1032 3704
rect 752 3658 1032 3689
rect 11230 3689 11356 3704
rect 11402 3689 11510 4769
rect 11230 3658 11510 3689
rect 752 3550 11510 3658
rect 752 3504 891 3550
rect 11371 3504 11510 3550
rect 752 3396 11510 3504
rect 752 3365 1032 3396
rect 752 2285 860 3365
rect 906 3350 1032 3365
rect 11230 3365 11510 3396
rect 11230 3350 11356 3365
rect 906 3328 11356 3350
rect 906 2322 928 3328
rect 11334 2322 11356 3328
rect 906 2300 11356 2322
rect 906 2285 1032 2300
rect 752 2254 1032 2285
rect 11230 2285 11356 2300
rect 11402 2285 11510 3365
rect 11230 2254 11510 2285
rect 752 2146 11510 2254
rect 752 2100 891 2146
rect 11371 2100 11510 2146
rect 752 1992 11510 2100
rect 752 1961 1032 1992
rect 752 881 860 1961
rect 906 1946 1032 1961
rect 11230 1961 11510 1992
rect 11230 1946 11356 1961
rect 906 1924 11356 1946
rect 906 918 928 1924
rect 11334 918 11356 1924
rect 906 896 11356 918
rect 906 881 1032 896
rect 752 872 1032 881
rect 684 850 1032 872
rect 11230 881 11356 896
rect 11402 881 11510 1961
rect 11230 872 11510 881
rect 11556 872 11578 6182
rect 11230 850 11578 872
rect 684 742 11578 850
rect 684 696 750 742
rect 11512 696 11578 742
rect 684 674 11578 696
<< psubdiffcont >>
rect 750 13719 11512 13765
rect 706 8279 752 13589
rect 860 12500 906 13580
rect 1032 13565 11230 13611
rect 1032 12469 11230 12515
rect 11356 12500 11402 13580
rect 891 12315 11371 12361
rect 860 11096 906 12176
rect 1032 12161 11230 12207
rect 1032 11065 11230 11111
rect 11356 11096 11402 12176
rect 891 10911 11371 10957
rect 860 9692 906 10772
rect 1032 10757 11230 10803
rect 1032 9661 11230 9707
rect 11356 9692 11402 10772
rect 891 9507 11371 9553
rect 860 8288 906 9368
rect 1032 9353 11230 9399
rect 1032 8257 11230 8303
rect 11356 8288 11402 9368
rect 11510 8279 11556 13589
rect 750 8103 11512 8149
rect 54 54 500 7000
rect 608 6554 11654 7000
rect 608 54 11654 500
rect 11762 54 12208 7000
<< nsubdiffcont >>
rect 54 7461 500 14407
rect 608 13961 11654 14407
rect 608 7461 11654 7907
rect 11762 7461 12208 14407
rect 750 6312 11512 6358
rect 706 872 752 6182
rect 860 5093 906 6173
rect 1032 6158 11230 6204
rect 1032 5062 11230 5108
rect 11356 5093 11402 6173
rect 891 4908 11371 4954
rect 860 3689 906 4769
rect 1032 4754 11230 4800
rect 1032 3658 11230 3704
rect 11356 3689 11402 4769
rect 891 3504 11371 3550
rect 860 2285 906 3365
rect 1032 3350 11230 3396
rect 1032 2254 11230 2300
rect 11356 2285 11402 3365
rect 891 2100 11371 2146
rect 860 881 906 1961
rect 1032 1946 11230 1992
rect 1032 850 11230 896
rect 11356 881 11402 1961
rect 11510 872 11556 6182
rect 750 696 11512 742
<< mvpdiode >>
rect 1131 5920 11131 5933
rect 1131 5874 1144 5920
rect 11118 5874 11131 5920
rect 1131 5815 11131 5874
rect 1131 5769 1144 5815
rect 11118 5769 11131 5815
rect 1131 5710 11131 5769
rect 1131 5664 1144 5710
rect 11118 5664 11131 5710
rect 1131 5604 11131 5664
rect 1131 5558 1144 5604
rect 11118 5558 11131 5604
rect 1131 5498 11131 5558
rect 1131 5452 1144 5498
rect 11118 5452 11131 5498
rect 1131 5392 11131 5452
rect 1131 5346 1144 5392
rect 11118 5346 11131 5392
rect 1131 5333 11131 5346
rect 1131 4516 11131 4529
rect 1131 4470 1144 4516
rect 11118 4470 11131 4516
rect 1131 4411 11131 4470
rect 1131 4365 1144 4411
rect 11118 4365 11131 4411
rect 1131 4306 11131 4365
rect 1131 4260 1144 4306
rect 11118 4260 11131 4306
rect 1131 4200 11131 4260
rect 1131 4154 1144 4200
rect 11118 4154 11131 4200
rect 1131 4094 11131 4154
rect 1131 4048 1144 4094
rect 11118 4048 11131 4094
rect 1131 3988 11131 4048
rect 1131 3942 1144 3988
rect 11118 3942 11131 3988
rect 1131 3929 11131 3942
rect 1131 3112 11131 3125
rect 1131 3066 1144 3112
rect 11118 3066 11131 3112
rect 1131 3007 11131 3066
rect 1131 2961 1144 3007
rect 11118 2961 11131 3007
rect 1131 2902 11131 2961
rect 1131 2856 1144 2902
rect 11118 2856 11131 2902
rect 1131 2796 11131 2856
rect 1131 2750 1144 2796
rect 11118 2750 11131 2796
rect 1131 2690 11131 2750
rect 1131 2644 1144 2690
rect 11118 2644 11131 2690
rect 1131 2584 11131 2644
rect 1131 2538 1144 2584
rect 11118 2538 11131 2584
rect 1131 2525 11131 2538
rect 1131 1708 11131 1721
rect 1131 1662 1144 1708
rect 11118 1662 11131 1708
rect 1131 1603 11131 1662
rect 1131 1557 1144 1603
rect 11118 1557 11131 1603
rect 1131 1498 11131 1557
rect 1131 1452 1144 1498
rect 11118 1452 11131 1498
rect 1131 1392 11131 1452
rect 1131 1346 1144 1392
rect 11118 1346 11131 1392
rect 1131 1286 11131 1346
rect 1131 1240 1144 1286
rect 11118 1240 11131 1286
rect 1131 1180 11131 1240
rect 1131 1134 1144 1180
rect 11118 1134 11131 1180
rect 1131 1121 11131 1134
<< mvndiode >>
rect 1131 13327 11131 13340
rect 1131 13281 1144 13327
rect 11118 13281 11131 13327
rect 1131 13222 11131 13281
rect 1131 13176 1144 13222
rect 11118 13176 11131 13222
rect 1131 13117 11131 13176
rect 1131 13071 1144 13117
rect 11118 13071 11131 13117
rect 1131 13011 11131 13071
rect 1131 12965 1144 13011
rect 11118 12965 11131 13011
rect 1131 12905 11131 12965
rect 1131 12859 1144 12905
rect 11118 12859 11131 12905
rect 1131 12799 11131 12859
rect 1131 12753 1144 12799
rect 11118 12753 11131 12799
rect 1131 12740 11131 12753
rect 1131 11923 11131 11936
rect 1131 11877 1144 11923
rect 11118 11877 11131 11923
rect 1131 11818 11131 11877
rect 1131 11772 1144 11818
rect 11118 11772 11131 11818
rect 1131 11713 11131 11772
rect 1131 11667 1144 11713
rect 11118 11667 11131 11713
rect 1131 11607 11131 11667
rect 1131 11561 1144 11607
rect 11118 11561 11131 11607
rect 1131 11501 11131 11561
rect 1131 11455 1144 11501
rect 11118 11455 11131 11501
rect 1131 11395 11131 11455
rect 1131 11349 1144 11395
rect 11118 11349 11131 11395
rect 1131 11336 11131 11349
rect 1131 10519 11131 10532
rect 1131 10473 1144 10519
rect 11118 10473 11131 10519
rect 1131 10414 11131 10473
rect 1131 10368 1144 10414
rect 11118 10368 11131 10414
rect 1131 10309 11131 10368
rect 1131 10263 1144 10309
rect 11118 10263 11131 10309
rect 1131 10203 11131 10263
rect 1131 10157 1144 10203
rect 11118 10157 11131 10203
rect 1131 10097 11131 10157
rect 1131 10051 1144 10097
rect 11118 10051 11131 10097
rect 1131 9991 11131 10051
rect 1131 9945 1144 9991
rect 11118 9945 11131 9991
rect 1131 9932 11131 9945
rect 1131 9115 11131 9128
rect 1131 9069 1144 9115
rect 11118 9069 11131 9115
rect 1131 9010 11131 9069
rect 1131 8964 1144 9010
rect 11118 8964 11131 9010
rect 1131 8905 11131 8964
rect 1131 8859 1144 8905
rect 11118 8859 11131 8905
rect 1131 8799 11131 8859
rect 1131 8753 1144 8799
rect 11118 8753 11131 8799
rect 1131 8693 11131 8753
rect 1131 8647 1144 8693
rect 11118 8647 11131 8693
rect 1131 8587 11131 8647
rect 1131 8541 1144 8587
rect 11118 8541 11131 8587
rect 1131 8528 11131 8541
<< mvpdiodec >>
rect 1144 5874 11118 5920
rect 1144 5769 11118 5815
rect 1144 5664 11118 5710
rect 1144 5558 11118 5604
rect 1144 5452 11118 5498
rect 1144 5346 11118 5392
rect 1144 4470 11118 4516
rect 1144 4365 11118 4411
rect 1144 4260 11118 4306
rect 1144 4154 11118 4200
rect 1144 4048 11118 4094
rect 1144 3942 11118 3988
rect 1144 3066 11118 3112
rect 1144 2961 11118 3007
rect 1144 2856 11118 2902
rect 1144 2750 11118 2796
rect 1144 2644 11118 2690
rect 1144 2538 11118 2584
rect 1144 1662 11118 1708
rect 1144 1557 11118 1603
rect 1144 1452 11118 1498
rect 1144 1346 11118 1392
rect 1144 1240 11118 1286
rect 1144 1134 11118 1180
<< mvndiodec >>
rect 1144 13281 11118 13327
rect 1144 13176 11118 13222
rect 1144 13071 11118 13117
rect 1144 12965 11118 13011
rect 1144 12859 11118 12905
rect 1144 12753 11118 12799
rect 1144 11877 11118 11923
rect 1144 11772 11118 11818
rect 1144 11667 11118 11713
rect 1144 11561 11118 11607
rect 1144 11455 11118 11501
rect 1144 11349 11118 11395
rect 1144 10473 11118 10519
rect 1144 10368 11118 10414
rect 1144 10263 11118 10309
rect 1144 10157 11118 10203
rect 1144 10051 11118 10097
rect 1144 9945 11118 9991
rect 1144 9069 11118 9115
rect 1144 8964 11118 9010
rect 1144 8859 11118 8905
rect 1144 8753 11118 8799
rect 1144 8647 11118 8693
rect 1144 8541 11118 8587
<< metal1 >>
rect 43 14407 12219 14418
rect 43 7461 54 14407
rect 500 14396 608 14407
rect 11654 14396 11762 14407
rect 500 14344 605 14396
rect 11657 14344 11762 14396
rect 500 14272 608 14344
rect 11654 14272 11762 14344
rect 500 14220 605 14272
rect 11657 14220 11762 14272
rect 500 14148 608 14220
rect 11654 14148 11762 14220
rect 500 14096 605 14148
rect 11657 14096 11762 14148
rect 500 14024 608 14096
rect 11654 14024 11762 14096
rect 500 13972 605 14024
rect 11657 13972 11762 14024
rect 500 13961 608 13972
rect 11654 13961 11762 13972
rect 500 13950 11762 13961
rect 500 7918 511 13950
rect 695 13765 11567 13776
rect 695 13719 750 13765
rect 11512 13719 11567 13765
rect 695 13693 1143 13719
rect 1195 13693 1251 13719
rect 1303 13693 1359 13719
rect 1411 13693 1467 13719
rect 1519 13693 1575 13719
rect 1627 13693 3415 13719
rect 3467 13693 3523 13719
rect 3575 13693 3631 13719
rect 3683 13693 3739 13719
rect 3791 13693 3847 13719
rect 3899 13693 5700 13719
rect 5752 13693 5808 13719
rect 5860 13693 5916 13719
rect 5968 13693 6024 13719
rect 6076 13693 6186 13719
rect 6238 13693 6294 13719
rect 6346 13693 6402 13719
rect 6454 13693 6510 13719
rect 6562 13693 8363 13719
rect 8415 13693 8471 13719
rect 8523 13693 8579 13719
rect 8631 13693 8687 13719
rect 8739 13693 8795 13719
rect 8847 13693 10635 13719
rect 10687 13693 10743 13719
rect 10795 13693 10851 13719
rect 10903 13693 10959 13719
rect 11011 13693 11067 13719
rect 11119 13693 11567 13719
rect 695 13637 11567 13693
rect 695 13611 1143 13637
rect 1195 13611 1251 13637
rect 1303 13611 1359 13637
rect 1411 13611 1467 13637
rect 1519 13611 1575 13637
rect 1627 13611 3415 13637
rect 3467 13611 3523 13637
rect 3575 13611 3631 13637
rect 3683 13611 3739 13637
rect 3791 13611 3847 13637
rect 3899 13611 5700 13637
rect 5752 13611 5808 13637
rect 5860 13611 5916 13637
rect 5968 13611 6024 13637
rect 6076 13611 6186 13637
rect 6238 13611 6294 13637
rect 6346 13611 6402 13637
rect 6454 13611 6510 13637
rect 6562 13611 8363 13637
rect 8415 13611 8471 13637
rect 8523 13611 8579 13637
rect 8631 13611 8687 13637
rect 8739 13611 8795 13637
rect 8847 13611 10635 13637
rect 10687 13611 10743 13637
rect 10795 13611 10851 13637
rect 10903 13611 10959 13637
rect 11011 13611 11067 13637
rect 11119 13611 11567 13637
rect 695 13589 1032 13611
rect 695 8279 706 13589
rect 752 13580 1032 13589
rect 11230 13589 11567 13611
rect 752 12500 860 13580
rect 906 13565 1032 13580
rect 11230 13580 11510 13589
rect 11230 13565 11356 13580
rect 906 13554 11356 13565
rect 906 12526 917 13554
rect 1131 13327 11131 13340
rect 1131 13281 1144 13327
rect 11118 13281 11131 13327
rect 1131 13262 1741 13281
rect 1793 13262 1865 13281
rect 1917 13262 1989 13281
rect 2041 13262 2113 13281
rect 2165 13262 2877 13281
rect 2929 13262 3001 13281
rect 3053 13262 3125 13281
rect 3177 13262 3249 13281
rect 3301 13262 4013 13281
rect 4065 13262 4137 13281
rect 4189 13262 4261 13281
rect 4313 13262 4385 13281
rect 4437 13262 5149 13281
rect 5201 13262 5273 13281
rect 5325 13262 5397 13281
rect 5449 13262 5521 13281
rect 5573 13262 6689 13281
rect 6741 13262 6813 13281
rect 6865 13262 6937 13281
rect 6989 13262 7061 13281
rect 7113 13262 7825 13281
rect 7877 13262 7949 13281
rect 8001 13262 8073 13281
rect 8125 13262 8197 13281
rect 8249 13262 8961 13281
rect 9013 13262 9085 13281
rect 9137 13262 9209 13281
rect 9261 13262 9333 13281
rect 9385 13262 10097 13281
rect 10149 13262 10221 13281
rect 10273 13262 10345 13281
rect 10397 13262 10469 13281
rect 10521 13262 11131 13281
rect 1131 13222 11131 13262
rect 1131 13176 1144 13222
rect 11118 13176 11131 13222
rect 1131 13138 1741 13176
rect 1793 13138 1865 13176
rect 1917 13138 1989 13176
rect 2041 13138 2113 13176
rect 2165 13138 2877 13176
rect 2929 13138 3001 13176
rect 3053 13138 3125 13176
rect 3177 13138 3249 13176
rect 3301 13138 4013 13176
rect 4065 13138 4137 13176
rect 4189 13138 4261 13176
rect 4313 13138 4385 13176
rect 4437 13138 5149 13176
rect 5201 13138 5273 13176
rect 5325 13138 5397 13176
rect 5449 13138 5521 13176
rect 5573 13138 6689 13176
rect 6741 13138 6813 13176
rect 6865 13138 6937 13176
rect 6989 13138 7061 13176
rect 7113 13138 7825 13176
rect 7877 13138 7949 13176
rect 8001 13138 8073 13176
rect 8125 13138 8197 13176
rect 8249 13138 8961 13176
rect 9013 13138 9085 13176
rect 9137 13138 9209 13176
rect 9261 13138 9333 13176
rect 9385 13138 10097 13176
rect 10149 13138 10221 13176
rect 10273 13138 10345 13176
rect 10397 13138 10469 13176
rect 10521 13138 11131 13176
rect 1131 13117 11131 13138
rect 1131 13071 1144 13117
rect 11118 13071 11131 13117
rect 1131 13066 11131 13071
rect 1131 13014 1741 13066
rect 1793 13014 1865 13066
rect 1917 13014 1989 13066
rect 2041 13014 2113 13066
rect 2165 13014 2877 13066
rect 2929 13014 3001 13066
rect 3053 13014 3125 13066
rect 3177 13014 3249 13066
rect 3301 13014 4013 13066
rect 4065 13014 4137 13066
rect 4189 13014 4261 13066
rect 4313 13014 4385 13066
rect 4437 13014 5149 13066
rect 5201 13014 5273 13066
rect 5325 13014 5397 13066
rect 5449 13014 5521 13066
rect 5573 13014 6689 13066
rect 6741 13014 6813 13066
rect 6865 13014 6937 13066
rect 6989 13014 7061 13066
rect 7113 13014 7825 13066
rect 7877 13014 7949 13066
rect 8001 13014 8073 13066
rect 8125 13014 8197 13066
rect 8249 13014 8961 13066
rect 9013 13014 9085 13066
rect 9137 13014 9209 13066
rect 9261 13014 9333 13066
rect 9385 13014 10097 13066
rect 10149 13014 10221 13066
rect 10273 13014 10345 13066
rect 10397 13014 10469 13066
rect 10521 13014 11131 13066
rect 1131 13011 11131 13014
rect 1131 12965 1144 13011
rect 11118 12965 11131 13011
rect 1131 12942 11131 12965
rect 1131 12905 1741 12942
rect 1793 12905 1865 12942
rect 1917 12905 1989 12942
rect 2041 12905 2113 12942
rect 2165 12905 2877 12942
rect 2929 12905 3001 12942
rect 3053 12905 3125 12942
rect 3177 12905 3249 12942
rect 3301 12905 4013 12942
rect 4065 12905 4137 12942
rect 4189 12905 4261 12942
rect 4313 12905 4385 12942
rect 4437 12905 5149 12942
rect 5201 12905 5273 12942
rect 5325 12905 5397 12942
rect 5449 12905 5521 12942
rect 5573 12905 6689 12942
rect 6741 12905 6813 12942
rect 6865 12905 6937 12942
rect 6989 12905 7061 12942
rect 7113 12905 7825 12942
rect 7877 12905 7949 12942
rect 8001 12905 8073 12942
rect 8125 12905 8197 12942
rect 8249 12905 8961 12942
rect 9013 12905 9085 12942
rect 9137 12905 9209 12942
rect 9261 12905 9333 12942
rect 9385 12905 10097 12942
rect 10149 12905 10221 12942
rect 10273 12905 10345 12942
rect 10397 12905 10469 12942
rect 10521 12905 11131 12942
rect 1131 12859 1144 12905
rect 11118 12859 11131 12905
rect 1131 12818 11131 12859
rect 1131 12799 1741 12818
rect 1793 12799 1865 12818
rect 1917 12799 1989 12818
rect 2041 12799 2113 12818
rect 2165 12799 2877 12818
rect 2929 12799 3001 12818
rect 3053 12799 3125 12818
rect 3177 12799 3249 12818
rect 3301 12799 4013 12818
rect 4065 12799 4137 12818
rect 4189 12799 4261 12818
rect 4313 12799 4385 12818
rect 4437 12799 5149 12818
rect 5201 12799 5273 12818
rect 5325 12799 5397 12818
rect 5449 12799 5521 12818
rect 5573 12799 6689 12818
rect 6741 12799 6813 12818
rect 6865 12799 6937 12818
rect 6989 12799 7061 12818
rect 7113 12799 7825 12818
rect 7877 12799 7949 12818
rect 8001 12799 8073 12818
rect 8125 12799 8197 12818
rect 8249 12799 8961 12818
rect 9013 12799 9085 12818
rect 9137 12799 9209 12818
rect 9261 12799 9333 12818
rect 9385 12799 10097 12818
rect 10149 12799 10221 12818
rect 10273 12799 10345 12818
rect 10397 12799 10469 12818
rect 10521 12799 11131 12818
rect 1131 12753 1144 12799
rect 11118 12753 11131 12799
rect 1131 12740 11131 12753
rect 11345 12526 11356 13554
rect 906 12515 11356 12526
rect 906 12500 1032 12515
rect 752 12469 1032 12500
rect 11230 12500 11356 12515
rect 11402 12500 11510 13580
rect 11230 12469 11510 12500
rect 752 12420 1143 12469
rect 1195 12420 1251 12469
rect 1303 12420 1359 12469
rect 1411 12420 1467 12469
rect 1519 12420 1575 12469
rect 1627 12420 3415 12469
rect 3467 12420 3523 12469
rect 3575 12420 3631 12469
rect 3683 12420 3739 12469
rect 3791 12420 3847 12469
rect 3899 12420 5700 12469
rect 5752 12420 5808 12469
rect 5860 12420 5916 12469
rect 5968 12420 6024 12469
rect 6076 12420 6186 12469
rect 6238 12420 6294 12469
rect 6346 12420 6402 12469
rect 6454 12420 6510 12469
rect 6562 12420 8363 12469
rect 8415 12420 8471 12469
rect 8523 12420 8579 12469
rect 8631 12420 8687 12469
rect 8739 12420 8795 12469
rect 8847 12420 10635 12469
rect 10687 12420 10743 12469
rect 10795 12420 10851 12469
rect 10903 12420 10959 12469
rect 11011 12420 11067 12469
rect 11119 12420 11510 12469
rect 752 12364 11510 12420
rect 752 12361 1143 12364
rect 1195 12361 1251 12364
rect 1303 12361 1359 12364
rect 1411 12361 1467 12364
rect 1519 12361 1575 12364
rect 1627 12361 3415 12364
rect 3467 12361 3523 12364
rect 3575 12361 3631 12364
rect 3683 12361 3739 12364
rect 3791 12361 3847 12364
rect 3899 12361 5700 12364
rect 5752 12361 5808 12364
rect 5860 12361 5916 12364
rect 5968 12361 6024 12364
rect 6076 12361 6186 12364
rect 6238 12361 6294 12364
rect 6346 12361 6402 12364
rect 6454 12361 6510 12364
rect 6562 12361 8363 12364
rect 8415 12361 8471 12364
rect 8523 12361 8579 12364
rect 8631 12361 8687 12364
rect 8739 12361 8795 12364
rect 8847 12361 10635 12364
rect 10687 12361 10743 12364
rect 10795 12361 10851 12364
rect 10903 12361 10959 12364
rect 11011 12361 11067 12364
rect 11119 12361 11510 12364
rect 752 12315 891 12361
rect 11371 12315 11510 12361
rect 752 12312 1143 12315
rect 1195 12312 1251 12315
rect 1303 12312 1359 12315
rect 1411 12312 1467 12315
rect 1519 12312 1575 12315
rect 1627 12312 3415 12315
rect 3467 12312 3523 12315
rect 3575 12312 3631 12315
rect 3683 12312 3739 12315
rect 3791 12312 3847 12315
rect 3899 12312 5700 12315
rect 5752 12312 5808 12315
rect 5860 12312 5916 12315
rect 5968 12312 6024 12315
rect 6076 12312 6186 12315
rect 6238 12312 6294 12315
rect 6346 12312 6402 12315
rect 6454 12312 6510 12315
rect 6562 12312 8363 12315
rect 8415 12312 8471 12315
rect 8523 12312 8579 12315
rect 8631 12312 8687 12315
rect 8739 12312 8795 12315
rect 8847 12312 10635 12315
rect 10687 12312 10743 12315
rect 10795 12312 10851 12315
rect 10903 12312 10959 12315
rect 11011 12312 11067 12315
rect 11119 12312 11510 12315
rect 752 12256 11510 12312
rect 752 12207 1143 12256
rect 1195 12207 1251 12256
rect 1303 12207 1359 12256
rect 1411 12207 1467 12256
rect 1519 12207 1575 12256
rect 1627 12207 3415 12256
rect 3467 12207 3523 12256
rect 3575 12207 3631 12256
rect 3683 12207 3739 12256
rect 3791 12207 3847 12256
rect 3899 12207 5700 12256
rect 5752 12207 5808 12256
rect 5860 12207 5916 12256
rect 5968 12207 6024 12256
rect 6076 12207 6186 12256
rect 6238 12207 6294 12256
rect 6346 12207 6402 12256
rect 6454 12207 6510 12256
rect 6562 12207 8363 12256
rect 8415 12207 8471 12256
rect 8523 12207 8579 12256
rect 8631 12207 8687 12256
rect 8739 12207 8795 12256
rect 8847 12207 10635 12256
rect 10687 12207 10743 12256
rect 10795 12207 10851 12256
rect 10903 12207 10959 12256
rect 11011 12207 11067 12256
rect 11119 12207 11510 12256
rect 752 12176 1032 12207
rect 752 11096 860 12176
rect 906 12161 1032 12176
rect 11230 12176 11510 12207
rect 11230 12161 11356 12176
rect 906 12150 11356 12161
rect 906 11122 917 12150
rect 1131 11923 11131 11936
rect 1131 11877 1144 11923
rect 11118 11877 11131 11923
rect 1131 11858 1741 11877
rect 1793 11858 1865 11877
rect 1917 11858 1989 11877
rect 2041 11858 2113 11877
rect 2165 11858 2877 11877
rect 2929 11858 3001 11877
rect 3053 11858 3125 11877
rect 3177 11858 3249 11877
rect 3301 11858 4013 11877
rect 4065 11858 4137 11877
rect 4189 11858 4261 11877
rect 4313 11858 4385 11877
rect 4437 11858 5149 11877
rect 5201 11858 5273 11877
rect 5325 11858 5397 11877
rect 5449 11858 5521 11877
rect 5573 11858 6689 11877
rect 6741 11858 6813 11877
rect 6865 11858 6937 11877
rect 6989 11858 7061 11877
rect 7113 11858 7825 11877
rect 7877 11858 7949 11877
rect 8001 11858 8073 11877
rect 8125 11858 8197 11877
rect 8249 11858 8961 11877
rect 9013 11858 9085 11877
rect 9137 11858 9209 11877
rect 9261 11858 9333 11877
rect 9385 11858 10097 11877
rect 10149 11858 10221 11877
rect 10273 11858 10345 11877
rect 10397 11858 10469 11877
rect 10521 11858 11131 11877
rect 1131 11818 11131 11858
rect 1131 11772 1144 11818
rect 11118 11772 11131 11818
rect 1131 11734 1741 11772
rect 1793 11734 1865 11772
rect 1917 11734 1989 11772
rect 2041 11734 2113 11772
rect 2165 11734 2877 11772
rect 2929 11734 3001 11772
rect 3053 11734 3125 11772
rect 3177 11734 3249 11772
rect 3301 11734 4013 11772
rect 4065 11734 4137 11772
rect 4189 11734 4261 11772
rect 4313 11734 4385 11772
rect 4437 11734 5149 11772
rect 5201 11734 5273 11772
rect 5325 11734 5397 11772
rect 5449 11734 5521 11772
rect 5573 11734 6689 11772
rect 6741 11734 6813 11772
rect 6865 11734 6937 11772
rect 6989 11734 7061 11772
rect 7113 11734 7825 11772
rect 7877 11734 7949 11772
rect 8001 11734 8073 11772
rect 8125 11734 8197 11772
rect 8249 11734 8961 11772
rect 9013 11734 9085 11772
rect 9137 11734 9209 11772
rect 9261 11734 9333 11772
rect 9385 11734 10097 11772
rect 10149 11734 10221 11772
rect 10273 11734 10345 11772
rect 10397 11734 10469 11772
rect 10521 11734 11131 11772
rect 1131 11713 11131 11734
rect 1131 11667 1144 11713
rect 11118 11667 11131 11713
rect 1131 11662 11131 11667
rect 1131 11610 1741 11662
rect 1793 11610 1865 11662
rect 1917 11610 1989 11662
rect 2041 11610 2113 11662
rect 2165 11610 2877 11662
rect 2929 11610 3001 11662
rect 3053 11610 3125 11662
rect 3177 11610 3249 11662
rect 3301 11610 4013 11662
rect 4065 11610 4137 11662
rect 4189 11610 4261 11662
rect 4313 11610 4385 11662
rect 4437 11610 5149 11662
rect 5201 11610 5273 11662
rect 5325 11610 5397 11662
rect 5449 11610 5521 11662
rect 5573 11610 6689 11662
rect 6741 11610 6813 11662
rect 6865 11610 6937 11662
rect 6989 11610 7061 11662
rect 7113 11610 7825 11662
rect 7877 11610 7949 11662
rect 8001 11610 8073 11662
rect 8125 11610 8197 11662
rect 8249 11610 8961 11662
rect 9013 11610 9085 11662
rect 9137 11610 9209 11662
rect 9261 11610 9333 11662
rect 9385 11610 10097 11662
rect 10149 11610 10221 11662
rect 10273 11610 10345 11662
rect 10397 11610 10469 11662
rect 10521 11610 11131 11662
rect 1131 11607 11131 11610
rect 1131 11561 1144 11607
rect 11118 11561 11131 11607
rect 1131 11538 11131 11561
rect 1131 11501 1741 11538
rect 1793 11501 1865 11538
rect 1917 11501 1989 11538
rect 2041 11501 2113 11538
rect 2165 11501 2877 11538
rect 2929 11501 3001 11538
rect 3053 11501 3125 11538
rect 3177 11501 3249 11538
rect 3301 11501 4013 11538
rect 4065 11501 4137 11538
rect 4189 11501 4261 11538
rect 4313 11501 4385 11538
rect 4437 11501 5149 11538
rect 5201 11501 5273 11538
rect 5325 11501 5397 11538
rect 5449 11501 5521 11538
rect 5573 11501 6689 11538
rect 6741 11501 6813 11538
rect 6865 11501 6937 11538
rect 6989 11501 7061 11538
rect 7113 11501 7825 11538
rect 7877 11501 7949 11538
rect 8001 11501 8073 11538
rect 8125 11501 8197 11538
rect 8249 11501 8961 11538
rect 9013 11501 9085 11538
rect 9137 11501 9209 11538
rect 9261 11501 9333 11538
rect 9385 11501 10097 11538
rect 10149 11501 10221 11538
rect 10273 11501 10345 11538
rect 10397 11501 10469 11538
rect 10521 11501 11131 11538
rect 1131 11455 1144 11501
rect 11118 11455 11131 11501
rect 1131 11414 11131 11455
rect 1131 11395 1741 11414
rect 1793 11395 1865 11414
rect 1917 11395 1989 11414
rect 2041 11395 2113 11414
rect 2165 11395 2877 11414
rect 2929 11395 3001 11414
rect 3053 11395 3125 11414
rect 3177 11395 3249 11414
rect 3301 11395 4013 11414
rect 4065 11395 4137 11414
rect 4189 11395 4261 11414
rect 4313 11395 4385 11414
rect 4437 11395 5149 11414
rect 5201 11395 5273 11414
rect 5325 11395 5397 11414
rect 5449 11395 5521 11414
rect 5573 11395 6689 11414
rect 6741 11395 6813 11414
rect 6865 11395 6937 11414
rect 6989 11395 7061 11414
rect 7113 11395 7825 11414
rect 7877 11395 7949 11414
rect 8001 11395 8073 11414
rect 8125 11395 8197 11414
rect 8249 11395 8961 11414
rect 9013 11395 9085 11414
rect 9137 11395 9209 11414
rect 9261 11395 9333 11414
rect 9385 11395 10097 11414
rect 10149 11395 10221 11414
rect 10273 11395 10345 11414
rect 10397 11395 10469 11414
rect 10521 11395 11131 11414
rect 1131 11349 1144 11395
rect 11118 11349 11131 11395
rect 1131 11336 11131 11349
rect 11345 11122 11356 12150
rect 906 11111 11356 11122
rect 906 11096 1032 11111
rect 752 11065 1032 11096
rect 11230 11096 11356 11111
rect 11402 11096 11510 12176
rect 11230 11065 11510 11096
rect 752 11016 1143 11065
rect 1195 11016 1251 11065
rect 1303 11016 1359 11065
rect 1411 11016 1467 11065
rect 1519 11016 1575 11065
rect 1627 11016 3415 11065
rect 3467 11016 3523 11065
rect 3575 11016 3631 11065
rect 3683 11016 3739 11065
rect 3791 11016 3847 11065
rect 3899 11016 5700 11065
rect 5752 11016 5808 11065
rect 5860 11016 5916 11065
rect 5968 11016 6024 11065
rect 6076 11016 6186 11065
rect 6238 11016 6294 11065
rect 6346 11016 6402 11065
rect 6454 11016 6510 11065
rect 6562 11016 8363 11065
rect 8415 11016 8471 11065
rect 8523 11016 8579 11065
rect 8631 11016 8687 11065
rect 8739 11016 8795 11065
rect 8847 11016 10635 11065
rect 10687 11016 10743 11065
rect 10795 11016 10851 11065
rect 10903 11016 10959 11065
rect 11011 11016 11067 11065
rect 11119 11016 11510 11065
rect 752 10960 11510 11016
rect 752 10957 1143 10960
rect 1195 10957 1251 10960
rect 1303 10957 1359 10960
rect 1411 10957 1467 10960
rect 1519 10957 1575 10960
rect 1627 10957 3415 10960
rect 3467 10957 3523 10960
rect 3575 10957 3631 10960
rect 3683 10957 3739 10960
rect 3791 10957 3847 10960
rect 3899 10957 5700 10960
rect 5752 10957 5808 10960
rect 5860 10957 5916 10960
rect 5968 10957 6024 10960
rect 6076 10957 6186 10960
rect 6238 10957 6294 10960
rect 6346 10957 6402 10960
rect 6454 10957 6510 10960
rect 6562 10957 8363 10960
rect 8415 10957 8471 10960
rect 8523 10957 8579 10960
rect 8631 10957 8687 10960
rect 8739 10957 8795 10960
rect 8847 10957 10635 10960
rect 10687 10957 10743 10960
rect 10795 10957 10851 10960
rect 10903 10957 10959 10960
rect 11011 10957 11067 10960
rect 11119 10957 11510 10960
rect 752 10911 891 10957
rect 11371 10911 11510 10957
rect 752 10908 1143 10911
rect 1195 10908 1251 10911
rect 1303 10908 1359 10911
rect 1411 10908 1467 10911
rect 1519 10908 1575 10911
rect 1627 10908 3415 10911
rect 3467 10908 3523 10911
rect 3575 10908 3631 10911
rect 3683 10908 3739 10911
rect 3791 10908 3847 10911
rect 3899 10908 5700 10911
rect 5752 10908 5808 10911
rect 5860 10908 5916 10911
rect 5968 10908 6024 10911
rect 6076 10908 6186 10911
rect 6238 10908 6294 10911
rect 6346 10908 6402 10911
rect 6454 10908 6510 10911
rect 6562 10908 8363 10911
rect 8415 10908 8471 10911
rect 8523 10908 8579 10911
rect 8631 10908 8687 10911
rect 8739 10908 8795 10911
rect 8847 10908 10635 10911
rect 10687 10908 10743 10911
rect 10795 10908 10851 10911
rect 10903 10908 10959 10911
rect 11011 10908 11067 10911
rect 11119 10908 11510 10911
rect 752 10852 11510 10908
rect 752 10803 1143 10852
rect 1195 10803 1251 10852
rect 1303 10803 1359 10852
rect 1411 10803 1467 10852
rect 1519 10803 1575 10852
rect 1627 10803 3415 10852
rect 3467 10803 3523 10852
rect 3575 10803 3631 10852
rect 3683 10803 3739 10852
rect 3791 10803 3847 10852
rect 3899 10803 5700 10852
rect 5752 10803 5808 10852
rect 5860 10803 5916 10852
rect 5968 10803 6024 10852
rect 6076 10803 6186 10852
rect 6238 10803 6294 10852
rect 6346 10803 6402 10852
rect 6454 10803 6510 10852
rect 6562 10803 8363 10852
rect 8415 10803 8471 10852
rect 8523 10803 8579 10852
rect 8631 10803 8687 10852
rect 8739 10803 8795 10852
rect 8847 10803 10635 10852
rect 10687 10803 10743 10852
rect 10795 10803 10851 10852
rect 10903 10803 10959 10852
rect 11011 10803 11067 10852
rect 11119 10803 11510 10852
rect 752 10772 1032 10803
rect 752 9692 860 10772
rect 906 10757 1032 10772
rect 11230 10772 11510 10803
rect 11230 10757 11356 10772
rect 906 10746 11356 10757
rect 906 9718 917 10746
rect 1131 10519 11131 10532
rect 1131 10473 1144 10519
rect 11118 10473 11131 10519
rect 1131 10454 1741 10473
rect 1793 10454 1865 10473
rect 1917 10454 1989 10473
rect 2041 10454 2113 10473
rect 2165 10454 2877 10473
rect 2929 10454 3001 10473
rect 3053 10454 3125 10473
rect 3177 10454 3249 10473
rect 3301 10454 4013 10473
rect 4065 10454 4137 10473
rect 4189 10454 4261 10473
rect 4313 10454 4385 10473
rect 4437 10454 5149 10473
rect 5201 10454 5273 10473
rect 5325 10454 5397 10473
rect 5449 10454 5521 10473
rect 5573 10454 6689 10473
rect 6741 10454 6813 10473
rect 6865 10454 6937 10473
rect 6989 10454 7061 10473
rect 7113 10454 7825 10473
rect 7877 10454 7949 10473
rect 8001 10454 8073 10473
rect 8125 10454 8197 10473
rect 8249 10454 8961 10473
rect 9013 10454 9085 10473
rect 9137 10454 9209 10473
rect 9261 10454 9333 10473
rect 9385 10454 10097 10473
rect 10149 10454 10221 10473
rect 10273 10454 10345 10473
rect 10397 10454 10469 10473
rect 10521 10454 11131 10473
rect 1131 10414 11131 10454
rect 1131 10368 1144 10414
rect 11118 10368 11131 10414
rect 1131 10330 1741 10368
rect 1793 10330 1865 10368
rect 1917 10330 1989 10368
rect 2041 10330 2113 10368
rect 2165 10330 2877 10368
rect 2929 10330 3001 10368
rect 3053 10330 3125 10368
rect 3177 10330 3249 10368
rect 3301 10330 4013 10368
rect 4065 10330 4137 10368
rect 4189 10330 4261 10368
rect 4313 10330 4385 10368
rect 4437 10330 5149 10368
rect 5201 10330 5273 10368
rect 5325 10330 5397 10368
rect 5449 10330 5521 10368
rect 5573 10330 6689 10368
rect 6741 10330 6813 10368
rect 6865 10330 6937 10368
rect 6989 10330 7061 10368
rect 7113 10330 7825 10368
rect 7877 10330 7949 10368
rect 8001 10330 8073 10368
rect 8125 10330 8197 10368
rect 8249 10330 8961 10368
rect 9013 10330 9085 10368
rect 9137 10330 9209 10368
rect 9261 10330 9333 10368
rect 9385 10330 10097 10368
rect 10149 10330 10221 10368
rect 10273 10330 10345 10368
rect 10397 10330 10469 10368
rect 10521 10330 11131 10368
rect 1131 10309 11131 10330
rect 1131 10263 1144 10309
rect 11118 10263 11131 10309
rect 1131 10258 11131 10263
rect 1131 10206 1741 10258
rect 1793 10206 1865 10258
rect 1917 10206 1989 10258
rect 2041 10206 2113 10258
rect 2165 10206 2877 10258
rect 2929 10206 3001 10258
rect 3053 10206 3125 10258
rect 3177 10206 3249 10258
rect 3301 10206 4013 10258
rect 4065 10206 4137 10258
rect 4189 10206 4261 10258
rect 4313 10206 4385 10258
rect 4437 10206 5149 10258
rect 5201 10206 5273 10258
rect 5325 10206 5397 10258
rect 5449 10206 5521 10258
rect 5573 10206 6689 10258
rect 6741 10206 6813 10258
rect 6865 10206 6937 10258
rect 6989 10206 7061 10258
rect 7113 10206 7825 10258
rect 7877 10206 7949 10258
rect 8001 10206 8073 10258
rect 8125 10206 8197 10258
rect 8249 10206 8961 10258
rect 9013 10206 9085 10258
rect 9137 10206 9209 10258
rect 9261 10206 9333 10258
rect 9385 10206 10097 10258
rect 10149 10206 10221 10258
rect 10273 10206 10345 10258
rect 10397 10206 10469 10258
rect 10521 10206 11131 10258
rect 1131 10203 11131 10206
rect 1131 10157 1144 10203
rect 11118 10157 11131 10203
rect 1131 10134 11131 10157
rect 1131 10097 1741 10134
rect 1793 10097 1865 10134
rect 1917 10097 1989 10134
rect 2041 10097 2113 10134
rect 2165 10097 2877 10134
rect 2929 10097 3001 10134
rect 3053 10097 3125 10134
rect 3177 10097 3249 10134
rect 3301 10097 4013 10134
rect 4065 10097 4137 10134
rect 4189 10097 4261 10134
rect 4313 10097 4385 10134
rect 4437 10097 5149 10134
rect 5201 10097 5273 10134
rect 5325 10097 5397 10134
rect 5449 10097 5521 10134
rect 5573 10097 6689 10134
rect 6741 10097 6813 10134
rect 6865 10097 6937 10134
rect 6989 10097 7061 10134
rect 7113 10097 7825 10134
rect 7877 10097 7949 10134
rect 8001 10097 8073 10134
rect 8125 10097 8197 10134
rect 8249 10097 8961 10134
rect 9013 10097 9085 10134
rect 9137 10097 9209 10134
rect 9261 10097 9333 10134
rect 9385 10097 10097 10134
rect 10149 10097 10221 10134
rect 10273 10097 10345 10134
rect 10397 10097 10469 10134
rect 10521 10097 11131 10134
rect 1131 10051 1144 10097
rect 11118 10051 11131 10097
rect 1131 10010 11131 10051
rect 1131 9991 1741 10010
rect 1793 9991 1865 10010
rect 1917 9991 1989 10010
rect 2041 9991 2113 10010
rect 2165 9991 2877 10010
rect 2929 9991 3001 10010
rect 3053 9991 3125 10010
rect 3177 9991 3249 10010
rect 3301 9991 4013 10010
rect 4065 9991 4137 10010
rect 4189 9991 4261 10010
rect 4313 9991 4385 10010
rect 4437 9991 5149 10010
rect 5201 9991 5273 10010
rect 5325 9991 5397 10010
rect 5449 9991 5521 10010
rect 5573 9991 6689 10010
rect 6741 9991 6813 10010
rect 6865 9991 6937 10010
rect 6989 9991 7061 10010
rect 7113 9991 7825 10010
rect 7877 9991 7949 10010
rect 8001 9991 8073 10010
rect 8125 9991 8197 10010
rect 8249 9991 8961 10010
rect 9013 9991 9085 10010
rect 9137 9991 9209 10010
rect 9261 9991 9333 10010
rect 9385 9991 10097 10010
rect 10149 9991 10221 10010
rect 10273 9991 10345 10010
rect 10397 9991 10469 10010
rect 10521 9991 11131 10010
rect 1131 9945 1144 9991
rect 11118 9945 11131 9991
rect 1131 9932 11131 9945
rect 11345 9718 11356 10746
rect 906 9707 11356 9718
rect 906 9692 1032 9707
rect 752 9661 1032 9692
rect 11230 9692 11356 9707
rect 11402 9692 11510 10772
rect 11230 9661 11510 9692
rect 752 9612 1143 9661
rect 1195 9612 1251 9661
rect 1303 9612 1359 9661
rect 1411 9612 1467 9661
rect 1519 9612 1575 9661
rect 1627 9612 3415 9661
rect 3467 9612 3523 9661
rect 3575 9612 3631 9661
rect 3683 9612 3739 9661
rect 3791 9612 3847 9661
rect 3899 9612 5700 9661
rect 5752 9612 5808 9661
rect 5860 9612 5916 9661
rect 5968 9612 6024 9661
rect 6076 9612 6186 9661
rect 6238 9612 6294 9661
rect 6346 9612 6402 9661
rect 6454 9612 6510 9661
rect 6562 9612 8363 9661
rect 8415 9612 8471 9661
rect 8523 9612 8579 9661
rect 8631 9612 8687 9661
rect 8739 9612 8795 9661
rect 8847 9612 10635 9661
rect 10687 9612 10743 9661
rect 10795 9612 10851 9661
rect 10903 9612 10959 9661
rect 11011 9612 11067 9661
rect 11119 9612 11510 9661
rect 752 9556 11510 9612
rect 752 9553 1143 9556
rect 1195 9553 1251 9556
rect 1303 9553 1359 9556
rect 1411 9553 1467 9556
rect 1519 9553 1575 9556
rect 1627 9553 3415 9556
rect 3467 9553 3523 9556
rect 3575 9553 3631 9556
rect 3683 9553 3739 9556
rect 3791 9553 3847 9556
rect 3899 9553 5700 9556
rect 5752 9553 5808 9556
rect 5860 9553 5916 9556
rect 5968 9553 6024 9556
rect 6076 9553 6186 9556
rect 6238 9553 6294 9556
rect 6346 9553 6402 9556
rect 6454 9553 6510 9556
rect 6562 9553 8363 9556
rect 8415 9553 8471 9556
rect 8523 9553 8579 9556
rect 8631 9553 8687 9556
rect 8739 9553 8795 9556
rect 8847 9553 10635 9556
rect 10687 9553 10743 9556
rect 10795 9553 10851 9556
rect 10903 9553 10959 9556
rect 11011 9553 11067 9556
rect 11119 9553 11510 9556
rect 752 9507 891 9553
rect 11371 9507 11510 9553
rect 752 9504 1143 9507
rect 1195 9504 1251 9507
rect 1303 9504 1359 9507
rect 1411 9504 1467 9507
rect 1519 9504 1575 9507
rect 1627 9504 3415 9507
rect 3467 9504 3523 9507
rect 3575 9504 3631 9507
rect 3683 9504 3739 9507
rect 3791 9504 3847 9507
rect 3899 9504 5700 9507
rect 5752 9504 5808 9507
rect 5860 9504 5916 9507
rect 5968 9504 6024 9507
rect 6076 9504 6186 9507
rect 6238 9504 6294 9507
rect 6346 9504 6402 9507
rect 6454 9504 6510 9507
rect 6562 9504 8363 9507
rect 8415 9504 8471 9507
rect 8523 9504 8579 9507
rect 8631 9504 8687 9507
rect 8739 9504 8795 9507
rect 8847 9504 10635 9507
rect 10687 9504 10743 9507
rect 10795 9504 10851 9507
rect 10903 9504 10959 9507
rect 11011 9504 11067 9507
rect 11119 9504 11510 9507
rect 752 9448 11510 9504
rect 752 9399 1143 9448
rect 1195 9399 1251 9448
rect 1303 9399 1359 9448
rect 1411 9399 1467 9448
rect 1519 9399 1575 9448
rect 1627 9399 3415 9448
rect 3467 9399 3523 9448
rect 3575 9399 3631 9448
rect 3683 9399 3739 9448
rect 3791 9399 3847 9448
rect 3899 9399 5700 9448
rect 5752 9399 5808 9448
rect 5860 9399 5916 9448
rect 5968 9399 6024 9448
rect 6076 9399 6186 9448
rect 6238 9399 6294 9448
rect 6346 9399 6402 9448
rect 6454 9399 6510 9448
rect 6562 9399 8363 9448
rect 8415 9399 8471 9448
rect 8523 9399 8579 9448
rect 8631 9399 8687 9448
rect 8739 9399 8795 9448
rect 8847 9399 10635 9448
rect 10687 9399 10743 9448
rect 10795 9399 10851 9448
rect 10903 9399 10959 9448
rect 11011 9399 11067 9448
rect 11119 9399 11510 9448
rect 752 9368 1032 9399
rect 752 8288 860 9368
rect 906 9353 1032 9368
rect 11230 9368 11510 9399
rect 11230 9353 11356 9368
rect 906 9342 11356 9353
rect 906 8314 917 9342
rect 1131 9115 11131 9128
rect 1131 9069 1144 9115
rect 11118 9069 11131 9115
rect 1131 9050 1741 9069
rect 1793 9050 1865 9069
rect 1917 9050 1989 9069
rect 2041 9050 2113 9069
rect 2165 9050 2877 9069
rect 2929 9050 3001 9069
rect 3053 9050 3125 9069
rect 3177 9050 3249 9069
rect 3301 9050 4013 9069
rect 4065 9050 4137 9069
rect 4189 9050 4261 9069
rect 4313 9050 4385 9069
rect 4437 9050 5149 9069
rect 5201 9050 5273 9069
rect 5325 9050 5397 9069
rect 5449 9050 5521 9069
rect 5573 9050 6689 9069
rect 6741 9050 6813 9069
rect 6865 9050 6937 9069
rect 6989 9050 7061 9069
rect 7113 9050 7825 9069
rect 7877 9050 7949 9069
rect 8001 9050 8073 9069
rect 8125 9050 8197 9069
rect 8249 9050 8961 9069
rect 9013 9050 9085 9069
rect 9137 9050 9209 9069
rect 9261 9050 9333 9069
rect 9385 9050 10097 9069
rect 10149 9050 10221 9069
rect 10273 9050 10345 9069
rect 10397 9050 10469 9069
rect 10521 9050 11131 9069
rect 1131 9010 11131 9050
rect 1131 8964 1144 9010
rect 11118 8964 11131 9010
rect 1131 8926 1741 8964
rect 1793 8926 1865 8964
rect 1917 8926 1989 8964
rect 2041 8926 2113 8964
rect 2165 8926 2877 8964
rect 2929 8926 3001 8964
rect 3053 8926 3125 8964
rect 3177 8926 3249 8964
rect 3301 8926 4013 8964
rect 4065 8926 4137 8964
rect 4189 8926 4261 8964
rect 4313 8926 4385 8964
rect 4437 8926 5149 8964
rect 5201 8926 5273 8964
rect 5325 8926 5397 8964
rect 5449 8926 5521 8964
rect 5573 8926 6689 8964
rect 6741 8926 6813 8964
rect 6865 8926 6937 8964
rect 6989 8926 7061 8964
rect 7113 8926 7825 8964
rect 7877 8926 7949 8964
rect 8001 8926 8073 8964
rect 8125 8926 8197 8964
rect 8249 8926 8961 8964
rect 9013 8926 9085 8964
rect 9137 8926 9209 8964
rect 9261 8926 9333 8964
rect 9385 8926 10097 8964
rect 10149 8926 10221 8964
rect 10273 8926 10345 8964
rect 10397 8926 10469 8964
rect 10521 8926 11131 8964
rect 1131 8905 11131 8926
rect 1131 8859 1144 8905
rect 11118 8859 11131 8905
rect 1131 8854 11131 8859
rect 1131 8802 1741 8854
rect 1793 8802 1865 8854
rect 1917 8802 1989 8854
rect 2041 8802 2113 8854
rect 2165 8802 2877 8854
rect 2929 8802 3001 8854
rect 3053 8802 3125 8854
rect 3177 8802 3249 8854
rect 3301 8802 4013 8854
rect 4065 8802 4137 8854
rect 4189 8802 4261 8854
rect 4313 8802 4385 8854
rect 4437 8802 5149 8854
rect 5201 8802 5273 8854
rect 5325 8802 5397 8854
rect 5449 8802 5521 8854
rect 5573 8802 6689 8854
rect 6741 8802 6813 8854
rect 6865 8802 6937 8854
rect 6989 8802 7061 8854
rect 7113 8802 7825 8854
rect 7877 8802 7949 8854
rect 8001 8802 8073 8854
rect 8125 8802 8197 8854
rect 8249 8802 8961 8854
rect 9013 8802 9085 8854
rect 9137 8802 9209 8854
rect 9261 8802 9333 8854
rect 9385 8802 10097 8854
rect 10149 8802 10221 8854
rect 10273 8802 10345 8854
rect 10397 8802 10469 8854
rect 10521 8802 11131 8854
rect 1131 8799 11131 8802
rect 1131 8753 1144 8799
rect 11118 8753 11131 8799
rect 1131 8730 11131 8753
rect 1131 8693 1741 8730
rect 1793 8693 1865 8730
rect 1917 8693 1989 8730
rect 2041 8693 2113 8730
rect 2165 8693 2877 8730
rect 2929 8693 3001 8730
rect 3053 8693 3125 8730
rect 3177 8693 3249 8730
rect 3301 8693 4013 8730
rect 4065 8693 4137 8730
rect 4189 8693 4261 8730
rect 4313 8693 4385 8730
rect 4437 8693 5149 8730
rect 5201 8693 5273 8730
rect 5325 8693 5397 8730
rect 5449 8693 5521 8730
rect 5573 8693 6689 8730
rect 6741 8693 6813 8730
rect 6865 8693 6937 8730
rect 6989 8693 7061 8730
rect 7113 8693 7825 8730
rect 7877 8693 7949 8730
rect 8001 8693 8073 8730
rect 8125 8693 8197 8730
rect 8249 8693 8961 8730
rect 9013 8693 9085 8730
rect 9137 8693 9209 8730
rect 9261 8693 9333 8730
rect 9385 8693 10097 8730
rect 10149 8693 10221 8730
rect 10273 8693 10345 8730
rect 10397 8693 10469 8730
rect 10521 8693 11131 8730
rect 1131 8647 1144 8693
rect 11118 8647 11131 8693
rect 1131 8606 11131 8647
rect 1131 8587 1741 8606
rect 1793 8587 1865 8606
rect 1917 8587 1989 8606
rect 2041 8587 2113 8606
rect 2165 8587 2877 8606
rect 2929 8587 3001 8606
rect 3053 8587 3125 8606
rect 3177 8587 3249 8606
rect 3301 8587 4013 8606
rect 4065 8587 4137 8606
rect 4189 8587 4261 8606
rect 4313 8587 4385 8606
rect 4437 8587 5149 8606
rect 5201 8587 5273 8606
rect 5325 8587 5397 8606
rect 5449 8587 5521 8606
rect 5573 8587 6689 8606
rect 6741 8587 6813 8606
rect 6865 8587 6937 8606
rect 6989 8587 7061 8606
rect 7113 8587 7825 8606
rect 7877 8587 7949 8606
rect 8001 8587 8073 8606
rect 8125 8587 8197 8606
rect 8249 8587 8961 8606
rect 9013 8587 9085 8606
rect 9137 8587 9209 8606
rect 9261 8587 9333 8606
rect 9385 8587 10097 8606
rect 10149 8587 10221 8606
rect 10273 8587 10345 8606
rect 10397 8587 10469 8606
rect 10521 8587 11131 8606
rect 1131 8541 1144 8587
rect 11118 8541 11131 8587
rect 1131 8528 11131 8541
rect 11345 8314 11356 9342
rect 906 8303 11356 8314
rect 906 8288 1032 8303
rect 752 8279 1032 8288
rect 11230 8288 11356 8303
rect 11402 8288 11510 9368
rect 695 8257 1032 8279
rect 11230 8279 11510 8288
rect 11556 8279 11567 13589
rect 11230 8257 11567 8279
rect 695 8231 1143 8257
rect 1195 8231 1251 8257
rect 1303 8231 1359 8257
rect 1411 8231 1467 8257
rect 1519 8231 1575 8257
rect 1627 8231 3415 8257
rect 3467 8231 3523 8257
rect 3575 8231 3631 8257
rect 3683 8231 3739 8257
rect 3791 8231 3847 8257
rect 3899 8231 5700 8257
rect 5752 8231 5808 8257
rect 5860 8231 5916 8257
rect 5968 8231 6024 8257
rect 6076 8231 6186 8257
rect 6238 8231 6294 8257
rect 6346 8231 6402 8257
rect 6454 8231 6510 8257
rect 6562 8231 8363 8257
rect 8415 8231 8471 8257
rect 8523 8231 8579 8257
rect 8631 8231 8687 8257
rect 8739 8231 8795 8257
rect 8847 8231 10635 8257
rect 10687 8231 10743 8257
rect 10795 8231 10851 8257
rect 10903 8231 10959 8257
rect 11011 8231 11067 8257
rect 11119 8231 11567 8257
rect 695 8175 11567 8231
rect 695 8149 1143 8175
rect 1195 8149 1251 8175
rect 1303 8149 1359 8175
rect 1411 8149 1467 8175
rect 1519 8149 1575 8175
rect 1627 8149 3415 8175
rect 3467 8149 3523 8175
rect 3575 8149 3631 8175
rect 3683 8149 3739 8175
rect 3791 8149 3847 8175
rect 3899 8149 5700 8175
rect 5752 8149 5808 8175
rect 5860 8149 5916 8175
rect 5968 8149 6024 8175
rect 6076 8149 6186 8175
rect 6238 8149 6294 8175
rect 6346 8149 6402 8175
rect 6454 8149 6510 8175
rect 6562 8149 8363 8175
rect 8415 8149 8471 8175
rect 8523 8149 8579 8175
rect 8631 8149 8687 8175
rect 8739 8149 8795 8175
rect 8847 8149 10635 8175
rect 10687 8149 10743 8175
rect 10795 8149 10851 8175
rect 10903 8149 10959 8175
rect 11011 8149 11067 8175
rect 11119 8149 11567 8175
rect 695 8103 750 8149
rect 11512 8103 11567 8149
rect 695 8092 11567 8103
rect 11751 7918 11762 13950
rect 500 7907 11762 7918
rect 500 7896 608 7907
rect 11654 7896 11762 7907
rect 500 7844 605 7896
rect 11657 7844 11762 7896
rect 500 7772 608 7844
rect 11654 7772 11762 7844
rect 500 7720 605 7772
rect 11657 7720 11762 7772
rect 500 7648 608 7720
rect 11654 7648 11762 7720
rect 500 7596 605 7648
rect 11657 7596 11762 7648
rect 500 7524 608 7596
rect 11654 7524 11762 7596
rect 500 7472 605 7524
rect 11657 7472 11762 7524
rect 500 7461 608 7472
rect 11654 7461 11762 7472
rect 12208 7461 12219 14407
rect 43 7450 12219 7461
rect 43 7000 12219 7011
rect 43 54 54 7000
rect 500 6554 608 7000
rect 11654 6554 11762 7000
rect 500 6543 11762 6554
rect 500 511 511 6543
rect 695 6358 11567 6369
rect 695 6312 750 6358
rect 11512 6312 11567 6358
rect 695 6307 2279 6312
rect 695 6255 737 6307
rect 789 6255 845 6307
rect 897 6286 2279 6307
rect 2331 6286 2387 6312
rect 2439 6286 2495 6312
rect 2547 6286 2603 6312
rect 2655 6286 2711 6312
rect 2763 6286 4551 6312
rect 4603 6286 4659 6312
rect 4711 6286 4767 6312
rect 4819 6286 4875 6312
rect 4927 6286 4983 6312
rect 5035 6286 7227 6312
rect 7279 6286 7335 6312
rect 7387 6286 7443 6312
rect 7495 6286 7551 6312
rect 7603 6286 7659 6312
rect 7711 6286 9499 6312
rect 9551 6286 9607 6312
rect 9659 6286 9715 6312
rect 9767 6286 9823 6312
rect 9875 6286 9931 6312
rect 9983 6307 11567 6312
rect 9983 6286 11365 6307
rect 897 6255 11365 6286
rect 11417 6255 11473 6307
rect 11525 6255 11567 6307
rect 695 6230 11567 6255
rect 695 6204 2279 6230
rect 2331 6204 2387 6230
rect 2439 6204 2495 6230
rect 2547 6204 2603 6230
rect 2655 6204 2711 6230
rect 2763 6204 4551 6230
rect 4603 6204 4659 6230
rect 4711 6204 4767 6230
rect 4819 6204 4875 6230
rect 4927 6204 4983 6230
rect 5035 6204 7227 6230
rect 7279 6204 7335 6230
rect 7387 6204 7443 6230
rect 7495 6204 7551 6230
rect 7603 6204 7659 6230
rect 7711 6204 9499 6230
rect 9551 6204 9607 6230
rect 9659 6204 9715 6230
rect 9767 6204 9823 6230
rect 9875 6204 9931 6230
rect 9983 6204 11567 6230
rect 695 6199 1032 6204
rect 695 6182 737 6199
rect 695 872 706 6182
rect 789 6147 845 6199
rect 897 6173 1032 6199
rect 11230 6199 11567 6204
rect 906 6158 1032 6173
rect 11230 6173 11365 6199
rect 11230 6158 11356 6173
rect 906 6147 11356 6158
rect 11417 6147 11473 6199
rect 11525 6182 11567 6199
rect 752 6091 860 6147
rect 789 6039 845 6091
rect 752 5983 860 6039
rect 789 5931 845 5983
rect 752 5875 860 5931
rect 789 5823 845 5875
rect 752 5767 860 5823
rect 789 5715 845 5767
rect 752 5659 860 5715
rect 789 5607 845 5659
rect 752 5551 860 5607
rect 789 5499 845 5551
rect 752 5443 860 5499
rect 789 5391 845 5443
rect 752 5335 860 5391
rect 789 5283 845 5335
rect 752 5227 860 5283
rect 789 5175 845 5227
rect 752 5119 860 5175
rect 906 5119 917 6147
rect 1131 5920 11131 5933
rect 1131 5874 1144 5920
rect 11118 5874 11131 5920
rect 1131 5855 1741 5874
rect 1793 5855 1865 5874
rect 1917 5855 1989 5874
rect 2041 5855 2113 5874
rect 2165 5855 2877 5874
rect 2929 5855 3001 5874
rect 3053 5855 3125 5874
rect 3177 5855 3249 5874
rect 3301 5855 4013 5874
rect 4065 5855 4137 5874
rect 4189 5855 4261 5874
rect 4313 5855 4385 5874
rect 4437 5855 5149 5874
rect 5201 5855 5273 5874
rect 5325 5855 5397 5874
rect 5449 5855 5521 5874
rect 5573 5855 6689 5874
rect 6741 5855 6813 5874
rect 6865 5855 6937 5874
rect 6989 5855 7061 5874
rect 7113 5855 7825 5874
rect 7877 5855 7949 5874
rect 8001 5855 8073 5874
rect 8125 5855 8197 5874
rect 8249 5855 8961 5874
rect 9013 5855 9085 5874
rect 9137 5855 9209 5874
rect 9261 5855 9333 5874
rect 9385 5855 10097 5874
rect 10149 5855 10221 5874
rect 10273 5855 10345 5874
rect 10397 5855 10469 5874
rect 10521 5855 11131 5874
rect 1131 5815 11131 5855
rect 1131 5769 1144 5815
rect 11118 5769 11131 5815
rect 1131 5731 1741 5769
rect 1793 5731 1865 5769
rect 1917 5731 1989 5769
rect 2041 5731 2113 5769
rect 2165 5731 2877 5769
rect 2929 5731 3001 5769
rect 3053 5731 3125 5769
rect 3177 5731 3249 5769
rect 3301 5731 4013 5769
rect 4065 5731 4137 5769
rect 4189 5731 4261 5769
rect 4313 5731 4385 5769
rect 4437 5731 5149 5769
rect 5201 5731 5273 5769
rect 5325 5731 5397 5769
rect 5449 5731 5521 5769
rect 5573 5731 6689 5769
rect 6741 5731 6813 5769
rect 6865 5731 6937 5769
rect 6989 5731 7061 5769
rect 7113 5731 7825 5769
rect 7877 5731 7949 5769
rect 8001 5731 8073 5769
rect 8125 5731 8197 5769
rect 8249 5731 8961 5769
rect 9013 5731 9085 5769
rect 9137 5731 9209 5769
rect 9261 5731 9333 5769
rect 9385 5731 10097 5769
rect 10149 5731 10221 5769
rect 10273 5731 10345 5769
rect 10397 5731 10469 5769
rect 10521 5731 11131 5769
rect 1131 5710 11131 5731
rect 1131 5664 1144 5710
rect 11118 5664 11131 5710
rect 1131 5659 11131 5664
rect 1131 5607 1741 5659
rect 1793 5607 1865 5659
rect 1917 5607 1989 5659
rect 2041 5607 2113 5659
rect 2165 5607 2877 5659
rect 2929 5607 3001 5659
rect 3053 5607 3125 5659
rect 3177 5607 3249 5659
rect 3301 5607 4013 5659
rect 4065 5607 4137 5659
rect 4189 5607 4261 5659
rect 4313 5607 4385 5659
rect 4437 5607 5149 5659
rect 5201 5607 5273 5659
rect 5325 5607 5397 5659
rect 5449 5607 5521 5659
rect 5573 5607 6689 5659
rect 6741 5607 6813 5659
rect 6865 5607 6937 5659
rect 6989 5607 7061 5659
rect 7113 5607 7825 5659
rect 7877 5607 7949 5659
rect 8001 5607 8073 5659
rect 8125 5607 8197 5659
rect 8249 5607 8961 5659
rect 9013 5607 9085 5659
rect 9137 5607 9209 5659
rect 9261 5607 9333 5659
rect 9385 5607 10097 5659
rect 10149 5607 10221 5659
rect 10273 5607 10345 5659
rect 10397 5607 10469 5659
rect 10521 5607 11131 5659
rect 1131 5604 11131 5607
rect 1131 5558 1144 5604
rect 11118 5558 11131 5604
rect 1131 5535 11131 5558
rect 1131 5498 1741 5535
rect 1793 5498 1865 5535
rect 1917 5498 1989 5535
rect 2041 5498 2113 5535
rect 2165 5498 2877 5535
rect 2929 5498 3001 5535
rect 3053 5498 3125 5535
rect 3177 5498 3249 5535
rect 3301 5498 4013 5535
rect 4065 5498 4137 5535
rect 4189 5498 4261 5535
rect 4313 5498 4385 5535
rect 4437 5498 5149 5535
rect 5201 5498 5273 5535
rect 5325 5498 5397 5535
rect 5449 5498 5521 5535
rect 5573 5498 6689 5535
rect 6741 5498 6813 5535
rect 6865 5498 6937 5535
rect 6989 5498 7061 5535
rect 7113 5498 7825 5535
rect 7877 5498 7949 5535
rect 8001 5498 8073 5535
rect 8125 5498 8197 5535
rect 8249 5498 8961 5535
rect 9013 5498 9085 5535
rect 9137 5498 9209 5535
rect 9261 5498 9333 5535
rect 9385 5498 10097 5535
rect 10149 5498 10221 5535
rect 10273 5498 10345 5535
rect 10397 5498 10469 5535
rect 10521 5498 11131 5535
rect 1131 5452 1144 5498
rect 11118 5452 11131 5498
rect 1131 5411 11131 5452
rect 1131 5392 1741 5411
rect 1793 5392 1865 5411
rect 1917 5392 1989 5411
rect 2041 5392 2113 5411
rect 2165 5392 2877 5411
rect 2929 5392 3001 5411
rect 3053 5392 3125 5411
rect 3177 5392 3249 5411
rect 3301 5392 4013 5411
rect 4065 5392 4137 5411
rect 4189 5392 4261 5411
rect 4313 5392 4385 5411
rect 4437 5392 5149 5411
rect 5201 5392 5273 5411
rect 5325 5392 5397 5411
rect 5449 5392 5521 5411
rect 5573 5392 6689 5411
rect 6741 5392 6813 5411
rect 6865 5392 6937 5411
rect 6989 5392 7061 5411
rect 7113 5392 7825 5411
rect 7877 5392 7949 5411
rect 8001 5392 8073 5411
rect 8125 5392 8197 5411
rect 8249 5392 8961 5411
rect 9013 5392 9085 5411
rect 9137 5392 9209 5411
rect 9261 5392 9333 5411
rect 9385 5392 10097 5411
rect 10149 5392 10221 5411
rect 10273 5392 10345 5411
rect 10397 5392 10469 5411
rect 10521 5392 11131 5411
rect 1131 5346 1144 5392
rect 11118 5346 11131 5392
rect 1131 5333 11131 5346
rect 11345 5119 11356 6147
rect 11402 6091 11510 6147
rect 11417 6039 11473 6091
rect 11402 5983 11510 6039
rect 11417 5931 11473 5983
rect 11402 5875 11510 5931
rect 11417 5823 11473 5875
rect 11402 5767 11510 5823
rect 11417 5715 11473 5767
rect 11402 5659 11510 5715
rect 11417 5607 11473 5659
rect 11402 5551 11510 5607
rect 11417 5499 11473 5551
rect 11402 5443 11510 5499
rect 11417 5391 11473 5443
rect 11402 5335 11510 5391
rect 11417 5283 11473 5335
rect 11402 5227 11510 5283
rect 11417 5175 11473 5227
rect 11402 5119 11510 5175
rect 789 5067 845 5119
rect 906 5108 11356 5119
rect 906 5093 1032 5108
rect 897 5067 1032 5093
rect 752 5062 1032 5067
rect 11230 5093 11356 5108
rect 11230 5067 11365 5093
rect 11417 5067 11473 5119
rect 11230 5062 11510 5067
rect 752 5013 2279 5062
rect 2331 5013 2387 5062
rect 2439 5013 2495 5062
rect 2547 5013 2603 5062
rect 2655 5013 2711 5062
rect 2763 5013 4551 5062
rect 4603 5013 4659 5062
rect 4711 5013 4767 5062
rect 4819 5013 4875 5062
rect 4927 5013 4983 5062
rect 5035 5013 7227 5062
rect 7279 5013 7335 5062
rect 7387 5013 7443 5062
rect 7495 5013 7551 5062
rect 7603 5013 7659 5062
rect 7711 5013 9499 5062
rect 9551 5013 9607 5062
rect 9659 5013 9715 5062
rect 9767 5013 9823 5062
rect 9875 5013 9931 5062
rect 9983 5013 11510 5062
rect 752 5011 11510 5013
rect 789 4959 845 5011
rect 897 4959 11365 5011
rect 11417 4959 11473 5011
rect 752 4957 11510 4959
rect 752 4954 2279 4957
rect 2331 4954 2387 4957
rect 2439 4954 2495 4957
rect 2547 4954 2603 4957
rect 2655 4954 2711 4957
rect 2763 4954 4551 4957
rect 4603 4954 4659 4957
rect 4711 4954 4767 4957
rect 4819 4954 4875 4957
rect 4927 4954 4983 4957
rect 5035 4954 7227 4957
rect 7279 4954 7335 4957
rect 7387 4954 7443 4957
rect 7495 4954 7551 4957
rect 7603 4954 7659 4957
rect 7711 4954 9499 4957
rect 9551 4954 9607 4957
rect 9659 4954 9715 4957
rect 9767 4954 9823 4957
rect 9875 4954 9931 4957
rect 9983 4954 11510 4957
rect 752 4908 891 4954
rect 11371 4908 11510 4954
rect 752 4905 2279 4908
rect 2331 4905 2387 4908
rect 2439 4905 2495 4908
rect 2547 4905 2603 4908
rect 2655 4905 2711 4908
rect 2763 4905 4551 4908
rect 4603 4905 4659 4908
rect 4711 4905 4767 4908
rect 4819 4905 4875 4908
rect 4927 4905 4983 4908
rect 5035 4905 7227 4908
rect 7279 4905 7335 4908
rect 7387 4905 7443 4908
rect 7495 4905 7551 4908
rect 7603 4905 7659 4908
rect 7711 4905 9499 4908
rect 9551 4905 9607 4908
rect 9659 4905 9715 4908
rect 9767 4905 9823 4908
rect 9875 4905 9931 4908
rect 9983 4905 11510 4908
rect 752 4903 11510 4905
rect 789 4851 845 4903
rect 897 4851 11365 4903
rect 11417 4851 11473 4903
rect 752 4849 11510 4851
rect 752 4800 2279 4849
rect 2331 4800 2387 4849
rect 2439 4800 2495 4849
rect 2547 4800 2603 4849
rect 2655 4800 2711 4849
rect 2763 4800 4551 4849
rect 4603 4800 4659 4849
rect 4711 4800 4767 4849
rect 4819 4800 4875 4849
rect 4927 4800 4983 4849
rect 5035 4800 7227 4849
rect 7279 4800 7335 4849
rect 7387 4800 7443 4849
rect 7495 4800 7551 4849
rect 7603 4800 7659 4849
rect 7711 4800 9499 4849
rect 9551 4800 9607 4849
rect 9659 4800 9715 4849
rect 9767 4800 9823 4849
rect 9875 4800 9931 4849
rect 9983 4800 11510 4849
rect 752 4795 1032 4800
rect 789 4743 845 4795
rect 897 4769 1032 4795
rect 906 4754 1032 4769
rect 11230 4795 11510 4800
rect 11230 4769 11365 4795
rect 11230 4754 11356 4769
rect 906 4743 11356 4754
rect 11417 4743 11473 4795
rect 752 4687 860 4743
rect 789 4635 845 4687
rect 752 4579 860 4635
rect 789 4527 845 4579
rect 752 4471 860 4527
rect 789 4419 845 4471
rect 752 4363 860 4419
rect 789 4311 845 4363
rect 752 4255 860 4311
rect 789 4203 845 4255
rect 752 4147 860 4203
rect 789 4095 845 4147
rect 752 4039 860 4095
rect 789 3987 845 4039
rect 752 3931 860 3987
rect 789 3879 845 3931
rect 752 3823 860 3879
rect 789 3771 845 3823
rect 752 3715 860 3771
rect 906 3715 917 4743
rect 1131 4516 11131 4529
rect 1131 4470 1144 4516
rect 11118 4470 11131 4516
rect 1131 4451 1741 4470
rect 1793 4451 1865 4470
rect 1917 4451 1989 4470
rect 2041 4451 2113 4470
rect 2165 4451 2877 4470
rect 2929 4451 3001 4470
rect 3053 4451 3125 4470
rect 3177 4451 3249 4470
rect 3301 4451 4013 4470
rect 4065 4451 4137 4470
rect 4189 4451 4261 4470
rect 4313 4451 4385 4470
rect 4437 4451 5149 4470
rect 5201 4451 5273 4470
rect 5325 4451 5397 4470
rect 5449 4451 5521 4470
rect 5573 4451 6689 4470
rect 6741 4451 6813 4470
rect 6865 4451 6937 4470
rect 6989 4451 7061 4470
rect 7113 4451 7825 4470
rect 7877 4451 7949 4470
rect 8001 4451 8073 4470
rect 8125 4451 8197 4470
rect 8249 4451 8961 4470
rect 9013 4451 9085 4470
rect 9137 4451 9209 4470
rect 9261 4451 9333 4470
rect 9385 4451 10097 4470
rect 10149 4451 10221 4470
rect 10273 4451 10345 4470
rect 10397 4451 10469 4470
rect 10521 4451 11131 4470
rect 1131 4411 11131 4451
rect 1131 4365 1144 4411
rect 11118 4365 11131 4411
rect 1131 4327 1741 4365
rect 1793 4327 1865 4365
rect 1917 4327 1989 4365
rect 2041 4327 2113 4365
rect 2165 4327 2877 4365
rect 2929 4327 3001 4365
rect 3053 4327 3125 4365
rect 3177 4327 3249 4365
rect 3301 4327 4013 4365
rect 4065 4327 4137 4365
rect 4189 4327 4261 4365
rect 4313 4327 4385 4365
rect 4437 4327 5149 4365
rect 5201 4327 5273 4365
rect 5325 4327 5397 4365
rect 5449 4327 5521 4365
rect 5573 4327 6689 4365
rect 6741 4327 6813 4365
rect 6865 4327 6937 4365
rect 6989 4327 7061 4365
rect 7113 4327 7825 4365
rect 7877 4327 7949 4365
rect 8001 4327 8073 4365
rect 8125 4327 8197 4365
rect 8249 4327 8961 4365
rect 9013 4327 9085 4365
rect 9137 4327 9209 4365
rect 9261 4327 9333 4365
rect 9385 4327 10097 4365
rect 10149 4327 10221 4365
rect 10273 4327 10345 4365
rect 10397 4327 10469 4365
rect 10521 4327 11131 4365
rect 1131 4306 11131 4327
rect 1131 4260 1144 4306
rect 11118 4260 11131 4306
rect 1131 4255 11131 4260
rect 1131 4203 1741 4255
rect 1793 4203 1865 4255
rect 1917 4203 1989 4255
rect 2041 4203 2113 4255
rect 2165 4203 2877 4255
rect 2929 4203 3001 4255
rect 3053 4203 3125 4255
rect 3177 4203 3249 4255
rect 3301 4203 4013 4255
rect 4065 4203 4137 4255
rect 4189 4203 4261 4255
rect 4313 4203 4385 4255
rect 4437 4203 5149 4255
rect 5201 4203 5273 4255
rect 5325 4203 5397 4255
rect 5449 4203 5521 4255
rect 5573 4203 6689 4255
rect 6741 4203 6813 4255
rect 6865 4203 6937 4255
rect 6989 4203 7061 4255
rect 7113 4203 7825 4255
rect 7877 4203 7949 4255
rect 8001 4203 8073 4255
rect 8125 4203 8197 4255
rect 8249 4203 8961 4255
rect 9013 4203 9085 4255
rect 9137 4203 9209 4255
rect 9261 4203 9333 4255
rect 9385 4203 10097 4255
rect 10149 4203 10221 4255
rect 10273 4203 10345 4255
rect 10397 4203 10469 4255
rect 10521 4203 11131 4255
rect 1131 4200 11131 4203
rect 1131 4154 1144 4200
rect 11118 4154 11131 4200
rect 1131 4131 11131 4154
rect 1131 4094 1741 4131
rect 1793 4094 1865 4131
rect 1917 4094 1989 4131
rect 2041 4094 2113 4131
rect 2165 4094 2877 4131
rect 2929 4094 3001 4131
rect 3053 4094 3125 4131
rect 3177 4094 3249 4131
rect 3301 4094 4013 4131
rect 4065 4094 4137 4131
rect 4189 4094 4261 4131
rect 4313 4094 4385 4131
rect 4437 4094 5149 4131
rect 5201 4094 5273 4131
rect 5325 4094 5397 4131
rect 5449 4094 5521 4131
rect 5573 4094 6689 4131
rect 6741 4094 6813 4131
rect 6865 4094 6937 4131
rect 6989 4094 7061 4131
rect 7113 4094 7825 4131
rect 7877 4094 7949 4131
rect 8001 4094 8073 4131
rect 8125 4094 8197 4131
rect 8249 4094 8961 4131
rect 9013 4094 9085 4131
rect 9137 4094 9209 4131
rect 9261 4094 9333 4131
rect 9385 4094 10097 4131
rect 10149 4094 10221 4131
rect 10273 4094 10345 4131
rect 10397 4094 10469 4131
rect 10521 4094 11131 4131
rect 1131 4048 1144 4094
rect 11118 4048 11131 4094
rect 1131 4007 11131 4048
rect 1131 3988 1741 4007
rect 1793 3988 1865 4007
rect 1917 3988 1989 4007
rect 2041 3988 2113 4007
rect 2165 3988 2877 4007
rect 2929 3988 3001 4007
rect 3053 3988 3125 4007
rect 3177 3988 3249 4007
rect 3301 3988 4013 4007
rect 4065 3988 4137 4007
rect 4189 3988 4261 4007
rect 4313 3988 4385 4007
rect 4437 3988 5149 4007
rect 5201 3988 5273 4007
rect 5325 3988 5397 4007
rect 5449 3988 5521 4007
rect 5573 3988 6689 4007
rect 6741 3988 6813 4007
rect 6865 3988 6937 4007
rect 6989 3988 7061 4007
rect 7113 3988 7825 4007
rect 7877 3988 7949 4007
rect 8001 3988 8073 4007
rect 8125 3988 8197 4007
rect 8249 3988 8961 4007
rect 9013 3988 9085 4007
rect 9137 3988 9209 4007
rect 9261 3988 9333 4007
rect 9385 3988 10097 4007
rect 10149 3988 10221 4007
rect 10273 3988 10345 4007
rect 10397 3988 10469 4007
rect 10521 3988 11131 4007
rect 1131 3942 1144 3988
rect 11118 3942 11131 3988
rect 1131 3929 11131 3942
rect 11345 3715 11356 4743
rect 11402 4687 11510 4743
rect 11417 4635 11473 4687
rect 11402 4579 11510 4635
rect 11417 4527 11473 4579
rect 11402 4471 11510 4527
rect 11417 4419 11473 4471
rect 11402 4363 11510 4419
rect 11417 4311 11473 4363
rect 11402 4255 11510 4311
rect 11417 4203 11473 4255
rect 11402 4147 11510 4203
rect 11417 4095 11473 4147
rect 11402 4039 11510 4095
rect 11417 3987 11473 4039
rect 11402 3931 11510 3987
rect 11417 3879 11473 3931
rect 11402 3823 11510 3879
rect 11417 3771 11473 3823
rect 11402 3715 11510 3771
rect 789 3663 845 3715
rect 906 3704 11356 3715
rect 906 3689 1032 3704
rect 897 3663 1032 3689
rect 752 3658 1032 3663
rect 11230 3689 11356 3704
rect 11230 3663 11365 3689
rect 11417 3663 11473 3715
rect 11230 3658 11510 3663
rect 752 3609 2279 3658
rect 2331 3609 2387 3658
rect 2439 3609 2495 3658
rect 2547 3609 2603 3658
rect 2655 3609 2711 3658
rect 2763 3609 4551 3658
rect 4603 3609 4659 3658
rect 4711 3609 4767 3658
rect 4819 3609 4875 3658
rect 4927 3609 4983 3658
rect 5035 3609 7227 3658
rect 7279 3609 7335 3658
rect 7387 3609 7443 3658
rect 7495 3609 7551 3658
rect 7603 3609 7659 3658
rect 7711 3609 9499 3658
rect 9551 3609 9607 3658
rect 9659 3609 9715 3658
rect 9767 3609 9823 3658
rect 9875 3609 9931 3658
rect 9983 3609 11510 3658
rect 752 3607 11510 3609
rect 789 3555 845 3607
rect 897 3555 11365 3607
rect 11417 3555 11473 3607
rect 752 3553 11510 3555
rect 752 3550 2279 3553
rect 2331 3550 2387 3553
rect 2439 3550 2495 3553
rect 2547 3550 2603 3553
rect 2655 3550 2711 3553
rect 2763 3550 4551 3553
rect 4603 3550 4659 3553
rect 4711 3550 4767 3553
rect 4819 3550 4875 3553
rect 4927 3550 4983 3553
rect 5035 3550 7227 3553
rect 7279 3550 7335 3553
rect 7387 3550 7443 3553
rect 7495 3550 7551 3553
rect 7603 3550 7659 3553
rect 7711 3550 9499 3553
rect 9551 3550 9607 3553
rect 9659 3550 9715 3553
rect 9767 3550 9823 3553
rect 9875 3550 9931 3553
rect 9983 3550 11510 3553
rect 752 3504 891 3550
rect 11371 3504 11510 3550
rect 752 3501 2279 3504
rect 2331 3501 2387 3504
rect 2439 3501 2495 3504
rect 2547 3501 2603 3504
rect 2655 3501 2711 3504
rect 2763 3501 4551 3504
rect 4603 3501 4659 3504
rect 4711 3501 4767 3504
rect 4819 3501 4875 3504
rect 4927 3501 4983 3504
rect 5035 3501 7227 3504
rect 7279 3501 7335 3504
rect 7387 3501 7443 3504
rect 7495 3501 7551 3504
rect 7603 3501 7659 3504
rect 7711 3501 9499 3504
rect 9551 3501 9607 3504
rect 9659 3501 9715 3504
rect 9767 3501 9823 3504
rect 9875 3501 9931 3504
rect 9983 3501 11510 3504
rect 752 3499 11510 3501
rect 789 3447 845 3499
rect 897 3447 11365 3499
rect 11417 3447 11473 3499
rect 752 3445 11510 3447
rect 752 3396 2279 3445
rect 2331 3396 2387 3445
rect 2439 3396 2495 3445
rect 2547 3396 2603 3445
rect 2655 3396 2711 3445
rect 2763 3396 4551 3445
rect 4603 3396 4659 3445
rect 4711 3396 4767 3445
rect 4819 3396 4875 3445
rect 4927 3396 4983 3445
rect 5035 3396 7227 3445
rect 7279 3396 7335 3445
rect 7387 3396 7443 3445
rect 7495 3396 7551 3445
rect 7603 3396 7659 3445
rect 7711 3396 9499 3445
rect 9551 3396 9607 3445
rect 9659 3396 9715 3445
rect 9767 3396 9823 3445
rect 9875 3396 9931 3445
rect 9983 3396 11510 3445
rect 752 3391 1032 3396
rect 789 3339 845 3391
rect 897 3365 1032 3391
rect 906 3350 1032 3365
rect 11230 3391 11510 3396
rect 11230 3365 11365 3391
rect 11230 3350 11356 3365
rect 906 3339 11356 3350
rect 11417 3339 11473 3391
rect 752 3283 860 3339
rect 789 3231 845 3283
rect 752 3175 860 3231
rect 789 3123 845 3175
rect 752 3067 860 3123
rect 789 3015 845 3067
rect 752 2959 860 3015
rect 789 2907 845 2959
rect 752 2851 860 2907
rect 789 2799 845 2851
rect 752 2743 860 2799
rect 789 2691 845 2743
rect 752 2635 860 2691
rect 789 2583 845 2635
rect 752 2527 860 2583
rect 789 2475 845 2527
rect 752 2419 860 2475
rect 789 2367 845 2419
rect 752 2311 860 2367
rect 906 2311 917 3339
rect 1131 3112 11131 3125
rect 1131 3066 1144 3112
rect 11118 3066 11131 3112
rect 1131 3047 1741 3066
rect 1793 3047 1865 3066
rect 1917 3047 1989 3066
rect 2041 3047 2113 3066
rect 2165 3047 2877 3066
rect 2929 3047 3001 3066
rect 3053 3047 3125 3066
rect 3177 3047 3249 3066
rect 3301 3047 4013 3066
rect 4065 3047 4137 3066
rect 4189 3047 4261 3066
rect 4313 3047 4385 3066
rect 4437 3047 5149 3066
rect 5201 3047 5273 3066
rect 5325 3047 5397 3066
rect 5449 3047 5521 3066
rect 5573 3047 6689 3066
rect 6741 3047 6813 3066
rect 6865 3047 6937 3066
rect 6989 3047 7061 3066
rect 7113 3047 7825 3066
rect 7877 3047 7949 3066
rect 8001 3047 8073 3066
rect 8125 3047 8197 3066
rect 8249 3047 8961 3066
rect 9013 3047 9085 3066
rect 9137 3047 9209 3066
rect 9261 3047 9333 3066
rect 9385 3047 10097 3066
rect 10149 3047 10221 3066
rect 10273 3047 10345 3066
rect 10397 3047 10469 3066
rect 10521 3047 11131 3066
rect 1131 3007 11131 3047
rect 1131 2961 1144 3007
rect 11118 2961 11131 3007
rect 1131 2923 1741 2961
rect 1793 2923 1865 2961
rect 1917 2923 1989 2961
rect 2041 2923 2113 2961
rect 2165 2923 2877 2961
rect 2929 2923 3001 2961
rect 3053 2923 3125 2961
rect 3177 2923 3249 2961
rect 3301 2923 4013 2961
rect 4065 2923 4137 2961
rect 4189 2923 4261 2961
rect 4313 2923 4385 2961
rect 4437 2923 5149 2961
rect 5201 2923 5273 2961
rect 5325 2923 5397 2961
rect 5449 2923 5521 2961
rect 5573 2923 6689 2961
rect 6741 2923 6813 2961
rect 6865 2923 6937 2961
rect 6989 2923 7061 2961
rect 7113 2923 7825 2961
rect 7877 2923 7949 2961
rect 8001 2923 8073 2961
rect 8125 2923 8197 2961
rect 8249 2923 8961 2961
rect 9013 2923 9085 2961
rect 9137 2923 9209 2961
rect 9261 2923 9333 2961
rect 9385 2923 10097 2961
rect 10149 2923 10221 2961
rect 10273 2923 10345 2961
rect 10397 2923 10469 2961
rect 10521 2923 11131 2961
rect 1131 2902 11131 2923
rect 1131 2856 1144 2902
rect 11118 2856 11131 2902
rect 1131 2851 11131 2856
rect 1131 2799 1741 2851
rect 1793 2799 1865 2851
rect 1917 2799 1989 2851
rect 2041 2799 2113 2851
rect 2165 2799 2877 2851
rect 2929 2799 3001 2851
rect 3053 2799 3125 2851
rect 3177 2799 3249 2851
rect 3301 2799 4013 2851
rect 4065 2799 4137 2851
rect 4189 2799 4261 2851
rect 4313 2799 4385 2851
rect 4437 2799 5149 2851
rect 5201 2799 5273 2851
rect 5325 2799 5397 2851
rect 5449 2799 5521 2851
rect 5573 2799 6689 2851
rect 6741 2799 6813 2851
rect 6865 2799 6937 2851
rect 6989 2799 7061 2851
rect 7113 2799 7825 2851
rect 7877 2799 7949 2851
rect 8001 2799 8073 2851
rect 8125 2799 8197 2851
rect 8249 2799 8961 2851
rect 9013 2799 9085 2851
rect 9137 2799 9209 2851
rect 9261 2799 9333 2851
rect 9385 2799 10097 2851
rect 10149 2799 10221 2851
rect 10273 2799 10345 2851
rect 10397 2799 10469 2851
rect 10521 2799 11131 2851
rect 1131 2796 11131 2799
rect 1131 2750 1144 2796
rect 11118 2750 11131 2796
rect 1131 2727 11131 2750
rect 1131 2690 1741 2727
rect 1793 2690 1865 2727
rect 1917 2690 1989 2727
rect 2041 2690 2113 2727
rect 2165 2690 2877 2727
rect 2929 2690 3001 2727
rect 3053 2690 3125 2727
rect 3177 2690 3249 2727
rect 3301 2690 4013 2727
rect 4065 2690 4137 2727
rect 4189 2690 4261 2727
rect 4313 2690 4385 2727
rect 4437 2690 5149 2727
rect 5201 2690 5273 2727
rect 5325 2690 5397 2727
rect 5449 2690 5521 2727
rect 5573 2690 6689 2727
rect 6741 2690 6813 2727
rect 6865 2690 6937 2727
rect 6989 2690 7061 2727
rect 7113 2690 7825 2727
rect 7877 2690 7949 2727
rect 8001 2690 8073 2727
rect 8125 2690 8197 2727
rect 8249 2690 8961 2727
rect 9013 2690 9085 2727
rect 9137 2690 9209 2727
rect 9261 2690 9333 2727
rect 9385 2690 10097 2727
rect 10149 2690 10221 2727
rect 10273 2690 10345 2727
rect 10397 2690 10469 2727
rect 10521 2690 11131 2727
rect 1131 2644 1144 2690
rect 11118 2644 11131 2690
rect 1131 2603 11131 2644
rect 1131 2584 1741 2603
rect 1793 2584 1865 2603
rect 1917 2584 1989 2603
rect 2041 2584 2113 2603
rect 2165 2584 2877 2603
rect 2929 2584 3001 2603
rect 3053 2584 3125 2603
rect 3177 2584 3249 2603
rect 3301 2584 4013 2603
rect 4065 2584 4137 2603
rect 4189 2584 4261 2603
rect 4313 2584 4385 2603
rect 4437 2584 5149 2603
rect 5201 2584 5273 2603
rect 5325 2584 5397 2603
rect 5449 2584 5521 2603
rect 5573 2584 6689 2603
rect 6741 2584 6813 2603
rect 6865 2584 6937 2603
rect 6989 2584 7061 2603
rect 7113 2584 7825 2603
rect 7877 2584 7949 2603
rect 8001 2584 8073 2603
rect 8125 2584 8197 2603
rect 8249 2584 8961 2603
rect 9013 2584 9085 2603
rect 9137 2584 9209 2603
rect 9261 2584 9333 2603
rect 9385 2584 10097 2603
rect 10149 2584 10221 2603
rect 10273 2584 10345 2603
rect 10397 2584 10469 2603
rect 10521 2584 11131 2603
rect 1131 2538 1144 2584
rect 11118 2538 11131 2584
rect 1131 2525 11131 2538
rect 11345 2311 11356 3339
rect 11402 3283 11510 3339
rect 11417 3231 11473 3283
rect 11402 3175 11510 3231
rect 11417 3123 11473 3175
rect 11402 3067 11510 3123
rect 11417 3015 11473 3067
rect 11402 2959 11510 3015
rect 11417 2907 11473 2959
rect 11402 2851 11510 2907
rect 11417 2799 11473 2851
rect 11402 2743 11510 2799
rect 11417 2691 11473 2743
rect 11402 2635 11510 2691
rect 11417 2583 11473 2635
rect 11402 2527 11510 2583
rect 11417 2475 11473 2527
rect 11402 2419 11510 2475
rect 11417 2367 11473 2419
rect 11402 2311 11510 2367
rect 789 2259 845 2311
rect 906 2300 11356 2311
rect 906 2285 1032 2300
rect 897 2259 1032 2285
rect 752 2254 1032 2259
rect 11230 2285 11356 2300
rect 11230 2259 11365 2285
rect 11417 2259 11473 2311
rect 11230 2254 11510 2259
rect 752 2205 2279 2254
rect 2331 2205 2387 2254
rect 2439 2205 2495 2254
rect 2547 2205 2603 2254
rect 2655 2205 2711 2254
rect 2763 2205 4551 2254
rect 4603 2205 4659 2254
rect 4711 2205 4767 2254
rect 4819 2205 4875 2254
rect 4927 2205 4983 2254
rect 5035 2205 7227 2254
rect 7279 2205 7335 2254
rect 7387 2205 7443 2254
rect 7495 2205 7551 2254
rect 7603 2205 7659 2254
rect 7711 2205 9499 2254
rect 9551 2205 9607 2254
rect 9659 2205 9715 2254
rect 9767 2205 9823 2254
rect 9875 2205 9931 2254
rect 9983 2205 11510 2254
rect 752 2203 11510 2205
rect 789 2151 845 2203
rect 897 2151 11365 2203
rect 11417 2151 11473 2203
rect 752 2149 11510 2151
rect 752 2146 2279 2149
rect 2331 2146 2387 2149
rect 2439 2146 2495 2149
rect 2547 2146 2603 2149
rect 2655 2146 2711 2149
rect 2763 2146 4551 2149
rect 4603 2146 4659 2149
rect 4711 2146 4767 2149
rect 4819 2146 4875 2149
rect 4927 2146 4983 2149
rect 5035 2146 7227 2149
rect 7279 2146 7335 2149
rect 7387 2146 7443 2149
rect 7495 2146 7551 2149
rect 7603 2146 7659 2149
rect 7711 2146 9499 2149
rect 9551 2146 9607 2149
rect 9659 2146 9715 2149
rect 9767 2146 9823 2149
rect 9875 2146 9931 2149
rect 9983 2146 11510 2149
rect 752 2100 891 2146
rect 11371 2100 11510 2146
rect 752 2097 2279 2100
rect 2331 2097 2387 2100
rect 2439 2097 2495 2100
rect 2547 2097 2603 2100
rect 2655 2097 2711 2100
rect 2763 2097 4551 2100
rect 4603 2097 4659 2100
rect 4711 2097 4767 2100
rect 4819 2097 4875 2100
rect 4927 2097 4983 2100
rect 5035 2097 7227 2100
rect 7279 2097 7335 2100
rect 7387 2097 7443 2100
rect 7495 2097 7551 2100
rect 7603 2097 7659 2100
rect 7711 2097 9499 2100
rect 9551 2097 9607 2100
rect 9659 2097 9715 2100
rect 9767 2097 9823 2100
rect 9875 2097 9931 2100
rect 9983 2097 11510 2100
rect 752 2095 11510 2097
rect 789 2043 845 2095
rect 897 2043 11365 2095
rect 11417 2043 11473 2095
rect 752 2041 11510 2043
rect 752 1992 2279 2041
rect 2331 1992 2387 2041
rect 2439 1992 2495 2041
rect 2547 1992 2603 2041
rect 2655 1992 2711 2041
rect 2763 1992 4551 2041
rect 4603 1992 4659 2041
rect 4711 1992 4767 2041
rect 4819 1992 4875 2041
rect 4927 1992 4983 2041
rect 5035 1992 7227 2041
rect 7279 1992 7335 2041
rect 7387 1992 7443 2041
rect 7495 1992 7551 2041
rect 7603 1992 7659 2041
rect 7711 1992 9499 2041
rect 9551 1992 9607 2041
rect 9659 1992 9715 2041
rect 9767 1992 9823 2041
rect 9875 1992 9931 2041
rect 9983 1992 11510 2041
rect 752 1987 1032 1992
rect 789 1935 845 1987
rect 897 1961 1032 1987
rect 906 1946 1032 1961
rect 11230 1987 11510 1992
rect 11230 1961 11365 1987
rect 11230 1946 11356 1961
rect 906 1935 11356 1946
rect 11417 1935 11473 1987
rect 752 1879 860 1935
rect 789 1827 845 1879
rect 752 1771 860 1827
rect 789 1719 845 1771
rect 752 1663 860 1719
rect 789 1611 845 1663
rect 752 1555 860 1611
rect 789 1503 845 1555
rect 752 1447 860 1503
rect 789 1395 845 1447
rect 752 1339 860 1395
rect 789 1287 845 1339
rect 752 1231 860 1287
rect 789 1179 845 1231
rect 752 1123 860 1179
rect 789 1071 845 1123
rect 752 1015 860 1071
rect 789 963 845 1015
rect 752 907 860 963
rect 906 907 917 1935
rect 1131 1708 11131 1721
rect 1131 1662 1144 1708
rect 11118 1662 11131 1708
rect 1131 1643 1741 1662
rect 1793 1643 1865 1662
rect 1917 1643 1989 1662
rect 2041 1643 2113 1662
rect 2165 1643 2877 1662
rect 2929 1643 3001 1662
rect 3053 1643 3125 1662
rect 3177 1643 3249 1662
rect 3301 1643 4013 1662
rect 4065 1643 4137 1662
rect 4189 1643 4261 1662
rect 4313 1643 4385 1662
rect 4437 1643 5149 1662
rect 5201 1643 5273 1662
rect 5325 1643 5397 1662
rect 5449 1643 5521 1662
rect 5573 1643 6689 1662
rect 6741 1643 6813 1662
rect 6865 1643 6937 1662
rect 6989 1643 7061 1662
rect 7113 1643 7825 1662
rect 7877 1643 7949 1662
rect 8001 1643 8073 1662
rect 8125 1643 8197 1662
rect 8249 1643 8961 1662
rect 9013 1643 9085 1662
rect 9137 1643 9209 1662
rect 9261 1643 9333 1662
rect 9385 1643 10097 1662
rect 10149 1643 10221 1662
rect 10273 1643 10345 1662
rect 10397 1643 10469 1662
rect 10521 1643 11131 1662
rect 1131 1603 11131 1643
rect 1131 1557 1144 1603
rect 11118 1557 11131 1603
rect 1131 1519 1741 1557
rect 1793 1519 1865 1557
rect 1917 1519 1989 1557
rect 2041 1519 2113 1557
rect 2165 1519 2877 1557
rect 2929 1519 3001 1557
rect 3053 1519 3125 1557
rect 3177 1519 3249 1557
rect 3301 1519 4013 1557
rect 4065 1519 4137 1557
rect 4189 1519 4261 1557
rect 4313 1519 4385 1557
rect 4437 1519 5149 1557
rect 5201 1519 5273 1557
rect 5325 1519 5397 1557
rect 5449 1519 5521 1557
rect 5573 1519 6689 1557
rect 6741 1519 6813 1557
rect 6865 1519 6937 1557
rect 6989 1519 7061 1557
rect 7113 1519 7825 1557
rect 7877 1519 7949 1557
rect 8001 1519 8073 1557
rect 8125 1519 8197 1557
rect 8249 1519 8961 1557
rect 9013 1519 9085 1557
rect 9137 1519 9209 1557
rect 9261 1519 9333 1557
rect 9385 1519 10097 1557
rect 10149 1519 10221 1557
rect 10273 1519 10345 1557
rect 10397 1519 10469 1557
rect 10521 1519 11131 1557
rect 1131 1498 11131 1519
rect 1131 1452 1144 1498
rect 11118 1452 11131 1498
rect 1131 1447 11131 1452
rect 1131 1395 1741 1447
rect 1793 1395 1865 1447
rect 1917 1395 1989 1447
rect 2041 1395 2113 1447
rect 2165 1395 2877 1447
rect 2929 1395 3001 1447
rect 3053 1395 3125 1447
rect 3177 1395 3249 1447
rect 3301 1395 4013 1447
rect 4065 1395 4137 1447
rect 4189 1395 4261 1447
rect 4313 1395 4385 1447
rect 4437 1395 5149 1447
rect 5201 1395 5273 1447
rect 5325 1395 5397 1447
rect 5449 1395 5521 1447
rect 5573 1395 6689 1447
rect 6741 1395 6813 1447
rect 6865 1395 6937 1447
rect 6989 1395 7061 1447
rect 7113 1395 7825 1447
rect 7877 1395 7949 1447
rect 8001 1395 8073 1447
rect 8125 1395 8197 1447
rect 8249 1395 8961 1447
rect 9013 1395 9085 1447
rect 9137 1395 9209 1447
rect 9261 1395 9333 1447
rect 9385 1395 10097 1447
rect 10149 1395 10221 1447
rect 10273 1395 10345 1447
rect 10397 1395 10469 1447
rect 10521 1395 11131 1447
rect 1131 1392 11131 1395
rect 1131 1346 1144 1392
rect 11118 1346 11131 1392
rect 1131 1323 11131 1346
rect 1131 1286 1741 1323
rect 1793 1286 1865 1323
rect 1917 1286 1989 1323
rect 2041 1286 2113 1323
rect 2165 1286 2877 1323
rect 2929 1286 3001 1323
rect 3053 1286 3125 1323
rect 3177 1286 3249 1323
rect 3301 1286 4013 1323
rect 4065 1286 4137 1323
rect 4189 1286 4261 1323
rect 4313 1286 4385 1323
rect 4437 1286 5149 1323
rect 5201 1286 5273 1323
rect 5325 1286 5397 1323
rect 5449 1286 5521 1323
rect 5573 1286 6689 1323
rect 6741 1286 6813 1323
rect 6865 1286 6937 1323
rect 6989 1286 7061 1323
rect 7113 1286 7825 1323
rect 7877 1286 7949 1323
rect 8001 1286 8073 1323
rect 8125 1286 8197 1323
rect 8249 1286 8961 1323
rect 9013 1286 9085 1323
rect 9137 1286 9209 1323
rect 9261 1286 9333 1323
rect 9385 1286 10097 1323
rect 10149 1286 10221 1323
rect 10273 1286 10345 1323
rect 10397 1286 10469 1323
rect 10521 1286 11131 1323
rect 1131 1240 1144 1286
rect 11118 1240 11131 1286
rect 1131 1199 11131 1240
rect 1131 1180 1741 1199
rect 1793 1180 1865 1199
rect 1917 1180 1989 1199
rect 2041 1180 2113 1199
rect 2165 1180 2877 1199
rect 2929 1180 3001 1199
rect 3053 1180 3125 1199
rect 3177 1180 3249 1199
rect 3301 1180 4013 1199
rect 4065 1180 4137 1199
rect 4189 1180 4261 1199
rect 4313 1180 4385 1199
rect 4437 1180 5149 1199
rect 5201 1180 5273 1199
rect 5325 1180 5397 1199
rect 5449 1180 5521 1199
rect 5573 1180 6689 1199
rect 6741 1180 6813 1199
rect 6865 1180 6937 1199
rect 6989 1180 7061 1199
rect 7113 1180 7825 1199
rect 7877 1180 7949 1199
rect 8001 1180 8073 1199
rect 8125 1180 8197 1199
rect 8249 1180 8961 1199
rect 9013 1180 9085 1199
rect 9137 1180 9209 1199
rect 9261 1180 9333 1199
rect 9385 1180 10097 1199
rect 10149 1180 10221 1199
rect 10273 1180 10345 1199
rect 10397 1180 10469 1199
rect 10521 1180 11131 1199
rect 1131 1134 1144 1180
rect 11118 1134 11131 1180
rect 1131 1121 11131 1134
rect 11345 907 11356 1935
rect 11402 1879 11510 1935
rect 11417 1827 11473 1879
rect 11402 1771 11510 1827
rect 11417 1719 11473 1771
rect 11402 1663 11510 1719
rect 11417 1611 11473 1663
rect 11402 1555 11510 1611
rect 11417 1503 11473 1555
rect 11402 1447 11510 1503
rect 11417 1395 11473 1447
rect 11402 1339 11510 1395
rect 11417 1287 11473 1339
rect 11402 1231 11510 1287
rect 11417 1179 11473 1231
rect 11402 1123 11510 1179
rect 11417 1071 11473 1123
rect 11402 1015 11510 1071
rect 11417 963 11473 1015
rect 11402 907 11510 963
rect 695 855 737 872
rect 789 855 845 907
rect 906 896 11356 907
rect 906 881 1032 896
rect 897 855 1032 881
rect 11230 881 11356 896
rect 695 850 1032 855
rect 11230 855 11365 881
rect 11417 855 11473 907
rect 11556 872 11567 6182
rect 11525 855 11567 872
rect 11230 850 11567 855
rect 695 824 2279 850
rect 2331 824 2387 850
rect 2439 824 2495 850
rect 2547 824 2603 850
rect 2655 824 2711 850
rect 2763 824 4551 850
rect 4603 824 4659 850
rect 4711 824 4767 850
rect 4819 824 4875 850
rect 4927 824 4983 850
rect 5035 824 7227 850
rect 7279 824 7335 850
rect 7387 824 7443 850
rect 7495 824 7551 850
rect 7603 824 7659 850
rect 7711 824 9499 850
rect 9551 824 9607 850
rect 9659 824 9715 850
rect 9767 824 9823 850
rect 9875 824 9931 850
rect 9983 824 11567 850
rect 695 799 11567 824
rect 695 747 737 799
rect 789 747 845 799
rect 897 768 11365 799
rect 897 747 2279 768
rect 695 742 2279 747
rect 2331 742 2387 768
rect 2439 742 2495 768
rect 2547 742 2603 768
rect 2655 742 2711 768
rect 2763 742 4551 768
rect 4603 742 4659 768
rect 4711 742 4767 768
rect 4819 742 4875 768
rect 4927 742 4983 768
rect 5035 742 7227 768
rect 7279 742 7335 768
rect 7387 742 7443 768
rect 7495 742 7551 768
rect 7603 742 7659 768
rect 7711 742 9499 768
rect 9551 742 9607 768
rect 9659 742 9715 768
rect 9767 742 9823 768
rect 9875 742 9931 768
rect 9983 747 11365 768
rect 11417 747 11473 799
rect 11525 747 11567 799
rect 9983 742 11567 747
rect 695 696 750 742
rect 11512 696 11567 742
rect 695 685 11567 696
rect 11751 511 11762 6543
rect 500 500 11762 511
rect 500 54 608 500
rect 11654 54 11762 500
rect 12208 54 12219 7000
rect 43 43 12219 54
<< via1 >>
rect 605 14344 608 14396
rect 608 14344 657 14396
rect 729 14344 781 14396
rect 853 14344 905 14396
rect 977 14344 1029 14396
rect 2309 14344 2361 14396
rect 2433 14344 2485 14396
rect 2557 14344 2609 14396
rect 2681 14344 2733 14396
rect 4581 14344 4633 14396
rect 4705 14344 4757 14396
rect 4829 14344 4881 14396
rect 4953 14344 5005 14396
rect 7257 14344 7309 14396
rect 7381 14344 7433 14396
rect 7505 14344 7557 14396
rect 7629 14344 7681 14396
rect 9529 14344 9581 14396
rect 9653 14344 9705 14396
rect 9777 14344 9829 14396
rect 9901 14344 9953 14396
rect 11233 14344 11285 14396
rect 11357 14344 11409 14396
rect 11481 14344 11533 14396
rect 11605 14344 11654 14396
rect 11654 14344 11657 14396
rect 605 14220 608 14272
rect 608 14220 657 14272
rect 729 14220 781 14272
rect 853 14220 905 14272
rect 977 14220 1029 14272
rect 2309 14220 2361 14272
rect 2433 14220 2485 14272
rect 2557 14220 2609 14272
rect 2681 14220 2733 14272
rect 4581 14220 4633 14272
rect 4705 14220 4757 14272
rect 4829 14220 4881 14272
rect 4953 14220 5005 14272
rect 7257 14220 7309 14272
rect 7381 14220 7433 14272
rect 7505 14220 7557 14272
rect 7629 14220 7681 14272
rect 9529 14220 9581 14272
rect 9653 14220 9705 14272
rect 9777 14220 9829 14272
rect 9901 14220 9953 14272
rect 11233 14220 11285 14272
rect 11357 14220 11409 14272
rect 11481 14220 11533 14272
rect 11605 14220 11654 14272
rect 11654 14220 11657 14272
rect 605 14096 608 14148
rect 608 14096 657 14148
rect 729 14096 781 14148
rect 853 14096 905 14148
rect 977 14096 1029 14148
rect 2309 14096 2361 14148
rect 2433 14096 2485 14148
rect 2557 14096 2609 14148
rect 2681 14096 2733 14148
rect 4581 14096 4633 14148
rect 4705 14096 4757 14148
rect 4829 14096 4881 14148
rect 4953 14096 5005 14148
rect 7257 14096 7309 14148
rect 7381 14096 7433 14148
rect 7505 14096 7557 14148
rect 7629 14096 7681 14148
rect 9529 14096 9581 14148
rect 9653 14096 9705 14148
rect 9777 14096 9829 14148
rect 9901 14096 9953 14148
rect 11233 14096 11285 14148
rect 11357 14096 11409 14148
rect 11481 14096 11533 14148
rect 11605 14096 11654 14148
rect 11654 14096 11657 14148
rect 605 13972 608 14024
rect 608 13972 657 14024
rect 729 13972 781 14024
rect 853 13972 905 14024
rect 977 13972 1029 14024
rect 2309 13972 2361 14024
rect 2433 13972 2485 14024
rect 2557 13972 2609 14024
rect 2681 13972 2733 14024
rect 4581 13972 4633 14024
rect 4705 13972 4757 14024
rect 4829 13972 4881 14024
rect 4953 13972 5005 14024
rect 7257 13972 7309 14024
rect 7381 13972 7433 14024
rect 7505 13972 7557 14024
rect 7629 13972 7681 14024
rect 9529 13972 9581 14024
rect 9653 13972 9705 14024
rect 9777 13972 9829 14024
rect 9901 13972 9953 14024
rect 11233 13972 11285 14024
rect 11357 13972 11409 14024
rect 11481 13972 11533 14024
rect 11605 13972 11654 14024
rect 11654 13972 11657 14024
rect 1143 13719 1195 13745
rect 1251 13719 1303 13745
rect 1359 13719 1411 13745
rect 1467 13719 1519 13745
rect 1575 13719 1627 13745
rect 3415 13719 3467 13745
rect 3523 13719 3575 13745
rect 3631 13719 3683 13745
rect 3739 13719 3791 13745
rect 3847 13719 3899 13745
rect 5700 13719 5752 13745
rect 5808 13719 5860 13745
rect 5916 13719 5968 13745
rect 6024 13719 6076 13745
rect 6186 13719 6238 13745
rect 6294 13719 6346 13745
rect 6402 13719 6454 13745
rect 6510 13719 6562 13745
rect 8363 13719 8415 13745
rect 8471 13719 8523 13745
rect 8579 13719 8631 13745
rect 8687 13719 8739 13745
rect 8795 13719 8847 13745
rect 10635 13719 10687 13745
rect 10743 13719 10795 13745
rect 10851 13719 10903 13745
rect 10959 13719 11011 13745
rect 11067 13719 11119 13745
rect 1143 13693 1195 13719
rect 1251 13693 1303 13719
rect 1359 13693 1411 13719
rect 1467 13693 1519 13719
rect 1575 13693 1627 13719
rect 3415 13693 3467 13719
rect 3523 13693 3575 13719
rect 3631 13693 3683 13719
rect 3739 13693 3791 13719
rect 3847 13693 3899 13719
rect 5700 13693 5752 13719
rect 5808 13693 5860 13719
rect 5916 13693 5968 13719
rect 6024 13693 6076 13719
rect 6186 13693 6238 13719
rect 6294 13693 6346 13719
rect 6402 13693 6454 13719
rect 6510 13693 6562 13719
rect 8363 13693 8415 13719
rect 8471 13693 8523 13719
rect 8579 13693 8631 13719
rect 8687 13693 8739 13719
rect 8795 13693 8847 13719
rect 10635 13693 10687 13719
rect 10743 13693 10795 13719
rect 10851 13693 10903 13719
rect 10959 13693 11011 13719
rect 11067 13693 11119 13719
rect 1143 13611 1195 13637
rect 1251 13611 1303 13637
rect 1359 13611 1411 13637
rect 1467 13611 1519 13637
rect 1575 13611 1627 13637
rect 3415 13611 3467 13637
rect 3523 13611 3575 13637
rect 3631 13611 3683 13637
rect 3739 13611 3791 13637
rect 3847 13611 3899 13637
rect 5700 13611 5752 13637
rect 5808 13611 5860 13637
rect 5916 13611 5968 13637
rect 6024 13611 6076 13637
rect 6186 13611 6238 13637
rect 6294 13611 6346 13637
rect 6402 13611 6454 13637
rect 6510 13611 6562 13637
rect 8363 13611 8415 13637
rect 8471 13611 8523 13637
rect 8579 13611 8631 13637
rect 8687 13611 8739 13637
rect 8795 13611 8847 13637
rect 10635 13611 10687 13637
rect 10743 13611 10795 13637
rect 10851 13611 10903 13637
rect 10959 13611 11011 13637
rect 11067 13611 11119 13637
rect 1143 13585 1195 13611
rect 1251 13585 1303 13611
rect 1359 13585 1411 13611
rect 1467 13585 1519 13611
rect 1575 13585 1627 13611
rect 3415 13585 3467 13611
rect 3523 13585 3575 13611
rect 3631 13585 3683 13611
rect 3739 13585 3791 13611
rect 3847 13585 3899 13611
rect 5700 13585 5752 13611
rect 5808 13585 5860 13611
rect 5916 13585 5968 13611
rect 6024 13585 6076 13611
rect 6186 13585 6238 13611
rect 6294 13585 6346 13611
rect 6402 13585 6454 13611
rect 6510 13585 6562 13611
rect 8363 13585 8415 13611
rect 8471 13585 8523 13611
rect 8579 13585 8631 13611
rect 8687 13585 8739 13611
rect 8795 13585 8847 13611
rect 10635 13585 10687 13611
rect 10743 13585 10795 13611
rect 10851 13585 10903 13611
rect 10959 13585 11011 13611
rect 11067 13585 11119 13611
rect 1741 13281 1793 13314
rect 1865 13281 1917 13314
rect 1989 13281 2041 13314
rect 2113 13281 2165 13314
rect 2877 13281 2929 13314
rect 3001 13281 3053 13314
rect 3125 13281 3177 13314
rect 3249 13281 3301 13314
rect 4013 13281 4065 13314
rect 4137 13281 4189 13314
rect 4261 13281 4313 13314
rect 4385 13281 4437 13314
rect 5149 13281 5201 13314
rect 5273 13281 5325 13314
rect 5397 13281 5449 13314
rect 5521 13281 5573 13314
rect 6689 13281 6741 13314
rect 6813 13281 6865 13314
rect 6937 13281 6989 13314
rect 7061 13281 7113 13314
rect 7825 13281 7877 13314
rect 7949 13281 8001 13314
rect 8073 13281 8125 13314
rect 8197 13281 8249 13314
rect 8961 13281 9013 13314
rect 9085 13281 9137 13314
rect 9209 13281 9261 13314
rect 9333 13281 9385 13314
rect 10097 13281 10149 13314
rect 10221 13281 10273 13314
rect 10345 13281 10397 13314
rect 10469 13281 10521 13314
rect 1741 13262 1793 13281
rect 1865 13262 1917 13281
rect 1989 13262 2041 13281
rect 2113 13262 2165 13281
rect 2877 13262 2929 13281
rect 3001 13262 3053 13281
rect 3125 13262 3177 13281
rect 3249 13262 3301 13281
rect 4013 13262 4065 13281
rect 4137 13262 4189 13281
rect 4261 13262 4313 13281
rect 4385 13262 4437 13281
rect 5149 13262 5201 13281
rect 5273 13262 5325 13281
rect 5397 13262 5449 13281
rect 5521 13262 5573 13281
rect 6689 13262 6741 13281
rect 6813 13262 6865 13281
rect 6937 13262 6989 13281
rect 7061 13262 7113 13281
rect 7825 13262 7877 13281
rect 7949 13262 8001 13281
rect 8073 13262 8125 13281
rect 8197 13262 8249 13281
rect 8961 13262 9013 13281
rect 9085 13262 9137 13281
rect 9209 13262 9261 13281
rect 9333 13262 9385 13281
rect 10097 13262 10149 13281
rect 10221 13262 10273 13281
rect 10345 13262 10397 13281
rect 10469 13262 10521 13281
rect 1741 13176 1793 13190
rect 1865 13176 1917 13190
rect 1989 13176 2041 13190
rect 2113 13176 2165 13190
rect 2877 13176 2929 13190
rect 3001 13176 3053 13190
rect 3125 13176 3177 13190
rect 3249 13176 3301 13190
rect 4013 13176 4065 13190
rect 4137 13176 4189 13190
rect 4261 13176 4313 13190
rect 4385 13176 4437 13190
rect 5149 13176 5201 13190
rect 5273 13176 5325 13190
rect 5397 13176 5449 13190
rect 5521 13176 5573 13190
rect 6689 13176 6741 13190
rect 6813 13176 6865 13190
rect 6937 13176 6989 13190
rect 7061 13176 7113 13190
rect 7825 13176 7877 13190
rect 7949 13176 8001 13190
rect 8073 13176 8125 13190
rect 8197 13176 8249 13190
rect 8961 13176 9013 13190
rect 9085 13176 9137 13190
rect 9209 13176 9261 13190
rect 9333 13176 9385 13190
rect 10097 13176 10149 13190
rect 10221 13176 10273 13190
rect 10345 13176 10397 13190
rect 10469 13176 10521 13190
rect 1741 13138 1793 13176
rect 1865 13138 1917 13176
rect 1989 13138 2041 13176
rect 2113 13138 2165 13176
rect 2877 13138 2929 13176
rect 3001 13138 3053 13176
rect 3125 13138 3177 13176
rect 3249 13138 3301 13176
rect 4013 13138 4065 13176
rect 4137 13138 4189 13176
rect 4261 13138 4313 13176
rect 4385 13138 4437 13176
rect 5149 13138 5201 13176
rect 5273 13138 5325 13176
rect 5397 13138 5449 13176
rect 5521 13138 5573 13176
rect 6689 13138 6741 13176
rect 6813 13138 6865 13176
rect 6937 13138 6989 13176
rect 7061 13138 7113 13176
rect 7825 13138 7877 13176
rect 7949 13138 8001 13176
rect 8073 13138 8125 13176
rect 8197 13138 8249 13176
rect 8961 13138 9013 13176
rect 9085 13138 9137 13176
rect 9209 13138 9261 13176
rect 9333 13138 9385 13176
rect 10097 13138 10149 13176
rect 10221 13138 10273 13176
rect 10345 13138 10397 13176
rect 10469 13138 10521 13176
rect 1741 13014 1793 13066
rect 1865 13014 1917 13066
rect 1989 13014 2041 13066
rect 2113 13014 2165 13066
rect 2877 13014 2929 13066
rect 3001 13014 3053 13066
rect 3125 13014 3177 13066
rect 3249 13014 3301 13066
rect 4013 13014 4065 13066
rect 4137 13014 4189 13066
rect 4261 13014 4313 13066
rect 4385 13014 4437 13066
rect 5149 13014 5201 13066
rect 5273 13014 5325 13066
rect 5397 13014 5449 13066
rect 5521 13014 5573 13066
rect 6689 13014 6741 13066
rect 6813 13014 6865 13066
rect 6937 13014 6989 13066
rect 7061 13014 7113 13066
rect 7825 13014 7877 13066
rect 7949 13014 8001 13066
rect 8073 13014 8125 13066
rect 8197 13014 8249 13066
rect 8961 13014 9013 13066
rect 9085 13014 9137 13066
rect 9209 13014 9261 13066
rect 9333 13014 9385 13066
rect 10097 13014 10149 13066
rect 10221 13014 10273 13066
rect 10345 13014 10397 13066
rect 10469 13014 10521 13066
rect 1741 12905 1793 12942
rect 1865 12905 1917 12942
rect 1989 12905 2041 12942
rect 2113 12905 2165 12942
rect 2877 12905 2929 12942
rect 3001 12905 3053 12942
rect 3125 12905 3177 12942
rect 3249 12905 3301 12942
rect 4013 12905 4065 12942
rect 4137 12905 4189 12942
rect 4261 12905 4313 12942
rect 4385 12905 4437 12942
rect 5149 12905 5201 12942
rect 5273 12905 5325 12942
rect 5397 12905 5449 12942
rect 5521 12905 5573 12942
rect 6689 12905 6741 12942
rect 6813 12905 6865 12942
rect 6937 12905 6989 12942
rect 7061 12905 7113 12942
rect 7825 12905 7877 12942
rect 7949 12905 8001 12942
rect 8073 12905 8125 12942
rect 8197 12905 8249 12942
rect 8961 12905 9013 12942
rect 9085 12905 9137 12942
rect 9209 12905 9261 12942
rect 9333 12905 9385 12942
rect 10097 12905 10149 12942
rect 10221 12905 10273 12942
rect 10345 12905 10397 12942
rect 10469 12905 10521 12942
rect 1741 12890 1793 12905
rect 1865 12890 1917 12905
rect 1989 12890 2041 12905
rect 2113 12890 2165 12905
rect 2877 12890 2929 12905
rect 3001 12890 3053 12905
rect 3125 12890 3177 12905
rect 3249 12890 3301 12905
rect 4013 12890 4065 12905
rect 4137 12890 4189 12905
rect 4261 12890 4313 12905
rect 4385 12890 4437 12905
rect 5149 12890 5201 12905
rect 5273 12890 5325 12905
rect 5397 12890 5449 12905
rect 5521 12890 5573 12905
rect 6689 12890 6741 12905
rect 6813 12890 6865 12905
rect 6937 12890 6989 12905
rect 7061 12890 7113 12905
rect 7825 12890 7877 12905
rect 7949 12890 8001 12905
rect 8073 12890 8125 12905
rect 8197 12890 8249 12905
rect 8961 12890 9013 12905
rect 9085 12890 9137 12905
rect 9209 12890 9261 12905
rect 9333 12890 9385 12905
rect 10097 12890 10149 12905
rect 10221 12890 10273 12905
rect 10345 12890 10397 12905
rect 10469 12890 10521 12905
rect 1741 12799 1793 12818
rect 1865 12799 1917 12818
rect 1989 12799 2041 12818
rect 2113 12799 2165 12818
rect 2877 12799 2929 12818
rect 3001 12799 3053 12818
rect 3125 12799 3177 12818
rect 3249 12799 3301 12818
rect 4013 12799 4065 12818
rect 4137 12799 4189 12818
rect 4261 12799 4313 12818
rect 4385 12799 4437 12818
rect 5149 12799 5201 12818
rect 5273 12799 5325 12818
rect 5397 12799 5449 12818
rect 5521 12799 5573 12818
rect 6689 12799 6741 12818
rect 6813 12799 6865 12818
rect 6937 12799 6989 12818
rect 7061 12799 7113 12818
rect 7825 12799 7877 12818
rect 7949 12799 8001 12818
rect 8073 12799 8125 12818
rect 8197 12799 8249 12818
rect 8961 12799 9013 12818
rect 9085 12799 9137 12818
rect 9209 12799 9261 12818
rect 9333 12799 9385 12818
rect 10097 12799 10149 12818
rect 10221 12799 10273 12818
rect 10345 12799 10397 12818
rect 10469 12799 10521 12818
rect 1741 12766 1793 12799
rect 1865 12766 1917 12799
rect 1989 12766 2041 12799
rect 2113 12766 2165 12799
rect 2877 12766 2929 12799
rect 3001 12766 3053 12799
rect 3125 12766 3177 12799
rect 3249 12766 3301 12799
rect 4013 12766 4065 12799
rect 4137 12766 4189 12799
rect 4261 12766 4313 12799
rect 4385 12766 4437 12799
rect 5149 12766 5201 12799
rect 5273 12766 5325 12799
rect 5397 12766 5449 12799
rect 5521 12766 5573 12799
rect 6689 12766 6741 12799
rect 6813 12766 6865 12799
rect 6937 12766 6989 12799
rect 7061 12766 7113 12799
rect 7825 12766 7877 12799
rect 7949 12766 8001 12799
rect 8073 12766 8125 12799
rect 8197 12766 8249 12799
rect 8961 12766 9013 12799
rect 9085 12766 9137 12799
rect 9209 12766 9261 12799
rect 9333 12766 9385 12799
rect 10097 12766 10149 12799
rect 10221 12766 10273 12799
rect 10345 12766 10397 12799
rect 10469 12766 10521 12799
rect 1143 12469 1195 12472
rect 1251 12469 1303 12472
rect 1359 12469 1411 12472
rect 1467 12469 1519 12472
rect 1575 12469 1627 12472
rect 3415 12469 3467 12472
rect 3523 12469 3575 12472
rect 3631 12469 3683 12472
rect 3739 12469 3791 12472
rect 3847 12469 3899 12472
rect 5700 12469 5752 12472
rect 5808 12469 5860 12472
rect 5916 12469 5968 12472
rect 6024 12469 6076 12472
rect 6186 12469 6238 12472
rect 6294 12469 6346 12472
rect 6402 12469 6454 12472
rect 6510 12469 6562 12472
rect 8363 12469 8415 12472
rect 8471 12469 8523 12472
rect 8579 12469 8631 12472
rect 8687 12469 8739 12472
rect 8795 12469 8847 12472
rect 10635 12469 10687 12472
rect 10743 12469 10795 12472
rect 10851 12469 10903 12472
rect 10959 12469 11011 12472
rect 11067 12469 11119 12472
rect 1143 12420 1195 12469
rect 1251 12420 1303 12469
rect 1359 12420 1411 12469
rect 1467 12420 1519 12469
rect 1575 12420 1627 12469
rect 3415 12420 3467 12469
rect 3523 12420 3575 12469
rect 3631 12420 3683 12469
rect 3739 12420 3791 12469
rect 3847 12420 3899 12469
rect 5700 12420 5752 12469
rect 5808 12420 5860 12469
rect 5916 12420 5968 12469
rect 6024 12420 6076 12469
rect 6186 12420 6238 12469
rect 6294 12420 6346 12469
rect 6402 12420 6454 12469
rect 6510 12420 6562 12469
rect 8363 12420 8415 12469
rect 8471 12420 8523 12469
rect 8579 12420 8631 12469
rect 8687 12420 8739 12469
rect 8795 12420 8847 12469
rect 10635 12420 10687 12469
rect 10743 12420 10795 12469
rect 10851 12420 10903 12469
rect 10959 12420 11011 12469
rect 11067 12420 11119 12469
rect 1143 12361 1195 12364
rect 1251 12361 1303 12364
rect 1359 12361 1411 12364
rect 1467 12361 1519 12364
rect 1575 12361 1627 12364
rect 3415 12361 3467 12364
rect 3523 12361 3575 12364
rect 3631 12361 3683 12364
rect 3739 12361 3791 12364
rect 3847 12361 3899 12364
rect 5700 12361 5752 12364
rect 5808 12361 5860 12364
rect 5916 12361 5968 12364
rect 6024 12361 6076 12364
rect 6186 12361 6238 12364
rect 6294 12361 6346 12364
rect 6402 12361 6454 12364
rect 6510 12361 6562 12364
rect 8363 12361 8415 12364
rect 8471 12361 8523 12364
rect 8579 12361 8631 12364
rect 8687 12361 8739 12364
rect 8795 12361 8847 12364
rect 10635 12361 10687 12364
rect 10743 12361 10795 12364
rect 10851 12361 10903 12364
rect 10959 12361 11011 12364
rect 11067 12361 11119 12364
rect 1143 12315 1195 12361
rect 1251 12315 1303 12361
rect 1359 12315 1411 12361
rect 1467 12315 1519 12361
rect 1575 12315 1627 12361
rect 3415 12315 3467 12361
rect 3523 12315 3575 12361
rect 3631 12315 3683 12361
rect 3739 12315 3791 12361
rect 3847 12315 3899 12361
rect 5700 12315 5752 12361
rect 5808 12315 5860 12361
rect 5916 12315 5968 12361
rect 6024 12315 6076 12361
rect 6186 12315 6238 12361
rect 6294 12315 6346 12361
rect 6402 12315 6454 12361
rect 6510 12315 6562 12361
rect 8363 12315 8415 12361
rect 8471 12315 8523 12361
rect 8579 12315 8631 12361
rect 8687 12315 8739 12361
rect 8795 12315 8847 12361
rect 10635 12315 10687 12361
rect 10743 12315 10795 12361
rect 10851 12315 10903 12361
rect 10959 12315 11011 12361
rect 11067 12315 11119 12361
rect 1143 12312 1195 12315
rect 1251 12312 1303 12315
rect 1359 12312 1411 12315
rect 1467 12312 1519 12315
rect 1575 12312 1627 12315
rect 3415 12312 3467 12315
rect 3523 12312 3575 12315
rect 3631 12312 3683 12315
rect 3739 12312 3791 12315
rect 3847 12312 3899 12315
rect 5700 12312 5752 12315
rect 5808 12312 5860 12315
rect 5916 12312 5968 12315
rect 6024 12312 6076 12315
rect 6186 12312 6238 12315
rect 6294 12312 6346 12315
rect 6402 12312 6454 12315
rect 6510 12312 6562 12315
rect 8363 12312 8415 12315
rect 8471 12312 8523 12315
rect 8579 12312 8631 12315
rect 8687 12312 8739 12315
rect 8795 12312 8847 12315
rect 10635 12312 10687 12315
rect 10743 12312 10795 12315
rect 10851 12312 10903 12315
rect 10959 12312 11011 12315
rect 11067 12312 11119 12315
rect 1143 12207 1195 12256
rect 1251 12207 1303 12256
rect 1359 12207 1411 12256
rect 1467 12207 1519 12256
rect 1575 12207 1627 12256
rect 3415 12207 3467 12256
rect 3523 12207 3575 12256
rect 3631 12207 3683 12256
rect 3739 12207 3791 12256
rect 3847 12207 3899 12256
rect 5700 12207 5752 12256
rect 5808 12207 5860 12256
rect 5916 12207 5968 12256
rect 6024 12207 6076 12256
rect 6186 12207 6238 12256
rect 6294 12207 6346 12256
rect 6402 12207 6454 12256
rect 6510 12207 6562 12256
rect 8363 12207 8415 12256
rect 8471 12207 8523 12256
rect 8579 12207 8631 12256
rect 8687 12207 8739 12256
rect 8795 12207 8847 12256
rect 10635 12207 10687 12256
rect 10743 12207 10795 12256
rect 10851 12207 10903 12256
rect 10959 12207 11011 12256
rect 11067 12207 11119 12256
rect 1143 12204 1195 12207
rect 1251 12204 1303 12207
rect 1359 12204 1411 12207
rect 1467 12204 1519 12207
rect 1575 12204 1627 12207
rect 3415 12204 3467 12207
rect 3523 12204 3575 12207
rect 3631 12204 3683 12207
rect 3739 12204 3791 12207
rect 3847 12204 3899 12207
rect 5700 12204 5752 12207
rect 5808 12204 5860 12207
rect 5916 12204 5968 12207
rect 6024 12204 6076 12207
rect 6186 12204 6238 12207
rect 6294 12204 6346 12207
rect 6402 12204 6454 12207
rect 6510 12204 6562 12207
rect 8363 12204 8415 12207
rect 8471 12204 8523 12207
rect 8579 12204 8631 12207
rect 8687 12204 8739 12207
rect 8795 12204 8847 12207
rect 10635 12204 10687 12207
rect 10743 12204 10795 12207
rect 10851 12204 10903 12207
rect 10959 12204 11011 12207
rect 11067 12204 11119 12207
rect 1741 11877 1793 11910
rect 1865 11877 1917 11910
rect 1989 11877 2041 11910
rect 2113 11877 2165 11910
rect 2877 11877 2929 11910
rect 3001 11877 3053 11910
rect 3125 11877 3177 11910
rect 3249 11877 3301 11910
rect 4013 11877 4065 11910
rect 4137 11877 4189 11910
rect 4261 11877 4313 11910
rect 4385 11877 4437 11910
rect 5149 11877 5201 11910
rect 5273 11877 5325 11910
rect 5397 11877 5449 11910
rect 5521 11877 5573 11910
rect 6689 11877 6741 11910
rect 6813 11877 6865 11910
rect 6937 11877 6989 11910
rect 7061 11877 7113 11910
rect 7825 11877 7877 11910
rect 7949 11877 8001 11910
rect 8073 11877 8125 11910
rect 8197 11877 8249 11910
rect 8961 11877 9013 11910
rect 9085 11877 9137 11910
rect 9209 11877 9261 11910
rect 9333 11877 9385 11910
rect 10097 11877 10149 11910
rect 10221 11877 10273 11910
rect 10345 11877 10397 11910
rect 10469 11877 10521 11910
rect 1741 11858 1793 11877
rect 1865 11858 1917 11877
rect 1989 11858 2041 11877
rect 2113 11858 2165 11877
rect 2877 11858 2929 11877
rect 3001 11858 3053 11877
rect 3125 11858 3177 11877
rect 3249 11858 3301 11877
rect 4013 11858 4065 11877
rect 4137 11858 4189 11877
rect 4261 11858 4313 11877
rect 4385 11858 4437 11877
rect 5149 11858 5201 11877
rect 5273 11858 5325 11877
rect 5397 11858 5449 11877
rect 5521 11858 5573 11877
rect 6689 11858 6741 11877
rect 6813 11858 6865 11877
rect 6937 11858 6989 11877
rect 7061 11858 7113 11877
rect 7825 11858 7877 11877
rect 7949 11858 8001 11877
rect 8073 11858 8125 11877
rect 8197 11858 8249 11877
rect 8961 11858 9013 11877
rect 9085 11858 9137 11877
rect 9209 11858 9261 11877
rect 9333 11858 9385 11877
rect 10097 11858 10149 11877
rect 10221 11858 10273 11877
rect 10345 11858 10397 11877
rect 10469 11858 10521 11877
rect 1741 11772 1793 11786
rect 1865 11772 1917 11786
rect 1989 11772 2041 11786
rect 2113 11772 2165 11786
rect 2877 11772 2929 11786
rect 3001 11772 3053 11786
rect 3125 11772 3177 11786
rect 3249 11772 3301 11786
rect 4013 11772 4065 11786
rect 4137 11772 4189 11786
rect 4261 11772 4313 11786
rect 4385 11772 4437 11786
rect 5149 11772 5201 11786
rect 5273 11772 5325 11786
rect 5397 11772 5449 11786
rect 5521 11772 5573 11786
rect 6689 11772 6741 11786
rect 6813 11772 6865 11786
rect 6937 11772 6989 11786
rect 7061 11772 7113 11786
rect 7825 11772 7877 11786
rect 7949 11772 8001 11786
rect 8073 11772 8125 11786
rect 8197 11772 8249 11786
rect 8961 11772 9013 11786
rect 9085 11772 9137 11786
rect 9209 11772 9261 11786
rect 9333 11772 9385 11786
rect 10097 11772 10149 11786
rect 10221 11772 10273 11786
rect 10345 11772 10397 11786
rect 10469 11772 10521 11786
rect 1741 11734 1793 11772
rect 1865 11734 1917 11772
rect 1989 11734 2041 11772
rect 2113 11734 2165 11772
rect 2877 11734 2929 11772
rect 3001 11734 3053 11772
rect 3125 11734 3177 11772
rect 3249 11734 3301 11772
rect 4013 11734 4065 11772
rect 4137 11734 4189 11772
rect 4261 11734 4313 11772
rect 4385 11734 4437 11772
rect 5149 11734 5201 11772
rect 5273 11734 5325 11772
rect 5397 11734 5449 11772
rect 5521 11734 5573 11772
rect 6689 11734 6741 11772
rect 6813 11734 6865 11772
rect 6937 11734 6989 11772
rect 7061 11734 7113 11772
rect 7825 11734 7877 11772
rect 7949 11734 8001 11772
rect 8073 11734 8125 11772
rect 8197 11734 8249 11772
rect 8961 11734 9013 11772
rect 9085 11734 9137 11772
rect 9209 11734 9261 11772
rect 9333 11734 9385 11772
rect 10097 11734 10149 11772
rect 10221 11734 10273 11772
rect 10345 11734 10397 11772
rect 10469 11734 10521 11772
rect 1741 11610 1793 11662
rect 1865 11610 1917 11662
rect 1989 11610 2041 11662
rect 2113 11610 2165 11662
rect 2877 11610 2929 11662
rect 3001 11610 3053 11662
rect 3125 11610 3177 11662
rect 3249 11610 3301 11662
rect 4013 11610 4065 11662
rect 4137 11610 4189 11662
rect 4261 11610 4313 11662
rect 4385 11610 4437 11662
rect 5149 11610 5201 11662
rect 5273 11610 5325 11662
rect 5397 11610 5449 11662
rect 5521 11610 5573 11662
rect 6689 11610 6741 11662
rect 6813 11610 6865 11662
rect 6937 11610 6989 11662
rect 7061 11610 7113 11662
rect 7825 11610 7877 11662
rect 7949 11610 8001 11662
rect 8073 11610 8125 11662
rect 8197 11610 8249 11662
rect 8961 11610 9013 11662
rect 9085 11610 9137 11662
rect 9209 11610 9261 11662
rect 9333 11610 9385 11662
rect 10097 11610 10149 11662
rect 10221 11610 10273 11662
rect 10345 11610 10397 11662
rect 10469 11610 10521 11662
rect 1741 11501 1793 11538
rect 1865 11501 1917 11538
rect 1989 11501 2041 11538
rect 2113 11501 2165 11538
rect 2877 11501 2929 11538
rect 3001 11501 3053 11538
rect 3125 11501 3177 11538
rect 3249 11501 3301 11538
rect 4013 11501 4065 11538
rect 4137 11501 4189 11538
rect 4261 11501 4313 11538
rect 4385 11501 4437 11538
rect 5149 11501 5201 11538
rect 5273 11501 5325 11538
rect 5397 11501 5449 11538
rect 5521 11501 5573 11538
rect 6689 11501 6741 11538
rect 6813 11501 6865 11538
rect 6937 11501 6989 11538
rect 7061 11501 7113 11538
rect 7825 11501 7877 11538
rect 7949 11501 8001 11538
rect 8073 11501 8125 11538
rect 8197 11501 8249 11538
rect 8961 11501 9013 11538
rect 9085 11501 9137 11538
rect 9209 11501 9261 11538
rect 9333 11501 9385 11538
rect 10097 11501 10149 11538
rect 10221 11501 10273 11538
rect 10345 11501 10397 11538
rect 10469 11501 10521 11538
rect 1741 11486 1793 11501
rect 1865 11486 1917 11501
rect 1989 11486 2041 11501
rect 2113 11486 2165 11501
rect 2877 11486 2929 11501
rect 3001 11486 3053 11501
rect 3125 11486 3177 11501
rect 3249 11486 3301 11501
rect 4013 11486 4065 11501
rect 4137 11486 4189 11501
rect 4261 11486 4313 11501
rect 4385 11486 4437 11501
rect 5149 11486 5201 11501
rect 5273 11486 5325 11501
rect 5397 11486 5449 11501
rect 5521 11486 5573 11501
rect 6689 11486 6741 11501
rect 6813 11486 6865 11501
rect 6937 11486 6989 11501
rect 7061 11486 7113 11501
rect 7825 11486 7877 11501
rect 7949 11486 8001 11501
rect 8073 11486 8125 11501
rect 8197 11486 8249 11501
rect 8961 11486 9013 11501
rect 9085 11486 9137 11501
rect 9209 11486 9261 11501
rect 9333 11486 9385 11501
rect 10097 11486 10149 11501
rect 10221 11486 10273 11501
rect 10345 11486 10397 11501
rect 10469 11486 10521 11501
rect 1741 11395 1793 11414
rect 1865 11395 1917 11414
rect 1989 11395 2041 11414
rect 2113 11395 2165 11414
rect 2877 11395 2929 11414
rect 3001 11395 3053 11414
rect 3125 11395 3177 11414
rect 3249 11395 3301 11414
rect 4013 11395 4065 11414
rect 4137 11395 4189 11414
rect 4261 11395 4313 11414
rect 4385 11395 4437 11414
rect 5149 11395 5201 11414
rect 5273 11395 5325 11414
rect 5397 11395 5449 11414
rect 5521 11395 5573 11414
rect 6689 11395 6741 11414
rect 6813 11395 6865 11414
rect 6937 11395 6989 11414
rect 7061 11395 7113 11414
rect 7825 11395 7877 11414
rect 7949 11395 8001 11414
rect 8073 11395 8125 11414
rect 8197 11395 8249 11414
rect 8961 11395 9013 11414
rect 9085 11395 9137 11414
rect 9209 11395 9261 11414
rect 9333 11395 9385 11414
rect 10097 11395 10149 11414
rect 10221 11395 10273 11414
rect 10345 11395 10397 11414
rect 10469 11395 10521 11414
rect 1741 11362 1793 11395
rect 1865 11362 1917 11395
rect 1989 11362 2041 11395
rect 2113 11362 2165 11395
rect 2877 11362 2929 11395
rect 3001 11362 3053 11395
rect 3125 11362 3177 11395
rect 3249 11362 3301 11395
rect 4013 11362 4065 11395
rect 4137 11362 4189 11395
rect 4261 11362 4313 11395
rect 4385 11362 4437 11395
rect 5149 11362 5201 11395
rect 5273 11362 5325 11395
rect 5397 11362 5449 11395
rect 5521 11362 5573 11395
rect 6689 11362 6741 11395
rect 6813 11362 6865 11395
rect 6937 11362 6989 11395
rect 7061 11362 7113 11395
rect 7825 11362 7877 11395
rect 7949 11362 8001 11395
rect 8073 11362 8125 11395
rect 8197 11362 8249 11395
rect 8961 11362 9013 11395
rect 9085 11362 9137 11395
rect 9209 11362 9261 11395
rect 9333 11362 9385 11395
rect 10097 11362 10149 11395
rect 10221 11362 10273 11395
rect 10345 11362 10397 11395
rect 10469 11362 10521 11395
rect 1143 11065 1195 11068
rect 1251 11065 1303 11068
rect 1359 11065 1411 11068
rect 1467 11065 1519 11068
rect 1575 11065 1627 11068
rect 3415 11065 3467 11068
rect 3523 11065 3575 11068
rect 3631 11065 3683 11068
rect 3739 11065 3791 11068
rect 3847 11065 3899 11068
rect 5700 11065 5752 11068
rect 5808 11065 5860 11068
rect 5916 11065 5968 11068
rect 6024 11065 6076 11068
rect 6186 11065 6238 11068
rect 6294 11065 6346 11068
rect 6402 11065 6454 11068
rect 6510 11065 6562 11068
rect 8363 11065 8415 11068
rect 8471 11065 8523 11068
rect 8579 11065 8631 11068
rect 8687 11065 8739 11068
rect 8795 11065 8847 11068
rect 10635 11065 10687 11068
rect 10743 11065 10795 11068
rect 10851 11065 10903 11068
rect 10959 11065 11011 11068
rect 11067 11065 11119 11068
rect 1143 11016 1195 11065
rect 1251 11016 1303 11065
rect 1359 11016 1411 11065
rect 1467 11016 1519 11065
rect 1575 11016 1627 11065
rect 3415 11016 3467 11065
rect 3523 11016 3575 11065
rect 3631 11016 3683 11065
rect 3739 11016 3791 11065
rect 3847 11016 3899 11065
rect 5700 11016 5752 11065
rect 5808 11016 5860 11065
rect 5916 11016 5968 11065
rect 6024 11016 6076 11065
rect 6186 11016 6238 11065
rect 6294 11016 6346 11065
rect 6402 11016 6454 11065
rect 6510 11016 6562 11065
rect 8363 11016 8415 11065
rect 8471 11016 8523 11065
rect 8579 11016 8631 11065
rect 8687 11016 8739 11065
rect 8795 11016 8847 11065
rect 10635 11016 10687 11065
rect 10743 11016 10795 11065
rect 10851 11016 10903 11065
rect 10959 11016 11011 11065
rect 11067 11016 11119 11065
rect 1143 10957 1195 10960
rect 1251 10957 1303 10960
rect 1359 10957 1411 10960
rect 1467 10957 1519 10960
rect 1575 10957 1627 10960
rect 3415 10957 3467 10960
rect 3523 10957 3575 10960
rect 3631 10957 3683 10960
rect 3739 10957 3791 10960
rect 3847 10957 3899 10960
rect 5700 10957 5752 10960
rect 5808 10957 5860 10960
rect 5916 10957 5968 10960
rect 6024 10957 6076 10960
rect 6186 10957 6238 10960
rect 6294 10957 6346 10960
rect 6402 10957 6454 10960
rect 6510 10957 6562 10960
rect 8363 10957 8415 10960
rect 8471 10957 8523 10960
rect 8579 10957 8631 10960
rect 8687 10957 8739 10960
rect 8795 10957 8847 10960
rect 10635 10957 10687 10960
rect 10743 10957 10795 10960
rect 10851 10957 10903 10960
rect 10959 10957 11011 10960
rect 11067 10957 11119 10960
rect 1143 10911 1195 10957
rect 1251 10911 1303 10957
rect 1359 10911 1411 10957
rect 1467 10911 1519 10957
rect 1575 10911 1627 10957
rect 3415 10911 3467 10957
rect 3523 10911 3575 10957
rect 3631 10911 3683 10957
rect 3739 10911 3791 10957
rect 3847 10911 3899 10957
rect 5700 10911 5752 10957
rect 5808 10911 5860 10957
rect 5916 10911 5968 10957
rect 6024 10911 6076 10957
rect 6186 10911 6238 10957
rect 6294 10911 6346 10957
rect 6402 10911 6454 10957
rect 6510 10911 6562 10957
rect 8363 10911 8415 10957
rect 8471 10911 8523 10957
rect 8579 10911 8631 10957
rect 8687 10911 8739 10957
rect 8795 10911 8847 10957
rect 10635 10911 10687 10957
rect 10743 10911 10795 10957
rect 10851 10911 10903 10957
rect 10959 10911 11011 10957
rect 11067 10911 11119 10957
rect 1143 10908 1195 10911
rect 1251 10908 1303 10911
rect 1359 10908 1411 10911
rect 1467 10908 1519 10911
rect 1575 10908 1627 10911
rect 3415 10908 3467 10911
rect 3523 10908 3575 10911
rect 3631 10908 3683 10911
rect 3739 10908 3791 10911
rect 3847 10908 3899 10911
rect 5700 10908 5752 10911
rect 5808 10908 5860 10911
rect 5916 10908 5968 10911
rect 6024 10908 6076 10911
rect 6186 10908 6238 10911
rect 6294 10908 6346 10911
rect 6402 10908 6454 10911
rect 6510 10908 6562 10911
rect 8363 10908 8415 10911
rect 8471 10908 8523 10911
rect 8579 10908 8631 10911
rect 8687 10908 8739 10911
rect 8795 10908 8847 10911
rect 10635 10908 10687 10911
rect 10743 10908 10795 10911
rect 10851 10908 10903 10911
rect 10959 10908 11011 10911
rect 11067 10908 11119 10911
rect 1143 10803 1195 10852
rect 1251 10803 1303 10852
rect 1359 10803 1411 10852
rect 1467 10803 1519 10852
rect 1575 10803 1627 10852
rect 3415 10803 3467 10852
rect 3523 10803 3575 10852
rect 3631 10803 3683 10852
rect 3739 10803 3791 10852
rect 3847 10803 3899 10852
rect 5700 10803 5752 10852
rect 5808 10803 5860 10852
rect 5916 10803 5968 10852
rect 6024 10803 6076 10852
rect 6186 10803 6238 10852
rect 6294 10803 6346 10852
rect 6402 10803 6454 10852
rect 6510 10803 6562 10852
rect 8363 10803 8415 10852
rect 8471 10803 8523 10852
rect 8579 10803 8631 10852
rect 8687 10803 8739 10852
rect 8795 10803 8847 10852
rect 10635 10803 10687 10852
rect 10743 10803 10795 10852
rect 10851 10803 10903 10852
rect 10959 10803 11011 10852
rect 11067 10803 11119 10852
rect 1143 10800 1195 10803
rect 1251 10800 1303 10803
rect 1359 10800 1411 10803
rect 1467 10800 1519 10803
rect 1575 10800 1627 10803
rect 3415 10800 3467 10803
rect 3523 10800 3575 10803
rect 3631 10800 3683 10803
rect 3739 10800 3791 10803
rect 3847 10800 3899 10803
rect 5700 10800 5752 10803
rect 5808 10800 5860 10803
rect 5916 10800 5968 10803
rect 6024 10800 6076 10803
rect 6186 10800 6238 10803
rect 6294 10800 6346 10803
rect 6402 10800 6454 10803
rect 6510 10800 6562 10803
rect 8363 10800 8415 10803
rect 8471 10800 8523 10803
rect 8579 10800 8631 10803
rect 8687 10800 8739 10803
rect 8795 10800 8847 10803
rect 10635 10800 10687 10803
rect 10743 10800 10795 10803
rect 10851 10800 10903 10803
rect 10959 10800 11011 10803
rect 11067 10800 11119 10803
rect 1741 10473 1793 10506
rect 1865 10473 1917 10506
rect 1989 10473 2041 10506
rect 2113 10473 2165 10506
rect 2877 10473 2929 10506
rect 3001 10473 3053 10506
rect 3125 10473 3177 10506
rect 3249 10473 3301 10506
rect 4013 10473 4065 10506
rect 4137 10473 4189 10506
rect 4261 10473 4313 10506
rect 4385 10473 4437 10506
rect 5149 10473 5201 10506
rect 5273 10473 5325 10506
rect 5397 10473 5449 10506
rect 5521 10473 5573 10506
rect 6689 10473 6741 10506
rect 6813 10473 6865 10506
rect 6937 10473 6989 10506
rect 7061 10473 7113 10506
rect 7825 10473 7877 10506
rect 7949 10473 8001 10506
rect 8073 10473 8125 10506
rect 8197 10473 8249 10506
rect 8961 10473 9013 10506
rect 9085 10473 9137 10506
rect 9209 10473 9261 10506
rect 9333 10473 9385 10506
rect 10097 10473 10149 10506
rect 10221 10473 10273 10506
rect 10345 10473 10397 10506
rect 10469 10473 10521 10506
rect 1741 10454 1793 10473
rect 1865 10454 1917 10473
rect 1989 10454 2041 10473
rect 2113 10454 2165 10473
rect 2877 10454 2929 10473
rect 3001 10454 3053 10473
rect 3125 10454 3177 10473
rect 3249 10454 3301 10473
rect 4013 10454 4065 10473
rect 4137 10454 4189 10473
rect 4261 10454 4313 10473
rect 4385 10454 4437 10473
rect 5149 10454 5201 10473
rect 5273 10454 5325 10473
rect 5397 10454 5449 10473
rect 5521 10454 5573 10473
rect 6689 10454 6741 10473
rect 6813 10454 6865 10473
rect 6937 10454 6989 10473
rect 7061 10454 7113 10473
rect 7825 10454 7877 10473
rect 7949 10454 8001 10473
rect 8073 10454 8125 10473
rect 8197 10454 8249 10473
rect 8961 10454 9013 10473
rect 9085 10454 9137 10473
rect 9209 10454 9261 10473
rect 9333 10454 9385 10473
rect 10097 10454 10149 10473
rect 10221 10454 10273 10473
rect 10345 10454 10397 10473
rect 10469 10454 10521 10473
rect 1741 10368 1793 10382
rect 1865 10368 1917 10382
rect 1989 10368 2041 10382
rect 2113 10368 2165 10382
rect 2877 10368 2929 10382
rect 3001 10368 3053 10382
rect 3125 10368 3177 10382
rect 3249 10368 3301 10382
rect 4013 10368 4065 10382
rect 4137 10368 4189 10382
rect 4261 10368 4313 10382
rect 4385 10368 4437 10382
rect 5149 10368 5201 10382
rect 5273 10368 5325 10382
rect 5397 10368 5449 10382
rect 5521 10368 5573 10382
rect 6689 10368 6741 10382
rect 6813 10368 6865 10382
rect 6937 10368 6989 10382
rect 7061 10368 7113 10382
rect 7825 10368 7877 10382
rect 7949 10368 8001 10382
rect 8073 10368 8125 10382
rect 8197 10368 8249 10382
rect 8961 10368 9013 10382
rect 9085 10368 9137 10382
rect 9209 10368 9261 10382
rect 9333 10368 9385 10382
rect 10097 10368 10149 10382
rect 10221 10368 10273 10382
rect 10345 10368 10397 10382
rect 10469 10368 10521 10382
rect 1741 10330 1793 10368
rect 1865 10330 1917 10368
rect 1989 10330 2041 10368
rect 2113 10330 2165 10368
rect 2877 10330 2929 10368
rect 3001 10330 3053 10368
rect 3125 10330 3177 10368
rect 3249 10330 3301 10368
rect 4013 10330 4065 10368
rect 4137 10330 4189 10368
rect 4261 10330 4313 10368
rect 4385 10330 4437 10368
rect 5149 10330 5201 10368
rect 5273 10330 5325 10368
rect 5397 10330 5449 10368
rect 5521 10330 5573 10368
rect 6689 10330 6741 10368
rect 6813 10330 6865 10368
rect 6937 10330 6989 10368
rect 7061 10330 7113 10368
rect 7825 10330 7877 10368
rect 7949 10330 8001 10368
rect 8073 10330 8125 10368
rect 8197 10330 8249 10368
rect 8961 10330 9013 10368
rect 9085 10330 9137 10368
rect 9209 10330 9261 10368
rect 9333 10330 9385 10368
rect 10097 10330 10149 10368
rect 10221 10330 10273 10368
rect 10345 10330 10397 10368
rect 10469 10330 10521 10368
rect 1741 10206 1793 10258
rect 1865 10206 1917 10258
rect 1989 10206 2041 10258
rect 2113 10206 2165 10258
rect 2877 10206 2929 10258
rect 3001 10206 3053 10258
rect 3125 10206 3177 10258
rect 3249 10206 3301 10258
rect 4013 10206 4065 10258
rect 4137 10206 4189 10258
rect 4261 10206 4313 10258
rect 4385 10206 4437 10258
rect 5149 10206 5201 10258
rect 5273 10206 5325 10258
rect 5397 10206 5449 10258
rect 5521 10206 5573 10258
rect 6689 10206 6741 10258
rect 6813 10206 6865 10258
rect 6937 10206 6989 10258
rect 7061 10206 7113 10258
rect 7825 10206 7877 10258
rect 7949 10206 8001 10258
rect 8073 10206 8125 10258
rect 8197 10206 8249 10258
rect 8961 10206 9013 10258
rect 9085 10206 9137 10258
rect 9209 10206 9261 10258
rect 9333 10206 9385 10258
rect 10097 10206 10149 10258
rect 10221 10206 10273 10258
rect 10345 10206 10397 10258
rect 10469 10206 10521 10258
rect 1741 10097 1793 10134
rect 1865 10097 1917 10134
rect 1989 10097 2041 10134
rect 2113 10097 2165 10134
rect 2877 10097 2929 10134
rect 3001 10097 3053 10134
rect 3125 10097 3177 10134
rect 3249 10097 3301 10134
rect 4013 10097 4065 10134
rect 4137 10097 4189 10134
rect 4261 10097 4313 10134
rect 4385 10097 4437 10134
rect 5149 10097 5201 10134
rect 5273 10097 5325 10134
rect 5397 10097 5449 10134
rect 5521 10097 5573 10134
rect 6689 10097 6741 10134
rect 6813 10097 6865 10134
rect 6937 10097 6989 10134
rect 7061 10097 7113 10134
rect 7825 10097 7877 10134
rect 7949 10097 8001 10134
rect 8073 10097 8125 10134
rect 8197 10097 8249 10134
rect 8961 10097 9013 10134
rect 9085 10097 9137 10134
rect 9209 10097 9261 10134
rect 9333 10097 9385 10134
rect 10097 10097 10149 10134
rect 10221 10097 10273 10134
rect 10345 10097 10397 10134
rect 10469 10097 10521 10134
rect 1741 10082 1793 10097
rect 1865 10082 1917 10097
rect 1989 10082 2041 10097
rect 2113 10082 2165 10097
rect 2877 10082 2929 10097
rect 3001 10082 3053 10097
rect 3125 10082 3177 10097
rect 3249 10082 3301 10097
rect 4013 10082 4065 10097
rect 4137 10082 4189 10097
rect 4261 10082 4313 10097
rect 4385 10082 4437 10097
rect 5149 10082 5201 10097
rect 5273 10082 5325 10097
rect 5397 10082 5449 10097
rect 5521 10082 5573 10097
rect 6689 10082 6741 10097
rect 6813 10082 6865 10097
rect 6937 10082 6989 10097
rect 7061 10082 7113 10097
rect 7825 10082 7877 10097
rect 7949 10082 8001 10097
rect 8073 10082 8125 10097
rect 8197 10082 8249 10097
rect 8961 10082 9013 10097
rect 9085 10082 9137 10097
rect 9209 10082 9261 10097
rect 9333 10082 9385 10097
rect 10097 10082 10149 10097
rect 10221 10082 10273 10097
rect 10345 10082 10397 10097
rect 10469 10082 10521 10097
rect 1741 9991 1793 10010
rect 1865 9991 1917 10010
rect 1989 9991 2041 10010
rect 2113 9991 2165 10010
rect 2877 9991 2929 10010
rect 3001 9991 3053 10010
rect 3125 9991 3177 10010
rect 3249 9991 3301 10010
rect 4013 9991 4065 10010
rect 4137 9991 4189 10010
rect 4261 9991 4313 10010
rect 4385 9991 4437 10010
rect 5149 9991 5201 10010
rect 5273 9991 5325 10010
rect 5397 9991 5449 10010
rect 5521 9991 5573 10010
rect 6689 9991 6741 10010
rect 6813 9991 6865 10010
rect 6937 9991 6989 10010
rect 7061 9991 7113 10010
rect 7825 9991 7877 10010
rect 7949 9991 8001 10010
rect 8073 9991 8125 10010
rect 8197 9991 8249 10010
rect 8961 9991 9013 10010
rect 9085 9991 9137 10010
rect 9209 9991 9261 10010
rect 9333 9991 9385 10010
rect 10097 9991 10149 10010
rect 10221 9991 10273 10010
rect 10345 9991 10397 10010
rect 10469 9991 10521 10010
rect 1741 9958 1793 9991
rect 1865 9958 1917 9991
rect 1989 9958 2041 9991
rect 2113 9958 2165 9991
rect 2877 9958 2929 9991
rect 3001 9958 3053 9991
rect 3125 9958 3177 9991
rect 3249 9958 3301 9991
rect 4013 9958 4065 9991
rect 4137 9958 4189 9991
rect 4261 9958 4313 9991
rect 4385 9958 4437 9991
rect 5149 9958 5201 9991
rect 5273 9958 5325 9991
rect 5397 9958 5449 9991
rect 5521 9958 5573 9991
rect 6689 9958 6741 9991
rect 6813 9958 6865 9991
rect 6937 9958 6989 9991
rect 7061 9958 7113 9991
rect 7825 9958 7877 9991
rect 7949 9958 8001 9991
rect 8073 9958 8125 9991
rect 8197 9958 8249 9991
rect 8961 9958 9013 9991
rect 9085 9958 9137 9991
rect 9209 9958 9261 9991
rect 9333 9958 9385 9991
rect 10097 9958 10149 9991
rect 10221 9958 10273 9991
rect 10345 9958 10397 9991
rect 10469 9958 10521 9991
rect 1143 9661 1195 9664
rect 1251 9661 1303 9664
rect 1359 9661 1411 9664
rect 1467 9661 1519 9664
rect 1575 9661 1627 9664
rect 3415 9661 3467 9664
rect 3523 9661 3575 9664
rect 3631 9661 3683 9664
rect 3739 9661 3791 9664
rect 3847 9661 3899 9664
rect 5700 9661 5752 9664
rect 5808 9661 5860 9664
rect 5916 9661 5968 9664
rect 6024 9661 6076 9664
rect 6186 9661 6238 9664
rect 6294 9661 6346 9664
rect 6402 9661 6454 9664
rect 6510 9661 6562 9664
rect 8363 9661 8415 9664
rect 8471 9661 8523 9664
rect 8579 9661 8631 9664
rect 8687 9661 8739 9664
rect 8795 9661 8847 9664
rect 10635 9661 10687 9664
rect 10743 9661 10795 9664
rect 10851 9661 10903 9664
rect 10959 9661 11011 9664
rect 11067 9661 11119 9664
rect 1143 9612 1195 9661
rect 1251 9612 1303 9661
rect 1359 9612 1411 9661
rect 1467 9612 1519 9661
rect 1575 9612 1627 9661
rect 3415 9612 3467 9661
rect 3523 9612 3575 9661
rect 3631 9612 3683 9661
rect 3739 9612 3791 9661
rect 3847 9612 3899 9661
rect 5700 9612 5752 9661
rect 5808 9612 5860 9661
rect 5916 9612 5968 9661
rect 6024 9612 6076 9661
rect 6186 9612 6238 9661
rect 6294 9612 6346 9661
rect 6402 9612 6454 9661
rect 6510 9612 6562 9661
rect 8363 9612 8415 9661
rect 8471 9612 8523 9661
rect 8579 9612 8631 9661
rect 8687 9612 8739 9661
rect 8795 9612 8847 9661
rect 10635 9612 10687 9661
rect 10743 9612 10795 9661
rect 10851 9612 10903 9661
rect 10959 9612 11011 9661
rect 11067 9612 11119 9661
rect 1143 9553 1195 9556
rect 1251 9553 1303 9556
rect 1359 9553 1411 9556
rect 1467 9553 1519 9556
rect 1575 9553 1627 9556
rect 3415 9553 3467 9556
rect 3523 9553 3575 9556
rect 3631 9553 3683 9556
rect 3739 9553 3791 9556
rect 3847 9553 3899 9556
rect 5700 9553 5752 9556
rect 5808 9553 5860 9556
rect 5916 9553 5968 9556
rect 6024 9553 6076 9556
rect 6186 9553 6238 9556
rect 6294 9553 6346 9556
rect 6402 9553 6454 9556
rect 6510 9553 6562 9556
rect 8363 9553 8415 9556
rect 8471 9553 8523 9556
rect 8579 9553 8631 9556
rect 8687 9553 8739 9556
rect 8795 9553 8847 9556
rect 10635 9553 10687 9556
rect 10743 9553 10795 9556
rect 10851 9553 10903 9556
rect 10959 9553 11011 9556
rect 11067 9553 11119 9556
rect 1143 9507 1195 9553
rect 1251 9507 1303 9553
rect 1359 9507 1411 9553
rect 1467 9507 1519 9553
rect 1575 9507 1627 9553
rect 3415 9507 3467 9553
rect 3523 9507 3575 9553
rect 3631 9507 3683 9553
rect 3739 9507 3791 9553
rect 3847 9507 3899 9553
rect 5700 9507 5752 9553
rect 5808 9507 5860 9553
rect 5916 9507 5968 9553
rect 6024 9507 6076 9553
rect 6186 9507 6238 9553
rect 6294 9507 6346 9553
rect 6402 9507 6454 9553
rect 6510 9507 6562 9553
rect 8363 9507 8415 9553
rect 8471 9507 8523 9553
rect 8579 9507 8631 9553
rect 8687 9507 8739 9553
rect 8795 9507 8847 9553
rect 10635 9507 10687 9553
rect 10743 9507 10795 9553
rect 10851 9507 10903 9553
rect 10959 9507 11011 9553
rect 11067 9507 11119 9553
rect 1143 9504 1195 9507
rect 1251 9504 1303 9507
rect 1359 9504 1411 9507
rect 1467 9504 1519 9507
rect 1575 9504 1627 9507
rect 3415 9504 3467 9507
rect 3523 9504 3575 9507
rect 3631 9504 3683 9507
rect 3739 9504 3791 9507
rect 3847 9504 3899 9507
rect 5700 9504 5752 9507
rect 5808 9504 5860 9507
rect 5916 9504 5968 9507
rect 6024 9504 6076 9507
rect 6186 9504 6238 9507
rect 6294 9504 6346 9507
rect 6402 9504 6454 9507
rect 6510 9504 6562 9507
rect 8363 9504 8415 9507
rect 8471 9504 8523 9507
rect 8579 9504 8631 9507
rect 8687 9504 8739 9507
rect 8795 9504 8847 9507
rect 10635 9504 10687 9507
rect 10743 9504 10795 9507
rect 10851 9504 10903 9507
rect 10959 9504 11011 9507
rect 11067 9504 11119 9507
rect 1143 9399 1195 9448
rect 1251 9399 1303 9448
rect 1359 9399 1411 9448
rect 1467 9399 1519 9448
rect 1575 9399 1627 9448
rect 3415 9399 3467 9448
rect 3523 9399 3575 9448
rect 3631 9399 3683 9448
rect 3739 9399 3791 9448
rect 3847 9399 3899 9448
rect 5700 9399 5752 9448
rect 5808 9399 5860 9448
rect 5916 9399 5968 9448
rect 6024 9399 6076 9448
rect 6186 9399 6238 9448
rect 6294 9399 6346 9448
rect 6402 9399 6454 9448
rect 6510 9399 6562 9448
rect 8363 9399 8415 9448
rect 8471 9399 8523 9448
rect 8579 9399 8631 9448
rect 8687 9399 8739 9448
rect 8795 9399 8847 9448
rect 10635 9399 10687 9448
rect 10743 9399 10795 9448
rect 10851 9399 10903 9448
rect 10959 9399 11011 9448
rect 11067 9399 11119 9448
rect 1143 9396 1195 9399
rect 1251 9396 1303 9399
rect 1359 9396 1411 9399
rect 1467 9396 1519 9399
rect 1575 9396 1627 9399
rect 3415 9396 3467 9399
rect 3523 9396 3575 9399
rect 3631 9396 3683 9399
rect 3739 9396 3791 9399
rect 3847 9396 3899 9399
rect 5700 9396 5752 9399
rect 5808 9396 5860 9399
rect 5916 9396 5968 9399
rect 6024 9396 6076 9399
rect 6186 9396 6238 9399
rect 6294 9396 6346 9399
rect 6402 9396 6454 9399
rect 6510 9396 6562 9399
rect 8363 9396 8415 9399
rect 8471 9396 8523 9399
rect 8579 9396 8631 9399
rect 8687 9396 8739 9399
rect 8795 9396 8847 9399
rect 10635 9396 10687 9399
rect 10743 9396 10795 9399
rect 10851 9396 10903 9399
rect 10959 9396 11011 9399
rect 11067 9396 11119 9399
rect 1741 9069 1793 9102
rect 1865 9069 1917 9102
rect 1989 9069 2041 9102
rect 2113 9069 2165 9102
rect 2877 9069 2929 9102
rect 3001 9069 3053 9102
rect 3125 9069 3177 9102
rect 3249 9069 3301 9102
rect 4013 9069 4065 9102
rect 4137 9069 4189 9102
rect 4261 9069 4313 9102
rect 4385 9069 4437 9102
rect 5149 9069 5201 9102
rect 5273 9069 5325 9102
rect 5397 9069 5449 9102
rect 5521 9069 5573 9102
rect 6689 9069 6741 9102
rect 6813 9069 6865 9102
rect 6937 9069 6989 9102
rect 7061 9069 7113 9102
rect 7825 9069 7877 9102
rect 7949 9069 8001 9102
rect 8073 9069 8125 9102
rect 8197 9069 8249 9102
rect 8961 9069 9013 9102
rect 9085 9069 9137 9102
rect 9209 9069 9261 9102
rect 9333 9069 9385 9102
rect 10097 9069 10149 9102
rect 10221 9069 10273 9102
rect 10345 9069 10397 9102
rect 10469 9069 10521 9102
rect 1741 9050 1793 9069
rect 1865 9050 1917 9069
rect 1989 9050 2041 9069
rect 2113 9050 2165 9069
rect 2877 9050 2929 9069
rect 3001 9050 3053 9069
rect 3125 9050 3177 9069
rect 3249 9050 3301 9069
rect 4013 9050 4065 9069
rect 4137 9050 4189 9069
rect 4261 9050 4313 9069
rect 4385 9050 4437 9069
rect 5149 9050 5201 9069
rect 5273 9050 5325 9069
rect 5397 9050 5449 9069
rect 5521 9050 5573 9069
rect 6689 9050 6741 9069
rect 6813 9050 6865 9069
rect 6937 9050 6989 9069
rect 7061 9050 7113 9069
rect 7825 9050 7877 9069
rect 7949 9050 8001 9069
rect 8073 9050 8125 9069
rect 8197 9050 8249 9069
rect 8961 9050 9013 9069
rect 9085 9050 9137 9069
rect 9209 9050 9261 9069
rect 9333 9050 9385 9069
rect 10097 9050 10149 9069
rect 10221 9050 10273 9069
rect 10345 9050 10397 9069
rect 10469 9050 10521 9069
rect 1741 8964 1793 8978
rect 1865 8964 1917 8978
rect 1989 8964 2041 8978
rect 2113 8964 2165 8978
rect 2877 8964 2929 8978
rect 3001 8964 3053 8978
rect 3125 8964 3177 8978
rect 3249 8964 3301 8978
rect 4013 8964 4065 8978
rect 4137 8964 4189 8978
rect 4261 8964 4313 8978
rect 4385 8964 4437 8978
rect 5149 8964 5201 8978
rect 5273 8964 5325 8978
rect 5397 8964 5449 8978
rect 5521 8964 5573 8978
rect 6689 8964 6741 8978
rect 6813 8964 6865 8978
rect 6937 8964 6989 8978
rect 7061 8964 7113 8978
rect 7825 8964 7877 8978
rect 7949 8964 8001 8978
rect 8073 8964 8125 8978
rect 8197 8964 8249 8978
rect 8961 8964 9013 8978
rect 9085 8964 9137 8978
rect 9209 8964 9261 8978
rect 9333 8964 9385 8978
rect 10097 8964 10149 8978
rect 10221 8964 10273 8978
rect 10345 8964 10397 8978
rect 10469 8964 10521 8978
rect 1741 8926 1793 8964
rect 1865 8926 1917 8964
rect 1989 8926 2041 8964
rect 2113 8926 2165 8964
rect 2877 8926 2929 8964
rect 3001 8926 3053 8964
rect 3125 8926 3177 8964
rect 3249 8926 3301 8964
rect 4013 8926 4065 8964
rect 4137 8926 4189 8964
rect 4261 8926 4313 8964
rect 4385 8926 4437 8964
rect 5149 8926 5201 8964
rect 5273 8926 5325 8964
rect 5397 8926 5449 8964
rect 5521 8926 5573 8964
rect 6689 8926 6741 8964
rect 6813 8926 6865 8964
rect 6937 8926 6989 8964
rect 7061 8926 7113 8964
rect 7825 8926 7877 8964
rect 7949 8926 8001 8964
rect 8073 8926 8125 8964
rect 8197 8926 8249 8964
rect 8961 8926 9013 8964
rect 9085 8926 9137 8964
rect 9209 8926 9261 8964
rect 9333 8926 9385 8964
rect 10097 8926 10149 8964
rect 10221 8926 10273 8964
rect 10345 8926 10397 8964
rect 10469 8926 10521 8964
rect 1741 8802 1793 8854
rect 1865 8802 1917 8854
rect 1989 8802 2041 8854
rect 2113 8802 2165 8854
rect 2877 8802 2929 8854
rect 3001 8802 3053 8854
rect 3125 8802 3177 8854
rect 3249 8802 3301 8854
rect 4013 8802 4065 8854
rect 4137 8802 4189 8854
rect 4261 8802 4313 8854
rect 4385 8802 4437 8854
rect 5149 8802 5201 8854
rect 5273 8802 5325 8854
rect 5397 8802 5449 8854
rect 5521 8802 5573 8854
rect 6689 8802 6741 8854
rect 6813 8802 6865 8854
rect 6937 8802 6989 8854
rect 7061 8802 7113 8854
rect 7825 8802 7877 8854
rect 7949 8802 8001 8854
rect 8073 8802 8125 8854
rect 8197 8802 8249 8854
rect 8961 8802 9013 8854
rect 9085 8802 9137 8854
rect 9209 8802 9261 8854
rect 9333 8802 9385 8854
rect 10097 8802 10149 8854
rect 10221 8802 10273 8854
rect 10345 8802 10397 8854
rect 10469 8802 10521 8854
rect 1741 8693 1793 8730
rect 1865 8693 1917 8730
rect 1989 8693 2041 8730
rect 2113 8693 2165 8730
rect 2877 8693 2929 8730
rect 3001 8693 3053 8730
rect 3125 8693 3177 8730
rect 3249 8693 3301 8730
rect 4013 8693 4065 8730
rect 4137 8693 4189 8730
rect 4261 8693 4313 8730
rect 4385 8693 4437 8730
rect 5149 8693 5201 8730
rect 5273 8693 5325 8730
rect 5397 8693 5449 8730
rect 5521 8693 5573 8730
rect 6689 8693 6741 8730
rect 6813 8693 6865 8730
rect 6937 8693 6989 8730
rect 7061 8693 7113 8730
rect 7825 8693 7877 8730
rect 7949 8693 8001 8730
rect 8073 8693 8125 8730
rect 8197 8693 8249 8730
rect 8961 8693 9013 8730
rect 9085 8693 9137 8730
rect 9209 8693 9261 8730
rect 9333 8693 9385 8730
rect 10097 8693 10149 8730
rect 10221 8693 10273 8730
rect 10345 8693 10397 8730
rect 10469 8693 10521 8730
rect 1741 8678 1793 8693
rect 1865 8678 1917 8693
rect 1989 8678 2041 8693
rect 2113 8678 2165 8693
rect 2877 8678 2929 8693
rect 3001 8678 3053 8693
rect 3125 8678 3177 8693
rect 3249 8678 3301 8693
rect 4013 8678 4065 8693
rect 4137 8678 4189 8693
rect 4261 8678 4313 8693
rect 4385 8678 4437 8693
rect 5149 8678 5201 8693
rect 5273 8678 5325 8693
rect 5397 8678 5449 8693
rect 5521 8678 5573 8693
rect 6689 8678 6741 8693
rect 6813 8678 6865 8693
rect 6937 8678 6989 8693
rect 7061 8678 7113 8693
rect 7825 8678 7877 8693
rect 7949 8678 8001 8693
rect 8073 8678 8125 8693
rect 8197 8678 8249 8693
rect 8961 8678 9013 8693
rect 9085 8678 9137 8693
rect 9209 8678 9261 8693
rect 9333 8678 9385 8693
rect 10097 8678 10149 8693
rect 10221 8678 10273 8693
rect 10345 8678 10397 8693
rect 10469 8678 10521 8693
rect 1741 8587 1793 8606
rect 1865 8587 1917 8606
rect 1989 8587 2041 8606
rect 2113 8587 2165 8606
rect 2877 8587 2929 8606
rect 3001 8587 3053 8606
rect 3125 8587 3177 8606
rect 3249 8587 3301 8606
rect 4013 8587 4065 8606
rect 4137 8587 4189 8606
rect 4261 8587 4313 8606
rect 4385 8587 4437 8606
rect 5149 8587 5201 8606
rect 5273 8587 5325 8606
rect 5397 8587 5449 8606
rect 5521 8587 5573 8606
rect 6689 8587 6741 8606
rect 6813 8587 6865 8606
rect 6937 8587 6989 8606
rect 7061 8587 7113 8606
rect 7825 8587 7877 8606
rect 7949 8587 8001 8606
rect 8073 8587 8125 8606
rect 8197 8587 8249 8606
rect 8961 8587 9013 8606
rect 9085 8587 9137 8606
rect 9209 8587 9261 8606
rect 9333 8587 9385 8606
rect 10097 8587 10149 8606
rect 10221 8587 10273 8606
rect 10345 8587 10397 8606
rect 10469 8587 10521 8606
rect 1741 8554 1793 8587
rect 1865 8554 1917 8587
rect 1989 8554 2041 8587
rect 2113 8554 2165 8587
rect 2877 8554 2929 8587
rect 3001 8554 3053 8587
rect 3125 8554 3177 8587
rect 3249 8554 3301 8587
rect 4013 8554 4065 8587
rect 4137 8554 4189 8587
rect 4261 8554 4313 8587
rect 4385 8554 4437 8587
rect 5149 8554 5201 8587
rect 5273 8554 5325 8587
rect 5397 8554 5449 8587
rect 5521 8554 5573 8587
rect 6689 8554 6741 8587
rect 6813 8554 6865 8587
rect 6937 8554 6989 8587
rect 7061 8554 7113 8587
rect 7825 8554 7877 8587
rect 7949 8554 8001 8587
rect 8073 8554 8125 8587
rect 8197 8554 8249 8587
rect 8961 8554 9013 8587
rect 9085 8554 9137 8587
rect 9209 8554 9261 8587
rect 9333 8554 9385 8587
rect 10097 8554 10149 8587
rect 10221 8554 10273 8587
rect 10345 8554 10397 8587
rect 10469 8554 10521 8587
rect 1143 8257 1195 8283
rect 1251 8257 1303 8283
rect 1359 8257 1411 8283
rect 1467 8257 1519 8283
rect 1575 8257 1627 8283
rect 3415 8257 3467 8283
rect 3523 8257 3575 8283
rect 3631 8257 3683 8283
rect 3739 8257 3791 8283
rect 3847 8257 3899 8283
rect 5700 8257 5752 8283
rect 5808 8257 5860 8283
rect 5916 8257 5968 8283
rect 6024 8257 6076 8283
rect 6186 8257 6238 8283
rect 6294 8257 6346 8283
rect 6402 8257 6454 8283
rect 6510 8257 6562 8283
rect 8363 8257 8415 8283
rect 8471 8257 8523 8283
rect 8579 8257 8631 8283
rect 8687 8257 8739 8283
rect 8795 8257 8847 8283
rect 10635 8257 10687 8283
rect 10743 8257 10795 8283
rect 10851 8257 10903 8283
rect 10959 8257 11011 8283
rect 11067 8257 11119 8283
rect 1143 8231 1195 8257
rect 1251 8231 1303 8257
rect 1359 8231 1411 8257
rect 1467 8231 1519 8257
rect 1575 8231 1627 8257
rect 3415 8231 3467 8257
rect 3523 8231 3575 8257
rect 3631 8231 3683 8257
rect 3739 8231 3791 8257
rect 3847 8231 3899 8257
rect 5700 8231 5752 8257
rect 5808 8231 5860 8257
rect 5916 8231 5968 8257
rect 6024 8231 6076 8257
rect 6186 8231 6238 8257
rect 6294 8231 6346 8257
rect 6402 8231 6454 8257
rect 6510 8231 6562 8257
rect 8363 8231 8415 8257
rect 8471 8231 8523 8257
rect 8579 8231 8631 8257
rect 8687 8231 8739 8257
rect 8795 8231 8847 8257
rect 10635 8231 10687 8257
rect 10743 8231 10795 8257
rect 10851 8231 10903 8257
rect 10959 8231 11011 8257
rect 11067 8231 11119 8257
rect 1143 8149 1195 8175
rect 1251 8149 1303 8175
rect 1359 8149 1411 8175
rect 1467 8149 1519 8175
rect 1575 8149 1627 8175
rect 3415 8149 3467 8175
rect 3523 8149 3575 8175
rect 3631 8149 3683 8175
rect 3739 8149 3791 8175
rect 3847 8149 3899 8175
rect 5700 8149 5752 8175
rect 5808 8149 5860 8175
rect 5916 8149 5968 8175
rect 6024 8149 6076 8175
rect 6186 8149 6238 8175
rect 6294 8149 6346 8175
rect 6402 8149 6454 8175
rect 6510 8149 6562 8175
rect 8363 8149 8415 8175
rect 8471 8149 8523 8175
rect 8579 8149 8631 8175
rect 8687 8149 8739 8175
rect 8795 8149 8847 8175
rect 10635 8149 10687 8175
rect 10743 8149 10795 8175
rect 10851 8149 10903 8175
rect 10959 8149 11011 8175
rect 11067 8149 11119 8175
rect 1143 8123 1195 8149
rect 1251 8123 1303 8149
rect 1359 8123 1411 8149
rect 1467 8123 1519 8149
rect 1575 8123 1627 8149
rect 3415 8123 3467 8149
rect 3523 8123 3575 8149
rect 3631 8123 3683 8149
rect 3739 8123 3791 8149
rect 3847 8123 3899 8149
rect 5700 8123 5752 8149
rect 5808 8123 5860 8149
rect 5916 8123 5968 8149
rect 6024 8123 6076 8149
rect 6186 8123 6238 8149
rect 6294 8123 6346 8149
rect 6402 8123 6454 8149
rect 6510 8123 6562 8149
rect 8363 8123 8415 8149
rect 8471 8123 8523 8149
rect 8579 8123 8631 8149
rect 8687 8123 8739 8149
rect 8795 8123 8847 8149
rect 10635 8123 10687 8149
rect 10743 8123 10795 8149
rect 10851 8123 10903 8149
rect 10959 8123 11011 8149
rect 11067 8123 11119 8149
rect 605 7844 608 7896
rect 608 7844 657 7896
rect 729 7844 781 7896
rect 853 7844 905 7896
rect 977 7844 1029 7896
rect 2309 7844 2361 7896
rect 2433 7844 2485 7896
rect 2557 7844 2609 7896
rect 2681 7844 2733 7896
rect 4581 7844 4633 7896
rect 4705 7844 4757 7896
rect 4829 7844 4881 7896
rect 4953 7844 5005 7896
rect 7257 7844 7309 7896
rect 7381 7844 7433 7896
rect 7505 7844 7557 7896
rect 7629 7844 7681 7896
rect 9529 7844 9581 7896
rect 9653 7844 9705 7896
rect 9777 7844 9829 7896
rect 9901 7844 9953 7896
rect 11233 7844 11285 7896
rect 11357 7844 11409 7896
rect 11481 7844 11533 7896
rect 11605 7844 11654 7896
rect 11654 7844 11657 7896
rect 605 7720 608 7772
rect 608 7720 657 7772
rect 729 7720 781 7772
rect 853 7720 905 7772
rect 977 7720 1029 7772
rect 2309 7720 2361 7772
rect 2433 7720 2485 7772
rect 2557 7720 2609 7772
rect 2681 7720 2733 7772
rect 4581 7720 4633 7772
rect 4705 7720 4757 7772
rect 4829 7720 4881 7772
rect 4953 7720 5005 7772
rect 7257 7720 7309 7772
rect 7381 7720 7433 7772
rect 7505 7720 7557 7772
rect 7629 7720 7681 7772
rect 9529 7720 9581 7772
rect 9653 7720 9705 7772
rect 9777 7720 9829 7772
rect 9901 7720 9953 7772
rect 11233 7720 11285 7772
rect 11357 7720 11409 7772
rect 11481 7720 11533 7772
rect 11605 7720 11654 7772
rect 11654 7720 11657 7772
rect 605 7596 608 7648
rect 608 7596 657 7648
rect 729 7596 781 7648
rect 853 7596 905 7648
rect 977 7596 1029 7648
rect 2309 7596 2361 7648
rect 2433 7596 2485 7648
rect 2557 7596 2609 7648
rect 2681 7596 2733 7648
rect 4581 7596 4633 7648
rect 4705 7596 4757 7648
rect 4829 7596 4881 7648
rect 4953 7596 5005 7648
rect 7257 7596 7309 7648
rect 7381 7596 7433 7648
rect 7505 7596 7557 7648
rect 7629 7596 7681 7648
rect 9529 7596 9581 7648
rect 9653 7596 9705 7648
rect 9777 7596 9829 7648
rect 9901 7596 9953 7648
rect 11233 7596 11285 7648
rect 11357 7596 11409 7648
rect 11481 7596 11533 7648
rect 11605 7596 11654 7648
rect 11654 7596 11657 7648
rect 605 7472 608 7524
rect 608 7472 657 7524
rect 729 7472 781 7524
rect 853 7472 905 7524
rect 977 7472 1029 7524
rect 2309 7472 2361 7524
rect 2433 7472 2485 7524
rect 2557 7472 2609 7524
rect 2681 7472 2733 7524
rect 4581 7472 4633 7524
rect 4705 7472 4757 7524
rect 4829 7472 4881 7524
rect 4953 7472 5005 7524
rect 7257 7472 7309 7524
rect 7381 7472 7433 7524
rect 7505 7472 7557 7524
rect 7629 7472 7681 7524
rect 9529 7472 9581 7524
rect 9653 7472 9705 7524
rect 9777 7472 9829 7524
rect 9901 7472 9953 7524
rect 11233 7472 11285 7524
rect 11357 7472 11409 7524
rect 11481 7472 11533 7524
rect 11605 7472 11654 7524
rect 11654 7472 11657 7524
rect 189 6903 241 6955
rect 297 6903 349 6955
rect 405 6903 457 6955
rect 189 6795 241 6847
rect 297 6795 349 6847
rect 405 6795 457 6847
rect 189 6687 241 6739
rect 297 6687 349 6739
rect 405 6687 457 6739
rect 189 6579 241 6631
rect 297 6579 349 6631
rect 405 6579 457 6631
rect 1173 6937 1225 6989
rect 1297 6937 1349 6989
rect 1421 6937 1473 6989
rect 1545 6937 1597 6989
rect 3445 6937 3497 6989
rect 3569 6937 3621 6989
rect 3693 6937 3745 6989
rect 3817 6937 3869 6989
rect 5738 6937 5790 6989
rect 5862 6937 5914 6989
rect 5986 6937 6038 6989
rect 6224 6937 6276 6989
rect 6348 6937 6400 6989
rect 6472 6937 6524 6989
rect 8393 6937 8445 6989
rect 8517 6937 8569 6989
rect 8641 6937 8693 6989
rect 8765 6937 8817 6989
rect 10665 6937 10717 6989
rect 10789 6937 10841 6989
rect 10913 6937 10965 6989
rect 11037 6937 11089 6989
rect 1173 6813 1225 6865
rect 1297 6813 1349 6865
rect 1421 6813 1473 6865
rect 1545 6813 1597 6865
rect 3445 6813 3497 6865
rect 3569 6813 3621 6865
rect 3693 6813 3745 6865
rect 3817 6813 3869 6865
rect 5738 6813 5790 6865
rect 5862 6813 5914 6865
rect 5986 6813 6038 6865
rect 6224 6813 6276 6865
rect 6348 6813 6400 6865
rect 6472 6813 6524 6865
rect 8393 6813 8445 6865
rect 8517 6813 8569 6865
rect 8641 6813 8693 6865
rect 8765 6813 8817 6865
rect 10665 6813 10717 6865
rect 10789 6813 10841 6865
rect 10913 6813 10965 6865
rect 11037 6813 11089 6865
rect 1173 6689 1225 6741
rect 1297 6689 1349 6741
rect 1421 6689 1473 6741
rect 1545 6689 1597 6741
rect 3445 6689 3497 6741
rect 3569 6689 3621 6741
rect 3693 6689 3745 6741
rect 3817 6689 3869 6741
rect 5738 6689 5790 6741
rect 5862 6689 5914 6741
rect 5986 6689 6038 6741
rect 6224 6689 6276 6741
rect 6348 6689 6400 6741
rect 6472 6689 6524 6741
rect 8393 6689 8445 6741
rect 8517 6689 8569 6741
rect 8641 6689 8693 6741
rect 8765 6689 8817 6741
rect 10665 6689 10717 6741
rect 10789 6689 10841 6741
rect 10913 6689 10965 6741
rect 11037 6689 11089 6741
rect 1173 6565 1225 6617
rect 1297 6565 1349 6617
rect 1421 6565 1473 6617
rect 1545 6565 1597 6617
rect 3445 6565 3497 6617
rect 3569 6565 3621 6617
rect 3693 6565 3745 6617
rect 3817 6565 3869 6617
rect 5738 6565 5790 6617
rect 5862 6565 5914 6617
rect 5986 6565 6038 6617
rect 6224 6565 6276 6617
rect 6348 6565 6400 6617
rect 6472 6565 6524 6617
rect 8393 6565 8445 6617
rect 8517 6565 8569 6617
rect 8641 6565 8693 6617
rect 8765 6565 8817 6617
rect 10665 6565 10717 6617
rect 10789 6565 10841 6617
rect 10913 6565 10965 6617
rect 11037 6565 11089 6617
rect 11805 6903 11857 6955
rect 11913 6903 11965 6955
rect 12021 6903 12073 6955
rect 11805 6795 11857 6847
rect 11913 6795 11965 6847
rect 12021 6795 12073 6847
rect 11805 6687 11857 6739
rect 11913 6687 11965 6739
rect 12021 6687 12073 6739
rect 11805 6579 11857 6631
rect 11913 6579 11965 6631
rect 12021 6579 12073 6631
rect 189 6471 241 6523
rect 297 6471 349 6523
rect 405 6471 457 6523
rect 189 6363 241 6415
rect 297 6363 349 6415
rect 405 6363 457 6415
rect 189 6255 241 6307
rect 297 6255 349 6307
rect 405 6255 457 6307
rect 189 6147 241 6199
rect 297 6147 349 6199
rect 405 6147 457 6199
rect 189 6039 241 6091
rect 297 6039 349 6091
rect 405 6039 457 6091
rect 189 5931 241 5983
rect 297 5931 349 5983
rect 405 5931 457 5983
rect 189 5823 241 5875
rect 297 5823 349 5875
rect 405 5823 457 5875
rect 189 5715 241 5767
rect 297 5715 349 5767
rect 405 5715 457 5767
rect 189 5607 241 5659
rect 297 5607 349 5659
rect 405 5607 457 5659
rect 189 5499 241 5551
rect 297 5499 349 5551
rect 405 5499 457 5551
rect 189 5391 241 5443
rect 297 5391 349 5443
rect 405 5391 457 5443
rect 189 5283 241 5335
rect 297 5283 349 5335
rect 405 5283 457 5335
rect 189 5175 241 5227
rect 297 5175 349 5227
rect 405 5175 457 5227
rect 189 5067 241 5119
rect 297 5067 349 5119
rect 405 5067 457 5119
rect 189 4959 241 5011
rect 297 4959 349 5011
rect 405 4959 457 5011
rect 189 4851 241 4903
rect 297 4851 349 4903
rect 405 4851 457 4903
rect 189 4743 241 4795
rect 297 4743 349 4795
rect 405 4743 457 4795
rect 189 4635 241 4687
rect 297 4635 349 4687
rect 405 4635 457 4687
rect 189 4527 241 4579
rect 297 4527 349 4579
rect 405 4527 457 4579
rect 189 4419 241 4471
rect 297 4419 349 4471
rect 405 4419 457 4471
rect 189 4311 241 4363
rect 297 4311 349 4363
rect 405 4311 457 4363
rect 189 4203 241 4255
rect 297 4203 349 4255
rect 405 4203 457 4255
rect 189 4095 241 4147
rect 297 4095 349 4147
rect 405 4095 457 4147
rect 189 3987 241 4039
rect 297 3987 349 4039
rect 405 3987 457 4039
rect 189 3879 241 3931
rect 297 3879 349 3931
rect 405 3879 457 3931
rect 189 3771 241 3823
rect 297 3771 349 3823
rect 405 3771 457 3823
rect 189 3663 241 3715
rect 297 3663 349 3715
rect 405 3663 457 3715
rect 189 3555 241 3607
rect 297 3555 349 3607
rect 405 3555 457 3607
rect 189 3447 241 3499
rect 297 3447 349 3499
rect 405 3447 457 3499
rect 189 3339 241 3391
rect 297 3339 349 3391
rect 405 3339 457 3391
rect 189 3231 241 3283
rect 297 3231 349 3283
rect 405 3231 457 3283
rect 189 3123 241 3175
rect 297 3123 349 3175
rect 405 3123 457 3175
rect 189 3015 241 3067
rect 297 3015 349 3067
rect 405 3015 457 3067
rect 189 2907 241 2959
rect 297 2907 349 2959
rect 405 2907 457 2959
rect 189 2799 241 2851
rect 297 2799 349 2851
rect 405 2799 457 2851
rect 189 2691 241 2743
rect 297 2691 349 2743
rect 405 2691 457 2743
rect 189 2583 241 2635
rect 297 2583 349 2635
rect 405 2583 457 2635
rect 189 2475 241 2527
rect 297 2475 349 2527
rect 405 2475 457 2527
rect 189 2367 241 2419
rect 297 2367 349 2419
rect 405 2367 457 2419
rect 189 2259 241 2311
rect 297 2259 349 2311
rect 405 2259 457 2311
rect 189 2151 241 2203
rect 297 2151 349 2203
rect 405 2151 457 2203
rect 189 2043 241 2095
rect 297 2043 349 2095
rect 405 2043 457 2095
rect 189 1935 241 1987
rect 297 1935 349 1987
rect 405 1935 457 1987
rect 189 1827 241 1879
rect 297 1827 349 1879
rect 405 1827 457 1879
rect 189 1719 241 1771
rect 297 1719 349 1771
rect 405 1719 457 1771
rect 189 1611 241 1663
rect 297 1611 349 1663
rect 405 1611 457 1663
rect 189 1503 241 1555
rect 297 1503 349 1555
rect 405 1503 457 1555
rect 189 1395 241 1447
rect 297 1395 349 1447
rect 405 1395 457 1447
rect 189 1287 241 1339
rect 297 1287 349 1339
rect 405 1287 457 1339
rect 189 1179 241 1231
rect 297 1179 349 1231
rect 405 1179 457 1231
rect 189 1071 241 1123
rect 297 1071 349 1123
rect 405 1071 457 1123
rect 189 963 241 1015
rect 297 963 349 1015
rect 405 963 457 1015
rect 189 855 241 907
rect 297 855 349 907
rect 405 855 457 907
rect 189 747 241 799
rect 297 747 349 799
rect 405 747 457 799
rect 189 639 241 691
rect 297 639 349 691
rect 405 639 457 691
rect 189 531 241 583
rect 297 531 349 583
rect 405 531 457 583
rect 2279 6312 2331 6338
rect 2387 6312 2439 6338
rect 2495 6312 2547 6338
rect 2603 6312 2655 6338
rect 2711 6312 2763 6338
rect 4551 6312 4603 6338
rect 4659 6312 4711 6338
rect 4767 6312 4819 6338
rect 4875 6312 4927 6338
rect 4983 6312 5035 6338
rect 7227 6312 7279 6338
rect 7335 6312 7387 6338
rect 7443 6312 7495 6338
rect 7551 6312 7603 6338
rect 7659 6312 7711 6338
rect 9499 6312 9551 6338
rect 9607 6312 9659 6338
rect 9715 6312 9767 6338
rect 9823 6312 9875 6338
rect 9931 6312 9983 6338
rect 737 6255 789 6307
rect 845 6255 897 6307
rect 2279 6286 2331 6312
rect 2387 6286 2439 6312
rect 2495 6286 2547 6312
rect 2603 6286 2655 6312
rect 2711 6286 2763 6312
rect 4551 6286 4603 6312
rect 4659 6286 4711 6312
rect 4767 6286 4819 6312
rect 4875 6286 4927 6312
rect 4983 6286 5035 6312
rect 7227 6286 7279 6312
rect 7335 6286 7387 6312
rect 7443 6286 7495 6312
rect 7551 6286 7603 6312
rect 7659 6286 7711 6312
rect 9499 6286 9551 6312
rect 9607 6286 9659 6312
rect 9715 6286 9767 6312
rect 9823 6286 9875 6312
rect 9931 6286 9983 6312
rect 11365 6255 11417 6307
rect 11473 6255 11525 6307
rect 2279 6204 2331 6230
rect 2387 6204 2439 6230
rect 2495 6204 2547 6230
rect 2603 6204 2655 6230
rect 2711 6204 2763 6230
rect 4551 6204 4603 6230
rect 4659 6204 4711 6230
rect 4767 6204 4819 6230
rect 4875 6204 4927 6230
rect 4983 6204 5035 6230
rect 7227 6204 7279 6230
rect 7335 6204 7387 6230
rect 7443 6204 7495 6230
rect 7551 6204 7603 6230
rect 7659 6204 7711 6230
rect 9499 6204 9551 6230
rect 9607 6204 9659 6230
rect 9715 6204 9767 6230
rect 9823 6204 9875 6230
rect 9931 6204 9983 6230
rect 737 6182 789 6199
rect 737 6147 752 6182
rect 752 6147 789 6182
rect 845 6173 897 6199
rect 2279 6178 2331 6204
rect 2387 6178 2439 6204
rect 2495 6178 2547 6204
rect 2603 6178 2655 6204
rect 2711 6178 2763 6204
rect 4551 6178 4603 6204
rect 4659 6178 4711 6204
rect 4767 6178 4819 6204
rect 4875 6178 4927 6204
rect 4983 6178 5035 6204
rect 7227 6178 7279 6204
rect 7335 6178 7387 6204
rect 7443 6178 7495 6204
rect 7551 6178 7603 6204
rect 7659 6178 7711 6204
rect 9499 6178 9551 6204
rect 9607 6178 9659 6204
rect 9715 6178 9767 6204
rect 9823 6178 9875 6204
rect 9931 6178 9983 6204
rect 845 6147 860 6173
rect 860 6147 897 6173
rect 11365 6173 11417 6199
rect 11365 6147 11402 6173
rect 11402 6147 11417 6173
rect 11473 6182 11525 6199
rect 11473 6147 11510 6182
rect 11510 6147 11525 6182
rect 737 6039 752 6091
rect 752 6039 789 6091
rect 845 6039 860 6091
rect 860 6039 897 6091
rect 737 5931 752 5983
rect 752 5931 789 5983
rect 845 5931 860 5983
rect 860 5931 897 5983
rect 737 5823 752 5875
rect 752 5823 789 5875
rect 845 5823 860 5875
rect 860 5823 897 5875
rect 737 5715 752 5767
rect 752 5715 789 5767
rect 845 5715 860 5767
rect 860 5715 897 5767
rect 737 5607 752 5659
rect 752 5607 789 5659
rect 845 5607 860 5659
rect 860 5607 897 5659
rect 737 5499 752 5551
rect 752 5499 789 5551
rect 845 5499 860 5551
rect 860 5499 897 5551
rect 737 5391 752 5443
rect 752 5391 789 5443
rect 845 5391 860 5443
rect 860 5391 897 5443
rect 737 5283 752 5335
rect 752 5283 789 5335
rect 845 5283 860 5335
rect 860 5283 897 5335
rect 737 5175 752 5227
rect 752 5175 789 5227
rect 845 5175 860 5227
rect 860 5175 897 5227
rect 1741 5874 1793 5907
rect 1865 5874 1917 5907
rect 1989 5874 2041 5907
rect 2113 5874 2165 5907
rect 2877 5874 2929 5907
rect 3001 5874 3053 5907
rect 3125 5874 3177 5907
rect 3249 5874 3301 5907
rect 4013 5874 4065 5907
rect 4137 5874 4189 5907
rect 4261 5874 4313 5907
rect 4385 5874 4437 5907
rect 5149 5874 5201 5907
rect 5273 5874 5325 5907
rect 5397 5874 5449 5907
rect 5521 5874 5573 5907
rect 6689 5874 6741 5907
rect 6813 5874 6865 5907
rect 6937 5874 6989 5907
rect 7061 5874 7113 5907
rect 7825 5874 7877 5907
rect 7949 5874 8001 5907
rect 8073 5874 8125 5907
rect 8197 5874 8249 5907
rect 8961 5874 9013 5907
rect 9085 5874 9137 5907
rect 9209 5874 9261 5907
rect 9333 5874 9385 5907
rect 10097 5874 10149 5907
rect 10221 5874 10273 5907
rect 10345 5874 10397 5907
rect 10469 5874 10521 5907
rect 1741 5855 1793 5874
rect 1865 5855 1917 5874
rect 1989 5855 2041 5874
rect 2113 5855 2165 5874
rect 2877 5855 2929 5874
rect 3001 5855 3053 5874
rect 3125 5855 3177 5874
rect 3249 5855 3301 5874
rect 4013 5855 4065 5874
rect 4137 5855 4189 5874
rect 4261 5855 4313 5874
rect 4385 5855 4437 5874
rect 5149 5855 5201 5874
rect 5273 5855 5325 5874
rect 5397 5855 5449 5874
rect 5521 5855 5573 5874
rect 6689 5855 6741 5874
rect 6813 5855 6865 5874
rect 6937 5855 6989 5874
rect 7061 5855 7113 5874
rect 7825 5855 7877 5874
rect 7949 5855 8001 5874
rect 8073 5855 8125 5874
rect 8197 5855 8249 5874
rect 8961 5855 9013 5874
rect 9085 5855 9137 5874
rect 9209 5855 9261 5874
rect 9333 5855 9385 5874
rect 10097 5855 10149 5874
rect 10221 5855 10273 5874
rect 10345 5855 10397 5874
rect 10469 5855 10521 5874
rect 1741 5769 1793 5783
rect 1865 5769 1917 5783
rect 1989 5769 2041 5783
rect 2113 5769 2165 5783
rect 2877 5769 2929 5783
rect 3001 5769 3053 5783
rect 3125 5769 3177 5783
rect 3249 5769 3301 5783
rect 4013 5769 4065 5783
rect 4137 5769 4189 5783
rect 4261 5769 4313 5783
rect 4385 5769 4437 5783
rect 5149 5769 5201 5783
rect 5273 5769 5325 5783
rect 5397 5769 5449 5783
rect 5521 5769 5573 5783
rect 6689 5769 6741 5783
rect 6813 5769 6865 5783
rect 6937 5769 6989 5783
rect 7061 5769 7113 5783
rect 7825 5769 7877 5783
rect 7949 5769 8001 5783
rect 8073 5769 8125 5783
rect 8197 5769 8249 5783
rect 8961 5769 9013 5783
rect 9085 5769 9137 5783
rect 9209 5769 9261 5783
rect 9333 5769 9385 5783
rect 10097 5769 10149 5783
rect 10221 5769 10273 5783
rect 10345 5769 10397 5783
rect 10469 5769 10521 5783
rect 1741 5731 1793 5769
rect 1865 5731 1917 5769
rect 1989 5731 2041 5769
rect 2113 5731 2165 5769
rect 2877 5731 2929 5769
rect 3001 5731 3053 5769
rect 3125 5731 3177 5769
rect 3249 5731 3301 5769
rect 4013 5731 4065 5769
rect 4137 5731 4189 5769
rect 4261 5731 4313 5769
rect 4385 5731 4437 5769
rect 5149 5731 5201 5769
rect 5273 5731 5325 5769
rect 5397 5731 5449 5769
rect 5521 5731 5573 5769
rect 6689 5731 6741 5769
rect 6813 5731 6865 5769
rect 6937 5731 6989 5769
rect 7061 5731 7113 5769
rect 7825 5731 7877 5769
rect 7949 5731 8001 5769
rect 8073 5731 8125 5769
rect 8197 5731 8249 5769
rect 8961 5731 9013 5769
rect 9085 5731 9137 5769
rect 9209 5731 9261 5769
rect 9333 5731 9385 5769
rect 10097 5731 10149 5769
rect 10221 5731 10273 5769
rect 10345 5731 10397 5769
rect 10469 5731 10521 5769
rect 1741 5607 1793 5659
rect 1865 5607 1917 5659
rect 1989 5607 2041 5659
rect 2113 5607 2165 5659
rect 2877 5607 2929 5659
rect 3001 5607 3053 5659
rect 3125 5607 3177 5659
rect 3249 5607 3301 5659
rect 4013 5607 4065 5659
rect 4137 5607 4189 5659
rect 4261 5607 4313 5659
rect 4385 5607 4437 5659
rect 5149 5607 5201 5659
rect 5273 5607 5325 5659
rect 5397 5607 5449 5659
rect 5521 5607 5573 5659
rect 6689 5607 6741 5659
rect 6813 5607 6865 5659
rect 6937 5607 6989 5659
rect 7061 5607 7113 5659
rect 7825 5607 7877 5659
rect 7949 5607 8001 5659
rect 8073 5607 8125 5659
rect 8197 5607 8249 5659
rect 8961 5607 9013 5659
rect 9085 5607 9137 5659
rect 9209 5607 9261 5659
rect 9333 5607 9385 5659
rect 10097 5607 10149 5659
rect 10221 5607 10273 5659
rect 10345 5607 10397 5659
rect 10469 5607 10521 5659
rect 1741 5498 1793 5535
rect 1865 5498 1917 5535
rect 1989 5498 2041 5535
rect 2113 5498 2165 5535
rect 2877 5498 2929 5535
rect 3001 5498 3053 5535
rect 3125 5498 3177 5535
rect 3249 5498 3301 5535
rect 4013 5498 4065 5535
rect 4137 5498 4189 5535
rect 4261 5498 4313 5535
rect 4385 5498 4437 5535
rect 5149 5498 5201 5535
rect 5273 5498 5325 5535
rect 5397 5498 5449 5535
rect 5521 5498 5573 5535
rect 6689 5498 6741 5535
rect 6813 5498 6865 5535
rect 6937 5498 6989 5535
rect 7061 5498 7113 5535
rect 7825 5498 7877 5535
rect 7949 5498 8001 5535
rect 8073 5498 8125 5535
rect 8197 5498 8249 5535
rect 8961 5498 9013 5535
rect 9085 5498 9137 5535
rect 9209 5498 9261 5535
rect 9333 5498 9385 5535
rect 10097 5498 10149 5535
rect 10221 5498 10273 5535
rect 10345 5498 10397 5535
rect 10469 5498 10521 5535
rect 1741 5483 1793 5498
rect 1865 5483 1917 5498
rect 1989 5483 2041 5498
rect 2113 5483 2165 5498
rect 2877 5483 2929 5498
rect 3001 5483 3053 5498
rect 3125 5483 3177 5498
rect 3249 5483 3301 5498
rect 4013 5483 4065 5498
rect 4137 5483 4189 5498
rect 4261 5483 4313 5498
rect 4385 5483 4437 5498
rect 5149 5483 5201 5498
rect 5273 5483 5325 5498
rect 5397 5483 5449 5498
rect 5521 5483 5573 5498
rect 6689 5483 6741 5498
rect 6813 5483 6865 5498
rect 6937 5483 6989 5498
rect 7061 5483 7113 5498
rect 7825 5483 7877 5498
rect 7949 5483 8001 5498
rect 8073 5483 8125 5498
rect 8197 5483 8249 5498
rect 8961 5483 9013 5498
rect 9085 5483 9137 5498
rect 9209 5483 9261 5498
rect 9333 5483 9385 5498
rect 10097 5483 10149 5498
rect 10221 5483 10273 5498
rect 10345 5483 10397 5498
rect 10469 5483 10521 5498
rect 1741 5392 1793 5411
rect 1865 5392 1917 5411
rect 1989 5392 2041 5411
rect 2113 5392 2165 5411
rect 2877 5392 2929 5411
rect 3001 5392 3053 5411
rect 3125 5392 3177 5411
rect 3249 5392 3301 5411
rect 4013 5392 4065 5411
rect 4137 5392 4189 5411
rect 4261 5392 4313 5411
rect 4385 5392 4437 5411
rect 5149 5392 5201 5411
rect 5273 5392 5325 5411
rect 5397 5392 5449 5411
rect 5521 5392 5573 5411
rect 6689 5392 6741 5411
rect 6813 5392 6865 5411
rect 6937 5392 6989 5411
rect 7061 5392 7113 5411
rect 7825 5392 7877 5411
rect 7949 5392 8001 5411
rect 8073 5392 8125 5411
rect 8197 5392 8249 5411
rect 8961 5392 9013 5411
rect 9085 5392 9137 5411
rect 9209 5392 9261 5411
rect 9333 5392 9385 5411
rect 10097 5392 10149 5411
rect 10221 5392 10273 5411
rect 10345 5392 10397 5411
rect 10469 5392 10521 5411
rect 1741 5359 1793 5392
rect 1865 5359 1917 5392
rect 1989 5359 2041 5392
rect 2113 5359 2165 5392
rect 2877 5359 2929 5392
rect 3001 5359 3053 5392
rect 3125 5359 3177 5392
rect 3249 5359 3301 5392
rect 4013 5359 4065 5392
rect 4137 5359 4189 5392
rect 4261 5359 4313 5392
rect 4385 5359 4437 5392
rect 5149 5359 5201 5392
rect 5273 5359 5325 5392
rect 5397 5359 5449 5392
rect 5521 5359 5573 5392
rect 6689 5359 6741 5392
rect 6813 5359 6865 5392
rect 6937 5359 6989 5392
rect 7061 5359 7113 5392
rect 7825 5359 7877 5392
rect 7949 5359 8001 5392
rect 8073 5359 8125 5392
rect 8197 5359 8249 5392
rect 8961 5359 9013 5392
rect 9085 5359 9137 5392
rect 9209 5359 9261 5392
rect 9333 5359 9385 5392
rect 10097 5359 10149 5392
rect 10221 5359 10273 5392
rect 10345 5359 10397 5392
rect 10469 5359 10521 5392
rect 11365 6039 11402 6091
rect 11402 6039 11417 6091
rect 11473 6039 11510 6091
rect 11510 6039 11525 6091
rect 11365 5931 11402 5983
rect 11402 5931 11417 5983
rect 11473 5931 11510 5983
rect 11510 5931 11525 5983
rect 11365 5823 11402 5875
rect 11402 5823 11417 5875
rect 11473 5823 11510 5875
rect 11510 5823 11525 5875
rect 11365 5715 11402 5767
rect 11402 5715 11417 5767
rect 11473 5715 11510 5767
rect 11510 5715 11525 5767
rect 11365 5607 11402 5659
rect 11402 5607 11417 5659
rect 11473 5607 11510 5659
rect 11510 5607 11525 5659
rect 11365 5499 11402 5551
rect 11402 5499 11417 5551
rect 11473 5499 11510 5551
rect 11510 5499 11525 5551
rect 11365 5391 11402 5443
rect 11402 5391 11417 5443
rect 11473 5391 11510 5443
rect 11510 5391 11525 5443
rect 11365 5283 11402 5335
rect 11402 5283 11417 5335
rect 11473 5283 11510 5335
rect 11510 5283 11525 5335
rect 11365 5175 11402 5227
rect 11402 5175 11417 5227
rect 11473 5175 11510 5227
rect 11510 5175 11525 5227
rect 737 5067 752 5119
rect 752 5067 789 5119
rect 845 5093 860 5119
rect 860 5093 897 5119
rect 845 5067 897 5093
rect 11365 5093 11402 5119
rect 11402 5093 11417 5119
rect 11365 5067 11417 5093
rect 11473 5067 11510 5119
rect 11510 5067 11525 5119
rect 2279 5062 2331 5065
rect 2387 5062 2439 5065
rect 2495 5062 2547 5065
rect 2603 5062 2655 5065
rect 2711 5062 2763 5065
rect 4551 5062 4603 5065
rect 4659 5062 4711 5065
rect 4767 5062 4819 5065
rect 4875 5062 4927 5065
rect 4983 5062 5035 5065
rect 7227 5062 7279 5065
rect 7335 5062 7387 5065
rect 7443 5062 7495 5065
rect 7551 5062 7603 5065
rect 7659 5062 7711 5065
rect 9499 5062 9551 5065
rect 9607 5062 9659 5065
rect 9715 5062 9767 5065
rect 9823 5062 9875 5065
rect 9931 5062 9983 5065
rect 2279 5013 2331 5062
rect 2387 5013 2439 5062
rect 2495 5013 2547 5062
rect 2603 5013 2655 5062
rect 2711 5013 2763 5062
rect 4551 5013 4603 5062
rect 4659 5013 4711 5062
rect 4767 5013 4819 5062
rect 4875 5013 4927 5062
rect 4983 5013 5035 5062
rect 7227 5013 7279 5062
rect 7335 5013 7387 5062
rect 7443 5013 7495 5062
rect 7551 5013 7603 5062
rect 7659 5013 7711 5062
rect 9499 5013 9551 5062
rect 9607 5013 9659 5062
rect 9715 5013 9767 5062
rect 9823 5013 9875 5062
rect 9931 5013 9983 5062
rect 737 4959 752 5011
rect 752 4959 789 5011
rect 845 4959 897 5011
rect 11365 4959 11417 5011
rect 11473 4959 11510 5011
rect 11510 4959 11525 5011
rect 2279 4954 2331 4957
rect 2387 4954 2439 4957
rect 2495 4954 2547 4957
rect 2603 4954 2655 4957
rect 2711 4954 2763 4957
rect 4551 4954 4603 4957
rect 4659 4954 4711 4957
rect 4767 4954 4819 4957
rect 4875 4954 4927 4957
rect 4983 4954 5035 4957
rect 7227 4954 7279 4957
rect 7335 4954 7387 4957
rect 7443 4954 7495 4957
rect 7551 4954 7603 4957
rect 7659 4954 7711 4957
rect 9499 4954 9551 4957
rect 9607 4954 9659 4957
rect 9715 4954 9767 4957
rect 9823 4954 9875 4957
rect 9931 4954 9983 4957
rect 2279 4908 2331 4954
rect 2387 4908 2439 4954
rect 2495 4908 2547 4954
rect 2603 4908 2655 4954
rect 2711 4908 2763 4954
rect 4551 4908 4603 4954
rect 4659 4908 4711 4954
rect 4767 4908 4819 4954
rect 4875 4908 4927 4954
rect 4983 4908 5035 4954
rect 7227 4908 7279 4954
rect 7335 4908 7387 4954
rect 7443 4908 7495 4954
rect 7551 4908 7603 4954
rect 7659 4908 7711 4954
rect 9499 4908 9551 4954
rect 9607 4908 9659 4954
rect 9715 4908 9767 4954
rect 9823 4908 9875 4954
rect 9931 4908 9983 4954
rect 2279 4905 2331 4908
rect 2387 4905 2439 4908
rect 2495 4905 2547 4908
rect 2603 4905 2655 4908
rect 2711 4905 2763 4908
rect 4551 4905 4603 4908
rect 4659 4905 4711 4908
rect 4767 4905 4819 4908
rect 4875 4905 4927 4908
rect 4983 4905 5035 4908
rect 7227 4905 7279 4908
rect 7335 4905 7387 4908
rect 7443 4905 7495 4908
rect 7551 4905 7603 4908
rect 7659 4905 7711 4908
rect 9499 4905 9551 4908
rect 9607 4905 9659 4908
rect 9715 4905 9767 4908
rect 9823 4905 9875 4908
rect 9931 4905 9983 4908
rect 737 4851 752 4903
rect 752 4851 789 4903
rect 845 4851 897 4903
rect 11365 4851 11417 4903
rect 11473 4851 11510 4903
rect 11510 4851 11525 4903
rect 2279 4800 2331 4849
rect 2387 4800 2439 4849
rect 2495 4800 2547 4849
rect 2603 4800 2655 4849
rect 2711 4800 2763 4849
rect 4551 4800 4603 4849
rect 4659 4800 4711 4849
rect 4767 4800 4819 4849
rect 4875 4800 4927 4849
rect 4983 4800 5035 4849
rect 7227 4800 7279 4849
rect 7335 4800 7387 4849
rect 7443 4800 7495 4849
rect 7551 4800 7603 4849
rect 7659 4800 7711 4849
rect 9499 4800 9551 4849
rect 9607 4800 9659 4849
rect 9715 4800 9767 4849
rect 9823 4800 9875 4849
rect 9931 4800 9983 4849
rect 2279 4797 2331 4800
rect 2387 4797 2439 4800
rect 2495 4797 2547 4800
rect 2603 4797 2655 4800
rect 2711 4797 2763 4800
rect 4551 4797 4603 4800
rect 4659 4797 4711 4800
rect 4767 4797 4819 4800
rect 4875 4797 4927 4800
rect 4983 4797 5035 4800
rect 7227 4797 7279 4800
rect 7335 4797 7387 4800
rect 7443 4797 7495 4800
rect 7551 4797 7603 4800
rect 7659 4797 7711 4800
rect 9499 4797 9551 4800
rect 9607 4797 9659 4800
rect 9715 4797 9767 4800
rect 9823 4797 9875 4800
rect 9931 4797 9983 4800
rect 737 4743 752 4795
rect 752 4743 789 4795
rect 845 4769 897 4795
rect 845 4743 860 4769
rect 860 4743 897 4769
rect 11365 4769 11417 4795
rect 11365 4743 11402 4769
rect 11402 4743 11417 4769
rect 11473 4743 11510 4795
rect 11510 4743 11525 4795
rect 737 4635 752 4687
rect 752 4635 789 4687
rect 845 4635 860 4687
rect 860 4635 897 4687
rect 737 4527 752 4579
rect 752 4527 789 4579
rect 845 4527 860 4579
rect 860 4527 897 4579
rect 737 4419 752 4471
rect 752 4419 789 4471
rect 845 4419 860 4471
rect 860 4419 897 4471
rect 737 4311 752 4363
rect 752 4311 789 4363
rect 845 4311 860 4363
rect 860 4311 897 4363
rect 737 4203 752 4255
rect 752 4203 789 4255
rect 845 4203 860 4255
rect 860 4203 897 4255
rect 737 4095 752 4147
rect 752 4095 789 4147
rect 845 4095 860 4147
rect 860 4095 897 4147
rect 737 3987 752 4039
rect 752 3987 789 4039
rect 845 3987 860 4039
rect 860 3987 897 4039
rect 737 3879 752 3931
rect 752 3879 789 3931
rect 845 3879 860 3931
rect 860 3879 897 3931
rect 737 3771 752 3823
rect 752 3771 789 3823
rect 845 3771 860 3823
rect 860 3771 897 3823
rect 1741 4470 1793 4503
rect 1865 4470 1917 4503
rect 1989 4470 2041 4503
rect 2113 4470 2165 4503
rect 2877 4470 2929 4503
rect 3001 4470 3053 4503
rect 3125 4470 3177 4503
rect 3249 4470 3301 4503
rect 4013 4470 4065 4503
rect 4137 4470 4189 4503
rect 4261 4470 4313 4503
rect 4385 4470 4437 4503
rect 5149 4470 5201 4503
rect 5273 4470 5325 4503
rect 5397 4470 5449 4503
rect 5521 4470 5573 4503
rect 6689 4470 6741 4503
rect 6813 4470 6865 4503
rect 6937 4470 6989 4503
rect 7061 4470 7113 4503
rect 7825 4470 7877 4503
rect 7949 4470 8001 4503
rect 8073 4470 8125 4503
rect 8197 4470 8249 4503
rect 8961 4470 9013 4503
rect 9085 4470 9137 4503
rect 9209 4470 9261 4503
rect 9333 4470 9385 4503
rect 10097 4470 10149 4503
rect 10221 4470 10273 4503
rect 10345 4470 10397 4503
rect 10469 4470 10521 4503
rect 1741 4451 1793 4470
rect 1865 4451 1917 4470
rect 1989 4451 2041 4470
rect 2113 4451 2165 4470
rect 2877 4451 2929 4470
rect 3001 4451 3053 4470
rect 3125 4451 3177 4470
rect 3249 4451 3301 4470
rect 4013 4451 4065 4470
rect 4137 4451 4189 4470
rect 4261 4451 4313 4470
rect 4385 4451 4437 4470
rect 5149 4451 5201 4470
rect 5273 4451 5325 4470
rect 5397 4451 5449 4470
rect 5521 4451 5573 4470
rect 6689 4451 6741 4470
rect 6813 4451 6865 4470
rect 6937 4451 6989 4470
rect 7061 4451 7113 4470
rect 7825 4451 7877 4470
rect 7949 4451 8001 4470
rect 8073 4451 8125 4470
rect 8197 4451 8249 4470
rect 8961 4451 9013 4470
rect 9085 4451 9137 4470
rect 9209 4451 9261 4470
rect 9333 4451 9385 4470
rect 10097 4451 10149 4470
rect 10221 4451 10273 4470
rect 10345 4451 10397 4470
rect 10469 4451 10521 4470
rect 1741 4365 1793 4379
rect 1865 4365 1917 4379
rect 1989 4365 2041 4379
rect 2113 4365 2165 4379
rect 2877 4365 2929 4379
rect 3001 4365 3053 4379
rect 3125 4365 3177 4379
rect 3249 4365 3301 4379
rect 4013 4365 4065 4379
rect 4137 4365 4189 4379
rect 4261 4365 4313 4379
rect 4385 4365 4437 4379
rect 5149 4365 5201 4379
rect 5273 4365 5325 4379
rect 5397 4365 5449 4379
rect 5521 4365 5573 4379
rect 6689 4365 6741 4379
rect 6813 4365 6865 4379
rect 6937 4365 6989 4379
rect 7061 4365 7113 4379
rect 7825 4365 7877 4379
rect 7949 4365 8001 4379
rect 8073 4365 8125 4379
rect 8197 4365 8249 4379
rect 8961 4365 9013 4379
rect 9085 4365 9137 4379
rect 9209 4365 9261 4379
rect 9333 4365 9385 4379
rect 10097 4365 10149 4379
rect 10221 4365 10273 4379
rect 10345 4365 10397 4379
rect 10469 4365 10521 4379
rect 1741 4327 1793 4365
rect 1865 4327 1917 4365
rect 1989 4327 2041 4365
rect 2113 4327 2165 4365
rect 2877 4327 2929 4365
rect 3001 4327 3053 4365
rect 3125 4327 3177 4365
rect 3249 4327 3301 4365
rect 4013 4327 4065 4365
rect 4137 4327 4189 4365
rect 4261 4327 4313 4365
rect 4385 4327 4437 4365
rect 5149 4327 5201 4365
rect 5273 4327 5325 4365
rect 5397 4327 5449 4365
rect 5521 4327 5573 4365
rect 6689 4327 6741 4365
rect 6813 4327 6865 4365
rect 6937 4327 6989 4365
rect 7061 4327 7113 4365
rect 7825 4327 7877 4365
rect 7949 4327 8001 4365
rect 8073 4327 8125 4365
rect 8197 4327 8249 4365
rect 8961 4327 9013 4365
rect 9085 4327 9137 4365
rect 9209 4327 9261 4365
rect 9333 4327 9385 4365
rect 10097 4327 10149 4365
rect 10221 4327 10273 4365
rect 10345 4327 10397 4365
rect 10469 4327 10521 4365
rect 1741 4203 1793 4255
rect 1865 4203 1917 4255
rect 1989 4203 2041 4255
rect 2113 4203 2165 4255
rect 2877 4203 2929 4255
rect 3001 4203 3053 4255
rect 3125 4203 3177 4255
rect 3249 4203 3301 4255
rect 4013 4203 4065 4255
rect 4137 4203 4189 4255
rect 4261 4203 4313 4255
rect 4385 4203 4437 4255
rect 5149 4203 5201 4255
rect 5273 4203 5325 4255
rect 5397 4203 5449 4255
rect 5521 4203 5573 4255
rect 6689 4203 6741 4255
rect 6813 4203 6865 4255
rect 6937 4203 6989 4255
rect 7061 4203 7113 4255
rect 7825 4203 7877 4255
rect 7949 4203 8001 4255
rect 8073 4203 8125 4255
rect 8197 4203 8249 4255
rect 8961 4203 9013 4255
rect 9085 4203 9137 4255
rect 9209 4203 9261 4255
rect 9333 4203 9385 4255
rect 10097 4203 10149 4255
rect 10221 4203 10273 4255
rect 10345 4203 10397 4255
rect 10469 4203 10521 4255
rect 1741 4094 1793 4131
rect 1865 4094 1917 4131
rect 1989 4094 2041 4131
rect 2113 4094 2165 4131
rect 2877 4094 2929 4131
rect 3001 4094 3053 4131
rect 3125 4094 3177 4131
rect 3249 4094 3301 4131
rect 4013 4094 4065 4131
rect 4137 4094 4189 4131
rect 4261 4094 4313 4131
rect 4385 4094 4437 4131
rect 5149 4094 5201 4131
rect 5273 4094 5325 4131
rect 5397 4094 5449 4131
rect 5521 4094 5573 4131
rect 6689 4094 6741 4131
rect 6813 4094 6865 4131
rect 6937 4094 6989 4131
rect 7061 4094 7113 4131
rect 7825 4094 7877 4131
rect 7949 4094 8001 4131
rect 8073 4094 8125 4131
rect 8197 4094 8249 4131
rect 8961 4094 9013 4131
rect 9085 4094 9137 4131
rect 9209 4094 9261 4131
rect 9333 4094 9385 4131
rect 10097 4094 10149 4131
rect 10221 4094 10273 4131
rect 10345 4094 10397 4131
rect 10469 4094 10521 4131
rect 1741 4079 1793 4094
rect 1865 4079 1917 4094
rect 1989 4079 2041 4094
rect 2113 4079 2165 4094
rect 2877 4079 2929 4094
rect 3001 4079 3053 4094
rect 3125 4079 3177 4094
rect 3249 4079 3301 4094
rect 4013 4079 4065 4094
rect 4137 4079 4189 4094
rect 4261 4079 4313 4094
rect 4385 4079 4437 4094
rect 5149 4079 5201 4094
rect 5273 4079 5325 4094
rect 5397 4079 5449 4094
rect 5521 4079 5573 4094
rect 6689 4079 6741 4094
rect 6813 4079 6865 4094
rect 6937 4079 6989 4094
rect 7061 4079 7113 4094
rect 7825 4079 7877 4094
rect 7949 4079 8001 4094
rect 8073 4079 8125 4094
rect 8197 4079 8249 4094
rect 8961 4079 9013 4094
rect 9085 4079 9137 4094
rect 9209 4079 9261 4094
rect 9333 4079 9385 4094
rect 10097 4079 10149 4094
rect 10221 4079 10273 4094
rect 10345 4079 10397 4094
rect 10469 4079 10521 4094
rect 1741 3988 1793 4007
rect 1865 3988 1917 4007
rect 1989 3988 2041 4007
rect 2113 3988 2165 4007
rect 2877 3988 2929 4007
rect 3001 3988 3053 4007
rect 3125 3988 3177 4007
rect 3249 3988 3301 4007
rect 4013 3988 4065 4007
rect 4137 3988 4189 4007
rect 4261 3988 4313 4007
rect 4385 3988 4437 4007
rect 5149 3988 5201 4007
rect 5273 3988 5325 4007
rect 5397 3988 5449 4007
rect 5521 3988 5573 4007
rect 6689 3988 6741 4007
rect 6813 3988 6865 4007
rect 6937 3988 6989 4007
rect 7061 3988 7113 4007
rect 7825 3988 7877 4007
rect 7949 3988 8001 4007
rect 8073 3988 8125 4007
rect 8197 3988 8249 4007
rect 8961 3988 9013 4007
rect 9085 3988 9137 4007
rect 9209 3988 9261 4007
rect 9333 3988 9385 4007
rect 10097 3988 10149 4007
rect 10221 3988 10273 4007
rect 10345 3988 10397 4007
rect 10469 3988 10521 4007
rect 1741 3955 1793 3988
rect 1865 3955 1917 3988
rect 1989 3955 2041 3988
rect 2113 3955 2165 3988
rect 2877 3955 2929 3988
rect 3001 3955 3053 3988
rect 3125 3955 3177 3988
rect 3249 3955 3301 3988
rect 4013 3955 4065 3988
rect 4137 3955 4189 3988
rect 4261 3955 4313 3988
rect 4385 3955 4437 3988
rect 5149 3955 5201 3988
rect 5273 3955 5325 3988
rect 5397 3955 5449 3988
rect 5521 3955 5573 3988
rect 6689 3955 6741 3988
rect 6813 3955 6865 3988
rect 6937 3955 6989 3988
rect 7061 3955 7113 3988
rect 7825 3955 7877 3988
rect 7949 3955 8001 3988
rect 8073 3955 8125 3988
rect 8197 3955 8249 3988
rect 8961 3955 9013 3988
rect 9085 3955 9137 3988
rect 9209 3955 9261 3988
rect 9333 3955 9385 3988
rect 10097 3955 10149 3988
rect 10221 3955 10273 3988
rect 10345 3955 10397 3988
rect 10469 3955 10521 3988
rect 11365 4635 11402 4687
rect 11402 4635 11417 4687
rect 11473 4635 11510 4687
rect 11510 4635 11525 4687
rect 11365 4527 11402 4579
rect 11402 4527 11417 4579
rect 11473 4527 11510 4579
rect 11510 4527 11525 4579
rect 11365 4419 11402 4471
rect 11402 4419 11417 4471
rect 11473 4419 11510 4471
rect 11510 4419 11525 4471
rect 11365 4311 11402 4363
rect 11402 4311 11417 4363
rect 11473 4311 11510 4363
rect 11510 4311 11525 4363
rect 11365 4203 11402 4255
rect 11402 4203 11417 4255
rect 11473 4203 11510 4255
rect 11510 4203 11525 4255
rect 11365 4095 11402 4147
rect 11402 4095 11417 4147
rect 11473 4095 11510 4147
rect 11510 4095 11525 4147
rect 11365 3987 11402 4039
rect 11402 3987 11417 4039
rect 11473 3987 11510 4039
rect 11510 3987 11525 4039
rect 11365 3879 11402 3931
rect 11402 3879 11417 3931
rect 11473 3879 11510 3931
rect 11510 3879 11525 3931
rect 11365 3771 11402 3823
rect 11402 3771 11417 3823
rect 11473 3771 11510 3823
rect 11510 3771 11525 3823
rect 737 3663 752 3715
rect 752 3663 789 3715
rect 845 3689 860 3715
rect 860 3689 897 3715
rect 845 3663 897 3689
rect 11365 3689 11402 3715
rect 11402 3689 11417 3715
rect 11365 3663 11417 3689
rect 11473 3663 11510 3715
rect 11510 3663 11525 3715
rect 2279 3658 2331 3661
rect 2387 3658 2439 3661
rect 2495 3658 2547 3661
rect 2603 3658 2655 3661
rect 2711 3658 2763 3661
rect 4551 3658 4603 3661
rect 4659 3658 4711 3661
rect 4767 3658 4819 3661
rect 4875 3658 4927 3661
rect 4983 3658 5035 3661
rect 7227 3658 7279 3661
rect 7335 3658 7387 3661
rect 7443 3658 7495 3661
rect 7551 3658 7603 3661
rect 7659 3658 7711 3661
rect 9499 3658 9551 3661
rect 9607 3658 9659 3661
rect 9715 3658 9767 3661
rect 9823 3658 9875 3661
rect 9931 3658 9983 3661
rect 2279 3609 2331 3658
rect 2387 3609 2439 3658
rect 2495 3609 2547 3658
rect 2603 3609 2655 3658
rect 2711 3609 2763 3658
rect 4551 3609 4603 3658
rect 4659 3609 4711 3658
rect 4767 3609 4819 3658
rect 4875 3609 4927 3658
rect 4983 3609 5035 3658
rect 7227 3609 7279 3658
rect 7335 3609 7387 3658
rect 7443 3609 7495 3658
rect 7551 3609 7603 3658
rect 7659 3609 7711 3658
rect 9499 3609 9551 3658
rect 9607 3609 9659 3658
rect 9715 3609 9767 3658
rect 9823 3609 9875 3658
rect 9931 3609 9983 3658
rect 737 3555 752 3607
rect 752 3555 789 3607
rect 845 3555 897 3607
rect 11365 3555 11417 3607
rect 11473 3555 11510 3607
rect 11510 3555 11525 3607
rect 2279 3550 2331 3553
rect 2387 3550 2439 3553
rect 2495 3550 2547 3553
rect 2603 3550 2655 3553
rect 2711 3550 2763 3553
rect 4551 3550 4603 3553
rect 4659 3550 4711 3553
rect 4767 3550 4819 3553
rect 4875 3550 4927 3553
rect 4983 3550 5035 3553
rect 7227 3550 7279 3553
rect 7335 3550 7387 3553
rect 7443 3550 7495 3553
rect 7551 3550 7603 3553
rect 7659 3550 7711 3553
rect 9499 3550 9551 3553
rect 9607 3550 9659 3553
rect 9715 3550 9767 3553
rect 9823 3550 9875 3553
rect 9931 3550 9983 3553
rect 2279 3504 2331 3550
rect 2387 3504 2439 3550
rect 2495 3504 2547 3550
rect 2603 3504 2655 3550
rect 2711 3504 2763 3550
rect 4551 3504 4603 3550
rect 4659 3504 4711 3550
rect 4767 3504 4819 3550
rect 4875 3504 4927 3550
rect 4983 3504 5035 3550
rect 7227 3504 7279 3550
rect 7335 3504 7387 3550
rect 7443 3504 7495 3550
rect 7551 3504 7603 3550
rect 7659 3504 7711 3550
rect 9499 3504 9551 3550
rect 9607 3504 9659 3550
rect 9715 3504 9767 3550
rect 9823 3504 9875 3550
rect 9931 3504 9983 3550
rect 2279 3501 2331 3504
rect 2387 3501 2439 3504
rect 2495 3501 2547 3504
rect 2603 3501 2655 3504
rect 2711 3501 2763 3504
rect 4551 3501 4603 3504
rect 4659 3501 4711 3504
rect 4767 3501 4819 3504
rect 4875 3501 4927 3504
rect 4983 3501 5035 3504
rect 7227 3501 7279 3504
rect 7335 3501 7387 3504
rect 7443 3501 7495 3504
rect 7551 3501 7603 3504
rect 7659 3501 7711 3504
rect 9499 3501 9551 3504
rect 9607 3501 9659 3504
rect 9715 3501 9767 3504
rect 9823 3501 9875 3504
rect 9931 3501 9983 3504
rect 737 3447 752 3499
rect 752 3447 789 3499
rect 845 3447 897 3499
rect 11365 3447 11417 3499
rect 11473 3447 11510 3499
rect 11510 3447 11525 3499
rect 2279 3396 2331 3445
rect 2387 3396 2439 3445
rect 2495 3396 2547 3445
rect 2603 3396 2655 3445
rect 2711 3396 2763 3445
rect 4551 3396 4603 3445
rect 4659 3396 4711 3445
rect 4767 3396 4819 3445
rect 4875 3396 4927 3445
rect 4983 3396 5035 3445
rect 7227 3396 7279 3445
rect 7335 3396 7387 3445
rect 7443 3396 7495 3445
rect 7551 3396 7603 3445
rect 7659 3396 7711 3445
rect 9499 3396 9551 3445
rect 9607 3396 9659 3445
rect 9715 3396 9767 3445
rect 9823 3396 9875 3445
rect 9931 3396 9983 3445
rect 2279 3393 2331 3396
rect 2387 3393 2439 3396
rect 2495 3393 2547 3396
rect 2603 3393 2655 3396
rect 2711 3393 2763 3396
rect 4551 3393 4603 3396
rect 4659 3393 4711 3396
rect 4767 3393 4819 3396
rect 4875 3393 4927 3396
rect 4983 3393 5035 3396
rect 7227 3393 7279 3396
rect 7335 3393 7387 3396
rect 7443 3393 7495 3396
rect 7551 3393 7603 3396
rect 7659 3393 7711 3396
rect 9499 3393 9551 3396
rect 9607 3393 9659 3396
rect 9715 3393 9767 3396
rect 9823 3393 9875 3396
rect 9931 3393 9983 3396
rect 737 3339 752 3391
rect 752 3339 789 3391
rect 845 3365 897 3391
rect 845 3339 860 3365
rect 860 3339 897 3365
rect 11365 3365 11417 3391
rect 11365 3339 11402 3365
rect 11402 3339 11417 3365
rect 11473 3339 11510 3391
rect 11510 3339 11525 3391
rect 737 3231 752 3283
rect 752 3231 789 3283
rect 845 3231 860 3283
rect 860 3231 897 3283
rect 737 3123 752 3175
rect 752 3123 789 3175
rect 845 3123 860 3175
rect 860 3123 897 3175
rect 737 3015 752 3067
rect 752 3015 789 3067
rect 845 3015 860 3067
rect 860 3015 897 3067
rect 737 2907 752 2959
rect 752 2907 789 2959
rect 845 2907 860 2959
rect 860 2907 897 2959
rect 737 2799 752 2851
rect 752 2799 789 2851
rect 845 2799 860 2851
rect 860 2799 897 2851
rect 737 2691 752 2743
rect 752 2691 789 2743
rect 845 2691 860 2743
rect 860 2691 897 2743
rect 737 2583 752 2635
rect 752 2583 789 2635
rect 845 2583 860 2635
rect 860 2583 897 2635
rect 737 2475 752 2527
rect 752 2475 789 2527
rect 845 2475 860 2527
rect 860 2475 897 2527
rect 737 2367 752 2419
rect 752 2367 789 2419
rect 845 2367 860 2419
rect 860 2367 897 2419
rect 1741 3066 1793 3099
rect 1865 3066 1917 3099
rect 1989 3066 2041 3099
rect 2113 3066 2165 3099
rect 2877 3066 2929 3099
rect 3001 3066 3053 3099
rect 3125 3066 3177 3099
rect 3249 3066 3301 3099
rect 4013 3066 4065 3099
rect 4137 3066 4189 3099
rect 4261 3066 4313 3099
rect 4385 3066 4437 3099
rect 5149 3066 5201 3099
rect 5273 3066 5325 3099
rect 5397 3066 5449 3099
rect 5521 3066 5573 3099
rect 6689 3066 6741 3099
rect 6813 3066 6865 3099
rect 6937 3066 6989 3099
rect 7061 3066 7113 3099
rect 7825 3066 7877 3099
rect 7949 3066 8001 3099
rect 8073 3066 8125 3099
rect 8197 3066 8249 3099
rect 8961 3066 9013 3099
rect 9085 3066 9137 3099
rect 9209 3066 9261 3099
rect 9333 3066 9385 3099
rect 10097 3066 10149 3099
rect 10221 3066 10273 3099
rect 10345 3066 10397 3099
rect 10469 3066 10521 3099
rect 1741 3047 1793 3066
rect 1865 3047 1917 3066
rect 1989 3047 2041 3066
rect 2113 3047 2165 3066
rect 2877 3047 2929 3066
rect 3001 3047 3053 3066
rect 3125 3047 3177 3066
rect 3249 3047 3301 3066
rect 4013 3047 4065 3066
rect 4137 3047 4189 3066
rect 4261 3047 4313 3066
rect 4385 3047 4437 3066
rect 5149 3047 5201 3066
rect 5273 3047 5325 3066
rect 5397 3047 5449 3066
rect 5521 3047 5573 3066
rect 6689 3047 6741 3066
rect 6813 3047 6865 3066
rect 6937 3047 6989 3066
rect 7061 3047 7113 3066
rect 7825 3047 7877 3066
rect 7949 3047 8001 3066
rect 8073 3047 8125 3066
rect 8197 3047 8249 3066
rect 8961 3047 9013 3066
rect 9085 3047 9137 3066
rect 9209 3047 9261 3066
rect 9333 3047 9385 3066
rect 10097 3047 10149 3066
rect 10221 3047 10273 3066
rect 10345 3047 10397 3066
rect 10469 3047 10521 3066
rect 1741 2961 1793 2975
rect 1865 2961 1917 2975
rect 1989 2961 2041 2975
rect 2113 2961 2165 2975
rect 2877 2961 2929 2975
rect 3001 2961 3053 2975
rect 3125 2961 3177 2975
rect 3249 2961 3301 2975
rect 4013 2961 4065 2975
rect 4137 2961 4189 2975
rect 4261 2961 4313 2975
rect 4385 2961 4437 2975
rect 5149 2961 5201 2975
rect 5273 2961 5325 2975
rect 5397 2961 5449 2975
rect 5521 2961 5573 2975
rect 6689 2961 6741 2975
rect 6813 2961 6865 2975
rect 6937 2961 6989 2975
rect 7061 2961 7113 2975
rect 7825 2961 7877 2975
rect 7949 2961 8001 2975
rect 8073 2961 8125 2975
rect 8197 2961 8249 2975
rect 8961 2961 9013 2975
rect 9085 2961 9137 2975
rect 9209 2961 9261 2975
rect 9333 2961 9385 2975
rect 10097 2961 10149 2975
rect 10221 2961 10273 2975
rect 10345 2961 10397 2975
rect 10469 2961 10521 2975
rect 1741 2923 1793 2961
rect 1865 2923 1917 2961
rect 1989 2923 2041 2961
rect 2113 2923 2165 2961
rect 2877 2923 2929 2961
rect 3001 2923 3053 2961
rect 3125 2923 3177 2961
rect 3249 2923 3301 2961
rect 4013 2923 4065 2961
rect 4137 2923 4189 2961
rect 4261 2923 4313 2961
rect 4385 2923 4437 2961
rect 5149 2923 5201 2961
rect 5273 2923 5325 2961
rect 5397 2923 5449 2961
rect 5521 2923 5573 2961
rect 6689 2923 6741 2961
rect 6813 2923 6865 2961
rect 6937 2923 6989 2961
rect 7061 2923 7113 2961
rect 7825 2923 7877 2961
rect 7949 2923 8001 2961
rect 8073 2923 8125 2961
rect 8197 2923 8249 2961
rect 8961 2923 9013 2961
rect 9085 2923 9137 2961
rect 9209 2923 9261 2961
rect 9333 2923 9385 2961
rect 10097 2923 10149 2961
rect 10221 2923 10273 2961
rect 10345 2923 10397 2961
rect 10469 2923 10521 2961
rect 1741 2799 1793 2851
rect 1865 2799 1917 2851
rect 1989 2799 2041 2851
rect 2113 2799 2165 2851
rect 2877 2799 2929 2851
rect 3001 2799 3053 2851
rect 3125 2799 3177 2851
rect 3249 2799 3301 2851
rect 4013 2799 4065 2851
rect 4137 2799 4189 2851
rect 4261 2799 4313 2851
rect 4385 2799 4437 2851
rect 5149 2799 5201 2851
rect 5273 2799 5325 2851
rect 5397 2799 5449 2851
rect 5521 2799 5573 2851
rect 6689 2799 6741 2851
rect 6813 2799 6865 2851
rect 6937 2799 6989 2851
rect 7061 2799 7113 2851
rect 7825 2799 7877 2851
rect 7949 2799 8001 2851
rect 8073 2799 8125 2851
rect 8197 2799 8249 2851
rect 8961 2799 9013 2851
rect 9085 2799 9137 2851
rect 9209 2799 9261 2851
rect 9333 2799 9385 2851
rect 10097 2799 10149 2851
rect 10221 2799 10273 2851
rect 10345 2799 10397 2851
rect 10469 2799 10521 2851
rect 1741 2690 1793 2727
rect 1865 2690 1917 2727
rect 1989 2690 2041 2727
rect 2113 2690 2165 2727
rect 2877 2690 2929 2727
rect 3001 2690 3053 2727
rect 3125 2690 3177 2727
rect 3249 2690 3301 2727
rect 4013 2690 4065 2727
rect 4137 2690 4189 2727
rect 4261 2690 4313 2727
rect 4385 2690 4437 2727
rect 5149 2690 5201 2727
rect 5273 2690 5325 2727
rect 5397 2690 5449 2727
rect 5521 2690 5573 2727
rect 6689 2690 6741 2727
rect 6813 2690 6865 2727
rect 6937 2690 6989 2727
rect 7061 2690 7113 2727
rect 7825 2690 7877 2727
rect 7949 2690 8001 2727
rect 8073 2690 8125 2727
rect 8197 2690 8249 2727
rect 8961 2690 9013 2727
rect 9085 2690 9137 2727
rect 9209 2690 9261 2727
rect 9333 2690 9385 2727
rect 10097 2690 10149 2727
rect 10221 2690 10273 2727
rect 10345 2690 10397 2727
rect 10469 2690 10521 2727
rect 1741 2675 1793 2690
rect 1865 2675 1917 2690
rect 1989 2675 2041 2690
rect 2113 2675 2165 2690
rect 2877 2675 2929 2690
rect 3001 2675 3053 2690
rect 3125 2675 3177 2690
rect 3249 2675 3301 2690
rect 4013 2675 4065 2690
rect 4137 2675 4189 2690
rect 4261 2675 4313 2690
rect 4385 2675 4437 2690
rect 5149 2675 5201 2690
rect 5273 2675 5325 2690
rect 5397 2675 5449 2690
rect 5521 2675 5573 2690
rect 6689 2675 6741 2690
rect 6813 2675 6865 2690
rect 6937 2675 6989 2690
rect 7061 2675 7113 2690
rect 7825 2675 7877 2690
rect 7949 2675 8001 2690
rect 8073 2675 8125 2690
rect 8197 2675 8249 2690
rect 8961 2675 9013 2690
rect 9085 2675 9137 2690
rect 9209 2675 9261 2690
rect 9333 2675 9385 2690
rect 10097 2675 10149 2690
rect 10221 2675 10273 2690
rect 10345 2675 10397 2690
rect 10469 2675 10521 2690
rect 1741 2584 1793 2603
rect 1865 2584 1917 2603
rect 1989 2584 2041 2603
rect 2113 2584 2165 2603
rect 2877 2584 2929 2603
rect 3001 2584 3053 2603
rect 3125 2584 3177 2603
rect 3249 2584 3301 2603
rect 4013 2584 4065 2603
rect 4137 2584 4189 2603
rect 4261 2584 4313 2603
rect 4385 2584 4437 2603
rect 5149 2584 5201 2603
rect 5273 2584 5325 2603
rect 5397 2584 5449 2603
rect 5521 2584 5573 2603
rect 6689 2584 6741 2603
rect 6813 2584 6865 2603
rect 6937 2584 6989 2603
rect 7061 2584 7113 2603
rect 7825 2584 7877 2603
rect 7949 2584 8001 2603
rect 8073 2584 8125 2603
rect 8197 2584 8249 2603
rect 8961 2584 9013 2603
rect 9085 2584 9137 2603
rect 9209 2584 9261 2603
rect 9333 2584 9385 2603
rect 10097 2584 10149 2603
rect 10221 2584 10273 2603
rect 10345 2584 10397 2603
rect 10469 2584 10521 2603
rect 1741 2551 1793 2584
rect 1865 2551 1917 2584
rect 1989 2551 2041 2584
rect 2113 2551 2165 2584
rect 2877 2551 2929 2584
rect 3001 2551 3053 2584
rect 3125 2551 3177 2584
rect 3249 2551 3301 2584
rect 4013 2551 4065 2584
rect 4137 2551 4189 2584
rect 4261 2551 4313 2584
rect 4385 2551 4437 2584
rect 5149 2551 5201 2584
rect 5273 2551 5325 2584
rect 5397 2551 5449 2584
rect 5521 2551 5573 2584
rect 6689 2551 6741 2584
rect 6813 2551 6865 2584
rect 6937 2551 6989 2584
rect 7061 2551 7113 2584
rect 7825 2551 7877 2584
rect 7949 2551 8001 2584
rect 8073 2551 8125 2584
rect 8197 2551 8249 2584
rect 8961 2551 9013 2584
rect 9085 2551 9137 2584
rect 9209 2551 9261 2584
rect 9333 2551 9385 2584
rect 10097 2551 10149 2584
rect 10221 2551 10273 2584
rect 10345 2551 10397 2584
rect 10469 2551 10521 2584
rect 11365 3231 11402 3283
rect 11402 3231 11417 3283
rect 11473 3231 11510 3283
rect 11510 3231 11525 3283
rect 11365 3123 11402 3175
rect 11402 3123 11417 3175
rect 11473 3123 11510 3175
rect 11510 3123 11525 3175
rect 11365 3015 11402 3067
rect 11402 3015 11417 3067
rect 11473 3015 11510 3067
rect 11510 3015 11525 3067
rect 11365 2907 11402 2959
rect 11402 2907 11417 2959
rect 11473 2907 11510 2959
rect 11510 2907 11525 2959
rect 11365 2799 11402 2851
rect 11402 2799 11417 2851
rect 11473 2799 11510 2851
rect 11510 2799 11525 2851
rect 11365 2691 11402 2743
rect 11402 2691 11417 2743
rect 11473 2691 11510 2743
rect 11510 2691 11525 2743
rect 11365 2583 11402 2635
rect 11402 2583 11417 2635
rect 11473 2583 11510 2635
rect 11510 2583 11525 2635
rect 11365 2475 11402 2527
rect 11402 2475 11417 2527
rect 11473 2475 11510 2527
rect 11510 2475 11525 2527
rect 11365 2367 11402 2419
rect 11402 2367 11417 2419
rect 11473 2367 11510 2419
rect 11510 2367 11525 2419
rect 737 2259 752 2311
rect 752 2259 789 2311
rect 845 2285 860 2311
rect 860 2285 897 2311
rect 845 2259 897 2285
rect 11365 2285 11402 2311
rect 11402 2285 11417 2311
rect 11365 2259 11417 2285
rect 11473 2259 11510 2311
rect 11510 2259 11525 2311
rect 2279 2254 2331 2257
rect 2387 2254 2439 2257
rect 2495 2254 2547 2257
rect 2603 2254 2655 2257
rect 2711 2254 2763 2257
rect 4551 2254 4603 2257
rect 4659 2254 4711 2257
rect 4767 2254 4819 2257
rect 4875 2254 4927 2257
rect 4983 2254 5035 2257
rect 7227 2254 7279 2257
rect 7335 2254 7387 2257
rect 7443 2254 7495 2257
rect 7551 2254 7603 2257
rect 7659 2254 7711 2257
rect 9499 2254 9551 2257
rect 9607 2254 9659 2257
rect 9715 2254 9767 2257
rect 9823 2254 9875 2257
rect 9931 2254 9983 2257
rect 2279 2205 2331 2254
rect 2387 2205 2439 2254
rect 2495 2205 2547 2254
rect 2603 2205 2655 2254
rect 2711 2205 2763 2254
rect 4551 2205 4603 2254
rect 4659 2205 4711 2254
rect 4767 2205 4819 2254
rect 4875 2205 4927 2254
rect 4983 2205 5035 2254
rect 7227 2205 7279 2254
rect 7335 2205 7387 2254
rect 7443 2205 7495 2254
rect 7551 2205 7603 2254
rect 7659 2205 7711 2254
rect 9499 2205 9551 2254
rect 9607 2205 9659 2254
rect 9715 2205 9767 2254
rect 9823 2205 9875 2254
rect 9931 2205 9983 2254
rect 737 2151 752 2203
rect 752 2151 789 2203
rect 845 2151 897 2203
rect 11365 2151 11417 2203
rect 11473 2151 11510 2203
rect 11510 2151 11525 2203
rect 2279 2146 2331 2149
rect 2387 2146 2439 2149
rect 2495 2146 2547 2149
rect 2603 2146 2655 2149
rect 2711 2146 2763 2149
rect 4551 2146 4603 2149
rect 4659 2146 4711 2149
rect 4767 2146 4819 2149
rect 4875 2146 4927 2149
rect 4983 2146 5035 2149
rect 7227 2146 7279 2149
rect 7335 2146 7387 2149
rect 7443 2146 7495 2149
rect 7551 2146 7603 2149
rect 7659 2146 7711 2149
rect 9499 2146 9551 2149
rect 9607 2146 9659 2149
rect 9715 2146 9767 2149
rect 9823 2146 9875 2149
rect 9931 2146 9983 2149
rect 2279 2100 2331 2146
rect 2387 2100 2439 2146
rect 2495 2100 2547 2146
rect 2603 2100 2655 2146
rect 2711 2100 2763 2146
rect 4551 2100 4603 2146
rect 4659 2100 4711 2146
rect 4767 2100 4819 2146
rect 4875 2100 4927 2146
rect 4983 2100 5035 2146
rect 7227 2100 7279 2146
rect 7335 2100 7387 2146
rect 7443 2100 7495 2146
rect 7551 2100 7603 2146
rect 7659 2100 7711 2146
rect 9499 2100 9551 2146
rect 9607 2100 9659 2146
rect 9715 2100 9767 2146
rect 9823 2100 9875 2146
rect 9931 2100 9983 2146
rect 2279 2097 2331 2100
rect 2387 2097 2439 2100
rect 2495 2097 2547 2100
rect 2603 2097 2655 2100
rect 2711 2097 2763 2100
rect 4551 2097 4603 2100
rect 4659 2097 4711 2100
rect 4767 2097 4819 2100
rect 4875 2097 4927 2100
rect 4983 2097 5035 2100
rect 7227 2097 7279 2100
rect 7335 2097 7387 2100
rect 7443 2097 7495 2100
rect 7551 2097 7603 2100
rect 7659 2097 7711 2100
rect 9499 2097 9551 2100
rect 9607 2097 9659 2100
rect 9715 2097 9767 2100
rect 9823 2097 9875 2100
rect 9931 2097 9983 2100
rect 737 2043 752 2095
rect 752 2043 789 2095
rect 845 2043 897 2095
rect 11365 2043 11417 2095
rect 11473 2043 11510 2095
rect 11510 2043 11525 2095
rect 2279 1992 2331 2041
rect 2387 1992 2439 2041
rect 2495 1992 2547 2041
rect 2603 1992 2655 2041
rect 2711 1992 2763 2041
rect 4551 1992 4603 2041
rect 4659 1992 4711 2041
rect 4767 1992 4819 2041
rect 4875 1992 4927 2041
rect 4983 1992 5035 2041
rect 7227 1992 7279 2041
rect 7335 1992 7387 2041
rect 7443 1992 7495 2041
rect 7551 1992 7603 2041
rect 7659 1992 7711 2041
rect 9499 1992 9551 2041
rect 9607 1992 9659 2041
rect 9715 1992 9767 2041
rect 9823 1992 9875 2041
rect 9931 1992 9983 2041
rect 2279 1989 2331 1992
rect 2387 1989 2439 1992
rect 2495 1989 2547 1992
rect 2603 1989 2655 1992
rect 2711 1989 2763 1992
rect 4551 1989 4603 1992
rect 4659 1989 4711 1992
rect 4767 1989 4819 1992
rect 4875 1989 4927 1992
rect 4983 1989 5035 1992
rect 7227 1989 7279 1992
rect 7335 1989 7387 1992
rect 7443 1989 7495 1992
rect 7551 1989 7603 1992
rect 7659 1989 7711 1992
rect 9499 1989 9551 1992
rect 9607 1989 9659 1992
rect 9715 1989 9767 1992
rect 9823 1989 9875 1992
rect 9931 1989 9983 1992
rect 737 1935 752 1987
rect 752 1935 789 1987
rect 845 1961 897 1987
rect 845 1935 860 1961
rect 860 1935 897 1961
rect 11365 1961 11417 1987
rect 11365 1935 11402 1961
rect 11402 1935 11417 1961
rect 11473 1935 11510 1987
rect 11510 1935 11525 1987
rect 737 1827 752 1879
rect 752 1827 789 1879
rect 845 1827 860 1879
rect 860 1827 897 1879
rect 737 1719 752 1771
rect 752 1719 789 1771
rect 845 1719 860 1771
rect 860 1719 897 1771
rect 737 1611 752 1663
rect 752 1611 789 1663
rect 845 1611 860 1663
rect 860 1611 897 1663
rect 737 1503 752 1555
rect 752 1503 789 1555
rect 845 1503 860 1555
rect 860 1503 897 1555
rect 737 1395 752 1447
rect 752 1395 789 1447
rect 845 1395 860 1447
rect 860 1395 897 1447
rect 737 1287 752 1339
rect 752 1287 789 1339
rect 845 1287 860 1339
rect 860 1287 897 1339
rect 737 1179 752 1231
rect 752 1179 789 1231
rect 845 1179 860 1231
rect 860 1179 897 1231
rect 737 1071 752 1123
rect 752 1071 789 1123
rect 845 1071 860 1123
rect 860 1071 897 1123
rect 737 963 752 1015
rect 752 963 789 1015
rect 845 963 860 1015
rect 860 963 897 1015
rect 1741 1662 1793 1695
rect 1865 1662 1917 1695
rect 1989 1662 2041 1695
rect 2113 1662 2165 1695
rect 2877 1662 2929 1695
rect 3001 1662 3053 1695
rect 3125 1662 3177 1695
rect 3249 1662 3301 1695
rect 4013 1662 4065 1695
rect 4137 1662 4189 1695
rect 4261 1662 4313 1695
rect 4385 1662 4437 1695
rect 5149 1662 5201 1695
rect 5273 1662 5325 1695
rect 5397 1662 5449 1695
rect 5521 1662 5573 1695
rect 6689 1662 6741 1695
rect 6813 1662 6865 1695
rect 6937 1662 6989 1695
rect 7061 1662 7113 1695
rect 7825 1662 7877 1695
rect 7949 1662 8001 1695
rect 8073 1662 8125 1695
rect 8197 1662 8249 1695
rect 8961 1662 9013 1695
rect 9085 1662 9137 1695
rect 9209 1662 9261 1695
rect 9333 1662 9385 1695
rect 10097 1662 10149 1695
rect 10221 1662 10273 1695
rect 10345 1662 10397 1695
rect 10469 1662 10521 1695
rect 1741 1643 1793 1662
rect 1865 1643 1917 1662
rect 1989 1643 2041 1662
rect 2113 1643 2165 1662
rect 2877 1643 2929 1662
rect 3001 1643 3053 1662
rect 3125 1643 3177 1662
rect 3249 1643 3301 1662
rect 4013 1643 4065 1662
rect 4137 1643 4189 1662
rect 4261 1643 4313 1662
rect 4385 1643 4437 1662
rect 5149 1643 5201 1662
rect 5273 1643 5325 1662
rect 5397 1643 5449 1662
rect 5521 1643 5573 1662
rect 6689 1643 6741 1662
rect 6813 1643 6865 1662
rect 6937 1643 6989 1662
rect 7061 1643 7113 1662
rect 7825 1643 7877 1662
rect 7949 1643 8001 1662
rect 8073 1643 8125 1662
rect 8197 1643 8249 1662
rect 8961 1643 9013 1662
rect 9085 1643 9137 1662
rect 9209 1643 9261 1662
rect 9333 1643 9385 1662
rect 10097 1643 10149 1662
rect 10221 1643 10273 1662
rect 10345 1643 10397 1662
rect 10469 1643 10521 1662
rect 1741 1557 1793 1571
rect 1865 1557 1917 1571
rect 1989 1557 2041 1571
rect 2113 1557 2165 1571
rect 2877 1557 2929 1571
rect 3001 1557 3053 1571
rect 3125 1557 3177 1571
rect 3249 1557 3301 1571
rect 4013 1557 4065 1571
rect 4137 1557 4189 1571
rect 4261 1557 4313 1571
rect 4385 1557 4437 1571
rect 5149 1557 5201 1571
rect 5273 1557 5325 1571
rect 5397 1557 5449 1571
rect 5521 1557 5573 1571
rect 6689 1557 6741 1571
rect 6813 1557 6865 1571
rect 6937 1557 6989 1571
rect 7061 1557 7113 1571
rect 7825 1557 7877 1571
rect 7949 1557 8001 1571
rect 8073 1557 8125 1571
rect 8197 1557 8249 1571
rect 8961 1557 9013 1571
rect 9085 1557 9137 1571
rect 9209 1557 9261 1571
rect 9333 1557 9385 1571
rect 10097 1557 10149 1571
rect 10221 1557 10273 1571
rect 10345 1557 10397 1571
rect 10469 1557 10521 1571
rect 1741 1519 1793 1557
rect 1865 1519 1917 1557
rect 1989 1519 2041 1557
rect 2113 1519 2165 1557
rect 2877 1519 2929 1557
rect 3001 1519 3053 1557
rect 3125 1519 3177 1557
rect 3249 1519 3301 1557
rect 4013 1519 4065 1557
rect 4137 1519 4189 1557
rect 4261 1519 4313 1557
rect 4385 1519 4437 1557
rect 5149 1519 5201 1557
rect 5273 1519 5325 1557
rect 5397 1519 5449 1557
rect 5521 1519 5573 1557
rect 6689 1519 6741 1557
rect 6813 1519 6865 1557
rect 6937 1519 6989 1557
rect 7061 1519 7113 1557
rect 7825 1519 7877 1557
rect 7949 1519 8001 1557
rect 8073 1519 8125 1557
rect 8197 1519 8249 1557
rect 8961 1519 9013 1557
rect 9085 1519 9137 1557
rect 9209 1519 9261 1557
rect 9333 1519 9385 1557
rect 10097 1519 10149 1557
rect 10221 1519 10273 1557
rect 10345 1519 10397 1557
rect 10469 1519 10521 1557
rect 1741 1395 1793 1447
rect 1865 1395 1917 1447
rect 1989 1395 2041 1447
rect 2113 1395 2165 1447
rect 2877 1395 2929 1447
rect 3001 1395 3053 1447
rect 3125 1395 3177 1447
rect 3249 1395 3301 1447
rect 4013 1395 4065 1447
rect 4137 1395 4189 1447
rect 4261 1395 4313 1447
rect 4385 1395 4437 1447
rect 5149 1395 5201 1447
rect 5273 1395 5325 1447
rect 5397 1395 5449 1447
rect 5521 1395 5573 1447
rect 6689 1395 6741 1447
rect 6813 1395 6865 1447
rect 6937 1395 6989 1447
rect 7061 1395 7113 1447
rect 7825 1395 7877 1447
rect 7949 1395 8001 1447
rect 8073 1395 8125 1447
rect 8197 1395 8249 1447
rect 8961 1395 9013 1447
rect 9085 1395 9137 1447
rect 9209 1395 9261 1447
rect 9333 1395 9385 1447
rect 10097 1395 10149 1447
rect 10221 1395 10273 1447
rect 10345 1395 10397 1447
rect 10469 1395 10521 1447
rect 1741 1286 1793 1323
rect 1865 1286 1917 1323
rect 1989 1286 2041 1323
rect 2113 1286 2165 1323
rect 2877 1286 2929 1323
rect 3001 1286 3053 1323
rect 3125 1286 3177 1323
rect 3249 1286 3301 1323
rect 4013 1286 4065 1323
rect 4137 1286 4189 1323
rect 4261 1286 4313 1323
rect 4385 1286 4437 1323
rect 5149 1286 5201 1323
rect 5273 1286 5325 1323
rect 5397 1286 5449 1323
rect 5521 1286 5573 1323
rect 6689 1286 6741 1323
rect 6813 1286 6865 1323
rect 6937 1286 6989 1323
rect 7061 1286 7113 1323
rect 7825 1286 7877 1323
rect 7949 1286 8001 1323
rect 8073 1286 8125 1323
rect 8197 1286 8249 1323
rect 8961 1286 9013 1323
rect 9085 1286 9137 1323
rect 9209 1286 9261 1323
rect 9333 1286 9385 1323
rect 10097 1286 10149 1323
rect 10221 1286 10273 1323
rect 10345 1286 10397 1323
rect 10469 1286 10521 1323
rect 1741 1271 1793 1286
rect 1865 1271 1917 1286
rect 1989 1271 2041 1286
rect 2113 1271 2165 1286
rect 2877 1271 2929 1286
rect 3001 1271 3053 1286
rect 3125 1271 3177 1286
rect 3249 1271 3301 1286
rect 4013 1271 4065 1286
rect 4137 1271 4189 1286
rect 4261 1271 4313 1286
rect 4385 1271 4437 1286
rect 5149 1271 5201 1286
rect 5273 1271 5325 1286
rect 5397 1271 5449 1286
rect 5521 1271 5573 1286
rect 6689 1271 6741 1286
rect 6813 1271 6865 1286
rect 6937 1271 6989 1286
rect 7061 1271 7113 1286
rect 7825 1271 7877 1286
rect 7949 1271 8001 1286
rect 8073 1271 8125 1286
rect 8197 1271 8249 1286
rect 8961 1271 9013 1286
rect 9085 1271 9137 1286
rect 9209 1271 9261 1286
rect 9333 1271 9385 1286
rect 10097 1271 10149 1286
rect 10221 1271 10273 1286
rect 10345 1271 10397 1286
rect 10469 1271 10521 1286
rect 1741 1180 1793 1199
rect 1865 1180 1917 1199
rect 1989 1180 2041 1199
rect 2113 1180 2165 1199
rect 2877 1180 2929 1199
rect 3001 1180 3053 1199
rect 3125 1180 3177 1199
rect 3249 1180 3301 1199
rect 4013 1180 4065 1199
rect 4137 1180 4189 1199
rect 4261 1180 4313 1199
rect 4385 1180 4437 1199
rect 5149 1180 5201 1199
rect 5273 1180 5325 1199
rect 5397 1180 5449 1199
rect 5521 1180 5573 1199
rect 6689 1180 6741 1199
rect 6813 1180 6865 1199
rect 6937 1180 6989 1199
rect 7061 1180 7113 1199
rect 7825 1180 7877 1199
rect 7949 1180 8001 1199
rect 8073 1180 8125 1199
rect 8197 1180 8249 1199
rect 8961 1180 9013 1199
rect 9085 1180 9137 1199
rect 9209 1180 9261 1199
rect 9333 1180 9385 1199
rect 10097 1180 10149 1199
rect 10221 1180 10273 1199
rect 10345 1180 10397 1199
rect 10469 1180 10521 1199
rect 1741 1147 1793 1180
rect 1865 1147 1917 1180
rect 1989 1147 2041 1180
rect 2113 1147 2165 1180
rect 2877 1147 2929 1180
rect 3001 1147 3053 1180
rect 3125 1147 3177 1180
rect 3249 1147 3301 1180
rect 4013 1147 4065 1180
rect 4137 1147 4189 1180
rect 4261 1147 4313 1180
rect 4385 1147 4437 1180
rect 5149 1147 5201 1180
rect 5273 1147 5325 1180
rect 5397 1147 5449 1180
rect 5521 1147 5573 1180
rect 6689 1147 6741 1180
rect 6813 1147 6865 1180
rect 6937 1147 6989 1180
rect 7061 1147 7113 1180
rect 7825 1147 7877 1180
rect 7949 1147 8001 1180
rect 8073 1147 8125 1180
rect 8197 1147 8249 1180
rect 8961 1147 9013 1180
rect 9085 1147 9137 1180
rect 9209 1147 9261 1180
rect 9333 1147 9385 1180
rect 10097 1147 10149 1180
rect 10221 1147 10273 1180
rect 10345 1147 10397 1180
rect 10469 1147 10521 1180
rect 11365 1827 11402 1879
rect 11402 1827 11417 1879
rect 11473 1827 11510 1879
rect 11510 1827 11525 1879
rect 11365 1719 11402 1771
rect 11402 1719 11417 1771
rect 11473 1719 11510 1771
rect 11510 1719 11525 1771
rect 11365 1611 11402 1663
rect 11402 1611 11417 1663
rect 11473 1611 11510 1663
rect 11510 1611 11525 1663
rect 11365 1503 11402 1555
rect 11402 1503 11417 1555
rect 11473 1503 11510 1555
rect 11510 1503 11525 1555
rect 11365 1395 11402 1447
rect 11402 1395 11417 1447
rect 11473 1395 11510 1447
rect 11510 1395 11525 1447
rect 11365 1287 11402 1339
rect 11402 1287 11417 1339
rect 11473 1287 11510 1339
rect 11510 1287 11525 1339
rect 11365 1179 11402 1231
rect 11402 1179 11417 1231
rect 11473 1179 11510 1231
rect 11510 1179 11525 1231
rect 11365 1071 11402 1123
rect 11402 1071 11417 1123
rect 11473 1071 11510 1123
rect 11510 1071 11525 1123
rect 11365 963 11402 1015
rect 11402 963 11417 1015
rect 11473 963 11510 1015
rect 11510 963 11525 1015
rect 737 872 752 907
rect 752 872 789 907
rect 737 855 789 872
rect 845 881 860 907
rect 860 881 897 907
rect 845 855 897 881
rect 11365 881 11402 907
rect 11402 881 11417 907
rect 2279 850 2331 876
rect 2387 850 2439 876
rect 2495 850 2547 876
rect 2603 850 2655 876
rect 2711 850 2763 876
rect 4551 850 4603 876
rect 4659 850 4711 876
rect 4767 850 4819 876
rect 4875 850 4927 876
rect 4983 850 5035 876
rect 7227 850 7279 876
rect 7335 850 7387 876
rect 7443 850 7495 876
rect 7551 850 7603 876
rect 7659 850 7711 876
rect 9499 850 9551 876
rect 9607 850 9659 876
rect 9715 850 9767 876
rect 9823 850 9875 876
rect 9931 850 9983 876
rect 11365 855 11417 881
rect 11473 872 11510 907
rect 11510 872 11525 907
rect 11473 855 11525 872
rect 2279 824 2331 850
rect 2387 824 2439 850
rect 2495 824 2547 850
rect 2603 824 2655 850
rect 2711 824 2763 850
rect 4551 824 4603 850
rect 4659 824 4711 850
rect 4767 824 4819 850
rect 4875 824 4927 850
rect 4983 824 5035 850
rect 7227 824 7279 850
rect 7335 824 7387 850
rect 7443 824 7495 850
rect 7551 824 7603 850
rect 7659 824 7711 850
rect 9499 824 9551 850
rect 9607 824 9659 850
rect 9715 824 9767 850
rect 9823 824 9875 850
rect 9931 824 9983 850
rect 737 747 789 799
rect 845 747 897 799
rect 2279 742 2331 768
rect 2387 742 2439 768
rect 2495 742 2547 768
rect 2603 742 2655 768
rect 2711 742 2763 768
rect 4551 742 4603 768
rect 4659 742 4711 768
rect 4767 742 4819 768
rect 4875 742 4927 768
rect 4983 742 5035 768
rect 7227 742 7279 768
rect 7335 742 7387 768
rect 7443 742 7495 768
rect 7551 742 7603 768
rect 7659 742 7711 768
rect 9499 742 9551 768
rect 9607 742 9659 768
rect 9715 742 9767 768
rect 9823 742 9875 768
rect 9931 742 9983 768
rect 11365 747 11417 799
rect 11473 747 11525 799
rect 2279 716 2331 742
rect 2387 716 2439 742
rect 2495 716 2547 742
rect 2603 716 2655 742
rect 2711 716 2763 742
rect 4551 716 4603 742
rect 4659 716 4711 742
rect 4767 716 4819 742
rect 4875 716 4927 742
rect 4983 716 5035 742
rect 7227 716 7279 742
rect 7335 716 7387 742
rect 7443 716 7495 742
rect 7551 716 7603 742
rect 7659 716 7711 742
rect 9499 716 9551 742
rect 9607 716 9659 742
rect 9715 716 9767 742
rect 9823 716 9875 742
rect 9931 716 9983 742
rect 11805 6471 11857 6523
rect 11913 6471 11965 6523
rect 12021 6471 12073 6523
rect 11805 6363 11857 6415
rect 11913 6363 11965 6415
rect 12021 6363 12073 6415
rect 11805 6255 11857 6307
rect 11913 6255 11965 6307
rect 12021 6255 12073 6307
rect 11805 6147 11857 6199
rect 11913 6147 11965 6199
rect 12021 6147 12073 6199
rect 11805 6039 11857 6091
rect 11913 6039 11965 6091
rect 12021 6039 12073 6091
rect 11805 5931 11857 5983
rect 11913 5931 11965 5983
rect 12021 5931 12073 5983
rect 11805 5823 11857 5875
rect 11913 5823 11965 5875
rect 12021 5823 12073 5875
rect 11805 5715 11857 5767
rect 11913 5715 11965 5767
rect 12021 5715 12073 5767
rect 11805 5607 11857 5659
rect 11913 5607 11965 5659
rect 12021 5607 12073 5659
rect 11805 5499 11857 5551
rect 11913 5499 11965 5551
rect 12021 5499 12073 5551
rect 11805 5391 11857 5443
rect 11913 5391 11965 5443
rect 12021 5391 12073 5443
rect 11805 5283 11857 5335
rect 11913 5283 11965 5335
rect 12021 5283 12073 5335
rect 11805 5175 11857 5227
rect 11913 5175 11965 5227
rect 12021 5175 12073 5227
rect 11805 5067 11857 5119
rect 11913 5067 11965 5119
rect 12021 5067 12073 5119
rect 11805 4959 11857 5011
rect 11913 4959 11965 5011
rect 12021 4959 12073 5011
rect 11805 4851 11857 4903
rect 11913 4851 11965 4903
rect 12021 4851 12073 4903
rect 11805 4743 11857 4795
rect 11913 4743 11965 4795
rect 12021 4743 12073 4795
rect 11805 4635 11857 4687
rect 11913 4635 11965 4687
rect 12021 4635 12073 4687
rect 11805 4527 11857 4579
rect 11913 4527 11965 4579
rect 12021 4527 12073 4579
rect 11805 4419 11857 4471
rect 11913 4419 11965 4471
rect 12021 4419 12073 4471
rect 11805 4311 11857 4363
rect 11913 4311 11965 4363
rect 12021 4311 12073 4363
rect 11805 4203 11857 4255
rect 11913 4203 11965 4255
rect 12021 4203 12073 4255
rect 11805 4095 11857 4147
rect 11913 4095 11965 4147
rect 12021 4095 12073 4147
rect 11805 3987 11857 4039
rect 11913 3987 11965 4039
rect 12021 3987 12073 4039
rect 11805 3879 11857 3931
rect 11913 3879 11965 3931
rect 12021 3879 12073 3931
rect 11805 3771 11857 3823
rect 11913 3771 11965 3823
rect 12021 3771 12073 3823
rect 11805 3663 11857 3715
rect 11913 3663 11965 3715
rect 12021 3663 12073 3715
rect 11805 3555 11857 3607
rect 11913 3555 11965 3607
rect 12021 3555 12073 3607
rect 11805 3447 11857 3499
rect 11913 3447 11965 3499
rect 12021 3447 12073 3499
rect 11805 3339 11857 3391
rect 11913 3339 11965 3391
rect 12021 3339 12073 3391
rect 11805 3231 11857 3283
rect 11913 3231 11965 3283
rect 12021 3231 12073 3283
rect 11805 3123 11857 3175
rect 11913 3123 11965 3175
rect 12021 3123 12073 3175
rect 11805 3015 11857 3067
rect 11913 3015 11965 3067
rect 12021 3015 12073 3067
rect 11805 2907 11857 2959
rect 11913 2907 11965 2959
rect 12021 2907 12073 2959
rect 11805 2799 11857 2851
rect 11913 2799 11965 2851
rect 12021 2799 12073 2851
rect 11805 2691 11857 2743
rect 11913 2691 11965 2743
rect 12021 2691 12073 2743
rect 11805 2583 11857 2635
rect 11913 2583 11965 2635
rect 12021 2583 12073 2635
rect 11805 2475 11857 2527
rect 11913 2475 11965 2527
rect 12021 2475 12073 2527
rect 11805 2367 11857 2419
rect 11913 2367 11965 2419
rect 12021 2367 12073 2419
rect 11805 2259 11857 2311
rect 11913 2259 11965 2311
rect 12021 2259 12073 2311
rect 11805 2151 11857 2203
rect 11913 2151 11965 2203
rect 12021 2151 12073 2203
rect 11805 2043 11857 2095
rect 11913 2043 11965 2095
rect 12021 2043 12073 2095
rect 11805 1935 11857 1987
rect 11913 1935 11965 1987
rect 12021 1935 12073 1987
rect 11805 1827 11857 1879
rect 11913 1827 11965 1879
rect 12021 1827 12073 1879
rect 11805 1719 11857 1771
rect 11913 1719 11965 1771
rect 12021 1719 12073 1771
rect 11805 1611 11857 1663
rect 11913 1611 11965 1663
rect 12021 1611 12073 1663
rect 11805 1503 11857 1555
rect 11913 1503 11965 1555
rect 12021 1503 12073 1555
rect 11805 1395 11857 1447
rect 11913 1395 11965 1447
rect 12021 1395 12073 1447
rect 11805 1287 11857 1339
rect 11913 1287 11965 1339
rect 12021 1287 12073 1339
rect 11805 1179 11857 1231
rect 11913 1179 11965 1231
rect 12021 1179 12073 1231
rect 11805 1071 11857 1123
rect 11913 1071 11965 1123
rect 12021 1071 12073 1123
rect 11805 963 11857 1015
rect 11913 963 11965 1015
rect 12021 963 12073 1015
rect 11805 855 11857 907
rect 11913 855 11965 907
rect 12021 855 12073 907
rect 11805 747 11857 799
rect 11913 747 11965 799
rect 12021 747 12073 799
rect 11805 639 11857 691
rect 11913 639 11965 691
rect 12021 639 12073 691
rect 11805 531 11857 583
rect 11913 531 11965 583
rect 12021 531 12073 583
rect 189 423 241 475
rect 297 423 349 475
rect 405 423 457 475
rect 189 315 241 367
rect 297 315 349 367
rect 405 315 457 367
rect 189 207 241 259
rect 297 207 349 259
rect 405 207 457 259
rect 189 99 241 151
rect 297 99 349 151
rect 405 99 457 151
rect 1173 437 1225 489
rect 1297 437 1349 489
rect 1421 437 1473 489
rect 1545 437 1597 489
rect 3445 437 3497 489
rect 3569 437 3621 489
rect 3693 437 3745 489
rect 3817 437 3869 489
rect 5738 437 5790 489
rect 5862 437 5914 489
rect 5986 437 6038 489
rect 6224 437 6276 489
rect 6348 437 6400 489
rect 6472 437 6524 489
rect 8393 437 8445 489
rect 8517 437 8569 489
rect 8641 437 8693 489
rect 8765 437 8817 489
rect 10665 437 10717 489
rect 10789 437 10841 489
rect 10913 437 10965 489
rect 11037 437 11089 489
rect 1173 313 1225 365
rect 1297 313 1349 365
rect 1421 313 1473 365
rect 1545 313 1597 365
rect 3445 313 3497 365
rect 3569 313 3621 365
rect 3693 313 3745 365
rect 3817 313 3869 365
rect 5738 313 5790 365
rect 5862 313 5914 365
rect 5986 313 6038 365
rect 6224 313 6276 365
rect 6348 313 6400 365
rect 6472 313 6524 365
rect 8393 313 8445 365
rect 8517 313 8569 365
rect 8641 313 8693 365
rect 8765 313 8817 365
rect 10665 313 10717 365
rect 10789 313 10841 365
rect 10913 313 10965 365
rect 11037 313 11089 365
rect 1173 189 1225 241
rect 1297 189 1349 241
rect 1421 189 1473 241
rect 1545 189 1597 241
rect 3445 189 3497 241
rect 3569 189 3621 241
rect 3693 189 3745 241
rect 3817 189 3869 241
rect 5738 189 5790 241
rect 5862 189 5914 241
rect 5986 189 6038 241
rect 6224 189 6276 241
rect 6348 189 6400 241
rect 6472 189 6524 241
rect 8393 189 8445 241
rect 8517 189 8569 241
rect 8641 189 8693 241
rect 8765 189 8817 241
rect 10665 189 10717 241
rect 10789 189 10841 241
rect 10913 189 10965 241
rect 11037 189 11089 241
rect 1173 65 1225 117
rect 1297 65 1349 117
rect 1421 65 1473 117
rect 1545 65 1597 117
rect 3445 65 3497 117
rect 3569 65 3621 117
rect 3693 65 3745 117
rect 3817 65 3869 117
rect 5738 65 5790 117
rect 5862 65 5914 117
rect 5986 65 6038 117
rect 6224 65 6276 117
rect 6348 65 6400 117
rect 6472 65 6524 117
rect 8393 65 8445 117
rect 8517 65 8569 117
rect 8641 65 8693 117
rect 8765 65 8817 117
rect 10665 65 10717 117
rect 10789 65 10841 117
rect 10913 65 10965 117
rect 11037 65 11089 117
rect 11805 423 11857 475
rect 11913 423 11965 475
rect 12021 423 12073 475
rect 11805 315 11857 367
rect 11913 315 11965 367
rect 12021 315 12073 367
rect 11805 207 11857 259
rect 11913 207 11965 259
rect 12021 207 12073 259
rect 11805 99 11857 151
rect 11913 99 11965 151
rect 12021 99 12073 151
<< metal2 >>
rect -5 6955 503 14905
rect -5 6903 189 6955
rect 241 6903 297 6955
rect 349 6903 405 6955
rect 457 6903 503 6955
rect -5 6847 503 6903
rect -5 6795 189 6847
rect 241 6795 297 6847
rect 349 6795 405 6847
rect 457 6795 503 6847
rect -5 6739 503 6795
rect -5 6687 189 6739
rect 241 6687 297 6739
rect 349 6687 405 6739
rect 457 6687 503 6739
rect -5 6631 503 6687
rect -5 6579 189 6631
rect 241 6579 297 6631
rect 349 6579 405 6631
rect 457 6579 503 6631
rect -5 6523 503 6579
rect -5 6471 189 6523
rect 241 6471 297 6523
rect 349 6471 405 6523
rect 457 6471 503 6523
rect -5 6415 503 6471
rect -5 6363 189 6415
rect 241 6363 297 6415
rect 349 6363 405 6415
rect 457 6363 503 6415
rect -5 6307 503 6363
rect -5 6255 189 6307
rect 241 6255 297 6307
rect 349 6255 405 6307
rect 457 6255 503 6307
rect -5 6199 503 6255
rect -5 6147 189 6199
rect 241 6147 297 6199
rect 349 6147 405 6199
rect 457 6147 503 6199
rect -5 6091 503 6147
rect -5 6039 189 6091
rect 241 6039 297 6091
rect 349 6039 405 6091
rect 457 6039 503 6091
rect -5 5983 503 6039
rect -5 5931 189 5983
rect 241 5931 297 5983
rect 349 5931 405 5983
rect 457 5931 503 5983
rect -5 5875 503 5931
rect -5 5823 189 5875
rect 241 5823 297 5875
rect 349 5823 405 5875
rect 457 5823 503 5875
rect -5 5767 503 5823
rect -5 5715 189 5767
rect 241 5715 297 5767
rect 349 5715 405 5767
rect 457 5715 503 5767
rect -5 5659 503 5715
rect -5 5607 189 5659
rect 241 5607 297 5659
rect 349 5607 405 5659
rect 457 5607 503 5659
rect -5 5551 503 5607
rect -5 5499 189 5551
rect 241 5499 297 5551
rect 349 5499 405 5551
rect 457 5499 503 5551
rect -5 5443 503 5499
rect -5 5391 189 5443
rect 241 5391 297 5443
rect 349 5391 405 5443
rect 457 5391 503 5443
rect -5 5335 503 5391
rect -5 5283 189 5335
rect 241 5283 297 5335
rect 349 5283 405 5335
rect 457 5283 503 5335
rect -5 5227 503 5283
rect -5 5175 189 5227
rect 241 5175 297 5227
rect 349 5175 405 5227
rect 457 5175 503 5227
rect -5 5119 503 5175
rect -5 5067 189 5119
rect 241 5067 297 5119
rect 349 5067 405 5119
rect 457 5067 503 5119
rect -5 5011 503 5067
rect -5 4959 189 5011
rect 241 4959 297 5011
rect 349 4959 405 5011
rect 457 4959 503 5011
rect -5 4903 503 4959
rect -5 4851 189 4903
rect 241 4851 297 4903
rect 349 4851 405 4903
rect 457 4851 503 4903
rect -5 4795 503 4851
rect -5 4743 189 4795
rect 241 4743 297 4795
rect 349 4743 405 4795
rect 457 4743 503 4795
rect -5 4687 503 4743
rect -5 4635 189 4687
rect 241 4635 297 4687
rect 349 4635 405 4687
rect 457 4635 503 4687
rect -5 4579 503 4635
rect -5 4527 189 4579
rect 241 4527 297 4579
rect 349 4527 405 4579
rect 457 4527 503 4579
rect -5 4471 503 4527
rect -5 4419 189 4471
rect 241 4419 297 4471
rect 349 4419 405 4471
rect 457 4419 503 4471
rect -5 4363 503 4419
rect -5 4311 189 4363
rect 241 4311 297 4363
rect 349 4311 405 4363
rect 457 4311 503 4363
rect -5 4255 503 4311
rect -5 4203 189 4255
rect 241 4203 297 4255
rect 349 4203 405 4255
rect 457 4203 503 4255
rect -5 4147 503 4203
rect -5 4095 189 4147
rect 241 4095 297 4147
rect 349 4095 405 4147
rect 457 4095 503 4147
rect -5 4039 503 4095
rect -5 3987 189 4039
rect 241 3987 297 4039
rect 349 3987 405 4039
rect 457 3987 503 4039
rect -5 3931 503 3987
rect -5 3879 189 3931
rect 241 3879 297 3931
rect 349 3879 405 3931
rect 457 3879 503 3931
rect -5 3823 503 3879
rect -5 3771 189 3823
rect 241 3771 297 3823
rect 349 3771 405 3823
rect 457 3771 503 3823
rect -5 3715 503 3771
rect -5 3663 189 3715
rect 241 3663 297 3715
rect 349 3663 405 3715
rect 457 3663 503 3715
rect -5 3607 503 3663
rect -5 3555 189 3607
rect 241 3555 297 3607
rect 349 3555 405 3607
rect 457 3555 503 3607
rect -5 3499 503 3555
rect -5 3447 189 3499
rect 241 3447 297 3499
rect 349 3447 405 3499
rect 457 3447 503 3499
rect -5 3391 503 3447
rect -5 3339 189 3391
rect 241 3339 297 3391
rect 349 3339 405 3391
rect 457 3339 503 3391
rect -5 3283 503 3339
rect -5 3231 189 3283
rect 241 3231 297 3283
rect 349 3231 405 3283
rect 457 3231 503 3283
rect -5 3175 503 3231
rect -5 3123 189 3175
rect 241 3123 297 3175
rect 349 3123 405 3175
rect 457 3123 503 3175
rect -5 3067 503 3123
rect -5 3015 189 3067
rect 241 3015 297 3067
rect 349 3015 405 3067
rect 457 3015 503 3067
rect -5 2959 503 3015
rect -5 2907 189 2959
rect 241 2907 297 2959
rect 349 2907 405 2959
rect 457 2907 503 2959
rect -5 2851 503 2907
rect -5 2799 189 2851
rect 241 2799 297 2851
rect 349 2799 405 2851
rect 457 2799 503 2851
rect -5 2743 503 2799
rect -5 2691 189 2743
rect 241 2691 297 2743
rect 349 2691 405 2743
rect 457 2691 503 2743
rect -5 2635 503 2691
rect -5 2583 189 2635
rect 241 2583 297 2635
rect 349 2583 405 2635
rect 457 2583 503 2635
rect -5 2527 503 2583
rect -5 2475 189 2527
rect 241 2475 297 2527
rect 349 2475 405 2527
rect 457 2475 503 2527
rect -5 2419 503 2475
rect -5 2367 189 2419
rect 241 2367 297 2419
rect 349 2367 405 2419
rect 457 2367 503 2419
rect -5 2311 503 2367
rect -5 2259 189 2311
rect 241 2259 297 2311
rect 349 2259 405 2311
rect 457 2259 503 2311
rect -5 2203 503 2259
rect -5 2151 189 2203
rect 241 2151 297 2203
rect 349 2151 405 2203
rect 457 2151 503 2203
rect -5 2095 503 2151
rect -5 2043 189 2095
rect 241 2043 297 2095
rect 349 2043 405 2095
rect 457 2043 503 2095
rect -5 1987 503 2043
rect -5 1935 189 1987
rect 241 1935 297 1987
rect 349 1935 405 1987
rect 457 1935 503 1987
rect -5 1879 503 1935
rect -5 1827 189 1879
rect 241 1827 297 1879
rect 349 1827 405 1879
rect 457 1827 503 1879
rect -5 1771 503 1827
rect -5 1719 189 1771
rect 241 1719 297 1771
rect 349 1719 405 1771
rect 457 1719 503 1771
rect -5 1663 503 1719
rect -5 1611 189 1663
rect 241 1611 297 1663
rect 349 1611 405 1663
rect 457 1611 503 1663
rect -5 1555 503 1611
rect -5 1503 189 1555
rect 241 1503 297 1555
rect 349 1503 405 1555
rect 457 1503 503 1555
rect -5 1447 503 1503
rect -5 1395 189 1447
rect 241 1395 297 1447
rect 349 1395 405 1447
rect 457 1395 503 1447
rect -5 1339 503 1395
rect -5 1287 189 1339
rect 241 1287 297 1339
rect 349 1287 405 1339
rect 457 1287 503 1339
rect -5 1231 503 1287
rect -5 1179 189 1231
rect 241 1179 297 1231
rect 349 1179 405 1231
rect 457 1179 503 1231
rect -5 1123 503 1179
rect -5 1071 189 1123
rect 241 1071 297 1123
rect 349 1071 405 1123
rect 457 1071 503 1123
rect -5 1015 503 1071
rect -5 963 189 1015
rect 241 963 297 1015
rect 349 963 405 1015
rect 457 963 503 1015
rect -5 907 503 963
rect -5 855 189 907
rect 241 855 297 907
rect 349 855 405 907
rect 457 855 503 907
rect -5 799 503 855
rect -5 747 189 799
rect 241 747 297 799
rect 349 747 405 799
rect 457 747 503 799
rect -5 691 503 747
rect -5 639 189 691
rect 241 639 297 691
rect 349 639 405 691
rect 457 639 503 691
rect -5 583 503 639
rect -5 531 189 583
rect 241 531 297 583
rect 349 531 405 583
rect 457 531 503 583
rect -5 475 503 531
rect -5 423 189 475
rect 241 423 297 475
rect 349 423 405 475
rect 457 423 503 475
rect -5 367 503 423
rect -5 315 189 367
rect 241 315 297 367
rect 349 315 405 367
rect 457 315 503 367
rect -5 259 503 315
rect -5 207 189 259
rect 241 207 297 259
rect 349 207 405 259
rect 457 207 503 259
rect -5 151 503 207
rect -5 99 189 151
rect 241 99 297 151
rect 349 99 405 151
rect 457 99 503 151
rect -5 43 503 99
rect 563 14396 1071 14905
rect 563 14344 605 14396
rect 657 14344 729 14396
rect 781 14344 853 14396
rect 905 14344 977 14396
rect 1029 14344 1071 14396
rect 563 14272 1071 14344
rect 563 14220 605 14272
rect 657 14220 729 14272
rect 781 14220 853 14272
rect 905 14220 977 14272
rect 1029 14220 1071 14272
rect 563 14148 1071 14220
rect 563 14096 605 14148
rect 657 14096 729 14148
rect 781 14096 853 14148
rect 905 14096 977 14148
rect 1029 14096 1071 14148
rect 563 14024 1071 14096
rect 563 13972 605 14024
rect 657 13972 729 14024
rect 781 13972 853 14024
rect 905 13972 977 14024
rect 1029 13972 1071 14024
rect 563 7896 1071 13972
rect 563 7844 605 7896
rect 657 7844 729 7896
rect 781 7844 853 7896
rect 905 7844 977 7896
rect 1029 7844 1071 7896
rect 563 7772 1071 7844
rect 563 7720 605 7772
rect 657 7720 729 7772
rect 781 7720 853 7772
rect 905 7720 977 7772
rect 1029 7720 1071 7772
rect 563 7648 1071 7720
rect 563 7596 605 7648
rect 657 7596 729 7648
rect 781 7596 853 7648
rect 905 7596 977 7648
rect 1029 7596 1071 7648
rect 563 7524 1071 7596
rect 563 7472 605 7524
rect 657 7472 729 7524
rect 781 7472 853 7524
rect 905 7472 977 7524
rect 1029 7472 1071 7524
rect 563 6307 1071 7472
rect 563 6255 737 6307
rect 789 6255 845 6307
rect 897 6255 1071 6307
rect 563 6199 1071 6255
rect 563 6147 737 6199
rect 789 6147 845 6199
rect 897 6147 1071 6199
rect 563 6091 1071 6147
rect 563 6039 737 6091
rect 789 6039 845 6091
rect 897 6039 1071 6091
rect 563 5983 1071 6039
rect 563 5931 737 5983
rect 789 5931 845 5983
rect 897 5931 1071 5983
rect 563 5875 1071 5931
rect 563 5823 737 5875
rect 789 5823 845 5875
rect 897 5823 1071 5875
rect 563 5767 1071 5823
rect 563 5715 737 5767
rect 789 5715 845 5767
rect 897 5715 1071 5767
rect 563 5659 1071 5715
rect 563 5607 737 5659
rect 789 5607 845 5659
rect 897 5607 1071 5659
rect 563 5551 1071 5607
rect 563 5499 737 5551
rect 789 5499 845 5551
rect 897 5499 1071 5551
rect 563 5443 1071 5499
rect 563 5391 737 5443
rect 789 5391 845 5443
rect 897 5391 1071 5443
rect 563 5335 1071 5391
rect 563 5283 737 5335
rect 789 5283 845 5335
rect 897 5283 1071 5335
rect 563 5227 1071 5283
rect 563 5175 737 5227
rect 789 5175 845 5227
rect 897 5175 1071 5227
rect 563 5119 1071 5175
rect 563 5067 737 5119
rect 789 5067 845 5119
rect 897 5067 1071 5119
rect 563 5011 1071 5067
rect 563 4959 737 5011
rect 789 4959 845 5011
rect 897 4959 1071 5011
rect 563 4903 1071 4959
rect 563 4851 737 4903
rect 789 4851 845 4903
rect 897 4851 1071 4903
rect 563 4795 1071 4851
rect 563 4743 737 4795
rect 789 4743 845 4795
rect 897 4743 1071 4795
rect 563 4687 1071 4743
rect 563 4635 737 4687
rect 789 4635 845 4687
rect 897 4635 1071 4687
rect 563 4579 1071 4635
rect 563 4527 737 4579
rect 789 4527 845 4579
rect 897 4527 1071 4579
rect 563 4471 1071 4527
rect 563 4419 737 4471
rect 789 4419 845 4471
rect 897 4419 1071 4471
rect 563 4363 1071 4419
rect 563 4311 737 4363
rect 789 4311 845 4363
rect 897 4311 1071 4363
rect 563 4255 1071 4311
rect 563 4203 737 4255
rect 789 4203 845 4255
rect 897 4203 1071 4255
rect 563 4147 1071 4203
rect 563 4095 737 4147
rect 789 4095 845 4147
rect 897 4095 1071 4147
rect 563 4039 1071 4095
rect 563 3987 737 4039
rect 789 3987 845 4039
rect 897 3987 1071 4039
rect 563 3931 1071 3987
rect 563 3879 737 3931
rect 789 3879 845 3931
rect 897 3879 1071 3931
rect 563 3823 1071 3879
rect 563 3771 737 3823
rect 789 3771 845 3823
rect 897 3771 1071 3823
rect 563 3715 1071 3771
rect 563 3663 737 3715
rect 789 3663 845 3715
rect 897 3663 1071 3715
rect 563 3607 1071 3663
rect 563 3555 737 3607
rect 789 3555 845 3607
rect 897 3555 1071 3607
rect 563 3499 1071 3555
rect 563 3447 737 3499
rect 789 3447 845 3499
rect 897 3447 1071 3499
rect 563 3391 1071 3447
rect 563 3339 737 3391
rect 789 3339 845 3391
rect 897 3339 1071 3391
rect 563 3283 1071 3339
rect 563 3231 737 3283
rect 789 3231 845 3283
rect 897 3231 1071 3283
rect 563 3175 1071 3231
rect 563 3123 737 3175
rect 789 3123 845 3175
rect 897 3123 1071 3175
rect 563 3067 1071 3123
rect 563 3015 737 3067
rect 789 3015 845 3067
rect 897 3015 1071 3067
rect 563 2959 1071 3015
rect 563 2907 737 2959
rect 789 2907 845 2959
rect 897 2907 1071 2959
rect 563 2851 1071 2907
rect 563 2799 737 2851
rect 789 2799 845 2851
rect 897 2799 1071 2851
rect 563 2743 1071 2799
rect 563 2691 737 2743
rect 789 2691 845 2743
rect 897 2691 1071 2743
rect 563 2635 1071 2691
rect 563 2583 737 2635
rect 789 2583 845 2635
rect 897 2583 1071 2635
rect 563 2527 1071 2583
rect 563 2475 737 2527
rect 789 2475 845 2527
rect 897 2475 1071 2527
rect 563 2419 1071 2475
rect 563 2367 737 2419
rect 789 2367 845 2419
rect 897 2367 1071 2419
rect 563 2311 1071 2367
rect 563 2259 737 2311
rect 789 2259 845 2311
rect 897 2259 1071 2311
rect 563 2203 1071 2259
rect 563 2151 737 2203
rect 789 2151 845 2203
rect 897 2151 1071 2203
rect 563 2095 1071 2151
rect 563 2043 737 2095
rect 789 2043 845 2095
rect 897 2043 1071 2095
rect 563 1987 1071 2043
rect 563 1935 737 1987
rect 789 1935 845 1987
rect 897 1935 1071 1987
rect 563 1879 1071 1935
rect 563 1827 737 1879
rect 789 1827 845 1879
rect 897 1827 1071 1879
rect 563 1771 1071 1827
rect 563 1719 737 1771
rect 789 1719 845 1771
rect 897 1719 1071 1771
rect 563 1663 1071 1719
rect 563 1611 737 1663
rect 789 1611 845 1663
rect 897 1611 1071 1663
rect 563 1555 1071 1611
rect 563 1503 737 1555
rect 789 1503 845 1555
rect 897 1503 1071 1555
rect 563 1447 1071 1503
rect 563 1395 737 1447
rect 789 1395 845 1447
rect 897 1395 1071 1447
rect 563 1339 1071 1395
rect 563 1287 737 1339
rect 789 1287 845 1339
rect 897 1287 1071 1339
rect 563 1231 1071 1287
rect 563 1179 737 1231
rect 789 1179 845 1231
rect 897 1179 1071 1231
rect 563 1123 1071 1179
rect 563 1071 737 1123
rect 789 1071 845 1123
rect 897 1071 1071 1123
rect 563 1015 1071 1071
rect 563 963 737 1015
rect 789 963 845 1015
rect 897 963 1071 1015
rect 563 907 1071 963
rect 563 855 737 907
rect 789 855 845 907
rect 897 855 1071 907
rect 563 799 1071 855
rect 563 747 737 799
rect 789 747 845 799
rect 897 747 1071 799
rect 563 43 1071 747
rect 1131 13745 1639 14905
rect 1131 13693 1143 13745
rect 1195 13693 1251 13745
rect 1303 13693 1359 13745
rect 1411 13693 1467 13745
rect 1519 13693 1575 13745
rect 1627 13693 1639 13745
rect 1131 13637 1639 13693
rect 1131 13585 1143 13637
rect 1195 13585 1251 13637
rect 1303 13585 1359 13637
rect 1411 13585 1467 13637
rect 1519 13585 1575 13637
rect 1627 13585 1639 13637
rect 1131 12472 1639 13585
rect 1131 12420 1143 12472
rect 1195 12420 1251 12472
rect 1303 12420 1359 12472
rect 1411 12420 1467 12472
rect 1519 12420 1575 12472
rect 1627 12420 1639 12472
rect 1131 12364 1639 12420
rect 1131 12312 1143 12364
rect 1195 12312 1251 12364
rect 1303 12312 1359 12364
rect 1411 12312 1467 12364
rect 1519 12312 1575 12364
rect 1627 12312 1639 12364
rect 1131 12256 1639 12312
rect 1131 12204 1143 12256
rect 1195 12204 1251 12256
rect 1303 12204 1359 12256
rect 1411 12204 1467 12256
rect 1519 12204 1575 12256
rect 1627 12204 1639 12256
rect 1131 11068 1639 12204
rect 1131 11016 1143 11068
rect 1195 11016 1251 11068
rect 1303 11016 1359 11068
rect 1411 11016 1467 11068
rect 1519 11016 1575 11068
rect 1627 11016 1639 11068
rect 1131 10960 1639 11016
rect 1131 10908 1143 10960
rect 1195 10908 1251 10960
rect 1303 10908 1359 10960
rect 1411 10908 1467 10960
rect 1519 10908 1575 10960
rect 1627 10908 1639 10960
rect 1131 10852 1639 10908
rect 1131 10800 1143 10852
rect 1195 10800 1251 10852
rect 1303 10800 1359 10852
rect 1411 10800 1467 10852
rect 1519 10800 1575 10852
rect 1627 10800 1639 10852
rect 1131 9664 1639 10800
rect 1131 9612 1143 9664
rect 1195 9612 1251 9664
rect 1303 9612 1359 9664
rect 1411 9612 1467 9664
rect 1519 9612 1575 9664
rect 1627 9612 1639 9664
rect 1131 9556 1639 9612
rect 1131 9504 1143 9556
rect 1195 9504 1251 9556
rect 1303 9504 1359 9556
rect 1411 9504 1467 9556
rect 1519 9504 1575 9556
rect 1627 9504 1639 9556
rect 1131 9448 1639 9504
rect 1131 9396 1143 9448
rect 1195 9396 1251 9448
rect 1303 9396 1359 9448
rect 1411 9396 1467 9448
rect 1519 9396 1575 9448
rect 1627 9396 1639 9448
rect 1131 8283 1639 9396
rect 1131 8231 1143 8283
rect 1195 8231 1251 8283
rect 1303 8231 1359 8283
rect 1411 8231 1467 8283
rect 1519 8231 1575 8283
rect 1627 8231 1639 8283
rect 1131 8175 1639 8231
rect 1131 8123 1143 8175
rect 1195 8123 1251 8175
rect 1303 8123 1359 8175
rect 1411 8123 1467 8175
rect 1519 8123 1575 8175
rect 1627 8123 1639 8175
rect 1131 6989 1639 8123
rect 1131 6937 1173 6989
rect 1225 6937 1297 6989
rect 1349 6937 1421 6989
rect 1473 6937 1545 6989
rect 1597 6937 1639 6989
rect 1131 6865 1639 6937
rect 1131 6813 1173 6865
rect 1225 6813 1297 6865
rect 1349 6813 1421 6865
rect 1473 6813 1545 6865
rect 1597 6813 1639 6865
rect 1131 6741 1639 6813
rect 1131 6689 1173 6741
rect 1225 6689 1297 6741
rect 1349 6689 1421 6741
rect 1473 6689 1545 6741
rect 1597 6689 1639 6741
rect 1131 6617 1639 6689
rect 1131 6565 1173 6617
rect 1225 6565 1297 6617
rect 1349 6565 1421 6617
rect 1473 6565 1545 6617
rect 1597 6565 1639 6617
rect 1131 489 1639 6565
rect 1131 437 1173 489
rect 1225 437 1297 489
rect 1349 437 1421 489
rect 1473 437 1545 489
rect 1597 437 1639 489
rect 1131 365 1639 437
rect 1131 313 1173 365
rect 1225 313 1297 365
rect 1349 313 1421 365
rect 1473 313 1545 365
rect 1597 313 1639 365
rect 1131 241 1639 313
rect 1131 189 1173 241
rect 1225 189 1297 241
rect 1349 189 1421 241
rect 1473 189 1545 241
rect 1597 189 1639 241
rect 1131 117 1639 189
rect 1131 65 1173 117
rect 1225 65 1297 117
rect 1349 65 1421 117
rect 1473 65 1545 117
rect 1597 65 1639 117
rect 1131 43 1639 65
rect 1699 13314 2207 56440
rect 1699 13262 1741 13314
rect 1793 13262 1865 13314
rect 1917 13262 1989 13314
rect 2041 13262 2113 13314
rect 2165 13262 2207 13314
rect 1699 13190 2207 13262
rect 1699 13138 1741 13190
rect 1793 13138 1865 13190
rect 1917 13138 1989 13190
rect 2041 13138 2113 13190
rect 2165 13138 2207 13190
rect 1699 13066 2207 13138
rect 1699 13014 1741 13066
rect 1793 13014 1865 13066
rect 1917 13014 1989 13066
rect 2041 13014 2113 13066
rect 2165 13014 2207 13066
rect 1699 12942 2207 13014
rect 1699 12890 1741 12942
rect 1793 12890 1865 12942
rect 1917 12890 1989 12942
rect 2041 12890 2113 12942
rect 2165 12890 2207 12942
rect 1699 12818 2207 12890
rect 1699 12766 1741 12818
rect 1793 12766 1865 12818
rect 1917 12766 1989 12818
rect 2041 12766 2113 12818
rect 2165 12766 2207 12818
rect 1699 11910 2207 12766
rect 1699 11858 1741 11910
rect 1793 11858 1865 11910
rect 1917 11858 1989 11910
rect 2041 11858 2113 11910
rect 2165 11858 2207 11910
rect 1699 11786 2207 11858
rect 1699 11734 1741 11786
rect 1793 11734 1865 11786
rect 1917 11734 1989 11786
rect 2041 11734 2113 11786
rect 2165 11734 2207 11786
rect 1699 11662 2207 11734
rect 1699 11610 1741 11662
rect 1793 11610 1865 11662
rect 1917 11610 1989 11662
rect 2041 11610 2113 11662
rect 2165 11610 2207 11662
rect 1699 11538 2207 11610
rect 1699 11486 1741 11538
rect 1793 11486 1865 11538
rect 1917 11486 1989 11538
rect 2041 11486 2113 11538
rect 2165 11486 2207 11538
rect 1699 11414 2207 11486
rect 1699 11362 1741 11414
rect 1793 11362 1865 11414
rect 1917 11362 1989 11414
rect 2041 11362 2113 11414
rect 2165 11362 2207 11414
rect 1699 10506 2207 11362
rect 1699 10454 1741 10506
rect 1793 10454 1865 10506
rect 1917 10454 1989 10506
rect 2041 10454 2113 10506
rect 2165 10454 2207 10506
rect 1699 10382 2207 10454
rect 1699 10330 1741 10382
rect 1793 10330 1865 10382
rect 1917 10330 1989 10382
rect 2041 10330 2113 10382
rect 2165 10330 2207 10382
rect 1699 10258 2207 10330
rect 1699 10206 1741 10258
rect 1793 10206 1865 10258
rect 1917 10206 1989 10258
rect 2041 10206 2113 10258
rect 2165 10206 2207 10258
rect 1699 10134 2207 10206
rect 1699 10082 1741 10134
rect 1793 10082 1865 10134
rect 1917 10082 1989 10134
rect 2041 10082 2113 10134
rect 2165 10082 2207 10134
rect 1699 10010 2207 10082
rect 1699 9958 1741 10010
rect 1793 9958 1865 10010
rect 1917 9958 1989 10010
rect 2041 9958 2113 10010
rect 2165 9958 2207 10010
rect 1699 9102 2207 9958
rect 1699 9050 1741 9102
rect 1793 9050 1865 9102
rect 1917 9050 1989 9102
rect 2041 9050 2113 9102
rect 2165 9050 2207 9102
rect 1699 8978 2207 9050
rect 1699 8926 1741 8978
rect 1793 8926 1865 8978
rect 1917 8926 1989 8978
rect 2041 8926 2113 8978
rect 2165 8926 2207 8978
rect 1699 8854 2207 8926
rect 1699 8802 1741 8854
rect 1793 8802 1865 8854
rect 1917 8802 1989 8854
rect 2041 8802 2113 8854
rect 2165 8802 2207 8854
rect 1699 8730 2207 8802
rect 1699 8678 1741 8730
rect 1793 8678 1865 8730
rect 1917 8678 1989 8730
rect 2041 8678 2113 8730
rect 2165 8678 2207 8730
rect 1699 8606 2207 8678
rect 1699 8554 1741 8606
rect 1793 8554 1865 8606
rect 1917 8554 1989 8606
rect 2041 8554 2113 8606
rect 2165 8554 2207 8606
rect 1699 5907 2207 8554
rect 1699 5855 1741 5907
rect 1793 5855 1865 5907
rect 1917 5855 1989 5907
rect 2041 5855 2113 5907
rect 2165 5855 2207 5907
rect 1699 5783 2207 5855
rect 1699 5731 1741 5783
rect 1793 5731 1865 5783
rect 1917 5731 1989 5783
rect 2041 5731 2113 5783
rect 2165 5731 2207 5783
rect 1699 5659 2207 5731
rect 1699 5607 1741 5659
rect 1793 5607 1865 5659
rect 1917 5607 1989 5659
rect 2041 5607 2113 5659
rect 2165 5607 2207 5659
rect 1699 5535 2207 5607
rect 1699 5483 1741 5535
rect 1793 5483 1865 5535
rect 1917 5483 1989 5535
rect 2041 5483 2113 5535
rect 2165 5483 2207 5535
rect 1699 5411 2207 5483
rect 1699 5359 1741 5411
rect 1793 5359 1865 5411
rect 1917 5359 1989 5411
rect 2041 5359 2113 5411
rect 2165 5359 2207 5411
rect 1699 4503 2207 5359
rect 1699 4451 1741 4503
rect 1793 4451 1865 4503
rect 1917 4451 1989 4503
rect 2041 4451 2113 4503
rect 2165 4451 2207 4503
rect 1699 4379 2207 4451
rect 1699 4327 1741 4379
rect 1793 4327 1865 4379
rect 1917 4327 1989 4379
rect 2041 4327 2113 4379
rect 2165 4327 2207 4379
rect 1699 4255 2207 4327
rect 1699 4203 1741 4255
rect 1793 4203 1865 4255
rect 1917 4203 1989 4255
rect 2041 4203 2113 4255
rect 2165 4203 2207 4255
rect 1699 4131 2207 4203
rect 1699 4079 1741 4131
rect 1793 4079 1865 4131
rect 1917 4079 1989 4131
rect 2041 4079 2113 4131
rect 2165 4079 2207 4131
rect 1699 4007 2207 4079
rect 1699 3955 1741 4007
rect 1793 3955 1865 4007
rect 1917 3955 1989 4007
rect 2041 3955 2113 4007
rect 2165 3955 2207 4007
rect 1699 3099 2207 3955
rect 1699 3047 1741 3099
rect 1793 3047 1865 3099
rect 1917 3047 1989 3099
rect 2041 3047 2113 3099
rect 2165 3047 2207 3099
rect 1699 2975 2207 3047
rect 1699 2923 1741 2975
rect 1793 2923 1865 2975
rect 1917 2923 1989 2975
rect 2041 2923 2113 2975
rect 2165 2923 2207 2975
rect 1699 2851 2207 2923
rect 1699 2799 1741 2851
rect 1793 2799 1865 2851
rect 1917 2799 1989 2851
rect 2041 2799 2113 2851
rect 2165 2799 2207 2851
rect 1699 2727 2207 2799
rect 1699 2675 1741 2727
rect 1793 2675 1865 2727
rect 1917 2675 1989 2727
rect 2041 2675 2113 2727
rect 2165 2675 2207 2727
rect 1699 2603 2207 2675
rect 1699 2551 1741 2603
rect 1793 2551 1865 2603
rect 1917 2551 1989 2603
rect 2041 2551 2113 2603
rect 2165 2551 2207 2603
rect 1699 1695 2207 2551
rect 1699 1643 1741 1695
rect 1793 1643 1865 1695
rect 1917 1643 1989 1695
rect 2041 1643 2113 1695
rect 2165 1643 2207 1695
rect 1699 1571 2207 1643
rect 1699 1519 1741 1571
rect 1793 1519 1865 1571
rect 1917 1519 1989 1571
rect 2041 1519 2113 1571
rect 2165 1519 2207 1571
rect 1699 1447 2207 1519
rect 1699 1395 1741 1447
rect 1793 1395 1865 1447
rect 1917 1395 1989 1447
rect 2041 1395 2113 1447
rect 2165 1395 2207 1447
rect 1699 1323 2207 1395
rect 1699 1271 1741 1323
rect 1793 1271 1865 1323
rect 1917 1271 1989 1323
rect 2041 1271 2113 1323
rect 2165 1271 2207 1323
rect 1699 1199 2207 1271
rect 1699 1147 1741 1199
rect 1793 1147 1865 1199
rect 1917 1147 1989 1199
rect 2041 1147 2113 1199
rect 2165 1147 2207 1199
rect 1699 -857 2207 1147
rect 2267 14396 2775 14905
rect 2267 14344 2309 14396
rect 2361 14344 2433 14396
rect 2485 14344 2557 14396
rect 2609 14344 2681 14396
rect 2733 14344 2775 14396
rect 2267 14272 2775 14344
rect 2267 14220 2309 14272
rect 2361 14220 2433 14272
rect 2485 14220 2557 14272
rect 2609 14220 2681 14272
rect 2733 14220 2775 14272
rect 2267 14148 2775 14220
rect 2267 14096 2309 14148
rect 2361 14096 2433 14148
rect 2485 14096 2557 14148
rect 2609 14096 2681 14148
rect 2733 14096 2775 14148
rect 2267 14024 2775 14096
rect 2267 13972 2309 14024
rect 2361 13972 2433 14024
rect 2485 13972 2557 14024
rect 2609 13972 2681 14024
rect 2733 13972 2775 14024
rect 2267 7896 2775 13972
rect 2267 7844 2309 7896
rect 2361 7844 2433 7896
rect 2485 7844 2557 7896
rect 2609 7844 2681 7896
rect 2733 7844 2775 7896
rect 2267 7772 2775 7844
rect 2267 7720 2309 7772
rect 2361 7720 2433 7772
rect 2485 7720 2557 7772
rect 2609 7720 2681 7772
rect 2733 7720 2775 7772
rect 2267 7648 2775 7720
rect 2267 7596 2309 7648
rect 2361 7596 2433 7648
rect 2485 7596 2557 7648
rect 2609 7596 2681 7648
rect 2733 7596 2775 7648
rect 2267 7524 2775 7596
rect 2267 7472 2309 7524
rect 2361 7472 2433 7524
rect 2485 7472 2557 7524
rect 2609 7472 2681 7524
rect 2733 7472 2775 7524
rect 2267 6338 2775 7472
rect 2267 6286 2279 6338
rect 2331 6286 2387 6338
rect 2439 6286 2495 6338
rect 2547 6286 2603 6338
rect 2655 6286 2711 6338
rect 2763 6286 2775 6338
rect 2267 6230 2775 6286
rect 2267 6178 2279 6230
rect 2331 6178 2387 6230
rect 2439 6178 2495 6230
rect 2547 6178 2603 6230
rect 2655 6178 2711 6230
rect 2763 6178 2775 6230
rect 2267 5065 2775 6178
rect 2267 5013 2279 5065
rect 2331 5013 2387 5065
rect 2439 5013 2495 5065
rect 2547 5013 2603 5065
rect 2655 5013 2711 5065
rect 2763 5013 2775 5065
rect 2267 4957 2775 5013
rect 2267 4905 2279 4957
rect 2331 4905 2387 4957
rect 2439 4905 2495 4957
rect 2547 4905 2603 4957
rect 2655 4905 2711 4957
rect 2763 4905 2775 4957
rect 2267 4849 2775 4905
rect 2267 4797 2279 4849
rect 2331 4797 2387 4849
rect 2439 4797 2495 4849
rect 2547 4797 2603 4849
rect 2655 4797 2711 4849
rect 2763 4797 2775 4849
rect 2267 3661 2775 4797
rect 2267 3609 2279 3661
rect 2331 3609 2387 3661
rect 2439 3609 2495 3661
rect 2547 3609 2603 3661
rect 2655 3609 2711 3661
rect 2763 3609 2775 3661
rect 2267 3553 2775 3609
rect 2267 3501 2279 3553
rect 2331 3501 2387 3553
rect 2439 3501 2495 3553
rect 2547 3501 2603 3553
rect 2655 3501 2711 3553
rect 2763 3501 2775 3553
rect 2267 3445 2775 3501
rect 2267 3393 2279 3445
rect 2331 3393 2387 3445
rect 2439 3393 2495 3445
rect 2547 3393 2603 3445
rect 2655 3393 2711 3445
rect 2763 3393 2775 3445
rect 2267 2257 2775 3393
rect 2267 2205 2279 2257
rect 2331 2205 2387 2257
rect 2439 2205 2495 2257
rect 2547 2205 2603 2257
rect 2655 2205 2711 2257
rect 2763 2205 2775 2257
rect 2267 2149 2775 2205
rect 2267 2097 2279 2149
rect 2331 2097 2387 2149
rect 2439 2097 2495 2149
rect 2547 2097 2603 2149
rect 2655 2097 2711 2149
rect 2763 2097 2775 2149
rect 2267 2041 2775 2097
rect 2267 1989 2279 2041
rect 2331 1989 2387 2041
rect 2439 1989 2495 2041
rect 2547 1989 2603 2041
rect 2655 1989 2711 2041
rect 2763 1989 2775 2041
rect 2267 876 2775 1989
rect 2267 824 2279 876
rect 2331 824 2387 876
rect 2439 824 2495 876
rect 2547 824 2603 876
rect 2655 824 2711 876
rect 2763 824 2775 876
rect 2267 768 2775 824
rect 2267 716 2279 768
rect 2331 716 2387 768
rect 2439 716 2495 768
rect 2547 716 2603 768
rect 2655 716 2711 768
rect 2763 716 2775 768
rect 2267 43 2775 716
rect 2835 13314 3343 56440
rect 2835 13262 2877 13314
rect 2929 13262 3001 13314
rect 3053 13262 3125 13314
rect 3177 13262 3249 13314
rect 3301 13262 3343 13314
rect 2835 13190 3343 13262
rect 2835 13138 2877 13190
rect 2929 13138 3001 13190
rect 3053 13138 3125 13190
rect 3177 13138 3249 13190
rect 3301 13138 3343 13190
rect 2835 13066 3343 13138
rect 2835 13014 2877 13066
rect 2929 13014 3001 13066
rect 3053 13014 3125 13066
rect 3177 13014 3249 13066
rect 3301 13014 3343 13066
rect 2835 12942 3343 13014
rect 2835 12890 2877 12942
rect 2929 12890 3001 12942
rect 3053 12890 3125 12942
rect 3177 12890 3249 12942
rect 3301 12890 3343 12942
rect 2835 12818 3343 12890
rect 2835 12766 2877 12818
rect 2929 12766 3001 12818
rect 3053 12766 3125 12818
rect 3177 12766 3249 12818
rect 3301 12766 3343 12818
rect 2835 11910 3343 12766
rect 2835 11858 2877 11910
rect 2929 11858 3001 11910
rect 3053 11858 3125 11910
rect 3177 11858 3249 11910
rect 3301 11858 3343 11910
rect 2835 11786 3343 11858
rect 2835 11734 2877 11786
rect 2929 11734 3001 11786
rect 3053 11734 3125 11786
rect 3177 11734 3249 11786
rect 3301 11734 3343 11786
rect 2835 11662 3343 11734
rect 2835 11610 2877 11662
rect 2929 11610 3001 11662
rect 3053 11610 3125 11662
rect 3177 11610 3249 11662
rect 3301 11610 3343 11662
rect 2835 11538 3343 11610
rect 2835 11486 2877 11538
rect 2929 11486 3001 11538
rect 3053 11486 3125 11538
rect 3177 11486 3249 11538
rect 3301 11486 3343 11538
rect 2835 11414 3343 11486
rect 2835 11362 2877 11414
rect 2929 11362 3001 11414
rect 3053 11362 3125 11414
rect 3177 11362 3249 11414
rect 3301 11362 3343 11414
rect 2835 10506 3343 11362
rect 2835 10454 2877 10506
rect 2929 10454 3001 10506
rect 3053 10454 3125 10506
rect 3177 10454 3249 10506
rect 3301 10454 3343 10506
rect 2835 10382 3343 10454
rect 2835 10330 2877 10382
rect 2929 10330 3001 10382
rect 3053 10330 3125 10382
rect 3177 10330 3249 10382
rect 3301 10330 3343 10382
rect 2835 10258 3343 10330
rect 2835 10206 2877 10258
rect 2929 10206 3001 10258
rect 3053 10206 3125 10258
rect 3177 10206 3249 10258
rect 3301 10206 3343 10258
rect 2835 10134 3343 10206
rect 2835 10082 2877 10134
rect 2929 10082 3001 10134
rect 3053 10082 3125 10134
rect 3177 10082 3249 10134
rect 3301 10082 3343 10134
rect 2835 10010 3343 10082
rect 2835 9958 2877 10010
rect 2929 9958 3001 10010
rect 3053 9958 3125 10010
rect 3177 9958 3249 10010
rect 3301 9958 3343 10010
rect 2835 9102 3343 9958
rect 2835 9050 2877 9102
rect 2929 9050 3001 9102
rect 3053 9050 3125 9102
rect 3177 9050 3249 9102
rect 3301 9050 3343 9102
rect 2835 8978 3343 9050
rect 2835 8926 2877 8978
rect 2929 8926 3001 8978
rect 3053 8926 3125 8978
rect 3177 8926 3249 8978
rect 3301 8926 3343 8978
rect 2835 8854 3343 8926
rect 2835 8802 2877 8854
rect 2929 8802 3001 8854
rect 3053 8802 3125 8854
rect 3177 8802 3249 8854
rect 3301 8802 3343 8854
rect 2835 8730 3343 8802
rect 2835 8678 2877 8730
rect 2929 8678 3001 8730
rect 3053 8678 3125 8730
rect 3177 8678 3249 8730
rect 3301 8678 3343 8730
rect 2835 8606 3343 8678
rect 2835 8554 2877 8606
rect 2929 8554 3001 8606
rect 3053 8554 3125 8606
rect 3177 8554 3249 8606
rect 3301 8554 3343 8606
rect 2835 5907 3343 8554
rect 2835 5855 2877 5907
rect 2929 5855 3001 5907
rect 3053 5855 3125 5907
rect 3177 5855 3249 5907
rect 3301 5855 3343 5907
rect 2835 5783 3343 5855
rect 2835 5731 2877 5783
rect 2929 5731 3001 5783
rect 3053 5731 3125 5783
rect 3177 5731 3249 5783
rect 3301 5731 3343 5783
rect 2835 5659 3343 5731
rect 2835 5607 2877 5659
rect 2929 5607 3001 5659
rect 3053 5607 3125 5659
rect 3177 5607 3249 5659
rect 3301 5607 3343 5659
rect 2835 5535 3343 5607
rect 2835 5483 2877 5535
rect 2929 5483 3001 5535
rect 3053 5483 3125 5535
rect 3177 5483 3249 5535
rect 3301 5483 3343 5535
rect 2835 5411 3343 5483
rect 2835 5359 2877 5411
rect 2929 5359 3001 5411
rect 3053 5359 3125 5411
rect 3177 5359 3249 5411
rect 3301 5359 3343 5411
rect 2835 4503 3343 5359
rect 2835 4451 2877 4503
rect 2929 4451 3001 4503
rect 3053 4451 3125 4503
rect 3177 4451 3249 4503
rect 3301 4451 3343 4503
rect 2835 4379 3343 4451
rect 2835 4327 2877 4379
rect 2929 4327 3001 4379
rect 3053 4327 3125 4379
rect 3177 4327 3249 4379
rect 3301 4327 3343 4379
rect 2835 4255 3343 4327
rect 2835 4203 2877 4255
rect 2929 4203 3001 4255
rect 3053 4203 3125 4255
rect 3177 4203 3249 4255
rect 3301 4203 3343 4255
rect 2835 4131 3343 4203
rect 2835 4079 2877 4131
rect 2929 4079 3001 4131
rect 3053 4079 3125 4131
rect 3177 4079 3249 4131
rect 3301 4079 3343 4131
rect 2835 4007 3343 4079
rect 2835 3955 2877 4007
rect 2929 3955 3001 4007
rect 3053 3955 3125 4007
rect 3177 3955 3249 4007
rect 3301 3955 3343 4007
rect 2835 3099 3343 3955
rect 2835 3047 2877 3099
rect 2929 3047 3001 3099
rect 3053 3047 3125 3099
rect 3177 3047 3249 3099
rect 3301 3047 3343 3099
rect 2835 2975 3343 3047
rect 2835 2923 2877 2975
rect 2929 2923 3001 2975
rect 3053 2923 3125 2975
rect 3177 2923 3249 2975
rect 3301 2923 3343 2975
rect 2835 2851 3343 2923
rect 2835 2799 2877 2851
rect 2929 2799 3001 2851
rect 3053 2799 3125 2851
rect 3177 2799 3249 2851
rect 3301 2799 3343 2851
rect 2835 2727 3343 2799
rect 2835 2675 2877 2727
rect 2929 2675 3001 2727
rect 3053 2675 3125 2727
rect 3177 2675 3249 2727
rect 3301 2675 3343 2727
rect 2835 2603 3343 2675
rect 2835 2551 2877 2603
rect 2929 2551 3001 2603
rect 3053 2551 3125 2603
rect 3177 2551 3249 2603
rect 3301 2551 3343 2603
rect 2835 1695 3343 2551
rect 2835 1643 2877 1695
rect 2929 1643 3001 1695
rect 3053 1643 3125 1695
rect 3177 1643 3249 1695
rect 3301 1643 3343 1695
rect 2835 1571 3343 1643
rect 2835 1519 2877 1571
rect 2929 1519 3001 1571
rect 3053 1519 3125 1571
rect 3177 1519 3249 1571
rect 3301 1519 3343 1571
rect 2835 1447 3343 1519
rect 2835 1395 2877 1447
rect 2929 1395 3001 1447
rect 3053 1395 3125 1447
rect 3177 1395 3249 1447
rect 3301 1395 3343 1447
rect 2835 1323 3343 1395
rect 2835 1271 2877 1323
rect 2929 1271 3001 1323
rect 3053 1271 3125 1323
rect 3177 1271 3249 1323
rect 3301 1271 3343 1323
rect 2835 1199 3343 1271
rect 2835 1147 2877 1199
rect 2929 1147 3001 1199
rect 3053 1147 3125 1199
rect 3177 1147 3249 1199
rect 3301 1147 3343 1199
rect 2835 -857 3343 1147
rect 3403 13745 3911 14905
rect 3403 13693 3415 13745
rect 3467 13693 3523 13745
rect 3575 13693 3631 13745
rect 3683 13693 3739 13745
rect 3791 13693 3847 13745
rect 3899 13693 3911 13745
rect 3403 13637 3911 13693
rect 3403 13585 3415 13637
rect 3467 13585 3523 13637
rect 3575 13585 3631 13637
rect 3683 13585 3739 13637
rect 3791 13585 3847 13637
rect 3899 13585 3911 13637
rect 3403 12472 3911 13585
rect 3403 12420 3415 12472
rect 3467 12420 3523 12472
rect 3575 12420 3631 12472
rect 3683 12420 3739 12472
rect 3791 12420 3847 12472
rect 3899 12420 3911 12472
rect 3403 12364 3911 12420
rect 3403 12312 3415 12364
rect 3467 12312 3523 12364
rect 3575 12312 3631 12364
rect 3683 12312 3739 12364
rect 3791 12312 3847 12364
rect 3899 12312 3911 12364
rect 3403 12256 3911 12312
rect 3403 12204 3415 12256
rect 3467 12204 3523 12256
rect 3575 12204 3631 12256
rect 3683 12204 3739 12256
rect 3791 12204 3847 12256
rect 3899 12204 3911 12256
rect 3403 11068 3911 12204
rect 3403 11016 3415 11068
rect 3467 11016 3523 11068
rect 3575 11016 3631 11068
rect 3683 11016 3739 11068
rect 3791 11016 3847 11068
rect 3899 11016 3911 11068
rect 3403 10960 3911 11016
rect 3403 10908 3415 10960
rect 3467 10908 3523 10960
rect 3575 10908 3631 10960
rect 3683 10908 3739 10960
rect 3791 10908 3847 10960
rect 3899 10908 3911 10960
rect 3403 10852 3911 10908
rect 3403 10800 3415 10852
rect 3467 10800 3523 10852
rect 3575 10800 3631 10852
rect 3683 10800 3739 10852
rect 3791 10800 3847 10852
rect 3899 10800 3911 10852
rect 3403 9664 3911 10800
rect 3403 9612 3415 9664
rect 3467 9612 3523 9664
rect 3575 9612 3631 9664
rect 3683 9612 3739 9664
rect 3791 9612 3847 9664
rect 3899 9612 3911 9664
rect 3403 9556 3911 9612
rect 3403 9504 3415 9556
rect 3467 9504 3523 9556
rect 3575 9504 3631 9556
rect 3683 9504 3739 9556
rect 3791 9504 3847 9556
rect 3899 9504 3911 9556
rect 3403 9448 3911 9504
rect 3403 9396 3415 9448
rect 3467 9396 3523 9448
rect 3575 9396 3631 9448
rect 3683 9396 3739 9448
rect 3791 9396 3847 9448
rect 3899 9396 3911 9448
rect 3403 8283 3911 9396
rect 3403 8231 3415 8283
rect 3467 8231 3523 8283
rect 3575 8231 3631 8283
rect 3683 8231 3739 8283
rect 3791 8231 3847 8283
rect 3899 8231 3911 8283
rect 3403 8175 3911 8231
rect 3403 8123 3415 8175
rect 3467 8123 3523 8175
rect 3575 8123 3631 8175
rect 3683 8123 3739 8175
rect 3791 8123 3847 8175
rect 3899 8123 3911 8175
rect 3403 6989 3911 8123
rect 3403 6937 3445 6989
rect 3497 6937 3569 6989
rect 3621 6937 3693 6989
rect 3745 6937 3817 6989
rect 3869 6937 3911 6989
rect 3403 6865 3911 6937
rect 3403 6813 3445 6865
rect 3497 6813 3569 6865
rect 3621 6813 3693 6865
rect 3745 6813 3817 6865
rect 3869 6813 3911 6865
rect 3403 6741 3911 6813
rect 3403 6689 3445 6741
rect 3497 6689 3569 6741
rect 3621 6689 3693 6741
rect 3745 6689 3817 6741
rect 3869 6689 3911 6741
rect 3403 6617 3911 6689
rect 3403 6565 3445 6617
rect 3497 6565 3569 6617
rect 3621 6565 3693 6617
rect 3745 6565 3817 6617
rect 3869 6565 3911 6617
rect 3403 489 3911 6565
rect 3403 437 3445 489
rect 3497 437 3569 489
rect 3621 437 3693 489
rect 3745 437 3817 489
rect 3869 437 3911 489
rect 3403 365 3911 437
rect 3403 313 3445 365
rect 3497 313 3569 365
rect 3621 313 3693 365
rect 3745 313 3817 365
rect 3869 313 3911 365
rect 3403 241 3911 313
rect 3403 189 3445 241
rect 3497 189 3569 241
rect 3621 189 3693 241
rect 3745 189 3817 241
rect 3869 189 3911 241
rect 3403 117 3911 189
rect 3403 65 3445 117
rect 3497 65 3569 117
rect 3621 65 3693 117
rect 3745 65 3817 117
rect 3869 65 3911 117
rect 3403 43 3911 65
rect 3971 13314 4479 56440
rect 3971 13262 4013 13314
rect 4065 13262 4137 13314
rect 4189 13262 4261 13314
rect 4313 13262 4385 13314
rect 4437 13262 4479 13314
rect 3971 13190 4479 13262
rect 3971 13138 4013 13190
rect 4065 13138 4137 13190
rect 4189 13138 4261 13190
rect 4313 13138 4385 13190
rect 4437 13138 4479 13190
rect 3971 13066 4479 13138
rect 3971 13014 4013 13066
rect 4065 13014 4137 13066
rect 4189 13014 4261 13066
rect 4313 13014 4385 13066
rect 4437 13014 4479 13066
rect 3971 12942 4479 13014
rect 3971 12890 4013 12942
rect 4065 12890 4137 12942
rect 4189 12890 4261 12942
rect 4313 12890 4385 12942
rect 4437 12890 4479 12942
rect 3971 12818 4479 12890
rect 3971 12766 4013 12818
rect 4065 12766 4137 12818
rect 4189 12766 4261 12818
rect 4313 12766 4385 12818
rect 4437 12766 4479 12818
rect 3971 11910 4479 12766
rect 3971 11858 4013 11910
rect 4065 11858 4137 11910
rect 4189 11858 4261 11910
rect 4313 11858 4385 11910
rect 4437 11858 4479 11910
rect 3971 11786 4479 11858
rect 3971 11734 4013 11786
rect 4065 11734 4137 11786
rect 4189 11734 4261 11786
rect 4313 11734 4385 11786
rect 4437 11734 4479 11786
rect 3971 11662 4479 11734
rect 3971 11610 4013 11662
rect 4065 11610 4137 11662
rect 4189 11610 4261 11662
rect 4313 11610 4385 11662
rect 4437 11610 4479 11662
rect 3971 11538 4479 11610
rect 3971 11486 4013 11538
rect 4065 11486 4137 11538
rect 4189 11486 4261 11538
rect 4313 11486 4385 11538
rect 4437 11486 4479 11538
rect 3971 11414 4479 11486
rect 3971 11362 4013 11414
rect 4065 11362 4137 11414
rect 4189 11362 4261 11414
rect 4313 11362 4385 11414
rect 4437 11362 4479 11414
rect 3971 10506 4479 11362
rect 3971 10454 4013 10506
rect 4065 10454 4137 10506
rect 4189 10454 4261 10506
rect 4313 10454 4385 10506
rect 4437 10454 4479 10506
rect 3971 10382 4479 10454
rect 3971 10330 4013 10382
rect 4065 10330 4137 10382
rect 4189 10330 4261 10382
rect 4313 10330 4385 10382
rect 4437 10330 4479 10382
rect 3971 10258 4479 10330
rect 3971 10206 4013 10258
rect 4065 10206 4137 10258
rect 4189 10206 4261 10258
rect 4313 10206 4385 10258
rect 4437 10206 4479 10258
rect 3971 10134 4479 10206
rect 3971 10082 4013 10134
rect 4065 10082 4137 10134
rect 4189 10082 4261 10134
rect 4313 10082 4385 10134
rect 4437 10082 4479 10134
rect 3971 10010 4479 10082
rect 3971 9958 4013 10010
rect 4065 9958 4137 10010
rect 4189 9958 4261 10010
rect 4313 9958 4385 10010
rect 4437 9958 4479 10010
rect 3971 9102 4479 9958
rect 3971 9050 4013 9102
rect 4065 9050 4137 9102
rect 4189 9050 4261 9102
rect 4313 9050 4385 9102
rect 4437 9050 4479 9102
rect 3971 8978 4479 9050
rect 3971 8926 4013 8978
rect 4065 8926 4137 8978
rect 4189 8926 4261 8978
rect 4313 8926 4385 8978
rect 4437 8926 4479 8978
rect 3971 8854 4479 8926
rect 3971 8802 4013 8854
rect 4065 8802 4137 8854
rect 4189 8802 4261 8854
rect 4313 8802 4385 8854
rect 4437 8802 4479 8854
rect 3971 8730 4479 8802
rect 3971 8678 4013 8730
rect 4065 8678 4137 8730
rect 4189 8678 4261 8730
rect 4313 8678 4385 8730
rect 4437 8678 4479 8730
rect 3971 8606 4479 8678
rect 3971 8554 4013 8606
rect 4065 8554 4137 8606
rect 4189 8554 4261 8606
rect 4313 8554 4385 8606
rect 4437 8554 4479 8606
rect 3971 5907 4479 8554
rect 3971 5855 4013 5907
rect 4065 5855 4137 5907
rect 4189 5855 4261 5907
rect 4313 5855 4385 5907
rect 4437 5855 4479 5907
rect 3971 5783 4479 5855
rect 3971 5731 4013 5783
rect 4065 5731 4137 5783
rect 4189 5731 4261 5783
rect 4313 5731 4385 5783
rect 4437 5731 4479 5783
rect 3971 5659 4479 5731
rect 3971 5607 4013 5659
rect 4065 5607 4137 5659
rect 4189 5607 4261 5659
rect 4313 5607 4385 5659
rect 4437 5607 4479 5659
rect 3971 5535 4479 5607
rect 3971 5483 4013 5535
rect 4065 5483 4137 5535
rect 4189 5483 4261 5535
rect 4313 5483 4385 5535
rect 4437 5483 4479 5535
rect 3971 5411 4479 5483
rect 3971 5359 4013 5411
rect 4065 5359 4137 5411
rect 4189 5359 4261 5411
rect 4313 5359 4385 5411
rect 4437 5359 4479 5411
rect 3971 4503 4479 5359
rect 3971 4451 4013 4503
rect 4065 4451 4137 4503
rect 4189 4451 4261 4503
rect 4313 4451 4385 4503
rect 4437 4451 4479 4503
rect 3971 4379 4479 4451
rect 3971 4327 4013 4379
rect 4065 4327 4137 4379
rect 4189 4327 4261 4379
rect 4313 4327 4385 4379
rect 4437 4327 4479 4379
rect 3971 4255 4479 4327
rect 3971 4203 4013 4255
rect 4065 4203 4137 4255
rect 4189 4203 4261 4255
rect 4313 4203 4385 4255
rect 4437 4203 4479 4255
rect 3971 4131 4479 4203
rect 3971 4079 4013 4131
rect 4065 4079 4137 4131
rect 4189 4079 4261 4131
rect 4313 4079 4385 4131
rect 4437 4079 4479 4131
rect 3971 4007 4479 4079
rect 3971 3955 4013 4007
rect 4065 3955 4137 4007
rect 4189 3955 4261 4007
rect 4313 3955 4385 4007
rect 4437 3955 4479 4007
rect 3971 3099 4479 3955
rect 3971 3047 4013 3099
rect 4065 3047 4137 3099
rect 4189 3047 4261 3099
rect 4313 3047 4385 3099
rect 4437 3047 4479 3099
rect 3971 2975 4479 3047
rect 3971 2923 4013 2975
rect 4065 2923 4137 2975
rect 4189 2923 4261 2975
rect 4313 2923 4385 2975
rect 4437 2923 4479 2975
rect 3971 2851 4479 2923
rect 3971 2799 4013 2851
rect 4065 2799 4137 2851
rect 4189 2799 4261 2851
rect 4313 2799 4385 2851
rect 4437 2799 4479 2851
rect 3971 2727 4479 2799
rect 3971 2675 4013 2727
rect 4065 2675 4137 2727
rect 4189 2675 4261 2727
rect 4313 2675 4385 2727
rect 4437 2675 4479 2727
rect 3971 2603 4479 2675
rect 3971 2551 4013 2603
rect 4065 2551 4137 2603
rect 4189 2551 4261 2603
rect 4313 2551 4385 2603
rect 4437 2551 4479 2603
rect 3971 1695 4479 2551
rect 3971 1643 4013 1695
rect 4065 1643 4137 1695
rect 4189 1643 4261 1695
rect 4313 1643 4385 1695
rect 4437 1643 4479 1695
rect 3971 1571 4479 1643
rect 3971 1519 4013 1571
rect 4065 1519 4137 1571
rect 4189 1519 4261 1571
rect 4313 1519 4385 1571
rect 4437 1519 4479 1571
rect 3971 1447 4479 1519
rect 3971 1395 4013 1447
rect 4065 1395 4137 1447
rect 4189 1395 4261 1447
rect 4313 1395 4385 1447
rect 4437 1395 4479 1447
rect 3971 1323 4479 1395
rect 3971 1271 4013 1323
rect 4065 1271 4137 1323
rect 4189 1271 4261 1323
rect 4313 1271 4385 1323
rect 4437 1271 4479 1323
rect 3971 1199 4479 1271
rect 3971 1147 4013 1199
rect 4065 1147 4137 1199
rect 4189 1147 4261 1199
rect 4313 1147 4385 1199
rect 4437 1147 4479 1199
rect 3971 -857 4479 1147
rect 4539 14396 5047 14905
rect 4539 14344 4581 14396
rect 4633 14344 4705 14396
rect 4757 14344 4829 14396
rect 4881 14344 4953 14396
rect 5005 14344 5047 14396
rect 4539 14272 5047 14344
rect 4539 14220 4581 14272
rect 4633 14220 4705 14272
rect 4757 14220 4829 14272
rect 4881 14220 4953 14272
rect 5005 14220 5047 14272
rect 4539 14148 5047 14220
rect 4539 14096 4581 14148
rect 4633 14096 4705 14148
rect 4757 14096 4829 14148
rect 4881 14096 4953 14148
rect 5005 14096 5047 14148
rect 4539 14024 5047 14096
rect 4539 13972 4581 14024
rect 4633 13972 4705 14024
rect 4757 13972 4829 14024
rect 4881 13972 4953 14024
rect 5005 13972 5047 14024
rect 4539 7896 5047 13972
rect 4539 7844 4581 7896
rect 4633 7844 4705 7896
rect 4757 7844 4829 7896
rect 4881 7844 4953 7896
rect 5005 7844 5047 7896
rect 4539 7772 5047 7844
rect 4539 7720 4581 7772
rect 4633 7720 4705 7772
rect 4757 7720 4829 7772
rect 4881 7720 4953 7772
rect 5005 7720 5047 7772
rect 4539 7648 5047 7720
rect 4539 7596 4581 7648
rect 4633 7596 4705 7648
rect 4757 7596 4829 7648
rect 4881 7596 4953 7648
rect 5005 7596 5047 7648
rect 4539 7524 5047 7596
rect 4539 7472 4581 7524
rect 4633 7472 4705 7524
rect 4757 7472 4829 7524
rect 4881 7472 4953 7524
rect 5005 7472 5047 7524
rect 4539 6338 5047 7472
rect 4539 6286 4551 6338
rect 4603 6286 4659 6338
rect 4711 6286 4767 6338
rect 4819 6286 4875 6338
rect 4927 6286 4983 6338
rect 5035 6286 5047 6338
rect 4539 6230 5047 6286
rect 4539 6178 4551 6230
rect 4603 6178 4659 6230
rect 4711 6178 4767 6230
rect 4819 6178 4875 6230
rect 4927 6178 4983 6230
rect 5035 6178 5047 6230
rect 4539 5065 5047 6178
rect 4539 5013 4551 5065
rect 4603 5013 4659 5065
rect 4711 5013 4767 5065
rect 4819 5013 4875 5065
rect 4927 5013 4983 5065
rect 5035 5013 5047 5065
rect 4539 4957 5047 5013
rect 4539 4905 4551 4957
rect 4603 4905 4659 4957
rect 4711 4905 4767 4957
rect 4819 4905 4875 4957
rect 4927 4905 4983 4957
rect 5035 4905 5047 4957
rect 4539 4849 5047 4905
rect 4539 4797 4551 4849
rect 4603 4797 4659 4849
rect 4711 4797 4767 4849
rect 4819 4797 4875 4849
rect 4927 4797 4983 4849
rect 5035 4797 5047 4849
rect 4539 3661 5047 4797
rect 4539 3609 4551 3661
rect 4603 3609 4659 3661
rect 4711 3609 4767 3661
rect 4819 3609 4875 3661
rect 4927 3609 4983 3661
rect 5035 3609 5047 3661
rect 4539 3553 5047 3609
rect 4539 3501 4551 3553
rect 4603 3501 4659 3553
rect 4711 3501 4767 3553
rect 4819 3501 4875 3553
rect 4927 3501 4983 3553
rect 5035 3501 5047 3553
rect 4539 3445 5047 3501
rect 4539 3393 4551 3445
rect 4603 3393 4659 3445
rect 4711 3393 4767 3445
rect 4819 3393 4875 3445
rect 4927 3393 4983 3445
rect 5035 3393 5047 3445
rect 4539 2257 5047 3393
rect 4539 2205 4551 2257
rect 4603 2205 4659 2257
rect 4711 2205 4767 2257
rect 4819 2205 4875 2257
rect 4927 2205 4983 2257
rect 5035 2205 5047 2257
rect 4539 2149 5047 2205
rect 4539 2097 4551 2149
rect 4603 2097 4659 2149
rect 4711 2097 4767 2149
rect 4819 2097 4875 2149
rect 4927 2097 4983 2149
rect 5035 2097 5047 2149
rect 4539 2041 5047 2097
rect 4539 1989 4551 2041
rect 4603 1989 4659 2041
rect 4711 1989 4767 2041
rect 4819 1989 4875 2041
rect 4927 1989 4983 2041
rect 5035 1989 5047 2041
rect 4539 876 5047 1989
rect 4539 824 4551 876
rect 4603 824 4659 876
rect 4711 824 4767 876
rect 4819 824 4875 876
rect 4927 824 4983 876
rect 5035 824 5047 876
rect 4539 768 5047 824
rect 4539 716 4551 768
rect 4603 716 4659 768
rect 4711 716 4767 768
rect 4819 716 4875 768
rect 4927 716 4983 768
rect 5035 716 5047 768
rect 4539 43 5047 716
rect 5107 13314 5615 56440
rect 5107 13262 5149 13314
rect 5201 13262 5273 13314
rect 5325 13262 5397 13314
rect 5449 13262 5521 13314
rect 5573 13262 5615 13314
rect 5107 13190 5615 13262
rect 5107 13138 5149 13190
rect 5201 13138 5273 13190
rect 5325 13138 5397 13190
rect 5449 13138 5521 13190
rect 5573 13138 5615 13190
rect 5107 13066 5615 13138
rect 5107 13014 5149 13066
rect 5201 13014 5273 13066
rect 5325 13014 5397 13066
rect 5449 13014 5521 13066
rect 5573 13014 5615 13066
rect 5107 12942 5615 13014
rect 5107 12890 5149 12942
rect 5201 12890 5273 12942
rect 5325 12890 5397 12942
rect 5449 12890 5521 12942
rect 5573 12890 5615 12942
rect 5107 12818 5615 12890
rect 5107 12766 5149 12818
rect 5201 12766 5273 12818
rect 5325 12766 5397 12818
rect 5449 12766 5521 12818
rect 5573 12766 5615 12818
rect 5107 11910 5615 12766
rect 5107 11858 5149 11910
rect 5201 11858 5273 11910
rect 5325 11858 5397 11910
rect 5449 11858 5521 11910
rect 5573 11858 5615 11910
rect 5107 11786 5615 11858
rect 5107 11734 5149 11786
rect 5201 11734 5273 11786
rect 5325 11734 5397 11786
rect 5449 11734 5521 11786
rect 5573 11734 5615 11786
rect 5107 11662 5615 11734
rect 5107 11610 5149 11662
rect 5201 11610 5273 11662
rect 5325 11610 5397 11662
rect 5449 11610 5521 11662
rect 5573 11610 5615 11662
rect 5107 11538 5615 11610
rect 5107 11486 5149 11538
rect 5201 11486 5273 11538
rect 5325 11486 5397 11538
rect 5449 11486 5521 11538
rect 5573 11486 5615 11538
rect 5107 11414 5615 11486
rect 5107 11362 5149 11414
rect 5201 11362 5273 11414
rect 5325 11362 5397 11414
rect 5449 11362 5521 11414
rect 5573 11362 5615 11414
rect 5107 10506 5615 11362
rect 5107 10454 5149 10506
rect 5201 10454 5273 10506
rect 5325 10454 5397 10506
rect 5449 10454 5521 10506
rect 5573 10454 5615 10506
rect 5107 10382 5615 10454
rect 5107 10330 5149 10382
rect 5201 10330 5273 10382
rect 5325 10330 5397 10382
rect 5449 10330 5521 10382
rect 5573 10330 5615 10382
rect 5107 10258 5615 10330
rect 5107 10206 5149 10258
rect 5201 10206 5273 10258
rect 5325 10206 5397 10258
rect 5449 10206 5521 10258
rect 5573 10206 5615 10258
rect 5107 10134 5615 10206
rect 5107 10082 5149 10134
rect 5201 10082 5273 10134
rect 5325 10082 5397 10134
rect 5449 10082 5521 10134
rect 5573 10082 5615 10134
rect 5107 10010 5615 10082
rect 5107 9958 5149 10010
rect 5201 9958 5273 10010
rect 5325 9958 5397 10010
rect 5449 9958 5521 10010
rect 5573 9958 5615 10010
rect 5107 9102 5615 9958
rect 5107 9050 5149 9102
rect 5201 9050 5273 9102
rect 5325 9050 5397 9102
rect 5449 9050 5521 9102
rect 5573 9050 5615 9102
rect 5107 8978 5615 9050
rect 5107 8926 5149 8978
rect 5201 8926 5273 8978
rect 5325 8926 5397 8978
rect 5449 8926 5521 8978
rect 5573 8926 5615 8978
rect 5107 8854 5615 8926
rect 5107 8802 5149 8854
rect 5201 8802 5273 8854
rect 5325 8802 5397 8854
rect 5449 8802 5521 8854
rect 5573 8802 5615 8854
rect 5107 8730 5615 8802
rect 5107 8678 5149 8730
rect 5201 8678 5273 8730
rect 5325 8678 5397 8730
rect 5449 8678 5521 8730
rect 5573 8678 5615 8730
rect 5107 8606 5615 8678
rect 5107 8554 5149 8606
rect 5201 8554 5273 8606
rect 5325 8554 5397 8606
rect 5449 8554 5521 8606
rect 5573 8554 5615 8606
rect 5107 5907 5615 8554
rect 5107 5855 5149 5907
rect 5201 5855 5273 5907
rect 5325 5855 5397 5907
rect 5449 5855 5521 5907
rect 5573 5855 5615 5907
rect 5107 5783 5615 5855
rect 5107 5731 5149 5783
rect 5201 5731 5273 5783
rect 5325 5731 5397 5783
rect 5449 5731 5521 5783
rect 5573 5731 5615 5783
rect 5107 5659 5615 5731
rect 5107 5607 5149 5659
rect 5201 5607 5273 5659
rect 5325 5607 5397 5659
rect 5449 5607 5521 5659
rect 5573 5607 5615 5659
rect 5107 5535 5615 5607
rect 5107 5483 5149 5535
rect 5201 5483 5273 5535
rect 5325 5483 5397 5535
rect 5449 5483 5521 5535
rect 5573 5483 5615 5535
rect 5107 5411 5615 5483
rect 5107 5359 5149 5411
rect 5201 5359 5273 5411
rect 5325 5359 5397 5411
rect 5449 5359 5521 5411
rect 5573 5359 5615 5411
rect 5107 4503 5615 5359
rect 5107 4451 5149 4503
rect 5201 4451 5273 4503
rect 5325 4451 5397 4503
rect 5449 4451 5521 4503
rect 5573 4451 5615 4503
rect 5107 4379 5615 4451
rect 5107 4327 5149 4379
rect 5201 4327 5273 4379
rect 5325 4327 5397 4379
rect 5449 4327 5521 4379
rect 5573 4327 5615 4379
rect 5107 4255 5615 4327
rect 5107 4203 5149 4255
rect 5201 4203 5273 4255
rect 5325 4203 5397 4255
rect 5449 4203 5521 4255
rect 5573 4203 5615 4255
rect 5107 4131 5615 4203
rect 5107 4079 5149 4131
rect 5201 4079 5273 4131
rect 5325 4079 5397 4131
rect 5449 4079 5521 4131
rect 5573 4079 5615 4131
rect 5107 4007 5615 4079
rect 5107 3955 5149 4007
rect 5201 3955 5273 4007
rect 5325 3955 5397 4007
rect 5449 3955 5521 4007
rect 5573 3955 5615 4007
rect 5107 3099 5615 3955
rect 5107 3047 5149 3099
rect 5201 3047 5273 3099
rect 5325 3047 5397 3099
rect 5449 3047 5521 3099
rect 5573 3047 5615 3099
rect 5107 2975 5615 3047
rect 5107 2923 5149 2975
rect 5201 2923 5273 2975
rect 5325 2923 5397 2975
rect 5449 2923 5521 2975
rect 5573 2923 5615 2975
rect 5107 2851 5615 2923
rect 5107 2799 5149 2851
rect 5201 2799 5273 2851
rect 5325 2799 5397 2851
rect 5449 2799 5521 2851
rect 5573 2799 5615 2851
rect 5107 2727 5615 2799
rect 5107 2675 5149 2727
rect 5201 2675 5273 2727
rect 5325 2675 5397 2727
rect 5449 2675 5521 2727
rect 5573 2675 5615 2727
rect 5107 2603 5615 2675
rect 5107 2551 5149 2603
rect 5201 2551 5273 2603
rect 5325 2551 5397 2603
rect 5449 2551 5521 2603
rect 5573 2551 5615 2603
rect 5107 1695 5615 2551
rect 5107 1643 5149 1695
rect 5201 1643 5273 1695
rect 5325 1643 5397 1695
rect 5449 1643 5521 1695
rect 5573 1643 5615 1695
rect 5107 1571 5615 1643
rect 5107 1519 5149 1571
rect 5201 1519 5273 1571
rect 5325 1519 5397 1571
rect 5449 1519 5521 1571
rect 5573 1519 5615 1571
rect 5107 1447 5615 1519
rect 5107 1395 5149 1447
rect 5201 1395 5273 1447
rect 5325 1395 5397 1447
rect 5449 1395 5521 1447
rect 5573 1395 5615 1447
rect 5107 1323 5615 1395
rect 5107 1271 5149 1323
rect 5201 1271 5273 1323
rect 5325 1271 5397 1323
rect 5449 1271 5521 1323
rect 5573 1271 5615 1323
rect 5107 1199 5615 1271
rect 5107 1147 5149 1199
rect 5201 1147 5273 1199
rect 5325 1147 5397 1199
rect 5449 1147 5521 1199
rect 5573 1147 5615 1199
rect 5107 -857 5615 1147
rect 5675 13745 6101 14905
rect 5675 13693 5700 13745
rect 5752 13693 5808 13745
rect 5860 13693 5916 13745
rect 5968 13693 6024 13745
rect 6076 13693 6101 13745
rect 5675 13637 6101 13693
rect 5675 13585 5700 13637
rect 5752 13585 5808 13637
rect 5860 13585 5916 13637
rect 5968 13585 6024 13637
rect 6076 13585 6101 13637
rect 5675 12472 6101 13585
rect 5675 12420 5700 12472
rect 5752 12420 5808 12472
rect 5860 12420 5916 12472
rect 5968 12420 6024 12472
rect 6076 12420 6101 12472
rect 5675 12364 6101 12420
rect 5675 12312 5700 12364
rect 5752 12312 5808 12364
rect 5860 12312 5916 12364
rect 5968 12312 6024 12364
rect 6076 12312 6101 12364
rect 5675 12256 6101 12312
rect 5675 12204 5700 12256
rect 5752 12204 5808 12256
rect 5860 12204 5916 12256
rect 5968 12204 6024 12256
rect 6076 12204 6101 12256
rect 5675 11068 6101 12204
rect 5675 11016 5700 11068
rect 5752 11016 5808 11068
rect 5860 11016 5916 11068
rect 5968 11016 6024 11068
rect 6076 11016 6101 11068
rect 5675 10960 6101 11016
rect 5675 10908 5700 10960
rect 5752 10908 5808 10960
rect 5860 10908 5916 10960
rect 5968 10908 6024 10960
rect 6076 10908 6101 10960
rect 5675 10852 6101 10908
rect 5675 10800 5700 10852
rect 5752 10800 5808 10852
rect 5860 10800 5916 10852
rect 5968 10800 6024 10852
rect 6076 10800 6101 10852
rect 5675 9664 6101 10800
rect 5675 9612 5700 9664
rect 5752 9612 5808 9664
rect 5860 9612 5916 9664
rect 5968 9612 6024 9664
rect 6076 9612 6101 9664
rect 5675 9556 6101 9612
rect 5675 9504 5700 9556
rect 5752 9504 5808 9556
rect 5860 9504 5916 9556
rect 5968 9504 6024 9556
rect 6076 9504 6101 9556
rect 5675 9448 6101 9504
rect 5675 9396 5700 9448
rect 5752 9396 5808 9448
rect 5860 9396 5916 9448
rect 5968 9396 6024 9448
rect 6076 9396 6101 9448
rect 5675 8283 6101 9396
rect 5675 8231 5700 8283
rect 5752 8231 5808 8283
rect 5860 8231 5916 8283
rect 5968 8231 6024 8283
rect 6076 8231 6101 8283
rect 5675 8175 6101 8231
rect 5675 8123 5700 8175
rect 5752 8123 5808 8175
rect 5860 8123 5916 8175
rect 5968 8123 6024 8175
rect 6076 8123 6101 8175
rect 5675 6989 6101 8123
rect 5675 6937 5738 6989
rect 5790 6937 5862 6989
rect 5914 6937 5986 6989
rect 6038 6937 6101 6989
rect 5675 6865 6101 6937
rect 5675 6813 5738 6865
rect 5790 6813 5862 6865
rect 5914 6813 5986 6865
rect 6038 6813 6101 6865
rect 5675 6741 6101 6813
rect 5675 6689 5738 6741
rect 5790 6689 5862 6741
rect 5914 6689 5986 6741
rect 6038 6689 6101 6741
rect 5675 6617 6101 6689
rect 5675 6565 5738 6617
rect 5790 6565 5862 6617
rect 5914 6565 5986 6617
rect 6038 6565 6101 6617
rect 5675 489 6101 6565
rect 5675 437 5738 489
rect 5790 437 5862 489
rect 5914 437 5986 489
rect 6038 437 6101 489
rect 5675 365 6101 437
rect 5675 313 5738 365
rect 5790 313 5862 365
rect 5914 313 5986 365
rect 6038 313 6101 365
rect 5675 241 6101 313
rect 5675 189 5738 241
rect 5790 189 5862 241
rect 5914 189 5986 241
rect 6038 189 6101 241
rect 5675 117 6101 189
rect 5675 65 5738 117
rect 5790 65 5862 117
rect 5914 65 5986 117
rect 6038 65 6101 117
rect 5675 43 6101 65
rect 6161 13745 6587 14905
rect 6161 13693 6186 13745
rect 6238 13693 6294 13745
rect 6346 13693 6402 13745
rect 6454 13693 6510 13745
rect 6562 13693 6587 13745
rect 6161 13637 6587 13693
rect 6161 13585 6186 13637
rect 6238 13585 6294 13637
rect 6346 13585 6402 13637
rect 6454 13585 6510 13637
rect 6562 13585 6587 13637
rect 6161 12472 6587 13585
rect 6161 12420 6186 12472
rect 6238 12420 6294 12472
rect 6346 12420 6402 12472
rect 6454 12420 6510 12472
rect 6562 12420 6587 12472
rect 6161 12364 6587 12420
rect 6161 12312 6186 12364
rect 6238 12312 6294 12364
rect 6346 12312 6402 12364
rect 6454 12312 6510 12364
rect 6562 12312 6587 12364
rect 6161 12256 6587 12312
rect 6161 12204 6186 12256
rect 6238 12204 6294 12256
rect 6346 12204 6402 12256
rect 6454 12204 6510 12256
rect 6562 12204 6587 12256
rect 6161 11068 6587 12204
rect 6161 11016 6186 11068
rect 6238 11016 6294 11068
rect 6346 11016 6402 11068
rect 6454 11016 6510 11068
rect 6562 11016 6587 11068
rect 6161 10960 6587 11016
rect 6161 10908 6186 10960
rect 6238 10908 6294 10960
rect 6346 10908 6402 10960
rect 6454 10908 6510 10960
rect 6562 10908 6587 10960
rect 6161 10852 6587 10908
rect 6161 10800 6186 10852
rect 6238 10800 6294 10852
rect 6346 10800 6402 10852
rect 6454 10800 6510 10852
rect 6562 10800 6587 10852
rect 6161 9664 6587 10800
rect 6161 9612 6186 9664
rect 6238 9612 6294 9664
rect 6346 9612 6402 9664
rect 6454 9612 6510 9664
rect 6562 9612 6587 9664
rect 6161 9556 6587 9612
rect 6161 9504 6186 9556
rect 6238 9504 6294 9556
rect 6346 9504 6402 9556
rect 6454 9504 6510 9556
rect 6562 9504 6587 9556
rect 6161 9448 6587 9504
rect 6161 9396 6186 9448
rect 6238 9396 6294 9448
rect 6346 9396 6402 9448
rect 6454 9396 6510 9448
rect 6562 9396 6587 9448
rect 6161 8283 6587 9396
rect 6161 8231 6186 8283
rect 6238 8231 6294 8283
rect 6346 8231 6402 8283
rect 6454 8231 6510 8283
rect 6562 8231 6587 8283
rect 6161 8175 6587 8231
rect 6161 8123 6186 8175
rect 6238 8123 6294 8175
rect 6346 8123 6402 8175
rect 6454 8123 6510 8175
rect 6562 8123 6587 8175
rect 6161 6989 6587 8123
rect 6161 6937 6224 6989
rect 6276 6937 6348 6989
rect 6400 6937 6472 6989
rect 6524 6937 6587 6989
rect 6161 6865 6587 6937
rect 6161 6813 6224 6865
rect 6276 6813 6348 6865
rect 6400 6813 6472 6865
rect 6524 6813 6587 6865
rect 6161 6741 6587 6813
rect 6161 6689 6224 6741
rect 6276 6689 6348 6741
rect 6400 6689 6472 6741
rect 6524 6689 6587 6741
rect 6161 6617 6587 6689
rect 6161 6565 6224 6617
rect 6276 6565 6348 6617
rect 6400 6565 6472 6617
rect 6524 6565 6587 6617
rect 6161 489 6587 6565
rect 6161 437 6224 489
rect 6276 437 6348 489
rect 6400 437 6472 489
rect 6524 437 6587 489
rect 6161 365 6587 437
rect 6161 313 6224 365
rect 6276 313 6348 365
rect 6400 313 6472 365
rect 6524 313 6587 365
rect 6161 241 6587 313
rect 6161 189 6224 241
rect 6276 189 6348 241
rect 6400 189 6472 241
rect 6524 189 6587 241
rect 6161 117 6587 189
rect 6161 65 6224 117
rect 6276 65 6348 117
rect 6400 65 6472 117
rect 6524 65 6587 117
rect 6161 43 6587 65
rect 6647 13314 7155 56440
rect 6647 13262 6689 13314
rect 6741 13262 6813 13314
rect 6865 13262 6937 13314
rect 6989 13262 7061 13314
rect 7113 13262 7155 13314
rect 6647 13190 7155 13262
rect 6647 13138 6689 13190
rect 6741 13138 6813 13190
rect 6865 13138 6937 13190
rect 6989 13138 7061 13190
rect 7113 13138 7155 13190
rect 6647 13066 7155 13138
rect 6647 13014 6689 13066
rect 6741 13014 6813 13066
rect 6865 13014 6937 13066
rect 6989 13014 7061 13066
rect 7113 13014 7155 13066
rect 6647 12942 7155 13014
rect 6647 12890 6689 12942
rect 6741 12890 6813 12942
rect 6865 12890 6937 12942
rect 6989 12890 7061 12942
rect 7113 12890 7155 12942
rect 6647 12818 7155 12890
rect 6647 12766 6689 12818
rect 6741 12766 6813 12818
rect 6865 12766 6937 12818
rect 6989 12766 7061 12818
rect 7113 12766 7155 12818
rect 6647 11910 7155 12766
rect 6647 11858 6689 11910
rect 6741 11858 6813 11910
rect 6865 11858 6937 11910
rect 6989 11858 7061 11910
rect 7113 11858 7155 11910
rect 6647 11786 7155 11858
rect 6647 11734 6689 11786
rect 6741 11734 6813 11786
rect 6865 11734 6937 11786
rect 6989 11734 7061 11786
rect 7113 11734 7155 11786
rect 6647 11662 7155 11734
rect 6647 11610 6689 11662
rect 6741 11610 6813 11662
rect 6865 11610 6937 11662
rect 6989 11610 7061 11662
rect 7113 11610 7155 11662
rect 6647 11538 7155 11610
rect 6647 11486 6689 11538
rect 6741 11486 6813 11538
rect 6865 11486 6937 11538
rect 6989 11486 7061 11538
rect 7113 11486 7155 11538
rect 6647 11414 7155 11486
rect 6647 11362 6689 11414
rect 6741 11362 6813 11414
rect 6865 11362 6937 11414
rect 6989 11362 7061 11414
rect 7113 11362 7155 11414
rect 6647 10506 7155 11362
rect 6647 10454 6689 10506
rect 6741 10454 6813 10506
rect 6865 10454 6937 10506
rect 6989 10454 7061 10506
rect 7113 10454 7155 10506
rect 6647 10382 7155 10454
rect 6647 10330 6689 10382
rect 6741 10330 6813 10382
rect 6865 10330 6937 10382
rect 6989 10330 7061 10382
rect 7113 10330 7155 10382
rect 6647 10258 7155 10330
rect 6647 10206 6689 10258
rect 6741 10206 6813 10258
rect 6865 10206 6937 10258
rect 6989 10206 7061 10258
rect 7113 10206 7155 10258
rect 6647 10134 7155 10206
rect 6647 10082 6689 10134
rect 6741 10082 6813 10134
rect 6865 10082 6937 10134
rect 6989 10082 7061 10134
rect 7113 10082 7155 10134
rect 6647 10010 7155 10082
rect 6647 9958 6689 10010
rect 6741 9958 6813 10010
rect 6865 9958 6937 10010
rect 6989 9958 7061 10010
rect 7113 9958 7155 10010
rect 6647 9102 7155 9958
rect 6647 9050 6689 9102
rect 6741 9050 6813 9102
rect 6865 9050 6937 9102
rect 6989 9050 7061 9102
rect 7113 9050 7155 9102
rect 6647 8978 7155 9050
rect 6647 8926 6689 8978
rect 6741 8926 6813 8978
rect 6865 8926 6937 8978
rect 6989 8926 7061 8978
rect 7113 8926 7155 8978
rect 6647 8854 7155 8926
rect 6647 8802 6689 8854
rect 6741 8802 6813 8854
rect 6865 8802 6937 8854
rect 6989 8802 7061 8854
rect 7113 8802 7155 8854
rect 6647 8730 7155 8802
rect 6647 8678 6689 8730
rect 6741 8678 6813 8730
rect 6865 8678 6937 8730
rect 6989 8678 7061 8730
rect 7113 8678 7155 8730
rect 6647 8606 7155 8678
rect 6647 8554 6689 8606
rect 6741 8554 6813 8606
rect 6865 8554 6937 8606
rect 6989 8554 7061 8606
rect 7113 8554 7155 8606
rect 6647 5907 7155 8554
rect 6647 5855 6689 5907
rect 6741 5855 6813 5907
rect 6865 5855 6937 5907
rect 6989 5855 7061 5907
rect 7113 5855 7155 5907
rect 6647 5783 7155 5855
rect 6647 5731 6689 5783
rect 6741 5731 6813 5783
rect 6865 5731 6937 5783
rect 6989 5731 7061 5783
rect 7113 5731 7155 5783
rect 6647 5659 7155 5731
rect 6647 5607 6689 5659
rect 6741 5607 6813 5659
rect 6865 5607 6937 5659
rect 6989 5607 7061 5659
rect 7113 5607 7155 5659
rect 6647 5535 7155 5607
rect 6647 5483 6689 5535
rect 6741 5483 6813 5535
rect 6865 5483 6937 5535
rect 6989 5483 7061 5535
rect 7113 5483 7155 5535
rect 6647 5411 7155 5483
rect 6647 5359 6689 5411
rect 6741 5359 6813 5411
rect 6865 5359 6937 5411
rect 6989 5359 7061 5411
rect 7113 5359 7155 5411
rect 6647 4503 7155 5359
rect 6647 4451 6689 4503
rect 6741 4451 6813 4503
rect 6865 4451 6937 4503
rect 6989 4451 7061 4503
rect 7113 4451 7155 4503
rect 6647 4379 7155 4451
rect 6647 4327 6689 4379
rect 6741 4327 6813 4379
rect 6865 4327 6937 4379
rect 6989 4327 7061 4379
rect 7113 4327 7155 4379
rect 6647 4255 7155 4327
rect 6647 4203 6689 4255
rect 6741 4203 6813 4255
rect 6865 4203 6937 4255
rect 6989 4203 7061 4255
rect 7113 4203 7155 4255
rect 6647 4131 7155 4203
rect 6647 4079 6689 4131
rect 6741 4079 6813 4131
rect 6865 4079 6937 4131
rect 6989 4079 7061 4131
rect 7113 4079 7155 4131
rect 6647 4007 7155 4079
rect 6647 3955 6689 4007
rect 6741 3955 6813 4007
rect 6865 3955 6937 4007
rect 6989 3955 7061 4007
rect 7113 3955 7155 4007
rect 6647 3099 7155 3955
rect 6647 3047 6689 3099
rect 6741 3047 6813 3099
rect 6865 3047 6937 3099
rect 6989 3047 7061 3099
rect 7113 3047 7155 3099
rect 6647 2975 7155 3047
rect 6647 2923 6689 2975
rect 6741 2923 6813 2975
rect 6865 2923 6937 2975
rect 6989 2923 7061 2975
rect 7113 2923 7155 2975
rect 6647 2851 7155 2923
rect 6647 2799 6689 2851
rect 6741 2799 6813 2851
rect 6865 2799 6937 2851
rect 6989 2799 7061 2851
rect 7113 2799 7155 2851
rect 6647 2727 7155 2799
rect 6647 2675 6689 2727
rect 6741 2675 6813 2727
rect 6865 2675 6937 2727
rect 6989 2675 7061 2727
rect 7113 2675 7155 2727
rect 6647 2603 7155 2675
rect 6647 2551 6689 2603
rect 6741 2551 6813 2603
rect 6865 2551 6937 2603
rect 6989 2551 7061 2603
rect 7113 2551 7155 2603
rect 6647 1695 7155 2551
rect 6647 1643 6689 1695
rect 6741 1643 6813 1695
rect 6865 1643 6937 1695
rect 6989 1643 7061 1695
rect 7113 1643 7155 1695
rect 6647 1571 7155 1643
rect 6647 1519 6689 1571
rect 6741 1519 6813 1571
rect 6865 1519 6937 1571
rect 6989 1519 7061 1571
rect 7113 1519 7155 1571
rect 6647 1447 7155 1519
rect 6647 1395 6689 1447
rect 6741 1395 6813 1447
rect 6865 1395 6937 1447
rect 6989 1395 7061 1447
rect 7113 1395 7155 1447
rect 6647 1323 7155 1395
rect 6647 1271 6689 1323
rect 6741 1271 6813 1323
rect 6865 1271 6937 1323
rect 6989 1271 7061 1323
rect 7113 1271 7155 1323
rect 6647 1199 7155 1271
rect 6647 1147 6689 1199
rect 6741 1147 6813 1199
rect 6865 1147 6937 1199
rect 6989 1147 7061 1199
rect 7113 1147 7155 1199
rect 6647 -857 7155 1147
rect 7215 14396 7723 14905
rect 7215 14344 7257 14396
rect 7309 14344 7381 14396
rect 7433 14344 7505 14396
rect 7557 14344 7629 14396
rect 7681 14344 7723 14396
rect 7215 14272 7723 14344
rect 7215 14220 7257 14272
rect 7309 14220 7381 14272
rect 7433 14220 7505 14272
rect 7557 14220 7629 14272
rect 7681 14220 7723 14272
rect 7215 14148 7723 14220
rect 7215 14096 7257 14148
rect 7309 14096 7381 14148
rect 7433 14096 7505 14148
rect 7557 14096 7629 14148
rect 7681 14096 7723 14148
rect 7215 14024 7723 14096
rect 7215 13972 7257 14024
rect 7309 13972 7381 14024
rect 7433 13972 7505 14024
rect 7557 13972 7629 14024
rect 7681 13972 7723 14024
rect 7215 7896 7723 13972
rect 7215 7844 7257 7896
rect 7309 7844 7381 7896
rect 7433 7844 7505 7896
rect 7557 7844 7629 7896
rect 7681 7844 7723 7896
rect 7215 7772 7723 7844
rect 7215 7720 7257 7772
rect 7309 7720 7381 7772
rect 7433 7720 7505 7772
rect 7557 7720 7629 7772
rect 7681 7720 7723 7772
rect 7215 7648 7723 7720
rect 7215 7596 7257 7648
rect 7309 7596 7381 7648
rect 7433 7596 7505 7648
rect 7557 7596 7629 7648
rect 7681 7596 7723 7648
rect 7215 7524 7723 7596
rect 7215 7472 7257 7524
rect 7309 7472 7381 7524
rect 7433 7472 7505 7524
rect 7557 7472 7629 7524
rect 7681 7472 7723 7524
rect 7215 6338 7723 7472
rect 7215 6286 7227 6338
rect 7279 6286 7335 6338
rect 7387 6286 7443 6338
rect 7495 6286 7551 6338
rect 7603 6286 7659 6338
rect 7711 6286 7723 6338
rect 7215 6230 7723 6286
rect 7215 6178 7227 6230
rect 7279 6178 7335 6230
rect 7387 6178 7443 6230
rect 7495 6178 7551 6230
rect 7603 6178 7659 6230
rect 7711 6178 7723 6230
rect 7215 5065 7723 6178
rect 7215 5013 7227 5065
rect 7279 5013 7335 5065
rect 7387 5013 7443 5065
rect 7495 5013 7551 5065
rect 7603 5013 7659 5065
rect 7711 5013 7723 5065
rect 7215 4957 7723 5013
rect 7215 4905 7227 4957
rect 7279 4905 7335 4957
rect 7387 4905 7443 4957
rect 7495 4905 7551 4957
rect 7603 4905 7659 4957
rect 7711 4905 7723 4957
rect 7215 4849 7723 4905
rect 7215 4797 7227 4849
rect 7279 4797 7335 4849
rect 7387 4797 7443 4849
rect 7495 4797 7551 4849
rect 7603 4797 7659 4849
rect 7711 4797 7723 4849
rect 7215 3661 7723 4797
rect 7215 3609 7227 3661
rect 7279 3609 7335 3661
rect 7387 3609 7443 3661
rect 7495 3609 7551 3661
rect 7603 3609 7659 3661
rect 7711 3609 7723 3661
rect 7215 3553 7723 3609
rect 7215 3501 7227 3553
rect 7279 3501 7335 3553
rect 7387 3501 7443 3553
rect 7495 3501 7551 3553
rect 7603 3501 7659 3553
rect 7711 3501 7723 3553
rect 7215 3445 7723 3501
rect 7215 3393 7227 3445
rect 7279 3393 7335 3445
rect 7387 3393 7443 3445
rect 7495 3393 7551 3445
rect 7603 3393 7659 3445
rect 7711 3393 7723 3445
rect 7215 2257 7723 3393
rect 7215 2205 7227 2257
rect 7279 2205 7335 2257
rect 7387 2205 7443 2257
rect 7495 2205 7551 2257
rect 7603 2205 7659 2257
rect 7711 2205 7723 2257
rect 7215 2149 7723 2205
rect 7215 2097 7227 2149
rect 7279 2097 7335 2149
rect 7387 2097 7443 2149
rect 7495 2097 7551 2149
rect 7603 2097 7659 2149
rect 7711 2097 7723 2149
rect 7215 2041 7723 2097
rect 7215 1989 7227 2041
rect 7279 1989 7335 2041
rect 7387 1989 7443 2041
rect 7495 1989 7551 2041
rect 7603 1989 7659 2041
rect 7711 1989 7723 2041
rect 7215 876 7723 1989
rect 7215 824 7227 876
rect 7279 824 7335 876
rect 7387 824 7443 876
rect 7495 824 7551 876
rect 7603 824 7659 876
rect 7711 824 7723 876
rect 7215 768 7723 824
rect 7215 716 7227 768
rect 7279 716 7335 768
rect 7387 716 7443 768
rect 7495 716 7551 768
rect 7603 716 7659 768
rect 7711 716 7723 768
rect 7215 43 7723 716
rect 7783 13314 8291 56440
rect 7783 13262 7825 13314
rect 7877 13262 7949 13314
rect 8001 13262 8073 13314
rect 8125 13262 8197 13314
rect 8249 13262 8291 13314
rect 7783 13190 8291 13262
rect 7783 13138 7825 13190
rect 7877 13138 7949 13190
rect 8001 13138 8073 13190
rect 8125 13138 8197 13190
rect 8249 13138 8291 13190
rect 7783 13066 8291 13138
rect 7783 13014 7825 13066
rect 7877 13014 7949 13066
rect 8001 13014 8073 13066
rect 8125 13014 8197 13066
rect 8249 13014 8291 13066
rect 7783 12942 8291 13014
rect 7783 12890 7825 12942
rect 7877 12890 7949 12942
rect 8001 12890 8073 12942
rect 8125 12890 8197 12942
rect 8249 12890 8291 12942
rect 7783 12818 8291 12890
rect 7783 12766 7825 12818
rect 7877 12766 7949 12818
rect 8001 12766 8073 12818
rect 8125 12766 8197 12818
rect 8249 12766 8291 12818
rect 7783 11910 8291 12766
rect 7783 11858 7825 11910
rect 7877 11858 7949 11910
rect 8001 11858 8073 11910
rect 8125 11858 8197 11910
rect 8249 11858 8291 11910
rect 7783 11786 8291 11858
rect 7783 11734 7825 11786
rect 7877 11734 7949 11786
rect 8001 11734 8073 11786
rect 8125 11734 8197 11786
rect 8249 11734 8291 11786
rect 7783 11662 8291 11734
rect 7783 11610 7825 11662
rect 7877 11610 7949 11662
rect 8001 11610 8073 11662
rect 8125 11610 8197 11662
rect 8249 11610 8291 11662
rect 7783 11538 8291 11610
rect 7783 11486 7825 11538
rect 7877 11486 7949 11538
rect 8001 11486 8073 11538
rect 8125 11486 8197 11538
rect 8249 11486 8291 11538
rect 7783 11414 8291 11486
rect 7783 11362 7825 11414
rect 7877 11362 7949 11414
rect 8001 11362 8073 11414
rect 8125 11362 8197 11414
rect 8249 11362 8291 11414
rect 7783 10506 8291 11362
rect 7783 10454 7825 10506
rect 7877 10454 7949 10506
rect 8001 10454 8073 10506
rect 8125 10454 8197 10506
rect 8249 10454 8291 10506
rect 7783 10382 8291 10454
rect 7783 10330 7825 10382
rect 7877 10330 7949 10382
rect 8001 10330 8073 10382
rect 8125 10330 8197 10382
rect 8249 10330 8291 10382
rect 7783 10258 8291 10330
rect 7783 10206 7825 10258
rect 7877 10206 7949 10258
rect 8001 10206 8073 10258
rect 8125 10206 8197 10258
rect 8249 10206 8291 10258
rect 7783 10134 8291 10206
rect 7783 10082 7825 10134
rect 7877 10082 7949 10134
rect 8001 10082 8073 10134
rect 8125 10082 8197 10134
rect 8249 10082 8291 10134
rect 7783 10010 8291 10082
rect 7783 9958 7825 10010
rect 7877 9958 7949 10010
rect 8001 9958 8073 10010
rect 8125 9958 8197 10010
rect 8249 9958 8291 10010
rect 7783 9102 8291 9958
rect 7783 9050 7825 9102
rect 7877 9050 7949 9102
rect 8001 9050 8073 9102
rect 8125 9050 8197 9102
rect 8249 9050 8291 9102
rect 7783 8978 8291 9050
rect 7783 8926 7825 8978
rect 7877 8926 7949 8978
rect 8001 8926 8073 8978
rect 8125 8926 8197 8978
rect 8249 8926 8291 8978
rect 7783 8854 8291 8926
rect 7783 8802 7825 8854
rect 7877 8802 7949 8854
rect 8001 8802 8073 8854
rect 8125 8802 8197 8854
rect 8249 8802 8291 8854
rect 7783 8730 8291 8802
rect 7783 8678 7825 8730
rect 7877 8678 7949 8730
rect 8001 8678 8073 8730
rect 8125 8678 8197 8730
rect 8249 8678 8291 8730
rect 7783 8606 8291 8678
rect 7783 8554 7825 8606
rect 7877 8554 7949 8606
rect 8001 8554 8073 8606
rect 8125 8554 8197 8606
rect 8249 8554 8291 8606
rect 7783 5907 8291 8554
rect 7783 5855 7825 5907
rect 7877 5855 7949 5907
rect 8001 5855 8073 5907
rect 8125 5855 8197 5907
rect 8249 5855 8291 5907
rect 7783 5783 8291 5855
rect 7783 5731 7825 5783
rect 7877 5731 7949 5783
rect 8001 5731 8073 5783
rect 8125 5731 8197 5783
rect 8249 5731 8291 5783
rect 7783 5659 8291 5731
rect 7783 5607 7825 5659
rect 7877 5607 7949 5659
rect 8001 5607 8073 5659
rect 8125 5607 8197 5659
rect 8249 5607 8291 5659
rect 7783 5535 8291 5607
rect 7783 5483 7825 5535
rect 7877 5483 7949 5535
rect 8001 5483 8073 5535
rect 8125 5483 8197 5535
rect 8249 5483 8291 5535
rect 7783 5411 8291 5483
rect 7783 5359 7825 5411
rect 7877 5359 7949 5411
rect 8001 5359 8073 5411
rect 8125 5359 8197 5411
rect 8249 5359 8291 5411
rect 7783 4503 8291 5359
rect 7783 4451 7825 4503
rect 7877 4451 7949 4503
rect 8001 4451 8073 4503
rect 8125 4451 8197 4503
rect 8249 4451 8291 4503
rect 7783 4379 8291 4451
rect 7783 4327 7825 4379
rect 7877 4327 7949 4379
rect 8001 4327 8073 4379
rect 8125 4327 8197 4379
rect 8249 4327 8291 4379
rect 7783 4255 8291 4327
rect 7783 4203 7825 4255
rect 7877 4203 7949 4255
rect 8001 4203 8073 4255
rect 8125 4203 8197 4255
rect 8249 4203 8291 4255
rect 7783 4131 8291 4203
rect 7783 4079 7825 4131
rect 7877 4079 7949 4131
rect 8001 4079 8073 4131
rect 8125 4079 8197 4131
rect 8249 4079 8291 4131
rect 7783 4007 8291 4079
rect 7783 3955 7825 4007
rect 7877 3955 7949 4007
rect 8001 3955 8073 4007
rect 8125 3955 8197 4007
rect 8249 3955 8291 4007
rect 7783 3099 8291 3955
rect 7783 3047 7825 3099
rect 7877 3047 7949 3099
rect 8001 3047 8073 3099
rect 8125 3047 8197 3099
rect 8249 3047 8291 3099
rect 7783 2975 8291 3047
rect 7783 2923 7825 2975
rect 7877 2923 7949 2975
rect 8001 2923 8073 2975
rect 8125 2923 8197 2975
rect 8249 2923 8291 2975
rect 7783 2851 8291 2923
rect 7783 2799 7825 2851
rect 7877 2799 7949 2851
rect 8001 2799 8073 2851
rect 8125 2799 8197 2851
rect 8249 2799 8291 2851
rect 7783 2727 8291 2799
rect 7783 2675 7825 2727
rect 7877 2675 7949 2727
rect 8001 2675 8073 2727
rect 8125 2675 8197 2727
rect 8249 2675 8291 2727
rect 7783 2603 8291 2675
rect 7783 2551 7825 2603
rect 7877 2551 7949 2603
rect 8001 2551 8073 2603
rect 8125 2551 8197 2603
rect 8249 2551 8291 2603
rect 7783 1695 8291 2551
rect 7783 1643 7825 1695
rect 7877 1643 7949 1695
rect 8001 1643 8073 1695
rect 8125 1643 8197 1695
rect 8249 1643 8291 1695
rect 7783 1571 8291 1643
rect 7783 1519 7825 1571
rect 7877 1519 7949 1571
rect 8001 1519 8073 1571
rect 8125 1519 8197 1571
rect 8249 1519 8291 1571
rect 7783 1447 8291 1519
rect 7783 1395 7825 1447
rect 7877 1395 7949 1447
rect 8001 1395 8073 1447
rect 8125 1395 8197 1447
rect 8249 1395 8291 1447
rect 7783 1323 8291 1395
rect 7783 1271 7825 1323
rect 7877 1271 7949 1323
rect 8001 1271 8073 1323
rect 8125 1271 8197 1323
rect 8249 1271 8291 1323
rect 7783 1199 8291 1271
rect 7783 1147 7825 1199
rect 7877 1147 7949 1199
rect 8001 1147 8073 1199
rect 8125 1147 8197 1199
rect 8249 1147 8291 1199
rect 7783 -857 8291 1147
rect 8351 13745 8859 14905
rect 8351 13693 8363 13745
rect 8415 13693 8471 13745
rect 8523 13693 8579 13745
rect 8631 13693 8687 13745
rect 8739 13693 8795 13745
rect 8847 13693 8859 13745
rect 8351 13637 8859 13693
rect 8351 13585 8363 13637
rect 8415 13585 8471 13637
rect 8523 13585 8579 13637
rect 8631 13585 8687 13637
rect 8739 13585 8795 13637
rect 8847 13585 8859 13637
rect 8351 12472 8859 13585
rect 8351 12420 8363 12472
rect 8415 12420 8471 12472
rect 8523 12420 8579 12472
rect 8631 12420 8687 12472
rect 8739 12420 8795 12472
rect 8847 12420 8859 12472
rect 8351 12364 8859 12420
rect 8351 12312 8363 12364
rect 8415 12312 8471 12364
rect 8523 12312 8579 12364
rect 8631 12312 8687 12364
rect 8739 12312 8795 12364
rect 8847 12312 8859 12364
rect 8351 12256 8859 12312
rect 8351 12204 8363 12256
rect 8415 12204 8471 12256
rect 8523 12204 8579 12256
rect 8631 12204 8687 12256
rect 8739 12204 8795 12256
rect 8847 12204 8859 12256
rect 8351 11068 8859 12204
rect 8351 11016 8363 11068
rect 8415 11016 8471 11068
rect 8523 11016 8579 11068
rect 8631 11016 8687 11068
rect 8739 11016 8795 11068
rect 8847 11016 8859 11068
rect 8351 10960 8859 11016
rect 8351 10908 8363 10960
rect 8415 10908 8471 10960
rect 8523 10908 8579 10960
rect 8631 10908 8687 10960
rect 8739 10908 8795 10960
rect 8847 10908 8859 10960
rect 8351 10852 8859 10908
rect 8351 10800 8363 10852
rect 8415 10800 8471 10852
rect 8523 10800 8579 10852
rect 8631 10800 8687 10852
rect 8739 10800 8795 10852
rect 8847 10800 8859 10852
rect 8351 9664 8859 10800
rect 8351 9612 8363 9664
rect 8415 9612 8471 9664
rect 8523 9612 8579 9664
rect 8631 9612 8687 9664
rect 8739 9612 8795 9664
rect 8847 9612 8859 9664
rect 8351 9556 8859 9612
rect 8351 9504 8363 9556
rect 8415 9504 8471 9556
rect 8523 9504 8579 9556
rect 8631 9504 8687 9556
rect 8739 9504 8795 9556
rect 8847 9504 8859 9556
rect 8351 9448 8859 9504
rect 8351 9396 8363 9448
rect 8415 9396 8471 9448
rect 8523 9396 8579 9448
rect 8631 9396 8687 9448
rect 8739 9396 8795 9448
rect 8847 9396 8859 9448
rect 8351 8283 8859 9396
rect 8351 8231 8363 8283
rect 8415 8231 8471 8283
rect 8523 8231 8579 8283
rect 8631 8231 8687 8283
rect 8739 8231 8795 8283
rect 8847 8231 8859 8283
rect 8351 8175 8859 8231
rect 8351 8123 8363 8175
rect 8415 8123 8471 8175
rect 8523 8123 8579 8175
rect 8631 8123 8687 8175
rect 8739 8123 8795 8175
rect 8847 8123 8859 8175
rect 8351 6989 8859 8123
rect 8351 6937 8393 6989
rect 8445 6937 8517 6989
rect 8569 6937 8641 6989
rect 8693 6937 8765 6989
rect 8817 6937 8859 6989
rect 8351 6865 8859 6937
rect 8351 6813 8393 6865
rect 8445 6813 8517 6865
rect 8569 6813 8641 6865
rect 8693 6813 8765 6865
rect 8817 6813 8859 6865
rect 8351 6741 8859 6813
rect 8351 6689 8393 6741
rect 8445 6689 8517 6741
rect 8569 6689 8641 6741
rect 8693 6689 8765 6741
rect 8817 6689 8859 6741
rect 8351 6617 8859 6689
rect 8351 6565 8393 6617
rect 8445 6565 8517 6617
rect 8569 6565 8641 6617
rect 8693 6565 8765 6617
rect 8817 6565 8859 6617
rect 8351 489 8859 6565
rect 8351 437 8393 489
rect 8445 437 8517 489
rect 8569 437 8641 489
rect 8693 437 8765 489
rect 8817 437 8859 489
rect 8351 365 8859 437
rect 8351 313 8393 365
rect 8445 313 8517 365
rect 8569 313 8641 365
rect 8693 313 8765 365
rect 8817 313 8859 365
rect 8351 241 8859 313
rect 8351 189 8393 241
rect 8445 189 8517 241
rect 8569 189 8641 241
rect 8693 189 8765 241
rect 8817 189 8859 241
rect 8351 117 8859 189
rect 8351 65 8393 117
rect 8445 65 8517 117
rect 8569 65 8641 117
rect 8693 65 8765 117
rect 8817 65 8859 117
rect 8351 43 8859 65
rect 8919 13314 9427 56440
rect 8919 13262 8961 13314
rect 9013 13262 9085 13314
rect 9137 13262 9209 13314
rect 9261 13262 9333 13314
rect 9385 13262 9427 13314
rect 8919 13190 9427 13262
rect 8919 13138 8961 13190
rect 9013 13138 9085 13190
rect 9137 13138 9209 13190
rect 9261 13138 9333 13190
rect 9385 13138 9427 13190
rect 8919 13066 9427 13138
rect 8919 13014 8961 13066
rect 9013 13014 9085 13066
rect 9137 13014 9209 13066
rect 9261 13014 9333 13066
rect 9385 13014 9427 13066
rect 8919 12942 9427 13014
rect 8919 12890 8961 12942
rect 9013 12890 9085 12942
rect 9137 12890 9209 12942
rect 9261 12890 9333 12942
rect 9385 12890 9427 12942
rect 8919 12818 9427 12890
rect 8919 12766 8961 12818
rect 9013 12766 9085 12818
rect 9137 12766 9209 12818
rect 9261 12766 9333 12818
rect 9385 12766 9427 12818
rect 8919 11910 9427 12766
rect 8919 11858 8961 11910
rect 9013 11858 9085 11910
rect 9137 11858 9209 11910
rect 9261 11858 9333 11910
rect 9385 11858 9427 11910
rect 8919 11786 9427 11858
rect 8919 11734 8961 11786
rect 9013 11734 9085 11786
rect 9137 11734 9209 11786
rect 9261 11734 9333 11786
rect 9385 11734 9427 11786
rect 8919 11662 9427 11734
rect 8919 11610 8961 11662
rect 9013 11610 9085 11662
rect 9137 11610 9209 11662
rect 9261 11610 9333 11662
rect 9385 11610 9427 11662
rect 8919 11538 9427 11610
rect 8919 11486 8961 11538
rect 9013 11486 9085 11538
rect 9137 11486 9209 11538
rect 9261 11486 9333 11538
rect 9385 11486 9427 11538
rect 8919 11414 9427 11486
rect 8919 11362 8961 11414
rect 9013 11362 9085 11414
rect 9137 11362 9209 11414
rect 9261 11362 9333 11414
rect 9385 11362 9427 11414
rect 8919 10506 9427 11362
rect 8919 10454 8961 10506
rect 9013 10454 9085 10506
rect 9137 10454 9209 10506
rect 9261 10454 9333 10506
rect 9385 10454 9427 10506
rect 8919 10382 9427 10454
rect 8919 10330 8961 10382
rect 9013 10330 9085 10382
rect 9137 10330 9209 10382
rect 9261 10330 9333 10382
rect 9385 10330 9427 10382
rect 8919 10258 9427 10330
rect 8919 10206 8961 10258
rect 9013 10206 9085 10258
rect 9137 10206 9209 10258
rect 9261 10206 9333 10258
rect 9385 10206 9427 10258
rect 8919 10134 9427 10206
rect 8919 10082 8961 10134
rect 9013 10082 9085 10134
rect 9137 10082 9209 10134
rect 9261 10082 9333 10134
rect 9385 10082 9427 10134
rect 8919 10010 9427 10082
rect 8919 9958 8961 10010
rect 9013 9958 9085 10010
rect 9137 9958 9209 10010
rect 9261 9958 9333 10010
rect 9385 9958 9427 10010
rect 8919 9102 9427 9958
rect 8919 9050 8961 9102
rect 9013 9050 9085 9102
rect 9137 9050 9209 9102
rect 9261 9050 9333 9102
rect 9385 9050 9427 9102
rect 8919 8978 9427 9050
rect 8919 8926 8961 8978
rect 9013 8926 9085 8978
rect 9137 8926 9209 8978
rect 9261 8926 9333 8978
rect 9385 8926 9427 8978
rect 8919 8854 9427 8926
rect 8919 8802 8961 8854
rect 9013 8802 9085 8854
rect 9137 8802 9209 8854
rect 9261 8802 9333 8854
rect 9385 8802 9427 8854
rect 8919 8730 9427 8802
rect 8919 8678 8961 8730
rect 9013 8678 9085 8730
rect 9137 8678 9209 8730
rect 9261 8678 9333 8730
rect 9385 8678 9427 8730
rect 8919 8606 9427 8678
rect 8919 8554 8961 8606
rect 9013 8554 9085 8606
rect 9137 8554 9209 8606
rect 9261 8554 9333 8606
rect 9385 8554 9427 8606
rect 8919 5907 9427 8554
rect 8919 5855 8961 5907
rect 9013 5855 9085 5907
rect 9137 5855 9209 5907
rect 9261 5855 9333 5907
rect 9385 5855 9427 5907
rect 8919 5783 9427 5855
rect 8919 5731 8961 5783
rect 9013 5731 9085 5783
rect 9137 5731 9209 5783
rect 9261 5731 9333 5783
rect 9385 5731 9427 5783
rect 8919 5659 9427 5731
rect 8919 5607 8961 5659
rect 9013 5607 9085 5659
rect 9137 5607 9209 5659
rect 9261 5607 9333 5659
rect 9385 5607 9427 5659
rect 8919 5535 9427 5607
rect 8919 5483 8961 5535
rect 9013 5483 9085 5535
rect 9137 5483 9209 5535
rect 9261 5483 9333 5535
rect 9385 5483 9427 5535
rect 8919 5411 9427 5483
rect 8919 5359 8961 5411
rect 9013 5359 9085 5411
rect 9137 5359 9209 5411
rect 9261 5359 9333 5411
rect 9385 5359 9427 5411
rect 8919 4503 9427 5359
rect 8919 4451 8961 4503
rect 9013 4451 9085 4503
rect 9137 4451 9209 4503
rect 9261 4451 9333 4503
rect 9385 4451 9427 4503
rect 8919 4379 9427 4451
rect 8919 4327 8961 4379
rect 9013 4327 9085 4379
rect 9137 4327 9209 4379
rect 9261 4327 9333 4379
rect 9385 4327 9427 4379
rect 8919 4255 9427 4327
rect 8919 4203 8961 4255
rect 9013 4203 9085 4255
rect 9137 4203 9209 4255
rect 9261 4203 9333 4255
rect 9385 4203 9427 4255
rect 8919 4131 9427 4203
rect 8919 4079 8961 4131
rect 9013 4079 9085 4131
rect 9137 4079 9209 4131
rect 9261 4079 9333 4131
rect 9385 4079 9427 4131
rect 8919 4007 9427 4079
rect 8919 3955 8961 4007
rect 9013 3955 9085 4007
rect 9137 3955 9209 4007
rect 9261 3955 9333 4007
rect 9385 3955 9427 4007
rect 8919 3099 9427 3955
rect 8919 3047 8961 3099
rect 9013 3047 9085 3099
rect 9137 3047 9209 3099
rect 9261 3047 9333 3099
rect 9385 3047 9427 3099
rect 8919 2975 9427 3047
rect 8919 2923 8961 2975
rect 9013 2923 9085 2975
rect 9137 2923 9209 2975
rect 9261 2923 9333 2975
rect 9385 2923 9427 2975
rect 8919 2851 9427 2923
rect 8919 2799 8961 2851
rect 9013 2799 9085 2851
rect 9137 2799 9209 2851
rect 9261 2799 9333 2851
rect 9385 2799 9427 2851
rect 8919 2727 9427 2799
rect 8919 2675 8961 2727
rect 9013 2675 9085 2727
rect 9137 2675 9209 2727
rect 9261 2675 9333 2727
rect 9385 2675 9427 2727
rect 8919 2603 9427 2675
rect 8919 2551 8961 2603
rect 9013 2551 9085 2603
rect 9137 2551 9209 2603
rect 9261 2551 9333 2603
rect 9385 2551 9427 2603
rect 8919 1695 9427 2551
rect 8919 1643 8961 1695
rect 9013 1643 9085 1695
rect 9137 1643 9209 1695
rect 9261 1643 9333 1695
rect 9385 1643 9427 1695
rect 8919 1571 9427 1643
rect 8919 1519 8961 1571
rect 9013 1519 9085 1571
rect 9137 1519 9209 1571
rect 9261 1519 9333 1571
rect 9385 1519 9427 1571
rect 8919 1447 9427 1519
rect 8919 1395 8961 1447
rect 9013 1395 9085 1447
rect 9137 1395 9209 1447
rect 9261 1395 9333 1447
rect 9385 1395 9427 1447
rect 8919 1323 9427 1395
rect 8919 1271 8961 1323
rect 9013 1271 9085 1323
rect 9137 1271 9209 1323
rect 9261 1271 9333 1323
rect 9385 1271 9427 1323
rect 8919 1199 9427 1271
rect 8919 1147 8961 1199
rect 9013 1147 9085 1199
rect 9137 1147 9209 1199
rect 9261 1147 9333 1199
rect 9385 1147 9427 1199
rect 8919 -857 9427 1147
rect 9487 14396 9995 14905
rect 9487 14344 9529 14396
rect 9581 14344 9653 14396
rect 9705 14344 9777 14396
rect 9829 14344 9901 14396
rect 9953 14344 9995 14396
rect 9487 14272 9995 14344
rect 9487 14220 9529 14272
rect 9581 14220 9653 14272
rect 9705 14220 9777 14272
rect 9829 14220 9901 14272
rect 9953 14220 9995 14272
rect 9487 14148 9995 14220
rect 9487 14096 9529 14148
rect 9581 14096 9653 14148
rect 9705 14096 9777 14148
rect 9829 14096 9901 14148
rect 9953 14096 9995 14148
rect 9487 14024 9995 14096
rect 9487 13972 9529 14024
rect 9581 13972 9653 14024
rect 9705 13972 9777 14024
rect 9829 13972 9901 14024
rect 9953 13972 9995 14024
rect 9487 7896 9995 13972
rect 9487 7844 9529 7896
rect 9581 7844 9653 7896
rect 9705 7844 9777 7896
rect 9829 7844 9901 7896
rect 9953 7844 9995 7896
rect 9487 7772 9995 7844
rect 9487 7720 9529 7772
rect 9581 7720 9653 7772
rect 9705 7720 9777 7772
rect 9829 7720 9901 7772
rect 9953 7720 9995 7772
rect 9487 7648 9995 7720
rect 9487 7596 9529 7648
rect 9581 7596 9653 7648
rect 9705 7596 9777 7648
rect 9829 7596 9901 7648
rect 9953 7596 9995 7648
rect 9487 7524 9995 7596
rect 9487 7472 9529 7524
rect 9581 7472 9653 7524
rect 9705 7472 9777 7524
rect 9829 7472 9901 7524
rect 9953 7472 9995 7524
rect 9487 6338 9995 7472
rect 9487 6286 9499 6338
rect 9551 6286 9607 6338
rect 9659 6286 9715 6338
rect 9767 6286 9823 6338
rect 9875 6286 9931 6338
rect 9983 6286 9995 6338
rect 9487 6230 9995 6286
rect 9487 6178 9499 6230
rect 9551 6178 9607 6230
rect 9659 6178 9715 6230
rect 9767 6178 9823 6230
rect 9875 6178 9931 6230
rect 9983 6178 9995 6230
rect 9487 5065 9995 6178
rect 9487 5013 9499 5065
rect 9551 5013 9607 5065
rect 9659 5013 9715 5065
rect 9767 5013 9823 5065
rect 9875 5013 9931 5065
rect 9983 5013 9995 5065
rect 9487 4957 9995 5013
rect 9487 4905 9499 4957
rect 9551 4905 9607 4957
rect 9659 4905 9715 4957
rect 9767 4905 9823 4957
rect 9875 4905 9931 4957
rect 9983 4905 9995 4957
rect 9487 4849 9995 4905
rect 9487 4797 9499 4849
rect 9551 4797 9607 4849
rect 9659 4797 9715 4849
rect 9767 4797 9823 4849
rect 9875 4797 9931 4849
rect 9983 4797 9995 4849
rect 9487 3661 9995 4797
rect 9487 3609 9499 3661
rect 9551 3609 9607 3661
rect 9659 3609 9715 3661
rect 9767 3609 9823 3661
rect 9875 3609 9931 3661
rect 9983 3609 9995 3661
rect 9487 3553 9995 3609
rect 9487 3501 9499 3553
rect 9551 3501 9607 3553
rect 9659 3501 9715 3553
rect 9767 3501 9823 3553
rect 9875 3501 9931 3553
rect 9983 3501 9995 3553
rect 9487 3445 9995 3501
rect 9487 3393 9499 3445
rect 9551 3393 9607 3445
rect 9659 3393 9715 3445
rect 9767 3393 9823 3445
rect 9875 3393 9931 3445
rect 9983 3393 9995 3445
rect 9487 2257 9995 3393
rect 9487 2205 9499 2257
rect 9551 2205 9607 2257
rect 9659 2205 9715 2257
rect 9767 2205 9823 2257
rect 9875 2205 9931 2257
rect 9983 2205 9995 2257
rect 9487 2149 9995 2205
rect 9487 2097 9499 2149
rect 9551 2097 9607 2149
rect 9659 2097 9715 2149
rect 9767 2097 9823 2149
rect 9875 2097 9931 2149
rect 9983 2097 9995 2149
rect 9487 2041 9995 2097
rect 9487 1989 9499 2041
rect 9551 1989 9607 2041
rect 9659 1989 9715 2041
rect 9767 1989 9823 2041
rect 9875 1989 9931 2041
rect 9983 1989 9995 2041
rect 9487 876 9995 1989
rect 9487 824 9499 876
rect 9551 824 9607 876
rect 9659 824 9715 876
rect 9767 824 9823 876
rect 9875 824 9931 876
rect 9983 824 9995 876
rect 9487 768 9995 824
rect 9487 716 9499 768
rect 9551 716 9607 768
rect 9659 716 9715 768
rect 9767 716 9823 768
rect 9875 716 9931 768
rect 9983 716 9995 768
rect 9487 43 9995 716
rect 10055 13314 10563 56440
rect 10055 13262 10097 13314
rect 10149 13262 10221 13314
rect 10273 13262 10345 13314
rect 10397 13262 10469 13314
rect 10521 13262 10563 13314
rect 10055 13190 10563 13262
rect 10055 13138 10097 13190
rect 10149 13138 10221 13190
rect 10273 13138 10345 13190
rect 10397 13138 10469 13190
rect 10521 13138 10563 13190
rect 10055 13066 10563 13138
rect 10055 13014 10097 13066
rect 10149 13014 10221 13066
rect 10273 13014 10345 13066
rect 10397 13014 10469 13066
rect 10521 13014 10563 13066
rect 10055 12942 10563 13014
rect 10055 12890 10097 12942
rect 10149 12890 10221 12942
rect 10273 12890 10345 12942
rect 10397 12890 10469 12942
rect 10521 12890 10563 12942
rect 10055 12818 10563 12890
rect 10055 12766 10097 12818
rect 10149 12766 10221 12818
rect 10273 12766 10345 12818
rect 10397 12766 10469 12818
rect 10521 12766 10563 12818
rect 10055 11910 10563 12766
rect 10055 11858 10097 11910
rect 10149 11858 10221 11910
rect 10273 11858 10345 11910
rect 10397 11858 10469 11910
rect 10521 11858 10563 11910
rect 10055 11786 10563 11858
rect 10055 11734 10097 11786
rect 10149 11734 10221 11786
rect 10273 11734 10345 11786
rect 10397 11734 10469 11786
rect 10521 11734 10563 11786
rect 10055 11662 10563 11734
rect 10055 11610 10097 11662
rect 10149 11610 10221 11662
rect 10273 11610 10345 11662
rect 10397 11610 10469 11662
rect 10521 11610 10563 11662
rect 10055 11538 10563 11610
rect 10055 11486 10097 11538
rect 10149 11486 10221 11538
rect 10273 11486 10345 11538
rect 10397 11486 10469 11538
rect 10521 11486 10563 11538
rect 10055 11414 10563 11486
rect 10055 11362 10097 11414
rect 10149 11362 10221 11414
rect 10273 11362 10345 11414
rect 10397 11362 10469 11414
rect 10521 11362 10563 11414
rect 10055 10506 10563 11362
rect 10055 10454 10097 10506
rect 10149 10454 10221 10506
rect 10273 10454 10345 10506
rect 10397 10454 10469 10506
rect 10521 10454 10563 10506
rect 10055 10382 10563 10454
rect 10055 10330 10097 10382
rect 10149 10330 10221 10382
rect 10273 10330 10345 10382
rect 10397 10330 10469 10382
rect 10521 10330 10563 10382
rect 10055 10258 10563 10330
rect 10055 10206 10097 10258
rect 10149 10206 10221 10258
rect 10273 10206 10345 10258
rect 10397 10206 10469 10258
rect 10521 10206 10563 10258
rect 10055 10134 10563 10206
rect 10055 10082 10097 10134
rect 10149 10082 10221 10134
rect 10273 10082 10345 10134
rect 10397 10082 10469 10134
rect 10521 10082 10563 10134
rect 10055 10010 10563 10082
rect 10055 9958 10097 10010
rect 10149 9958 10221 10010
rect 10273 9958 10345 10010
rect 10397 9958 10469 10010
rect 10521 9958 10563 10010
rect 10055 9102 10563 9958
rect 10055 9050 10097 9102
rect 10149 9050 10221 9102
rect 10273 9050 10345 9102
rect 10397 9050 10469 9102
rect 10521 9050 10563 9102
rect 10055 8978 10563 9050
rect 10055 8926 10097 8978
rect 10149 8926 10221 8978
rect 10273 8926 10345 8978
rect 10397 8926 10469 8978
rect 10521 8926 10563 8978
rect 10055 8854 10563 8926
rect 10055 8802 10097 8854
rect 10149 8802 10221 8854
rect 10273 8802 10345 8854
rect 10397 8802 10469 8854
rect 10521 8802 10563 8854
rect 10055 8730 10563 8802
rect 10055 8678 10097 8730
rect 10149 8678 10221 8730
rect 10273 8678 10345 8730
rect 10397 8678 10469 8730
rect 10521 8678 10563 8730
rect 10055 8606 10563 8678
rect 10055 8554 10097 8606
rect 10149 8554 10221 8606
rect 10273 8554 10345 8606
rect 10397 8554 10469 8606
rect 10521 8554 10563 8606
rect 10055 5907 10563 8554
rect 10055 5855 10097 5907
rect 10149 5855 10221 5907
rect 10273 5855 10345 5907
rect 10397 5855 10469 5907
rect 10521 5855 10563 5907
rect 10055 5783 10563 5855
rect 10055 5731 10097 5783
rect 10149 5731 10221 5783
rect 10273 5731 10345 5783
rect 10397 5731 10469 5783
rect 10521 5731 10563 5783
rect 10055 5659 10563 5731
rect 10055 5607 10097 5659
rect 10149 5607 10221 5659
rect 10273 5607 10345 5659
rect 10397 5607 10469 5659
rect 10521 5607 10563 5659
rect 10055 5535 10563 5607
rect 10055 5483 10097 5535
rect 10149 5483 10221 5535
rect 10273 5483 10345 5535
rect 10397 5483 10469 5535
rect 10521 5483 10563 5535
rect 10055 5411 10563 5483
rect 10055 5359 10097 5411
rect 10149 5359 10221 5411
rect 10273 5359 10345 5411
rect 10397 5359 10469 5411
rect 10521 5359 10563 5411
rect 10055 4503 10563 5359
rect 10055 4451 10097 4503
rect 10149 4451 10221 4503
rect 10273 4451 10345 4503
rect 10397 4451 10469 4503
rect 10521 4451 10563 4503
rect 10055 4379 10563 4451
rect 10055 4327 10097 4379
rect 10149 4327 10221 4379
rect 10273 4327 10345 4379
rect 10397 4327 10469 4379
rect 10521 4327 10563 4379
rect 10055 4255 10563 4327
rect 10055 4203 10097 4255
rect 10149 4203 10221 4255
rect 10273 4203 10345 4255
rect 10397 4203 10469 4255
rect 10521 4203 10563 4255
rect 10055 4131 10563 4203
rect 10055 4079 10097 4131
rect 10149 4079 10221 4131
rect 10273 4079 10345 4131
rect 10397 4079 10469 4131
rect 10521 4079 10563 4131
rect 10055 4007 10563 4079
rect 10055 3955 10097 4007
rect 10149 3955 10221 4007
rect 10273 3955 10345 4007
rect 10397 3955 10469 4007
rect 10521 3955 10563 4007
rect 10055 3099 10563 3955
rect 10055 3047 10097 3099
rect 10149 3047 10221 3099
rect 10273 3047 10345 3099
rect 10397 3047 10469 3099
rect 10521 3047 10563 3099
rect 10055 2975 10563 3047
rect 10055 2923 10097 2975
rect 10149 2923 10221 2975
rect 10273 2923 10345 2975
rect 10397 2923 10469 2975
rect 10521 2923 10563 2975
rect 10055 2851 10563 2923
rect 10055 2799 10097 2851
rect 10149 2799 10221 2851
rect 10273 2799 10345 2851
rect 10397 2799 10469 2851
rect 10521 2799 10563 2851
rect 10055 2727 10563 2799
rect 10055 2675 10097 2727
rect 10149 2675 10221 2727
rect 10273 2675 10345 2727
rect 10397 2675 10469 2727
rect 10521 2675 10563 2727
rect 10055 2603 10563 2675
rect 10055 2551 10097 2603
rect 10149 2551 10221 2603
rect 10273 2551 10345 2603
rect 10397 2551 10469 2603
rect 10521 2551 10563 2603
rect 10055 1695 10563 2551
rect 10055 1643 10097 1695
rect 10149 1643 10221 1695
rect 10273 1643 10345 1695
rect 10397 1643 10469 1695
rect 10521 1643 10563 1695
rect 10055 1571 10563 1643
rect 10055 1519 10097 1571
rect 10149 1519 10221 1571
rect 10273 1519 10345 1571
rect 10397 1519 10469 1571
rect 10521 1519 10563 1571
rect 10055 1447 10563 1519
rect 10055 1395 10097 1447
rect 10149 1395 10221 1447
rect 10273 1395 10345 1447
rect 10397 1395 10469 1447
rect 10521 1395 10563 1447
rect 10055 1323 10563 1395
rect 10055 1271 10097 1323
rect 10149 1271 10221 1323
rect 10273 1271 10345 1323
rect 10397 1271 10469 1323
rect 10521 1271 10563 1323
rect 10055 1199 10563 1271
rect 10055 1147 10097 1199
rect 10149 1147 10221 1199
rect 10273 1147 10345 1199
rect 10397 1147 10469 1199
rect 10521 1147 10563 1199
rect 10055 -857 10563 1147
rect 10623 13745 11131 14905
rect 10623 13693 10635 13745
rect 10687 13693 10743 13745
rect 10795 13693 10851 13745
rect 10903 13693 10959 13745
rect 11011 13693 11067 13745
rect 11119 13693 11131 13745
rect 10623 13637 11131 13693
rect 10623 13585 10635 13637
rect 10687 13585 10743 13637
rect 10795 13585 10851 13637
rect 10903 13585 10959 13637
rect 11011 13585 11067 13637
rect 11119 13585 11131 13637
rect 10623 12472 11131 13585
rect 10623 12420 10635 12472
rect 10687 12420 10743 12472
rect 10795 12420 10851 12472
rect 10903 12420 10959 12472
rect 11011 12420 11067 12472
rect 11119 12420 11131 12472
rect 10623 12364 11131 12420
rect 10623 12312 10635 12364
rect 10687 12312 10743 12364
rect 10795 12312 10851 12364
rect 10903 12312 10959 12364
rect 11011 12312 11067 12364
rect 11119 12312 11131 12364
rect 10623 12256 11131 12312
rect 10623 12204 10635 12256
rect 10687 12204 10743 12256
rect 10795 12204 10851 12256
rect 10903 12204 10959 12256
rect 11011 12204 11067 12256
rect 11119 12204 11131 12256
rect 10623 11068 11131 12204
rect 10623 11016 10635 11068
rect 10687 11016 10743 11068
rect 10795 11016 10851 11068
rect 10903 11016 10959 11068
rect 11011 11016 11067 11068
rect 11119 11016 11131 11068
rect 10623 10960 11131 11016
rect 10623 10908 10635 10960
rect 10687 10908 10743 10960
rect 10795 10908 10851 10960
rect 10903 10908 10959 10960
rect 11011 10908 11067 10960
rect 11119 10908 11131 10960
rect 10623 10852 11131 10908
rect 10623 10800 10635 10852
rect 10687 10800 10743 10852
rect 10795 10800 10851 10852
rect 10903 10800 10959 10852
rect 11011 10800 11067 10852
rect 11119 10800 11131 10852
rect 10623 9664 11131 10800
rect 10623 9612 10635 9664
rect 10687 9612 10743 9664
rect 10795 9612 10851 9664
rect 10903 9612 10959 9664
rect 11011 9612 11067 9664
rect 11119 9612 11131 9664
rect 10623 9556 11131 9612
rect 10623 9504 10635 9556
rect 10687 9504 10743 9556
rect 10795 9504 10851 9556
rect 10903 9504 10959 9556
rect 11011 9504 11067 9556
rect 11119 9504 11131 9556
rect 10623 9448 11131 9504
rect 10623 9396 10635 9448
rect 10687 9396 10743 9448
rect 10795 9396 10851 9448
rect 10903 9396 10959 9448
rect 11011 9396 11067 9448
rect 11119 9396 11131 9448
rect 10623 8283 11131 9396
rect 10623 8231 10635 8283
rect 10687 8231 10743 8283
rect 10795 8231 10851 8283
rect 10903 8231 10959 8283
rect 11011 8231 11067 8283
rect 11119 8231 11131 8283
rect 10623 8175 11131 8231
rect 10623 8123 10635 8175
rect 10687 8123 10743 8175
rect 10795 8123 10851 8175
rect 10903 8123 10959 8175
rect 11011 8123 11067 8175
rect 11119 8123 11131 8175
rect 10623 6989 11131 8123
rect 10623 6937 10665 6989
rect 10717 6937 10789 6989
rect 10841 6937 10913 6989
rect 10965 6937 11037 6989
rect 11089 6937 11131 6989
rect 10623 6865 11131 6937
rect 10623 6813 10665 6865
rect 10717 6813 10789 6865
rect 10841 6813 10913 6865
rect 10965 6813 11037 6865
rect 11089 6813 11131 6865
rect 10623 6741 11131 6813
rect 10623 6689 10665 6741
rect 10717 6689 10789 6741
rect 10841 6689 10913 6741
rect 10965 6689 11037 6741
rect 11089 6689 11131 6741
rect 10623 6617 11131 6689
rect 10623 6565 10665 6617
rect 10717 6565 10789 6617
rect 10841 6565 10913 6617
rect 10965 6565 11037 6617
rect 11089 6565 11131 6617
rect 10623 489 11131 6565
rect 10623 437 10665 489
rect 10717 437 10789 489
rect 10841 437 10913 489
rect 10965 437 11037 489
rect 11089 437 11131 489
rect 10623 365 11131 437
rect 10623 313 10665 365
rect 10717 313 10789 365
rect 10841 313 10913 365
rect 10965 313 11037 365
rect 11089 313 11131 365
rect 10623 241 11131 313
rect 10623 189 10665 241
rect 10717 189 10789 241
rect 10841 189 10913 241
rect 10965 189 11037 241
rect 11089 189 11131 241
rect 10623 117 11131 189
rect 10623 65 10665 117
rect 10717 65 10789 117
rect 10841 65 10913 117
rect 10965 65 11037 117
rect 11089 65 11131 117
rect 10623 43 11131 65
rect 11191 14396 11699 14905
rect 11191 14344 11233 14396
rect 11285 14344 11357 14396
rect 11409 14344 11481 14396
rect 11533 14344 11605 14396
rect 11657 14344 11699 14396
rect 11191 14272 11699 14344
rect 11191 14220 11233 14272
rect 11285 14220 11357 14272
rect 11409 14220 11481 14272
rect 11533 14220 11605 14272
rect 11657 14220 11699 14272
rect 11191 14148 11699 14220
rect 11191 14096 11233 14148
rect 11285 14096 11357 14148
rect 11409 14096 11481 14148
rect 11533 14096 11605 14148
rect 11657 14096 11699 14148
rect 11191 14024 11699 14096
rect 11191 13972 11233 14024
rect 11285 13972 11357 14024
rect 11409 13972 11481 14024
rect 11533 13972 11605 14024
rect 11657 13972 11699 14024
rect 11191 7896 11699 13972
rect 11191 7844 11233 7896
rect 11285 7844 11357 7896
rect 11409 7844 11481 7896
rect 11533 7844 11605 7896
rect 11657 7844 11699 7896
rect 11191 7772 11699 7844
rect 11191 7720 11233 7772
rect 11285 7720 11357 7772
rect 11409 7720 11481 7772
rect 11533 7720 11605 7772
rect 11657 7720 11699 7772
rect 11191 7648 11699 7720
rect 11191 7596 11233 7648
rect 11285 7596 11357 7648
rect 11409 7596 11481 7648
rect 11533 7596 11605 7648
rect 11657 7596 11699 7648
rect 11191 7524 11699 7596
rect 11191 7472 11233 7524
rect 11285 7472 11357 7524
rect 11409 7472 11481 7524
rect 11533 7472 11605 7524
rect 11657 7472 11699 7524
rect 11191 6307 11699 7472
rect 11191 6255 11365 6307
rect 11417 6255 11473 6307
rect 11525 6255 11699 6307
rect 11191 6199 11699 6255
rect 11191 6147 11365 6199
rect 11417 6147 11473 6199
rect 11525 6147 11699 6199
rect 11191 6091 11699 6147
rect 11191 6039 11365 6091
rect 11417 6039 11473 6091
rect 11525 6039 11699 6091
rect 11191 5983 11699 6039
rect 11191 5931 11365 5983
rect 11417 5931 11473 5983
rect 11525 5931 11699 5983
rect 11191 5875 11699 5931
rect 11191 5823 11365 5875
rect 11417 5823 11473 5875
rect 11525 5823 11699 5875
rect 11191 5767 11699 5823
rect 11191 5715 11365 5767
rect 11417 5715 11473 5767
rect 11525 5715 11699 5767
rect 11191 5659 11699 5715
rect 11191 5607 11365 5659
rect 11417 5607 11473 5659
rect 11525 5607 11699 5659
rect 11191 5551 11699 5607
rect 11191 5499 11365 5551
rect 11417 5499 11473 5551
rect 11525 5499 11699 5551
rect 11191 5443 11699 5499
rect 11191 5391 11365 5443
rect 11417 5391 11473 5443
rect 11525 5391 11699 5443
rect 11191 5335 11699 5391
rect 11191 5283 11365 5335
rect 11417 5283 11473 5335
rect 11525 5283 11699 5335
rect 11191 5227 11699 5283
rect 11191 5175 11365 5227
rect 11417 5175 11473 5227
rect 11525 5175 11699 5227
rect 11191 5119 11699 5175
rect 11191 5067 11365 5119
rect 11417 5067 11473 5119
rect 11525 5067 11699 5119
rect 11191 5011 11699 5067
rect 11191 4959 11365 5011
rect 11417 4959 11473 5011
rect 11525 4959 11699 5011
rect 11191 4903 11699 4959
rect 11191 4851 11365 4903
rect 11417 4851 11473 4903
rect 11525 4851 11699 4903
rect 11191 4795 11699 4851
rect 11191 4743 11365 4795
rect 11417 4743 11473 4795
rect 11525 4743 11699 4795
rect 11191 4687 11699 4743
rect 11191 4635 11365 4687
rect 11417 4635 11473 4687
rect 11525 4635 11699 4687
rect 11191 4579 11699 4635
rect 11191 4527 11365 4579
rect 11417 4527 11473 4579
rect 11525 4527 11699 4579
rect 11191 4471 11699 4527
rect 11191 4419 11365 4471
rect 11417 4419 11473 4471
rect 11525 4419 11699 4471
rect 11191 4363 11699 4419
rect 11191 4311 11365 4363
rect 11417 4311 11473 4363
rect 11525 4311 11699 4363
rect 11191 4255 11699 4311
rect 11191 4203 11365 4255
rect 11417 4203 11473 4255
rect 11525 4203 11699 4255
rect 11191 4147 11699 4203
rect 11191 4095 11365 4147
rect 11417 4095 11473 4147
rect 11525 4095 11699 4147
rect 11191 4039 11699 4095
rect 11191 3987 11365 4039
rect 11417 3987 11473 4039
rect 11525 3987 11699 4039
rect 11191 3931 11699 3987
rect 11191 3879 11365 3931
rect 11417 3879 11473 3931
rect 11525 3879 11699 3931
rect 11191 3823 11699 3879
rect 11191 3771 11365 3823
rect 11417 3771 11473 3823
rect 11525 3771 11699 3823
rect 11191 3715 11699 3771
rect 11191 3663 11365 3715
rect 11417 3663 11473 3715
rect 11525 3663 11699 3715
rect 11191 3607 11699 3663
rect 11191 3555 11365 3607
rect 11417 3555 11473 3607
rect 11525 3555 11699 3607
rect 11191 3499 11699 3555
rect 11191 3447 11365 3499
rect 11417 3447 11473 3499
rect 11525 3447 11699 3499
rect 11191 3391 11699 3447
rect 11191 3339 11365 3391
rect 11417 3339 11473 3391
rect 11525 3339 11699 3391
rect 11191 3283 11699 3339
rect 11191 3231 11365 3283
rect 11417 3231 11473 3283
rect 11525 3231 11699 3283
rect 11191 3175 11699 3231
rect 11191 3123 11365 3175
rect 11417 3123 11473 3175
rect 11525 3123 11699 3175
rect 11191 3067 11699 3123
rect 11191 3015 11365 3067
rect 11417 3015 11473 3067
rect 11525 3015 11699 3067
rect 11191 2959 11699 3015
rect 11191 2907 11365 2959
rect 11417 2907 11473 2959
rect 11525 2907 11699 2959
rect 11191 2851 11699 2907
rect 11191 2799 11365 2851
rect 11417 2799 11473 2851
rect 11525 2799 11699 2851
rect 11191 2743 11699 2799
rect 11191 2691 11365 2743
rect 11417 2691 11473 2743
rect 11525 2691 11699 2743
rect 11191 2635 11699 2691
rect 11191 2583 11365 2635
rect 11417 2583 11473 2635
rect 11525 2583 11699 2635
rect 11191 2527 11699 2583
rect 11191 2475 11365 2527
rect 11417 2475 11473 2527
rect 11525 2475 11699 2527
rect 11191 2419 11699 2475
rect 11191 2367 11365 2419
rect 11417 2367 11473 2419
rect 11525 2367 11699 2419
rect 11191 2311 11699 2367
rect 11191 2259 11365 2311
rect 11417 2259 11473 2311
rect 11525 2259 11699 2311
rect 11191 2203 11699 2259
rect 11191 2151 11365 2203
rect 11417 2151 11473 2203
rect 11525 2151 11699 2203
rect 11191 2095 11699 2151
rect 11191 2043 11365 2095
rect 11417 2043 11473 2095
rect 11525 2043 11699 2095
rect 11191 1987 11699 2043
rect 11191 1935 11365 1987
rect 11417 1935 11473 1987
rect 11525 1935 11699 1987
rect 11191 1879 11699 1935
rect 11191 1827 11365 1879
rect 11417 1827 11473 1879
rect 11525 1827 11699 1879
rect 11191 1771 11699 1827
rect 11191 1719 11365 1771
rect 11417 1719 11473 1771
rect 11525 1719 11699 1771
rect 11191 1663 11699 1719
rect 11191 1611 11365 1663
rect 11417 1611 11473 1663
rect 11525 1611 11699 1663
rect 11191 1555 11699 1611
rect 11191 1503 11365 1555
rect 11417 1503 11473 1555
rect 11525 1503 11699 1555
rect 11191 1447 11699 1503
rect 11191 1395 11365 1447
rect 11417 1395 11473 1447
rect 11525 1395 11699 1447
rect 11191 1339 11699 1395
rect 11191 1287 11365 1339
rect 11417 1287 11473 1339
rect 11525 1287 11699 1339
rect 11191 1231 11699 1287
rect 11191 1179 11365 1231
rect 11417 1179 11473 1231
rect 11525 1179 11699 1231
rect 11191 1123 11699 1179
rect 11191 1071 11365 1123
rect 11417 1071 11473 1123
rect 11525 1071 11699 1123
rect 11191 1015 11699 1071
rect 11191 963 11365 1015
rect 11417 963 11473 1015
rect 11525 963 11699 1015
rect 11191 907 11699 963
rect 11191 855 11365 907
rect 11417 855 11473 907
rect 11525 855 11699 907
rect 11191 799 11699 855
rect 11191 747 11365 799
rect 11417 747 11473 799
rect 11525 747 11699 799
rect 11191 43 11699 747
rect 11759 6955 12267 14905
rect 11759 6903 11805 6955
rect 11857 6903 11913 6955
rect 11965 6903 12021 6955
rect 12073 6903 12267 6955
rect 11759 6847 12267 6903
rect 11759 6795 11805 6847
rect 11857 6795 11913 6847
rect 11965 6795 12021 6847
rect 12073 6795 12267 6847
rect 11759 6739 12267 6795
rect 11759 6687 11805 6739
rect 11857 6687 11913 6739
rect 11965 6687 12021 6739
rect 12073 6687 12267 6739
rect 11759 6631 12267 6687
rect 11759 6579 11805 6631
rect 11857 6579 11913 6631
rect 11965 6579 12021 6631
rect 12073 6579 12267 6631
rect 11759 6523 12267 6579
rect 11759 6471 11805 6523
rect 11857 6471 11913 6523
rect 11965 6471 12021 6523
rect 12073 6471 12267 6523
rect 11759 6415 12267 6471
rect 11759 6363 11805 6415
rect 11857 6363 11913 6415
rect 11965 6363 12021 6415
rect 12073 6363 12267 6415
rect 11759 6307 12267 6363
rect 11759 6255 11805 6307
rect 11857 6255 11913 6307
rect 11965 6255 12021 6307
rect 12073 6255 12267 6307
rect 11759 6199 12267 6255
rect 11759 6147 11805 6199
rect 11857 6147 11913 6199
rect 11965 6147 12021 6199
rect 12073 6147 12267 6199
rect 11759 6091 12267 6147
rect 11759 6039 11805 6091
rect 11857 6039 11913 6091
rect 11965 6039 12021 6091
rect 12073 6039 12267 6091
rect 11759 5983 12267 6039
rect 11759 5931 11805 5983
rect 11857 5931 11913 5983
rect 11965 5931 12021 5983
rect 12073 5931 12267 5983
rect 11759 5875 12267 5931
rect 11759 5823 11805 5875
rect 11857 5823 11913 5875
rect 11965 5823 12021 5875
rect 12073 5823 12267 5875
rect 11759 5767 12267 5823
rect 11759 5715 11805 5767
rect 11857 5715 11913 5767
rect 11965 5715 12021 5767
rect 12073 5715 12267 5767
rect 11759 5659 12267 5715
rect 11759 5607 11805 5659
rect 11857 5607 11913 5659
rect 11965 5607 12021 5659
rect 12073 5607 12267 5659
rect 11759 5551 12267 5607
rect 11759 5499 11805 5551
rect 11857 5499 11913 5551
rect 11965 5499 12021 5551
rect 12073 5499 12267 5551
rect 11759 5443 12267 5499
rect 11759 5391 11805 5443
rect 11857 5391 11913 5443
rect 11965 5391 12021 5443
rect 12073 5391 12267 5443
rect 11759 5335 12267 5391
rect 11759 5283 11805 5335
rect 11857 5283 11913 5335
rect 11965 5283 12021 5335
rect 12073 5283 12267 5335
rect 11759 5227 12267 5283
rect 11759 5175 11805 5227
rect 11857 5175 11913 5227
rect 11965 5175 12021 5227
rect 12073 5175 12267 5227
rect 11759 5119 12267 5175
rect 11759 5067 11805 5119
rect 11857 5067 11913 5119
rect 11965 5067 12021 5119
rect 12073 5067 12267 5119
rect 11759 5011 12267 5067
rect 11759 4959 11805 5011
rect 11857 4959 11913 5011
rect 11965 4959 12021 5011
rect 12073 4959 12267 5011
rect 11759 4903 12267 4959
rect 11759 4851 11805 4903
rect 11857 4851 11913 4903
rect 11965 4851 12021 4903
rect 12073 4851 12267 4903
rect 11759 4795 12267 4851
rect 11759 4743 11805 4795
rect 11857 4743 11913 4795
rect 11965 4743 12021 4795
rect 12073 4743 12267 4795
rect 11759 4687 12267 4743
rect 11759 4635 11805 4687
rect 11857 4635 11913 4687
rect 11965 4635 12021 4687
rect 12073 4635 12267 4687
rect 11759 4579 12267 4635
rect 11759 4527 11805 4579
rect 11857 4527 11913 4579
rect 11965 4527 12021 4579
rect 12073 4527 12267 4579
rect 11759 4471 12267 4527
rect 11759 4419 11805 4471
rect 11857 4419 11913 4471
rect 11965 4419 12021 4471
rect 12073 4419 12267 4471
rect 11759 4363 12267 4419
rect 11759 4311 11805 4363
rect 11857 4311 11913 4363
rect 11965 4311 12021 4363
rect 12073 4311 12267 4363
rect 11759 4255 12267 4311
rect 11759 4203 11805 4255
rect 11857 4203 11913 4255
rect 11965 4203 12021 4255
rect 12073 4203 12267 4255
rect 11759 4147 12267 4203
rect 11759 4095 11805 4147
rect 11857 4095 11913 4147
rect 11965 4095 12021 4147
rect 12073 4095 12267 4147
rect 11759 4039 12267 4095
rect 11759 3987 11805 4039
rect 11857 3987 11913 4039
rect 11965 3987 12021 4039
rect 12073 3987 12267 4039
rect 11759 3931 12267 3987
rect 11759 3879 11805 3931
rect 11857 3879 11913 3931
rect 11965 3879 12021 3931
rect 12073 3879 12267 3931
rect 11759 3823 12267 3879
rect 11759 3771 11805 3823
rect 11857 3771 11913 3823
rect 11965 3771 12021 3823
rect 12073 3771 12267 3823
rect 11759 3715 12267 3771
rect 11759 3663 11805 3715
rect 11857 3663 11913 3715
rect 11965 3663 12021 3715
rect 12073 3663 12267 3715
rect 11759 3607 12267 3663
rect 11759 3555 11805 3607
rect 11857 3555 11913 3607
rect 11965 3555 12021 3607
rect 12073 3555 12267 3607
rect 11759 3499 12267 3555
rect 11759 3447 11805 3499
rect 11857 3447 11913 3499
rect 11965 3447 12021 3499
rect 12073 3447 12267 3499
rect 11759 3391 12267 3447
rect 11759 3339 11805 3391
rect 11857 3339 11913 3391
rect 11965 3339 12021 3391
rect 12073 3339 12267 3391
rect 11759 3283 12267 3339
rect 11759 3231 11805 3283
rect 11857 3231 11913 3283
rect 11965 3231 12021 3283
rect 12073 3231 12267 3283
rect 11759 3175 12267 3231
rect 11759 3123 11805 3175
rect 11857 3123 11913 3175
rect 11965 3123 12021 3175
rect 12073 3123 12267 3175
rect 11759 3067 12267 3123
rect 11759 3015 11805 3067
rect 11857 3015 11913 3067
rect 11965 3015 12021 3067
rect 12073 3015 12267 3067
rect 11759 2959 12267 3015
rect 11759 2907 11805 2959
rect 11857 2907 11913 2959
rect 11965 2907 12021 2959
rect 12073 2907 12267 2959
rect 11759 2851 12267 2907
rect 11759 2799 11805 2851
rect 11857 2799 11913 2851
rect 11965 2799 12021 2851
rect 12073 2799 12267 2851
rect 11759 2743 12267 2799
rect 11759 2691 11805 2743
rect 11857 2691 11913 2743
rect 11965 2691 12021 2743
rect 12073 2691 12267 2743
rect 11759 2635 12267 2691
rect 11759 2583 11805 2635
rect 11857 2583 11913 2635
rect 11965 2583 12021 2635
rect 12073 2583 12267 2635
rect 11759 2527 12267 2583
rect 11759 2475 11805 2527
rect 11857 2475 11913 2527
rect 11965 2475 12021 2527
rect 12073 2475 12267 2527
rect 11759 2419 12267 2475
rect 11759 2367 11805 2419
rect 11857 2367 11913 2419
rect 11965 2367 12021 2419
rect 12073 2367 12267 2419
rect 11759 2311 12267 2367
rect 11759 2259 11805 2311
rect 11857 2259 11913 2311
rect 11965 2259 12021 2311
rect 12073 2259 12267 2311
rect 11759 2203 12267 2259
rect 11759 2151 11805 2203
rect 11857 2151 11913 2203
rect 11965 2151 12021 2203
rect 12073 2151 12267 2203
rect 11759 2095 12267 2151
rect 11759 2043 11805 2095
rect 11857 2043 11913 2095
rect 11965 2043 12021 2095
rect 12073 2043 12267 2095
rect 11759 1987 12267 2043
rect 11759 1935 11805 1987
rect 11857 1935 11913 1987
rect 11965 1935 12021 1987
rect 12073 1935 12267 1987
rect 11759 1879 12267 1935
rect 11759 1827 11805 1879
rect 11857 1827 11913 1879
rect 11965 1827 12021 1879
rect 12073 1827 12267 1879
rect 11759 1771 12267 1827
rect 11759 1719 11805 1771
rect 11857 1719 11913 1771
rect 11965 1719 12021 1771
rect 12073 1719 12267 1771
rect 11759 1663 12267 1719
rect 11759 1611 11805 1663
rect 11857 1611 11913 1663
rect 11965 1611 12021 1663
rect 12073 1611 12267 1663
rect 11759 1555 12267 1611
rect 11759 1503 11805 1555
rect 11857 1503 11913 1555
rect 11965 1503 12021 1555
rect 12073 1503 12267 1555
rect 11759 1447 12267 1503
rect 11759 1395 11805 1447
rect 11857 1395 11913 1447
rect 11965 1395 12021 1447
rect 12073 1395 12267 1447
rect 11759 1339 12267 1395
rect 11759 1287 11805 1339
rect 11857 1287 11913 1339
rect 11965 1287 12021 1339
rect 12073 1287 12267 1339
rect 11759 1231 12267 1287
rect 11759 1179 11805 1231
rect 11857 1179 11913 1231
rect 11965 1179 12021 1231
rect 12073 1179 12267 1231
rect 11759 1123 12267 1179
rect 11759 1071 11805 1123
rect 11857 1071 11913 1123
rect 11965 1071 12021 1123
rect 12073 1071 12267 1123
rect 11759 1015 12267 1071
rect 11759 963 11805 1015
rect 11857 963 11913 1015
rect 11965 963 12021 1015
rect 12073 963 12267 1015
rect 11759 907 12267 963
rect 11759 855 11805 907
rect 11857 855 11913 907
rect 11965 855 12021 907
rect 12073 855 12267 907
rect 11759 799 12267 855
rect 11759 747 11805 799
rect 11857 747 11913 799
rect 11965 747 12021 799
rect 12073 747 12267 799
rect 11759 691 12267 747
rect 11759 639 11805 691
rect 11857 639 11913 691
rect 11965 639 12021 691
rect 12073 639 12267 691
rect 11759 583 12267 639
rect 11759 531 11805 583
rect 11857 531 11913 583
rect 11965 531 12021 583
rect 12073 531 12267 583
rect 11759 475 12267 531
rect 11759 423 11805 475
rect 11857 423 11913 475
rect 11965 423 12021 475
rect 12073 423 12267 475
rect 11759 367 12267 423
rect 11759 315 11805 367
rect 11857 315 11913 367
rect 11965 315 12021 367
rect 12073 315 12267 367
rect 11759 259 12267 315
rect 11759 207 11805 259
rect 11857 207 11913 259
rect 11965 207 12021 259
rect 12073 207 12267 259
rect 11759 151 12267 207
rect 11759 99 11805 151
rect 11857 99 11913 151
rect 11965 99 12021 151
rect 12073 99 12267 151
rect 11759 43 12267 99
use M1_NWELL_CDNS_40661953145217  M1_NWELL_CDNS_40661953145217_0
timestamp 1698431365
transform 1 0 11379 0 1 2825
box 0 0 1 1
use M1_NWELL_CDNS_40661953145217  M1_NWELL_CDNS_40661953145217_1
timestamp 1698431365
transform 1 0 11379 0 1 1421
box 0 0 1 1
use M1_NWELL_CDNS_40661953145217  M1_NWELL_CDNS_40661953145217_2
timestamp 1698431365
transform 1 0 11379 0 1 4229
box 0 0 1 1
use M1_NWELL_CDNS_40661953145217  M1_NWELL_CDNS_40661953145217_3
timestamp 1698431365
transform 1 0 11379 0 1 5633
box 0 0 1 1
use M1_NWELL_CDNS_40661953145217  M1_NWELL_CDNS_40661953145217_4
timestamp 1698431365
transform 1 0 883 0 1 1421
box 0 0 1 1
use M1_NWELL_CDNS_40661953145217  M1_NWELL_CDNS_40661953145217_5
timestamp 1698431365
transform 1 0 883 0 1 2825
box 0 0 1 1
use M1_NWELL_CDNS_40661953145217  M1_NWELL_CDNS_40661953145217_6
timestamp 1698431365
transform 1 0 883 0 1 4229
box 0 0 1 1
use M1_NWELL_CDNS_40661953145217  M1_NWELL_CDNS_40661953145217_7
timestamp 1698431365
transform 1 0 883 0 1 5633
box 0 0 1 1
use M1_NWELL_CDNS_40661953145397  M1_NWELL_CDNS_40661953145397_0
timestamp 1698431365
transform 1 0 6131 0 1 4931
box 0 0 1 1
use M1_NWELL_CDNS_40661953145397  M1_NWELL_CDNS_40661953145397_1
timestamp 1698431365
transform 1 0 6131 0 1 3527
box 0 0 1 1
use M1_NWELL_CDNS_40661953145397  M1_NWELL_CDNS_40661953145397_2
timestamp 1698431365
transform 1 0 6131 0 1 2123
box 0 0 1 1
use M1_NWELL_CDNS_40661953145398  M1_NWELL_CDNS_40661953145398_0
timestamp 1698431365
transform 1 0 6131 0 1 6335
box 0 0 1 1
use M1_NWELL_CDNS_40661953145398  M1_NWELL_CDNS_40661953145398_1
timestamp 1698431365
transform 1 0 6131 0 1 719
box 0 0 1 1
use M1_NWELL_CDNS_40661953145399  M1_NWELL_CDNS_40661953145399_0
timestamp 1698431365
transform 1 0 6131 0 1 3373
box 0 0 1 1
use M1_NWELL_CDNS_40661953145399  M1_NWELL_CDNS_40661953145399_1
timestamp 1698431365
transform 1 0 6131 0 1 873
box 0 0 1 1
use M1_NWELL_CDNS_40661953145399  M1_NWELL_CDNS_40661953145399_2
timestamp 1698431365
transform 1 0 6131 0 1 2277
box 0 0 1 1
use M1_NWELL_CDNS_40661953145399  M1_NWELL_CDNS_40661953145399_3
timestamp 1698431365
transform 1 0 6131 0 1 1969
box 0 0 1 1
use M1_NWELL_CDNS_40661953145399  M1_NWELL_CDNS_40661953145399_4
timestamp 1698431365
transform 1 0 6131 0 1 3681
box 0 0 1 1
use M1_NWELL_CDNS_40661953145399  M1_NWELL_CDNS_40661953145399_5
timestamp 1698431365
transform 1 0 6131 0 1 5085
box 0 0 1 1
use M1_NWELL_CDNS_40661953145399  M1_NWELL_CDNS_40661953145399_6
timestamp 1698431365
transform 1 0 6131 0 1 6181
box 0 0 1 1
use M1_NWELL_CDNS_40661953145399  M1_NWELL_CDNS_40661953145399_7
timestamp 1698431365
transform 1 0 6131 0 1 4777
box 0 0 1 1
use M1_NWELL_CDNS_40661953145400  M1_NWELL_CDNS_40661953145400_0
timestamp 1698431365
transform 1 0 11533 0 1 3527
box 0 0 1 1
use M1_NWELL_CDNS_40661953145400  M1_NWELL_CDNS_40661953145400_1
timestamp 1698431365
transform 1 0 729 0 1 3527
box 0 0 1 1
use M1_NWELL_CDNS_40661953145407  M1_NWELL_CDNS_40661953145407_0
timestamp 1698431365
transform 1 0 6131 0 1 7684
box 0 0 1 1
use M1_NWELL_CDNS_40661953145407  M1_NWELL_CDNS_40661953145407_1
timestamp 1698431365
transform 1 0 6131 0 1 14184
box 0 0 1 1
use M1_NWELL_CDNS_40661953145412  M1_NWELL_CDNS_40661953145412_0
timestamp 1698431365
transform 1 0 277 0 1 10934
box 0 0 1 1
use M1_NWELL_CDNS_40661953145412  M1_NWELL_CDNS_40661953145412_1
timestamp 1698431365
transform 1 0 11985 0 1 10934
box 0 0 1 1
use M1_PSUB_CDNS_40661953145401  M1_PSUB_CDNS_40661953145401_0
timestamp 1698431365
transform 1 0 6131 0 1 8126
box 0 0 1 1
use M1_PSUB_CDNS_40661953145401  M1_PSUB_CDNS_40661953145401_1
timestamp 1698431365
transform 1 0 6131 0 1 13742
box 0 0 1 1
use M1_PSUB_CDNS_40661953145402  M1_PSUB_CDNS_40661953145402_0
timestamp 1698431365
transform 1 0 729 0 1 10934
box 0 0 1 1
use M1_PSUB_CDNS_40661953145402  M1_PSUB_CDNS_40661953145402_1
timestamp 1698431365
transform 1 0 11533 0 1 10934
box 0 0 1 1
use M1_PSUB_CDNS_40661953145403  M1_PSUB_CDNS_40661953145403_0
timestamp 1698431365
transform 1 0 6131 0 1 13588
box 0 0 1 1
use M1_PSUB_CDNS_40661953145403  M1_PSUB_CDNS_40661953145403_1
timestamp 1698431365
transform 1 0 6131 0 1 12184
box 0 0 1 1
use M1_PSUB_CDNS_40661953145403  M1_PSUB_CDNS_40661953145403_2
timestamp 1698431365
transform 1 0 6131 0 1 11088
box 0 0 1 1
use M1_PSUB_CDNS_40661953145403  M1_PSUB_CDNS_40661953145403_3
timestamp 1698431365
transform 1 0 6131 0 1 10780
box 0 0 1 1
use M1_PSUB_CDNS_40661953145403  M1_PSUB_CDNS_40661953145403_4
timestamp 1698431365
transform 1 0 6131 0 1 9684
box 0 0 1 1
use M1_PSUB_CDNS_40661953145403  M1_PSUB_CDNS_40661953145403_5
timestamp 1698431365
transform 1 0 6131 0 1 9376
box 0 0 1 1
use M1_PSUB_CDNS_40661953145403  M1_PSUB_CDNS_40661953145403_6
timestamp 1698431365
transform 1 0 6131 0 1 12492
box 0 0 1 1
use M1_PSUB_CDNS_40661953145403  M1_PSUB_CDNS_40661953145403_7
timestamp 1698431365
transform 1 0 6131 0 1 8280
box 0 0 1 1
use M1_PSUB_CDNS_40661953145404  M1_PSUB_CDNS_40661953145404_0
timestamp 1698431365
transform 1 0 883 0 1 13040
box 0 0 1 1
use M1_PSUB_CDNS_40661953145404  M1_PSUB_CDNS_40661953145404_1
timestamp 1698431365
transform 1 0 883 0 1 11636
box 0 0 1 1
use M1_PSUB_CDNS_40661953145404  M1_PSUB_CDNS_40661953145404_2
timestamp 1698431365
transform 1 0 883 0 1 10232
box 0 0 1 1
use M1_PSUB_CDNS_40661953145404  M1_PSUB_CDNS_40661953145404_3
timestamp 1698431365
transform 1 0 883 0 1 8828
box 0 0 1 1
use M1_PSUB_CDNS_40661953145404  M1_PSUB_CDNS_40661953145404_4
timestamp 1698431365
transform 1 0 11379 0 1 13040
box 0 0 1 1
use M1_PSUB_CDNS_40661953145404  M1_PSUB_CDNS_40661953145404_5
timestamp 1698431365
transform 1 0 11379 0 1 11636
box 0 0 1 1
use M1_PSUB_CDNS_40661953145404  M1_PSUB_CDNS_40661953145404_6
timestamp 1698431365
transform 1 0 11379 0 1 10232
box 0 0 1 1
use M1_PSUB_CDNS_40661953145404  M1_PSUB_CDNS_40661953145404_7
timestamp 1698431365
transform 1 0 11379 0 1 8828
box 0 0 1 1
use M1_PSUB_CDNS_40661953145405  M1_PSUB_CDNS_40661953145405_0
timestamp 1698431365
transform 1 0 6131 0 1 12338
box 0 0 1 1
use M1_PSUB_CDNS_40661953145405  M1_PSUB_CDNS_40661953145405_1
timestamp 1698431365
transform 1 0 6131 0 1 10934
box 0 0 1 1
use M1_PSUB_CDNS_40661953145405  M1_PSUB_CDNS_40661953145405_2
timestamp 1698431365
transform 1 0 6131 0 1 9530
box 0 0 1 1
use M1_PSUB_CDNS_40661953145409  M1_PSUB_CDNS_40661953145409_0
timestamp 1698431365
transform 1 0 11985 0 1 3527
box 0 0 1 1
use M1_PSUB_CDNS_40661953145409  M1_PSUB_CDNS_40661953145409_1
timestamp 1698431365
transform 1 0 277 0 1 3527
box 0 0 1 1
use M1_PSUB_CDNS_40661953145411  M1_PSUB_CDNS_40661953145411_0
timestamp 1698431365
transform 1 0 6131 0 1 6777
box 0 0 1 1
use M1_PSUB_CDNS_40661953145411  M1_PSUB_CDNS_40661953145411_1
timestamp 1698431365
transform 1 0 6131 0 1 277
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_0
timestamp 1698431365
transform -1 0 9741 0 1 2123
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_1
timestamp 1698431365
transform -1 0 7469 0 1 2123
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_2
timestamp 1698431365
transform -1 0 7469 0 1 3527
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_3
timestamp 1698431365
transform -1 0 9741 0 1 4931
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_4
timestamp 1698431365
transform -1 0 7469 0 1 4931
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_5
timestamp 1698431365
transform -1 0 9741 0 1 3527
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_6
timestamp 1698431365
transform 1 0 4793 0 1 4931
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_7
timestamp 1698431365
transform 1 0 4793 0 1 3527
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_8
timestamp 1698431365
transform 1 0 4793 0 1 2123
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_9
timestamp 1698431365
transform 1 0 2521 0 1 4931
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_10
timestamp 1698431365
transform 1 0 2521 0 1 3527
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_11
timestamp 1698431365
transform 1 0 2521 0 1 2123
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_12
timestamp 1698431365
transform 1 0 1385 0 1 12338
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_13
timestamp 1698431365
transform 1 0 1385 0 1 9530
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_14
timestamp 1698431365
transform 1 0 3657 0 1 12338
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_15
timestamp 1698431365
transform 1 0 3657 0 1 10934
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_16
timestamp 1698431365
transform 1 0 3657 0 1 9530
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_17
timestamp 1698431365
transform 1 0 1385 0 1 10934
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_18
timestamp 1698431365
transform -1 0 8605 0 1 9530
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_19
timestamp 1698431365
transform -1 0 8605 0 1 12338
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_20
timestamp 1698431365
transform -1 0 10877 0 1 10934
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_21
timestamp 1698431365
transform -1 0 10877 0 1 12338
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_22
timestamp 1698431365
transform -1 0 8605 0 1 10934
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_23
timestamp 1698431365
transform -1 0 10877 0 1 9530
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_0
timestamp 1698431365
transform -1 0 7469 0 1 6258
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_1
timestamp 1698431365
transform -1 0 9741 0 1 796
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_2
timestamp 1698431365
transform -1 0 7469 0 1 796
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_3
timestamp 1698431365
transform -1 0 9741 0 1 6258
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_4
timestamp 1698431365
transform 1 0 2521 0 1 6258
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_5
timestamp 1698431365
transform 1 0 4793 0 1 796
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_6
timestamp 1698431365
transform 1 0 4793 0 1 6258
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_7
timestamp 1698431365
transform 1 0 2521 0 1 796
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_8
timestamp 1698431365
transform 1 0 1385 0 1 8203
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_9
timestamp 1698431365
transform 1 0 1385 0 1 13665
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_10
timestamp 1698431365
transform 1 0 3657 0 1 8203
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_11
timestamp 1698431365
transform 1 0 3657 0 1 13665
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_12
timestamp 1698431365
transform -1 0 8605 0 1 13665
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_13
timestamp 1698431365
transform -1 0 10877 0 1 8203
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_14
timestamp 1698431365
transform -1 0 8605 0 1 8203
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_15
timestamp 1698431365
transform -1 0 10877 0 1 13665
box 0 0 1 1
use M2_M1_CDNS_40661953145385  M2_M1_CDNS_40661953145385_0
timestamp 1698431365
transform 1 0 5888 0 1 8203
box 0 0 1 1
use M2_M1_CDNS_40661953145385  M2_M1_CDNS_40661953145385_1
timestamp 1698431365
transform 1 0 5888 0 1 13665
box 0 0 1 1
use M2_M1_CDNS_40661953145385  M2_M1_CDNS_40661953145385_2
timestamp 1698431365
transform -1 0 6374 0 1 8203
box 0 0 1 1
use M2_M1_CDNS_40661953145385  M2_M1_CDNS_40661953145385_3
timestamp 1698431365
transform -1 0 6374 0 1 13665
box 0 0 1 1
use M2_M1_CDNS_40661953145386  M2_M1_CDNS_40661953145386_0
timestamp 1698431365
transform 1 0 5888 0 1 10934
box 0 0 1 1
use M2_M1_CDNS_40661953145386  M2_M1_CDNS_40661953145386_1
timestamp 1698431365
transform 1 0 5888 0 1 12338
box 0 0 1 1
use M2_M1_CDNS_40661953145386  M2_M1_CDNS_40661953145386_2
timestamp 1698431365
transform 1 0 5888 0 1 9530
box 0 0 1 1
use M2_M1_CDNS_40661953145386  M2_M1_CDNS_40661953145386_3
timestamp 1698431365
transform -1 0 6374 0 1 9530
box 0 0 1 1
use M2_M1_CDNS_40661953145386  M2_M1_CDNS_40661953145386_4
timestamp 1698431365
transform -1 0 6374 0 1 12338
box 0 0 1 1
use M2_M1_CDNS_40661953145386  M2_M1_CDNS_40661953145386_5
timestamp 1698431365
transform -1 0 6374 0 1 10934
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_0
timestamp 1698431365
transform 1 0 6901 0 1 1421
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_1
timestamp 1698431365
transform 1 0 10309 0 1 4229
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_2
timestamp 1698431365
transform 1 0 8037 0 1 4229
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_3
timestamp 1698431365
transform 1 0 9173 0 1 4229
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_4
timestamp 1698431365
transform 1 0 6901 0 1 2825
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_5
timestamp 1698431365
transform 1 0 10309 0 1 2825
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_6
timestamp 1698431365
transform 1 0 8037 0 1 2825
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_7
timestamp 1698431365
transform 1 0 9173 0 1 2825
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_8
timestamp 1698431365
transform 1 0 9173 0 1 5633
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_9
timestamp 1698431365
transform 1 0 8037 0 1 5633
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_10
timestamp 1698431365
transform 1 0 10309 0 1 5633
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_11
timestamp 1698431365
transform 1 0 6901 0 1 5633
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_12
timestamp 1698431365
transform 1 0 6901 0 1 4229
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_13
timestamp 1698431365
transform 1 0 9173 0 1 1421
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_14
timestamp 1698431365
transform 1 0 8037 0 1 1421
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_15
timestamp 1698431365
transform 1 0 10309 0 1 1421
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_16
timestamp 1698431365
transform 1 0 4225 0 1 4229
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_17
timestamp 1698431365
transform 1 0 5361 0 1 4229
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_18
timestamp 1698431365
transform 1 0 1953 0 1 4229
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_19
timestamp 1698431365
transform 1 0 3089 0 1 5633
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_20
timestamp 1698431365
transform 1 0 5361 0 1 5633
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_21
timestamp 1698431365
transform 1 0 1953 0 1 5633
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_22
timestamp 1698431365
transform 1 0 4225 0 1 5633
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_23
timestamp 1698431365
transform 1 0 4225 0 1 1421
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_24
timestamp 1698431365
transform 1 0 3089 0 1 1421
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_25
timestamp 1698431365
transform 1 0 5361 0 1 1421
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_26
timestamp 1698431365
transform 1 0 1953 0 1 2825
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_27
timestamp 1698431365
transform 1 0 5361 0 1 2825
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_28
timestamp 1698431365
transform 1 0 3089 0 1 2825
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_29
timestamp 1698431365
transform 1 0 3089 0 1 4229
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_30
timestamp 1698431365
transform 1 0 4225 0 1 2825
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_31
timestamp 1698431365
transform 1 0 1953 0 1 1421
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_32
timestamp 1698431365
transform 1 0 4225 0 1 8828
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_33
timestamp 1698431365
transform 1 0 1953 0 1 11636
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_34
timestamp 1698431365
transform 1 0 5361 0 1 11636
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_35
timestamp 1698431365
transform 1 0 3089 0 1 11636
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_36
timestamp 1698431365
transform 1 0 4225 0 1 11636
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_37
timestamp 1698431365
transform 1 0 1953 0 1 10232
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_38
timestamp 1698431365
transform 1 0 5361 0 1 10232
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_39
timestamp 1698431365
transform 1 0 3089 0 1 10232
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_40
timestamp 1698431365
transform 1 0 4225 0 1 10232
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_41
timestamp 1698431365
transform 1 0 1953 0 1 8828
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_42
timestamp 1698431365
transform 1 0 1953 0 1 13040
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_43
timestamp 1698431365
transform 1 0 5361 0 1 13040
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_44
timestamp 1698431365
transform 1 0 3089 0 1 13040
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_45
timestamp 1698431365
transform 1 0 4225 0 1 13040
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_46
timestamp 1698431365
transform 1 0 5361 0 1 8828
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_47
timestamp 1698431365
transform 1 0 3089 0 1 8828
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_48
timestamp 1698431365
transform 1 0 9173 0 1 8828
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_49
timestamp 1698431365
transform 1 0 8037 0 1 8828
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_50
timestamp 1698431365
transform 1 0 10309 0 1 8828
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_51
timestamp 1698431365
transform 1 0 6901 0 1 8828
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_52
timestamp 1698431365
transform 1 0 8037 0 1 13040
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_53
timestamp 1698431365
transform 1 0 6901 0 1 11636
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_54
timestamp 1698431365
transform 1 0 10309 0 1 11636
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_55
timestamp 1698431365
transform 1 0 8037 0 1 11636
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_56
timestamp 1698431365
transform 1 0 6901 0 1 10232
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_57
timestamp 1698431365
transform 1 0 10309 0 1 10232
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_58
timestamp 1698431365
transform 1 0 8037 0 1 10232
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_59
timestamp 1698431365
transform 1 0 9173 0 1 10232
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_60
timestamp 1698431365
transform 1 0 9173 0 1 11636
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_61
timestamp 1698431365
transform 1 0 6901 0 1 13040
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_62
timestamp 1698431365
transform 1 0 10309 0 1 13040
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_63
timestamp 1698431365
transform 1 0 9173 0 1 13040
box 0 0 1 1
use M2_M1_CDNS_40661953145406  M2_M1_CDNS_40661953145406_0
timestamp 1698431365
transform -1 0 11939 0 1 3527
box 0 0 1 1
use M2_M1_CDNS_40661953145406  M2_M1_CDNS_40661953145406_1
timestamp 1698431365
transform 1 0 323 0 1 3527
box 0 0 1 1
use M2_M1_CDNS_40661953145408  M2_M1_CDNS_40661953145408_0
timestamp 1698431365
transform -1 0 11445 0 1 3527
box 0 0 1 1
use M2_M1_CDNS_40661953145408  M2_M1_CDNS_40661953145408_1
timestamp 1698431365
transform 1 0 817 0 1 3527
box 0 0 1 1
use M2_M1_CDNS_40661953145410  M2_M1_CDNS_40661953145410_0
timestamp 1698431365
transform 1 0 11939 0 1 3527
box 0 0 1 1
use M2_M1_CDNS_40661953145413  M2_M1_CDNS_40661953145413_0
timestamp 1698431365
transform -1 0 8605 0 1 277
box 0 0 1 1
use M2_M1_CDNS_40661953145413  M2_M1_CDNS_40661953145413_1
timestamp 1698431365
transform -1 0 10877 0 1 277
box 0 0 1 1
use M2_M1_CDNS_40661953145413  M2_M1_CDNS_40661953145413_2
timestamp 1698431365
transform -1 0 8605 0 1 6777
box 0 0 1 1
use M2_M1_CDNS_40661953145413  M2_M1_CDNS_40661953145413_3
timestamp 1698431365
transform -1 0 10877 0 1 6777
box 0 0 1 1
use M2_M1_CDNS_40661953145413  M2_M1_CDNS_40661953145413_4
timestamp 1698431365
transform 1 0 3657 0 1 6777
box 0 0 1 1
use M2_M1_CDNS_40661953145413  M2_M1_CDNS_40661953145413_5
timestamp 1698431365
transform 1 0 3657 0 1 277
box 0 0 1 1
use M2_M1_CDNS_40661953145413  M2_M1_CDNS_40661953145413_6
timestamp 1698431365
transform 1 0 1385 0 1 6777
box 0 0 1 1
use M2_M1_CDNS_40661953145413  M2_M1_CDNS_40661953145413_7
timestamp 1698431365
transform 1 0 1385 0 1 277
box 0 0 1 1
use M2_M1_CDNS_40661953145413  M2_M1_CDNS_40661953145413_8
timestamp 1698431365
transform 1 0 817 0 1 14184
box 0 0 1 1
use M2_M1_CDNS_40661953145413  M2_M1_CDNS_40661953145413_9
timestamp 1698431365
transform 1 0 817 0 1 7684
box 0 0 1 1
use M2_M1_CDNS_40661953145413  M2_M1_CDNS_40661953145413_10
timestamp 1698431365
transform 1 0 2521 0 1 14184
box 0 0 1 1
use M2_M1_CDNS_40661953145413  M2_M1_CDNS_40661953145413_11
timestamp 1698431365
transform 1 0 2521 0 1 7684
box 0 0 1 1
use M2_M1_CDNS_40661953145413  M2_M1_CDNS_40661953145413_12
timestamp 1698431365
transform 1 0 4793 0 1 14184
box 0 0 1 1
use M2_M1_CDNS_40661953145413  M2_M1_CDNS_40661953145413_13
timestamp 1698431365
transform 1 0 4793 0 1 7684
box 0 0 1 1
use M2_M1_CDNS_40661953145413  M2_M1_CDNS_40661953145413_14
timestamp 1698431365
transform -1 0 7469 0 1 7684
box 0 0 1 1
use M2_M1_CDNS_40661953145413  M2_M1_CDNS_40661953145413_15
timestamp 1698431365
transform -1 0 9741 0 1 7684
box 0 0 1 1
use M2_M1_CDNS_40661953145413  M2_M1_CDNS_40661953145413_16
timestamp 1698431365
transform -1 0 11445 0 1 7684
box 0 0 1 1
use M2_M1_CDNS_40661953145413  M2_M1_CDNS_40661953145413_17
timestamp 1698431365
transform -1 0 7469 0 1 14184
box 0 0 1 1
use M2_M1_CDNS_40661953145413  M2_M1_CDNS_40661953145413_18
timestamp 1698431365
transform -1 0 11445 0 1 14184
box 0 0 1 1
use M2_M1_CDNS_40661953145413  M2_M1_CDNS_40661953145413_19
timestamp 1698431365
transform -1 0 9741 0 1 14184
box 0 0 1 1
use M2_M1_CDNS_40661953145414  M2_M1_CDNS_40661953145414_0
timestamp 1698431365
transform -1 0 6374 0 1 277
box 0 0 1 1
use M2_M1_CDNS_40661953145414  M2_M1_CDNS_40661953145414_1
timestamp 1698431365
transform -1 0 6374 0 1 6777
box 0 0 1 1
use M2_M1_CDNS_40661953145414  M2_M1_CDNS_40661953145414_2
timestamp 1698431365
transform 1 0 5888 0 1 277
box 0 0 1 1
use M2_M1_CDNS_40661953145414  M2_M1_CDNS_40661953145414_3
timestamp 1698431365
transform 1 0 5888 0 1 6777
box 0 0 1 1
use np_6p0_CDNS_4066195314553  np_6p0_CDNS_4066195314553_0
timestamp 1698431365
transform 0 -1 11131 1 0 9932
box 0 0 1 1
use np_6p0_CDNS_4066195314553  np_6p0_CDNS_4066195314553_1
timestamp 1698431365
transform 0 -1 11131 1 0 11336
box 0 0 1 1
use np_6p0_CDNS_4066195314553  np_6p0_CDNS_4066195314553_2
timestamp 1698431365
transform 0 -1 11131 1 0 12740
box 0 0 1 1
use np_6p0_CDNS_4066195314553  np_6p0_CDNS_4066195314553_3
timestamp 1698431365
transform 0 -1 11131 1 0 8528
box 0 0 1 1
use pn_6p0_CDNS_4066195314552  pn_6p0_CDNS_4066195314552_0
timestamp 1698431365
transform 0 -1 11131 1 0 5333
box 0 0 1 1
use pn_6p0_CDNS_4066195314552  pn_6p0_CDNS_4066195314552_1
timestamp 1698431365
transform 0 -1 11131 1 0 3929
box 0 0 1 1
use pn_6p0_CDNS_4066195314552  pn_6p0_CDNS_4066195314552_2
timestamp 1698431365
transform 0 -1 11131 1 0 2525
box 0 0 1 1
use pn_6p0_CDNS_4066195314552  pn_6p0_CDNS_4066195314552_3
timestamp 1698431365
transform 0 -1 11131 1 0 1121
box 0 0 1 1
<< properties >>
string GDS_END 1402478
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 1386050
string path 257.725 1411.000 257.725 -21.425 
<< end >>
