magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 352 534 870
<< pwell >>
rect -86 -86 534 352
<< metal1 >>
rect 0 724 448 844
rect 49 496 95 724
rect 49 60 95 208
rect 141 194 206 590
rect 252 120 319 674
rect 0 -60 448 60
<< labels >>
rlabel metal1 s 141 194 206 590 6 I
port 1 nsew default input
rlabel metal1 s 252 120 319 674 6 ZN
port 2 nsew default output
rlabel metal1 s 49 496 95 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 724 448 844 6 VDD
port 3 nsew power bidirectional abutment
rlabel nwell s -86 352 534 870 6 VNW
port 4 nsew power bidirectional
rlabel pwell s -86 -86 534 352 6 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 0 -60 448 60 8 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 208 6 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 448 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 817360
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 815228
<< end >>
