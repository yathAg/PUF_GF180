magic
tech gf180mcuD
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 352 2438 870
<< pwell >>
rect -86 -86 2438 352
<< mvnmos >>
rect 124 79 244 172
rect 384 93 504 172
rect 552 93 672 172
rect 776 93 896 172
rect 944 93 1064 172
rect 1204 79 1324 172
rect 1388 79 1508 172
rect 1796 139 1916 232
rect 2056 68 2176 232
<< mvpmos >>
rect 124 531 224 716
rect 384 590 484 716
rect 532 590 632 716
rect 736 590 836 716
rect 944 590 1044 716
rect 1204 531 1304 716
rect 1408 531 1508 716
rect 1796 531 1896 716
rect 2076 472 2176 716
<< mvndiff >>
rect 1708 204 1796 232
rect 36 152 124 172
rect 36 106 49 152
rect 95 106 124 152
rect 36 79 124 106
rect 244 152 384 172
rect 244 106 273 152
rect 319 106 384 152
rect 244 93 384 106
rect 504 93 552 172
rect 672 152 776 172
rect 672 106 701 152
rect 747 106 776 152
rect 672 93 776 106
rect 896 93 944 172
rect 1064 152 1204 172
rect 1064 106 1093 152
rect 1139 106 1204 152
rect 1064 93 1204 106
rect 244 79 324 93
rect 1124 79 1204 93
rect 1324 79 1388 172
rect 1508 152 1596 172
rect 1508 106 1537 152
rect 1583 106 1596 152
rect 1708 158 1721 204
rect 1767 158 1796 204
rect 1708 139 1796 158
rect 1916 204 2056 232
rect 1916 158 1945 204
rect 1991 158 2056 204
rect 1916 139 2056 158
rect 1508 79 1596 106
rect 1976 68 2056 139
rect 2176 204 2264 232
rect 2176 158 2205 204
rect 2251 158 2264 204
rect 2176 68 2264 158
<< mvpdiff >>
rect 36 665 124 716
rect 36 619 49 665
rect 95 619 124 665
rect 36 531 124 619
rect 224 703 384 716
rect 224 563 253 703
rect 299 590 384 703
rect 484 590 532 716
rect 632 665 736 716
rect 632 619 661 665
rect 707 619 736 665
rect 632 590 736 619
rect 836 590 944 716
rect 1044 665 1204 716
rect 1044 619 1073 665
rect 1119 619 1204 665
rect 1044 590 1204 619
rect 299 563 324 590
rect 224 531 324 563
rect 1124 531 1204 590
rect 1304 665 1408 716
rect 1304 619 1333 665
rect 1379 619 1408 665
rect 1304 531 1408 619
rect 1508 703 1596 716
rect 1508 563 1537 703
rect 1583 563 1596 703
rect 1508 531 1596 563
rect 1708 639 1796 716
rect 1708 593 1721 639
rect 1767 593 1796 639
rect 1708 531 1796 593
rect 1896 665 2076 716
rect 1896 531 2001 665
rect 1976 525 2001 531
rect 2047 525 2076 665
rect 1976 472 2076 525
rect 2176 665 2264 716
rect 2176 525 2205 665
rect 2251 525 2264 665
rect 2176 472 2264 525
<< mvndiffc >>
rect 49 106 95 152
rect 273 106 319 152
rect 701 106 747 152
rect 1093 106 1139 152
rect 1537 106 1583 152
rect 1721 158 1767 204
rect 1945 158 1991 204
rect 2205 158 2251 204
<< mvpdiffc >>
rect 49 619 95 665
rect 253 563 299 703
rect 661 619 707 665
rect 1073 619 1119 665
rect 1333 619 1379 665
rect 1537 563 1583 703
rect 1721 593 1767 639
rect 2001 525 2047 665
rect 2205 525 2251 665
<< polysilicon >>
rect 124 716 224 760
rect 384 716 484 760
rect 532 716 632 760
rect 736 716 836 760
rect 944 716 1044 760
rect 1204 716 1304 760
rect 1408 716 1508 760
rect 1796 716 1896 760
rect 2076 716 2176 760
rect 124 413 224 531
rect 384 414 484 590
rect 124 302 244 413
rect 124 256 175 302
rect 221 256 244 302
rect 124 172 244 256
rect 384 368 411 414
rect 457 368 484 414
rect 384 268 484 368
rect 532 516 632 590
rect 532 470 559 516
rect 605 470 632 516
rect 532 409 632 470
rect 736 516 836 590
rect 736 470 763 516
rect 809 470 836 516
rect 736 457 836 470
rect 944 516 1044 590
rect 944 470 981 516
rect 1027 470 1044 516
rect 944 467 1044 470
rect 532 363 896 409
rect 552 302 672 315
rect 384 172 504 268
rect 552 256 593 302
rect 639 256 672 302
rect 552 172 672 256
rect 776 172 896 363
rect 944 172 1064 467
rect 1204 444 1304 531
rect 1408 444 1508 531
rect 1204 291 1324 444
rect 1204 245 1241 291
rect 1287 245 1324 291
rect 1204 172 1324 245
rect 1388 415 1508 444
rect 1388 369 1411 415
rect 1457 369 1508 415
rect 1388 172 1508 369
rect 1796 418 1896 531
rect 1796 372 1809 418
rect 1855 404 1896 418
rect 2076 404 2176 472
rect 1855 372 1916 404
rect 1796 232 1916 372
rect 2056 358 2093 404
rect 2139 358 2176 404
rect 2056 232 2176 358
rect 124 35 244 79
rect 384 35 504 93
rect 552 35 672 93
rect 776 35 896 93
rect 944 35 1064 93
rect 1204 35 1324 79
rect 1388 35 1508 79
rect 1796 24 1916 139
rect 2056 24 2176 68
<< polycontact >>
rect 175 256 221 302
rect 411 368 457 414
rect 559 470 605 516
rect 763 470 809 516
rect 981 470 1027 516
rect 593 256 639 302
rect 1241 245 1287 291
rect 1411 369 1457 415
rect 1809 372 1855 418
rect 2093 358 2139 404
<< metal1 >>
rect 0 724 2352 844
rect 242 703 310 724
rect 38 665 106 676
rect 38 619 49 665
rect 95 619 106 665
rect 38 516 106 619
rect 242 563 253 703
rect 299 563 310 703
rect 1073 665 1119 724
rect 1526 703 1594 724
rect 632 619 661 665
rect 707 619 912 665
rect 700 516 809 559
rect 38 470 559 516
rect 605 470 632 516
rect 700 470 763 516
rect 38 152 106 470
rect 193 414 654 424
rect 193 368 411 414
rect 457 368 654 414
rect 193 358 654 368
rect 700 312 809 470
rect 156 302 809 312
rect 156 256 175 302
rect 221 256 593 302
rect 639 256 809 302
rect 156 248 809 256
rect 864 291 912 619
rect 1073 600 1119 619
rect 1333 665 1379 676
rect 1333 516 1379 619
rect 1526 563 1537 703
rect 1583 563 1594 703
rect 2001 665 2047 724
rect 1721 639 1767 650
rect 1721 525 1767 593
rect 962 470 981 516
rect 1027 470 1594 516
rect 1721 479 1951 525
rect 2001 506 2047 525
rect 2179 665 2326 676
rect 2179 525 2205 665
rect 2251 525 2326 665
rect 2179 506 2326 525
rect 1526 429 1594 470
rect 1008 415 1476 424
rect 1008 369 1411 415
rect 1457 369 1476 415
rect 1008 360 1476 369
rect 1526 418 1857 429
rect 1526 372 1809 418
rect 1855 372 1857 418
rect 1526 361 1857 372
rect 1905 404 1951 479
rect 864 245 1241 291
rect 1287 245 1306 291
rect 38 106 49 152
rect 95 106 106 152
rect 273 152 319 172
rect 864 152 912 245
rect 682 106 701 152
rect 747 106 912 152
rect 1093 152 1139 172
rect 1526 152 1594 361
rect 1905 358 2093 404
rect 2139 358 2150 404
rect 1905 311 1951 358
rect 1526 106 1537 152
rect 1583 106 1594 152
rect 1721 265 1951 311
rect 1721 204 1767 265
rect 1721 147 1767 158
rect 1945 204 1991 215
rect 2264 213 2326 506
rect 273 60 319 106
rect 1093 60 1139 106
rect 1945 60 1991 158
rect 2150 204 2326 213
rect 2150 158 2205 204
rect 2251 158 2326 204
rect 2150 120 2326 158
rect 0 -60 2352 60
<< labels >>
flabel metal1 s 2179 506 2326 676 0 FreeSans 400 0 0 0 Q
port 4 nsew default output
flabel metal1 s 1945 172 1991 215 0 FreeSans 400 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel metal1 s 1008 360 1476 424 0 FreeSans 400 0 0 0 SETN
port 3 nsew default input
flabel metal1 s 0 724 2352 844 0 FreeSans 400 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 193 358 654 424 0 FreeSans 400 0 0 0 D
port 1 nsew default input
flabel metal1 s 700 312 809 559 0 FreeSans 400 0 0 0 E
port 2 nsew clock input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 6 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 156 248 809 312 1 E
port 2 nsew clock input
rlabel metal1 s 2264 213 2326 506 1 Q
port 4 nsew default output
rlabel metal1 s 2150 120 2326 213 1 Q
port 4 nsew default output
rlabel metal1 s 2001 600 2047 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1526 600 1594 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1073 600 1119 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 242 600 310 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2001 563 2047 600 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1526 563 1594 600 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 242 563 310 600 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2001 506 2047 563 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1945 60 1991 172 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1093 60 1139 172 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 60 319 172 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 2352 60 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2352 784
string GDS_END 646628
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 641042
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
