magic
tech gf180mcuB
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 453 1206 1094
<< pwell >>
rect -86 -86 1206 453
<< mvnmos >>
rect 125 96 245 333
rect 293 96 413 333
rect 553 96 673 254
rect 777 96 897 254
<< mvpmos >>
rect 125 573 225 939
rect 329 573 429 939
rect 553 573 653 939
rect 777 573 877 939
<< mvndiff >>
rect 37 249 125 333
rect 37 109 50 249
rect 96 109 125 249
rect 37 96 125 109
rect 245 96 293 333
rect 413 254 493 333
rect 413 196 553 254
rect 413 150 442 196
rect 488 150 553 196
rect 413 96 553 150
rect 673 155 777 254
rect 673 109 702 155
rect 748 109 777 155
rect 673 96 777 109
rect 897 241 985 254
rect 897 195 926 241
rect 972 195 985 241
rect 897 96 985 195
<< mvpdiff >>
rect 37 861 125 939
rect 37 721 50 861
rect 96 721 125 861
rect 37 573 125 721
rect 225 726 329 939
rect 225 586 254 726
rect 300 586 329 726
rect 225 573 329 586
rect 429 861 553 939
rect 429 721 458 861
rect 504 721 553 861
rect 429 573 553 721
rect 653 573 777 939
rect 877 926 965 939
rect 877 786 906 926
rect 952 786 965 926
rect 877 573 965 786
<< mvndiffc >>
rect 50 109 96 249
rect 442 150 488 196
rect 702 109 748 155
rect 926 195 972 241
<< mvpdiffc >>
rect 50 721 96 861
rect 254 586 300 726
rect 458 721 504 861
rect 906 786 952 926
<< polysilicon >>
rect 125 939 225 983
rect 329 939 429 983
rect 553 939 653 983
rect 777 939 877 983
rect 125 508 225 573
rect 125 462 142 508
rect 188 462 225 508
rect 125 377 225 462
rect 329 412 429 573
rect 329 393 354 412
rect 125 333 245 377
rect 293 366 354 393
rect 400 393 429 412
rect 400 366 413 393
rect 293 333 413 366
rect 553 380 653 573
rect 553 334 585 380
rect 631 334 653 380
rect 553 298 653 334
rect 777 380 877 573
rect 777 334 809 380
rect 855 334 877 380
rect 777 298 877 334
rect 553 254 673 298
rect 777 254 897 298
rect 125 52 245 96
rect 293 52 413 96
rect 553 52 673 96
rect 777 52 897 96
<< polycontact >>
rect 142 462 188 508
rect 354 366 400 412
rect 585 334 631 380
rect 809 334 855 380
<< metal1 >>
rect 0 926 1120 1098
rect 0 918 906 926
rect 50 861 504 872
rect 96 826 458 861
rect 50 710 96 721
rect 254 726 306 766
rect 300 586 306 726
rect 952 918 1120 926
rect 906 775 952 786
rect 458 710 504 721
rect 23 508 194 519
rect 23 462 142 508
rect 188 462 194 508
rect 23 341 194 462
rect 50 249 96 260
rect 254 196 306 586
rect 354 412 539 423
rect 400 366 539 412
rect 354 242 539 366
rect 585 380 763 430
rect 631 334 763 380
rect 585 323 763 334
rect 809 380 983 430
rect 855 334 983 380
rect 809 323 983 334
rect 610 241 972 258
rect 610 212 926 241
rect 610 196 656 212
rect 254 150 442 196
rect 488 150 656 196
rect 926 184 972 195
rect 702 155 748 166
rect 50 90 96 109
rect 702 90 748 109
rect 0 -90 1120 90
<< labels >>
flabel metal1 s 354 242 539 423 0 FreeSans 200 0 0 0 A1
port 1 nsew default input
flabel metal1 s 23 341 194 519 0 FreeSans 200 0 0 0 A2
port 2 nsew default input
flabel metal1 s 585 323 763 430 0 FreeSans 200 0 0 0 B
port 3 nsew default input
flabel metal1 s 809 323 983 430 0 FreeSans 200 0 0 0 C
port 4 nsew default input
flabel metal1 s 0 918 1120 1098 0 FreeSans 200 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 50 166 96 260 0 FreeSans 200 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel metal1 s 254 258 306 766 0 FreeSans 200 0 0 0 ZN
port 5 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 7 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 8 nsew ground bidirectional
rlabel metal1 s 610 212 972 258 1 ZN
port 5 nsew default output
rlabel metal1 s 254 212 306 258 1 ZN
port 5 nsew default output
rlabel metal1 s 926 196 972 212 1 ZN
port 5 nsew default output
rlabel metal1 s 610 196 656 212 1 ZN
port 5 nsew default output
rlabel metal1 s 254 196 306 212 1 ZN
port 5 nsew default output
rlabel metal1 s 926 184 972 196 1 ZN
port 5 nsew default output
rlabel metal1 s 254 184 656 196 1 ZN
port 5 nsew default output
rlabel metal1 s 254 150 656 184 1 ZN
port 5 nsew default output
rlabel metal1 s 906 775 952 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 702 90 748 166 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 50 90 96 166 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 1120 90 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1120 1008
string GDS_END 1202566
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1198950
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
