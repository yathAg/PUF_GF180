magic
tech gf180mcuA
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 453 4790 1094
<< pwell >>
rect -86 -86 4790 453
<< mvnmos >>
rect 124 175 244 333
rect 348 175 468 333
rect 720 215 840 333
rect 964 215 1084 333
rect 1188 215 1308 333
rect 1356 215 1476 333
rect 1588 215 1708 333
rect 1816 215 1936 333
rect 2040 215 2160 333
rect 2300 183 2420 333
rect 2896 183 3016 333
rect 3156 215 3276 333
rect 3416 183 3536 333
rect 3784 69 3904 333
rect 4008 69 4128 333
rect 4232 69 4352 333
rect 4456 69 4576 333
<< mvpmos >>
rect 144 573 244 849
rect 348 573 448 849
rect 740 582 840 782
rect 944 582 1044 782
rect 1148 582 1248 782
rect 1296 582 1396 782
rect 1588 573 1688 773
rect 1836 651 1936 851
rect 2300 573 2400 773
rect 2568 573 2668 793
rect 2916 633 3016 853
rect 3176 575 3276 775
rect 3424 575 3524 795
rect 3804 573 3904 939
rect 4008 573 4108 939
rect 4212 573 4312 939
rect 4416 573 4516 939
<< mvndiff >>
rect 36 320 124 333
rect 36 274 49 320
rect 95 274 124 320
rect 36 175 124 274
rect 244 234 348 333
rect 244 188 273 234
rect 319 188 348 234
rect 244 175 348 188
rect 468 320 556 333
rect 468 274 497 320
rect 543 274 556 320
rect 468 175 556 274
rect 632 274 720 333
rect 632 228 645 274
rect 691 228 720 274
rect 632 215 720 228
rect 840 320 964 333
rect 840 274 869 320
rect 915 274 964 320
rect 840 215 964 274
rect 1084 320 1188 333
rect 1084 274 1113 320
rect 1159 274 1188 320
rect 1084 215 1188 274
rect 1308 215 1356 333
rect 1476 274 1588 333
rect 1476 228 1505 274
rect 1551 228 1588 274
rect 1476 215 1588 228
rect 1708 215 1816 333
rect 1936 320 2040 333
rect 1936 274 1965 320
rect 2011 274 2040 320
rect 1936 215 2040 274
rect 2160 320 2300 333
rect 2160 274 2225 320
rect 2271 274 2300 320
rect 2160 215 2300 274
rect 2220 183 2300 215
rect 2420 298 2508 333
rect 2420 252 2449 298
rect 2495 252 2508 298
rect 2420 183 2508 252
rect 2808 320 2896 333
rect 2808 274 2821 320
rect 2867 274 2896 320
rect 2808 183 2896 274
rect 3016 215 3156 333
rect 3276 274 3416 333
rect 3276 228 3305 274
rect 3351 228 3416 274
rect 3276 215 3416 228
rect 3016 183 3096 215
rect 3336 183 3416 215
rect 3536 320 3624 333
rect 3536 274 3565 320
rect 3611 274 3624 320
rect 3536 183 3624 274
rect 3696 222 3784 333
rect 3696 82 3709 222
rect 3755 82 3784 222
rect 3696 69 3784 82
rect 3904 320 4008 333
rect 3904 180 3933 320
rect 3979 180 4008 320
rect 3904 69 4008 180
rect 4128 222 4232 333
rect 4128 82 4157 222
rect 4203 82 4232 222
rect 4128 69 4232 82
rect 4352 314 4456 333
rect 4352 174 4381 314
rect 4427 174 4456 314
rect 4352 69 4456 174
rect 4576 222 4664 333
rect 4576 82 4605 222
rect 4651 82 4664 222
rect 4576 69 4664 82
<< mvpdiff >>
rect 56 739 144 849
rect 56 599 69 739
rect 115 599 144 739
rect 56 573 144 599
rect 244 836 348 849
rect 244 696 273 836
rect 319 696 348 836
rect 244 573 348 696
rect 448 726 536 849
rect 448 586 477 726
rect 523 586 536 726
rect 448 573 536 586
rect 608 829 680 842
rect 608 783 621 829
rect 667 783 680 829
rect 608 782 680 783
rect 1456 932 1528 945
rect 1456 792 1469 932
rect 1515 792 1528 932
rect 3716 926 3804 939
rect 1456 782 1528 792
rect 608 582 740 782
rect 840 641 944 782
rect 840 595 869 641
rect 915 595 944 641
rect 840 582 944 595
rect 1044 641 1148 782
rect 1044 595 1073 641
rect 1119 595 1148 641
rect 1044 582 1148 595
rect 1248 582 1296 782
rect 1396 773 1528 782
rect 1756 773 1836 851
rect 1396 582 1588 773
rect 1508 573 1588 582
rect 1688 651 1836 773
rect 1936 838 2024 851
rect 1936 792 1965 838
rect 2011 792 2024 838
rect 1936 651 2024 792
rect 2828 840 2916 853
rect 2828 794 2841 840
rect 2887 794 2916 840
rect 2488 773 2568 793
rect 1688 632 1776 651
rect 1688 586 1717 632
rect 1763 586 1776 632
rect 1688 573 1776 586
rect 2212 632 2300 773
rect 2212 586 2225 632
rect 2271 586 2300 632
rect 2212 573 2300 586
rect 2400 726 2568 773
rect 2400 586 2429 726
rect 2475 586 2568 726
rect 2400 573 2568 586
rect 2668 632 2756 793
rect 2828 633 2916 794
rect 3016 775 3096 853
rect 3336 782 3424 795
rect 3336 775 3349 782
rect 3016 645 3176 775
rect 3016 633 3101 645
rect 2668 586 2697 632
rect 2743 586 2756 632
rect 2668 573 2756 586
rect 3088 599 3101 633
rect 3147 599 3176 645
rect 3088 575 3176 599
rect 3276 642 3349 775
rect 3395 642 3424 782
rect 3276 575 3424 642
rect 3524 728 3612 795
rect 3524 588 3553 728
rect 3599 588 3612 728
rect 3524 575 3612 588
rect 3716 786 3729 926
rect 3775 786 3804 926
rect 3716 573 3804 786
rect 3904 726 4008 939
rect 3904 586 3933 726
rect 3979 586 4008 726
rect 3904 573 4008 586
rect 4108 926 4212 939
rect 4108 786 4137 926
rect 4183 786 4212 926
rect 4108 573 4212 786
rect 4312 726 4416 939
rect 4312 586 4341 726
rect 4387 586 4416 726
rect 4312 573 4416 586
rect 4516 926 4604 939
rect 4516 786 4545 926
rect 4591 786 4604 926
rect 4516 573 4604 786
<< mvndiffc >>
rect 49 274 95 320
rect 273 188 319 234
rect 497 274 543 320
rect 645 228 691 274
rect 869 274 915 320
rect 1113 274 1159 320
rect 1505 228 1551 274
rect 1965 274 2011 320
rect 2225 274 2271 320
rect 2449 252 2495 298
rect 2821 274 2867 320
rect 3305 228 3351 274
rect 3565 274 3611 320
rect 3709 82 3755 222
rect 3933 180 3979 320
rect 4157 82 4203 222
rect 4381 174 4427 314
rect 4605 82 4651 222
<< mvpdiffc >>
rect 69 599 115 739
rect 273 696 319 836
rect 477 586 523 726
rect 621 783 667 829
rect 1469 792 1515 932
rect 869 595 915 641
rect 1073 595 1119 641
rect 1965 792 2011 838
rect 2841 794 2887 840
rect 1717 586 1763 632
rect 2225 586 2271 632
rect 2429 586 2475 726
rect 2697 586 2743 632
rect 3101 599 3147 645
rect 3349 642 3395 782
rect 3553 588 3599 728
rect 3729 786 3775 926
rect 3933 586 3979 726
rect 4137 786 4183 926
rect 4341 586 4387 726
rect 4545 786 4591 926
<< polysilicon >>
rect 348 909 1044 949
rect 144 849 244 893
rect 348 849 448 909
rect 740 782 840 826
rect 944 782 1044 909
rect 1148 861 1248 874
rect 1148 815 1161 861
rect 1207 815 1248 861
rect 1148 782 1248 815
rect 1296 782 1396 826
rect 1836 913 3016 953
rect 3804 939 3904 983
rect 4008 939 4108 983
rect 4212 939 4312 983
rect 4416 939 4516 983
rect 1836 851 1936 913
rect 2300 852 2400 865
rect 2916 853 3016 913
rect 1588 773 1688 817
rect 144 494 244 573
rect 144 448 157 494
rect 203 448 244 494
rect 144 377 244 448
rect 124 333 244 377
rect 348 412 448 573
rect 348 366 361 412
rect 407 377 448 412
rect 740 523 840 582
rect 944 538 1044 582
rect 740 477 753 523
rect 799 477 840 523
rect 1148 490 1248 582
rect 740 377 840 477
rect 407 366 468 377
rect 348 333 468 366
rect 720 333 840 377
rect 964 450 1248 490
rect 1296 549 1396 582
rect 2300 806 2313 852
rect 2359 806 2400 852
rect 2300 773 2400 806
rect 2568 793 2668 837
rect 1296 503 1337 549
rect 1383 503 1396 549
rect 964 333 1084 450
rect 1296 425 1396 503
rect 1188 333 1308 377
rect 1356 333 1476 425
rect 1588 412 1688 573
rect 1588 366 1601 412
rect 1647 377 1688 412
rect 1836 377 1936 651
rect 3176 775 3276 819
rect 3424 795 3524 839
rect 2300 377 2400 573
rect 1647 366 1708 377
rect 1588 333 1708 366
rect 1816 333 1936 377
rect 2040 333 2160 377
rect 2300 333 2420 377
rect 124 131 244 175
rect 348 91 468 175
rect 720 171 840 215
rect 964 171 1084 215
rect 1188 91 1308 215
rect 1356 171 1476 215
rect 1588 171 1708 215
rect 1816 171 1936 215
rect 2040 91 2160 215
rect 2300 139 2420 183
rect 2568 91 2668 573
rect 2916 487 3016 633
rect 2916 441 2942 487
rect 2988 441 3016 487
rect 2916 377 3016 441
rect 3176 412 3276 575
rect 3176 377 3217 412
rect 2896 333 3016 377
rect 3156 366 3217 377
rect 3263 366 3276 412
rect 3424 542 3524 575
rect 3424 496 3437 542
rect 3483 496 3524 542
rect 3424 377 3524 496
rect 3804 465 3904 573
rect 4008 465 4108 573
rect 4212 465 4312 573
rect 4416 465 4516 573
rect 3804 451 4516 465
rect 3804 405 3817 451
rect 3863 405 4037 451
rect 4083 405 4239 451
rect 4285 405 4516 451
rect 3804 393 4516 405
rect 3804 377 3904 393
rect 3156 333 3276 366
rect 3416 333 3536 377
rect 3784 333 3904 377
rect 4008 333 4128 393
rect 4232 333 4352 393
rect 4456 377 4516 393
rect 4456 333 4576 377
rect 2896 139 3016 183
rect 3156 171 3276 215
rect 3416 139 3536 183
rect 348 51 2668 91
rect 3784 25 3904 69
rect 4008 25 4128 69
rect 4232 25 4352 69
rect 4456 25 4576 69
<< polycontact >>
rect 1161 815 1207 861
rect 157 448 203 494
rect 361 366 407 412
rect 753 477 799 523
rect 2313 806 2359 852
rect 1337 503 1383 549
rect 1601 366 1647 412
rect 2942 441 2988 487
rect 3217 366 3263 412
rect 3437 496 3483 542
rect 3817 405 3863 451
rect 4037 405 4083 451
rect 4239 405 4285 451
<< metal1 >>
rect 0 932 4704 1098
rect 0 918 1469 932
rect 273 836 319 918
rect 69 739 115 750
rect 621 829 667 918
rect 621 772 667 783
rect 1161 861 1207 872
rect 1161 744 1207 815
rect 1515 926 4704 932
rect 1515 918 3729 926
rect 1469 781 1515 792
rect 1965 838 2011 918
rect 1965 781 2011 792
rect 2313 852 2359 863
rect 273 685 319 696
rect 477 726 523 737
rect 704 735 1207 744
rect 2313 735 2359 806
rect 2841 840 2887 918
rect 2841 783 2887 794
rect 3349 782 3395 918
rect 704 726 2359 735
rect 115 599 407 634
rect 69 588 407 599
rect 142 494 315 542
rect 142 448 157 494
rect 203 448 315 494
rect 361 412 407 588
rect 361 337 407 366
rect 49 320 407 337
rect 95 291 407 320
rect 523 698 2359 726
rect 523 680 741 698
rect 1179 689 2359 698
rect 2429 726 3303 737
rect 523 586 543 680
rect 1073 641 1119 652
rect 858 634 869 641
rect 477 320 543 586
rect 610 595 869 634
rect 915 595 926 641
rect 610 588 926 595
rect 610 420 656 588
rect 702 523 905 542
rect 702 477 753 523
rect 799 477 905 523
rect 702 466 905 477
rect 610 374 915 420
rect 49 263 95 274
rect 477 274 497 320
rect 869 320 915 374
rect 477 263 543 274
rect 645 274 691 285
rect 273 234 319 245
rect 273 90 319 188
rect 869 263 915 274
rect 1073 412 1119 595
rect 1717 632 1763 643
rect 1717 549 1763 586
rect 2225 632 2271 643
rect 2225 549 2271 586
rect 1326 503 1337 549
rect 1383 503 2271 549
rect 2475 691 3303 726
rect 1073 366 1601 412
rect 1647 366 1658 412
rect 1073 320 1159 366
rect 1073 274 1113 320
rect 1965 320 2011 503
rect 2429 401 2475 586
rect 2697 632 3101 645
rect 2743 599 3101 632
rect 3147 599 3158 645
rect 2743 586 2867 599
rect 2697 575 2867 586
rect 1073 263 1159 274
rect 1505 274 1551 285
rect 645 90 691 228
rect 1965 263 2011 274
rect 2225 355 2475 401
rect 2225 320 2271 355
rect 2821 320 2867 575
rect 3257 542 3303 691
rect 3775 918 4137 926
rect 3729 775 3775 786
rect 4183 918 4545 926
rect 4137 775 4183 786
rect 4591 918 4704 926
rect 4545 775 4591 786
rect 3349 631 3395 642
rect 3553 728 3599 739
rect 2942 487 3106 542
rect 3257 496 3437 542
rect 3483 496 3494 542
rect 2988 441 3106 487
rect 2942 430 3106 441
rect 3553 464 3599 588
rect 3933 726 3979 737
rect 4341 726 4427 737
rect 3979 586 4341 621
rect 4387 586 4427 726
rect 3933 575 4427 586
rect 3553 451 4285 464
rect 3553 423 3817 451
rect 3217 412 3817 423
rect 3263 405 3817 412
rect 3863 405 4037 451
rect 4083 405 4239 451
rect 3263 392 4285 405
rect 3263 366 3611 392
rect 3217 355 3611 366
rect 2225 263 2271 274
rect 2449 298 2821 309
rect 2495 274 2821 298
rect 3565 320 3611 355
rect 4331 331 4427 575
rect 2495 252 2867 274
rect 2449 241 2867 252
rect 3305 274 3351 285
rect 1505 90 1551 228
rect 3565 263 3611 274
rect 3933 320 4427 331
rect 3305 90 3351 228
rect 3709 222 3755 233
rect 0 82 3709 90
rect 3979 314 4427 320
rect 3979 279 4381 314
rect 3933 169 3979 180
rect 4157 222 4203 233
rect 3755 82 4157 90
rect 4286 174 4381 279
rect 4286 163 4427 174
rect 4605 222 4651 233
rect 4203 82 4605 90
rect 4651 82 4704 90
rect 0 -90 4704 82
<< labels >>
flabel metal1 s 142 448 315 542 0 FreeSans 200 0 0 0 CLKN
port 3 nsew clock input
flabel metal1 s 702 466 905 542 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 4341 621 4427 737 0 FreeSans 200 0 0 0 Q
port 4 nsew default output
flabel metal1 s 2942 430 3106 542 0 FreeSans 200 0 0 0 SETN
port 2 nsew default input
flabel metal1 s 0 918 4704 1098 0 FreeSans 200 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 3305 245 3351 285 0 FreeSans 200 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 6 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 3933 621 3979 737 1 Q
port 4 nsew default output
rlabel metal1 s 3933 575 4427 621 1 Q
port 4 nsew default output
rlabel metal1 s 4331 331 4427 575 1 Q
port 4 nsew default output
rlabel metal1 s 3933 279 4427 331 1 Q
port 4 nsew default output
rlabel metal1 s 4286 169 4427 279 1 Q
port 4 nsew default output
rlabel metal1 s 3933 169 3979 279 1 Q
port 4 nsew default output
rlabel metal1 s 4286 163 4427 169 1 Q
port 4 nsew default output
rlabel metal1 s 4545 783 4591 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4137 783 4183 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3729 783 3775 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3349 783 3395 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2841 783 2887 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1965 783 2011 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1469 783 1515 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 621 783 667 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 783 319 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4545 781 4591 783 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4137 781 4183 783 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3729 781 3775 783 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3349 781 3395 783 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1965 781 2011 783 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1469 781 1515 783 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 621 781 667 783 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 781 319 783 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4545 775 4591 781 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4137 775 4183 781 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3729 775 3775 781 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3349 775 3395 781 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 621 775 667 781 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 775 319 781 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3349 772 3395 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 621 772 667 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 772 319 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3349 685 3395 772 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 685 319 772 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3349 631 3395 685 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1505 245 1551 285 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 645 245 691 285 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3305 233 3351 245 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1505 233 1551 245 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 645 233 691 245 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 233 319 245 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4605 90 4651 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4157 90 4203 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3709 90 3755 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3305 90 3351 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1505 90 1551 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 645 90 691 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 4704 90 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4704 1008
string GDS_END 580260
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 570398
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
