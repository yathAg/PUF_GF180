magic
tech gf180mcuA
timestamp 1698431365
<< properties >>
string GDS_END 5137074
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 5136494
<< end >>
