magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 453 1878 1094
<< pwell >>
rect -86 -86 1878 453
<< mvnmos >>
rect 124 69 244 333
rect 308 69 428 333
rect 539 69 659 333
rect 716 69 836 333
rect 940 69 1060 333
rect 1124 69 1244 333
rect 1348 69 1468 333
rect 1532 69 1652 333
<< mvpmos >>
rect 124 573 224 939
rect 328 573 428 939
rect 532 573 632 939
rect 736 573 836 939
rect 940 573 1040 939
rect 1144 573 1244 939
rect 1348 573 1448 939
rect 1552 573 1652 939
<< mvndiff >>
rect 36 222 124 333
rect 36 82 49 222
rect 95 82 124 222
rect 36 69 124 82
rect 244 69 308 333
rect 428 287 539 333
rect 428 147 464 287
rect 510 147 539 287
rect 428 69 539 147
rect 659 69 716 333
rect 836 128 940 333
rect 836 82 865 128
rect 911 82 940 128
rect 836 69 940 82
rect 1060 69 1124 333
rect 1244 287 1348 333
rect 1244 147 1273 287
rect 1319 147 1348 287
rect 1244 69 1348 147
rect 1468 69 1532 333
rect 1652 222 1740 333
rect 1652 82 1681 222
rect 1727 82 1740 222
rect 1652 69 1740 82
<< mvpdiff >>
rect 36 834 124 939
rect 36 694 49 834
rect 95 694 124 834
rect 36 573 124 694
rect 224 926 328 939
rect 224 786 253 926
rect 299 786 328 926
rect 224 573 328 786
rect 428 834 532 939
rect 428 694 457 834
rect 503 694 532 834
rect 428 573 532 694
rect 632 926 736 939
rect 632 786 661 926
rect 707 786 736 926
rect 632 573 736 786
rect 836 858 940 939
rect 836 812 865 858
rect 911 812 940 858
rect 836 573 940 812
rect 1040 755 1144 939
rect 1040 615 1069 755
rect 1115 615 1144 755
rect 1040 573 1144 615
rect 1244 847 1348 939
rect 1244 707 1273 847
rect 1319 707 1348 847
rect 1244 573 1348 707
rect 1448 755 1552 939
rect 1448 615 1477 755
rect 1523 615 1552 755
rect 1448 573 1552 615
rect 1652 847 1740 939
rect 1652 707 1681 847
rect 1727 707 1740 847
rect 1652 573 1740 707
<< mvndiffc >>
rect 49 82 95 222
rect 464 147 510 287
rect 865 82 911 128
rect 1273 147 1319 287
rect 1681 82 1727 222
<< mvpdiffc >>
rect 49 694 95 834
rect 253 786 299 926
rect 457 694 503 834
rect 661 786 707 926
rect 865 812 911 858
rect 1069 615 1115 755
rect 1273 707 1319 847
rect 1477 615 1523 755
rect 1681 707 1727 847
<< polysilicon >>
rect 124 939 224 983
rect 328 939 428 983
rect 532 939 632 983
rect 736 939 836 983
rect 940 939 1040 983
rect 1144 939 1244 983
rect 1348 939 1448 983
rect 1552 939 1652 983
rect 124 412 224 573
rect 124 366 142 412
rect 188 377 224 412
rect 328 513 428 573
rect 532 513 632 573
rect 328 441 632 513
rect 328 412 428 441
rect 328 377 361 412
rect 188 366 244 377
rect 124 333 244 366
rect 308 366 361 377
rect 407 366 428 412
rect 308 333 428 366
rect 539 377 632 441
rect 736 504 836 573
rect 736 458 749 504
rect 795 458 836 504
rect 736 377 836 458
rect 539 333 659 377
rect 716 333 836 377
rect 940 425 1040 573
rect 1144 465 1244 573
rect 1348 465 1448 573
rect 1144 452 1448 465
rect 940 412 1060 425
rect 940 366 1001 412
rect 1047 366 1060 412
rect 1144 406 1157 452
rect 1391 406 1448 452
rect 1144 393 1448 406
rect 1144 377 1244 393
rect 940 333 1060 366
rect 1124 333 1244 377
rect 1348 377 1448 393
rect 1552 523 1652 573
rect 1552 477 1580 523
rect 1626 477 1652 523
rect 1552 377 1652 477
rect 1348 333 1468 377
rect 1532 333 1652 377
rect 124 25 244 69
rect 308 25 428 69
rect 539 25 659 69
rect 716 25 836 69
rect 940 25 1060 69
rect 1124 25 1244 69
rect 1348 25 1468 69
rect 1532 25 1652 69
<< polycontact >>
rect 142 366 188 412
rect 361 366 407 412
rect 749 458 795 504
rect 1001 366 1047 412
rect 1157 406 1391 452
rect 1580 477 1626 523
<< metal1 >>
rect 0 926 1792 1098
rect 0 918 253 926
rect 49 834 95 845
rect 299 918 661 926
rect 253 775 299 786
rect 457 834 503 845
rect 95 694 457 729
rect 707 918 1792 926
rect 661 775 707 786
rect 759 812 865 858
rect 911 847 1727 858
rect 911 812 1273 847
rect 759 729 805 812
rect 503 694 805 729
rect 49 683 805 694
rect 869 755 1115 766
rect 869 615 1069 755
rect 1319 812 1681 847
rect 1273 696 1319 707
rect 1477 755 1523 766
rect 1115 615 1477 650
rect 1681 696 1727 707
rect 869 604 1523 615
rect 138 458 749 504
rect 795 458 806 504
rect 138 412 194 458
rect 138 366 142 412
rect 188 366 194 412
rect 138 354 194 366
rect 330 366 361 412
rect 407 366 418 412
rect 330 326 418 366
rect 244 242 418 326
rect 869 298 944 604
rect 990 523 1654 558
rect 990 512 1580 523
rect 990 412 1102 512
rect 1572 477 1580 512
rect 1626 477 1654 523
rect 990 366 1001 412
rect 1047 366 1102 412
rect 1150 452 1442 463
rect 1150 406 1157 452
rect 1391 406 1442 452
rect 1572 436 1654 477
rect 1150 344 1442 406
rect 464 287 510 298
rect 49 222 95 233
rect 0 82 49 90
rect 868 221 944 298
rect 1273 287 1319 298
rect 510 175 1273 221
rect 464 136 510 147
rect 1273 136 1319 147
rect 1681 222 1727 233
rect 854 90 865 128
rect 95 82 865 90
rect 911 90 922 128
rect 911 82 1681 90
rect 1727 82 1792 90
rect 0 -90 1792 82
<< labels >>
flabel metal1 s 1150 344 1442 463 0 FreeSans 200 0 0 0 A1
port 1 nsew default input
flabel metal1 s 990 512 1654 558 0 FreeSans 200 0 0 0 A2
port 2 nsew default input
flabel metal1 s 330 326 418 412 0 FreeSans 200 0 0 0 B1
port 3 nsew default input
flabel metal1 s 138 458 806 504 0 FreeSans 200 0 0 0 B2
port 4 nsew default input
flabel metal1 s 0 918 1792 1098 0 FreeSans 200 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 1681 128 1727 233 0 FreeSans 200 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel metal1 s 1477 650 1523 766 0 FreeSans 200 0 0 0 ZN
port 5 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 7 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 8 nsew ground bidirectional
rlabel metal1 s 1572 436 1654 512 1 A2
port 2 nsew default input
rlabel metal1 s 990 436 1102 512 1 A2
port 2 nsew default input
rlabel metal1 s 990 366 1102 436 1 A2
port 2 nsew default input
rlabel metal1 s 244 242 418 326 1 B1
port 3 nsew default input
rlabel metal1 s 138 354 194 458 1 B2
port 4 nsew default input
rlabel metal1 s 869 650 1115 766 1 ZN
port 5 nsew default output
rlabel metal1 s 869 604 1523 650 1 ZN
port 5 nsew default output
rlabel metal1 s 869 298 944 604 1 ZN
port 5 nsew default output
rlabel metal1 s 1273 221 1319 298 1 ZN
port 5 nsew default output
rlabel metal1 s 868 221 944 298 1 ZN
port 5 nsew default output
rlabel metal1 s 464 221 510 298 1 ZN
port 5 nsew default output
rlabel metal1 s 464 175 1319 221 1 ZN
port 5 nsew default output
rlabel metal1 s 1273 136 1319 175 1 ZN
port 5 nsew default output
rlabel metal1 s 464 136 510 175 1 ZN
port 5 nsew default output
rlabel metal1 s 661 775 707 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 253 775 299 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 49 128 95 233 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1681 90 1727 128 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 854 90 922 128 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 49 90 95 128 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 1792 90 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1792 1008
string GDS_END 1190580
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1185268
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
