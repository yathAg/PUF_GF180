magic
tech gf180mcuD
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 453 3670 1094
<< pwell >>
rect -86 -86 3670 453
<< mvnmos >>
rect 124 69 244 333
rect 348 69 468 333
rect 572 69 692 333
rect 796 69 916 333
rect 1020 69 1140 333
rect 1244 69 1364 333
rect 1468 69 1588 333
rect 1692 69 1812 333
rect 1922 69 2042 333
rect 2116 69 2236 333
rect 2340 69 2460 333
rect 2524 69 2644 333
rect 2748 69 2868 333
rect 2932 69 3052 333
rect 3156 69 3276 333
rect 3340 69 3460 333
<< mvpmos >>
rect 144 573 244 939
rect 368 573 468 939
rect 582 573 682 939
rect 806 573 906 939
rect 1030 573 1130 939
rect 1254 573 1354 939
rect 1478 573 1578 939
rect 1692 573 1792 939
rect 1932 647 2032 939
rect 2136 647 2236 939
rect 2340 647 2440 939
rect 2544 647 2644 939
rect 2748 647 2848 939
rect 2952 647 3052 939
rect 3156 647 3256 939
rect 3360 647 3460 939
<< mvndiff >>
rect 36 287 124 333
rect 36 147 49 287
rect 95 147 124 287
rect 36 69 124 147
rect 244 285 348 333
rect 244 239 273 285
rect 319 239 348 285
rect 244 69 348 239
rect 468 193 572 333
rect 468 147 497 193
rect 543 147 572 193
rect 468 69 572 147
rect 692 274 796 333
rect 692 228 721 274
rect 767 228 796 274
rect 692 69 796 228
rect 916 193 1020 333
rect 916 147 945 193
rect 991 147 1020 193
rect 916 69 1020 147
rect 1140 285 1244 333
rect 1140 239 1169 285
rect 1215 239 1244 285
rect 1140 69 1244 239
rect 1364 193 1468 333
rect 1364 147 1393 193
rect 1439 147 1468 193
rect 1364 69 1468 147
rect 1588 285 1692 333
rect 1588 239 1617 285
rect 1663 239 1692 285
rect 1588 69 1692 239
rect 1812 287 1922 333
rect 1812 147 1841 287
rect 1887 147 1922 287
rect 1812 69 1922 147
rect 2042 69 2116 333
rect 2236 242 2340 333
rect 2236 102 2265 242
rect 2311 102 2340 242
rect 2236 69 2340 102
rect 2460 69 2524 333
rect 2644 287 2748 333
rect 2644 147 2673 287
rect 2719 147 2748 287
rect 2644 69 2748 147
rect 2868 69 2932 333
rect 3052 287 3156 333
rect 3052 147 3081 287
rect 3127 147 3156 287
rect 3052 69 3156 147
rect 3276 69 3340 333
rect 3460 287 3548 333
rect 3460 147 3489 287
rect 3535 147 3548 287
rect 3460 69 3548 147
<< mvpdiff >>
rect 56 905 144 939
rect 56 765 69 905
rect 115 765 144 905
rect 56 573 144 765
rect 244 573 368 939
rect 468 861 582 939
rect 468 721 497 861
rect 543 721 582 861
rect 468 573 582 721
rect 682 573 806 939
rect 906 905 1030 939
rect 906 765 935 905
rect 981 765 1030 905
rect 906 573 1030 765
rect 1130 573 1254 939
rect 1354 861 1478 939
rect 1354 721 1383 861
rect 1429 721 1478 861
rect 1354 573 1478 721
rect 1578 573 1692 939
rect 1792 905 1932 939
rect 1792 765 1821 905
rect 1867 765 1932 905
rect 1792 647 1932 765
rect 2032 813 2136 939
rect 2032 673 2061 813
rect 2107 673 2136 813
rect 2032 647 2136 673
rect 2236 905 2340 939
rect 2236 765 2265 905
rect 2311 765 2340 905
rect 2236 647 2340 765
rect 2440 861 2544 939
rect 2440 721 2469 861
rect 2515 721 2544 861
rect 2440 647 2544 721
rect 2644 905 2748 939
rect 2644 765 2673 905
rect 2719 765 2748 905
rect 2644 647 2748 765
rect 2848 858 2952 939
rect 2848 718 2877 858
rect 2923 718 2952 858
rect 2848 647 2952 718
rect 3052 905 3156 939
rect 3052 765 3081 905
rect 3127 765 3156 905
rect 3052 647 3156 765
rect 3256 861 3360 939
rect 3256 721 3285 861
rect 3331 721 3360 861
rect 3256 647 3360 721
rect 3460 905 3548 939
rect 3460 765 3489 905
rect 3535 765 3548 905
rect 3460 647 3548 765
rect 1792 573 1872 647
<< mvndiffc >>
rect 49 147 95 287
rect 273 239 319 285
rect 497 147 543 193
rect 721 228 767 274
rect 945 147 991 193
rect 1169 239 1215 285
rect 1393 147 1439 193
rect 1617 239 1663 285
rect 1841 147 1887 287
rect 2265 102 2311 242
rect 2673 147 2719 287
rect 3081 147 3127 287
rect 3489 147 3535 287
<< mvpdiffc >>
rect 69 765 115 905
rect 497 721 543 861
rect 935 765 981 905
rect 1383 721 1429 861
rect 1821 765 1867 905
rect 2061 673 2107 813
rect 2265 765 2311 905
rect 2469 721 2515 861
rect 2673 765 2719 905
rect 2877 718 2923 858
rect 3081 765 3127 905
rect 3285 721 3331 861
rect 3489 765 3535 905
<< polysilicon >>
rect 144 939 244 983
rect 368 939 468 983
rect 582 939 682 983
rect 806 939 906 983
rect 1030 939 1130 983
rect 1254 939 1354 983
rect 1478 939 1578 983
rect 1692 939 1792 983
rect 1932 939 2032 983
rect 2136 939 2236 983
rect 2340 939 2440 983
rect 2544 939 2644 983
rect 2748 939 2848 983
rect 2952 939 3052 983
rect 3156 939 3256 983
rect 3360 939 3460 983
rect 144 524 244 573
rect 144 478 185 524
rect 231 478 244 524
rect 144 377 244 478
rect 368 513 468 573
rect 582 524 682 573
rect 582 513 623 524
rect 368 478 623 513
rect 669 478 682 524
rect 368 441 682 478
rect 368 377 468 441
rect 124 333 244 377
rect 348 333 468 377
rect 572 377 682 441
rect 806 524 906 573
rect 806 478 819 524
rect 865 513 906 524
rect 1030 513 1130 573
rect 865 478 1130 513
rect 806 441 1130 478
rect 806 377 916 441
rect 572 333 692 377
rect 796 333 916 377
rect 1020 377 1130 441
rect 1254 524 1354 573
rect 1254 478 1267 524
rect 1313 513 1354 524
rect 1478 513 1578 573
rect 1313 478 1578 513
rect 1254 441 1578 478
rect 1254 377 1364 441
rect 1020 333 1140 377
rect 1244 333 1364 377
rect 1468 377 1578 441
rect 1692 524 1792 573
rect 1692 478 1705 524
rect 1751 478 1792 524
rect 1692 377 1792 478
rect 1932 524 2032 647
rect 1932 478 1945 524
rect 1991 478 2032 524
rect 1932 377 2032 478
rect 2136 513 2236 647
rect 2340 524 2440 647
rect 2340 513 2381 524
rect 2136 478 2381 513
rect 2427 478 2440 524
rect 2136 441 2440 478
rect 2136 377 2236 441
rect 1468 333 1588 377
rect 1692 333 1812 377
rect 1922 333 2042 377
rect 2116 333 2236 377
rect 2340 377 2440 441
rect 2544 524 2644 647
rect 2544 478 2575 524
rect 2621 513 2644 524
rect 2748 513 2848 647
rect 2952 537 3052 647
rect 2621 478 2848 513
rect 2544 441 2848 478
rect 2544 377 2644 441
rect 2340 333 2460 377
rect 2524 333 2644 377
rect 2748 377 2848 441
rect 2932 524 3052 537
rect 2932 478 2945 524
rect 2991 513 3052 524
rect 3156 513 3256 647
rect 2991 478 3256 513
rect 2932 441 3256 478
rect 2748 333 2868 377
rect 2932 333 3052 441
rect 3156 377 3256 441
rect 3360 524 3460 647
rect 3360 478 3373 524
rect 3419 478 3460 524
rect 3360 377 3460 478
rect 3156 333 3276 377
rect 3340 333 3460 377
rect 124 25 244 69
rect 348 25 468 69
rect 572 25 692 69
rect 796 25 916 69
rect 1020 25 1140 69
rect 1244 25 1364 69
rect 1468 25 1588 69
rect 1692 25 1812 69
rect 1922 25 2042 69
rect 2116 25 2236 69
rect 2340 25 2460 69
rect 2524 25 2644 69
rect 2748 25 2868 69
rect 2932 25 3052 69
rect 3156 25 3276 69
rect 3340 25 3460 69
<< polycontact >>
rect 185 478 231 524
rect 623 478 669 524
rect 819 478 865 524
rect 1267 478 1313 524
rect 1705 478 1751 524
rect 1945 478 1991 524
rect 2381 478 2427 524
rect 2575 478 2621 524
rect 2945 478 2991 524
rect 3373 478 3419 524
<< metal1 >>
rect 0 918 3584 1098
rect 69 905 115 918
rect 935 905 981 918
rect 69 754 115 765
rect 497 861 543 872
rect 1821 905 1867 918
rect 935 754 981 765
rect 1383 861 1429 872
rect 497 708 543 721
rect 2265 905 2311 918
rect 1821 754 1867 765
rect 2061 813 2107 824
rect 1383 708 1429 721
rect 82 673 2061 708
rect 2673 905 2719 918
rect 2469 861 2515 872
rect 2265 754 2311 765
rect 2382 721 2469 766
rect 3081 905 3127 918
rect 2673 754 2719 765
rect 2877 858 2923 869
rect 2382 708 2515 721
rect 3489 905 3535 918
rect 3081 754 3127 765
rect 3285 861 3331 872
rect 2877 708 2923 718
rect 3489 754 3535 765
rect 3285 708 3331 721
rect 2107 673 3331 708
rect 82 662 3331 673
rect 82 390 128 662
rect 174 570 1416 616
rect 174 524 242 570
rect 814 524 866 570
rect 1370 524 1416 570
rect 1934 570 3094 616
rect 1934 524 1991 570
rect 2575 524 2621 570
rect 3048 524 3094 570
rect 174 478 185 524
rect 231 478 242 524
rect 612 478 623 524
rect 669 478 754 524
rect 702 420 754 478
rect 814 478 819 524
rect 865 478 866 524
rect 814 466 866 478
rect 912 478 1267 524
rect 1313 478 1324 524
rect 1370 478 1705 524
rect 1751 478 1762 524
rect 1934 478 1945 524
rect 2370 478 2381 524
rect 2427 478 2500 524
rect 912 420 958 478
rect 1934 466 1991 478
rect 82 344 656 390
rect 702 374 958 420
rect 2454 431 2500 478
rect 2575 467 2621 478
rect 2667 478 2945 524
rect 2991 478 3002 524
rect 3048 478 3373 524
rect 3419 478 3430 524
rect 2454 400 2546 431
rect 2667 400 2713 478
rect 702 354 754 374
rect 49 287 95 298
rect 273 285 319 344
rect 273 228 319 239
rect 610 308 656 344
rect 1196 320 1663 366
rect 2466 354 2713 400
rect 1196 316 1242 320
rect 798 308 1242 316
rect 610 285 1242 308
rect 610 274 1169 285
rect 610 228 721 274
rect 767 270 1169 274
rect 767 228 824 270
rect 1215 239 1242 285
rect 1169 228 1242 239
rect 1617 285 1663 320
rect 1617 228 1663 239
rect 1841 308 2420 345
rect 2759 344 3535 390
rect 2759 308 2805 344
rect 1841 299 2805 308
rect 1841 287 1887 299
rect 486 182 497 193
rect 95 147 497 182
rect 543 182 554 193
rect 934 182 945 193
rect 543 147 945 182
rect 991 182 1002 193
rect 1382 182 1393 193
rect 991 147 1393 182
rect 1439 182 1450 193
rect 1439 147 1841 182
rect 2374 287 2805 299
rect 2374 262 2673 287
rect 49 136 1887 147
rect 2265 242 2311 253
rect 2719 262 2805 287
rect 3081 287 3127 298
rect 2673 136 2719 147
rect 2265 90 2311 102
rect 3081 90 3127 147
rect 3489 287 3535 344
rect 3489 136 3535 147
rect 0 -90 3584 90
<< labels >>
flabel metal1 s 912 478 1324 524 0 FreeSans 200 0 0 0 A1
port 1 nsew default input
flabel metal1 s 174 570 1416 616 0 FreeSans 200 0 0 0 A2
port 2 nsew default input
flabel metal1 s 1934 570 3094 616 0 FreeSans 200 0 0 0 B
port 3 nsew default input
flabel metal1 s 2667 478 3002 524 0 FreeSans 200 0 0 0 C
port 4 nsew default input
flabel metal1 s 0 918 3584 1098 0 FreeSans 200 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 3081 253 3127 298 0 FreeSans 200 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel metal1 s 3285 869 3331 872 0 FreeSans 200 0 0 0 ZN
port 5 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 7 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 8 nsew ground bidirectional
rlabel metal1 s 612 478 754 524 1 A1
port 1 nsew default input
rlabel metal1 s 912 420 958 478 1 A1
port 1 nsew default input
rlabel metal1 s 702 420 754 478 1 A1
port 1 nsew default input
rlabel metal1 s 702 374 958 420 1 A1
port 1 nsew default input
rlabel metal1 s 702 354 754 374 1 A1
port 1 nsew default input
rlabel metal1 s 1370 524 1416 570 1 A2
port 2 nsew default input
rlabel metal1 s 814 524 866 570 1 A2
port 2 nsew default input
rlabel metal1 s 174 524 242 570 1 A2
port 2 nsew default input
rlabel metal1 s 1370 478 1762 524 1 A2
port 2 nsew default input
rlabel metal1 s 814 478 866 524 1 A2
port 2 nsew default input
rlabel metal1 s 174 478 242 524 1 A2
port 2 nsew default input
rlabel metal1 s 814 466 866 478 1 A2
port 2 nsew default input
rlabel metal1 s 3048 524 3094 570 1 B
port 3 nsew default input
rlabel metal1 s 2575 524 2621 570 1 B
port 3 nsew default input
rlabel metal1 s 1934 524 1991 570 1 B
port 3 nsew default input
rlabel metal1 s 3048 478 3430 524 1 B
port 3 nsew default input
rlabel metal1 s 2575 478 2621 524 1 B
port 3 nsew default input
rlabel metal1 s 1934 478 1991 524 1 B
port 3 nsew default input
rlabel metal1 s 2575 467 2621 478 1 B
port 3 nsew default input
rlabel metal1 s 1934 467 1991 478 1 B
port 3 nsew default input
rlabel metal1 s 1934 466 1991 467 1 B
port 3 nsew default input
rlabel metal1 s 2370 478 2500 524 1 C
port 4 nsew default input
rlabel metal1 s 2667 431 2713 478 1 C
port 4 nsew default input
rlabel metal1 s 2454 431 2500 478 1 C
port 4 nsew default input
rlabel metal1 s 2667 400 2713 431 1 C
port 4 nsew default input
rlabel metal1 s 2454 400 2546 431 1 C
port 4 nsew default input
rlabel metal1 s 2466 354 2713 400 1 C
port 4 nsew default input
rlabel metal1 s 2469 869 2515 872 1 ZN
port 5 nsew default output
rlabel metal1 s 1383 869 1429 872 1 ZN
port 5 nsew default output
rlabel metal1 s 497 869 543 872 1 ZN
port 5 nsew default output
rlabel metal1 s 3285 824 3331 869 1 ZN
port 5 nsew default output
rlabel metal1 s 2877 824 2923 869 1 ZN
port 5 nsew default output
rlabel metal1 s 2469 824 2515 869 1 ZN
port 5 nsew default output
rlabel metal1 s 1383 824 1429 869 1 ZN
port 5 nsew default output
rlabel metal1 s 497 824 543 869 1 ZN
port 5 nsew default output
rlabel metal1 s 3285 766 3331 824 1 ZN
port 5 nsew default output
rlabel metal1 s 2877 766 2923 824 1 ZN
port 5 nsew default output
rlabel metal1 s 2469 766 2515 824 1 ZN
port 5 nsew default output
rlabel metal1 s 2061 766 2107 824 1 ZN
port 5 nsew default output
rlabel metal1 s 1383 766 1429 824 1 ZN
port 5 nsew default output
rlabel metal1 s 497 766 543 824 1 ZN
port 5 nsew default output
rlabel metal1 s 3285 708 3331 766 1 ZN
port 5 nsew default output
rlabel metal1 s 2877 708 2923 766 1 ZN
port 5 nsew default output
rlabel metal1 s 2382 708 2515 766 1 ZN
port 5 nsew default output
rlabel metal1 s 2061 708 2107 766 1 ZN
port 5 nsew default output
rlabel metal1 s 1383 708 1429 766 1 ZN
port 5 nsew default output
rlabel metal1 s 497 708 543 766 1 ZN
port 5 nsew default output
rlabel metal1 s 82 662 3331 708 1 ZN
port 5 nsew default output
rlabel metal1 s 82 390 128 662 1 ZN
port 5 nsew default output
rlabel metal1 s 82 366 656 390 1 ZN
port 5 nsew default output
rlabel metal1 s 1196 344 1663 366 1 ZN
port 5 nsew default output
rlabel metal1 s 82 344 656 366 1 ZN
port 5 nsew default output
rlabel metal1 s 1196 320 1663 344 1 ZN
port 5 nsew default output
rlabel metal1 s 610 320 656 344 1 ZN
port 5 nsew default output
rlabel metal1 s 273 320 319 344 1 ZN
port 5 nsew default output
rlabel metal1 s 1617 316 1663 320 1 ZN
port 5 nsew default output
rlabel metal1 s 1196 316 1242 320 1 ZN
port 5 nsew default output
rlabel metal1 s 610 316 656 320 1 ZN
port 5 nsew default output
rlabel metal1 s 273 316 319 320 1 ZN
port 5 nsew default output
rlabel metal1 s 1617 308 1663 316 1 ZN
port 5 nsew default output
rlabel metal1 s 798 308 1242 316 1 ZN
port 5 nsew default output
rlabel metal1 s 610 308 656 316 1 ZN
port 5 nsew default output
rlabel metal1 s 273 308 319 316 1 ZN
port 5 nsew default output
rlabel metal1 s 1617 270 1663 308 1 ZN
port 5 nsew default output
rlabel metal1 s 610 270 1242 308 1 ZN
port 5 nsew default output
rlabel metal1 s 273 270 319 308 1 ZN
port 5 nsew default output
rlabel metal1 s 1617 228 1663 270 1 ZN
port 5 nsew default output
rlabel metal1 s 1169 228 1242 270 1 ZN
port 5 nsew default output
rlabel metal1 s 610 228 824 270 1 ZN
port 5 nsew default output
rlabel metal1 s 273 228 319 270 1 ZN
port 5 nsew default output
rlabel metal1 s 3489 754 3535 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3081 754 3127 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2673 754 2719 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2265 754 2311 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1821 754 1867 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 935 754 981 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 69 754 115 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3081 90 3127 253 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2265 90 2311 253 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 3584 90 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3584 1008
string GDS_END 220710
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 212630
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
