magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 453 2774 1094
<< pwell >>
rect -86 -86 2774 453
<< mvnmos >>
rect 168 68 288 332
rect 336 68 456 332
rect 560 68 680 332
rect 728 68 848 332
rect 952 68 1072 332
rect 1120 68 1240 332
rect 1344 68 1464 332
rect 1512 68 1632 332
rect 1772 148 1892 332
rect 1996 148 2116 332
rect 2220 148 2340 332
rect 2444 148 2564 332
<< mvpmos >>
rect 164 574 264 940
rect 368 574 468 940
rect 572 574 672 940
rect 776 574 876 940
rect 980 574 1080 940
rect 1184 574 1284 940
rect 1388 574 1488 940
rect 1592 574 1692 940
rect 1852 574 1952 940
rect 2056 574 2156 940
rect 2260 574 2360 940
rect 2464 574 2564 940
<< mvndiff >>
rect 80 127 168 332
rect 80 81 93 127
rect 139 81 168 127
rect 80 68 168 81
rect 288 68 336 332
rect 456 219 560 332
rect 456 173 485 219
rect 531 173 560 219
rect 456 68 560 173
rect 680 68 728 332
rect 848 127 952 332
rect 848 81 877 127
rect 923 81 952 127
rect 848 68 952 81
rect 1072 68 1120 332
rect 1240 233 1344 332
rect 1240 187 1269 233
rect 1315 187 1344 233
rect 1240 68 1344 187
rect 1464 68 1512 332
rect 1632 206 1772 332
rect 1632 160 1661 206
rect 1707 160 1772 206
rect 1632 148 1772 160
rect 1892 319 1996 332
rect 1892 179 1921 319
rect 1967 179 1996 319
rect 1892 148 1996 179
rect 2116 301 2220 332
rect 2116 161 2145 301
rect 2191 161 2220 301
rect 2116 148 2220 161
rect 2340 319 2444 332
rect 2340 179 2369 319
rect 2415 179 2444 319
rect 2340 148 2444 179
rect 2564 301 2652 332
rect 2564 161 2593 301
rect 2639 161 2652 301
rect 2564 148 2652 161
rect 1632 68 1712 148
<< mvpdiff >>
rect 76 858 164 940
rect 76 718 89 858
rect 135 718 164 858
rect 76 574 164 718
rect 264 755 368 940
rect 264 615 293 755
rect 339 615 368 755
rect 264 574 368 615
rect 468 858 572 940
rect 468 718 497 858
rect 543 718 572 858
rect 468 574 572 718
rect 672 756 776 940
rect 672 616 701 756
rect 747 616 776 756
rect 672 574 776 616
rect 876 858 980 940
rect 876 718 905 858
rect 951 718 980 858
rect 876 574 980 718
rect 1080 766 1184 940
rect 1080 626 1109 766
rect 1155 626 1184 766
rect 1080 574 1184 626
rect 1284 858 1388 940
rect 1284 718 1313 858
rect 1359 718 1388 858
rect 1284 574 1388 718
rect 1488 766 1592 940
rect 1488 626 1517 766
rect 1563 626 1592 766
rect 1488 574 1592 626
rect 1692 835 1852 940
rect 1692 695 1721 835
rect 1767 695 1852 835
rect 1692 574 1852 695
rect 1952 927 2056 940
rect 1952 787 1981 927
rect 2027 787 2056 927
rect 1952 574 2056 787
rect 2156 835 2260 940
rect 2156 695 2185 835
rect 2231 695 2260 835
rect 2156 574 2260 695
rect 2360 927 2464 940
rect 2360 787 2389 927
rect 2435 787 2464 927
rect 2360 574 2464 787
rect 2564 835 2652 940
rect 2564 695 2593 835
rect 2639 695 2652 835
rect 2564 574 2652 695
<< mvndiffc >>
rect 93 81 139 127
rect 485 173 531 219
rect 877 81 923 127
rect 1269 187 1315 233
rect 1661 160 1707 206
rect 1921 179 1967 319
rect 2145 161 2191 301
rect 2369 179 2415 319
rect 2593 161 2639 301
<< mvpdiffc >>
rect 89 718 135 858
rect 293 615 339 755
rect 497 718 543 858
rect 701 616 747 756
rect 905 718 951 858
rect 1109 626 1155 766
rect 1313 718 1359 858
rect 1517 626 1563 766
rect 1721 695 1767 835
rect 1981 787 2027 927
rect 2185 695 2231 835
rect 2389 787 2435 927
rect 2593 695 2639 835
<< polysilicon >>
rect 164 940 264 984
rect 368 940 468 984
rect 572 940 672 984
rect 776 940 876 984
rect 980 940 1080 984
rect 1184 940 1284 984
rect 1388 940 1488 984
rect 1592 940 1692 984
rect 1852 940 1952 984
rect 2056 940 2156 984
rect 2260 940 2360 984
rect 2464 940 2564 984
rect 164 530 264 574
rect 168 479 264 530
rect 368 541 468 574
rect 368 495 381 541
rect 427 514 468 541
rect 572 514 672 574
rect 427 495 672 514
rect 168 466 299 479
rect 168 420 240 466
rect 286 420 299 466
rect 168 407 299 420
rect 368 442 672 495
rect 168 332 288 407
rect 368 376 456 442
rect 336 332 456 376
rect 560 376 672 442
rect 776 464 876 574
rect 980 530 1080 574
rect 980 464 1072 530
rect 1184 464 1284 574
rect 1388 530 1488 574
rect 1592 541 1692 574
rect 1388 464 1464 530
rect 776 449 1072 464
rect 776 403 789 449
rect 835 403 1072 449
rect 776 392 1072 403
rect 776 376 848 392
rect 560 332 680 376
rect 728 332 848 376
rect 952 332 1072 392
rect 1120 411 1464 464
rect 1120 365 1133 411
rect 1179 392 1464 411
rect 1179 365 1240 392
rect 1120 332 1240 365
rect 1344 332 1464 392
rect 1592 495 1605 541
rect 1651 495 1692 541
rect 1592 482 1692 495
rect 1592 376 1632 482
rect 1852 464 1952 574
rect 2056 539 2156 574
rect 2056 493 2084 539
rect 2130 493 2156 539
rect 2056 464 2156 493
rect 2260 540 2360 574
rect 2260 494 2288 540
rect 2334 494 2360 540
rect 2260 464 2360 494
rect 2464 487 2564 574
rect 2464 464 2494 487
rect 1512 332 1632 376
rect 1772 441 2494 464
rect 2540 441 2564 487
rect 1772 392 2564 441
rect 1772 332 1892 392
rect 1996 332 2116 392
rect 2220 332 2340 392
rect 2444 332 2564 392
rect 1772 104 1892 148
rect 1996 104 2116 148
rect 2220 104 2340 148
rect 2444 104 2564 148
rect 168 24 288 68
rect 336 24 456 68
rect 560 24 680 68
rect 728 24 848 68
rect 952 24 1072 68
rect 1120 24 1240 68
rect 1344 24 1464 68
rect 1512 24 1632 68
<< polycontact >>
rect 381 495 427 541
rect 240 420 286 466
rect 789 403 835 449
rect 1133 365 1179 411
rect 1605 495 1651 541
rect 2084 493 2130 539
rect 2288 494 2334 540
rect 2494 441 2540 487
<< metal1 >>
rect 0 927 2688 1098
rect 0 918 1981 927
rect 89 858 1776 869
rect 135 823 497 858
rect 89 707 135 718
rect 282 755 339 767
rect 282 615 293 755
rect 543 823 905 858
rect 497 707 543 718
rect 701 756 747 767
rect 339 616 701 661
rect 951 823 1313 858
rect 905 707 951 718
rect 1109 766 1155 777
rect 747 626 1109 661
rect 1359 835 1776 858
rect 1359 823 1721 835
rect 1313 707 1359 718
rect 1517 766 1563 777
rect 1155 626 1517 661
rect 1710 695 1721 823
rect 1767 741 1776 835
rect 1970 787 1981 918
rect 2027 918 2389 927
rect 2027 787 2038 918
rect 2174 835 2242 846
rect 2174 741 2185 835
rect 1767 695 2185 741
rect 2231 741 2242 835
rect 2378 787 2389 918
rect 2435 918 2688 927
rect 2435 787 2446 918
rect 2582 835 2650 846
rect 2582 741 2593 835
rect 2231 695 2593 741
rect 2639 695 2650 835
rect 1563 626 1766 649
rect 747 616 1766 626
rect 339 615 1766 616
rect 1516 603 1766 615
rect 142 541 427 569
rect 142 523 381 541
rect 142 314 194 523
rect 381 484 427 495
rect 686 541 1662 542
rect 686 495 1605 541
rect 1651 495 1662 541
rect 240 466 286 477
rect 686 449 873 495
rect 686 438 789 449
rect 286 420 789 438
rect 240 403 789 420
rect 835 403 873 449
rect 240 392 873 403
rect 1133 411 1179 422
rect 1710 404 1766 603
rect 1926 540 2547 550
rect 1926 539 2288 540
rect 1926 493 2084 539
rect 2130 494 2288 539
rect 2334 494 2547 540
rect 2130 493 2547 494
rect 1926 487 2547 493
rect 1926 466 2494 487
rect 2540 466 2547 487
rect 2540 441 2546 466
rect 2494 430 2546 441
rect 1710 400 2415 404
rect 1133 314 1179 365
rect 142 265 1179 314
rect 1269 358 2415 400
rect 1269 354 1967 358
rect 1269 233 1315 354
rect 474 173 485 219
rect 531 187 1269 219
rect 1921 319 1967 354
rect 531 173 1315 187
rect 1661 206 1707 217
rect 2369 319 2415 358
rect 1921 168 1967 179
rect 2145 301 2191 312
rect 93 127 139 138
rect 0 81 93 90
rect 866 90 877 127
rect 139 81 877 90
rect 923 90 934 127
rect 1661 90 1707 160
rect 2369 168 2415 179
rect 2593 301 2639 312
rect 2145 90 2191 161
rect 2593 90 2639 161
rect 923 81 2688 90
rect 0 -90 2688 81
<< labels >>
flabel metal1 s 142 523 427 569 0 FreeSans 200 0 0 0 A1
port 1 nsew default input
flabel metal1 s 686 495 1662 542 0 FreeSans 200 0 0 0 A2
port 2 nsew default input
flabel metal1 s 1926 466 2547 550 0 FreeSans 200 0 0 0 B
port 3 nsew default input
flabel metal1 s 0 918 2688 1098 0 FreeSans 200 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 2593 217 2639 312 0 FreeSans 200 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel metal1 s 1517 767 1563 777 0 FreeSans 200 0 0 0 ZN
port 4 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 6 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 381 484 427 523 1 A1
port 1 nsew default input
rlabel metal1 s 142 484 194 523 1 A1
port 1 nsew default input
rlabel metal1 s 142 422 194 484 1 A1
port 1 nsew default input
rlabel metal1 s 1133 314 1179 422 1 A1
port 1 nsew default input
rlabel metal1 s 142 314 194 422 1 A1
port 1 nsew default input
rlabel metal1 s 142 265 1179 314 1 A1
port 1 nsew default input
rlabel metal1 s 686 477 873 495 1 A2
port 2 nsew default input
rlabel metal1 s 686 438 873 477 1 A2
port 2 nsew default input
rlabel metal1 s 240 438 286 477 1 A2
port 2 nsew default input
rlabel metal1 s 240 392 873 438 1 A2
port 2 nsew default input
rlabel metal1 s 2494 430 2546 466 1 B
port 3 nsew default input
rlabel metal1 s 1109 767 1155 777 1 ZN
port 4 nsew default output
rlabel metal1 s 1517 661 1563 767 1 ZN
port 4 nsew default output
rlabel metal1 s 1109 661 1155 767 1 ZN
port 4 nsew default output
rlabel metal1 s 701 661 747 767 1 ZN
port 4 nsew default output
rlabel metal1 s 282 661 339 767 1 ZN
port 4 nsew default output
rlabel metal1 s 282 649 1563 661 1 ZN
port 4 nsew default output
rlabel metal1 s 282 615 1766 649 1 ZN
port 4 nsew default output
rlabel metal1 s 1516 603 1766 615 1 ZN
port 4 nsew default output
rlabel metal1 s 1710 404 1766 603 1 ZN
port 4 nsew default output
rlabel metal1 s 1710 400 2415 404 1 ZN
port 4 nsew default output
rlabel metal1 s 1269 358 2415 400 1 ZN
port 4 nsew default output
rlabel metal1 s 2369 354 2415 358 1 ZN
port 4 nsew default output
rlabel metal1 s 1269 354 1967 358 1 ZN
port 4 nsew default output
rlabel metal1 s 2369 219 2415 354 1 ZN
port 4 nsew default output
rlabel metal1 s 1921 219 1967 354 1 ZN
port 4 nsew default output
rlabel metal1 s 1269 219 1315 354 1 ZN
port 4 nsew default output
rlabel metal1 s 2369 173 2415 219 1 ZN
port 4 nsew default output
rlabel metal1 s 1921 173 1967 219 1 ZN
port 4 nsew default output
rlabel metal1 s 474 173 1315 219 1 ZN
port 4 nsew default output
rlabel metal1 s 2369 168 2415 173 1 ZN
port 4 nsew default output
rlabel metal1 s 1921 168 1967 173 1 ZN
port 4 nsew default output
rlabel metal1 s 2378 787 2446 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1970 787 2038 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2145 217 2191 312 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2593 138 2639 217 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2145 138 2191 217 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1661 138 1707 217 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2593 127 2639 138 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2145 127 2191 138 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1661 127 1707 138 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 93 127 139 138 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2593 90 2639 127 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2145 90 2191 127 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1661 90 1707 127 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 866 90 934 127 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 93 90 139 127 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 2688 90 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2688 1008
string GDS_END 1181428
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1174770
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
