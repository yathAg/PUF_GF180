magic
tech gf180mcuD
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 352 5686 870
<< pwell >>
rect -86 -86 5686 352
<< mvnmos >>
rect 124 68 244 232
rect 348 68 468 232
rect 572 68 692 232
rect 796 68 916 232
rect 1020 68 1140 232
rect 1244 68 1364 232
rect 1468 68 1588 232
rect 1692 68 1812 232
rect 1916 68 2036 232
rect 2140 68 2260 232
rect 2364 68 2484 232
rect 2588 68 2708 232
rect 2812 68 2932 232
rect 3036 68 3156 232
rect 3260 68 3380 232
rect 3484 68 3604 232
rect 3708 68 3828 232
rect 3932 68 4052 232
rect 4156 68 4276 232
rect 4380 68 4500 232
rect 4604 68 4724 232
rect 4828 68 4948 232
rect 5052 68 5172 232
rect 5276 68 5396 232
<< mvpmos >>
rect 124 472 224 716
rect 348 472 448 716
rect 572 472 672 716
rect 796 472 896 716
rect 1020 472 1120 716
rect 1244 472 1344 716
rect 1468 472 1568 716
rect 1692 472 1792 716
rect 1916 472 2016 716
rect 2140 472 2240 716
rect 2364 472 2464 716
rect 2588 472 2688 716
rect 2812 472 2912 716
rect 3036 472 3136 716
rect 3260 472 3360 716
rect 3484 472 3584 716
rect 3708 472 3808 716
rect 3932 472 4032 716
rect 4156 472 4256 716
rect 4380 472 4480 716
rect 4604 472 4704 716
rect 4828 472 4928 716
rect 5052 472 5152 716
rect 5276 472 5376 716
<< mvndiff >>
rect 36 142 124 232
rect 36 96 49 142
rect 95 96 124 142
rect 36 68 124 96
rect 244 192 348 232
rect 244 146 273 192
rect 319 146 348 192
rect 244 68 348 146
rect 468 142 572 232
rect 468 96 497 142
rect 543 96 572 142
rect 468 68 572 96
rect 692 192 796 232
rect 692 146 721 192
rect 767 146 796 192
rect 692 68 796 146
rect 916 142 1020 232
rect 916 96 945 142
rect 991 96 1020 142
rect 916 68 1020 96
rect 1140 192 1244 232
rect 1140 146 1169 192
rect 1215 146 1244 192
rect 1140 68 1244 146
rect 1364 142 1468 232
rect 1364 96 1393 142
rect 1439 96 1468 142
rect 1364 68 1468 96
rect 1588 192 1692 232
rect 1588 146 1617 192
rect 1663 146 1692 192
rect 1588 68 1692 146
rect 1812 142 1916 232
rect 1812 96 1841 142
rect 1887 96 1916 142
rect 1812 68 1916 96
rect 2036 192 2140 232
rect 2036 146 2065 192
rect 2111 146 2140 192
rect 2036 68 2140 146
rect 2260 140 2364 232
rect 2260 94 2289 140
rect 2335 94 2364 140
rect 2260 68 2364 94
rect 2484 192 2588 232
rect 2484 146 2513 192
rect 2559 146 2588 192
rect 2484 68 2588 146
rect 2708 140 2812 232
rect 2708 94 2737 140
rect 2783 94 2812 140
rect 2708 68 2812 94
rect 2932 192 3036 232
rect 2932 146 2961 192
rect 3007 146 3036 192
rect 2932 68 3036 146
rect 3156 140 3260 232
rect 3156 94 3185 140
rect 3231 94 3260 140
rect 3156 68 3260 94
rect 3380 192 3484 232
rect 3380 146 3409 192
rect 3455 146 3484 192
rect 3380 68 3484 146
rect 3604 140 3708 232
rect 3604 94 3633 140
rect 3679 94 3708 140
rect 3604 68 3708 94
rect 3828 192 3932 232
rect 3828 146 3857 192
rect 3903 146 3932 192
rect 3828 68 3932 146
rect 4052 140 4156 232
rect 4052 94 4081 140
rect 4127 94 4156 140
rect 4052 68 4156 94
rect 4276 192 4380 232
rect 4276 146 4305 192
rect 4351 146 4380 192
rect 4276 68 4380 146
rect 4500 140 4604 232
rect 4500 94 4529 140
rect 4575 94 4604 140
rect 4500 68 4604 94
rect 4724 192 4828 232
rect 4724 146 4753 192
rect 4799 146 4828 192
rect 4724 68 4828 146
rect 4948 140 5052 232
rect 4948 94 4977 140
rect 5023 94 5052 140
rect 4948 68 5052 94
rect 5172 192 5276 232
rect 5172 146 5201 192
rect 5247 146 5276 192
rect 5172 68 5276 146
rect 5396 142 5484 232
rect 5396 96 5425 142
rect 5471 96 5484 142
rect 5396 68 5484 96
<< mvpdiff >>
rect 36 665 124 716
rect 36 525 49 665
rect 95 525 124 665
rect 36 472 124 525
rect 224 665 348 716
rect 224 525 253 665
rect 299 525 348 665
rect 224 472 348 525
rect 448 665 572 716
rect 448 619 477 665
rect 523 619 572 665
rect 448 472 572 619
rect 672 665 796 716
rect 672 525 701 665
rect 747 525 796 665
rect 672 472 796 525
rect 896 665 1020 716
rect 896 619 925 665
rect 971 619 1020 665
rect 896 472 1020 619
rect 1120 665 1244 716
rect 1120 525 1149 665
rect 1195 525 1244 665
rect 1120 472 1244 525
rect 1344 665 1468 716
rect 1344 619 1373 665
rect 1419 619 1468 665
rect 1344 472 1468 619
rect 1568 665 1692 716
rect 1568 525 1597 665
rect 1643 525 1692 665
rect 1568 472 1692 525
rect 1792 665 1916 716
rect 1792 525 1821 665
rect 1867 525 1916 665
rect 1792 472 1916 525
rect 2016 665 2140 716
rect 2016 525 2065 665
rect 2111 525 2140 665
rect 2016 472 2140 525
rect 2240 665 2364 716
rect 2240 619 2269 665
rect 2315 619 2364 665
rect 2240 472 2364 619
rect 2464 665 2588 716
rect 2464 525 2493 665
rect 2539 525 2588 665
rect 2464 472 2588 525
rect 2688 665 2812 716
rect 2688 619 2717 665
rect 2763 619 2812 665
rect 2688 472 2812 619
rect 2912 665 3036 716
rect 2912 525 2941 665
rect 2987 525 3036 665
rect 2912 472 3036 525
rect 3136 665 3260 716
rect 3136 619 3165 665
rect 3211 619 3260 665
rect 3136 472 3260 619
rect 3360 665 3484 716
rect 3360 525 3389 665
rect 3435 525 3484 665
rect 3360 472 3484 525
rect 3584 665 3708 716
rect 3584 619 3613 665
rect 3659 619 3708 665
rect 3584 472 3708 619
rect 3808 665 3932 716
rect 3808 525 3837 665
rect 3883 525 3932 665
rect 3808 472 3932 525
rect 4032 665 4156 716
rect 4032 619 4061 665
rect 4107 619 4156 665
rect 4032 472 4156 619
rect 4256 665 4380 716
rect 4256 525 4285 665
rect 4331 525 4380 665
rect 4256 472 4380 525
rect 4480 665 4604 716
rect 4480 619 4509 665
rect 4555 619 4604 665
rect 4480 472 4604 619
rect 4704 665 4828 716
rect 4704 525 4733 665
rect 4779 525 4828 665
rect 4704 472 4828 525
rect 4928 665 5052 716
rect 4928 619 4957 665
rect 5003 619 5052 665
rect 4928 472 5052 619
rect 5152 665 5276 716
rect 5152 525 5181 665
rect 5227 525 5276 665
rect 5152 472 5276 525
rect 5376 665 5464 716
rect 5376 525 5405 665
rect 5451 525 5464 665
rect 5376 472 5464 525
<< mvndiffc >>
rect 49 96 95 142
rect 273 146 319 192
rect 497 96 543 142
rect 721 146 767 192
rect 945 96 991 142
rect 1169 146 1215 192
rect 1393 96 1439 142
rect 1617 146 1663 192
rect 1841 96 1887 142
rect 2065 146 2111 192
rect 2289 94 2335 140
rect 2513 146 2559 192
rect 2737 94 2783 140
rect 2961 146 3007 192
rect 3185 94 3231 140
rect 3409 146 3455 192
rect 3633 94 3679 140
rect 3857 146 3903 192
rect 4081 94 4127 140
rect 4305 146 4351 192
rect 4529 94 4575 140
rect 4753 146 4799 192
rect 4977 94 5023 140
rect 5201 146 5247 192
rect 5425 96 5471 142
<< mvpdiffc >>
rect 49 525 95 665
rect 253 525 299 665
rect 477 619 523 665
rect 701 525 747 665
rect 925 619 971 665
rect 1149 525 1195 665
rect 1373 619 1419 665
rect 1597 525 1643 665
rect 1821 525 1867 665
rect 2065 525 2111 665
rect 2269 619 2315 665
rect 2493 525 2539 665
rect 2717 619 2763 665
rect 2941 525 2987 665
rect 3165 619 3211 665
rect 3389 525 3435 665
rect 3613 619 3659 665
rect 3837 525 3883 665
rect 4061 619 4107 665
rect 4285 525 4331 665
rect 4509 619 4555 665
rect 4733 525 4779 665
rect 4957 619 5003 665
rect 5181 525 5227 665
rect 5405 525 5451 665
<< polysilicon >>
rect 124 716 224 760
rect 348 716 448 760
rect 572 716 672 760
rect 796 716 896 760
rect 1020 716 1120 760
rect 1244 716 1344 760
rect 1468 716 1568 760
rect 1692 716 1792 760
rect 1916 716 2016 760
rect 2140 716 2240 760
rect 2364 716 2464 760
rect 2588 716 2688 760
rect 2812 716 2912 760
rect 3036 716 3136 760
rect 3260 716 3360 760
rect 3484 716 3584 760
rect 3708 716 3808 760
rect 3932 716 4032 760
rect 4156 716 4256 760
rect 4380 716 4480 760
rect 4604 716 4704 760
rect 4828 716 4928 760
rect 5052 716 5152 760
rect 5276 716 5376 760
rect 124 402 224 472
rect 348 402 448 472
rect 572 402 672 472
rect 796 402 896 472
rect 1020 402 1120 472
rect 1244 402 1344 472
rect 1468 402 1568 472
rect 1692 402 1792 472
rect 1916 407 2016 472
rect 2140 407 2240 472
rect 2364 407 2464 472
rect 2588 407 2688 472
rect 2812 407 2912 472
rect 3036 407 3136 472
rect 3260 407 3360 472
rect 3484 407 3584 472
rect 3708 407 3808 472
rect 3932 407 4032 472
rect 4156 407 4256 472
rect 4380 407 4480 472
rect 4604 407 4704 472
rect 4828 407 4928 472
rect 5052 407 5152 472
rect 5276 407 5376 472
rect 124 389 1812 402
rect 124 343 159 389
rect 1615 343 1812 389
rect 124 330 1812 343
rect 124 232 244 330
rect 348 232 468 330
rect 572 232 692 330
rect 796 232 916 330
rect 1020 232 1140 330
rect 1244 232 1364 330
rect 1468 300 1812 330
rect 1468 232 1588 300
rect 1692 232 1812 300
rect 1916 394 5396 407
rect 1916 348 1929 394
rect 3291 348 3923 394
rect 5379 348 5396 394
rect 1916 335 5396 348
rect 1916 232 2036 335
rect 2140 232 2260 335
rect 2364 232 2484 335
rect 2588 232 2708 335
rect 2812 232 2932 335
rect 3036 232 3156 335
rect 3260 232 3380 335
rect 3484 232 3604 335
rect 3708 232 3828 335
rect 3932 232 4052 335
rect 4156 232 4276 335
rect 4380 232 4500 335
rect 4604 232 4724 335
rect 4828 232 4948 335
rect 5052 232 5172 335
rect 5276 232 5396 335
rect 124 24 244 68
rect 348 24 468 68
rect 572 24 692 68
rect 796 24 916 68
rect 1020 24 1140 68
rect 1244 24 1364 68
rect 1468 24 1588 68
rect 1692 24 1812 68
rect 1916 24 2036 68
rect 2140 24 2260 68
rect 2364 24 2484 68
rect 2588 24 2708 68
rect 2812 24 2932 68
rect 3036 24 3156 68
rect 3260 24 3380 68
rect 3484 24 3604 68
rect 3708 24 3828 68
rect 3932 24 4052 68
rect 4156 24 4276 68
rect 4380 24 4500 68
rect 4604 24 4724 68
rect 4828 24 4948 68
rect 5052 24 5172 68
rect 5276 24 5396 68
<< polycontact >>
rect 159 343 1615 389
rect 1929 348 3291 394
rect 3923 348 5379 394
<< metal1 >>
rect 0 724 5600 844
rect 49 665 95 724
rect 49 506 95 525
rect 253 665 299 676
rect 477 665 523 724
rect 477 600 523 619
rect 701 665 747 676
rect 299 525 701 552
rect 925 665 971 724
rect 925 600 971 619
rect 1149 665 1195 676
rect 747 525 1149 552
rect 1373 665 1419 724
rect 1373 600 1419 619
rect 1597 665 1643 676
rect 1195 525 1597 552
rect 1821 665 1867 724
rect 1643 525 1754 552
rect 253 506 1754 525
rect 1821 506 1867 525
rect 2065 665 2111 676
rect 2269 665 2315 724
rect 2269 608 2315 619
rect 2493 665 2539 676
rect 2111 525 2493 562
rect 2717 665 2763 724
rect 2717 608 2763 619
rect 2941 665 2987 676
rect 2539 525 2941 562
rect 3165 665 3211 724
rect 3165 608 3211 619
rect 3389 665 3435 676
rect 2987 525 3389 562
rect 3613 665 3659 724
rect 3613 608 3659 619
rect 3837 665 3883 676
rect 3435 525 3837 562
rect 4061 665 4107 724
rect 4061 608 4107 619
rect 4285 665 4331 676
rect 3883 525 4285 562
rect 4509 665 4555 724
rect 4509 608 4555 619
rect 4733 665 4779 676
rect 4331 525 4733 562
rect 4957 665 5003 724
rect 4957 608 5003 619
rect 5181 665 5227 676
rect 4779 525 5181 562
rect 124 389 1637 430
rect 124 343 159 389
rect 1615 343 1637 389
rect 124 342 1637 343
rect 1707 394 1754 506
rect 2065 446 5227 525
rect 5405 665 5451 724
rect 5405 506 5451 525
rect 1707 348 1929 394
rect 3291 348 3302 394
rect 1707 250 1754 348
rect 3550 302 3730 446
rect 3912 348 3923 394
rect 5379 348 5396 394
rect 273 203 1754 250
rect 273 192 319 203
rect 38 142 106 153
rect 38 96 49 142
rect 95 96 106 142
rect 721 192 767 203
rect 273 135 319 146
rect 486 142 554 153
rect 38 60 106 96
rect 486 96 497 142
rect 543 96 554 142
rect 1169 192 1215 203
rect 721 135 767 146
rect 934 142 1002 153
rect 486 60 554 96
rect 934 96 945 142
rect 991 96 1002 142
rect 1617 192 1663 203
rect 1169 135 1215 146
rect 1382 142 1450 153
rect 934 60 1002 96
rect 1382 96 1393 142
rect 1439 96 1450 142
rect 2065 192 5247 302
rect 1617 135 1663 146
rect 1830 142 1898 153
rect 1382 60 1450 96
rect 1830 96 1841 142
rect 1887 96 1898 142
rect 2111 186 2513 192
rect 2111 146 2117 186
rect 2065 135 2117 146
rect 2559 186 2961 192
rect 1830 60 1898 96
rect 2278 94 2289 140
rect 2335 94 2346 140
rect 2513 135 2559 146
rect 3007 186 3409 192
rect 2278 60 2346 94
rect 2726 94 2737 140
rect 2783 94 2794 140
rect 2961 135 3007 146
rect 3455 186 3857 192
rect 2726 60 2794 94
rect 3174 94 3185 140
rect 3231 94 3242 140
rect 3409 135 3455 146
rect 3903 186 4305 192
rect 3174 60 3242 94
rect 3622 94 3633 140
rect 3679 94 3690 140
rect 3857 135 3903 146
rect 4351 186 4753 192
rect 3622 60 3690 94
rect 4070 94 4081 140
rect 4127 94 4138 140
rect 4305 135 4351 146
rect 4799 186 5201 192
rect 4070 60 4138 94
rect 4518 94 4529 140
rect 4575 94 4586 140
rect 4753 135 4799 146
rect 4518 60 4586 94
rect 4966 94 4977 140
rect 5023 94 5034 140
rect 5201 135 5247 146
rect 5414 142 5482 153
rect 4966 60 5034 94
rect 5414 96 5425 142
rect 5471 96 5482 142
rect 5414 60 5482 96
rect 0 -60 5600 60
<< labels >>
flabel metal1 s 5181 562 5227 676 0 FreeSans 600 0 0 0 Z
port 2 nsew default output
flabel metal1 s 124 342 1637 430 0 FreeSans 600 0 0 0 I
port 1 nsew default input
flabel metal1 s 0 724 5600 844 0 FreeSans 400 0 0 0 VDD
port 3 nsew power bidirectional abutment
flabel metal1 s 5414 140 5482 153 0 FreeSans 400 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 4 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 4733 562 4779 676 1 Z
port 2 nsew default output
rlabel metal1 s 4285 562 4331 676 1 Z
port 2 nsew default output
rlabel metal1 s 3837 562 3883 676 1 Z
port 2 nsew default output
rlabel metal1 s 3389 562 3435 676 1 Z
port 2 nsew default output
rlabel metal1 s 2941 562 2987 676 1 Z
port 2 nsew default output
rlabel metal1 s 2493 562 2539 676 1 Z
port 2 nsew default output
rlabel metal1 s 2065 562 2111 676 1 Z
port 2 nsew default output
rlabel metal1 s 2065 446 5227 562 1 Z
port 2 nsew default output
rlabel metal1 s 3550 302 3730 446 1 Z
port 2 nsew default output
rlabel metal1 s 2065 186 5247 302 1 Z
port 2 nsew default output
rlabel metal1 s 5201 135 5247 186 1 Z
port 2 nsew default output
rlabel metal1 s 4753 135 4799 186 1 Z
port 2 nsew default output
rlabel metal1 s 4305 135 4351 186 1 Z
port 2 nsew default output
rlabel metal1 s 3857 135 3903 186 1 Z
port 2 nsew default output
rlabel metal1 s 3409 135 3455 186 1 Z
port 2 nsew default output
rlabel metal1 s 2961 135 3007 186 1 Z
port 2 nsew default output
rlabel metal1 s 2513 135 2559 186 1 Z
port 2 nsew default output
rlabel metal1 s 2065 135 2117 186 1 Z
port 2 nsew default output
rlabel metal1 s 5405 608 5451 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4957 608 5003 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4509 608 4555 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4061 608 4107 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3613 608 3659 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3165 608 3211 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2717 608 2763 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2269 608 2315 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1821 608 1867 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1373 608 1419 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 925 608 971 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 477 608 523 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 608 95 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 5405 600 5451 608 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1821 600 1867 608 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1373 600 1419 608 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 925 600 971 608 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 477 600 523 608 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 600 95 608 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 5405 506 5451 600 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1821 506 1867 600 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 506 95 600 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1830 140 1898 153 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1382 140 1450 153 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 934 140 1002 153 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 486 140 554 153 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 38 140 106 153 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 5414 60 5482 140 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 4966 60 5034 140 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 4518 60 4586 140 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 4070 60 4138 140 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3622 60 3690 140 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3174 60 3242 140 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2726 60 2794 140 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2278 60 2346 140 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1830 60 1898 140 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1382 60 1450 140 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 934 60 1002 140 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 486 60 554 140 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 38 60 106 140 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 5600 60 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 5600 784
string GDS_END 1372732
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1360696
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
