magic
tech gf180mcuA
magscale 1 10
timestamp 1698431365
<< nwell >>
rect 3728 2553 5177 2591
rect 2156 2431 3010 2432
rect 3726 2431 5177 2553
rect 2155 2302 5177 2431
rect -532 1217 5177 2302
rect -532 1196 4580 1217
rect -176 1137 4580 1196
rect -176 1096 1540 1137
rect 1813 1115 2349 1137
<< mvnmos >>
rect 2635 2569 2755 2761
rect 3030 2553 3150 2673
rect 79 533 199 957
rect 303 533 423 957
rect 527 533 647 957
rect 751 533 871 957
rect 975 533 1095 957
rect 1199 533 1319 957
rect 1629 544 1749 864
rect 2021 540 2141 980
rect 2491 544 2611 998
rect 2715 544 2835 998
rect 2939 544 3059 998
rect 3409 807 3529 999
rect 3981 389 4101 957
rect 4205 389 4325 957
rect 4429 389 4549 957
rect 4653 389 4773 957
<< mvpmos >>
rect 79 1238 199 1994
rect 303 1238 423 1994
rect 527 1238 647 1994
rect 751 1238 871 1994
rect 975 1238 1095 1994
rect 1199 1238 1319 1994
rect 1629 1279 1749 2079
rect 2021 1235 2141 2135
rect 2411 2062 2531 2290
rect 2635 2062 2755 2290
rect 3017 2050 3137 2290
rect 2491 1279 2611 1733
rect 2715 1279 2835 1733
rect 2939 1279 3059 1733
rect 3409 1406 3529 1860
rect 3936 1337 4056 2471
rect 4160 1337 4280 2471
rect 4384 1337 4504 2471
rect 4608 1337 4728 2471
<< mvndiff >>
rect 2547 2748 2635 2761
rect 2547 2702 2560 2748
rect 2606 2702 2635 2748
rect 2547 2628 2635 2702
rect 2547 2582 2560 2628
rect 2606 2582 2635 2628
rect 2547 2569 2635 2582
rect 2755 2748 2843 2761
rect 2755 2702 2784 2748
rect 2830 2702 2843 2748
rect 2755 2628 2843 2702
rect 2755 2582 2784 2628
rect 2830 2582 2843 2628
rect 2755 2569 2843 2582
rect 2942 2636 3030 2673
rect 2942 2590 2955 2636
rect 3001 2590 3030 2636
rect 2942 2553 3030 2590
rect 3150 2636 3238 2673
rect 3150 2590 3179 2636
rect 3225 2590 3238 2636
rect 3150 2553 3238 2590
rect -9 944 79 957
rect -9 898 4 944
rect 50 898 79 944
rect -9 826 79 898
rect -9 780 4 826
rect 50 780 79 826
rect -9 709 79 780
rect -9 663 4 709
rect 50 663 79 709
rect -9 592 79 663
rect -9 546 4 592
rect 50 546 79 592
rect -9 533 79 546
rect 199 944 303 957
rect 199 898 228 944
rect 274 898 303 944
rect 199 826 303 898
rect 199 780 228 826
rect 274 780 303 826
rect 199 709 303 780
rect 199 663 228 709
rect 274 663 303 709
rect 199 592 303 663
rect 199 546 228 592
rect 274 546 303 592
rect 199 533 303 546
rect 423 944 527 957
rect 423 898 452 944
rect 498 898 527 944
rect 423 826 527 898
rect 423 780 452 826
rect 498 780 527 826
rect 423 709 527 780
rect 423 663 452 709
rect 498 663 527 709
rect 423 592 527 663
rect 423 546 452 592
rect 498 546 527 592
rect 423 533 527 546
rect 647 944 751 957
rect 647 898 676 944
rect 722 898 751 944
rect 647 826 751 898
rect 647 780 676 826
rect 722 780 751 826
rect 647 709 751 780
rect 647 663 676 709
rect 722 663 751 709
rect 647 592 751 663
rect 647 546 676 592
rect 722 546 751 592
rect 647 533 751 546
rect 871 944 975 957
rect 871 898 900 944
rect 946 898 975 944
rect 871 826 975 898
rect 871 780 900 826
rect 946 780 975 826
rect 871 709 975 780
rect 871 663 900 709
rect 946 663 975 709
rect 871 592 975 663
rect 871 546 900 592
rect 946 546 975 592
rect 871 533 975 546
rect 1095 944 1199 957
rect 1095 898 1124 944
rect 1170 898 1199 944
rect 1095 826 1199 898
rect 1095 780 1124 826
rect 1170 780 1199 826
rect 1095 709 1199 780
rect 1095 663 1124 709
rect 1170 663 1199 709
rect 1095 592 1199 663
rect 1095 546 1124 592
rect 1170 546 1199 592
rect 1095 533 1199 546
rect 1319 944 1407 957
rect 1319 898 1348 944
rect 1394 898 1407 944
rect 1319 826 1407 898
rect 2403 985 2491 998
rect 1933 967 2021 980
rect 1933 921 1946 967
rect 1992 921 2021 967
rect 1319 780 1348 826
rect 1394 780 1407 826
rect 1319 709 1407 780
rect 1319 663 1348 709
rect 1394 663 1407 709
rect 1319 592 1407 663
rect 1319 546 1348 592
rect 1394 546 1407 592
rect 1319 533 1407 546
rect 1541 851 1629 864
rect 1541 805 1554 851
rect 1600 805 1629 851
rect 1541 727 1629 805
rect 1541 681 1554 727
rect 1600 681 1629 727
rect 1541 603 1629 681
rect 1541 557 1554 603
rect 1600 557 1629 603
rect 1541 544 1629 557
rect 1749 851 1837 864
rect 1749 805 1778 851
rect 1824 805 1837 851
rect 1749 727 1837 805
rect 1749 681 1778 727
rect 1824 681 1837 727
rect 1749 603 1837 681
rect 1749 557 1778 603
rect 1824 557 1837 603
rect 1749 544 1837 557
rect 1933 845 2021 921
rect 1933 799 1946 845
rect 1992 799 2021 845
rect 1933 722 2021 799
rect 1933 676 1946 722
rect 1992 676 2021 722
rect 1933 599 2021 676
rect 1933 553 1946 599
rect 1992 553 2021 599
rect 1933 540 2021 553
rect 2141 967 2229 980
rect 2141 921 2170 967
rect 2216 921 2229 967
rect 2141 845 2229 921
rect 2141 799 2170 845
rect 2216 799 2229 845
rect 2141 722 2229 799
rect 2141 676 2170 722
rect 2216 676 2229 722
rect 2141 599 2229 676
rect 2141 553 2170 599
rect 2216 553 2229 599
rect 2141 540 2229 553
rect 2403 939 2416 985
rect 2462 939 2491 985
rect 2403 858 2491 939
rect 2403 812 2416 858
rect 2462 812 2491 858
rect 2403 731 2491 812
rect 2403 685 2416 731
rect 2462 685 2491 731
rect 2403 603 2491 685
rect 2403 557 2416 603
rect 2462 557 2491 603
rect 2403 544 2491 557
rect 2611 985 2715 998
rect 2611 939 2640 985
rect 2686 939 2715 985
rect 2611 858 2715 939
rect 2611 812 2640 858
rect 2686 812 2715 858
rect 2611 731 2715 812
rect 2611 685 2640 731
rect 2686 685 2715 731
rect 2611 603 2715 685
rect 2611 557 2640 603
rect 2686 557 2715 603
rect 2611 544 2715 557
rect 2835 985 2939 998
rect 2835 939 2864 985
rect 2910 939 2939 985
rect 2835 858 2939 939
rect 2835 812 2864 858
rect 2910 812 2939 858
rect 2835 731 2939 812
rect 2835 685 2864 731
rect 2910 685 2939 731
rect 2835 603 2939 685
rect 2835 557 2864 603
rect 2910 557 2939 603
rect 2835 544 2939 557
rect 3059 985 3147 998
rect 3059 939 3088 985
rect 3134 939 3147 985
rect 3059 858 3147 939
rect 3059 812 3088 858
rect 3134 812 3147 858
rect 3059 731 3147 812
rect 3321 986 3409 999
rect 3321 940 3334 986
rect 3380 940 3409 986
rect 3321 866 3409 940
rect 3321 820 3334 866
rect 3380 820 3409 866
rect 3321 807 3409 820
rect 3529 986 3617 999
rect 3529 940 3558 986
rect 3604 940 3617 986
rect 3529 866 3617 940
rect 3529 820 3558 866
rect 3604 820 3617 866
rect 3529 807 3617 820
rect 3893 944 3981 957
rect 3893 898 3906 944
rect 3952 898 3981 944
rect 3893 820 3981 898
rect 3059 685 3088 731
rect 3134 685 3147 731
rect 3059 603 3147 685
rect 3059 557 3088 603
rect 3134 557 3147 603
rect 3059 544 3147 557
rect 3893 774 3906 820
rect 3952 774 3981 820
rect 3893 696 3981 774
rect 3893 650 3906 696
rect 3952 650 3981 696
rect 3893 572 3981 650
rect 3893 526 3906 572
rect 3952 526 3981 572
rect 3893 448 3981 526
rect 3893 402 3906 448
rect 3952 402 3981 448
rect 3893 389 3981 402
rect 4101 944 4205 957
rect 4101 898 4130 944
rect 4176 898 4205 944
rect 4101 820 4205 898
rect 4101 774 4130 820
rect 4176 774 4205 820
rect 4101 696 4205 774
rect 4101 650 4130 696
rect 4176 650 4205 696
rect 4101 572 4205 650
rect 4101 526 4130 572
rect 4176 526 4205 572
rect 4101 448 4205 526
rect 4101 402 4130 448
rect 4176 402 4205 448
rect 4101 389 4205 402
rect 4325 944 4429 957
rect 4325 898 4354 944
rect 4400 898 4429 944
rect 4325 820 4429 898
rect 4325 774 4354 820
rect 4400 774 4429 820
rect 4325 696 4429 774
rect 4325 650 4354 696
rect 4400 650 4429 696
rect 4325 572 4429 650
rect 4325 526 4354 572
rect 4400 526 4429 572
rect 4325 448 4429 526
rect 4325 402 4354 448
rect 4400 402 4429 448
rect 4325 389 4429 402
rect 4549 944 4653 957
rect 4549 898 4578 944
rect 4624 898 4653 944
rect 4549 820 4653 898
rect 4549 774 4578 820
rect 4624 774 4653 820
rect 4549 696 4653 774
rect 4549 650 4578 696
rect 4624 650 4653 696
rect 4549 572 4653 650
rect 4549 526 4578 572
rect 4624 526 4653 572
rect 4549 448 4653 526
rect 4549 402 4578 448
rect 4624 402 4653 448
rect 4549 389 4653 402
rect 4773 944 4861 957
rect 4773 898 4802 944
rect 4848 898 4861 944
rect 4773 820 4861 898
rect 4773 774 4802 820
rect 4848 774 4861 820
rect 4773 696 4861 774
rect 4773 650 4802 696
rect 4848 650 4861 696
rect 4773 572 4861 650
rect 4773 526 4802 572
rect 4848 526 4861 572
rect 4773 448 4861 526
rect 4773 402 4802 448
rect 4848 402 4861 448
rect 4773 389 4861 402
<< mvpdiff >>
rect 3848 2458 3936 2471
rect 3848 2412 3861 2458
rect 3907 2412 3936 2458
rect 3848 2352 3936 2412
rect 3848 2306 3861 2352
rect 3907 2306 3936 2352
rect 2323 2277 2411 2290
rect 2323 2231 2336 2277
rect 2382 2231 2411 2277
rect 1933 2122 2021 2135
rect 1541 2066 1629 2079
rect 1541 2020 1554 2066
rect 1600 2020 1629 2066
rect -9 1981 79 1994
rect -9 1935 4 1981
rect 50 1935 79 1981
rect -9 1867 79 1935
rect -9 1821 4 1867
rect 50 1821 79 1867
rect -9 1753 79 1821
rect -9 1707 4 1753
rect 50 1707 79 1753
rect -9 1639 79 1707
rect -9 1593 4 1639
rect 50 1593 79 1639
rect -9 1525 79 1593
rect -9 1479 4 1525
rect 50 1479 79 1525
rect -9 1411 79 1479
rect -9 1365 4 1411
rect 50 1365 79 1411
rect -9 1297 79 1365
rect -9 1251 4 1297
rect 50 1251 79 1297
rect -9 1238 79 1251
rect 199 1981 303 1994
rect 199 1935 228 1981
rect 274 1935 303 1981
rect 199 1867 303 1935
rect 199 1821 228 1867
rect 274 1821 303 1867
rect 199 1753 303 1821
rect 199 1707 228 1753
rect 274 1707 303 1753
rect 199 1639 303 1707
rect 199 1593 228 1639
rect 274 1593 303 1639
rect 199 1525 303 1593
rect 199 1479 228 1525
rect 274 1479 303 1525
rect 199 1411 303 1479
rect 199 1365 228 1411
rect 274 1365 303 1411
rect 199 1297 303 1365
rect 199 1251 228 1297
rect 274 1251 303 1297
rect 199 1238 303 1251
rect 423 1981 527 1994
rect 423 1935 452 1981
rect 498 1935 527 1981
rect 423 1867 527 1935
rect 423 1821 452 1867
rect 498 1821 527 1867
rect 423 1753 527 1821
rect 423 1707 452 1753
rect 498 1707 527 1753
rect 423 1639 527 1707
rect 423 1593 452 1639
rect 498 1593 527 1639
rect 423 1525 527 1593
rect 423 1479 452 1525
rect 498 1479 527 1525
rect 423 1411 527 1479
rect 423 1365 452 1411
rect 498 1365 527 1411
rect 423 1297 527 1365
rect 423 1251 452 1297
rect 498 1251 527 1297
rect 423 1238 527 1251
rect 647 1981 751 1994
rect 647 1935 676 1981
rect 722 1935 751 1981
rect 647 1867 751 1935
rect 647 1821 676 1867
rect 722 1821 751 1867
rect 647 1753 751 1821
rect 647 1707 676 1753
rect 722 1707 751 1753
rect 647 1639 751 1707
rect 647 1593 676 1639
rect 722 1593 751 1639
rect 647 1525 751 1593
rect 647 1479 676 1525
rect 722 1479 751 1525
rect 647 1411 751 1479
rect 647 1365 676 1411
rect 722 1365 751 1411
rect 647 1297 751 1365
rect 647 1251 676 1297
rect 722 1251 751 1297
rect 647 1238 751 1251
rect 871 1981 975 1994
rect 871 1935 900 1981
rect 946 1935 975 1981
rect 871 1867 975 1935
rect 871 1821 900 1867
rect 946 1821 975 1867
rect 871 1753 975 1821
rect 871 1707 900 1753
rect 946 1707 975 1753
rect 871 1639 975 1707
rect 871 1593 900 1639
rect 946 1593 975 1639
rect 871 1525 975 1593
rect 871 1479 900 1525
rect 946 1479 975 1525
rect 871 1411 975 1479
rect 871 1365 900 1411
rect 946 1365 975 1411
rect 871 1297 975 1365
rect 871 1251 900 1297
rect 946 1251 975 1297
rect 871 1238 975 1251
rect 1095 1981 1199 1994
rect 1095 1935 1124 1981
rect 1170 1935 1199 1981
rect 1095 1867 1199 1935
rect 1095 1821 1124 1867
rect 1170 1821 1199 1867
rect 1095 1753 1199 1821
rect 1095 1707 1124 1753
rect 1170 1707 1199 1753
rect 1095 1639 1199 1707
rect 1095 1593 1124 1639
rect 1170 1593 1199 1639
rect 1095 1525 1199 1593
rect 1095 1479 1124 1525
rect 1170 1479 1199 1525
rect 1095 1411 1199 1479
rect 1095 1365 1124 1411
rect 1170 1365 1199 1411
rect 1095 1297 1199 1365
rect 1095 1251 1124 1297
rect 1170 1251 1199 1297
rect 1095 1238 1199 1251
rect 1319 1981 1407 1994
rect 1319 1935 1348 1981
rect 1394 1935 1407 1981
rect 1319 1867 1407 1935
rect 1319 1821 1348 1867
rect 1394 1821 1407 1867
rect 1319 1753 1407 1821
rect 1319 1707 1348 1753
rect 1394 1707 1407 1753
rect 1319 1639 1407 1707
rect 1319 1593 1348 1639
rect 1394 1593 1407 1639
rect 1319 1525 1407 1593
rect 1319 1479 1348 1525
rect 1394 1479 1407 1525
rect 1319 1411 1407 1479
rect 1319 1365 1348 1411
rect 1394 1365 1407 1411
rect 1319 1297 1407 1365
rect 1319 1251 1348 1297
rect 1394 1251 1407 1297
rect 1541 1962 1629 2020
rect 1541 1916 1554 1962
rect 1600 1916 1629 1962
rect 1541 1858 1629 1916
rect 1541 1812 1554 1858
rect 1600 1812 1629 1858
rect 1541 1754 1629 1812
rect 1541 1708 1554 1754
rect 1600 1708 1629 1754
rect 1541 1650 1629 1708
rect 1541 1604 1554 1650
rect 1600 1604 1629 1650
rect 1541 1546 1629 1604
rect 1541 1500 1554 1546
rect 1600 1500 1629 1546
rect 1541 1442 1629 1500
rect 1541 1396 1554 1442
rect 1600 1396 1629 1442
rect 1541 1338 1629 1396
rect 1541 1292 1554 1338
rect 1600 1292 1629 1338
rect 1541 1279 1629 1292
rect 1749 2066 1837 2079
rect 1749 2020 1778 2066
rect 1824 2020 1837 2066
rect 1749 1962 1837 2020
rect 1749 1916 1778 1962
rect 1824 1916 1837 1962
rect 1749 1858 1837 1916
rect 1749 1812 1778 1858
rect 1824 1812 1837 1858
rect 1749 1754 1837 1812
rect 1749 1708 1778 1754
rect 1824 1708 1837 1754
rect 1749 1650 1837 1708
rect 1749 1604 1778 1650
rect 1824 1604 1837 1650
rect 1749 1546 1837 1604
rect 1749 1500 1778 1546
rect 1824 1500 1837 1546
rect 1749 1442 1837 1500
rect 1749 1396 1778 1442
rect 1824 1396 1837 1442
rect 1749 1338 1837 1396
rect 1749 1292 1778 1338
rect 1824 1292 1837 1338
rect 1749 1279 1837 1292
rect 1933 2076 1946 2122
rect 1992 2076 2021 2122
rect 1933 2019 2021 2076
rect 1933 1973 1946 2019
rect 1992 1973 2021 2019
rect 1933 1916 2021 1973
rect 1933 1870 1946 1916
rect 1992 1870 2021 1916
rect 1933 1813 2021 1870
rect 1933 1767 1946 1813
rect 1992 1767 2021 1813
rect 1933 1710 2021 1767
rect 1933 1664 1946 1710
rect 1992 1664 2021 1710
rect 1933 1606 2021 1664
rect 1933 1560 1946 1606
rect 1992 1560 2021 1606
rect 1933 1502 2021 1560
rect 1933 1456 1946 1502
rect 1992 1456 2021 1502
rect 1933 1398 2021 1456
rect 1933 1352 1946 1398
rect 1992 1352 2021 1398
rect 1933 1294 2021 1352
rect 1319 1238 1407 1251
rect 1933 1248 1946 1294
rect 1992 1248 2021 1294
rect 1933 1235 2021 1248
rect 2141 2122 2229 2135
rect 2141 2076 2170 2122
rect 2216 2076 2229 2122
rect 2141 2019 2229 2076
rect 2323 2121 2411 2231
rect 2323 2075 2336 2121
rect 2382 2075 2411 2121
rect 2323 2062 2411 2075
rect 2531 2277 2635 2290
rect 2531 2231 2560 2277
rect 2606 2231 2635 2277
rect 2531 2121 2635 2231
rect 2531 2075 2560 2121
rect 2606 2075 2635 2121
rect 2531 2062 2635 2075
rect 2755 2277 3017 2290
rect 2755 2231 2784 2277
rect 2830 2231 2942 2277
rect 2988 2231 3017 2277
rect 2755 2121 3017 2231
rect 2755 2075 2784 2121
rect 2830 2109 3017 2121
rect 2830 2075 2942 2109
rect 2755 2063 2942 2075
rect 2988 2063 3017 2109
rect 2755 2062 3017 2063
rect 2141 1973 2170 2019
rect 2216 1973 2229 2019
rect 2929 2050 3017 2062
rect 3137 2277 3225 2290
rect 3137 2231 3166 2277
rect 3212 2231 3225 2277
rect 3137 2109 3225 2231
rect 3137 2063 3166 2109
rect 3212 2063 3225 2109
rect 3137 2050 3225 2063
rect 3848 2246 3936 2306
rect 3848 2200 3861 2246
rect 3907 2200 3936 2246
rect 3848 2140 3936 2200
rect 3848 2094 3861 2140
rect 3907 2094 3936 2140
rect 3848 2034 3936 2094
rect 2141 1916 2229 1973
rect 2141 1870 2170 1916
rect 2216 1870 2229 1916
rect 2141 1813 2229 1870
rect 2141 1767 2170 1813
rect 2216 1767 2229 1813
rect 2141 1710 2229 1767
rect 3848 1988 3861 2034
rect 3907 1988 3936 2034
rect 3848 1928 3936 1988
rect 3848 1882 3861 1928
rect 3907 1882 3936 1928
rect 3321 1847 3409 1860
rect 3321 1801 3334 1847
rect 3380 1801 3409 1847
rect 2141 1664 2170 1710
rect 2216 1664 2229 1710
rect 2141 1606 2229 1664
rect 2141 1560 2170 1606
rect 2216 1560 2229 1606
rect 2141 1502 2229 1560
rect 2141 1456 2170 1502
rect 2216 1456 2229 1502
rect 2141 1398 2229 1456
rect 2141 1352 2170 1398
rect 2216 1352 2229 1398
rect 2141 1294 2229 1352
rect 2141 1248 2170 1294
rect 2216 1248 2229 1294
rect 2403 1720 2491 1733
rect 2403 1674 2416 1720
rect 2462 1674 2491 1720
rect 2403 1593 2491 1674
rect 2403 1547 2416 1593
rect 2462 1547 2491 1593
rect 2403 1466 2491 1547
rect 2403 1420 2416 1466
rect 2462 1420 2491 1466
rect 2403 1338 2491 1420
rect 2403 1292 2416 1338
rect 2462 1292 2491 1338
rect 2403 1279 2491 1292
rect 2611 1720 2715 1733
rect 2611 1674 2640 1720
rect 2686 1674 2715 1720
rect 2611 1593 2715 1674
rect 2611 1547 2640 1593
rect 2686 1547 2715 1593
rect 2611 1466 2715 1547
rect 2611 1420 2640 1466
rect 2686 1420 2715 1466
rect 2611 1338 2715 1420
rect 2611 1292 2640 1338
rect 2686 1292 2715 1338
rect 2611 1279 2715 1292
rect 2835 1720 2939 1733
rect 2835 1674 2864 1720
rect 2910 1674 2939 1720
rect 2835 1593 2939 1674
rect 2835 1547 2864 1593
rect 2910 1547 2939 1593
rect 2835 1466 2939 1547
rect 2835 1420 2864 1466
rect 2910 1420 2939 1466
rect 2835 1338 2939 1420
rect 2835 1292 2864 1338
rect 2910 1292 2939 1338
rect 2835 1279 2939 1292
rect 3059 1720 3147 1733
rect 3059 1674 3088 1720
rect 3134 1674 3147 1720
rect 3059 1593 3147 1674
rect 3059 1547 3088 1593
rect 3134 1547 3147 1593
rect 3059 1466 3147 1547
rect 3059 1420 3088 1466
rect 3134 1420 3147 1466
rect 3059 1338 3147 1420
rect 3321 1720 3409 1801
rect 3321 1674 3334 1720
rect 3380 1674 3409 1720
rect 3321 1593 3409 1674
rect 3321 1547 3334 1593
rect 3380 1547 3409 1593
rect 3321 1465 3409 1547
rect 3321 1419 3334 1465
rect 3380 1419 3409 1465
rect 3321 1406 3409 1419
rect 3529 1847 3617 1860
rect 3529 1801 3558 1847
rect 3604 1801 3617 1847
rect 3529 1720 3617 1801
rect 3529 1674 3558 1720
rect 3604 1674 3617 1720
rect 3529 1593 3617 1674
rect 3529 1547 3558 1593
rect 3604 1547 3617 1593
rect 3529 1465 3617 1547
rect 3529 1419 3558 1465
rect 3604 1419 3617 1465
rect 3529 1406 3617 1419
rect 3848 1822 3936 1882
rect 3848 1776 3861 1822
rect 3907 1776 3936 1822
rect 3848 1716 3936 1776
rect 3848 1670 3861 1716
rect 3907 1670 3936 1716
rect 3848 1610 3936 1670
rect 3848 1564 3861 1610
rect 3907 1564 3936 1610
rect 3848 1503 3936 1564
rect 3848 1457 3861 1503
rect 3907 1457 3936 1503
rect 3059 1292 3088 1338
rect 3134 1292 3147 1338
rect 3059 1279 3147 1292
rect 2141 1235 2229 1248
rect 3848 1396 3936 1457
rect 3848 1350 3861 1396
rect 3907 1350 3936 1396
rect 3848 1337 3936 1350
rect 4056 2458 4160 2471
rect 4056 2412 4085 2458
rect 4131 2412 4160 2458
rect 4056 2352 4160 2412
rect 4056 2306 4085 2352
rect 4131 2306 4160 2352
rect 4056 2246 4160 2306
rect 4056 2200 4085 2246
rect 4131 2200 4160 2246
rect 4056 2140 4160 2200
rect 4056 2094 4085 2140
rect 4131 2094 4160 2140
rect 4056 2034 4160 2094
rect 4056 1988 4085 2034
rect 4131 1988 4160 2034
rect 4056 1928 4160 1988
rect 4056 1882 4085 1928
rect 4131 1882 4160 1928
rect 4056 1822 4160 1882
rect 4056 1776 4085 1822
rect 4131 1776 4160 1822
rect 4056 1716 4160 1776
rect 4056 1670 4085 1716
rect 4131 1670 4160 1716
rect 4056 1610 4160 1670
rect 4056 1564 4085 1610
rect 4131 1564 4160 1610
rect 4056 1503 4160 1564
rect 4056 1457 4085 1503
rect 4131 1457 4160 1503
rect 4056 1396 4160 1457
rect 4056 1350 4085 1396
rect 4131 1350 4160 1396
rect 4056 1337 4160 1350
rect 4280 2458 4384 2471
rect 4280 2412 4309 2458
rect 4355 2412 4384 2458
rect 4280 2352 4384 2412
rect 4280 2306 4309 2352
rect 4355 2306 4384 2352
rect 4280 2246 4384 2306
rect 4280 2200 4309 2246
rect 4355 2200 4384 2246
rect 4280 2140 4384 2200
rect 4280 2094 4309 2140
rect 4355 2094 4384 2140
rect 4280 2034 4384 2094
rect 4280 1988 4309 2034
rect 4355 1988 4384 2034
rect 4280 1928 4384 1988
rect 4280 1882 4309 1928
rect 4355 1882 4384 1928
rect 4280 1822 4384 1882
rect 4280 1776 4309 1822
rect 4355 1776 4384 1822
rect 4280 1716 4384 1776
rect 4280 1670 4309 1716
rect 4355 1670 4384 1716
rect 4280 1610 4384 1670
rect 4280 1564 4309 1610
rect 4355 1564 4384 1610
rect 4280 1503 4384 1564
rect 4280 1457 4309 1503
rect 4355 1457 4384 1503
rect 4280 1396 4384 1457
rect 4280 1350 4309 1396
rect 4355 1350 4384 1396
rect 4280 1337 4384 1350
rect 4504 2458 4608 2471
rect 4504 2412 4533 2458
rect 4579 2412 4608 2458
rect 4504 2352 4608 2412
rect 4504 2306 4533 2352
rect 4579 2306 4608 2352
rect 4504 2246 4608 2306
rect 4504 2200 4533 2246
rect 4579 2200 4608 2246
rect 4504 2140 4608 2200
rect 4504 2094 4533 2140
rect 4579 2094 4608 2140
rect 4504 2034 4608 2094
rect 4504 1988 4533 2034
rect 4579 1988 4608 2034
rect 4504 1928 4608 1988
rect 4504 1882 4533 1928
rect 4579 1882 4608 1928
rect 4504 1822 4608 1882
rect 4504 1776 4533 1822
rect 4579 1776 4608 1822
rect 4504 1716 4608 1776
rect 4504 1670 4533 1716
rect 4579 1670 4608 1716
rect 4504 1610 4608 1670
rect 4504 1564 4533 1610
rect 4579 1564 4608 1610
rect 4504 1503 4608 1564
rect 4504 1457 4533 1503
rect 4579 1457 4608 1503
rect 4504 1396 4608 1457
rect 4504 1350 4533 1396
rect 4579 1350 4608 1396
rect 4504 1337 4608 1350
rect 4728 2458 4816 2471
rect 4728 2412 4757 2458
rect 4803 2412 4816 2458
rect 4728 2352 4816 2412
rect 4728 2306 4757 2352
rect 4803 2306 4816 2352
rect 4728 2246 4816 2306
rect 4728 2200 4757 2246
rect 4803 2200 4816 2246
rect 4728 2140 4816 2200
rect 4728 2094 4757 2140
rect 4803 2094 4816 2140
rect 4728 2034 4816 2094
rect 4728 1988 4757 2034
rect 4803 1988 4816 2034
rect 4728 1928 4816 1988
rect 4728 1882 4757 1928
rect 4803 1882 4816 1928
rect 4728 1822 4816 1882
rect 4728 1776 4757 1822
rect 4803 1776 4816 1822
rect 4728 1716 4816 1776
rect 4728 1670 4757 1716
rect 4803 1670 4816 1716
rect 4728 1610 4816 1670
rect 4728 1564 4757 1610
rect 4803 1564 4816 1610
rect 4728 1503 4816 1564
rect 4728 1457 4757 1503
rect 4803 1457 4816 1503
rect 4728 1396 4816 1457
rect 4728 1350 4757 1396
rect 4803 1350 4816 1396
rect 4728 1337 4816 1350
<< mvndiffc >>
rect 2560 2702 2606 2748
rect 2560 2582 2606 2628
rect 2784 2702 2830 2748
rect 2784 2582 2830 2628
rect 2955 2590 3001 2636
rect 3179 2590 3225 2636
rect 4 898 50 944
rect 4 780 50 826
rect 4 663 50 709
rect 4 546 50 592
rect 228 898 274 944
rect 228 780 274 826
rect 228 663 274 709
rect 228 546 274 592
rect 452 898 498 944
rect 452 780 498 826
rect 452 663 498 709
rect 452 546 498 592
rect 676 898 722 944
rect 676 780 722 826
rect 676 663 722 709
rect 676 546 722 592
rect 900 898 946 944
rect 900 780 946 826
rect 900 663 946 709
rect 900 546 946 592
rect 1124 898 1170 944
rect 1124 780 1170 826
rect 1124 663 1170 709
rect 1124 546 1170 592
rect 1348 898 1394 944
rect 1946 921 1992 967
rect 1348 780 1394 826
rect 1348 663 1394 709
rect 1348 546 1394 592
rect 1554 805 1600 851
rect 1554 681 1600 727
rect 1554 557 1600 603
rect 1778 805 1824 851
rect 1778 681 1824 727
rect 1778 557 1824 603
rect 1946 799 1992 845
rect 1946 676 1992 722
rect 1946 553 1992 599
rect 2170 921 2216 967
rect 2170 799 2216 845
rect 2170 676 2216 722
rect 2170 553 2216 599
rect 2416 939 2462 985
rect 2416 812 2462 858
rect 2416 685 2462 731
rect 2416 557 2462 603
rect 2640 939 2686 985
rect 2640 812 2686 858
rect 2640 685 2686 731
rect 2640 557 2686 603
rect 2864 939 2910 985
rect 2864 812 2910 858
rect 2864 685 2910 731
rect 2864 557 2910 603
rect 3088 939 3134 985
rect 3088 812 3134 858
rect 3334 940 3380 986
rect 3334 820 3380 866
rect 3558 940 3604 986
rect 3558 820 3604 866
rect 3906 898 3952 944
rect 3088 685 3134 731
rect 3088 557 3134 603
rect 3906 774 3952 820
rect 3906 650 3952 696
rect 3906 526 3952 572
rect 3906 402 3952 448
rect 4130 898 4176 944
rect 4130 774 4176 820
rect 4130 650 4176 696
rect 4130 526 4176 572
rect 4130 402 4176 448
rect 4354 898 4400 944
rect 4354 774 4400 820
rect 4354 650 4400 696
rect 4354 526 4400 572
rect 4354 402 4400 448
rect 4578 898 4624 944
rect 4578 774 4624 820
rect 4578 650 4624 696
rect 4578 526 4624 572
rect 4578 402 4624 448
rect 4802 898 4848 944
rect 4802 774 4848 820
rect 4802 650 4848 696
rect 4802 526 4848 572
rect 4802 402 4848 448
<< mvpdiffc >>
rect 3861 2412 3907 2458
rect 3861 2306 3907 2352
rect 2336 2231 2382 2277
rect 1554 2020 1600 2066
rect 4 1935 50 1981
rect 4 1821 50 1867
rect 4 1707 50 1753
rect 4 1593 50 1639
rect 4 1479 50 1525
rect 4 1365 50 1411
rect 4 1251 50 1297
rect 228 1935 274 1981
rect 228 1821 274 1867
rect 228 1707 274 1753
rect 228 1593 274 1639
rect 228 1479 274 1525
rect 228 1365 274 1411
rect 228 1251 274 1297
rect 452 1935 498 1981
rect 452 1821 498 1867
rect 452 1707 498 1753
rect 452 1593 498 1639
rect 452 1479 498 1525
rect 452 1365 498 1411
rect 452 1251 498 1297
rect 676 1935 722 1981
rect 676 1821 722 1867
rect 676 1707 722 1753
rect 676 1593 722 1639
rect 676 1479 722 1525
rect 676 1365 722 1411
rect 676 1251 722 1297
rect 900 1935 946 1981
rect 900 1821 946 1867
rect 900 1707 946 1753
rect 900 1593 946 1639
rect 900 1479 946 1525
rect 900 1365 946 1411
rect 900 1251 946 1297
rect 1124 1935 1170 1981
rect 1124 1821 1170 1867
rect 1124 1707 1170 1753
rect 1124 1593 1170 1639
rect 1124 1479 1170 1525
rect 1124 1365 1170 1411
rect 1124 1251 1170 1297
rect 1348 1935 1394 1981
rect 1348 1821 1394 1867
rect 1348 1707 1394 1753
rect 1348 1593 1394 1639
rect 1348 1479 1394 1525
rect 1348 1365 1394 1411
rect 1348 1251 1394 1297
rect 1554 1916 1600 1962
rect 1554 1812 1600 1858
rect 1554 1708 1600 1754
rect 1554 1604 1600 1650
rect 1554 1500 1600 1546
rect 1554 1396 1600 1442
rect 1554 1292 1600 1338
rect 1778 2020 1824 2066
rect 1778 1916 1824 1962
rect 1778 1812 1824 1858
rect 1778 1708 1824 1754
rect 1778 1604 1824 1650
rect 1778 1500 1824 1546
rect 1778 1396 1824 1442
rect 1778 1292 1824 1338
rect 1946 2076 1992 2122
rect 1946 1973 1992 2019
rect 1946 1870 1992 1916
rect 1946 1767 1992 1813
rect 1946 1664 1992 1710
rect 1946 1560 1992 1606
rect 1946 1456 1992 1502
rect 1946 1352 1992 1398
rect 1946 1248 1992 1294
rect 2170 2076 2216 2122
rect 2336 2075 2382 2121
rect 2560 2231 2606 2277
rect 2560 2075 2606 2121
rect 2784 2231 2830 2277
rect 2942 2231 2988 2277
rect 2784 2075 2830 2121
rect 2942 2063 2988 2109
rect 2170 1973 2216 2019
rect 3166 2231 3212 2277
rect 3166 2063 3212 2109
rect 3861 2200 3907 2246
rect 3861 2094 3907 2140
rect 2170 1870 2216 1916
rect 2170 1767 2216 1813
rect 3861 1988 3907 2034
rect 3861 1882 3907 1928
rect 3334 1801 3380 1847
rect 2170 1664 2216 1710
rect 2170 1560 2216 1606
rect 2170 1456 2216 1502
rect 2170 1352 2216 1398
rect 2170 1248 2216 1294
rect 2416 1674 2462 1720
rect 2416 1547 2462 1593
rect 2416 1420 2462 1466
rect 2416 1292 2462 1338
rect 2640 1674 2686 1720
rect 2640 1547 2686 1593
rect 2640 1420 2686 1466
rect 2640 1292 2686 1338
rect 2864 1674 2910 1720
rect 2864 1547 2910 1593
rect 2864 1420 2910 1466
rect 2864 1292 2910 1338
rect 3088 1674 3134 1720
rect 3088 1547 3134 1593
rect 3088 1420 3134 1466
rect 3334 1674 3380 1720
rect 3334 1547 3380 1593
rect 3334 1419 3380 1465
rect 3558 1801 3604 1847
rect 3558 1674 3604 1720
rect 3558 1547 3604 1593
rect 3558 1419 3604 1465
rect 3861 1776 3907 1822
rect 3861 1670 3907 1716
rect 3861 1564 3907 1610
rect 3861 1457 3907 1503
rect 3088 1292 3134 1338
rect 3861 1350 3907 1396
rect 4085 2412 4131 2458
rect 4085 2306 4131 2352
rect 4085 2200 4131 2246
rect 4085 2094 4131 2140
rect 4085 1988 4131 2034
rect 4085 1882 4131 1928
rect 4085 1776 4131 1822
rect 4085 1670 4131 1716
rect 4085 1564 4131 1610
rect 4085 1457 4131 1503
rect 4085 1350 4131 1396
rect 4309 2412 4355 2458
rect 4309 2306 4355 2352
rect 4309 2200 4355 2246
rect 4309 2094 4355 2140
rect 4309 1988 4355 2034
rect 4309 1882 4355 1928
rect 4309 1776 4355 1822
rect 4309 1670 4355 1716
rect 4309 1564 4355 1610
rect 4309 1457 4355 1503
rect 4309 1350 4355 1396
rect 4533 2412 4579 2458
rect 4533 2306 4579 2352
rect 4533 2200 4579 2246
rect 4533 2094 4579 2140
rect 4533 1988 4579 2034
rect 4533 1882 4579 1928
rect 4533 1776 4579 1822
rect 4533 1670 4579 1716
rect 4533 1564 4579 1610
rect 4533 1457 4579 1503
rect 4533 1350 4579 1396
rect 4757 2412 4803 2458
rect 4757 2306 4803 2352
rect 4757 2200 4803 2246
rect 4757 2094 4803 2140
rect 4757 1988 4803 2034
rect 4757 1882 4803 1928
rect 4757 1776 4803 1822
rect 4757 1670 4803 1716
rect 4757 1564 4803 1610
rect 4757 1457 4803 1503
rect 4757 1350 4803 1396
<< psubdiff >>
rect 3438 2700 3598 2760
rect 3438 2654 3495 2700
rect 3541 2654 3598 2700
rect 3438 2595 3598 2654
rect -352 891 -268 910
rect -352 563 -333 891
rect -287 563 -268 891
rect -352 544 -268 563
rect -64 361 1430 380
rect -64 315 -45 361
rect 1411 315 1430 361
rect -64 296 1430 315
rect 4913 -63 4997 -44
rect 4913 -297 4932 -63
rect 4978 -297 4997 -63
rect 4913 -316 4997 -297
<< nsubdiff >>
rect -222 2200 1178 2219
rect -222 2154 -203 2200
rect 1159 2154 1178 2200
rect -222 2135 1178 2154
rect -387 1773 -232 1830
rect -387 1727 -333 1773
rect -287 1727 -232 1773
rect -387 1610 -232 1727
rect -387 1564 -333 1610
rect -287 1564 -232 1610
rect -387 1447 -232 1564
rect -387 1401 -333 1447
rect -287 1401 -232 1447
rect -387 1343 -232 1401
rect 4913 2350 4997 2369
rect 4913 1552 4932 2350
rect 4978 1552 4997 2350
rect 4913 1533 4997 1552
<< psubdiffcont >>
rect 3495 2654 3541 2700
rect -333 563 -287 891
rect -45 315 1411 361
rect 4932 -297 4978 -63
<< nsubdiffcont >>
rect -203 2154 1159 2200
rect -333 1727 -287 1773
rect -333 1564 -287 1610
rect -333 1401 -287 1447
rect 4932 1552 4978 2350
<< polysilicon >>
rect 2635 2761 2755 2835
rect 3030 2673 3150 2746
rect 2635 2465 2755 2569
rect 4030 2722 4728 2741
rect 4030 2676 4049 2722
rect 4189 2676 4728 2722
rect 4030 2666 4728 2676
rect 4030 2657 4504 2666
rect 3714 2601 3798 2620
rect 3714 2555 3733 2601
rect 3779 2597 3798 2601
rect 3779 2555 4280 2597
rect 2635 2422 2678 2465
rect 2411 2419 2678 2422
rect 2724 2419 2755 2465
rect 3030 2445 3150 2553
rect 3714 2536 4280 2555
rect 3936 2471 4056 2536
rect 4160 2471 4280 2536
rect 4384 2471 4504 2657
rect 4608 2471 4728 2666
rect 3030 2426 3422 2445
rect 3030 2422 3357 2426
rect 2411 2361 2755 2419
rect 2411 2290 2531 2361
rect 2635 2290 2755 2361
rect 3017 2380 3357 2422
rect 3403 2380 3422 2426
rect 3017 2361 3422 2380
rect 3017 2290 3137 2361
rect 2021 2135 2141 2179
rect 1629 2079 1749 2123
rect 79 1994 199 2038
rect 303 1994 423 2038
rect 527 1994 647 2038
rect 751 1994 871 2038
rect 975 1994 1095 2038
rect 1199 1994 1319 2038
rect 79 1166 199 1238
rect 303 1166 423 1238
rect 527 1166 647 1238
rect 751 1166 871 1238
rect 975 1166 1095 1238
rect 1199 1166 1319 1238
rect 79 1147 1521 1166
rect 79 1105 1456 1147
rect 79 957 199 1105
rect 303 957 423 1105
rect 527 957 647 1105
rect 751 957 871 1105
rect 975 957 1095 1105
rect 1199 1101 1456 1105
rect 1502 1101 1521 1147
rect 1199 1082 1521 1101
rect 1199 957 1319 1082
rect 1629 864 1749 1279
rect 2411 1990 2531 2062
rect 2635 1990 2755 2062
rect 3017 2006 3137 2050
rect 3409 1998 3529 2017
rect 3409 1952 3444 1998
rect 3490 1952 3529 1998
rect 2491 1858 3154 1877
rect 3409 1860 3529 1952
rect 2491 1812 3089 1858
rect 3135 1812 3154 1858
rect 2491 1793 3154 1812
rect 2491 1733 2611 1793
rect 2715 1733 2835 1793
rect 2939 1733 3059 1793
rect 2491 1235 2611 1279
rect 2715 1235 2835 1279
rect 2939 1235 3059 1279
rect 2021 1124 2141 1235
rect 1853 1105 2141 1124
rect 1853 1059 1872 1105
rect 2012 1059 2141 1105
rect 1853 1040 2141 1059
rect 2021 980 2141 1040
rect 2491 998 2611 1042
rect 2715 998 2835 1042
rect 2939 998 3059 1042
rect 3409 999 3529 1406
rect 3936 1293 4056 1337
rect 4160 1293 4280 1337
rect 4384 1293 4504 1337
rect 4608 1293 4728 1337
rect 3981 1136 4462 1155
rect 3981 1090 4303 1136
rect 4443 1090 4462 1136
rect 3981 1071 4462 1090
rect 79 489 199 533
rect 303 489 423 533
rect 527 489 647 533
rect 751 489 871 533
rect 975 489 1095 533
rect 1199 489 1319 533
rect 1629 393 1749 544
rect 3981 957 4101 1071
rect 4205 957 4325 1071
rect 4429 957 4549 1001
rect 4653 957 4773 1001
rect 2021 480 2141 540
rect 2491 484 2611 544
rect 2715 484 2835 544
rect 2939 484 3059 544
rect 3409 511 3529 807
rect 3240 488 3324 507
rect 3240 484 3259 488
rect 2021 461 2214 480
rect 2021 415 2055 461
rect 2195 415 2214 461
rect 2491 442 3259 484
rect 3305 442 3324 488
rect 2491 423 3324 442
rect 3409 492 3588 511
rect 3409 446 3523 492
rect 3569 446 3588 492
rect 3409 427 3588 446
rect 2021 396 2214 415
rect 1597 374 1775 393
rect 1597 328 1616 374
rect 1756 328 1775 374
rect 3981 345 4101 389
rect 4205 345 4325 389
rect 1597 309 1775 328
rect 4429 216 4549 389
rect 4653 216 4773 389
rect 4429 197 4773 216
rect 4429 151 4525 197
rect 4665 151 4773 197
rect 4429 132 4773 151
<< polycontact >>
rect 4049 2676 4189 2722
rect 3733 2555 3779 2601
rect 2678 2419 2724 2465
rect 3357 2380 3403 2426
rect 1456 1101 1502 1147
rect 3444 1952 3490 1998
rect 3089 1812 3135 1858
rect 1872 1059 2012 1105
rect 4303 1090 4443 1136
rect 2055 415 2195 461
rect 3259 442 3305 488
rect 3523 446 3569 492
rect 1616 328 1756 374
rect 4525 151 4665 197
<< metal1 >>
rect 2784 2853 2941 3324
rect 2784 2778 3519 2853
rect 2560 2748 2606 2761
rect 2170 2727 2478 2747
rect 2170 2675 2200 2727
rect 2252 2675 2386 2727
rect 2438 2675 2478 2727
rect 2170 2655 2478 2675
rect 1124 2211 1170 2239
rect -214 2200 1170 2211
rect -214 2154 -203 2200
rect 1159 2154 1170 2200
rect -214 2143 1170 2154
rect 4 1981 50 1994
rect 4 1867 50 1935
rect -356 1810 -264 1811
rect -367 1781 -252 1810
rect -367 1729 -336 1781
rect -284 1729 -252 1781
rect -367 1727 -333 1729
rect -287 1727 -252 1729
rect -367 1610 -252 1727
rect -367 1595 -333 1610
rect -287 1595 -252 1610
rect -367 1543 -336 1595
rect -284 1543 -252 1595
rect -367 1447 -252 1543
rect -367 1401 -333 1447
rect -287 1401 -252 1447
rect -367 1364 -252 1401
rect 4 1753 50 1821
rect 4 1639 50 1707
rect 194 1981 310 2143
rect 194 1935 228 1981
rect 274 1935 310 1981
rect 194 1867 310 1935
rect 194 1821 228 1867
rect 274 1821 310 1867
rect 194 1781 310 1821
rect 194 1729 226 1781
rect 278 1729 310 1781
rect 194 1707 228 1729
rect 274 1707 310 1729
rect 194 1665 310 1707
rect 452 1981 498 1994
rect 452 1867 498 1935
rect 452 1753 498 1821
rect 4 1525 50 1593
rect 206 1639 298 1665
rect 206 1595 228 1639
rect 274 1595 298 1639
rect 206 1543 226 1595
rect 278 1543 298 1595
rect 206 1525 298 1543
rect 206 1503 228 1525
rect 4 1411 50 1479
rect 4 1297 50 1365
rect 4 1166 50 1251
rect 274 1503 298 1525
rect 452 1639 498 1707
rect 642 1981 758 2143
rect 642 1935 676 1981
rect 722 1935 758 1981
rect 642 1867 758 1935
rect 642 1821 676 1867
rect 722 1821 758 1867
rect 642 1781 758 1821
rect 642 1729 672 1781
rect 724 1729 758 1781
rect 642 1707 676 1729
rect 722 1707 758 1729
rect 642 1665 758 1707
rect 900 1981 946 1994
rect 900 1867 946 1935
rect 900 1753 946 1821
rect 1124 1981 1170 2143
rect 1946 2122 1992 2135
rect 1554 2066 1600 2079
rect 1124 1867 1170 1935
rect 1124 1811 1170 1821
rect 1348 1981 1394 1994
rect 1348 1867 1394 1935
rect 452 1525 498 1593
rect 228 1411 274 1479
rect 228 1297 274 1365
rect 228 1238 274 1251
rect 652 1639 744 1665
rect 652 1595 676 1639
rect 722 1595 744 1639
rect 652 1543 672 1595
rect 724 1543 744 1595
rect 652 1525 744 1543
rect 652 1503 676 1525
rect 452 1411 498 1479
rect 452 1297 498 1365
rect 452 1166 498 1251
rect 722 1503 744 1525
rect 900 1639 946 1707
rect 900 1525 946 1593
rect 676 1411 722 1479
rect 676 1297 722 1365
rect 676 1238 722 1251
rect 1100 1781 1192 1811
rect 1100 1729 1120 1781
rect 1172 1729 1192 1781
rect 1100 1707 1124 1729
rect 1170 1707 1192 1729
rect 1100 1639 1192 1707
rect 1100 1595 1124 1639
rect 1170 1595 1192 1639
rect 1100 1543 1120 1595
rect 1172 1543 1192 1595
rect 1100 1525 1192 1543
rect 1100 1503 1124 1525
rect 900 1411 946 1479
rect 900 1297 946 1365
rect 900 1166 946 1251
rect 1170 1503 1192 1525
rect 1348 1753 1394 1821
rect 1554 1962 1600 2020
rect 1554 1858 1600 1916
rect 1554 1811 1600 1812
rect 1778 2066 1824 2079
rect 1778 1962 1824 2020
rect 1778 1858 1824 1916
rect 1348 1639 1394 1707
rect 1348 1525 1394 1593
rect 1124 1411 1170 1479
rect 1124 1297 1170 1365
rect 1124 1238 1170 1251
rect 1531 1781 1623 1811
rect 1531 1729 1551 1781
rect 1603 1729 1623 1781
rect 1531 1708 1554 1729
rect 1600 1708 1623 1729
rect 1531 1650 1623 1708
rect 1531 1604 1554 1650
rect 1600 1604 1623 1650
rect 1531 1595 1623 1604
rect 1531 1543 1551 1595
rect 1603 1543 1623 1595
rect 1531 1503 1554 1543
rect 1348 1411 1394 1479
rect 1348 1297 1394 1365
rect 1600 1503 1623 1543
rect 1778 1754 1824 1812
rect 1946 2019 1992 2076
rect 1946 1916 1992 1973
rect 1946 1813 1992 1870
rect 1778 1650 1824 1708
rect 1778 1546 1824 1604
rect 1554 1442 1600 1500
rect 1554 1338 1600 1396
rect 1554 1279 1600 1292
rect 1923 1781 1946 1811
rect 2170 2122 2216 2655
rect 2560 2628 2606 2702
rect 2170 2019 2216 2076
rect 2312 2282 2404 2312
rect 2312 2230 2332 2282
rect 2384 2230 2404 2282
rect 2312 2121 2404 2230
rect 2312 2096 2336 2121
rect 2382 2096 2404 2121
rect 2312 2044 2332 2096
rect 2384 2044 2404 2096
rect 2312 2004 2404 2044
rect 2560 2277 2606 2582
rect 2784 2748 3001 2778
rect 2830 2702 3001 2748
rect 2784 2636 3001 2702
rect 3447 2751 3519 2778
rect 3709 2790 3801 2830
rect 3447 2700 3589 2751
rect 2784 2628 2955 2636
rect 2830 2590 2955 2628
rect 2830 2582 3001 2590
rect 2784 2553 3001 2582
rect 3131 2636 3247 2699
rect 3131 2590 3179 2636
rect 3225 2590 3247 2636
rect 3447 2654 3495 2700
rect 3541 2654 3589 2700
rect 3447 2604 3589 2654
rect 3709 2738 3729 2790
rect 3781 2738 3801 2790
rect 3709 2604 3801 2738
rect 3918 2727 4226 2747
rect 3918 2675 3948 2727
rect 4000 2722 4134 2727
rect 4186 2722 4226 2727
rect 4000 2676 4049 2722
rect 4189 2676 4226 2722
rect 4000 2675 4134 2676
rect 4186 2675 4226 2676
rect 3918 2655 4226 2675
rect 3131 2476 3247 2590
rect 3709 2552 3729 2604
rect 3781 2552 3801 2604
rect 3709 2511 3801 2552
rect 3861 2563 4803 2609
rect 2667 2465 3247 2476
rect 2667 2419 2678 2465
rect 2724 2419 3247 2465
rect 3861 2458 3907 2563
rect 2667 2402 3247 2419
rect 2560 2121 2606 2231
rect 2170 1916 2216 1973
rect 2560 1923 2606 2075
rect 2761 2282 2853 2312
rect 2761 2230 2781 2282
rect 2833 2230 2853 2282
rect 2761 2121 2853 2230
rect 2761 2096 2784 2121
rect 2830 2096 2853 2121
rect 2761 2044 2781 2096
rect 2833 2044 2853 2096
rect 2761 2004 2853 2044
rect 2919 2282 3011 2312
rect 2919 2230 2939 2282
rect 2991 2230 3011 2282
rect 2919 2109 3011 2230
rect 3131 2277 3247 2402
rect 3324 2426 3580 2445
rect 3324 2380 3357 2426
rect 3403 2415 3580 2426
rect 3324 2363 3363 2380
rect 3415 2363 3580 2415
rect 3324 2290 3580 2363
rect 3861 2352 3907 2412
rect 3131 2231 3166 2277
rect 3212 2231 3247 2277
rect 3131 2152 3247 2231
rect 3861 2246 3907 2306
rect 2919 2096 2942 2109
rect 2988 2096 3011 2109
rect 2919 2044 2939 2096
rect 2991 2044 3011 2096
rect 3166 2109 3212 2152
rect 3861 2140 3907 2200
rect 3166 2050 3212 2063
rect 2919 2004 3011 2044
rect 3263 2023 3602 2064
rect 3263 2004 3300 2023
rect 3098 1971 3300 2004
rect 3352 1998 3512 2023
rect 3352 1971 3444 1998
rect 3098 1952 3444 1971
rect 3490 1971 3512 1998
rect 3564 1971 3602 2023
rect 3490 1952 3602 1971
rect 3098 1929 3602 1952
rect 3861 2034 3907 2094
rect 2170 1813 2216 1870
rect 1992 1781 2015 1811
rect 1923 1729 1943 1781
rect 1995 1729 2015 1781
rect 1923 1710 2015 1729
rect 1923 1664 1946 1710
rect 1992 1664 2015 1710
rect 1923 1606 2015 1664
rect 1923 1595 1946 1606
rect 1992 1595 2015 1606
rect 1923 1543 1943 1595
rect 1995 1543 2015 1595
rect 1923 1503 2015 1543
rect 2170 1710 2216 1767
rect 2170 1606 2216 1664
rect 1778 1442 1824 1500
rect 1778 1338 1824 1396
rect 1348 1166 1394 1251
rect 4 1046 1394 1166
rect 1468 1158 1648 1166
rect 1445 1154 1648 1158
rect 1445 1147 1480 1154
rect 1445 1101 1456 1147
rect 1636 1102 1648 1154
rect 1502 1101 1648 1102
rect 1445 1090 1648 1101
rect 1778 1116 1824 1292
rect 1946 1502 1992 1503
rect 1946 1398 1992 1456
rect 1946 1294 1992 1352
rect 1946 1235 1992 1248
rect 2170 1502 2216 1560
rect 2170 1398 2216 1456
rect 2170 1294 2216 1352
rect 1778 1105 2023 1116
rect 4 944 50 1046
rect -356 908 -264 938
rect -356 856 -336 908
rect -284 856 -264 908
rect -356 722 -333 856
rect -287 722 -264 856
rect -356 670 -336 722
rect -284 670 -264 722
rect -356 630 -333 670
rect -344 563 -333 630
rect -287 630 -264 670
rect 228 944 274 957
rect 206 908 228 938
rect 452 944 498 1046
rect 274 908 298 938
rect 206 901 226 908
rect 4 826 50 898
rect 4 709 50 780
rect -287 563 -276 630
rect -344 552 -276 563
rect 4 592 50 663
rect 4 533 50 546
rect 194 856 226 901
rect 278 901 298 908
rect 278 856 310 901
rect 194 826 310 856
rect 194 780 228 826
rect 274 780 310 826
rect 194 722 310 780
rect 194 670 226 722
rect 278 670 310 722
rect 194 663 228 670
rect 274 663 310 670
rect 194 592 310 663
rect 194 546 228 592
rect 274 546 310 592
rect 194 372 310 546
rect 676 944 722 957
rect 652 908 676 938
rect 900 944 946 1046
rect 722 908 744 938
rect 652 901 672 908
rect 452 826 498 898
rect 452 709 498 780
rect 452 592 498 663
rect 452 533 498 546
rect 642 856 672 901
rect 724 901 744 908
rect 724 856 758 901
rect 642 826 758 856
rect 642 780 676 826
rect 722 780 758 826
rect 642 722 758 780
rect 642 670 672 722
rect 724 670 758 722
rect 642 663 676 670
rect 722 663 758 670
rect 642 592 758 663
rect 642 546 676 592
rect 722 546 758 592
rect 642 372 758 546
rect 1124 944 1170 957
rect 1102 908 1124 938
rect 1348 944 1394 1046
rect 1170 908 1194 938
rect 1102 901 1122 908
rect 900 826 946 898
rect 900 709 946 780
rect 900 592 946 663
rect 900 533 946 546
rect 1090 856 1122 901
rect 1174 901 1194 908
rect 1174 856 1206 901
rect 1090 826 1206 856
rect 1090 780 1124 826
rect 1170 780 1206 826
rect 1090 722 1206 780
rect 1090 670 1122 722
rect 1174 670 1206 722
rect 1090 663 1124 670
rect 1170 663 1206 670
rect 1090 592 1206 663
rect 1090 546 1124 592
rect 1170 546 1206 592
rect 1090 372 1206 546
rect 1348 826 1394 898
rect 1778 1059 1872 1105
rect 2012 1059 2023 1105
rect 1778 1048 2023 1059
rect 1554 851 1600 864
rect 1348 709 1394 780
rect 1348 592 1394 663
rect 1348 533 1394 546
rect 1531 815 1554 845
rect 1778 851 1824 1048
rect 1600 815 1623 845
rect 1531 763 1551 815
rect 1603 763 1623 815
rect 1531 727 1623 763
rect 1531 681 1554 727
rect 1600 681 1623 727
rect 1531 629 1623 681
rect 1531 577 1551 629
rect 1603 577 1623 629
rect 1531 557 1554 577
rect 1600 557 1623 577
rect 1531 537 1623 557
rect 1946 967 1992 980
rect 1946 845 1992 921
rect 2170 967 2216 1248
rect 2170 845 2216 921
rect 1778 727 1824 805
rect 1778 603 1824 681
rect 1778 544 1824 557
rect 1923 815 1946 845
rect 1992 815 2015 845
rect 1923 763 1943 815
rect 1995 763 2015 815
rect 1923 722 2015 763
rect 1923 676 1946 722
rect 1992 676 2015 722
rect 1923 629 2015 676
rect 1923 577 1943 629
rect 1995 577 2015 629
rect 1923 553 1946 577
rect 1992 553 2015 577
rect 1923 537 2015 553
rect 2170 722 2216 799
rect 2170 599 2216 676
rect 2170 540 2216 553
rect 2382 1804 2946 1923
rect 3098 1869 3170 1929
rect 2382 1720 2498 1804
rect 2640 1722 2686 1733
rect 2382 1674 2416 1720
rect 2462 1674 2498 1720
rect 2382 1593 2498 1674
rect 2382 1547 2416 1593
rect 2462 1547 2498 1593
rect 2382 1466 2498 1547
rect 2382 1420 2416 1466
rect 2462 1420 2498 1466
rect 2382 1338 2498 1420
rect 2382 1292 2416 1338
rect 2462 1292 2498 1338
rect 2382 985 2498 1292
rect 2382 939 2416 985
rect 2462 939 2498 985
rect 2382 858 2498 939
rect 2382 812 2416 858
rect 2462 812 2498 858
rect 2382 731 2498 812
rect 2382 685 2416 731
rect 2462 685 2498 731
rect 2382 603 2498 685
rect 2382 557 2416 603
rect 2462 557 2498 603
rect 2382 544 2498 557
rect 2606 1720 2722 1722
rect 2606 1674 2640 1720
rect 2686 1674 2722 1720
rect 2606 1593 2722 1674
rect 2606 1547 2640 1593
rect 2686 1547 2722 1593
rect 2606 1466 2722 1547
rect 2606 1420 2640 1466
rect 2686 1420 2722 1466
rect 2606 1364 2722 1420
rect 2606 1312 2638 1364
rect 2690 1312 2722 1364
rect 2606 1292 2640 1312
rect 2686 1292 2722 1312
rect 2606 1178 2722 1292
rect 2606 1126 2638 1178
rect 2690 1126 2722 1178
rect 2606 985 2722 1126
rect 2606 939 2640 985
rect 2686 939 2722 985
rect 2606 858 2722 939
rect 2606 812 2640 858
rect 2686 812 2722 858
rect 2606 731 2722 812
rect 2606 685 2640 731
rect 2686 685 2722 731
rect 2606 603 2722 685
rect 2606 557 2640 603
rect 2686 557 2722 603
rect 2160 472 2206 476
rect 2044 461 2206 472
rect 2044 415 2055 461
rect 2195 415 2206 461
rect 2044 404 2206 415
rect 1600 376 1780 388
rect -56 361 1422 372
rect -56 315 -45 361
rect 1411 315 1422 361
rect -56 304 1422 315
rect 1600 324 1612 376
rect 1768 324 1780 376
rect 1600 312 1780 324
rect 2160 237 2206 404
rect 2606 472 2722 557
rect 2830 1720 2946 1804
rect 3078 1858 3170 1869
rect 3861 1928 3907 1988
rect 3078 1812 3089 1858
rect 3135 1812 3170 1858
rect 3078 1801 3170 1812
rect 3334 1847 3380 1860
rect 3558 1847 3604 1860
rect 3088 1724 3134 1733
rect 2830 1674 2864 1720
rect 2910 1674 2946 1720
rect 2830 1593 2946 1674
rect 2830 1547 2864 1593
rect 2910 1547 2946 1593
rect 2830 1466 2946 1547
rect 2830 1420 2864 1466
rect 2910 1420 2946 1466
rect 2830 1338 2946 1420
rect 2830 1292 2864 1338
rect 2910 1292 2946 1338
rect 2830 985 2946 1292
rect 2830 939 2864 985
rect 2910 939 2946 985
rect 2830 858 2946 939
rect 2830 812 2864 858
rect 2910 812 2946 858
rect 2830 731 2946 812
rect 2830 685 2864 731
rect 2910 685 2946 731
rect 2830 603 2946 685
rect 2830 557 2864 603
rect 2910 557 2946 603
rect 2830 544 2946 557
rect 3054 1720 3170 1724
rect 3054 1674 3088 1720
rect 3134 1674 3170 1720
rect 3054 1593 3170 1674
rect 3054 1547 3088 1593
rect 3134 1547 3170 1593
rect 3054 1466 3170 1547
rect 3054 1420 3088 1466
rect 3134 1420 3170 1466
rect 3054 1364 3170 1420
rect 3054 1338 3097 1364
rect 3054 1292 3088 1338
rect 3149 1312 3170 1364
rect 3134 1292 3170 1312
rect 3054 1178 3170 1292
rect 3054 1126 3097 1178
rect 3149 1126 3170 1178
rect 3054 985 3170 1126
rect 3054 939 3088 985
rect 3134 939 3170 985
rect 3054 858 3170 939
rect 3334 1720 3380 1801
rect 3334 1593 3380 1674
rect 3334 1465 3380 1547
rect 3525 1801 3558 1811
rect 3861 1822 3907 1882
rect 3604 1801 3617 1811
rect 3525 1781 3617 1801
rect 3525 1729 3545 1781
rect 3597 1729 3617 1781
rect 3525 1720 3617 1729
rect 3525 1674 3558 1720
rect 3604 1674 3617 1720
rect 3525 1595 3617 1674
rect 3525 1543 3545 1595
rect 3597 1593 3617 1595
rect 3604 1547 3617 1593
rect 3597 1543 3617 1547
rect 3525 1503 3617 1543
rect 3861 1716 3907 1776
rect 3861 1610 3907 1670
rect 3861 1503 3907 1564
rect 3334 986 3380 1419
rect 3558 1465 3604 1503
rect 3558 1406 3604 1419
rect 3861 1396 3907 1457
rect 3861 1337 3907 1350
rect 4085 2458 4131 2471
rect 4085 2352 4131 2412
rect 4085 2246 4131 2306
rect 4085 2140 4131 2200
rect 4085 2034 4131 2094
rect 4085 1928 4131 1988
rect 4085 1822 4131 1882
rect 4085 1716 4131 1776
rect 4085 1610 4131 1670
rect 4085 1503 4131 1564
rect 4085 1396 4131 1457
rect 4085 1194 4131 1350
rect 4309 2458 4355 2563
rect 4309 2352 4355 2412
rect 4533 2458 4579 2471
rect 4533 2352 4579 2412
rect 4309 2246 4355 2306
rect 4309 2140 4355 2200
rect 4309 2034 4355 2094
rect 4510 2306 4533 2312
rect 4757 2458 4803 2563
rect 4757 2352 4803 2412
rect 4579 2306 4602 2312
rect 4510 2282 4602 2306
rect 4510 2230 4530 2282
rect 4582 2230 4602 2282
rect 4510 2200 4533 2230
rect 4579 2200 4602 2230
rect 4510 2140 4602 2200
rect 4510 2096 4533 2140
rect 4579 2096 4602 2140
rect 4510 2044 4530 2096
rect 4582 2044 4602 2096
rect 4510 2034 4602 2044
rect 4510 2004 4533 2034
rect 4309 1928 4355 1988
rect 4309 1822 4355 1882
rect 4579 2004 4602 2034
rect 4921 2350 4989 2361
rect 4921 2312 4932 2350
rect 4757 2246 4803 2306
rect 4757 2140 4803 2200
rect 4757 2034 4803 2094
rect 4533 1928 4579 1988
rect 4533 1822 4579 1882
rect 4309 1716 4355 1776
rect 4309 1610 4355 1670
rect 4309 1503 4355 1564
rect 4510 1781 4533 1811
rect 4909 2282 4932 2312
rect 4978 2312 4989 2350
rect 4978 2282 5001 2312
rect 4909 2230 4929 2282
rect 4981 2230 5001 2282
rect 4909 2096 4932 2230
rect 4978 2096 5001 2230
rect 4909 2044 4929 2096
rect 4981 2044 5001 2096
rect 4909 2004 4932 2044
rect 4757 1928 4803 1988
rect 4757 1822 4803 1882
rect 4579 1781 4602 1811
rect 4510 1729 4530 1781
rect 4582 1729 4602 1781
rect 4510 1716 4602 1729
rect 4510 1670 4533 1716
rect 4579 1670 4602 1716
rect 4510 1610 4602 1670
rect 4510 1595 4533 1610
rect 4579 1595 4602 1610
rect 4510 1543 4530 1595
rect 4582 1543 4602 1595
rect 4510 1503 4602 1543
rect 4921 1811 4932 2004
rect 4757 1716 4803 1776
rect 4757 1610 4803 1670
rect 4757 1503 4803 1564
rect 4909 1781 4932 1811
rect 4978 2004 5001 2044
rect 4978 1811 4989 2004
rect 4978 1781 5001 1811
rect 4909 1729 4929 1781
rect 4981 1729 5001 1781
rect 4909 1595 4932 1729
rect 4978 1595 5001 1729
rect 4909 1543 4929 1595
rect 4981 1543 5001 1595
rect 4909 1503 5001 1543
rect 4309 1396 4355 1457
rect 4309 1337 4355 1350
rect 4533 1396 4579 1457
rect 4533 1337 4579 1350
rect 4757 1396 4803 1457
rect 4757 1337 4803 1350
rect 3951 1182 4131 1194
rect 3951 1130 3963 1182
rect 4119 1130 4131 1182
rect 3951 1118 4131 1130
rect 3334 866 3380 940
rect 3558 986 3604 999
rect 4085 957 4131 1118
rect 4280 1139 4460 1151
rect 4280 1087 4292 1139
rect 4448 1087 4460 1139
rect 4280 1075 4460 1087
rect 3558 938 3604 940
rect 3906 944 3952 957
rect 3054 812 3088 858
rect 3134 812 3170 858
rect 3054 731 3170 812
rect 3054 685 3088 731
rect 3134 685 3170 731
rect 3054 603 3170 685
rect 3054 557 3088 603
rect 3134 557 3170 603
rect 3054 472 3170 557
rect 3282 820 3334 863
rect 3282 807 3380 820
rect 3547 908 3639 938
rect 3547 866 3567 908
rect 3547 820 3558 866
rect 3619 856 3639 908
rect 3604 820 3639 856
rect 3282 499 3354 807
rect 3547 722 3639 820
rect 3547 670 3567 722
rect 3619 670 3639 722
rect 3547 630 3639 670
rect 3906 820 3952 898
rect 4085 944 4176 957
rect 4085 898 4130 944
rect 4085 862 4176 898
rect 3906 696 3952 774
rect 3906 572 3952 650
rect 2606 353 3170 472
rect 3248 488 3354 499
rect 3248 442 3259 488
rect 3305 442 3354 488
rect 3248 432 3354 442
rect 3432 493 3771 534
rect 3432 441 3469 493
rect 3521 492 3681 493
rect 3521 446 3523 492
rect 3569 446 3681 492
rect 3521 441 3681 446
rect 3733 441 3771 493
rect 3248 431 3316 432
rect 3432 400 3771 441
rect 3906 448 3952 526
rect 3906 330 3952 402
rect 4130 820 4176 862
rect 4130 696 4176 774
rect 4130 572 4176 650
rect 4130 448 4176 526
rect 4130 389 4176 402
rect 4354 944 4400 957
rect 4578 944 4624 957
rect 4354 820 4400 898
rect 4354 696 4400 774
rect 4354 572 4400 650
rect 4555 908 4578 938
rect 4802 944 4848 957
rect 4624 908 4647 938
rect 4555 856 4575 908
rect 4627 856 4647 908
rect 4555 820 4647 856
rect 4555 774 4578 820
rect 4624 774 4647 820
rect 4555 722 4647 774
rect 4555 670 4575 722
rect 4627 670 4647 722
rect 4555 650 4578 670
rect 4624 650 4647 670
rect 4555 630 4647 650
rect 4802 820 4848 898
rect 4802 696 4848 774
rect 4354 448 4400 526
rect 4354 330 4400 402
rect 4578 572 4624 630
rect 4578 448 4624 526
rect 4578 389 4624 402
rect 4802 572 4848 650
rect 4802 448 4848 526
rect 4802 330 4848 402
rect 3906 284 4848 330
rect 2160 197 3783 237
rect 4514 197 4676 208
rect 2160 191 4525 197
rect 3702 151 4525 191
rect 4665 151 4676 197
rect 4514 140 4676 151
rect 4909 -62 5001 -32
rect 4909 -114 4929 -62
rect 4981 -114 5001 -62
rect 4909 -248 4932 -114
rect 4978 -248 5001 -114
rect 4909 -300 4929 -248
rect 4981 -300 5001 -248
rect 4909 -340 5001 -300
<< via1 >>
rect 2200 2675 2252 2727
rect 2386 2675 2438 2727
rect -336 1773 -284 1781
rect -336 1729 -333 1773
rect -333 1729 -287 1773
rect -287 1729 -284 1773
rect -336 1564 -333 1595
rect -333 1564 -287 1595
rect -287 1564 -284 1595
rect -336 1543 -284 1564
rect 226 1753 278 1781
rect 226 1729 228 1753
rect 228 1729 274 1753
rect 274 1729 278 1753
rect 226 1593 228 1595
rect 228 1593 274 1595
rect 274 1593 278 1595
rect 226 1543 278 1593
rect 672 1753 724 1781
rect 672 1729 676 1753
rect 676 1729 722 1753
rect 722 1729 724 1753
rect 672 1593 676 1595
rect 676 1593 722 1595
rect 722 1593 724 1595
rect 672 1543 724 1593
rect 1120 1753 1172 1781
rect 1120 1729 1124 1753
rect 1124 1729 1170 1753
rect 1170 1729 1172 1753
rect 1120 1593 1124 1595
rect 1124 1593 1170 1595
rect 1170 1593 1172 1595
rect 1120 1543 1172 1593
rect 1551 1754 1603 1781
rect 1551 1729 1554 1754
rect 1554 1729 1600 1754
rect 1600 1729 1603 1754
rect 1551 1546 1603 1595
rect 1551 1543 1554 1546
rect 1554 1543 1600 1546
rect 1600 1543 1603 1546
rect 2332 2277 2384 2282
rect 2332 2231 2336 2277
rect 2336 2231 2382 2277
rect 2382 2231 2384 2277
rect 2332 2230 2384 2231
rect 2332 2075 2336 2096
rect 2336 2075 2382 2096
rect 2382 2075 2384 2096
rect 2332 2044 2384 2075
rect 3729 2738 3781 2790
rect 3948 2675 4000 2727
rect 4134 2722 4186 2727
rect 4134 2676 4186 2722
rect 4134 2675 4186 2676
rect 3729 2601 3781 2604
rect 3729 2555 3733 2601
rect 3733 2555 3779 2601
rect 3779 2555 3781 2601
rect 3729 2552 3781 2555
rect 2781 2277 2833 2282
rect 2781 2231 2784 2277
rect 2784 2231 2830 2277
rect 2830 2231 2833 2277
rect 2781 2230 2833 2231
rect 2781 2075 2784 2096
rect 2784 2075 2830 2096
rect 2830 2075 2833 2096
rect 2781 2044 2833 2075
rect 2939 2277 2991 2282
rect 2939 2231 2942 2277
rect 2942 2231 2988 2277
rect 2988 2231 2991 2277
rect 2939 2230 2991 2231
rect 3363 2380 3403 2415
rect 3403 2380 3415 2415
rect 3363 2363 3415 2380
rect 2939 2063 2942 2096
rect 2942 2063 2988 2096
rect 2988 2063 2991 2096
rect 2939 2044 2991 2063
rect 3300 1971 3352 2023
rect 3512 1971 3564 2023
rect 1943 1767 1946 1781
rect 1946 1767 1992 1781
rect 1992 1767 1995 1781
rect 1943 1729 1995 1767
rect 1943 1560 1946 1595
rect 1946 1560 1992 1595
rect 1992 1560 1995 1595
rect 1943 1543 1995 1560
rect 1480 1147 1636 1154
rect 1480 1102 1502 1147
rect 1502 1102 1636 1147
rect -336 891 -284 908
rect -336 856 -333 891
rect -333 856 -287 891
rect -287 856 -284 891
rect -336 670 -333 722
rect -333 670 -287 722
rect -287 670 -284 722
rect 226 898 228 908
rect 228 898 274 908
rect 274 898 278 908
rect 226 856 278 898
rect 226 709 278 722
rect 226 670 228 709
rect 228 670 274 709
rect 274 670 278 709
rect 672 898 676 908
rect 676 898 722 908
rect 722 898 724 908
rect 672 856 724 898
rect 672 709 724 722
rect 672 670 676 709
rect 676 670 722 709
rect 722 670 724 709
rect 1122 898 1124 908
rect 1124 898 1170 908
rect 1170 898 1174 908
rect 1122 856 1174 898
rect 1122 709 1174 722
rect 1122 670 1124 709
rect 1124 670 1170 709
rect 1170 670 1174 709
rect 1551 805 1554 815
rect 1554 805 1600 815
rect 1600 805 1603 815
rect 1551 763 1603 805
rect 1551 603 1603 629
rect 1551 577 1554 603
rect 1554 577 1600 603
rect 1600 577 1603 603
rect 1943 799 1946 815
rect 1946 799 1992 815
rect 1992 799 1995 815
rect 1943 763 1995 799
rect 1943 599 1995 629
rect 1943 577 1946 599
rect 1946 577 1992 599
rect 1992 577 1995 599
rect 2638 1338 2690 1364
rect 2638 1312 2640 1338
rect 2640 1312 2686 1338
rect 2686 1312 2690 1338
rect 2638 1126 2690 1178
rect 1612 374 1768 376
rect 1612 328 1616 374
rect 1616 328 1756 374
rect 1756 328 1768 374
rect 1612 324 1768 328
rect 3097 1338 3149 1364
rect 3097 1312 3134 1338
rect 3134 1312 3149 1338
rect 3097 1126 3149 1178
rect 3545 1729 3597 1781
rect 3545 1593 3597 1595
rect 3545 1547 3558 1593
rect 3558 1547 3597 1593
rect 3545 1543 3597 1547
rect 4530 2246 4582 2282
rect 4530 2230 4533 2246
rect 4533 2230 4579 2246
rect 4579 2230 4582 2246
rect 4530 2094 4533 2096
rect 4533 2094 4579 2096
rect 4579 2094 4582 2096
rect 4530 2044 4582 2094
rect 4929 2230 4932 2282
rect 4932 2230 4978 2282
rect 4978 2230 4981 2282
rect 4929 2044 4932 2096
rect 4932 2044 4978 2096
rect 4978 2044 4981 2096
rect 4530 1776 4533 1781
rect 4533 1776 4579 1781
rect 4579 1776 4582 1781
rect 4530 1729 4582 1776
rect 4530 1564 4533 1595
rect 4533 1564 4579 1595
rect 4579 1564 4582 1595
rect 4530 1543 4582 1564
rect 4929 1729 4932 1781
rect 4932 1729 4978 1781
rect 4978 1729 4981 1781
rect 4929 1552 4932 1595
rect 4932 1552 4978 1595
rect 4978 1552 4981 1595
rect 4929 1543 4981 1552
rect 3963 1130 4119 1182
rect 4292 1136 4448 1139
rect 4292 1090 4303 1136
rect 4303 1090 4443 1136
rect 4443 1090 4448 1136
rect 4292 1087 4448 1090
rect 3567 866 3619 908
rect 3567 856 3604 866
rect 3604 856 3619 866
rect 3567 670 3619 722
rect 3469 441 3521 493
rect 3681 441 3733 493
rect 4575 898 4578 908
rect 4578 898 4624 908
rect 4624 898 4627 908
rect 4575 856 4627 898
rect 4575 696 4627 722
rect 4575 670 4578 696
rect 4578 670 4624 696
rect 4624 670 4627 696
rect 4929 -63 4981 -62
rect 4929 -114 4932 -63
rect 4932 -114 4978 -63
rect 4978 -114 4981 -63
rect 4929 -297 4932 -248
rect 4932 -297 4978 -248
rect 4978 -297 4981 -248
rect 4929 -300 4981 -297
<< metal2 >>
rect 3709 2790 3801 2830
rect 3709 2751 3729 2790
rect 2170 2729 2478 2747
rect 2170 2673 2198 2729
rect 2254 2673 2384 2729
rect 2440 2673 2478 2729
rect 2170 2655 2478 2673
rect 3708 2738 3729 2751
rect 3781 2751 3801 2790
rect 3781 2738 3802 2751
rect 3708 2604 3802 2738
rect 3918 2729 4226 2747
rect 3918 2673 3946 2729
rect 4002 2673 4132 2729
rect 4188 2673 4226 2729
rect 3918 2655 4226 2673
rect 3708 2552 3729 2604
rect 3781 2552 3802 2604
rect 3076 2415 3452 2438
rect 3076 2363 3363 2415
rect 3415 2363 3452 2415
rect 3076 2341 3452 2363
rect 2312 2284 2404 2312
rect 2312 2228 2330 2284
rect 2386 2228 2404 2284
rect 2312 2098 2404 2228
rect 2312 2042 2330 2098
rect 2386 2042 2404 2098
rect 2312 2004 2404 2042
rect 2761 2284 2853 2312
rect 2761 2228 2779 2284
rect 2835 2228 2853 2284
rect 2761 2098 2853 2228
rect 2761 2042 2779 2098
rect 2835 2042 2853 2098
rect 2761 2004 2853 2042
rect 2919 2284 3011 2312
rect 2919 2228 2937 2284
rect 2993 2228 3011 2284
rect 2919 2098 3011 2228
rect 2919 2042 2937 2098
rect 2993 2042 3011 2098
rect 2919 2004 3011 2042
rect -356 1783 -264 1811
rect -356 1727 -338 1783
rect -282 1727 -264 1783
rect -356 1597 -264 1727
rect -356 1541 -338 1597
rect -282 1541 -264 1597
rect -356 1503 -264 1541
rect 206 1783 298 1811
rect 206 1727 224 1783
rect 280 1727 298 1783
rect 206 1597 298 1727
rect 206 1541 224 1597
rect 280 1541 298 1597
rect 206 1503 298 1541
rect 652 1783 744 1811
rect 652 1727 670 1783
rect 726 1727 744 1783
rect 652 1597 744 1727
rect 652 1541 670 1597
rect 726 1541 744 1597
rect 652 1503 744 1541
rect 1100 1783 1192 1811
rect 1100 1727 1118 1783
rect 1174 1727 1192 1783
rect 1100 1597 1192 1727
rect 1100 1541 1118 1597
rect 1174 1541 1192 1597
rect 1100 1503 1192 1541
rect 1531 1783 1623 1811
rect 1531 1727 1549 1783
rect 1605 1727 1623 1783
rect 1531 1597 1623 1727
rect 1531 1541 1549 1597
rect 1605 1541 1623 1597
rect 1531 1503 1623 1541
rect 1923 1783 2015 1811
rect 1923 1727 1941 1783
rect 1997 1727 2015 1783
rect 1923 1597 2015 1727
rect 1923 1541 1941 1597
rect 1997 1541 2015 1597
rect 1923 1503 2015 1541
rect 2618 1366 2710 1394
rect 2618 1310 2636 1366
rect 2692 1310 2710 1366
rect 2618 1180 2710 1310
rect 1468 1165 1648 1166
rect 1468 1155 1671 1165
rect 1468 1154 1501 1155
rect 1468 1102 1480 1154
rect 1468 1099 1501 1102
rect 1661 1099 1671 1155
rect 1468 1090 1671 1099
rect 1491 1089 1671 1090
rect 2618 1124 2636 1180
rect 2692 1124 2710 1180
rect 2618 1086 2710 1124
rect 3076 1366 3170 2341
rect 3263 2023 3602 2064
rect 3263 1971 3300 2023
rect 3352 1971 3512 2023
rect 3564 1971 3602 2023
rect 3263 1930 3602 1971
rect 3076 1310 3095 1366
rect 3151 1310 3170 1366
rect 3076 1180 3170 1310
rect 3076 1124 3095 1180
rect 3151 1124 3170 1180
rect 3076 1103 3170 1124
rect 3077 1086 3169 1103
rect -356 910 -264 938
rect -356 854 -338 910
rect -282 854 -264 910
rect -356 724 -264 854
rect -356 668 -338 724
rect -282 668 -264 724
rect -356 630 -264 668
rect 206 910 298 938
rect 206 854 224 910
rect 280 854 298 910
rect 206 724 298 854
rect 206 668 224 724
rect 280 668 298 724
rect 206 630 298 668
rect 652 910 744 938
rect 652 854 670 910
rect 726 854 744 910
rect 652 724 744 854
rect 652 668 670 724
rect 726 668 744 724
rect 652 630 744 668
rect 1102 910 1194 938
rect 1102 854 1120 910
rect 1176 854 1194 910
rect 1102 724 1194 854
rect 1102 668 1120 724
rect 1176 668 1194 724
rect 1102 630 1194 668
rect 1531 817 1623 845
rect 1531 761 1549 817
rect 1605 761 1623 817
rect 1531 631 1623 761
rect 1531 575 1549 631
rect 1605 575 1623 631
rect 1531 537 1623 575
rect 1923 817 2015 845
rect 1923 761 1941 817
rect 1997 761 2015 817
rect 1923 631 2015 761
rect 1923 575 1941 631
rect 1997 575 2015 631
rect 1923 537 2015 575
rect 3344 534 3433 1930
rect 3525 1783 3617 1811
rect 3525 1727 3543 1783
rect 3599 1727 3617 1783
rect 3525 1597 3617 1727
rect 3525 1541 3543 1597
rect 3599 1541 3617 1597
rect 3525 1503 3617 1541
rect 3708 1060 3802 2552
rect 3951 1184 4131 1194
rect 3951 1128 3961 1184
rect 4121 1128 4131 1184
rect 4324 1151 4418 2751
rect 4510 2284 4602 2312
rect 4510 2228 4528 2284
rect 4584 2228 4602 2284
rect 4510 2098 4602 2228
rect 4510 2042 4528 2098
rect 4584 2042 4602 2098
rect 4510 2004 4602 2042
rect 4909 2284 5001 2312
rect 4909 2228 4927 2284
rect 4983 2228 5001 2284
rect 4909 2098 5001 2228
rect 4909 2042 4927 2098
rect 4983 2042 5001 2098
rect 4909 2004 5001 2042
rect 4510 1783 4602 1811
rect 4510 1727 4528 1783
rect 4584 1727 4602 1783
rect 4510 1597 4602 1727
rect 4510 1541 4528 1597
rect 4584 1541 4602 1597
rect 4510 1503 4602 1541
rect 4909 1783 5001 1811
rect 4909 1727 4927 1783
rect 4983 1727 5001 1783
rect 4909 1597 5001 1727
rect 4909 1541 4927 1597
rect 4983 1541 5001 1597
rect 4909 1503 5001 1541
rect 3951 1118 4131 1128
rect 4280 1139 4460 1151
rect 4280 1087 4292 1139
rect 4448 1087 4460 1139
rect 4280 1075 4460 1087
rect 3547 910 3639 938
rect 3547 854 3565 910
rect 3621 854 3639 910
rect 3547 724 3639 854
rect 3547 668 3565 724
rect 3621 668 3639 724
rect 3547 630 3639 668
rect 4555 910 4647 938
rect 4555 854 4573 910
rect 4629 854 4647 910
rect 4555 724 4647 854
rect 4555 668 4573 724
rect 4629 668 4647 724
rect 4555 630 4647 668
rect 3344 493 3771 534
rect 3344 441 3469 493
rect 3521 441 3681 493
rect 3733 441 3771 493
rect 3344 400 3771 441
rect 1600 376 1780 388
rect 1600 324 1612 376
rect 1768 324 1780 376
rect 1600 312 1780 324
rect 4909 -60 5001 -32
rect 4909 -116 4927 -60
rect 4983 -116 5001 -60
rect 4909 -246 5001 -116
rect 4909 -302 4927 -246
rect 4983 -302 5001 -246
rect 4909 -340 5001 -302
<< via2 >>
rect 2198 2727 2254 2729
rect 2198 2675 2200 2727
rect 2200 2675 2252 2727
rect 2252 2675 2254 2727
rect 2198 2673 2254 2675
rect 2384 2727 2440 2729
rect 2384 2675 2386 2727
rect 2386 2675 2438 2727
rect 2438 2675 2440 2727
rect 2384 2673 2440 2675
rect 3946 2727 4002 2729
rect 3946 2675 3948 2727
rect 3948 2675 4000 2727
rect 4000 2675 4002 2727
rect 3946 2673 4002 2675
rect 4132 2727 4188 2729
rect 4132 2675 4134 2727
rect 4134 2675 4186 2727
rect 4186 2675 4188 2727
rect 4132 2673 4188 2675
rect 2330 2282 2386 2284
rect 2330 2230 2332 2282
rect 2332 2230 2384 2282
rect 2384 2230 2386 2282
rect 2330 2228 2386 2230
rect 2330 2096 2386 2098
rect 2330 2044 2332 2096
rect 2332 2044 2384 2096
rect 2384 2044 2386 2096
rect 2330 2042 2386 2044
rect 2779 2282 2835 2284
rect 2779 2230 2781 2282
rect 2781 2230 2833 2282
rect 2833 2230 2835 2282
rect 2779 2228 2835 2230
rect 2779 2096 2835 2098
rect 2779 2044 2781 2096
rect 2781 2044 2833 2096
rect 2833 2044 2835 2096
rect 2779 2042 2835 2044
rect 2937 2282 2993 2284
rect 2937 2230 2939 2282
rect 2939 2230 2991 2282
rect 2991 2230 2993 2282
rect 2937 2228 2993 2230
rect 2937 2096 2993 2098
rect 2937 2044 2939 2096
rect 2939 2044 2991 2096
rect 2991 2044 2993 2096
rect 2937 2042 2993 2044
rect -338 1781 -282 1783
rect -338 1729 -336 1781
rect -336 1729 -284 1781
rect -284 1729 -282 1781
rect -338 1727 -282 1729
rect -338 1595 -282 1597
rect -338 1543 -336 1595
rect -336 1543 -284 1595
rect -284 1543 -282 1595
rect -338 1541 -282 1543
rect 224 1781 280 1783
rect 224 1729 226 1781
rect 226 1729 278 1781
rect 278 1729 280 1781
rect 224 1727 280 1729
rect 224 1595 280 1597
rect 224 1543 226 1595
rect 226 1543 278 1595
rect 278 1543 280 1595
rect 224 1541 280 1543
rect 670 1781 726 1783
rect 670 1729 672 1781
rect 672 1729 724 1781
rect 724 1729 726 1781
rect 670 1727 726 1729
rect 670 1595 726 1597
rect 670 1543 672 1595
rect 672 1543 724 1595
rect 724 1543 726 1595
rect 670 1541 726 1543
rect 1118 1781 1174 1783
rect 1118 1729 1120 1781
rect 1120 1729 1172 1781
rect 1172 1729 1174 1781
rect 1118 1727 1174 1729
rect 1118 1595 1174 1597
rect 1118 1543 1120 1595
rect 1120 1543 1172 1595
rect 1172 1543 1174 1595
rect 1118 1541 1174 1543
rect 1549 1781 1605 1783
rect 1549 1729 1551 1781
rect 1551 1729 1603 1781
rect 1603 1729 1605 1781
rect 1549 1727 1605 1729
rect 1549 1595 1605 1597
rect 1549 1543 1551 1595
rect 1551 1543 1603 1595
rect 1603 1543 1605 1595
rect 1549 1541 1605 1543
rect 1941 1781 1997 1783
rect 1941 1729 1943 1781
rect 1943 1729 1995 1781
rect 1995 1729 1997 1781
rect 1941 1727 1997 1729
rect 1941 1595 1997 1597
rect 1941 1543 1943 1595
rect 1943 1543 1995 1595
rect 1995 1543 1997 1595
rect 1941 1541 1997 1543
rect 2636 1364 2692 1366
rect 2636 1312 2638 1364
rect 2638 1312 2690 1364
rect 2690 1312 2692 1364
rect 2636 1310 2692 1312
rect 1501 1154 1661 1155
rect 1501 1102 1636 1154
rect 1636 1102 1661 1154
rect 1501 1099 1661 1102
rect 2636 1178 2692 1180
rect 2636 1126 2638 1178
rect 2638 1126 2690 1178
rect 2690 1126 2692 1178
rect 2636 1124 2692 1126
rect 3095 1364 3151 1366
rect 3095 1312 3097 1364
rect 3097 1312 3149 1364
rect 3149 1312 3151 1364
rect 3095 1310 3151 1312
rect 3095 1178 3151 1180
rect 3095 1126 3097 1178
rect 3097 1126 3149 1178
rect 3149 1126 3151 1178
rect 3095 1124 3151 1126
rect -338 908 -282 910
rect -338 856 -336 908
rect -336 856 -284 908
rect -284 856 -282 908
rect -338 854 -282 856
rect -338 722 -282 724
rect -338 670 -336 722
rect -336 670 -284 722
rect -284 670 -282 722
rect -338 668 -282 670
rect 224 908 280 910
rect 224 856 226 908
rect 226 856 278 908
rect 278 856 280 908
rect 224 854 280 856
rect 224 722 280 724
rect 224 670 226 722
rect 226 670 278 722
rect 278 670 280 722
rect 224 668 280 670
rect 670 908 726 910
rect 670 856 672 908
rect 672 856 724 908
rect 724 856 726 908
rect 670 854 726 856
rect 670 722 726 724
rect 670 670 672 722
rect 672 670 724 722
rect 724 670 726 722
rect 670 668 726 670
rect 1120 908 1176 910
rect 1120 856 1122 908
rect 1122 856 1174 908
rect 1174 856 1176 908
rect 1120 854 1176 856
rect 1120 722 1176 724
rect 1120 670 1122 722
rect 1122 670 1174 722
rect 1174 670 1176 722
rect 1120 668 1176 670
rect 1549 815 1605 817
rect 1549 763 1551 815
rect 1551 763 1603 815
rect 1603 763 1605 815
rect 1549 761 1605 763
rect 1549 629 1605 631
rect 1549 577 1551 629
rect 1551 577 1603 629
rect 1603 577 1605 629
rect 1549 575 1605 577
rect 1941 815 1997 817
rect 1941 763 1943 815
rect 1943 763 1995 815
rect 1995 763 1997 815
rect 1941 761 1997 763
rect 1941 629 1997 631
rect 1941 577 1943 629
rect 1943 577 1995 629
rect 1995 577 1997 629
rect 1941 575 1997 577
rect 3543 1781 3599 1783
rect 3543 1729 3545 1781
rect 3545 1729 3597 1781
rect 3597 1729 3599 1781
rect 3543 1727 3599 1729
rect 3543 1595 3599 1597
rect 3543 1543 3545 1595
rect 3545 1543 3597 1595
rect 3597 1543 3599 1595
rect 3543 1541 3599 1543
rect 3961 1182 4121 1184
rect 3961 1130 3963 1182
rect 3963 1130 4119 1182
rect 4119 1130 4121 1182
rect 3961 1128 4121 1130
rect 4528 2282 4584 2284
rect 4528 2230 4530 2282
rect 4530 2230 4582 2282
rect 4582 2230 4584 2282
rect 4528 2228 4584 2230
rect 4528 2096 4584 2098
rect 4528 2044 4530 2096
rect 4530 2044 4582 2096
rect 4582 2044 4584 2096
rect 4528 2042 4584 2044
rect 4927 2282 4983 2284
rect 4927 2230 4929 2282
rect 4929 2230 4981 2282
rect 4981 2230 4983 2282
rect 4927 2228 4983 2230
rect 4927 2096 4983 2098
rect 4927 2044 4929 2096
rect 4929 2044 4981 2096
rect 4981 2044 4983 2096
rect 4927 2042 4983 2044
rect 4528 1781 4584 1783
rect 4528 1729 4530 1781
rect 4530 1729 4582 1781
rect 4582 1729 4584 1781
rect 4528 1727 4584 1729
rect 4528 1595 4584 1597
rect 4528 1543 4530 1595
rect 4530 1543 4582 1595
rect 4582 1543 4584 1595
rect 4528 1541 4584 1543
rect 4927 1781 4983 1783
rect 4927 1729 4929 1781
rect 4929 1729 4981 1781
rect 4981 1729 4983 1781
rect 4927 1727 4983 1729
rect 4927 1595 4983 1597
rect 4927 1543 4929 1595
rect 4929 1543 4981 1595
rect 4981 1543 4983 1595
rect 4927 1541 4983 1543
rect 3565 908 3621 910
rect 3565 856 3567 908
rect 3567 856 3619 908
rect 3619 856 3621 908
rect 3565 854 3621 856
rect 3565 722 3621 724
rect 3565 670 3567 722
rect 3567 670 3619 722
rect 3619 670 3621 722
rect 3565 668 3621 670
rect 4573 908 4629 910
rect 4573 856 4575 908
rect 4575 856 4627 908
rect 4627 856 4629 908
rect 4573 854 4629 856
rect 4573 722 4629 724
rect 4573 670 4575 722
rect 4575 670 4627 722
rect 4627 670 4629 722
rect 4573 668 4629 670
rect 4927 -62 4983 -60
rect 4927 -114 4929 -62
rect 4929 -114 4981 -62
rect 4981 -114 4983 -62
rect 4927 -116 4983 -114
rect 4927 -248 4983 -246
rect 4927 -300 4929 -248
rect 4929 -300 4981 -248
rect 4981 -300 4983 -248
rect 4927 -302 4983 -300
<< metal3 >>
rect 2113 2729 4296 2748
rect 2113 2673 2198 2729
rect 2254 2673 2384 2729
rect 2440 2673 3946 2729
rect 4002 2673 4132 2729
rect 4188 2673 4296 2729
rect 2113 2655 4296 2673
rect -356 2284 5006 2312
rect -356 2228 2330 2284
rect 2386 2228 2779 2284
rect 2835 2228 2937 2284
rect 2993 2228 4528 2284
rect 4584 2228 4927 2284
rect 4983 2228 5006 2284
rect -356 2098 5006 2228
rect -356 2042 2330 2098
rect 2386 2042 2779 2098
rect 2835 2042 2937 2098
rect 2993 2042 4528 2098
rect 4584 2042 4927 2098
rect 4983 2042 5006 2098
rect -356 1783 5006 2042
rect -356 1727 -338 1783
rect -282 1727 224 1783
rect 280 1727 670 1783
rect 726 1727 1118 1783
rect 1174 1727 1549 1783
rect 1605 1727 1941 1783
rect 1997 1727 3543 1783
rect 3599 1727 4528 1783
rect 4584 1727 4927 1783
rect 4983 1727 5006 1783
rect -356 1597 5006 1727
rect -356 1541 -338 1597
rect -282 1541 224 1597
rect 280 1541 670 1597
rect 726 1541 1118 1597
rect 1174 1541 1549 1597
rect 1605 1541 1941 1597
rect 1997 1541 3543 1597
rect 3599 1541 4528 1597
rect 4584 1541 4927 1597
rect 4983 1541 5006 1597
rect -356 1502 5006 1541
rect 2617 1366 2710 1394
rect 2617 1310 2636 1366
rect 2692 1310 2710 1366
rect 2617 1203 2710 1310
rect 3076 1366 3169 1394
rect 3076 1310 3095 1366
rect 3151 1310 3169 1366
rect 3076 1203 3169 1310
rect 1491 1184 4131 1203
rect 1491 1180 3961 1184
rect 1491 1155 2636 1180
rect 1491 1099 1501 1155
rect 1661 1124 2636 1155
rect 2692 1124 3095 1180
rect 3151 1128 3961 1180
rect 4121 1128 4131 1184
rect 3151 1124 4131 1128
rect 1661 1106 4131 1124
rect 1661 1099 1671 1106
rect 1491 1089 1671 1099
rect 2617 1085 2710 1106
rect 3076 1085 3169 1106
rect -356 910 5028 957
rect -356 854 -338 910
rect -282 854 224 910
rect 280 854 670 910
rect 726 854 1120 910
rect 1176 854 3565 910
rect 3621 854 4573 910
rect 4629 854 5028 910
rect -356 817 5028 854
rect -356 761 1549 817
rect 1605 761 1941 817
rect 1997 761 5028 817
rect -356 724 5028 761
rect -356 668 -338 724
rect -282 668 224 724
rect 280 668 670 724
rect 726 668 1120 724
rect 1176 668 3565 724
rect 3621 668 4573 724
rect 4629 668 5028 724
rect -356 631 5028 668
rect -356 575 1549 631
rect 1605 575 1941 631
rect 1997 575 5028 631
rect -356 169 5028 575
rect -357 -60 5028 169
rect -357 -116 4927 -60
rect 4983 -116 5028 -60
rect -357 -246 5028 -116
rect -357 -302 4927 -246
rect 4983 -302 5028 -246
rect -357 -359 5028 -302
use M1_NACTIVE4310591302038_512x8m81  M1_NACTIVE4310591302038_512x8m81_0
timestamp 1698431365
transform 1 0 4955 0 1 1951
box 0 0 1 1
use M1_NACTIVE4310591302041_512x8m81  M1_NACTIVE4310591302041_512x8m81_0
timestamp 1698431365
transform 1 0 478 0 1 2177
box 0 0 1 1
use M1_NWELL_01_R270_512x8m81  M1_NWELL_01_R270_512x8m81_0
timestamp 1698431365
transform 0 1 -310 -1 0 1587
box 0 0 1 1
use M1_PACTIVE4310591302034_512x8m81  M1_PACTIVE4310591302034_512x8m81_0
timestamp 1698431365
transform 1 0 -310 0 1 727
box 0 0 1 1
use M1_PACTIVE4310591302039_512x8m81  M1_PACTIVE4310591302039_512x8m81_0
timestamp 1698431365
transform 1 0 4955 0 1 -180
box 0 0 1 1
use M1_PACTIVE4310591302040_512x8m81  M1_PACTIVE4310591302040_512x8m81_0
timestamp 1698431365
transform 1 0 683 0 1 338
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_0
timestamp 1698431365
transform 0 -1 1479 1 0 1124
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_1
timestamp 1698431365
transform 1 0 3546 0 1 469
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_2
timestamp 1698431365
transform 1 0 2701 0 1 2442
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_3
timestamp 1698431365
transform 1 0 3380 0 1 2403
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_4
timestamp 1698431365
transform 1 0 3112 0 1 1835
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_5
timestamp 1698431365
transform 1 0 3467 0 1 1975
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_6
timestamp 1698431365
transform 1 0 3756 0 1 2578
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_7
timestamp 1698431365
transform 1 0 3282 0 1 465
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_0
timestamp 1698431365
transform -1 0 2125 0 -1 438
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_1
timestamp 1698431365
transform -1 0 1942 0 -1 1082
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_2
timestamp 1698431365
transform 1 0 4119 0 -1 2699
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_3
timestamp 1698431365
transform 1 0 4595 0 1 174
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_4
timestamp 1698431365
transform 1 0 1686 0 1 351
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_5
timestamp 1698431365
transform 1 0 4373 0 1 1113
box 0 0 1 1
use M1_PSUB_02_512x8m81  M1_PSUB_02_512x8m81_0
timestamp 1698431365
transform 1 0 3518 0 1 2677
box 0 0 1 1
use M2_M1$$168351788_R90_512x8m81  M2_M1$$168351788_R90_512x8m81_0
timestamp 1698431365
transform 0 -1 3601 1 0 467
box 0 0 1 1
use M2_M1$$168351788_R90_512x8m81  M2_M1$$168351788_R90_512x8m81_1
timestamp 1698431365
transform 0 -1 3432 1 0 1997
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_0
timestamp 1698431365
transform 1 0 1690 0 1 350
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_1
timestamp 1698431365
transform 1 0 1558 0 1 1128
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_2
timestamp 1698431365
transform 1 0 4041 0 1 1156
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_3
timestamp 1698431365
transform 1 0 4370 0 1 1113
box 0 0 1 1
use M3_M2431059130207_512x8m81  M3_M2431059130207_512x8m81_0
timestamp 1698431365
transform 1 0 4041 0 1 1156
box 0 0 1 1
use M3_M2431059130207_512x8m81  M3_M2431059130207_512x8m81_1
timestamp 1698431365
transform 1 0 1581 0 1 1127
box 0 0 1 1
use nmos_5p0431059130208_512x8m81  nmos_5p0431059130208_512x8m81_0
timestamp 1698431365
transform -1 0 3529 0 1 807
box 0 0 1 1
use nmos_5p0431059130208_512x8m81  nmos_5p0431059130208_512x8m81_1
timestamp 1698431365
transform 1 0 2635 0 -1 2761
box 0 0 1 1
use nmos_5p04310591302033_512x8m81  nmos_5p04310591302033_512x8m81_0
timestamp 1698431365
transform 1 0 3030 0 -1 2673
box 0 0 1 1
use nmos_5p04310591302044_512x8m81  nmos_5p04310591302044_512x8m81_0
timestamp 1698431365
transform -1 0 2141 0 1 540
box 0 0 1 1
use nmos_5p04310591302045_512x8m81  nmos_5p04310591302045_512x8m81_0
timestamp 1698431365
transform 1 0 4429 0 -1 957
box 0 0 1 1
use nmos_5p04310591302045_512x8m81  nmos_5p04310591302045_512x8m81_1
timestamp 1698431365
transform 1 0 3981 0 -1 957
box 0 0 1 1
use nmos_5p04310591302046_512x8m81  nmos_5p04310591302046_512x8m81_0
timestamp 1698431365
transform -1 0 1319 0 -1 957
box 0 0 1 1
use nmos_5p04310591302050_512x8m81  nmos_5p04310591302050_512x8m81_0
timestamp 1698431365
transform -1 0 3059 0 1 544
box 0 0 1 1
use nmos_5p04310591302052_512x8m81  nmos_5p04310591302052_512x8m81_0
timestamp 1698431365
transform -1 0 1749 0 1 544
box 0 0 1 1
use pmos_1p2$$171625516_512x8m81  pmos_1p2$$171625516_512x8m81_0
timestamp 1698431365
transform 1 0 2442 0 -1 2290
box -31 0 -30 1
use pmos_5p04310591302013_512x8m81  pmos_5p04310591302013_512x8m81_0
timestamp 1698431365
transform -1 0 3059 0 1 1279
box 0 0 1 1
use pmos_5p04310591302014_512x8m81  pmos_5p04310591302014_512x8m81_0
timestamp 1698431365
transform -1 0 3529 0 1 1406
box 0 0 1 1
use pmos_5p04310591302038_512x8m81  pmos_5p04310591302038_512x8m81_0
timestamp 1698431365
transform 1 0 3017 0 -1 2290
box 0 0 1 1
use pmos_5p04310591302047_512x8m81  pmos_5p04310591302047_512x8m81_0
timestamp 1698431365
transform -1 0 1749 0 1 1279
box 0 0 1 1
use pmos_5p04310591302048_512x8m81  pmos_5p04310591302048_512x8m81_0
timestamp 1698431365
transform -1 0 2141 0 1 1235
box 0 0 1 1
use pmos_5p04310591302049_512x8m81  pmos_5p04310591302049_512x8m81_0
timestamp 1698431365
transform -1 0 1319 0 1 1238
box 0 0 1 1
use pmos_5p04310591302051_512x8m81  pmos_5p04310591302051_512x8m81_0
timestamp 1698431365
transform 1 0 3936 0 1 1337
box 0 0 1 1
use pmos_5p04310591302051_512x8m81  pmos_5p04310591302051_512x8m81_1
timestamp 1698431365
transform 1 0 4384 0 1 1337
box 0 0 1 1
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_0
timestamp 1698431365
transform -1 0 3169 0 1 1086
box 0 0 1 1
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_1
timestamp 1698431365
transform -1 0 2710 0 1 1086
box 0 0 1 1
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_2
timestamp 1698431365
transform 0 -1 4226 1 0 2655
box 0 0 1 1
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_3
timestamp 1698431365
transform 0 -1 2478 1 0 2655
box 0 0 1 1
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_4
timestamp 1698431365
transform 1 0 4909 0 1 -340
box 0 0 1 1
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_5
timestamp 1698431365
transform 1 0 206 0 1 1503
box 0 0 1 1
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_6
timestamp 1698431365
transform 1 0 652 0 1 1503
box 0 0 1 1
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_7
timestamp 1698431365
transform 1 0 1100 0 1 1503
box 0 0 1 1
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_8
timestamp 1698431365
transform 1 0 652 0 1 630
box 0 0 1 1
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_9
timestamp 1698431365
transform 1 0 206 0 1 630
box 0 0 1 1
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_10
timestamp 1698431365
transform 1 0 4510 0 1 1503
box 0 0 1 1
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_11
timestamp 1698431365
transform 1 0 4510 0 1 2004
box 0 0 1 1
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_12
timestamp 1698431365
transform 1 0 4555 0 1 630
box 0 0 1 1
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_13
timestamp 1698431365
transform 1 0 3525 0 1 1503
box 0 0 1 1
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_14
timestamp 1698431365
transform 1 0 3547 0 1 630
box 0 0 1 1
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_15
timestamp 1698431365
transform 1 0 1102 0 1 630
box 0 0 1 1
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_16
timestamp 1698431365
transform 1 0 2761 0 1 2004
box 0 0 1 1
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_17
timestamp 1698431365
transform 1 0 2312 0 1 2004
box 0 0 1 1
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_18
timestamp 1698431365
transform 1 0 -356 0 1 1503
box 0 0 1 1
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_19
timestamp 1698431365
transform 1 0 -356 0 1 630
box 0 0 1 1
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_20
timestamp 1698431365
transform 1 0 4909 0 1 1503
box 0 0 1 1
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_21
timestamp 1698431365
transform 1 0 4909 0 1 2004
box 0 0 1 1
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_22
timestamp 1698431365
transform 1 0 1531 0 1 1503
box 0 0 1 1
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_23
timestamp 1698431365
transform 1 0 1923 0 1 1503
box 0 0 1 1
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_24
timestamp 1698431365
transform 1 0 1531 0 1 537
box 0 0 1 1
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_25
timestamp 1698431365
transform 1 0 1923 0 1 537
box 0 0 1 1
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_26
timestamp 1698431365
transform 1 0 2919 0 1 2004
box 0 0 1 1
use via1_R270_512x8m81  via1_R270_512x8m81_0
timestamp 1698431365
transform 0 1 3325 -1 0 2437
box 0 0 1 1
use via1_x2_512x8m81  via1_x2_512x8m81_0
timestamp 1698431365
transform -1 0 3801 0 1 2512
box 0 0 1 1
<< labels >>
rlabel metal3 s -214 644 -214 644 4 vss
port 1 nsew
rlabel metal3 s -255 2131 -255 2131 4 vdd
port 2 nsew
rlabel metal2 s 3762 2693 3762 2693 4 qp
port 3 nsew
rlabel metal2 s 4401 2693 4401 2693 4 qn
port 4 nsew
rlabel metal1 s 3628 469 3628 469 4 se
port 5 nsew
rlabel metal1 s 467 1145 467 1145 4 q
port 6 nsew
rlabel metal1 s 3511 2689 3511 2689 4 vss
port 1 nsew
rlabel metal1 s 1613 361 1613 361 4 GWE
port 7 nsew
<< properties >>
string GDS_END 421608
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 410634
string path 21.660 12.815 21.660 12.970 
<< end >>
