magic
tech gf180mcuD
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 352 1654 870
<< pwell >>
rect -86 -86 1654 352
<< metal1 >>
rect 0 724 1568 844
rect 132 203 204 458
rect 356 296 428 678
rect 580 296 652 678
rect 804 296 876 678
rect 964 506 1010 724
rect 1194 536 1317 678
rect 1409 598 1455 724
rect 1194 472 1456 536
rect 1402 312 1456 472
rect 1205 248 1456 312
rect 38 60 106 131
rect 486 60 554 131
rect 934 60 1002 131
rect 1205 106 1317 248
rect 1429 60 1475 180
rect 0 -60 1568 60
<< obsm1 >>
rect 69 552 115 678
rect 69 506 308 552
rect 262 236 308 506
rect 1006 369 1350 415
rect 1006 236 1052 369
rect 262 189 1052 236
rect 262 106 330 189
rect 710 106 778 189
<< labels >>
rlabel metal1 s 132 203 204 458 6 A1
port 1 nsew default input
rlabel metal1 s 356 296 428 678 6 A2
port 2 nsew default input
rlabel metal1 s 580 296 652 678 6 A3
port 3 nsew default input
rlabel metal1 s 804 296 876 678 6 A4
port 4 nsew default input
rlabel metal1 s 1205 106 1317 248 6 Z
port 5 nsew default output
rlabel metal1 s 1205 248 1456 312 6 Z
port 5 nsew default output
rlabel metal1 s 1402 312 1456 472 6 Z
port 5 nsew default output
rlabel metal1 s 1194 472 1456 536 6 Z
port 5 nsew default output
rlabel metal1 s 1194 536 1317 678 6 Z
port 5 nsew default output
rlabel metal1 s 1409 598 1455 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 964 506 1010 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 724 1568 844 6 VDD
port 6 nsew power bidirectional abutment
rlabel nwell s -86 352 1654 870 6 VNW
port 7 nsew power bidirectional
rlabel pwell s -86 -86 1654 352 6 VPW
port 8 nsew ground bidirectional
rlabel metal1 s 0 -60 1568 60 8 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1429 60 1475 180 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 934 60 1002 131 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 486 60 554 131 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 38 60 106 131 6 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1568 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 175942
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 171784
<< end >>
