magic
tech gf180mcuC
timestamp 1698431365
<< properties >>
string GDS_END 7034088
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 7031972
<< end >>
