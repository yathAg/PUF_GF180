magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 377 3558 870
rect -86 352 973 377
rect 1224 352 3558 377
<< pwell >>
rect 973 352 1224 377
rect -86 -86 3558 352
<< mvnmos >>
rect 124 151 244 232
rect 348 151 468 232
rect 716 159 836 231
rect 884 159 1004 231
rect 1208 159 1328 231
rect 1376 159 1496 231
rect 1688 159 1808 231
rect 1912 159 2032 231
rect 2136 159 2256 231
rect 2304 159 2424 231
rect 2572 151 2692 231
rect 2960 68 3080 232
rect 3184 68 3304 232
<< mvpmos >>
rect 144 472 244 645
rect 348 472 448 645
rect 780 527 880 599
rect 940 527 1040 599
rect 1248 527 1348 599
rect 1396 527 1496 599
rect 1612 527 1712 599
rect 1911 527 2011 599
rect 2196 527 2296 599
rect 2352 527 2452 599
rect 2600 527 2700 687
rect 2948 472 3048 716
rect 3152 472 3252 716
<< mvndiff >>
rect 36 219 124 232
rect 36 173 49 219
rect 95 173 124 219
rect 36 151 124 173
rect 244 210 348 232
rect 244 164 273 210
rect 319 164 348 210
rect 244 151 348 164
rect 468 219 556 232
rect 1064 244 1136 257
rect 1064 231 1077 244
rect 468 173 497 219
rect 543 173 556 219
rect 468 151 556 173
rect 628 218 716 231
rect 628 172 641 218
rect 687 172 716 218
rect 628 159 716 172
rect 836 159 884 231
rect 1004 198 1077 231
rect 1123 231 1136 244
rect 1123 198 1208 231
rect 1004 159 1208 198
rect 1328 159 1376 231
rect 1496 159 1688 231
rect 1808 218 1912 231
rect 1808 172 1837 218
rect 1883 172 1912 218
rect 1808 159 1912 172
rect 2032 218 2136 231
rect 2032 172 2061 218
rect 2107 172 2136 218
rect 2032 159 2136 172
rect 2256 159 2304 231
rect 2424 210 2572 231
rect 2424 164 2497 210
rect 2543 164 2572 210
rect 2424 159 2572 164
rect 1556 117 1628 159
rect 1556 71 1569 117
rect 1615 71 1628 117
rect 2484 151 2572 159
rect 2692 218 2780 231
rect 2692 172 2721 218
rect 2767 172 2780 218
rect 2692 151 2780 172
rect 2872 167 2960 232
rect 1556 58 1628 71
rect 2872 121 2885 167
rect 2931 121 2960 167
rect 2872 68 2960 121
rect 3080 167 3184 232
rect 3080 121 3109 167
rect 3155 121 3184 167
rect 3080 68 3184 121
rect 3304 167 3392 232
rect 3304 121 3333 167
rect 3379 121 3392 167
rect 3304 68 3392 121
<< mvpdiff >>
rect 648 694 720 720
rect 648 648 661 694
rect 707 648 720 694
rect 56 619 144 645
rect 56 573 69 619
rect 115 573 144 619
rect 56 472 144 573
rect 244 632 348 645
rect 244 586 273 632
rect 319 586 348 632
rect 244 472 348 586
rect 448 531 536 645
rect 448 485 477 531
rect 523 485 536 531
rect 648 599 720 648
rect 2860 689 2948 716
rect 2512 599 2600 687
rect 648 527 780 599
rect 880 527 940 599
rect 1040 586 1248 599
rect 1040 540 1133 586
rect 1179 540 1248 586
rect 1040 527 1248 540
rect 1348 527 1396 599
rect 1496 586 1612 599
rect 1496 540 1537 586
rect 1583 540 1612 586
rect 1496 527 1612 540
rect 1712 586 1911 599
rect 1712 540 1836 586
rect 1882 540 1911 586
rect 1712 527 1911 540
rect 2011 586 2196 599
rect 2011 540 2061 586
rect 2107 540 2196 586
rect 2011 527 2196 540
rect 2296 527 2352 599
rect 2452 595 2600 599
rect 2452 549 2525 595
rect 2571 549 2600 595
rect 2452 527 2600 549
rect 2700 595 2788 687
rect 2700 549 2729 595
rect 2775 549 2788 595
rect 2700 527 2788 549
rect 2860 549 2873 689
rect 2919 549 2948 689
rect 448 472 536 485
rect 2860 472 2948 549
rect 3048 595 3152 716
rect 3048 549 3077 595
rect 3123 549 3152 595
rect 3048 472 3152 549
rect 3252 689 3392 716
rect 3252 549 3333 689
rect 3379 549 3392 689
rect 3252 472 3392 549
<< mvndiffc >>
rect 49 173 95 219
rect 273 164 319 210
rect 497 173 543 219
rect 641 172 687 218
rect 1077 198 1123 244
rect 1837 172 1883 218
rect 2061 172 2107 218
rect 2497 164 2543 210
rect 1569 71 1615 117
rect 2721 172 2767 218
rect 2885 121 2931 167
rect 3109 121 3155 167
rect 3333 121 3379 167
<< mvpdiffc >>
rect 661 648 707 694
rect 69 573 115 619
rect 273 586 319 632
rect 477 485 523 531
rect 1133 540 1179 586
rect 1537 540 1583 586
rect 1836 540 1882 586
rect 2061 540 2107 586
rect 2525 549 2571 595
rect 2729 549 2775 595
rect 2873 549 2919 689
rect 3077 549 3123 595
rect 3333 549 3379 689
<< polysilicon >>
rect 1248 720 2011 760
rect 144 645 244 690
rect 348 645 448 690
rect 1248 678 1348 720
rect 780 599 880 672
rect 940 599 1040 672
rect 1248 632 1261 678
rect 1307 632 1348 678
rect 1248 599 1348 632
rect 1396 599 1496 672
rect 1612 599 1712 672
rect 1911 599 2011 720
rect 2196 678 2296 691
rect 2600 687 2700 760
rect 2948 716 3048 760
rect 3152 716 3252 760
rect 2196 632 2209 678
rect 2255 632 2296 678
rect 2196 599 2296 632
rect 2352 599 2452 643
rect 144 416 244 472
rect 144 370 157 416
rect 203 370 244 416
rect 144 288 244 370
rect 124 232 244 288
rect 348 332 448 472
rect 780 467 880 527
rect 756 454 880 467
rect 756 408 769 454
rect 815 408 880 454
rect 756 395 880 408
rect 348 313 836 332
rect 940 324 1040 527
rect 1248 471 1348 527
rect 348 267 383 313
rect 429 292 836 313
rect 429 267 468 292
rect 348 232 468 267
rect 716 231 836 292
rect 884 317 1040 324
rect 884 311 1004 317
rect 884 265 926 311
rect 972 265 1004 311
rect 884 231 1004 265
rect 1208 311 1328 324
rect 1208 265 1233 311
rect 1279 265 1328 311
rect 1396 310 1496 527
rect 1612 494 1712 527
rect 1612 448 1625 494
rect 1671 448 1712 494
rect 1612 396 1712 448
rect 1911 412 2011 527
rect 2196 483 2296 527
rect 2352 416 2452 527
rect 2600 425 2700 527
rect 2948 428 3048 472
rect 1612 356 1808 396
rect 1911 372 2176 412
rect 1396 275 1437 310
rect 1208 231 1328 265
rect 1376 264 1437 275
rect 1483 264 1496 310
rect 1376 231 1496 264
rect 1688 231 1808 356
rect 1912 310 2032 323
rect 1912 264 1944 310
rect 1990 264 2032 310
rect 1912 231 2032 264
rect 2136 275 2176 372
rect 2352 326 2424 416
rect 2352 280 2365 326
rect 2411 280 2424 326
rect 2600 379 2613 425
rect 2659 379 2700 425
rect 2600 311 2700 379
rect 2960 370 3048 428
rect 3152 370 3252 472
rect 2960 357 3252 370
rect 2960 311 2973 357
rect 3113 311 3304 357
rect 2600 288 2692 311
rect 2352 275 2424 280
rect 2136 231 2256 275
rect 2304 231 2424 275
rect 2572 231 2692 288
rect 2960 298 3304 311
rect 2960 232 3080 298
rect 3184 232 3304 298
rect 124 107 244 151
rect 348 107 468 151
rect 716 115 836 159
rect 884 115 1004 159
rect 1208 115 1328 159
rect 1376 115 1496 159
rect 1688 115 1808 159
rect 1912 115 2032 159
rect 2136 115 2256 159
rect 2304 115 2424 159
rect 2572 24 2692 151
rect 2960 24 3080 68
rect 3184 24 3304 68
<< polycontact >>
rect 1261 632 1307 678
rect 2209 632 2255 678
rect 157 370 203 416
rect 769 408 815 454
rect 383 267 429 313
rect 926 265 972 311
rect 1233 265 1279 311
rect 1625 448 1671 494
rect 1437 264 1483 310
rect 1944 264 1990 310
rect 2365 280 2411 326
rect 2613 379 2659 425
rect 2973 311 3113 357
<< metal1 >>
rect 0 724 3472 844
rect 262 632 330 724
rect 661 694 707 724
rect 69 619 115 631
rect 262 586 273 632
rect 319 586 330 632
rect 383 596 615 643
rect 661 637 707 648
rect 69 540 115 573
rect 383 540 429 596
rect 569 577 615 596
rect 778 632 1261 678
rect 1307 632 1318 678
rect 778 577 824 632
rect 1526 586 1594 724
rect 69 494 429 540
rect 130 416 318 430
rect 130 370 157 416
rect 203 370 318 416
rect 130 354 318 370
rect 383 313 429 494
rect 477 531 523 542
rect 569 530 824 577
rect 477 465 523 485
rect 477 454 815 465
rect 477 418 769 454
rect 49 267 383 302
rect 769 311 815 408
rect 49 256 429 267
rect 497 265 815 311
rect 49 219 95 256
rect 497 219 543 265
rect 49 162 95 173
rect 262 164 273 210
rect 319 164 330 210
rect 262 60 330 164
rect 497 162 543 173
rect 630 172 641 218
rect 687 172 698 218
rect 630 60 698 172
rect 769 152 815 265
rect 914 311 995 542
rect 1122 540 1133 586
rect 1179 540 1190 586
rect 1526 540 1537 586
rect 1583 540 1594 586
rect 1728 632 2209 678
rect 2255 632 2266 678
rect 1122 494 1190 540
rect 914 265 926 311
rect 972 265 995 311
rect 914 242 995 265
rect 1065 448 1625 494
rect 1671 448 1682 494
rect 1065 244 1134 448
rect 1728 402 1774 632
rect 1065 198 1077 244
rect 1123 198 1134 244
rect 1233 356 1774 402
rect 1825 540 1836 586
rect 1882 540 1894 586
rect 1233 311 1279 356
rect 1825 310 1894 540
rect 1233 152 1279 265
rect 1426 264 1437 310
rect 1483 264 1894 310
rect 1826 218 1894 264
rect 1944 310 1990 632
rect 2525 595 2571 724
rect 2873 689 2919 724
rect 1944 245 1990 264
rect 2050 540 2061 586
rect 2107 540 2118 586
rect 2050 426 2118 540
rect 2525 527 2571 549
rect 2729 595 2775 606
rect 2050 425 2670 426
rect 2050 379 2613 425
rect 2659 379 2670 425
rect 1826 172 1837 218
rect 1883 172 1894 218
rect 2050 218 2118 379
rect 2729 368 2775 549
rect 3333 689 3379 724
rect 2873 527 2919 549
rect 3066 549 3077 595
rect 3123 549 3282 595
rect 3066 466 3282 549
rect 3333 527 3379 549
rect 2729 357 3113 368
rect 2729 326 2973 357
rect 2354 280 2365 326
rect 2411 311 2973 326
rect 2411 300 3113 311
rect 2411 280 2774 300
rect 2050 172 2061 218
rect 2107 172 2118 218
rect 2497 210 2543 221
rect 769 106 1279 152
rect 1558 71 1569 117
rect 1615 71 1626 117
rect 1558 60 1626 71
rect 2497 60 2543 164
rect 2721 218 2774 280
rect 2767 172 2774 218
rect 3206 204 3282 466
rect 2721 161 2774 172
rect 2885 167 2931 178
rect 2885 60 2931 121
rect 3090 167 3282 204
rect 3090 121 3109 167
rect 3155 121 3282 167
rect 3090 110 3282 121
rect 3333 167 3379 194
rect 3333 60 3379 121
rect 0 -60 3472 60
<< labels >>
flabel metal1 s 914 242 995 542 0 FreeSans 600 0 0 0 D
port 1 nsew default input
flabel metal1 s 0 724 3472 844 0 FreeSans 600 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 2497 218 2543 221 0 FreeSans 600 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel metal1 s 130 354 318 430 0 FreeSans 600 0 0 0 CLK
port 2 nsew clock input
flabel metal1 s 3066 466 3282 595 0 FreeSans 600 0 0 0 Q
port 3 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 5 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 6 nsew ground bidirectional
rlabel metal1 s 3206 204 3282 466 1 Q
port 3 nsew default output
rlabel metal1 s 3090 110 3282 204 1 Q
port 3 nsew default output
rlabel metal1 s 3333 637 3379 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2873 637 2919 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2525 637 2571 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1526 637 1594 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 661 637 707 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 262 637 330 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3333 586 3379 637 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2873 586 2919 637 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2525 586 2571 637 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1526 586 1594 637 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 262 586 330 637 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3333 540 3379 586 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2873 540 2919 586 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2525 540 2571 586 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1526 540 1594 586 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3333 527 3379 540 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2873 527 2919 540 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2525 527 2571 540 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2497 210 2543 218 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 630 210 698 218 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2497 194 2543 210 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 630 194 698 210 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 194 330 210 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3333 178 3379 194 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2497 178 2543 194 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 630 178 698 194 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 178 330 194 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3333 117 3379 178 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2885 117 2931 178 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2497 117 2543 178 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 630 117 698 178 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 117 330 178 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3333 60 3379 117 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2885 60 2931 117 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2497 60 2543 117 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1558 60 1626 117 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 630 60 698 117 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 60 330 117 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3472 60 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3472 784
string GDS_END 981854
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 974442
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
