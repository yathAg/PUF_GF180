magic
tech gf180mcuB
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -1789 9497 11222 10481
rect -1789 -266 -560 9497
rect 10028 -266 11222 9497
rect -1789 -834 11222 -266
<< psubdiff >>
rect -528 8756 9996 9430
rect -528 8372 9406 8756
rect -528 -174 -486 8372
rect -140 8195 9406 8372
rect 9586 8372 9996 8756
rect -140 -35 -118 8195
rect 9586 -35 9608 8372
rect -140 -57 9608 -35
rect -140 -174 208 -57
rect -528 -197 208 -174
rect 9278 -174 9608 -57
rect 9954 -174 9996 8372
rect 9278 -197 9996 -174
rect -528 -219 9996 -197
<< nsubdiff >>
rect -1707 10376 11139 10398
rect -1707 10330 -421 10376
rect 9925 10330 11139 10376
rect -1707 10272 11139 10330
rect -1707 10226 -421 10272
rect 9925 10226 11139 10272
rect -1707 10168 11139 10226
rect -1707 10122 -421 10168
rect 9925 10122 11139 10168
rect -1707 10064 11139 10122
rect -1707 10018 -421 10064
rect 9925 10018 11139 10064
rect -1707 9960 11139 10018
rect -1707 9914 -421 9960
rect 9925 9914 11139 9960
rect -1707 9856 11139 9914
rect -1707 9810 -421 9856
rect 9925 9810 11139 9856
rect -1707 9752 11139 9810
rect -1707 9706 -421 9752
rect 9925 9706 11139 9752
rect -1707 9648 11139 9706
rect -1707 9602 -421 9648
rect 9925 9602 11139 9648
rect -1707 9580 11139 9602
rect -1707 8368 -643 9580
rect -1707 22 -1647 8368
rect -1601 22 -1543 8368
rect -1497 22 -1439 8368
rect -1393 22 -1335 8368
rect -1289 22 -1231 8368
rect -1185 22 -1127 8368
rect -1081 22 -1023 8368
rect -977 22 -919 8368
rect -873 22 -815 8368
rect -769 22 -711 8368
rect -665 22 -643 8368
rect -1707 -83 -643 22
rect -1707 -729 -1647 -83
rect -1601 -729 -1543 -83
rect -1497 -729 -1439 -83
rect -1393 -729 -1335 -83
rect -1289 -729 -1231 -83
rect -1185 -729 -1127 -83
rect -1081 -729 -1023 -83
rect -977 -729 -919 -83
rect -873 -729 -815 -83
rect -769 -729 -711 -83
rect -665 -349 -643 -83
rect 10111 8368 11139 9580
rect 10111 22 10133 8368
rect 10179 22 10237 8368
rect 10283 22 10341 8368
rect 10387 22 10445 8368
rect 10491 22 10549 8368
rect 10595 22 10653 8368
rect 10699 22 10757 8368
rect 10803 22 10861 8368
rect 10907 22 10965 8368
rect 11011 22 11069 8368
rect 11115 22 11139 8368
rect 10111 -83 11139 22
rect 10111 -349 10133 -83
rect -665 -371 10133 -349
rect -665 -417 -413 -371
rect 9933 -417 10133 -371
rect -665 -475 10133 -417
rect -665 -521 -413 -475
rect 9933 -521 10133 -475
rect -665 -579 10133 -521
rect -665 -625 -413 -579
rect 9933 -625 10133 -579
rect -665 -683 10133 -625
rect -665 -729 -413 -683
rect 9933 -729 10133 -683
rect 10179 -729 10237 -83
rect 10283 -729 10341 -83
rect 10387 -729 10445 -83
rect 10491 -729 10549 -83
rect 10595 -729 10653 -83
rect 10699 -729 10757 -83
rect 10803 -729 10861 -83
rect 10907 -729 10965 -83
rect 11011 -729 11069 -83
rect 11115 -729 11139 -83
rect -1707 -751 11139 -729
<< psubdiffcont >>
rect -486 -174 -140 8372
rect 208 -197 9278 -57
rect 9608 -174 9954 8372
<< nsubdiffcont >>
rect -421 10330 9925 10376
rect -421 10226 9925 10272
rect -421 10122 9925 10168
rect -421 10018 9925 10064
rect -421 9914 9925 9960
rect -421 9810 9925 9856
rect -421 9706 9925 9752
rect -421 9602 9925 9648
rect -1647 22 -1601 8368
rect -1543 22 -1497 8368
rect -1439 22 -1393 8368
rect -1335 22 -1289 8368
rect -1231 22 -1185 8368
rect -1127 22 -1081 8368
rect -1023 22 -977 8368
rect -919 22 -873 8368
rect -815 22 -769 8368
rect -711 22 -665 8368
rect -1647 -729 -1601 -83
rect -1543 -729 -1497 -83
rect -1439 -729 -1393 -83
rect -1335 -729 -1289 -83
rect -1231 -729 -1185 -83
rect -1127 -729 -1081 -83
rect -1023 -729 -977 -83
rect -919 -729 -873 -83
rect -815 -729 -769 -83
rect -711 -729 -665 -83
rect 10133 22 10179 8368
rect 10237 22 10283 8368
rect 10341 22 10387 8368
rect 10445 22 10491 8368
rect 10549 22 10595 8368
rect 10653 22 10699 8368
rect 10757 22 10803 8368
rect 10861 22 10907 8368
rect 10965 22 11011 8368
rect 11069 22 11115 8368
rect -413 -417 9933 -371
rect -413 -521 9933 -475
rect -413 -625 9933 -579
rect -413 -729 9933 -683
rect 10133 -729 10179 -83
rect 10237 -729 10283 -83
rect 10341 -729 10387 -83
rect 10445 -729 10491 -83
rect 10549 -729 10595 -83
rect 10653 -729 10699 -83
rect 10757 -729 10803 -83
rect 10861 -729 10907 -83
rect 10965 -729 11011 -83
rect 11069 -729 11115 -83
<< metal1 >>
rect -432 10376 9936 10387
rect -432 10330 -421 10376
rect 9925 10330 9936 10376
rect -432 10272 9936 10330
rect -432 10226 -421 10272
rect 9925 10226 9936 10272
rect -432 10168 9936 10226
rect -432 10122 -421 10168
rect 9925 10122 9936 10168
rect -432 10064 9936 10122
rect -432 10018 -421 10064
rect 9925 10018 9936 10064
rect -432 9960 9936 10018
rect -432 9914 -421 9960
rect 9925 9914 9936 9960
rect -432 9856 9936 9914
rect -432 9810 -421 9856
rect 9925 9810 9936 9856
rect -432 9752 9936 9810
rect -432 9706 -421 9752
rect 9925 9706 9936 9752
rect -432 9648 9936 9706
rect -432 9602 -421 9648
rect 9925 9602 9936 9648
rect -432 9591 9936 9602
rect -1658 8368 -654 8388
rect -1658 22 -1647 8368
rect -1601 22 -1543 8368
rect -1497 22 -1439 8368
rect -1393 22 -1335 8368
rect -1289 22 -1231 8368
rect -1185 22 -1127 8368
rect -1081 22 -1023 8368
rect -977 22 -919 8368
rect -873 22 -815 8368
rect -769 22 -711 8368
rect -665 22 -654 8368
rect -1658 -83 -654 22
rect -1658 -729 -1647 -83
rect -1601 -729 -1543 -83
rect -1497 -729 -1439 -83
rect -1393 -729 -1335 -83
rect -1289 -729 -1231 -83
rect -1185 -729 -1127 -83
rect -1081 -729 -1023 -83
rect -977 -729 -919 -83
rect -873 -729 -815 -83
rect -769 -729 -711 -83
rect -665 -360 -654 -83
rect -517 8372 51 8396
rect -517 -174 -486 8372
rect -140 -46 51 8372
rect 9597 8372 9985 8383
rect 9597 -46 9608 8372
rect -140 -57 9608 -46
rect -140 -174 208 -57
rect -517 -197 208 -174
rect 9278 -174 9608 -57
rect 9954 -174 9985 8372
rect 9278 -197 9985 -174
rect -517 -208 9985 -197
rect 10122 8368 11126 8410
rect 10122 22 10133 8368
rect 10179 22 10237 8368
rect 10283 22 10341 8368
rect 10387 22 10445 8368
rect 10491 22 10549 8368
rect 10595 22 10653 8368
rect 10699 22 10757 8368
rect 10803 22 10861 8368
rect 10907 22 10965 8368
rect 11011 22 11069 8368
rect 11115 22 11126 8368
rect 10122 -83 11126 22
rect 10122 -360 10133 -83
rect -665 -371 10133 -360
rect -665 -417 -413 -371
rect 9933 -417 10133 -371
rect -665 -475 10133 -417
rect -665 -521 -413 -475
rect 9933 -521 10133 -475
rect -665 -579 10133 -521
rect -665 -625 -413 -579
rect 9933 -625 10133 -579
rect -665 -683 10133 -625
rect -665 -729 -413 -683
rect 9933 -729 10133 -683
rect 10179 -729 10237 -83
rect 10283 -729 10341 -83
rect 10387 -729 10445 -83
rect 10491 -729 10549 -83
rect 10595 -729 10653 -83
rect 10699 -729 10757 -83
rect 10803 -729 10861 -83
rect 10907 -729 10965 -83
rect 11011 -729 11069 -83
rect 11115 -729 11126 -83
rect -1658 -740 11126 -729
use M1_NWELL_CDNS_40661954729561  M1_NWELL_CDNS_40661954729561_0
timestamp 1698431365
transform 1 0 4752 0 1 9989
box 0 0 1 1
use M1_NWELL_CDNS_40661954729564  M1_NWELL_CDNS_40661954729564_0
timestamp 1698431365
transform 1 0 4760 0 1 -550
box 0 0 1 1
use M1_PSUB_CDNS_40661954729562  M1_PSUB_CDNS_40661954729562_0
timestamp 1698431365
transform 1 0 -313 0 1 4099
box 0 0 1 1
use M1_PSUB_CDNS_40661954729562  M1_PSUB_CDNS_40661954729562_1
timestamp 1698431365
transform 1 0 9781 0 1 4099
box 0 0 1 1
use M1_PSUB_CDNS_40661954729563  M1_PSUB_CDNS_40661954729563_0
timestamp 1698431365
transform 0 -1 4743 1 0 -127
box 0 0 1 1
<< properties >>
string GDS_END 1958388
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 1802970
<< end >>
