magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< obsm1 >>
rect 13108 13108 71000 71000
<< obsm2 >>
rect 13606 13594 70901 70890
<< metal3 >>
rect 14000 70800 17000 71000
rect 17200 70800 20200 71000
rect 20400 70800 23400 71000
rect 23600 70800 25000 71000
rect 25200 70800 26600 71000
rect 26800 70800 29800 71000
rect 30000 70800 33000 71000
rect 33200 70800 36200 71000
rect 36400 70800 39400 71000
rect 39600 70800 41000 71000
rect 41200 70800 42600 71000
rect 42800 70800 45800 71000
rect 46000 70800 49000 71000
rect 49200 70800 50600 71000
rect 50800 70800 52200 71000
rect 52400 70800 53800 71000
rect 54000 70800 55400 71000
rect 55600 70800 57000 71000
rect 57200 70800 58600 71000
rect 58800 70800 60200 71000
rect 60400 70800 61800 71000
rect 62000 70800 63400 71000
rect 63600 70800 65000 71000
rect 65200 70800 66600 71000
rect 66800 70800 68200 71000
rect 68400 70800 69678 71000
rect 70800 68400 71000 69678
rect 70800 66800 71000 68200
rect 70800 65200 71000 66600
rect 70800 63600 71000 65000
rect 70800 62000 71000 63400
rect 70800 60400 71000 61800
rect 70800 58800 71000 60200
rect 70800 57200 71000 58600
rect 70800 55600 71000 57000
rect 70800 54000 71000 55400
rect 70800 52400 71000 53800
rect 70800 50800 71000 52200
rect 70800 49200 71000 50600
rect 70800 46000 71000 49000
rect 70800 42800 71000 45800
rect 70800 41200 71000 42600
rect 70800 39600 71000 41000
rect 70800 36400 71000 39400
rect 70800 33200 71000 36200
rect 70800 30000 71000 33000
rect 70800 26800 71000 29800
rect 70800 25200 71000 26600
rect 70800 23600 71000 25000
rect 70800 20400 71000 23400
rect 70800 17200 71000 20200
rect 70800 14000 71000 17000
<< obsm3 >>
rect 17060 70740 17140 70890
rect 20260 70740 20340 70890
rect 23460 70740 23540 70890
rect 25060 70740 25140 70890
rect 26660 70740 26740 70890
rect 29860 70740 29940 70890
rect 33060 70740 33140 70890
rect 36260 70740 36340 70890
rect 39460 70740 39540 70890
rect 41060 70740 41140 70890
rect 42660 70740 42740 70890
rect 45860 70740 45940 70890
rect 49060 70740 49140 70890
rect 50660 70740 50740 70890
rect 52260 70740 52340 70890
rect 53860 70740 53940 70890
rect 55460 70740 55540 70890
rect 57060 70740 57140 70890
rect 58660 70740 58740 70890
rect 60260 70740 60340 70890
rect 61860 70740 61940 70890
rect 63460 70740 63540 70890
rect 65060 70740 65140 70890
rect 66660 70740 66740 70890
rect 68260 70740 68340 70890
rect 69738 70740 70800 70890
rect 14000 69738 70800 70740
rect 14000 68340 70740 69738
rect 14000 68260 70800 68340
rect 14000 66740 70740 68260
rect 14000 66660 70800 66740
rect 14000 65140 70740 66660
rect 14000 65060 70800 65140
rect 14000 63540 70740 65060
rect 14000 63460 70800 63540
rect 14000 61940 70740 63460
rect 14000 61860 70800 61940
rect 14000 60340 70740 61860
rect 14000 60260 70800 60340
rect 14000 58740 70740 60260
rect 14000 58660 70800 58740
rect 14000 57140 70740 58660
rect 14000 57060 70800 57140
rect 14000 55540 70740 57060
rect 14000 55460 70800 55540
rect 14000 53940 70740 55460
rect 14000 53860 70800 53940
rect 14000 52340 70740 53860
rect 14000 52260 70800 52340
rect 14000 50740 70740 52260
rect 14000 50660 70800 50740
rect 14000 49140 70740 50660
rect 14000 49060 70800 49140
rect 14000 45940 70740 49060
rect 14000 45860 70800 45940
rect 14000 42740 70740 45860
rect 14000 42660 70800 42740
rect 14000 41140 70740 42660
rect 14000 41060 70800 41140
rect 14000 39540 70740 41060
rect 14000 39460 70800 39540
rect 14000 36340 70740 39460
rect 14000 36260 70800 36340
rect 14000 33140 70740 36260
rect 14000 33060 70800 33140
rect 14000 29940 70740 33060
rect 14000 29860 70800 29940
rect 14000 26740 70740 29860
rect 14000 26660 70800 26740
rect 14000 25140 70740 26660
rect 14000 25060 70800 25140
rect 14000 23540 70740 25060
rect 14000 23460 70800 23540
rect 14000 20340 70740 23460
rect 14000 20260 70800 20340
rect 14000 17140 70740 20260
rect 14000 17060 70800 17140
rect 14000 14000 70740 17060
<< metal4 >>
rect 14000 70800 17000 71000
rect 17200 70800 20200 71000
rect 20400 70800 23400 71000
rect 23600 70800 25000 71000
rect 25200 70800 26600 71000
rect 26800 70800 29800 71000
rect 30000 70800 33000 71000
rect 33200 70800 36200 71000
rect 36400 70800 39400 71000
rect 39600 70800 41000 71000
rect 41200 70800 42600 71000
rect 42800 70800 45800 71000
rect 46000 70800 49000 71000
rect 49200 70800 50600 71000
rect 50800 70800 52200 71000
rect 52400 70800 53800 71000
rect 54000 70800 55400 71000
rect 55600 70800 57000 71000
rect 57200 70800 58600 71000
rect 58800 70800 60200 71000
rect 60400 70800 61800 71000
rect 62000 70800 63400 71000
rect 63600 70800 65000 71000
rect 65200 70800 66600 71000
rect 66800 70800 68200 71000
rect 68400 70800 69678 71000
rect 34408 70196 34464 70252
rect 70800 68400 71000 69678
rect 70800 66800 71000 68200
rect 70800 65200 71000 66600
rect 70800 63600 71000 65000
rect 70800 62000 71000 63400
rect 70800 60400 71000 61800
rect 70800 58800 71000 60200
rect 70800 57200 71000 58600
rect 70800 55600 71000 57000
rect 70800 54000 71000 55400
rect 70390 53138 70446 53194
rect 70800 52400 71000 53800
rect 70517 51406 70573 51462
rect 70800 50800 71000 52200
rect 70516 49938 70572 49994
rect 70800 49200 71000 50600
rect 70800 46000 71000 49000
rect 70800 42800 71000 45800
rect 70800 41200 71000 42600
rect 70800 39600 71000 41000
rect 70800 36400 71000 39400
rect 70800 33200 71000 36200
rect 70800 30000 71000 33000
rect 70800 26800 71000 29800
rect 70800 25200 71000 26600
rect 70800 23600 71000 25000
rect 70800 20400 71000 23400
rect 70800 17200 71000 20200
rect 70800 14000 71000 17000
<< obsm4 >>
rect 17060 70740 17140 70800
rect 20260 70740 20340 70800
rect 23460 70740 23540 70800
rect 25060 70740 25140 70800
rect 26660 70740 26740 70800
rect 29860 70740 29940 70800
rect 33060 70740 33140 70800
rect 36260 70740 36340 70800
rect 39460 70740 39540 70800
rect 41060 70740 41140 70800
rect 42660 70740 42740 70800
rect 45860 70740 45940 70800
rect 49060 70740 49140 70800
rect 50660 70740 50740 70800
rect 52260 70740 52340 70800
rect 53860 70740 53940 70800
rect 55460 70740 55540 70800
rect 57060 70740 57140 70800
rect 58660 70740 58740 70800
rect 60260 70740 60340 70800
rect 61860 70740 61940 70800
rect 63460 70740 63540 70800
rect 65060 70740 65140 70800
rect 66660 70740 66740 70800
rect 68260 70740 68340 70800
rect 69738 70740 70800 70800
rect 14000 70252 70800 70740
rect 14000 70196 34408 70252
rect 34464 70196 70800 70252
rect 14000 69738 70800 70196
rect 14000 68340 70740 69738
rect 14000 68260 70800 68340
rect 14000 66740 70740 68260
rect 14000 66660 70800 66740
rect 14000 65140 70740 66660
rect 14000 65060 70800 65140
rect 14000 63540 70740 65060
rect 14000 63460 70800 63540
rect 14000 61940 70740 63460
rect 14000 61860 70800 61940
rect 14000 60340 70740 61860
rect 14000 60260 70800 60340
rect 14000 58740 70740 60260
rect 14000 58660 70800 58740
rect 14000 57140 70740 58660
rect 14000 57060 70800 57140
rect 14000 55540 70740 57060
rect 14000 55460 70800 55540
rect 14000 53940 70740 55460
rect 14000 53860 70800 53940
rect 14000 53194 70740 53860
rect 14000 53138 70390 53194
rect 70446 53138 70740 53194
rect 14000 52340 70740 53138
rect 14000 52260 70800 52340
rect 14000 51462 70740 52260
rect 14000 51406 70517 51462
rect 70573 51406 70740 51462
rect 14000 50740 70740 51406
rect 14000 50660 70800 50740
rect 14000 49994 70740 50660
rect 14000 49938 70516 49994
rect 70572 49938 70740 49994
rect 14000 49140 70740 49938
rect 14000 49060 70800 49140
rect 14000 45940 70740 49060
rect 14000 45860 70800 45940
rect 14000 42740 70740 45860
rect 14000 42660 70800 42740
rect 14000 41140 70740 42660
rect 14000 41060 70800 41140
rect 14000 39540 70740 41060
rect 14000 39460 70800 39540
rect 14000 36340 70740 39460
rect 14000 36260 70800 36340
rect 14000 33140 70740 36260
rect 14000 33060 70800 33140
rect 14000 29940 70740 33060
rect 14000 29860 70800 29940
rect 14000 26740 70740 29860
rect 14000 26660 70800 26740
rect 14000 25140 70740 26660
rect 14000 25060 70800 25140
rect 14000 23540 70740 25060
rect 14000 23460 70800 23540
rect 14000 20340 70740 23460
rect 14000 20260 70800 20340
rect 14000 17140 70740 20260
rect 14000 17060 70800 17140
rect 14000 14000 70740 17060
<< metal5 >>
rect 14000 70800 17000 71000
rect 17200 70800 20200 71000
rect 20400 70800 23400 71000
rect 23600 70800 25000 71000
rect 25200 70800 26600 71000
rect 26800 70800 29800 71000
rect 30000 70800 33000 71000
rect 33200 70800 36200 71000
rect 36400 70800 39400 71000
rect 39600 70800 41000 71000
rect 41200 70800 42600 71000
rect 42800 70800 45800 71000
rect 46000 70800 49000 71000
rect 49200 70800 50600 71000
rect 50800 70800 52200 71000
rect 52400 70800 53800 71000
rect 54000 70800 55400 71000
rect 55600 70800 57000 71000
rect 57200 70800 58600 71000
rect 58800 70800 60200 71000
rect 60400 70800 61800 71000
rect 62000 70800 63400 71000
rect 63600 70800 65000 71000
rect 65200 70800 66600 71000
rect 66800 70800 68200 71000
rect 68400 70800 69678 71000
rect 15396 47287 15472 70800
rect 18596 48623 18672 70800
rect 20400 70151 23400 70227
rect 23600 70160 25000 70236
rect 25200 70164 26600 70240
rect 28064 52629 28140 70800
rect 31264 53967 31340 70800
rect 34408 70196 34464 70252
rect 37664 56640 37740 70800
rect 40262 57314 40338 70800
rect 41862 57986 41938 70800
rect 42800 70148 45800 70224
rect 46000 70171 49000 70247
rect 49200 70176 50600 70252
rect 51462 62015 51538 70800
rect 53062 62683 53138 70800
rect 54662 63349 54738 70800
rect 56262 64012 56338 70800
rect 57862 64675 57938 70800
rect 59462 65342 59538 70800
rect 61062 66007 61138 70800
rect 62662 66670 62738 70800
rect 64262 67342 64338 70800
rect 65867 68000 65943 70800
rect 67462 68669 67538 70800
rect 69001 69258 69077 70800
rect 70395 68400 70471 69678
rect 70800 68400 71000 69678
rect 70402 66800 70478 68200
rect 70800 66800 71000 68200
rect 70400 65200 70476 66600
rect 70800 65200 71000 66600
rect 70399 63600 70475 65000
rect 70800 63600 71000 65000
rect 70393 62000 70469 63400
rect 70800 62000 71000 63400
rect 70391 60400 70467 61800
rect 70800 60400 71000 61800
rect 70389 58800 70465 60200
rect 70800 58800 71000 60200
rect 70386 57200 70462 58600
rect 70800 57200 71000 58600
rect 70384 55600 70460 57000
rect 70800 55600 71000 57000
rect 70382 54000 70458 55400
rect 70800 54000 71000 55400
rect 70390 53138 70446 53194
rect 70800 52400 71000 53800
rect 70517 51406 70573 51462
rect 70800 50800 71000 52200
rect 70516 49938 70572 49994
rect 70800 49200 71000 50600
rect 70800 47604 71000 49000
rect 60617 47528 71000 47604
rect 70800 46000 71000 47528
rect 70412 42800 70488 45800
rect 70800 42800 71000 45800
rect 70407 41200 70483 42600
rect 70800 41200 71000 42600
rect 70401 39600 70477 41000
rect 70800 39600 71000 41000
rect 70394 36400 70470 39400
rect 70800 36400 71000 39400
rect 70384 33200 70460 36200
rect 70800 33200 71000 36200
rect 70800 31604 71000 33000
rect 58681 31528 71000 31604
rect 70800 30000 71000 31528
rect 70800 28404 71000 29800
rect 58681 28328 71000 28404
rect 70800 26800 71000 28328
rect 70800 26070 71000 26600
rect 51296 25994 71000 26070
rect 70800 25200 71000 25994
rect 70424 23600 70500 25000
rect 70800 23600 71000 25000
rect 70415 20400 70491 23400
rect 70800 20400 71000 23400
rect 70800 18936 71000 20200
rect 58405 18860 71000 18936
rect 70800 17200 71000 18860
rect 70404 14000 70480 17000
rect 70800 14000 71000 17000
<< obsm5 >>
rect 14000 47167 15276 70680
rect 15592 48503 18476 70680
rect 18792 70360 27944 70680
rect 18792 70356 25080 70360
rect 18792 70347 23480 70356
rect 18792 70031 20280 70347
rect 26720 70044 27944 70360
rect 25120 70040 27944 70044
rect 23520 70031 27944 70040
rect 18792 52509 27944 70031
rect 28260 53847 31144 70680
rect 31460 70372 37544 70680
rect 31460 70076 34288 70372
rect 34584 70076 37544 70372
rect 31460 56520 37544 70076
rect 37860 57194 40142 70680
rect 40458 57866 41742 70680
rect 42058 70372 51342 70680
rect 42058 70367 49080 70372
rect 42058 70344 45880 70367
rect 42058 70028 42680 70344
rect 50720 70056 51342 70372
rect 49120 70051 51342 70056
rect 45920 70028 51342 70051
rect 42058 61895 51342 70028
rect 51658 62563 52942 70680
rect 53258 63229 54542 70680
rect 54858 63892 56142 70680
rect 56458 64555 57742 70680
rect 58058 65222 59342 70680
rect 59658 65887 60942 70680
rect 61258 66550 62542 70680
rect 62858 67222 64142 70680
rect 64458 67880 65747 70680
rect 66063 68549 67342 70680
rect 67658 69138 68881 70680
rect 69798 70680 70800 70800
rect 69197 69798 70800 70680
rect 69197 69138 70275 69798
rect 67658 68549 70275 69138
rect 66063 68280 70275 68549
rect 70591 68320 70680 69798
rect 66063 67880 70282 68280
rect 64458 67222 70282 67880
rect 62858 66720 70282 67222
rect 62858 66550 70280 66720
rect 70598 66680 70680 68320
rect 61258 65887 70280 66550
rect 59658 65222 70280 65887
rect 58058 65120 70280 65222
rect 58058 64555 70279 65120
rect 70596 65080 70680 66680
rect 56458 63892 70279 64555
rect 54858 63520 70279 63892
rect 54858 63229 70273 63520
rect 70595 63480 70680 65080
rect 53258 62563 70273 63229
rect 51658 61920 70273 62563
rect 51658 61895 70271 61920
rect 42058 60320 70271 61895
rect 70589 61880 70680 63480
rect 42058 58720 70269 60320
rect 70587 60280 70680 61880
rect 42058 57866 70266 58720
rect 70585 58680 70680 60280
rect 40458 57194 70266 57866
rect 37860 57120 70266 57194
rect 37860 56520 70264 57120
rect 70582 57080 70680 58680
rect 31460 55520 70264 56520
rect 31460 53880 70262 55520
rect 70580 55480 70680 57080
rect 70578 53880 70680 55480
rect 31460 53847 70680 53880
rect 28260 53314 70680 53847
rect 28260 53018 70270 53314
rect 70566 53018 70680 53314
rect 28260 52509 70680 53018
rect 18792 51582 70680 52509
rect 18792 51286 70397 51582
rect 18792 50114 70680 51286
rect 18792 49818 70396 50114
rect 18792 48503 70680 49818
rect 15592 47724 70680 48503
rect 15592 47408 60497 47724
rect 15592 47167 70680 47408
rect 14000 45920 70680 47167
rect 14000 42720 70292 45920
rect 14000 41120 70287 42720
rect 70608 42680 70680 45920
rect 14000 39520 70281 41120
rect 70603 41080 70680 42680
rect 14000 36320 70274 39520
rect 70597 39480 70680 41080
rect 14000 33080 70264 36320
rect 70590 36280 70680 39480
rect 70580 33080 70680 36280
rect 14000 31724 70680 33080
rect 14000 31408 58561 31724
rect 14000 28524 70680 31408
rect 14000 28208 58561 28524
rect 14000 26190 70680 28208
rect 14000 25874 51176 26190
rect 14000 25120 70680 25874
rect 14000 23520 70304 25120
rect 14000 20280 70295 23520
rect 70620 23480 70680 25120
rect 70611 20280 70680 23480
rect 14000 19056 70680 20280
rect 14000 18740 58285 19056
rect 14000 17120 70680 18740
rect 14000 14000 70284 17120
rect 70600 14000 70680 17120
<< labels >>
rlabel metal3 s 66800 70800 68200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 66800 71000 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 58800 70800 60200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 58800 71000 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 55600 70800 57000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 55600 71000 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 54000 70800 55400 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 54000 71000 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 52400 70800 53800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 52400 71000 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 42800 70800 45800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 42800 71000 45800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 41200 70800 42600 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 41200 71000 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 36400 70800 39400 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 36400 71000 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 33200 70800 36200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 33200 71000 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 30000 70800 33000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 30000 71000 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 26800 70800 29800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 26800 71000 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 23600 70800 25000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 66800 70800 68200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 66800 71000 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 58800 70800 60200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 58800 71000 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 55600 70800 57000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 55600 71000 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 54000 70800 55400 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 54000 71000 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 52400 70800 53800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 52400 71000 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 42800 70800 45800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 42800 71000 45800 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 41200 70800 42600 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 41200 71000 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 36400 70800 39400 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 36400 71000 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 33200 70800 36200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 33200 71000 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 30000 70800 33000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 30000 71000 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 26800 70800 29800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 26800 71000 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 23600 70800 25000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 66800 70800 68200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 66800 71000 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 58800 70800 60200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 58800 71000 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 55600 70800 57000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 55600 71000 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 54000 70800 55400 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 54000 71000 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 52400 70800 53800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 52400 71000 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 42800 70800 45800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 42800 71000 45800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 41200 70800 42600 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 41200 71000 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 36400 70800 39400 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 36400 71000 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 33200 70800 36200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 33200 71000 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 30000 70800 33000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 30000 71000 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 26800 70800 29800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 26800 71000 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 23600 70800 25000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 23600 71000 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 23600 71000 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 23600 71000 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 67462 68669 67538 70800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70412 42800 70488 45800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70390 53138 70446 53194 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70390 53138 70446 53194 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70382 54000 70458 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70384 55600 70460 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70389 58800 70465 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70402 66800 70478 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 42800 70148 45800 70224 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 53062 62683 53138 70800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 54662 63349 54738 70800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 56262 64012 56338 70800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 59462 65342 59538 70800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 41862 57986 41938 70800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 37664 56640 37740 70800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 23600 70160 25000 70236 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 28064 52629 28140 70800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 31264 53967 31340 70800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 34408 70196 34464 70252 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 34408 70196 34464 70252 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70394 36400 70470 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70407 41200 70483 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 58681 31528 70800 31604 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70384 33200 70460 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70424 23600 70500 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 58681 28328 70800 28404 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 68400 70800 69678 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 68400 71000 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 65200 70800 66600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 65200 71000 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 60400 70800 61800 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 60400 71000 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 57200 70800 58600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 57200 71000 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 46000 70800 49000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 46000 71000 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 39600 70800 41000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 39600 71000 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 25200 70800 26600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 25200 71000 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 20400 70800 23400 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 20400 71000 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 17200 70800 20200 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 17200 71000 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 14000 70800 17000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 68400 70800 69678 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 68400 71000 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 65200 70800 66600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 65200 71000 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 60400 70800 61800 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 60400 71000 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 57200 70800 58600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 57200 71000 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 46000 70800 49000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 46000 71000 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 39600 70800 41000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 39600 71000 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 25200 70800 26600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 25200 71000 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 20400 70800 23400 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 20400 71000 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 17200 70800 20200 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 17200 71000 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 14000 70800 17000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 68400 70800 69678 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 68400 71000 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 65200 70800 66600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 65200 71000 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 60400 70800 61800 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 60400 71000 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 57200 70800 58600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 57200 71000 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 46000 70800 49000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 46000 71000 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 39600 70800 41000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 39600 71000 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 25200 70800 26600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 25200 71000 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 20400 70800 23400 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 20400 71000 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 17200 70800 20200 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 17200 71000 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 14000 70800 17000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 14000 71000 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 14000 71000 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 14000 71000 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 69001 69258 69077 70800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 60617 47528 70800 47604 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70386 57200 70462 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70391 60400 70467 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70400 65200 70476 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70395 68400 70471 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 46000 70171 49000 70247 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 57862 64675 57938 70800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 61062 66007 61138 70800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 65867 68000 65943 70800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 40262 57314 40338 70800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 15396 47287 15472 70800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 18596 48623 18672 70800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 20400 70151 23400 70227 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 25200 70164 26600 70240 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 58405 18860 70800 18936 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70404 14000 70480 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70415 20400 70491 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 51296 25994 70800 26070 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70401 39600 70477 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 62000 70800 63400 71000 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 70800 62000 71000 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 50800 70800 52200 71000 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 62000 70800 63400 71000 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 70800 62000 71000 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 50800 70800 52200 71000 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 62000 70800 63400 71000 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 70800 62000 71000 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 50800 70800 52200 71000 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 70800 50800 71000 52200 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 70800 50800 71000 52200 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 70800 50800 71000 52200 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 70517 51406 70573 51462 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 70517 51406 70573 51462 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 70393 62000 70469 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 51462 62015 51538 70800 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 62662 66670 62738 70800 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 63600 70800 65000 71000 6 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 70800 63600 71000 65000 6 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 49200 70800 50600 71000 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 63600 70800 65000 71000 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 70800 63600 71000 65000 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 49200 70800 50600 71000 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 63600 70800 65000 71000 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 70800 63600 71000 65000 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 49200 70800 50600 71000 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 70800 49200 71000 50600 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 70800 49200 71000 50600 6 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 70800 49200 71000 50600 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 70516 49938 70572 49994 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 70516 49938 70572 49994 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 70399 63600 70475 65000 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 49200 70176 50600 70252 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 64262 67342 64338 70800 6 VSS
port 4 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 71000 71000
string LEFclass ENDCAP BOTTOMLEFT
string LEFsite GF_COR_Site
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 17526672
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 17515934
<< end >>
