magic
tech gf180mcuA
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 453 2998 1094
<< pwell >>
rect -86 -86 2998 453
<< mvnmos >>
rect 124 69 244 333
rect 348 69 468 333
rect 572 69 692 333
rect 796 69 916 333
rect 1020 69 1140 333
rect 1244 69 1364 333
rect 1468 69 1588 333
rect 1692 69 1812 333
rect 1916 69 2036 333
rect 2140 69 2260 333
rect 2364 69 2484 333
rect 2588 69 2708 333
<< mvpmos >>
rect 124 573 224 939
rect 348 573 448 939
rect 572 573 672 939
rect 796 573 896 939
rect 1020 573 1120 939
rect 1244 573 1344 939
rect 1468 573 1568 939
rect 1692 573 1792 939
rect 1916 573 2016 939
rect 2140 573 2240 939
rect 2364 573 2464 939
rect 2588 573 2688 939
<< mvndiff >>
rect 36 287 124 333
rect 36 147 49 287
rect 95 147 124 287
rect 36 69 124 147
rect 244 287 348 333
rect 244 147 273 287
rect 319 147 348 287
rect 244 69 348 147
rect 468 287 572 333
rect 468 147 497 287
rect 543 147 572 287
rect 468 69 572 147
rect 692 287 796 333
rect 692 147 721 287
rect 767 147 796 287
rect 692 69 796 147
rect 916 287 1020 333
rect 916 147 945 287
rect 991 147 1020 287
rect 916 69 1020 147
rect 1140 287 1244 333
rect 1140 147 1169 287
rect 1215 147 1244 287
rect 1140 69 1244 147
rect 1364 287 1468 333
rect 1364 147 1393 287
rect 1439 147 1468 287
rect 1364 69 1468 147
rect 1588 287 1692 333
rect 1588 147 1617 287
rect 1663 147 1692 287
rect 1588 69 1692 147
rect 1812 222 1916 333
rect 1812 82 1841 222
rect 1887 82 1916 222
rect 1812 69 1916 82
rect 2036 287 2140 333
rect 2036 147 2065 287
rect 2111 147 2140 287
rect 2036 69 2140 147
rect 2260 287 2364 333
rect 2260 147 2289 287
rect 2335 147 2364 287
rect 2260 69 2364 147
rect 2484 287 2588 333
rect 2484 147 2513 287
rect 2559 147 2588 287
rect 2484 69 2588 147
rect 2708 287 2796 333
rect 2708 147 2737 287
rect 2783 147 2796 287
rect 2708 69 2796 147
<< mvpdiff >>
rect 36 861 124 939
rect 36 721 49 861
rect 95 721 124 861
rect 36 573 124 721
rect 224 861 348 939
rect 224 721 273 861
rect 319 721 348 861
rect 224 573 348 721
rect 448 861 572 939
rect 448 721 477 861
rect 523 721 572 861
rect 448 573 572 721
rect 672 861 796 939
rect 672 721 701 861
rect 747 721 796 861
rect 672 573 796 721
rect 896 861 1020 939
rect 896 721 925 861
rect 971 721 1020 861
rect 896 573 1020 721
rect 1120 861 1244 939
rect 1120 721 1169 861
rect 1215 721 1244 861
rect 1120 573 1244 721
rect 1344 861 1468 939
rect 1344 721 1373 861
rect 1419 721 1468 861
rect 1344 573 1468 721
rect 1568 861 1692 939
rect 1568 721 1597 861
rect 1643 721 1692 861
rect 1568 573 1692 721
rect 1792 861 1916 939
rect 1792 721 1821 861
rect 1867 721 1916 861
rect 1792 573 1916 721
rect 2016 861 2140 939
rect 2016 721 2045 861
rect 2091 721 2140 861
rect 2016 573 2140 721
rect 2240 861 2364 939
rect 2240 721 2269 861
rect 2315 721 2364 861
rect 2240 573 2364 721
rect 2464 861 2588 939
rect 2464 721 2493 861
rect 2539 721 2588 861
rect 2464 573 2588 721
rect 2688 861 2776 939
rect 2688 721 2717 861
rect 2763 721 2776 861
rect 2688 573 2776 721
<< mvndiffc >>
rect 49 147 95 287
rect 273 147 319 287
rect 497 147 543 287
rect 721 147 767 287
rect 945 147 991 287
rect 1169 147 1215 287
rect 1393 147 1439 287
rect 1617 147 1663 287
rect 1841 82 1887 222
rect 2065 147 2111 287
rect 2289 147 2335 287
rect 2513 147 2559 287
rect 2737 147 2783 287
<< mvpdiffc >>
rect 49 721 95 861
rect 273 721 319 861
rect 477 721 523 861
rect 701 721 747 861
rect 925 721 971 861
rect 1169 721 1215 861
rect 1373 721 1419 861
rect 1597 721 1643 861
rect 1821 721 1867 861
rect 2045 721 2091 861
rect 2269 721 2315 861
rect 2493 721 2539 861
rect 2717 721 2763 861
<< polysilicon >>
rect 124 939 224 983
rect 348 939 448 983
rect 572 939 672 983
rect 796 939 896 983
rect 1020 939 1120 983
rect 1244 939 1344 983
rect 1468 939 1568 983
rect 1692 939 1792 983
rect 1916 939 2016 983
rect 2140 939 2240 983
rect 2364 939 2464 983
rect 2588 939 2688 983
rect 124 513 224 573
rect 348 513 448 573
rect 572 513 672 573
rect 796 513 896 573
rect 124 500 896 513
rect 124 454 137 500
rect 841 454 896 500
rect 124 441 896 454
rect 124 333 244 441
rect 348 333 468 441
rect 572 333 692 441
rect 796 377 896 441
rect 1020 513 1120 573
rect 1244 513 1344 573
rect 1468 513 1568 573
rect 1692 513 1792 573
rect 1020 512 1792 513
rect 1916 513 2016 573
rect 2140 513 2240 573
rect 2364 513 2464 573
rect 2588 513 2688 573
rect 1916 512 2688 513
rect 1020 500 2688 512
rect 1020 454 1033 500
rect 1737 454 1940 500
rect 2644 454 2688 500
rect 1020 441 2688 454
rect 796 333 916 377
rect 1020 333 1140 441
rect 1244 333 1364 441
rect 1548 377 1588 441
rect 1468 333 1588 377
rect 1692 333 1812 441
rect 1916 333 2036 441
rect 2140 333 2260 441
rect 2364 333 2484 441
rect 2588 377 2688 441
rect 2588 333 2708 377
rect 124 25 244 69
rect 348 25 468 69
rect 572 25 692 69
rect 796 25 916 69
rect 1020 25 1140 69
rect 1244 25 1364 69
rect 1468 25 1588 69
rect 1692 25 1812 69
rect 1916 25 2036 69
rect 2140 25 2260 69
rect 2364 25 2484 69
rect 2588 25 2708 69
<< polycontact >>
rect 137 454 841 500
rect 1033 454 1737 500
rect 1940 454 2644 500
<< metal1 >>
rect 0 918 2912 1098
rect 49 861 95 918
rect 49 710 95 721
rect 273 861 319 872
rect 273 641 319 721
rect 477 861 523 918
rect 477 710 523 721
rect 701 861 747 872
rect 701 641 747 721
rect 925 861 971 918
rect 925 710 971 721
rect 1169 861 1215 872
rect 1169 664 1215 721
rect 1373 861 1419 918
rect 1373 710 1419 721
rect 1597 861 1643 872
rect 1597 664 1643 721
rect 1821 861 1867 918
rect 1821 710 1867 721
rect 2045 861 2091 872
rect 2045 664 2091 721
rect 2269 861 2315 918
rect 2269 710 2315 721
rect 2493 861 2539 872
rect 2493 664 2539 721
rect 2717 861 2763 918
rect 2717 710 2763 721
rect 273 595 933 641
rect 887 530 933 595
rect 1169 576 2539 664
rect 137 500 841 530
rect 137 443 841 454
rect 887 500 1748 530
rect 887 454 1033 500
rect 1737 454 1748 500
rect 887 397 933 454
rect 1794 408 1894 576
rect 1940 500 2644 530
rect 1940 443 2644 454
rect 273 351 933 397
rect 1169 397 1894 408
rect 49 287 95 298
rect 49 90 95 147
rect 273 287 319 351
rect 273 136 319 147
rect 497 287 543 298
rect 497 90 543 147
rect 721 287 767 351
rect 1169 344 2559 397
rect 721 136 767 147
rect 945 287 991 298
rect 945 90 991 147
rect 1169 287 1215 344
rect 1169 136 1215 147
rect 1393 287 1439 298
rect 1393 90 1439 147
rect 1611 287 1663 344
rect 1611 147 1617 287
rect 2065 287 2111 344
rect 1611 136 1663 147
rect 1841 222 1887 233
rect 0 82 1841 90
rect 2065 136 2111 147
rect 2289 287 2335 298
rect 2289 90 2335 147
rect 2513 287 2559 344
rect 2513 136 2559 147
rect 2737 287 2783 298
rect 2737 90 2783 147
rect 1887 82 2912 90
rect 0 -90 2912 82
<< labels >>
flabel metal1 s 137 443 841 530 0 FreeSans 200 0 0 0 I
port 1 nsew default input
flabel metal1 s 0 918 2912 1098 0 FreeSans 200 0 0 0 VDD
port 3 nsew power bidirectional abutment
flabel metal1 s 2737 233 2783 298 0 FreeSans 200 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel metal1 s 2493 664 2539 872 0 FreeSans 200 0 0 0 Z
port 2 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 4 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 2045 664 2091 872 1 Z
port 2 nsew default output
rlabel metal1 s 1597 664 1643 872 1 Z
port 2 nsew default output
rlabel metal1 s 1169 664 1215 872 1 Z
port 2 nsew default output
rlabel metal1 s 1169 576 2539 664 1 Z
port 2 nsew default output
rlabel metal1 s 1794 408 1894 576 1 Z
port 2 nsew default output
rlabel metal1 s 1169 397 1894 408 1 Z
port 2 nsew default output
rlabel metal1 s 1169 344 2559 397 1 Z
port 2 nsew default output
rlabel metal1 s 2513 136 2559 344 1 Z
port 2 nsew default output
rlabel metal1 s 2065 136 2111 344 1 Z
port 2 nsew default output
rlabel metal1 s 1611 136 1663 344 1 Z
port 2 nsew default output
rlabel metal1 s 1169 136 1215 344 1 Z
port 2 nsew default output
rlabel metal1 s 2717 710 2763 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2269 710 2315 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1821 710 1867 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1373 710 1419 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 925 710 971 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 477 710 523 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 710 95 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2289 233 2335 298 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1393 233 1439 298 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 945 233 991 298 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 497 233 543 298 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 49 233 95 298 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2737 90 2783 233 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2289 90 2335 233 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1841 90 1887 233 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1393 90 1439 233 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 945 90 991 233 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 497 90 543 233 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 49 90 95 233 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 2912 90 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2912 1008
string GDS_END 1282152
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1273938
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
