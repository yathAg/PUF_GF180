magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 352 4566 870
<< pwell >>
rect -86 -86 4566 352
<< metal1 >>
rect 0 724 4480 844
rect 297 657 365 724
rect 1293 657 1361 724
rect 2349 657 2417 724
rect 186 240 671 320
rect 3492 506 3538 724
rect 3696 479 3742 676
rect 3905 525 3973 724
rect 4144 479 4238 676
rect 4348 506 4394 724
rect 3696 433 4238 479
rect 4144 230 4238 433
rect 3685 184 4238 230
rect 3685 146 3753 184
rect 317 60 385 127
rect 1333 60 1401 127
rect 2389 60 2457 127
rect 3436 60 3482 138
rect 3920 60 3966 138
rect 4144 135 4238 184
rect 4368 60 4414 138
rect 0 -60 4480 60
<< obsm1 >>
rect 49 481 117 621
rect 49 413 653 481
rect 49 180 95 413
rect 744 361 790 632
rect 877 575 1158 621
rect 744 293 1066 361
rect 1112 350 1158 575
rect 1780 564 1857 632
rect 1933 575 2214 621
rect 1780 361 1826 564
rect 1112 304 1623 350
rect 49 134 117 180
rect 744 154 821 293
rect 1112 200 1158 304
rect 897 154 1158 200
rect 1780 293 2122 361
rect 2168 350 2214 575
rect 2836 564 2913 632
rect 2836 375 2882 564
rect 3000 493 3046 632
rect 3000 447 3376 493
rect 2168 304 2679 350
rect 2836 307 3272 375
rect 3330 364 3376 447
rect 3330 318 4013 364
rect 1780 143 1826 293
rect 2168 200 2214 304
rect 1953 154 2214 200
rect 2836 143 2882 307
rect 3330 200 3376 318
rect 2989 154 3376 200
<< labels >>
rlabel metal1 s 186 240 671 320 6 I
port 1 nsew default input
rlabel metal1 s 4144 135 4238 184 6 Z
port 2 nsew default output
rlabel metal1 s 3685 146 3753 184 6 Z
port 2 nsew default output
rlabel metal1 s 3685 184 4238 230 6 Z
port 2 nsew default output
rlabel metal1 s 4144 230 4238 433 6 Z
port 2 nsew default output
rlabel metal1 s 3696 433 4238 479 6 Z
port 2 nsew default output
rlabel metal1 s 4144 479 4238 676 6 Z
port 2 nsew default output
rlabel metal1 s 3696 479 3742 676 6 Z
port 2 nsew default output
rlabel metal1 s 4348 506 4394 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3905 525 3973 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3492 506 3538 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2349 657 2417 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1293 657 1361 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 297 657 365 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 724 4480 844 6 VDD
port 3 nsew power bidirectional abutment
rlabel nwell s -86 352 4566 870 6 VNW
port 4 nsew power bidirectional
rlabel pwell s -86 -86 4566 352 6 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 0 -60 4480 60 8 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 4368 60 4414 138 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3920 60 3966 138 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3436 60 3482 138 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2389 60 2457 127 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1333 60 1401 127 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 317 60 385 127 6 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4480 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1144252
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1136152
<< end >>
