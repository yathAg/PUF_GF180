magic
tech gf180mcuA
magscale 1 10
timestamp 1698431365
<< psubdiff >>
rect 0 69946 15000 69968
rect 0 69897 210 69946
rect 0 13151 25 69897
rect 71 69800 210 69897
rect 14856 69897 15000 69946
rect 14856 69800 14929 69897
rect 71 69778 14929 69800
rect 71 13287 93 69778
rect 14907 13287 14929 69778
rect 71 13265 14929 13287
rect 71 13151 210 13265
rect 0 13119 210 13151
rect 14856 13151 14929 13265
rect 14975 13151 15000 69897
rect 14856 13119 15000 13151
rect 0 13097 15000 13119
<< psubdiffcont >>
rect 25 13151 71 69897
rect 210 69800 14856 69946
rect 210 13119 14856 13265
rect 14929 13151 14975 69897
<< metal1 >>
rect -32 69946 15032 69957
rect -32 69897 210 69946
rect -32 13151 25 69897
rect 71 69800 210 69897
rect 14856 69897 15032 69946
rect 14856 69800 14929 69897
rect 71 69789 14929 69800
rect 71 13276 82 69789
rect 14918 13276 14929 69789
rect 71 13265 14929 13276
rect 71 13151 210 13265
rect -32 13119 210 13151
rect 14856 13151 14929 13265
rect 14975 13151 15032 69897
rect 14856 13119 15032 13151
rect -32 13108 15032 13119
<< metal3 >>
rect 0 68400 15000 69678
rect 0 66800 15000 68200
rect 0 65200 15000 66600
rect 0 63600 15000 65000
rect 0 62000 15000 63400
rect 0 60400 15000 61800
rect 0 58800 15000 60200
rect 0 57200 15000 58600
rect 0 55600 15000 57000
rect 937 55400 3937 55600
rect 4337 55400 7337 55600
rect 7737 55400 10737 55600
rect 11137 55400 14137 55600
rect 0 54000 15000 55400
rect 937 53800 3937 54000
rect 4337 53800 7337 54000
rect 7737 53800 10737 54000
rect 11137 53800 14137 54000
rect 0 52400 15000 53800
rect 0 50800 15000 52200
rect 0 49200 15000 50600
rect 0 46000 15000 49000
rect 0 42800 15000 45800
rect 937 42600 3937 42800
rect 4337 42600 7337 42800
rect 7737 42600 10737 42800
rect 11137 42600 14137 42800
rect 0 41200 15000 42600
rect 0 39600 15000 41000
rect 0 36400 15000 39400
rect 937 36200 3937 36400
rect 4337 36200 7337 36400
rect 7737 36200 10737 36400
rect 11137 36200 14137 36400
rect 0 33200 15000 36200
rect 937 33000 3937 33200
rect 4337 33000 7337 33200
rect 7737 33000 10737 33200
rect 11137 33000 14137 33200
rect 0 30000 15000 33000
rect 937 29800 3937 30000
rect 4337 29800 7337 30000
rect 7737 29800 10737 30000
rect 11137 29800 14137 30000
rect 0 26800 15000 29800
rect 0 25200 15000 26600
rect 0 23600 15000 25000
rect 0 20400 15000 23400
rect 937 20200 3937 20400
rect 4337 20200 7337 20400
rect 7737 20200 10737 20400
rect 11137 20200 14137 20400
rect 0 17200 15000 20200
rect 937 17000 3937 17200
rect 4337 17000 7337 17200
rect 7737 17000 10737 17200
rect 11137 17000 14137 17200
rect 0 14000 15000 17000
use M1_PSUB_CDNS_40661956134176  M1_PSUB_CDNS_40661956134176_0
timestamp 1698431365
transform 1 0 14952 0 1 41524
box 0 0 1 1
use M1_PSUB_CDNS_40661956134176  M1_PSUB_CDNS_40661956134176_1
timestamp 1698431365
transform 1 0 48 0 1 41524
box 0 0 1 1
use M1_PSUB_CDNS_40661956134192  M1_PSUB_CDNS_40661956134192_0
timestamp 1698431365
transform 1 0 7533 0 1 13192
box 0 0 1 1
use M1_PSUB_CDNS_40661956134192  M1_PSUB_CDNS_40661956134192_1
timestamp 1698431365
transform 1 0 7533 0 1 69873
box 0 0 1 1
<< labels >>
rlabel metal3 s 763 15661 763 15661 4 DVSS
port 1 nsew
rlabel metal3 s 716 18832 716 18832 4 DVSS
port 1 nsew
rlabel metal3 s 785 21818 785 21818 4 DVSS
port 1 nsew
rlabel metal3 s 785 49934 785 49934 4 VSS
port 2 nsew
rlabel metal3 s 785 64169 785 64169 4 VSS
port 2 nsew
rlabel metal3 s 785 62734 785 62734 4 VDD
port 3 nsew
rlabel metal3 s 785 51369 785 51369 4 VDD
port 3 nsew
rlabel metal3 s 785 68960 785 68960 4 DVSS
port 1 nsew
rlabel metal3 s 785 65934 785 65934 4 DVSS
port 1 nsew
rlabel metal3 s 785 60969 785 60969 4 DVSS
port 1 nsew
rlabel metal3 s 785 57769 785 57769 4 DVSS
port 1 nsew
rlabel metal3 s 785 26011 785 26011 4 DVSS
port 1 nsew
rlabel metal3 s 785 47506 785 47506 4 DVSS
port 1 nsew
rlabel metal3 s 785 40253 785 40253 4 DVSS
port 1 nsew
rlabel metal3 s 785 59534 785 59534 4 DVDD
port 4 nsew
rlabel metal3 s 785 53134 785 53134 4 DVDD
port 4 nsew
rlabel metal3 s 785 54569 785 54569 4 DVDD
port 4 nsew
rlabel metal3 s 785 56334 785 56334 4 DVDD
port 4 nsew
rlabel metal3 s 785 44279 785 44279 4 DVDD
port 4 nsew
rlabel metal3 s 785 41888 785 41888 4 DVDD
port 4 nsew
rlabel metal3 s 785 37870 785 37870 4 DVDD
port 4 nsew
rlabel metal3 s 785 34634 785 34634 4 DVDD
port 4 nsew
rlabel metal3 s 785 31520 785 31520 4 DVDD
port 4 nsew
rlabel metal3 s 785 28305 785 28305 4 DVDD
port 4 nsew
rlabel metal3 s 785 24195 785 24195 4 DVDD
port 4 nsew
rlabel metal3 s 785 67369 785 67369 4 DVDD
port 4 nsew
<< properties >>
string FIXED_BBOX 0 13097 15000 70000
string GDS_END 61768
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 55844
<< end >>
