magic
tech gf180mcuD
magscale 1 10
timestamp 1698431365
<< metal1 >>
rect 3621 37081 3945 37093
rect 3621 37029 3633 37081
rect 3685 37029 3757 37081
rect 3809 37029 3881 37081
rect 3933 37029 3945 37081
rect 3621 36957 3945 37029
rect 3621 36905 3633 36957
rect 3685 36905 3757 36957
rect 3809 36905 3881 36957
rect 3933 36905 3945 36957
rect 3621 36833 3945 36905
rect 3621 36781 3633 36833
rect 3685 36781 3757 36833
rect 3809 36781 3881 36833
rect 3933 36781 3945 36833
rect 3621 36709 3945 36781
rect 3621 36657 3633 36709
rect 3685 36657 3757 36709
rect 3809 36657 3881 36709
rect 3933 36657 3945 36709
rect 3621 36585 3945 36657
rect 3621 36533 3633 36585
rect 3685 36533 3757 36585
rect 3809 36533 3881 36585
rect 3933 36533 3945 36585
rect 3621 36461 3945 36533
rect 3621 36409 3633 36461
rect 3685 36409 3757 36461
rect 3809 36409 3881 36461
rect 3933 36409 3945 36461
rect 3621 36397 3945 36409
rect 3621 30157 3945 30169
rect 3621 30105 3633 30157
rect 3685 30105 3757 30157
rect 3809 30105 3881 30157
rect 3933 30105 3945 30157
rect 3621 30033 3945 30105
rect 3621 29981 3633 30033
rect 3685 29981 3757 30033
rect 3809 29981 3881 30033
rect 3933 29981 3945 30033
rect 3621 29909 3945 29981
rect 3621 29857 3633 29909
rect 3685 29857 3757 29909
rect 3809 29857 3881 29909
rect 3933 29857 3945 29909
rect 3621 29785 3945 29857
rect 3621 29733 3633 29785
rect 3685 29733 3757 29785
rect 3809 29733 3881 29785
rect 3933 29733 3945 29785
rect 3621 29661 3945 29733
rect 3621 29609 3633 29661
rect 3685 29609 3757 29661
rect 3809 29609 3881 29661
rect 3933 29609 3945 29661
rect 3621 29537 3945 29609
rect 3621 29485 3633 29537
rect 3685 29485 3757 29537
rect 3809 29485 3881 29537
rect 3933 29485 3945 29537
rect 3621 29413 3945 29485
rect 3621 29361 3633 29413
rect 3685 29361 3757 29413
rect 3809 29361 3881 29413
rect 3933 29361 3945 29413
rect 3621 29289 3945 29361
rect 3621 29237 3633 29289
rect 3685 29237 3757 29289
rect 3809 29237 3881 29289
rect 3933 29237 3945 29289
rect 3621 29165 3945 29237
rect 3621 29113 3633 29165
rect 3685 29113 3757 29165
rect 3809 29113 3881 29165
rect 3933 29113 3945 29165
rect 3621 29041 3945 29113
rect 3621 28989 3633 29041
rect 3685 28989 3757 29041
rect 3809 28989 3881 29041
rect 3933 28989 3945 29041
rect 3621 28917 3945 28989
rect 3621 28865 3633 28917
rect 3685 28865 3757 28917
rect 3809 28865 3881 28917
rect 3933 28903 3945 28917
rect 3933 28865 6188 28903
rect 3621 28793 6188 28865
rect 3621 28741 3633 28793
rect 3685 28741 3757 28793
rect 3809 28741 3881 28793
rect 3933 28769 6188 28793
rect 3933 28741 3945 28769
rect 3621 28669 3945 28741
rect 3621 28617 3633 28669
rect 3685 28617 3757 28669
rect 3809 28617 3881 28669
rect 3933 28617 3945 28669
rect 3621 28545 3945 28617
rect 3621 28493 3633 28545
rect 3685 28493 3757 28545
rect 3809 28493 3881 28545
rect 3933 28493 3945 28545
rect 3621 28421 3945 28493
rect 3621 28369 3633 28421
rect 3685 28369 3757 28421
rect 3809 28369 3881 28421
rect 3933 28369 3945 28421
rect 3621 28357 3945 28369
rect 3621 24062 3945 24074
rect 3621 24010 3633 24062
rect 3685 24010 3757 24062
rect 3809 24010 3881 24062
rect 3933 24010 3945 24062
rect 3621 23938 3945 24010
rect 3621 23886 3633 23938
rect 3685 23886 3757 23938
rect 3809 23886 3881 23938
rect 3933 23886 3945 23938
rect 3621 23868 3945 23886
rect 3621 23814 5873 23868
rect 3621 23762 3633 23814
rect 3685 23762 3757 23814
rect 3809 23762 3881 23814
rect 3933 23762 5873 23814
rect 3621 23690 5873 23762
rect 3621 23638 3633 23690
rect 3685 23638 3757 23690
rect 3809 23638 3881 23690
rect 3933 23673 5873 23690
rect 3933 23638 3945 23673
rect 3621 23566 3945 23638
rect 3621 23514 3633 23566
rect 3685 23514 3757 23566
rect 3809 23514 3881 23566
rect 3933 23514 3945 23566
rect 3621 23442 3945 23514
rect 3621 23390 3633 23442
rect 3685 23390 3757 23442
rect 3809 23390 3881 23442
rect 3933 23390 3945 23442
rect 3621 23318 3945 23390
rect 3621 23266 3633 23318
rect 3685 23266 3757 23318
rect 3809 23266 3881 23318
rect 3933 23266 3945 23318
rect 3621 23194 3945 23266
rect 3621 23142 3633 23194
rect 3685 23142 3757 23194
rect 3809 23142 3881 23194
rect 3933 23142 3945 23194
rect 3621 23130 3945 23142
rect 3621 19505 3945 19517
rect 3621 19453 3633 19505
rect 3685 19453 3757 19505
rect 3809 19453 3881 19505
rect 3933 19453 3945 19505
rect 3621 19381 3945 19453
rect 3621 19329 3633 19381
rect 3685 19329 3757 19381
rect 3809 19329 3881 19381
rect 3933 19329 3945 19381
rect 3621 19257 3945 19329
rect 3621 19205 3633 19257
rect 3685 19205 3757 19257
rect 3809 19205 3881 19257
rect 3933 19205 3945 19257
rect 3621 19133 3945 19205
rect 3621 19081 3633 19133
rect 3685 19081 3757 19133
rect 3809 19081 3881 19133
rect 3933 19081 3945 19133
rect 3621 19009 3945 19081
rect 3621 18957 3633 19009
rect 3685 18957 3757 19009
rect 3809 18957 3881 19009
rect 3933 18957 3945 19009
rect 3621 18885 3945 18957
rect 3621 18833 3633 18885
rect 3685 18833 3757 18885
rect 3809 18833 3881 18885
rect 3933 18833 3945 18885
rect 3621 18761 3945 18833
rect 3621 18709 3633 18761
rect 3685 18709 3757 18761
rect 3809 18709 3881 18761
rect 3933 18709 3945 18761
rect 3621 18637 3945 18709
rect 3621 18585 3633 18637
rect 3685 18585 3757 18637
rect 3809 18585 3881 18637
rect 3933 18585 3945 18637
rect 3621 18513 3945 18585
rect 3621 18461 3633 18513
rect 3685 18461 3757 18513
rect 3809 18461 3881 18513
rect 3933 18461 3945 18513
rect 3621 18389 3945 18461
rect 3621 18337 3633 18389
rect 3685 18337 3757 18389
rect 3809 18337 3881 18389
rect 3933 18337 3945 18389
rect 3621 18265 3945 18337
rect 3621 18213 3633 18265
rect 3685 18213 3757 18265
rect 3809 18213 3881 18265
rect 3933 18213 3945 18265
rect 3621 18141 3945 18213
rect 3621 18089 3633 18141
rect 3685 18089 3757 18141
rect 3809 18089 3881 18141
rect 3933 18089 3945 18141
rect 3621 18017 3945 18089
rect 3621 17965 3633 18017
rect 3685 17965 3757 18017
rect 3809 17965 3881 18017
rect 3933 17965 3945 18017
rect 3621 17893 3945 17965
rect 3621 17841 3633 17893
rect 3685 17841 3757 17893
rect 3809 17841 3881 17893
rect 3933 17841 3945 17893
rect 3621 17769 3945 17841
rect 3621 17717 3633 17769
rect 3685 17717 3757 17769
rect 3809 17717 3881 17769
rect 3933 17717 3945 17769
rect 3621 17645 3945 17717
rect 3621 17593 3633 17645
rect 3685 17593 3757 17645
rect 3809 17593 3881 17645
rect 3933 17593 3945 17645
rect 3621 17521 3945 17593
rect 3621 17469 3633 17521
rect 3685 17469 3757 17521
rect 3809 17469 3881 17521
rect 3933 17469 3945 17521
rect 3621 17397 3945 17469
rect 3621 17345 3633 17397
rect 3685 17345 3757 17397
rect 3809 17345 3881 17397
rect 3933 17345 3945 17397
rect 3621 17273 3945 17345
rect 3621 17221 3633 17273
rect 3685 17221 3757 17273
rect 3809 17221 3881 17273
rect 3933 17221 3945 17273
rect 3621 17149 3945 17221
rect 3621 17097 3633 17149
rect 3685 17097 3757 17149
rect 3809 17097 3881 17149
rect 3933 17097 3945 17149
rect 3621 17025 3945 17097
rect 3621 16973 3633 17025
rect 3685 16973 3757 17025
rect 3809 16973 3881 17025
rect 3933 16973 3945 17025
rect 3621 16901 3945 16973
rect 3621 16849 3633 16901
rect 3685 16849 3757 16901
rect 3809 16849 3881 16901
rect 3933 16849 3945 16901
rect 3621 16777 3945 16849
rect 3621 16725 3633 16777
rect 3685 16725 3757 16777
rect 3809 16725 3881 16777
rect 3933 16725 3945 16777
rect 3621 16653 3945 16725
rect 3621 16601 3633 16653
rect 3685 16601 3757 16653
rect 3809 16601 3881 16653
rect 3933 16601 3945 16653
rect 3621 16529 3945 16601
rect 3621 16477 3633 16529
rect 3685 16477 3757 16529
rect 3809 16477 3881 16529
rect 3933 16477 3945 16529
rect 3621 16405 3945 16477
rect 3621 16353 3633 16405
rect 3685 16353 3757 16405
rect 3809 16353 3881 16405
rect 3933 16353 3945 16405
rect 3621 16281 3945 16353
rect 3621 16229 3633 16281
rect 3685 16229 3757 16281
rect 3809 16229 3881 16281
rect 3933 16229 3945 16281
rect 3621 16217 3945 16229
rect 3621 13226 3945 13238
rect 3621 13174 3633 13226
rect 3685 13174 3757 13226
rect 3809 13174 3881 13226
rect 3933 13174 3945 13226
rect 3621 13102 3945 13174
rect 3621 13050 3633 13102
rect 3685 13050 3757 13102
rect 3809 13050 3881 13102
rect 3933 13050 3945 13102
rect 3621 12978 3945 13050
rect 3621 12926 3633 12978
rect 3685 12926 3757 12978
rect 3809 12926 3881 12978
rect 3933 12926 3945 12978
rect 3621 12854 3945 12926
rect 3621 12802 3633 12854
rect 3685 12802 3757 12854
rect 3809 12802 3881 12854
rect 3933 12802 3945 12854
rect 3621 12730 3945 12802
rect 3621 12678 3633 12730
rect 3685 12678 3757 12730
rect 3809 12678 3881 12730
rect 3933 12678 3945 12730
rect 3621 12606 3945 12678
rect 3621 12554 3633 12606
rect 3685 12554 3757 12606
rect 3809 12554 3881 12606
rect 3933 12554 3945 12606
rect 3621 12482 3945 12554
rect 3621 12430 3633 12482
rect 3685 12430 3757 12482
rect 3809 12430 3881 12482
rect 3933 12430 3945 12482
rect 3621 12358 3945 12430
rect 3621 12306 3633 12358
rect 3685 12306 3757 12358
rect 3809 12306 3881 12358
rect 3933 12306 3945 12358
rect 3621 12234 3945 12306
rect 3621 12182 3633 12234
rect 3685 12182 3757 12234
rect 3809 12182 3881 12234
rect 3933 12182 3945 12234
rect 3621 12110 3945 12182
rect 3621 12058 3633 12110
rect 3685 12058 3757 12110
rect 3809 12058 3881 12110
rect 3933 12058 3945 12110
rect 3621 12046 3945 12058
rect 3621 9390 3945 9402
rect 3621 9338 3633 9390
rect 3685 9338 3757 9390
rect 3809 9338 3881 9390
rect 3933 9338 3945 9390
rect 3621 9266 3945 9338
rect 3621 9214 3633 9266
rect 3685 9214 3757 9266
rect 3809 9214 3881 9266
rect 3933 9214 3945 9266
rect 3621 9142 3945 9214
rect 3621 9090 3633 9142
rect 3685 9090 3757 9142
rect 3809 9090 3881 9142
rect 3933 9090 3945 9142
rect 3621 9018 3945 9090
rect 3621 8966 3633 9018
rect 3685 8966 3757 9018
rect 3809 8966 3881 9018
rect 3933 8966 3945 9018
rect 3621 8894 3945 8966
rect 3621 8842 3633 8894
rect 3685 8842 3757 8894
rect 3809 8842 3881 8894
rect 3933 8842 3945 8894
rect 3621 8770 3945 8842
rect 3621 8718 3633 8770
rect 3685 8718 3757 8770
rect 3809 8718 3881 8770
rect 3933 8718 3945 8770
rect 3621 8646 3945 8718
rect 3621 8594 3633 8646
rect 3685 8594 3757 8646
rect 3809 8594 3881 8646
rect 3933 8594 3945 8646
rect 3621 8522 3945 8594
rect 3621 8470 3633 8522
rect 3685 8470 3757 8522
rect 3809 8470 3881 8522
rect 3933 8470 3945 8522
rect 3621 8398 3945 8470
rect 3621 8346 3633 8398
rect 3685 8346 3757 8398
rect 3809 8346 3881 8398
rect 3933 8346 3945 8398
rect 3621 8274 3945 8346
rect 3621 8222 3633 8274
rect 3685 8222 3757 8274
rect 3809 8222 3881 8274
rect 3933 8222 3945 8274
rect 3621 8150 3945 8222
rect 3621 8098 3633 8150
rect 3685 8098 3757 8150
rect 3809 8098 3881 8150
rect 3933 8098 3945 8150
rect 3621 8026 3945 8098
rect 3621 7974 3633 8026
rect 3685 7974 3757 8026
rect 3809 7974 3881 8026
rect 3933 7974 3945 8026
rect 3621 7902 3945 7974
rect 3621 7850 3633 7902
rect 3685 7850 3757 7902
rect 3809 7850 3881 7902
rect 3933 7850 3945 7902
rect 3621 7778 3945 7850
rect 3621 7726 3633 7778
rect 3685 7726 3757 7778
rect 3809 7726 3881 7778
rect 3933 7726 3945 7778
rect 3621 7654 3945 7726
rect 3621 7602 3633 7654
rect 3685 7602 3757 7654
rect 3809 7602 3881 7654
rect 3933 7602 3945 7654
rect 3621 7590 3945 7602
rect 3621 5526 3945 5538
rect 3621 5474 3633 5526
rect 3685 5474 3757 5526
rect 3809 5474 3881 5526
rect 3933 5474 3945 5526
rect 3621 5402 3945 5474
rect 3621 5350 3633 5402
rect 3685 5350 3757 5402
rect 3809 5350 3881 5402
rect 3933 5350 3945 5402
rect 3621 5278 3945 5350
rect 3621 5226 3633 5278
rect 3685 5226 3757 5278
rect 3809 5226 3881 5278
rect 3933 5226 3945 5278
rect 3621 5154 3945 5226
rect 3621 5102 3633 5154
rect 3685 5102 3757 5154
rect 3809 5102 3881 5154
rect 3933 5102 3945 5154
rect 3621 5030 3945 5102
rect 3621 4978 3633 5030
rect 3685 4978 3757 5030
rect 3809 4978 3881 5030
rect 3933 4978 3945 5030
rect 3621 4906 3945 4978
rect 3621 4854 3633 4906
rect 3685 4854 3757 4906
rect 3809 4854 3881 4906
rect 3933 4854 3945 4906
rect 3621 4782 3945 4854
rect 3621 4730 3633 4782
rect 3685 4730 3757 4782
rect 3809 4730 3881 4782
rect 3933 4730 3945 4782
rect 3621 4658 3945 4730
rect 3621 4606 3633 4658
rect 3685 4606 3757 4658
rect 3809 4606 3881 4658
rect 3933 4606 3945 4658
rect 3621 4534 3945 4606
rect 3621 4482 3633 4534
rect 3685 4482 3757 4534
rect 3809 4482 3881 4534
rect 3933 4482 3945 4534
rect 3621 4410 3945 4482
rect 3621 4358 3633 4410
rect 3685 4358 3757 4410
rect 3809 4358 3881 4410
rect 3933 4358 3945 4410
rect 3621 4346 3945 4358
<< via1 >>
rect 3633 37029 3685 37081
rect 3757 37029 3809 37081
rect 3881 37029 3933 37081
rect 3633 36905 3685 36957
rect 3757 36905 3809 36957
rect 3881 36905 3933 36957
rect 3633 36781 3685 36833
rect 3757 36781 3809 36833
rect 3881 36781 3933 36833
rect 3633 36657 3685 36709
rect 3757 36657 3809 36709
rect 3881 36657 3933 36709
rect 3633 36533 3685 36585
rect 3757 36533 3809 36585
rect 3881 36533 3933 36585
rect 3633 36409 3685 36461
rect 3757 36409 3809 36461
rect 3881 36409 3933 36461
rect 3633 30105 3685 30157
rect 3757 30105 3809 30157
rect 3881 30105 3933 30157
rect 3633 29981 3685 30033
rect 3757 29981 3809 30033
rect 3881 29981 3933 30033
rect 3633 29857 3685 29909
rect 3757 29857 3809 29909
rect 3881 29857 3933 29909
rect 3633 29733 3685 29785
rect 3757 29733 3809 29785
rect 3881 29733 3933 29785
rect 3633 29609 3685 29661
rect 3757 29609 3809 29661
rect 3881 29609 3933 29661
rect 3633 29485 3685 29537
rect 3757 29485 3809 29537
rect 3881 29485 3933 29537
rect 3633 29361 3685 29413
rect 3757 29361 3809 29413
rect 3881 29361 3933 29413
rect 3633 29237 3685 29289
rect 3757 29237 3809 29289
rect 3881 29237 3933 29289
rect 3633 29113 3685 29165
rect 3757 29113 3809 29165
rect 3881 29113 3933 29165
rect 3633 28989 3685 29041
rect 3757 28989 3809 29041
rect 3881 28989 3933 29041
rect 3633 28865 3685 28917
rect 3757 28865 3809 28917
rect 3881 28865 3933 28917
rect 3633 28741 3685 28793
rect 3757 28741 3809 28793
rect 3881 28741 3933 28793
rect 3633 28617 3685 28669
rect 3757 28617 3809 28669
rect 3881 28617 3933 28669
rect 3633 28493 3685 28545
rect 3757 28493 3809 28545
rect 3881 28493 3933 28545
rect 3633 28369 3685 28421
rect 3757 28369 3809 28421
rect 3881 28369 3933 28421
rect 3633 24010 3685 24062
rect 3757 24010 3809 24062
rect 3881 24010 3933 24062
rect 3633 23886 3685 23938
rect 3757 23886 3809 23938
rect 3881 23886 3933 23938
rect 3633 23762 3685 23814
rect 3757 23762 3809 23814
rect 3881 23762 3933 23814
rect 3633 23638 3685 23690
rect 3757 23638 3809 23690
rect 3881 23638 3933 23690
rect 3633 23514 3685 23566
rect 3757 23514 3809 23566
rect 3881 23514 3933 23566
rect 3633 23390 3685 23442
rect 3757 23390 3809 23442
rect 3881 23390 3933 23442
rect 3633 23266 3685 23318
rect 3757 23266 3809 23318
rect 3881 23266 3933 23318
rect 3633 23142 3685 23194
rect 3757 23142 3809 23194
rect 3881 23142 3933 23194
rect 3633 19453 3685 19505
rect 3757 19453 3809 19505
rect 3881 19453 3933 19505
rect 3633 19329 3685 19381
rect 3757 19329 3809 19381
rect 3881 19329 3933 19381
rect 3633 19205 3685 19257
rect 3757 19205 3809 19257
rect 3881 19205 3933 19257
rect 3633 19081 3685 19133
rect 3757 19081 3809 19133
rect 3881 19081 3933 19133
rect 3633 18957 3685 19009
rect 3757 18957 3809 19009
rect 3881 18957 3933 19009
rect 3633 18833 3685 18885
rect 3757 18833 3809 18885
rect 3881 18833 3933 18885
rect 3633 18709 3685 18761
rect 3757 18709 3809 18761
rect 3881 18709 3933 18761
rect 3633 18585 3685 18637
rect 3757 18585 3809 18637
rect 3881 18585 3933 18637
rect 3633 18461 3685 18513
rect 3757 18461 3809 18513
rect 3881 18461 3933 18513
rect 3633 18337 3685 18389
rect 3757 18337 3809 18389
rect 3881 18337 3933 18389
rect 3633 18213 3685 18265
rect 3757 18213 3809 18265
rect 3881 18213 3933 18265
rect 3633 18089 3685 18141
rect 3757 18089 3809 18141
rect 3881 18089 3933 18141
rect 3633 17965 3685 18017
rect 3757 17965 3809 18017
rect 3881 17965 3933 18017
rect 3633 17841 3685 17893
rect 3757 17841 3809 17893
rect 3881 17841 3933 17893
rect 3633 17717 3685 17769
rect 3757 17717 3809 17769
rect 3881 17717 3933 17769
rect 3633 17593 3685 17645
rect 3757 17593 3809 17645
rect 3881 17593 3933 17645
rect 3633 17469 3685 17521
rect 3757 17469 3809 17521
rect 3881 17469 3933 17521
rect 3633 17345 3685 17397
rect 3757 17345 3809 17397
rect 3881 17345 3933 17397
rect 3633 17221 3685 17273
rect 3757 17221 3809 17273
rect 3881 17221 3933 17273
rect 3633 17097 3685 17149
rect 3757 17097 3809 17149
rect 3881 17097 3933 17149
rect 3633 16973 3685 17025
rect 3757 16973 3809 17025
rect 3881 16973 3933 17025
rect 3633 16849 3685 16901
rect 3757 16849 3809 16901
rect 3881 16849 3933 16901
rect 3633 16725 3685 16777
rect 3757 16725 3809 16777
rect 3881 16725 3933 16777
rect 3633 16601 3685 16653
rect 3757 16601 3809 16653
rect 3881 16601 3933 16653
rect 3633 16477 3685 16529
rect 3757 16477 3809 16529
rect 3881 16477 3933 16529
rect 3633 16353 3685 16405
rect 3757 16353 3809 16405
rect 3881 16353 3933 16405
rect 3633 16229 3685 16281
rect 3757 16229 3809 16281
rect 3881 16229 3933 16281
rect 3633 13174 3685 13226
rect 3757 13174 3809 13226
rect 3881 13174 3933 13226
rect 3633 13050 3685 13102
rect 3757 13050 3809 13102
rect 3881 13050 3933 13102
rect 3633 12926 3685 12978
rect 3757 12926 3809 12978
rect 3881 12926 3933 12978
rect 3633 12802 3685 12854
rect 3757 12802 3809 12854
rect 3881 12802 3933 12854
rect 3633 12678 3685 12730
rect 3757 12678 3809 12730
rect 3881 12678 3933 12730
rect 3633 12554 3685 12606
rect 3757 12554 3809 12606
rect 3881 12554 3933 12606
rect 3633 12430 3685 12482
rect 3757 12430 3809 12482
rect 3881 12430 3933 12482
rect 3633 12306 3685 12358
rect 3757 12306 3809 12358
rect 3881 12306 3933 12358
rect 3633 12182 3685 12234
rect 3757 12182 3809 12234
rect 3881 12182 3933 12234
rect 3633 12058 3685 12110
rect 3757 12058 3809 12110
rect 3881 12058 3933 12110
rect 3633 9338 3685 9390
rect 3757 9338 3809 9390
rect 3881 9338 3933 9390
rect 3633 9214 3685 9266
rect 3757 9214 3809 9266
rect 3881 9214 3933 9266
rect 3633 9090 3685 9142
rect 3757 9090 3809 9142
rect 3881 9090 3933 9142
rect 3633 8966 3685 9018
rect 3757 8966 3809 9018
rect 3881 8966 3933 9018
rect 3633 8842 3685 8894
rect 3757 8842 3809 8894
rect 3881 8842 3933 8894
rect 3633 8718 3685 8770
rect 3757 8718 3809 8770
rect 3881 8718 3933 8770
rect 3633 8594 3685 8646
rect 3757 8594 3809 8646
rect 3881 8594 3933 8646
rect 3633 8470 3685 8522
rect 3757 8470 3809 8522
rect 3881 8470 3933 8522
rect 3633 8346 3685 8398
rect 3757 8346 3809 8398
rect 3881 8346 3933 8398
rect 3633 8222 3685 8274
rect 3757 8222 3809 8274
rect 3881 8222 3933 8274
rect 3633 8098 3685 8150
rect 3757 8098 3809 8150
rect 3881 8098 3933 8150
rect 3633 7974 3685 8026
rect 3757 7974 3809 8026
rect 3881 7974 3933 8026
rect 3633 7850 3685 7902
rect 3757 7850 3809 7902
rect 3881 7850 3933 7902
rect 3633 7726 3685 7778
rect 3757 7726 3809 7778
rect 3881 7726 3933 7778
rect 3633 7602 3685 7654
rect 3757 7602 3809 7654
rect 3881 7602 3933 7654
rect 3633 5474 3685 5526
rect 3757 5474 3809 5526
rect 3881 5474 3933 5526
rect 3633 5350 3685 5402
rect 3757 5350 3809 5402
rect 3881 5350 3933 5402
rect 3633 5226 3685 5278
rect 3757 5226 3809 5278
rect 3881 5226 3933 5278
rect 3633 5102 3685 5154
rect 3757 5102 3809 5154
rect 3881 5102 3933 5154
rect 3633 4978 3685 5030
rect 3757 4978 3809 5030
rect 3881 4978 3933 5030
rect 3633 4854 3685 4906
rect 3757 4854 3809 4906
rect 3881 4854 3933 4906
rect 3633 4730 3685 4782
rect 3757 4730 3809 4782
rect 3881 4730 3933 4782
rect 3633 4606 3685 4658
rect 3757 4606 3809 4658
rect 3881 4606 3933 4658
rect 3633 4482 3685 4534
rect 3757 4482 3809 4534
rect 3881 4482 3933 4534
rect 3633 4358 3685 4410
rect 3757 4358 3809 4410
rect 3881 4358 3933 4410
<< metal2 >>
rect 3621 37083 3945 37093
rect 3621 37027 3631 37083
rect 3687 37027 3755 37083
rect 3811 37027 3879 37083
rect 3935 37027 3945 37083
rect 3621 36959 3945 37027
rect 3621 36903 3631 36959
rect 3687 36903 3755 36959
rect 3811 36903 3879 36959
rect 3935 36903 3945 36959
rect 3621 36835 3945 36903
rect 3621 36779 3631 36835
rect 3687 36779 3755 36835
rect 3811 36779 3879 36835
rect 3935 36779 3945 36835
rect 3621 36711 3945 36779
rect 3621 36655 3631 36711
rect 3687 36655 3755 36711
rect 3811 36655 3879 36711
rect 3935 36655 3945 36711
rect 3621 36587 3945 36655
rect 3621 36531 3631 36587
rect 3687 36531 3755 36587
rect 3811 36531 3879 36587
rect 3935 36531 3945 36587
rect 3621 36463 3945 36531
rect 3621 36407 3631 36463
rect 3687 36407 3755 36463
rect 3811 36407 3879 36463
rect 3935 36407 3945 36463
rect 3621 36397 3945 36407
rect 4045 35929 5045 52645
rect 4045 35873 4095 35929
rect 4151 35873 4219 35929
rect 4275 35873 4343 35929
rect 4399 35873 4467 35929
rect 4523 35873 4591 35929
rect 4647 35873 4715 35929
rect 4771 35873 4839 35929
rect 4895 35873 4963 35929
rect 5019 35873 5045 35929
rect 4045 35805 5045 35873
rect 4045 35749 4095 35805
rect 4151 35749 4219 35805
rect 4275 35749 4343 35805
rect 4399 35749 4467 35805
rect 4523 35749 4591 35805
rect 4647 35749 4715 35805
rect 4771 35749 4839 35805
rect 4895 35749 4963 35805
rect 5019 35749 5045 35805
rect 4045 35681 5045 35749
rect 4045 35625 4095 35681
rect 4151 35625 4219 35681
rect 4275 35625 4343 35681
rect 4399 35625 4467 35681
rect 4523 35625 4591 35681
rect 4647 35625 4715 35681
rect 4771 35625 4839 35681
rect 4895 35625 4963 35681
rect 5019 35625 5045 35681
rect 4045 35557 5045 35625
rect 4045 35501 4095 35557
rect 4151 35501 4219 35557
rect 4275 35501 4343 35557
rect 4399 35501 4467 35557
rect 4523 35501 4591 35557
rect 4647 35501 4715 35557
rect 4771 35501 4839 35557
rect 4895 35501 4963 35557
rect 5019 35501 5045 35557
rect 4045 35433 5045 35501
rect 4045 35377 4095 35433
rect 4151 35377 4219 35433
rect 4275 35377 4343 35433
rect 4399 35377 4467 35433
rect 4523 35377 4591 35433
rect 4647 35377 4715 35433
rect 4771 35377 4839 35433
rect 4895 35377 4963 35433
rect 5019 35377 5045 35433
rect 4045 35309 5045 35377
rect 4045 35253 4095 35309
rect 4151 35253 4219 35309
rect 4275 35253 4343 35309
rect 4399 35253 4467 35309
rect 4523 35253 4591 35309
rect 4647 35253 4715 35309
rect 4771 35253 4839 35309
rect 4895 35253 4963 35309
rect 5019 35253 5045 35309
rect 4045 35185 5045 35253
rect 4045 35129 4095 35185
rect 4151 35129 4219 35185
rect 4275 35129 4343 35185
rect 4399 35129 4467 35185
rect 4523 35129 4591 35185
rect 4647 35129 4715 35185
rect 4771 35129 4839 35185
rect 4895 35129 4963 35185
rect 5019 35129 5045 35185
rect 4045 35061 5045 35129
rect 4045 35005 4095 35061
rect 4151 35005 4219 35061
rect 4275 35005 4343 35061
rect 4399 35005 4467 35061
rect 4523 35005 4591 35061
rect 4647 35005 4715 35061
rect 4771 35005 4839 35061
rect 4895 35005 4963 35061
rect 5019 35005 5045 35061
rect 4045 34937 5045 35005
rect 4045 34881 4095 34937
rect 4151 34881 4219 34937
rect 4275 34881 4343 34937
rect 4399 34881 4467 34937
rect 4523 34881 4591 34937
rect 4647 34881 4715 34937
rect 4771 34881 4839 34937
rect 4895 34881 4963 34937
rect 5019 34881 5045 34937
rect 4045 34813 5045 34881
rect 4045 34757 4095 34813
rect 4151 34757 4219 34813
rect 4275 34757 4343 34813
rect 4399 34757 4467 34813
rect 4523 34757 4591 34813
rect 4647 34757 4715 34813
rect 4771 34757 4839 34813
rect 4895 34757 4963 34813
rect 5019 34757 5045 34813
rect 4045 34689 5045 34757
rect 4045 34633 4095 34689
rect 4151 34633 4219 34689
rect 4275 34633 4343 34689
rect 4399 34633 4467 34689
rect 4523 34633 4591 34689
rect 4647 34633 4715 34689
rect 4771 34633 4839 34689
rect 4895 34633 4963 34689
rect 5019 34633 5045 34689
rect 4045 34565 5045 34633
rect 4045 34509 4095 34565
rect 4151 34509 4219 34565
rect 4275 34509 4343 34565
rect 4399 34509 4467 34565
rect 4523 34509 4591 34565
rect 4647 34509 4715 34565
rect 4771 34509 4839 34565
rect 4895 34509 4963 34565
rect 5019 34509 5045 34565
rect 4045 34441 5045 34509
rect 4045 34385 4095 34441
rect 4151 34385 4219 34441
rect 4275 34385 4343 34441
rect 4399 34385 4467 34441
rect 4523 34385 4591 34441
rect 4647 34385 4715 34441
rect 4771 34385 4839 34441
rect 4895 34385 4963 34441
rect 5019 34385 5045 34441
rect 4045 34317 5045 34385
rect 4045 34261 4095 34317
rect 4151 34261 4219 34317
rect 4275 34261 4343 34317
rect 4399 34261 4467 34317
rect 4523 34261 4591 34317
rect 4647 34261 4715 34317
rect 4771 34261 4839 34317
rect 4895 34261 4963 34317
rect 5019 34261 5045 34317
rect 4045 34193 5045 34261
rect 4045 34137 4095 34193
rect 4151 34137 4219 34193
rect 4275 34137 4343 34193
rect 4399 34137 4467 34193
rect 4523 34137 4591 34193
rect 4647 34137 4715 34193
rect 4771 34137 4839 34193
rect 4895 34137 4963 34193
rect 5019 34137 5045 34193
rect 4045 34069 5045 34137
rect 4045 34013 4095 34069
rect 4151 34013 4219 34069
rect 4275 34013 4343 34069
rect 4399 34013 4467 34069
rect 4523 34013 4591 34069
rect 4647 34013 4715 34069
rect 4771 34013 4839 34069
rect 4895 34013 4963 34069
rect 5019 34013 5045 34069
rect 4045 33945 5045 34013
rect 4045 33889 4095 33945
rect 4151 33889 4219 33945
rect 4275 33889 4343 33945
rect 4399 33889 4467 33945
rect 4523 33889 4591 33945
rect 4647 33889 4715 33945
rect 4771 33889 4839 33945
rect 4895 33889 4963 33945
rect 5019 33889 5045 33945
rect 4045 33821 5045 33889
rect 4045 33765 4095 33821
rect 4151 33765 4219 33821
rect 4275 33765 4343 33821
rect 4399 33765 4467 33821
rect 4523 33765 4591 33821
rect 4647 33765 4715 33821
rect 4771 33765 4839 33821
rect 4895 33765 4963 33821
rect 5019 33765 5045 33821
rect 4045 33697 5045 33765
rect 4045 33641 4095 33697
rect 4151 33641 4219 33697
rect 4275 33641 4343 33697
rect 4399 33641 4467 33697
rect 4523 33641 4591 33697
rect 4647 33641 4715 33697
rect 4771 33641 4839 33697
rect 4895 33641 4963 33697
rect 5019 33641 5045 33697
rect 4045 33573 5045 33641
rect 4045 33517 4095 33573
rect 4151 33517 4219 33573
rect 4275 33517 4343 33573
rect 4399 33517 4467 33573
rect 4523 33517 4591 33573
rect 4647 33517 4715 33573
rect 4771 33517 4839 33573
rect 4895 33517 4963 33573
rect 5019 33517 5045 33573
rect 4045 33449 5045 33517
rect 4045 33393 4095 33449
rect 4151 33393 4219 33449
rect 4275 33393 4343 33449
rect 4399 33393 4467 33449
rect 4523 33393 4591 33449
rect 4647 33393 4715 33449
rect 4771 33393 4839 33449
rect 4895 33393 4963 33449
rect 5019 33393 5045 33449
rect 4045 33325 5045 33393
rect 4045 33269 4095 33325
rect 4151 33269 4219 33325
rect 4275 33269 4343 33325
rect 4399 33269 4467 33325
rect 4523 33269 4591 33325
rect 4647 33269 4715 33325
rect 4771 33269 4839 33325
rect 4895 33269 4963 33325
rect 5019 33269 5045 33325
rect 4045 33201 5045 33269
rect 4045 33145 4095 33201
rect 4151 33145 4219 33201
rect 4275 33145 4343 33201
rect 4399 33145 4467 33201
rect 4523 33145 4591 33201
rect 4647 33145 4715 33201
rect 4771 33145 4839 33201
rect 4895 33145 4963 33201
rect 5019 33145 5045 33201
rect 4045 33077 5045 33145
rect 4045 33021 4095 33077
rect 4151 33021 4219 33077
rect 4275 33021 4343 33077
rect 4399 33021 4467 33077
rect 4523 33021 4591 33077
rect 4647 33021 4715 33077
rect 4771 33021 4839 33077
rect 4895 33021 4963 33077
rect 5019 33021 5045 33077
rect 4045 32953 5045 33021
rect 4045 32897 4095 32953
rect 4151 32897 4219 32953
rect 4275 32897 4343 32953
rect 4399 32897 4467 32953
rect 4523 32897 4591 32953
rect 4647 32897 4715 32953
rect 4771 32897 4839 32953
rect 4895 32897 4963 32953
rect 5019 32897 5045 32953
rect 4045 32829 5045 32897
rect 4045 32773 4095 32829
rect 4151 32773 4219 32829
rect 4275 32773 4343 32829
rect 4399 32773 4467 32829
rect 4523 32773 4591 32829
rect 4647 32773 4715 32829
rect 4771 32773 4839 32829
rect 4895 32773 4963 32829
rect 5019 32773 5045 32829
rect 4045 32705 5045 32773
rect 4045 32649 4095 32705
rect 4151 32649 4219 32705
rect 4275 32649 4343 32705
rect 4399 32649 4467 32705
rect 4523 32649 4591 32705
rect 4647 32649 4715 32705
rect 4771 32649 4839 32705
rect 4895 32649 4963 32705
rect 5019 32649 5045 32705
rect 4045 32581 5045 32649
rect 4045 32525 4095 32581
rect 4151 32525 4219 32581
rect 4275 32525 4343 32581
rect 4399 32525 4467 32581
rect 4523 32525 4591 32581
rect 4647 32525 4715 32581
rect 4771 32525 4839 32581
rect 4895 32525 4963 32581
rect 5019 32525 5045 32581
rect 4045 32457 5045 32525
rect 4045 32401 4095 32457
rect 4151 32401 4219 32457
rect 4275 32401 4343 32457
rect 4399 32401 4467 32457
rect 4523 32401 4591 32457
rect 4647 32401 4715 32457
rect 4771 32401 4839 32457
rect 4895 32401 4963 32457
rect 5019 32401 5045 32457
rect 4045 32333 5045 32401
rect 4045 32277 4095 32333
rect 4151 32277 4219 32333
rect 4275 32277 4343 32333
rect 4399 32277 4467 32333
rect 4523 32277 4591 32333
rect 4647 32277 4715 32333
rect 4771 32277 4839 32333
rect 4895 32277 4963 32333
rect 5019 32277 5045 32333
rect 4045 32209 5045 32277
rect 4045 32153 4095 32209
rect 4151 32153 4219 32209
rect 4275 32153 4343 32209
rect 4399 32153 4467 32209
rect 4523 32153 4591 32209
rect 4647 32153 4715 32209
rect 4771 32153 4839 32209
rect 4895 32153 4963 32209
rect 5019 32153 5045 32209
rect 4045 32085 5045 32153
rect 4045 32029 4095 32085
rect 4151 32029 4219 32085
rect 4275 32029 4343 32085
rect 4399 32029 4467 32085
rect 4523 32029 4591 32085
rect 4647 32029 4715 32085
rect 4771 32029 4839 32085
rect 4895 32029 4963 32085
rect 5019 32029 5045 32085
rect 4045 31961 5045 32029
rect 4045 31905 4095 31961
rect 4151 31905 4219 31961
rect 4275 31905 4343 31961
rect 4399 31905 4467 31961
rect 4523 31905 4591 31961
rect 4647 31905 4715 31961
rect 4771 31905 4839 31961
rect 4895 31905 4963 31961
rect 5019 31905 5045 31961
rect 4045 31837 5045 31905
rect 4045 31781 4095 31837
rect 4151 31781 4219 31837
rect 4275 31781 4343 31837
rect 4399 31781 4467 31837
rect 4523 31781 4591 31837
rect 4647 31781 4715 31837
rect 4771 31781 4839 31837
rect 4895 31781 4963 31837
rect 5019 31781 5045 31837
rect 4045 31713 5045 31781
rect 4045 31657 4095 31713
rect 4151 31657 4219 31713
rect 4275 31657 4343 31713
rect 4399 31657 4467 31713
rect 4523 31657 4591 31713
rect 4647 31657 4715 31713
rect 4771 31657 4839 31713
rect 4895 31657 4963 31713
rect 5019 31657 5045 31713
rect 4045 31589 5045 31657
rect 4045 31533 4095 31589
rect 4151 31533 4219 31589
rect 4275 31533 4343 31589
rect 4399 31533 4467 31589
rect 4523 31533 4591 31589
rect 4647 31533 4715 31589
rect 4771 31533 4839 31589
rect 4895 31533 4963 31589
rect 5019 31533 5045 31589
rect 4045 31465 5045 31533
rect 4045 31409 4095 31465
rect 4151 31409 4219 31465
rect 4275 31409 4343 31465
rect 4399 31409 4467 31465
rect 4523 31409 4591 31465
rect 4647 31409 4715 31465
rect 4771 31409 4839 31465
rect 4895 31409 4963 31465
rect 5019 31409 5045 31465
rect 4045 31341 5045 31409
rect 4045 31285 4095 31341
rect 4151 31285 4219 31341
rect 4275 31285 4343 31341
rect 4399 31285 4467 31341
rect 4523 31285 4591 31341
rect 4647 31285 4715 31341
rect 4771 31285 4839 31341
rect 4895 31285 4963 31341
rect 5019 31285 5045 31341
rect 3621 30159 3945 30169
rect 3621 30103 3631 30159
rect 3687 30103 3755 30159
rect 3811 30103 3879 30159
rect 3935 30103 3945 30159
rect 3621 30035 3945 30103
rect 3621 29979 3631 30035
rect 3687 29979 3755 30035
rect 3811 29979 3879 30035
rect 3935 29979 3945 30035
rect 3621 29911 3945 29979
rect 3621 29855 3631 29911
rect 3687 29855 3755 29911
rect 3811 29855 3879 29911
rect 3935 29855 3945 29911
rect 3621 29787 3945 29855
rect 3621 29731 3631 29787
rect 3687 29731 3755 29787
rect 3811 29731 3879 29787
rect 3935 29731 3945 29787
rect 3621 29663 3945 29731
rect 3621 29607 3631 29663
rect 3687 29607 3755 29663
rect 3811 29607 3879 29663
rect 3935 29607 3945 29663
rect 3621 29539 3945 29607
rect 3621 29483 3631 29539
rect 3687 29483 3755 29539
rect 3811 29483 3879 29539
rect 3935 29483 3945 29539
rect 3621 29415 3945 29483
rect 3621 29359 3631 29415
rect 3687 29359 3755 29415
rect 3811 29359 3879 29415
rect 3935 29359 3945 29415
rect 3621 29291 3945 29359
rect 3621 29235 3631 29291
rect 3687 29235 3755 29291
rect 3811 29235 3879 29291
rect 3935 29235 3945 29291
rect 3621 29167 3945 29235
rect 3621 29111 3631 29167
rect 3687 29111 3755 29167
rect 3811 29111 3879 29167
rect 3935 29111 3945 29167
rect 3621 29043 3945 29111
rect 3621 28987 3631 29043
rect 3687 28987 3755 29043
rect 3811 28987 3879 29043
rect 3935 28987 3945 29043
rect 3621 28919 3945 28987
rect 3621 28863 3631 28919
rect 3687 28863 3755 28919
rect 3811 28863 3879 28919
rect 3935 28863 3945 28919
rect 3621 28795 3945 28863
rect 3621 28739 3631 28795
rect 3687 28739 3755 28795
rect 3811 28739 3879 28795
rect 3935 28739 3945 28795
rect 3621 28671 3945 28739
rect 3621 28615 3631 28671
rect 3687 28615 3755 28671
rect 3811 28615 3879 28671
rect 3935 28615 3945 28671
rect 3621 28547 3945 28615
rect 3621 28491 3631 28547
rect 3687 28491 3755 28547
rect 3811 28491 3879 28547
rect 3935 28491 3945 28547
rect 3621 28423 3945 28491
rect 3621 28367 3631 28423
rect 3687 28367 3755 28423
rect 3811 28367 3879 28423
rect 3935 28367 3945 28423
rect 3621 28357 3945 28367
rect 4045 25691 5045 31285
rect 4045 25635 4095 25691
rect 4151 25635 4219 25691
rect 4275 25635 4343 25691
rect 4399 25635 4467 25691
rect 4523 25635 4591 25691
rect 4647 25635 4715 25691
rect 4771 25635 4839 25691
rect 4895 25635 4963 25691
rect 5019 25635 5045 25691
rect 4045 25567 5045 25635
rect 4045 25511 4095 25567
rect 4151 25511 4219 25567
rect 4275 25511 4343 25567
rect 4399 25511 4467 25567
rect 4523 25511 4591 25567
rect 4647 25511 4715 25567
rect 4771 25511 4839 25567
rect 4895 25511 4963 25567
rect 5019 25511 5045 25567
rect 4045 25443 5045 25511
rect 4045 25387 4095 25443
rect 4151 25387 4219 25443
rect 4275 25387 4343 25443
rect 4399 25387 4467 25443
rect 4523 25387 4591 25443
rect 4647 25387 4715 25443
rect 4771 25387 4839 25443
rect 4895 25387 4963 25443
rect 5019 25387 5045 25443
rect 4045 25319 5045 25387
rect 4045 25263 4095 25319
rect 4151 25263 4219 25319
rect 4275 25263 4343 25319
rect 4399 25263 4467 25319
rect 4523 25263 4591 25319
rect 4647 25263 4715 25319
rect 4771 25263 4839 25319
rect 4895 25263 4963 25319
rect 5019 25263 5045 25319
rect 4045 25195 5045 25263
rect 4045 25139 4095 25195
rect 4151 25139 4219 25195
rect 4275 25139 4343 25195
rect 4399 25139 4467 25195
rect 4523 25139 4591 25195
rect 4647 25139 4715 25195
rect 4771 25139 4839 25195
rect 4895 25139 4963 25195
rect 5019 25139 5045 25195
rect 4045 25071 5045 25139
rect 4045 25015 4095 25071
rect 4151 25015 4219 25071
rect 4275 25015 4343 25071
rect 4399 25015 4467 25071
rect 4523 25015 4591 25071
rect 4647 25015 4715 25071
rect 4771 25015 4839 25071
rect 4895 25015 4963 25071
rect 5019 25015 5045 25071
rect 4045 24947 5045 25015
rect 4045 24891 4095 24947
rect 4151 24891 4219 24947
rect 4275 24891 4343 24947
rect 4399 24891 4467 24947
rect 4523 24891 4591 24947
rect 4647 24891 4715 24947
rect 4771 24891 4839 24947
rect 4895 24891 4963 24947
rect 5019 24891 5045 24947
rect 4045 24823 5045 24891
rect 4045 24767 4095 24823
rect 4151 24767 4219 24823
rect 4275 24767 4343 24823
rect 4399 24767 4467 24823
rect 4523 24767 4591 24823
rect 4647 24767 4715 24823
rect 4771 24767 4839 24823
rect 4895 24767 4963 24823
rect 5019 24767 5045 24823
rect 3621 24064 3945 24074
rect 3621 24008 3631 24064
rect 3687 24008 3755 24064
rect 3811 24008 3879 24064
rect 3935 24008 3945 24064
rect 3621 23940 3945 24008
rect 3621 23884 3631 23940
rect 3687 23884 3755 23940
rect 3811 23884 3879 23940
rect 3935 23884 3945 23940
rect 3621 23816 3945 23884
rect 3621 23760 3631 23816
rect 3687 23760 3755 23816
rect 3811 23760 3879 23816
rect 3935 23760 3945 23816
rect 3621 23692 3945 23760
rect 3621 23636 3631 23692
rect 3687 23636 3755 23692
rect 3811 23636 3879 23692
rect 3935 23636 3945 23692
rect 3621 23568 3945 23636
rect 3621 23512 3631 23568
rect 3687 23512 3755 23568
rect 3811 23512 3879 23568
rect 3935 23512 3945 23568
rect 3621 23444 3945 23512
rect 3621 23388 3631 23444
rect 3687 23388 3755 23444
rect 3811 23388 3879 23444
rect 3935 23388 3945 23444
rect 3621 23320 3945 23388
rect 3621 23264 3631 23320
rect 3687 23264 3755 23320
rect 3811 23264 3879 23320
rect 3935 23264 3945 23320
rect 3621 23196 3945 23264
rect 3621 23140 3631 23196
rect 3687 23140 3755 23196
rect 3811 23140 3879 23196
rect 3935 23140 3945 23196
rect 3621 23130 3945 23140
rect 4045 22512 5045 24767
rect 4045 22456 4095 22512
rect 4151 22456 4219 22512
rect 4275 22456 4343 22512
rect 4399 22456 4467 22512
rect 4523 22456 4591 22512
rect 4647 22456 4715 22512
rect 4771 22456 4839 22512
rect 4895 22456 4963 22512
rect 5019 22456 5045 22512
rect 4045 22388 5045 22456
rect 4045 22332 4095 22388
rect 4151 22332 4219 22388
rect 4275 22332 4343 22388
rect 4399 22332 4467 22388
rect 4523 22332 4591 22388
rect 4647 22332 4715 22388
rect 4771 22332 4839 22388
rect 4895 22332 4963 22388
rect 5019 22332 5045 22388
rect 4045 22264 5045 22332
rect 4045 22208 4095 22264
rect 4151 22208 4219 22264
rect 4275 22208 4343 22264
rect 4399 22208 4467 22264
rect 4523 22208 4591 22264
rect 4647 22208 4715 22264
rect 4771 22208 4839 22264
rect 4895 22208 4963 22264
rect 5019 22208 5045 22264
rect 4045 22140 5045 22208
rect 4045 22084 4095 22140
rect 4151 22084 4219 22140
rect 4275 22084 4343 22140
rect 4399 22084 4467 22140
rect 4523 22084 4591 22140
rect 4647 22084 4715 22140
rect 4771 22084 4839 22140
rect 4895 22084 4963 22140
rect 5019 22084 5045 22140
rect 4045 22016 5045 22084
rect 4045 21960 4095 22016
rect 4151 21960 4219 22016
rect 4275 21960 4343 22016
rect 4399 21960 4467 22016
rect 4523 21960 4591 22016
rect 4647 21960 4715 22016
rect 4771 21960 4839 22016
rect 4895 21960 4963 22016
rect 5019 21960 5045 22016
rect 4045 21892 5045 21960
rect 4045 21836 4095 21892
rect 4151 21836 4219 21892
rect 4275 21836 4343 21892
rect 4399 21836 4467 21892
rect 4523 21836 4591 21892
rect 4647 21836 4715 21892
rect 4771 21836 4839 21892
rect 4895 21836 4963 21892
rect 5019 21836 5045 21892
rect 4045 21768 5045 21836
rect 4045 21712 4095 21768
rect 4151 21712 4219 21768
rect 4275 21712 4343 21768
rect 4399 21712 4467 21768
rect 4523 21712 4591 21768
rect 4647 21712 4715 21768
rect 4771 21712 4839 21768
rect 4895 21712 4963 21768
rect 5019 21712 5045 21768
rect 4045 21644 5045 21712
rect 4045 21588 4095 21644
rect 4151 21588 4219 21644
rect 4275 21588 4343 21644
rect 4399 21588 4467 21644
rect 4523 21588 4591 21644
rect 4647 21588 4715 21644
rect 4771 21588 4839 21644
rect 4895 21588 4963 21644
rect 5019 21588 5045 21644
rect 4045 21520 5045 21588
rect 4045 21464 4095 21520
rect 4151 21464 4219 21520
rect 4275 21464 4343 21520
rect 4399 21464 4467 21520
rect 4523 21464 4591 21520
rect 4647 21464 4715 21520
rect 4771 21464 4839 21520
rect 4895 21464 4963 21520
rect 5019 21464 5045 21520
rect 4045 21396 5045 21464
rect 4045 21340 4095 21396
rect 4151 21340 4219 21396
rect 4275 21340 4343 21396
rect 4399 21340 4467 21396
rect 4523 21340 4591 21396
rect 4647 21340 4715 21396
rect 4771 21340 4839 21396
rect 4895 21340 4963 21396
rect 5019 21340 5045 21396
rect 4045 21272 5045 21340
rect 4045 21216 4095 21272
rect 4151 21216 4219 21272
rect 4275 21216 4343 21272
rect 4399 21216 4467 21272
rect 4523 21216 4591 21272
rect 4647 21216 4715 21272
rect 4771 21216 4839 21272
rect 4895 21216 4963 21272
rect 5019 21216 5045 21272
rect 4045 21148 5045 21216
rect 4045 21092 4095 21148
rect 4151 21092 4219 21148
rect 4275 21092 4343 21148
rect 4399 21092 4467 21148
rect 4523 21092 4591 21148
rect 4647 21092 4715 21148
rect 4771 21092 4839 21148
rect 4895 21092 4963 21148
rect 5019 21092 5045 21148
rect 4045 21024 5045 21092
rect 4045 20968 4095 21024
rect 4151 20968 4219 21024
rect 4275 20968 4343 21024
rect 4399 20968 4467 21024
rect 4523 20968 4591 21024
rect 4647 20968 4715 21024
rect 4771 20968 4839 21024
rect 4895 20968 4963 21024
rect 5019 20968 5045 21024
rect 4045 20900 5045 20968
rect 4045 20844 4095 20900
rect 4151 20844 4219 20900
rect 4275 20844 4343 20900
rect 4399 20844 4467 20900
rect 4523 20844 4591 20900
rect 4647 20844 4715 20900
rect 4771 20844 4839 20900
rect 4895 20844 4963 20900
rect 5019 20844 5045 20900
rect 4045 20776 5045 20844
rect 4045 20720 4095 20776
rect 4151 20720 4219 20776
rect 4275 20720 4343 20776
rect 4399 20720 4467 20776
rect 4523 20720 4591 20776
rect 4647 20720 4715 20776
rect 4771 20720 4839 20776
rect 4895 20720 4963 20776
rect 5019 20720 5045 20776
rect 4045 20652 5045 20720
rect 4045 20596 4095 20652
rect 4151 20596 4219 20652
rect 4275 20596 4343 20652
rect 4399 20596 4467 20652
rect 4523 20596 4591 20652
rect 4647 20596 4715 20652
rect 4771 20596 4839 20652
rect 4895 20596 4963 20652
rect 5019 20596 5045 20652
rect 4045 20528 5045 20596
rect 4045 20472 4095 20528
rect 4151 20472 4219 20528
rect 4275 20472 4343 20528
rect 4399 20472 4467 20528
rect 4523 20472 4591 20528
rect 4647 20472 4715 20528
rect 4771 20472 4839 20528
rect 4895 20472 4963 20528
rect 5019 20472 5045 20528
rect 4045 20404 5045 20472
rect 4045 20348 4095 20404
rect 4151 20348 4219 20404
rect 4275 20348 4343 20404
rect 4399 20348 4467 20404
rect 4523 20348 4591 20404
rect 4647 20348 4715 20404
rect 4771 20348 4839 20404
rect 4895 20348 4963 20404
rect 5019 20348 5045 20404
rect 4045 20280 5045 20348
rect 4045 20224 4095 20280
rect 4151 20224 4219 20280
rect 4275 20224 4343 20280
rect 4399 20224 4467 20280
rect 4523 20224 4591 20280
rect 4647 20224 4715 20280
rect 4771 20224 4839 20280
rect 4895 20224 4963 20280
rect 5019 20224 5045 20280
rect 4045 20156 5045 20224
rect 4045 20100 4095 20156
rect 4151 20100 4219 20156
rect 4275 20100 4343 20156
rect 4399 20100 4467 20156
rect 4523 20100 4591 20156
rect 4647 20100 4715 20156
rect 4771 20100 4839 20156
rect 4895 20100 4963 20156
rect 5019 20100 5045 20156
rect 4045 20032 5045 20100
rect 4045 19976 4095 20032
rect 4151 19976 4219 20032
rect 4275 19976 4343 20032
rect 4399 19976 4467 20032
rect 4523 19976 4591 20032
rect 4647 19976 4715 20032
rect 4771 19976 4839 20032
rect 4895 19976 4963 20032
rect 5019 19976 5045 20032
rect 4045 19908 5045 19976
rect 4045 19852 4095 19908
rect 4151 19852 4219 19908
rect 4275 19852 4343 19908
rect 4399 19852 4467 19908
rect 4523 19852 4591 19908
rect 4647 19852 4715 19908
rect 4771 19852 4839 19908
rect 4895 19852 4963 19908
rect 5019 19852 5045 19908
rect 3621 19507 3945 19517
rect 3621 19451 3631 19507
rect 3687 19451 3755 19507
rect 3811 19451 3879 19507
rect 3935 19451 3945 19507
rect 3621 19383 3945 19451
rect 3621 19327 3631 19383
rect 3687 19327 3755 19383
rect 3811 19327 3879 19383
rect 3935 19327 3945 19383
rect 3621 19259 3945 19327
rect 3621 19203 3631 19259
rect 3687 19203 3755 19259
rect 3811 19203 3879 19259
rect 3935 19203 3945 19259
rect 3621 19135 3945 19203
rect 3621 19079 3631 19135
rect 3687 19079 3755 19135
rect 3811 19079 3879 19135
rect 3935 19079 3945 19135
rect 3621 19011 3945 19079
rect 3621 18955 3631 19011
rect 3687 18955 3755 19011
rect 3811 18955 3879 19011
rect 3935 18955 3945 19011
rect 3621 18887 3945 18955
rect 3621 18831 3631 18887
rect 3687 18831 3755 18887
rect 3811 18831 3879 18887
rect 3935 18831 3945 18887
rect 3621 18763 3945 18831
rect 3621 18707 3631 18763
rect 3687 18707 3755 18763
rect 3811 18707 3879 18763
rect 3935 18707 3945 18763
rect 3621 18639 3945 18707
rect 3621 18583 3631 18639
rect 3687 18583 3755 18639
rect 3811 18583 3879 18639
rect 3935 18583 3945 18639
rect 3621 18515 3945 18583
rect 3621 18459 3631 18515
rect 3687 18459 3755 18515
rect 3811 18459 3879 18515
rect 3935 18459 3945 18515
rect 3621 18391 3945 18459
rect 3621 18335 3631 18391
rect 3687 18335 3755 18391
rect 3811 18335 3879 18391
rect 3935 18335 3945 18391
rect 3621 18267 3945 18335
rect 3621 18211 3631 18267
rect 3687 18211 3755 18267
rect 3811 18211 3879 18267
rect 3935 18211 3945 18267
rect 3621 18143 3945 18211
rect 3621 18087 3631 18143
rect 3687 18087 3755 18143
rect 3811 18087 3879 18143
rect 3935 18087 3945 18143
rect 3621 18019 3945 18087
rect 3621 17963 3631 18019
rect 3687 17963 3755 18019
rect 3811 17963 3879 18019
rect 3935 17963 3945 18019
rect 3621 17895 3945 17963
rect 3621 17839 3631 17895
rect 3687 17839 3755 17895
rect 3811 17839 3879 17895
rect 3935 17839 3945 17895
rect 3621 17771 3945 17839
rect 3621 17715 3631 17771
rect 3687 17715 3755 17771
rect 3811 17715 3879 17771
rect 3935 17715 3945 17771
rect 3621 17647 3945 17715
rect 3621 17591 3631 17647
rect 3687 17591 3755 17647
rect 3811 17591 3879 17647
rect 3935 17591 3945 17647
rect 3621 17523 3945 17591
rect 3621 17467 3631 17523
rect 3687 17467 3755 17523
rect 3811 17467 3879 17523
rect 3935 17467 3945 17523
rect 3621 17399 3945 17467
rect 3621 17343 3631 17399
rect 3687 17343 3755 17399
rect 3811 17343 3879 17399
rect 3935 17343 3945 17399
rect 3621 17275 3945 17343
rect 3621 17219 3631 17275
rect 3687 17219 3755 17275
rect 3811 17219 3879 17275
rect 3935 17219 3945 17275
rect 3621 17151 3945 17219
rect 3621 17095 3631 17151
rect 3687 17095 3755 17151
rect 3811 17095 3879 17151
rect 3935 17095 3945 17151
rect 3621 17027 3945 17095
rect 3621 16971 3631 17027
rect 3687 16971 3755 17027
rect 3811 16971 3879 17027
rect 3935 16971 3945 17027
rect 3621 16903 3945 16971
rect 3621 16847 3631 16903
rect 3687 16847 3755 16903
rect 3811 16847 3879 16903
rect 3935 16847 3945 16903
rect 3621 16779 3945 16847
rect 3621 16723 3631 16779
rect 3687 16723 3755 16779
rect 3811 16723 3879 16779
rect 3935 16723 3945 16779
rect 3621 16655 3945 16723
rect 3621 16599 3631 16655
rect 3687 16599 3755 16655
rect 3811 16599 3879 16655
rect 3935 16599 3945 16655
rect 3621 16531 3945 16599
rect 3621 16475 3631 16531
rect 3687 16475 3755 16531
rect 3811 16475 3879 16531
rect 3935 16475 3945 16531
rect 3621 16407 3945 16475
rect 3621 16351 3631 16407
rect 3687 16351 3755 16407
rect 3811 16351 3879 16407
rect 3935 16351 3945 16407
rect 3621 16283 3945 16351
rect 3621 16227 3631 16283
rect 3687 16227 3755 16283
rect 3811 16227 3879 16283
rect 3935 16227 3945 16283
rect 3621 16217 3945 16227
rect 4045 15942 5045 19852
rect 4045 15886 4095 15942
rect 4151 15886 4219 15942
rect 4275 15886 4343 15942
rect 4399 15886 4467 15942
rect 4523 15886 4591 15942
rect 4647 15886 4715 15942
rect 4771 15886 4839 15942
rect 4895 15886 4963 15942
rect 5019 15886 5045 15942
rect 4045 15818 5045 15886
rect 4045 15762 4095 15818
rect 4151 15762 4219 15818
rect 4275 15762 4343 15818
rect 4399 15762 4467 15818
rect 4523 15762 4591 15818
rect 4647 15762 4715 15818
rect 4771 15762 4839 15818
rect 4895 15762 4963 15818
rect 5019 15762 5045 15818
rect 4045 15694 5045 15762
rect 4045 15638 4095 15694
rect 4151 15638 4219 15694
rect 4275 15638 4343 15694
rect 4399 15638 4467 15694
rect 4523 15638 4591 15694
rect 4647 15638 4715 15694
rect 4771 15638 4839 15694
rect 4895 15638 4963 15694
rect 5019 15638 5045 15694
rect 4045 15570 5045 15638
rect 4045 15514 4095 15570
rect 4151 15514 4219 15570
rect 4275 15514 4343 15570
rect 4399 15514 4467 15570
rect 4523 15514 4591 15570
rect 4647 15514 4715 15570
rect 4771 15514 4839 15570
rect 4895 15514 4963 15570
rect 5019 15514 5045 15570
rect 4045 15446 5045 15514
rect 4045 15390 4095 15446
rect 4151 15390 4219 15446
rect 4275 15390 4343 15446
rect 4399 15390 4467 15446
rect 4523 15390 4591 15446
rect 4647 15390 4715 15446
rect 4771 15390 4839 15446
rect 4895 15390 4963 15446
rect 5019 15390 5045 15446
rect 4045 15322 5045 15390
rect 4045 15266 4095 15322
rect 4151 15266 4219 15322
rect 4275 15266 4343 15322
rect 4399 15266 4467 15322
rect 4523 15266 4591 15322
rect 4647 15266 4715 15322
rect 4771 15266 4839 15322
rect 4895 15266 4963 15322
rect 5019 15266 5045 15322
rect 4045 15198 5045 15266
rect 4045 15142 4095 15198
rect 4151 15142 4219 15198
rect 4275 15142 4343 15198
rect 4399 15142 4467 15198
rect 4523 15142 4591 15198
rect 4647 15142 4715 15198
rect 4771 15142 4839 15198
rect 4895 15142 4963 15198
rect 5019 15142 5045 15198
rect 4045 15074 5045 15142
rect 4045 15018 4095 15074
rect 4151 15018 4219 15074
rect 4275 15018 4343 15074
rect 4399 15018 4467 15074
rect 4523 15018 4591 15074
rect 4647 15018 4715 15074
rect 4771 15018 4839 15074
rect 4895 15018 4963 15074
rect 5019 15018 5045 15074
rect 4045 14950 5045 15018
rect 4045 14894 4095 14950
rect 4151 14894 4219 14950
rect 4275 14894 4343 14950
rect 4399 14894 4467 14950
rect 4523 14894 4591 14950
rect 4647 14894 4715 14950
rect 4771 14894 4839 14950
rect 4895 14894 4963 14950
rect 5019 14894 5045 14950
rect 4045 14826 5045 14894
rect 4045 14770 4095 14826
rect 4151 14770 4219 14826
rect 4275 14770 4343 14826
rect 4399 14770 4467 14826
rect 4523 14770 4591 14826
rect 4647 14770 4715 14826
rect 4771 14770 4839 14826
rect 4895 14770 4963 14826
rect 5019 14770 5045 14826
rect 4045 14702 5045 14770
rect 4045 14646 4095 14702
rect 4151 14646 4219 14702
rect 4275 14646 4343 14702
rect 4399 14646 4467 14702
rect 4523 14646 4591 14702
rect 4647 14646 4715 14702
rect 4771 14646 4839 14702
rect 4895 14646 4963 14702
rect 5019 14646 5045 14702
rect 4045 14578 5045 14646
rect 4045 14522 4095 14578
rect 4151 14522 4219 14578
rect 4275 14522 4343 14578
rect 4399 14522 4467 14578
rect 4523 14522 4591 14578
rect 4647 14522 4715 14578
rect 4771 14522 4839 14578
rect 4895 14522 4963 14578
rect 5019 14522 5045 14578
rect 4045 14454 5045 14522
rect 4045 14398 4095 14454
rect 4151 14398 4219 14454
rect 4275 14398 4343 14454
rect 4399 14398 4467 14454
rect 4523 14398 4591 14454
rect 4647 14398 4715 14454
rect 4771 14398 4839 14454
rect 4895 14398 4963 14454
rect 5019 14398 5045 14454
rect 4045 14330 5045 14398
rect 4045 14274 4095 14330
rect 4151 14274 4219 14330
rect 4275 14274 4343 14330
rect 4399 14274 4467 14330
rect 4523 14274 4591 14330
rect 4647 14274 4715 14330
rect 4771 14274 4839 14330
rect 4895 14274 4963 14330
rect 5019 14274 5045 14330
rect 4045 14206 5045 14274
rect 4045 14150 4095 14206
rect 4151 14150 4219 14206
rect 4275 14150 4343 14206
rect 4399 14150 4467 14206
rect 4523 14150 4591 14206
rect 4647 14150 4715 14206
rect 4771 14150 4839 14206
rect 4895 14150 4963 14206
rect 5019 14150 5045 14206
rect 4045 14082 5045 14150
rect 4045 14026 4095 14082
rect 4151 14026 4219 14082
rect 4275 14026 4343 14082
rect 4399 14026 4467 14082
rect 4523 14026 4591 14082
rect 4647 14026 4715 14082
rect 4771 14026 4839 14082
rect 4895 14026 4963 14082
rect 5019 14026 5045 14082
rect 4045 13958 5045 14026
rect 4045 13902 4095 13958
rect 4151 13902 4219 13958
rect 4275 13902 4343 13958
rect 4399 13902 4467 13958
rect 4523 13902 4591 13958
rect 4647 13902 4715 13958
rect 4771 13902 4839 13958
rect 4895 13902 4963 13958
rect 5019 13902 5045 13958
rect 3621 13228 3945 13238
rect 3621 13172 3631 13228
rect 3687 13172 3755 13228
rect 3811 13172 3879 13228
rect 3935 13172 3945 13228
rect 3621 13104 3945 13172
rect 3621 13048 3631 13104
rect 3687 13048 3755 13104
rect 3811 13048 3879 13104
rect 3935 13048 3945 13104
rect 3621 12980 3945 13048
rect 3621 12924 3631 12980
rect 3687 12924 3755 12980
rect 3811 12924 3879 12980
rect 3935 12924 3945 12980
rect 3621 12856 3945 12924
rect 3621 12800 3631 12856
rect 3687 12800 3755 12856
rect 3811 12800 3879 12856
rect 3935 12800 3945 12856
rect 3621 12732 3945 12800
rect 3621 12676 3631 12732
rect 3687 12676 3755 12732
rect 3811 12676 3879 12732
rect 3935 12676 3945 12732
rect 3621 12608 3945 12676
rect 3621 12552 3631 12608
rect 3687 12552 3755 12608
rect 3811 12552 3879 12608
rect 3935 12552 3945 12608
rect 3621 12484 3945 12552
rect 3621 12428 3631 12484
rect 3687 12428 3755 12484
rect 3811 12428 3879 12484
rect 3935 12428 3945 12484
rect 3621 12360 3945 12428
rect 3621 12304 3631 12360
rect 3687 12304 3755 12360
rect 3811 12304 3879 12360
rect 3935 12304 3945 12360
rect 3621 12236 3945 12304
rect 3621 12180 3631 12236
rect 3687 12180 3755 12236
rect 3811 12180 3879 12236
rect 3935 12180 3945 12236
rect 3621 12112 3945 12180
rect 3621 12056 3631 12112
rect 3687 12056 3755 12112
rect 3811 12056 3879 12112
rect 3935 12056 3945 12112
rect 3621 12046 3945 12056
rect 4045 11292 5045 13902
rect 4045 11236 4095 11292
rect 4151 11236 4219 11292
rect 4275 11236 4343 11292
rect 4399 11236 4467 11292
rect 4523 11236 4591 11292
rect 4647 11236 4715 11292
rect 4771 11236 4839 11292
rect 4895 11236 4963 11292
rect 5019 11236 5045 11292
rect 4045 11168 5045 11236
rect 4045 11112 4095 11168
rect 4151 11112 4219 11168
rect 4275 11112 4343 11168
rect 4399 11112 4467 11168
rect 4523 11112 4591 11168
rect 4647 11112 4715 11168
rect 4771 11112 4839 11168
rect 4895 11112 4963 11168
rect 5019 11112 5045 11168
rect 4045 11044 5045 11112
rect 4045 10988 4095 11044
rect 4151 10988 4219 11044
rect 4275 10988 4343 11044
rect 4399 10988 4467 11044
rect 4523 10988 4591 11044
rect 4647 10988 4715 11044
rect 4771 10988 4839 11044
rect 4895 10988 4963 11044
rect 5019 10988 5045 11044
rect 4045 10920 5045 10988
rect 4045 10864 4095 10920
rect 4151 10864 4219 10920
rect 4275 10864 4343 10920
rect 4399 10864 4467 10920
rect 4523 10864 4591 10920
rect 4647 10864 4715 10920
rect 4771 10864 4839 10920
rect 4895 10864 4963 10920
rect 5019 10864 5045 10920
rect 4045 10796 5045 10864
rect 4045 10740 4095 10796
rect 4151 10740 4219 10796
rect 4275 10740 4343 10796
rect 4399 10740 4467 10796
rect 4523 10740 4591 10796
rect 4647 10740 4715 10796
rect 4771 10740 4839 10796
rect 4895 10740 4963 10796
rect 5019 10740 5045 10796
rect 4045 10672 5045 10740
rect 4045 10616 4095 10672
rect 4151 10616 4219 10672
rect 4275 10616 4343 10672
rect 4399 10616 4467 10672
rect 4523 10616 4591 10672
rect 4647 10616 4715 10672
rect 4771 10616 4839 10672
rect 4895 10616 4963 10672
rect 5019 10616 5045 10672
rect 4045 10548 5045 10616
rect 4045 10492 4095 10548
rect 4151 10492 4219 10548
rect 4275 10492 4343 10548
rect 4399 10492 4467 10548
rect 4523 10492 4591 10548
rect 4647 10492 4715 10548
rect 4771 10492 4839 10548
rect 4895 10492 4963 10548
rect 5019 10492 5045 10548
rect 4045 10424 5045 10492
rect 4045 10368 4095 10424
rect 4151 10368 4219 10424
rect 4275 10368 4343 10424
rect 4399 10368 4467 10424
rect 4523 10368 4591 10424
rect 4647 10368 4715 10424
rect 4771 10368 4839 10424
rect 4895 10368 4963 10424
rect 5019 10368 5045 10424
rect 4045 10300 5045 10368
rect 4045 10244 4095 10300
rect 4151 10244 4219 10300
rect 4275 10244 4343 10300
rect 4399 10244 4467 10300
rect 4523 10244 4591 10300
rect 4647 10244 4715 10300
rect 4771 10244 4839 10300
rect 4895 10244 4963 10300
rect 5019 10244 5045 10300
rect 4045 10176 5045 10244
rect 4045 10120 4095 10176
rect 4151 10120 4219 10176
rect 4275 10120 4343 10176
rect 4399 10120 4467 10176
rect 4523 10120 4591 10176
rect 4647 10120 4715 10176
rect 4771 10120 4839 10176
rect 4895 10120 4963 10176
rect 5019 10120 5045 10176
rect 4045 10052 5045 10120
rect 4045 9996 4095 10052
rect 4151 9996 4219 10052
rect 4275 9996 4343 10052
rect 4399 9996 4467 10052
rect 4523 9996 4591 10052
rect 4647 9996 4715 10052
rect 4771 9996 4839 10052
rect 4895 9996 4963 10052
rect 5019 9996 5045 10052
rect 3621 9392 3945 9402
rect 3621 9336 3631 9392
rect 3687 9336 3755 9392
rect 3811 9336 3879 9392
rect 3935 9336 3945 9392
rect 3621 9268 3945 9336
rect 3621 9212 3631 9268
rect 3687 9212 3755 9268
rect 3811 9212 3879 9268
rect 3935 9212 3945 9268
rect 3621 9144 3945 9212
rect 3621 9088 3631 9144
rect 3687 9088 3755 9144
rect 3811 9088 3879 9144
rect 3935 9088 3945 9144
rect 3621 9020 3945 9088
rect 3621 8964 3631 9020
rect 3687 8964 3755 9020
rect 3811 8964 3879 9020
rect 3935 8964 3945 9020
rect 3621 8896 3945 8964
rect 3621 8840 3631 8896
rect 3687 8840 3755 8896
rect 3811 8840 3879 8896
rect 3935 8840 3945 8896
rect 3621 8772 3945 8840
rect 3621 8716 3631 8772
rect 3687 8716 3755 8772
rect 3811 8716 3879 8772
rect 3935 8716 3945 8772
rect 3621 8648 3945 8716
rect 3621 8592 3631 8648
rect 3687 8592 3755 8648
rect 3811 8592 3879 8648
rect 3935 8592 3945 8648
rect 3621 8524 3945 8592
rect 3621 8468 3631 8524
rect 3687 8468 3755 8524
rect 3811 8468 3879 8524
rect 3935 8468 3945 8524
rect 3621 8400 3945 8468
rect 3621 8344 3631 8400
rect 3687 8344 3755 8400
rect 3811 8344 3879 8400
rect 3935 8344 3945 8400
rect 3621 8276 3945 8344
rect 3621 8220 3631 8276
rect 3687 8220 3755 8276
rect 3811 8220 3879 8276
rect 3935 8220 3945 8276
rect 3621 8152 3945 8220
rect 3621 8096 3631 8152
rect 3687 8096 3755 8152
rect 3811 8096 3879 8152
rect 3935 8096 3945 8152
rect 3621 8028 3945 8096
rect 3621 7972 3631 8028
rect 3687 7972 3755 8028
rect 3811 7972 3879 8028
rect 3935 7972 3945 8028
rect 3621 7904 3945 7972
rect 3621 7848 3631 7904
rect 3687 7848 3755 7904
rect 3811 7848 3879 7904
rect 3935 7848 3945 7904
rect 3621 7780 3945 7848
rect 3621 7724 3631 7780
rect 3687 7724 3755 7780
rect 3811 7724 3879 7780
rect 3935 7724 3945 7780
rect 3621 7656 3945 7724
rect 3621 7600 3631 7656
rect 3687 7600 3755 7656
rect 3811 7600 3879 7656
rect 3935 7600 3945 7656
rect 3621 7590 3945 7600
rect 4045 7435 5045 9996
rect 4045 7379 4095 7435
rect 4151 7379 4219 7435
rect 4275 7379 4343 7435
rect 4399 7379 4467 7435
rect 4523 7379 4591 7435
rect 4647 7379 4715 7435
rect 4771 7379 4839 7435
rect 4895 7379 4963 7435
rect 5019 7379 5045 7435
rect 4045 7311 5045 7379
rect 4045 7255 4095 7311
rect 4151 7255 4219 7311
rect 4275 7255 4343 7311
rect 4399 7255 4467 7311
rect 4523 7255 4591 7311
rect 4647 7255 4715 7311
rect 4771 7255 4839 7311
rect 4895 7255 4963 7311
rect 5019 7255 5045 7311
rect 4045 7187 5045 7255
rect 4045 7131 4095 7187
rect 4151 7131 4219 7187
rect 4275 7131 4343 7187
rect 4399 7131 4467 7187
rect 4523 7131 4591 7187
rect 4647 7131 4715 7187
rect 4771 7131 4839 7187
rect 4895 7131 4963 7187
rect 5019 7131 5045 7187
rect 4045 7063 5045 7131
rect 4045 7007 4095 7063
rect 4151 7007 4219 7063
rect 4275 7007 4343 7063
rect 4399 7007 4467 7063
rect 4523 7007 4591 7063
rect 4647 7007 4715 7063
rect 4771 7007 4839 7063
rect 4895 7007 4963 7063
rect 5019 7007 5045 7063
rect 4045 6939 5045 7007
rect 4045 6883 4095 6939
rect 4151 6883 4219 6939
rect 4275 6883 4343 6939
rect 4399 6883 4467 6939
rect 4523 6883 4591 6939
rect 4647 6883 4715 6939
rect 4771 6883 4839 6939
rect 4895 6883 4963 6939
rect 5019 6883 5045 6939
rect 4045 6815 5045 6883
rect 4045 6759 4095 6815
rect 4151 6759 4219 6815
rect 4275 6759 4343 6815
rect 4399 6759 4467 6815
rect 4523 6759 4591 6815
rect 4647 6759 4715 6815
rect 4771 6759 4839 6815
rect 4895 6759 4963 6815
rect 5019 6759 5045 6815
rect 4045 6691 5045 6759
rect 4045 6635 4095 6691
rect 4151 6635 4219 6691
rect 4275 6635 4343 6691
rect 4399 6635 4467 6691
rect 4523 6635 4591 6691
rect 4647 6635 4715 6691
rect 4771 6635 4839 6691
rect 4895 6635 4963 6691
rect 5019 6635 5045 6691
rect 4045 6567 5045 6635
rect 4045 6511 4095 6567
rect 4151 6511 4219 6567
rect 4275 6511 4343 6567
rect 4399 6511 4467 6567
rect 4523 6511 4591 6567
rect 4647 6511 4715 6567
rect 4771 6511 4839 6567
rect 4895 6511 4963 6567
rect 5019 6511 5045 6567
rect 4045 6443 5045 6511
rect 4045 6387 4095 6443
rect 4151 6387 4219 6443
rect 4275 6387 4343 6443
rect 4399 6387 4467 6443
rect 4523 6387 4591 6443
rect 4647 6387 4715 6443
rect 4771 6387 4839 6443
rect 4895 6387 4963 6443
rect 5019 6387 5045 6443
rect 4045 6319 5045 6387
rect 4045 6263 4095 6319
rect 4151 6263 4219 6319
rect 4275 6263 4343 6319
rect 4399 6263 4467 6319
rect 4523 6263 4591 6319
rect 4647 6263 4715 6319
rect 4771 6263 4839 6319
rect 4895 6263 4963 6319
rect 5019 6263 5045 6319
rect 4045 6195 5045 6263
rect 4045 6139 4095 6195
rect 4151 6139 4219 6195
rect 4275 6139 4343 6195
rect 4399 6139 4467 6195
rect 4523 6139 4591 6195
rect 4647 6139 4715 6195
rect 4771 6139 4839 6195
rect 4895 6139 4963 6195
rect 5019 6139 5045 6195
rect 4045 6071 5045 6139
rect 4045 6015 4095 6071
rect 4151 6015 4219 6071
rect 4275 6015 4343 6071
rect 4399 6015 4467 6071
rect 4523 6015 4591 6071
rect 4647 6015 4715 6071
rect 4771 6015 4839 6071
rect 4895 6015 4963 6071
rect 5019 6015 5045 6071
rect 4045 5947 5045 6015
rect 4045 5891 4095 5947
rect 4151 5891 4219 5947
rect 4275 5891 4343 5947
rect 4399 5891 4467 5947
rect 4523 5891 4591 5947
rect 4647 5891 4715 5947
rect 4771 5891 4839 5947
rect 4895 5891 4963 5947
rect 5019 5891 5045 5947
rect 3621 5528 3945 5538
rect 3621 5472 3631 5528
rect 3687 5472 3755 5528
rect 3811 5472 3879 5528
rect 3935 5472 3945 5528
rect 3621 5404 3945 5472
rect 3621 5348 3631 5404
rect 3687 5348 3755 5404
rect 3811 5348 3879 5404
rect 3935 5348 3945 5404
rect 3621 5280 3945 5348
rect 3621 5224 3631 5280
rect 3687 5224 3755 5280
rect 3811 5224 3879 5280
rect 3935 5224 3945 5280
rect 3621 5156 3945 5224
rect 3621 5100 3631 5156
rect 3687 5100 3755 5156
rect 3811 5100 3879 5156
rect 3935 5100 3945 5156
rect 3621 5032 3945 5100
rect 3621 4976 3631 5032
rect 3687 4976 3755 5032
rect 3811 4976 3879 5032
rect 3935 4976 3945 5032
rect 3621 4908 3945 4976
rect 3621 4852 3631 4908
rect 3687 4852 3755 4908
rect 3811 4852 3879 4908
rect 3935 4852 3945 4908
rect 3621 4784 3945 4852
rect 3621 4728 3631 4784
rect 3687 4728 3755 4784
rect 3811 4728 3879 4784
rect 3935 4728 3945 4784
rect 3621 4660 3945 4728
rect 3621 4604 3631 4660
rect 3687 4604 3755 4660
rect 3811 4604 3879 4660
rect 3935 4604 3945 4660
rect 3621 4536 3945 4604
rect 3621 4480 3631 4536
rect 3687 4480 3755 4536
rect 3811 4480 3879 4536
rect 3935 4480 3945 4536
rect 3621 4412 3945 4480
rect 3621 4356 3631 4412
rect 3687 4356 3755 4412
rect 3811 4356 3879 4412
rect 3935 4356 3945 4412
rect 3621 4346 3945 4356
rect 4045 4010 5045 5891
rect 4045 3954 4095 4010
rect 4151 3954 4219 4010
rect 4275 3954 4343 4010
rect 4399 3954 4467 4010
rect 4523 3954 4591 4010
rect 4647 3954 4715 4010
rect 4771 3954 4839 4010
rect 4895 3954 4963 4010
rect 5019 3954 5045 4010
rect 4045 3886 5045 3954
rect 4045 3830 4095 3886
rect 4151 3830 4219 3886
rect 4275 3830 4343 3886
rect 4399 3830 4467 3886
rect 4523 3830 4591 3886
rect 4647 3830 4715 3886
rect 4771 3830 4839 3886
rect 4895 3830 4963 3886
rect 5019 3830 5045 3886
rect 4045 3762 5045 3830
rect 4045 3706 4095 3762
rect 4151 3706 4219 3762
rect 4275 3706 4343 3762
rect 4399 3706 4467 3762
rect 4523 3706 4591 3762
rect 4647 3706 4715 3762
rect 4771 3706 4839 3762
rect 4895 3706 4963 3762
rect 5019 3706 5045 3762
rect 4045 3638 5045 3706
rect 4045 3582 4095 3638
rect 4151 3582 4219 3638
rect 4275 3582 4343 3638
rect 4399 3582 4467 3638
rect 4523 3582 4591 3638
rect 4647 3582 4715 3638
rect 4771 3582 4839 3638
rect 4895 3582 4963 3638
rect 5019 3582 5045 3638
rect 4045 3514 5045 3582
rect 4045 3458 4095 3514
rect 4151 3458 4219 3514
rect 4275 3458 4343 3514
rect 4399 3458 4467 3514
rect 4523 3458 4591 3514
rect 4647 3458 4715 3514
rect 4771 3458 4839 3514
rect 4895 3458 4963 3514
rect 5019 3458 5045 3514
rect 4045 3390 5045 3458
rect 4045 3334 4095 3390
rect 4151 3334 4219 3390
rect 4275 3334 4343 3390
rect 4399 3334 4467 3390
rect 4523 3334 4591 3390
rect 4647 3334 4715 3390
rect 4771 3334 4839 3390
rect 4895 3334 4963 3390
rect 5019 3334 5045 3390
rect 4045 3266 5045 3334
rect 4045 3210 4095 3266
rect 4151 3210 4219 3266
rect 4275 3210 4343 3266
rect 4399 3210 4467 3266
rect 4523 3210 4591 3266
rect 4647 3210 4715 3266
rect 4771 3210 4839 3266
rect 4895 3210 4963 3266
rect 5019 3210 5045 3266
rect 4045 3142 5045 3210
rect 4045 3086 4095 3142
rect 4151 3086 4219 3142
rect 4275 3086 4343 3142
rect 4399 3086 4467 3142
rect 4523 3086 4591 3142
rect 4647 3086 4715 3142
rect 4771 3086 4839 3142
rect 4895 3086 4963 3142
rect 5019 3086 5045 3142
rect 4045 2101 5045 3086
<< via2 >>
rect 3631 37081 3687 37083
rect 3631 37029 3633 37081
rect 3633 37029 3685 37081
rect 3685 37029 3687 37081
rect 3631 37027 3687 37029
rect 3755 37081 3811 37083
rect 3755 37029 3757 37081
rect 3757 37029 3809 37081
rect 3809 37029 3811 37081
rect 3755 37027 3811 37029
rect 3879 37081 3935 37083
rect 3879 37029 3881 37081
rect 3881 37029 3933 37081
rect 3933 37029 3935 37081
rect 3879 37027 3935 37029
rect 3631 36957 3687 36959
rect 3631 36905 3633 36957
rect 3633 36905 3685 36957
rect 3685 36905 3687 36957
rect 3631 36903 3687 36905
rect 3755 36957 3811 36959
rect 3755 36905 3757 36957
rect 3757 36905 3809 36957
rect 3809 36905 3811 36957
rect 3755 36903 3811 36905
rect 3879 36957 3935 36959
rect 3879 36905 3881 36957
rect 3881 36905 3933 36957
rect 3933 36905 3935 36957
rect 3879 36903 3935 36905
rect 3631 36833 3687 36835
rect 3631 36781 3633 36833
rect 3633 36781 3685 36833
rect 3685 36781 3687 36833
rect 3631 36779 3687 36781
rect 3755 36833 3811 36835
rect 3755 36781 3757 36833
rect 3757 36781 3809 36833
rect 3809 36781 3811 36833
rect 3755 36779 3811 36781
rect 3879 36833 3935 36835
rect 3879 36781 3881 36833
rect 3881 36781 3933 36833
rect 3933 36781 3935 36833
rect 3879 36779 3935 36781
rect 3631 36709 3687 36711
rect 3631 36657 3633 36709
rect 3633 36657 3685 36709
rect 3685 36657 3687 36709
rect 3631 36655 3687 36657
rect 3755 36709 3811 36711
rect 3755 36657 3757 36709
rect 3757 36657 3809 36709
rect 3809 36657 3811 36709
rect 3755 36655 3811 36657
rect 3879 36709 3935 36711
rect 3879 36657 3881 36709
rect 3881 36657 3933 36709
rect 3933 36657 3935 36709
rect 3879 36655 3935 36657
rect 3631 36585 3687 36587
rect 3631 36533 3633 36585
rect 3633 36533 3685 36585
rect 3685 36533 3687 36585
rect 3631 36531 3687 36533
rect 3755 36585 3811 36587
rect 3755 36533 3757 36585
rect 3757 36533 3809 36585
rect 3809 36533 3811 36585
rect 3755 36531 3811 36533
rect 3879 36585 3935 36587
rect 3879 36533 3881 36585
rect 3881 36533 3933 36585
rect 3933 36533 3935 36585
rect 3879 36531 3935 36533
rect 3631 36461 3687 36463
rect 3631 36409 3633 36461
rect 3633 36409 3685 36461
rect 3685 36409 3687 36461
rect 3631 36407 3687 36409
rect 3755 36461 3811 36463
rect 3755 36409 3757 36461
rect 3757 36409 3809 36461
rect 3809 36409 3811 36461
rect 3755 36407 3811 36409
rect 3879 36461 3935 36463
rect 3879 36409 3881 36461
rect 3881 36409 3933 36461
rect 3933 36409 3935 36461
rect 3879 36407 3935 36409
rect 4095 35873 4151 35929
rect 4219 35873 4275 35929
rect 4343 35873 4399 35929
rect 4467 35873 4523 35929
rect 4591 35873 4647 35929
rect 4715 35873 4771 35929
rect 4839 35873 4895 35929
rect 4963 35873 5019 35929
rect 4095 35749 4151 35805
rect 4219 35749 4275 35805
rect 4343 35749 4399 35805
rect 4467 35749 4523 35805
rect 4591 35749 4647 35805
rect 4715 35749 4771 35805
rect 4839 35749 4895 35805
rect 4963 35749 5019 35805
rect 4095 35625 4151 35681
rect 4219 35625 4275 35681
rect 4343 35625 4399 35681
rect 4467 35625 4523 35681
rect 4591 35625 4647 35681
rect 4715 35625 4771 35681
rect 4839 35625 4895 35681
rect 4963 35625 5019 35681
rect 4095 35501 4151 35557
rect 4219 35501 4275 35557
rect 4343 35501 4399 35557
rect 4467 35501 4523 35557
rect 4591 35501 4647 35557
rect 4715 35501 4771 35557
rect 4839 35501 4895 35557
rect 4963 35501 5019 35557
rect 4095 35377 4151 35433
rect 4219 35377 4275 35433
rect 4343 35377 4399 35433
rect 4467 35377 4523 35433
rect 4591 35377 4647 35433
rect 4715 35377 4771 35433
rect 4839 35377 4895 35433
rect 4963 35377 5019 35433
rect 4095 35253 4151 35309
rect 4219 35253 4275 35309
rect 4343 35253 4399 35309
rect 4467 35253 4523 35309
rect 4591 35253 4647 35309
rect 4715 35253 4771 35309
rect 4839 35253 4895 35309
rect 4963 35253 5019 35309
rect 4095 35129 4151 35185
rect 4219 35129 4275 35185
rect 4343 35129 4399 35185
rect 4467 35129 4523 35185
rect 4591 35129 4647 35185
rect 4715 35129 4771 35185
rect 4839 35129 4895 35185
rect 4963 35129 5019 35185
rect 4095 35005 4151 35061
rect 4219 35005 4275 35061
rect 4343 35005 4399 35061
rect 4467 35005 4523 35061
rect 4591 35005 4647 35061
rect 4715 35005 4771 35061
rect 4839 35005 4895 35061
rect 4963 35005 5019 35061
rect 4095 34881 4151 34937
rect 4219 34881 4275 34937
rect 4343 34881 4399 34937
rect 4467 34881 4523 34937
rect 4591 34881 4647 34937
rect 4715 34881 4771 34937
rect 4839 34881 4895 34937
rect 4963 34881 5019 34937
rect 4095 34757 4151 34813
rect 4219 34757 4275 34813
rect 4343 34757 4399 34813
rect 4467 34757 4523 34813
rect 4591 34757 4647 34813
rect 4715 34757 4771 34813
rect 4839 34757 4895 34813
rect 4963 34757 5019 34813
rect 4095 34633 4151 34689
rect 4219 34633 4275 34689
rect 4343 34633 4399 34689
rect 4467 34633 4523 34689
rect 4591 34633 4647 34689
rect 4715 34633 4771 34689
rect 4839 34633 4895 34689
rect 4963 34633 5019 34689
rect 4095 34509 4151 34565
rect 4219 34509 4275 34565
rect 4343 34509 4399 34565
rect 4467 34509 4523 34565
rect 4591 34509 4647 34565
rect 4715 34509 4771 34565
rect 4839 34509 4895 34565
rect 4963 34509 5019 34565
rect 4095 34385 4151 34441
rect 4219 34385 4275 34441
rect 4343 34385 4399 34441
rect 4467 34385 4523 34441
rect 4591 34385 4647 34441
rect 4715 34385 4771 34441
rect 4839 34385 4895 34441
rect 4963 34385 5019 34441
rect 4095 34261 4151 34317
rect 4219 34261 4275 34317
rect 4343 34261 4399 34317
rect 4467 34261 4523 34317
rect 4591 34261 4647 34317
rect 4715 34261 4771 34317
rect 4839 34261 4895 34317
rect 4963 34261 5019 34317
rect 4095 34137 4151 34193
rect 4219 34137 4275 34193
rect 4343 34137 4399 34193
rect 4467 34137 4523 34193
rect 4591 34137 4647 34193
rect 4715 34137 4771 34193
rect 4839 34137 4895 34193
rect 4963 34137 5019 34193
rect 4095 34013 4151 34069
rect 4219 34013 4275 34069
rect 4343 34013 4399 34069
rect 4467 34013 4523 34069
rect 4591 34013 4647 34069
rect 4715 34013 4771 34069
rect 4839 34013 4895 34069
rect 4963 34013 5019 34069
rect 4095 33889 4151 33945
rect 4219 33889 4275 33945
rect 4343 33889 4399 33945
rect 4467 33889 4523 33945
rect 4591 33889 4647 33945
rect 4715 33889 4771 33945
rect 4839 33889 4895 33945
rect 4963 33889 5019 33945
rect 4095 33765 4151 33821
rect 4219 33765 4275 33821
rect 4343 33765 4399 33821
rect 4467 33765 4523 33821
rect 4591 33765 4647 33821
rect 4715 33765 4771 33821
rect 4839 33765 4895 33821
rect 4963 33765 5019 33821
rect 4095 33641 4151 33697
rect 4219 33641 4275 33697
rect 4343 33641 4399 33697
rect 4467 33641 4523 33697
rect 4591 33641 4647 33697
rect 4715 33641 4771 33697
rect 4839 33641 4895 33697
rect 4963 33641 5019 33697
rect 4095 33517 4151 33573
rect 4219 33517 4275 33573
rect 4343 33517 4399 33573
rect 4467 33517 4523 33573
rect 4591 33517 4647 33573
rect 4715 33517 4771 33573
rect 4839 33517 4895 33573
rect 4963 33517 5019 33573
rect 4095 33393 4151 33449
rect 4219 33393 4275 33449
rect 4343 33393 4399 33449
rect 4467 33393 4523 33449
rect 4591 33393 4647 33449
rect 4715 33393 4771 33449
rect 4839 33393 4895 33449
rect 4963 33393 5019 33449
rect 4095 33269 4151 33325
rect 4219 33269 4275 33325
rect 4343 33269 4399 33325
rect 4467 33269 4523 33325
rect 4591 33269 4647 33325
rect 4715 33269 4771 33325
rect 4839 33269 4895 33325
rect 4963 33269 5019 33325
rect 4095 33145 4151 33201
rect 4219 33145 4275 33201
rect 4343 33145 4399 33201
rect 4467 33145 4523 33201
rect 4591 33145 4647 33201
rect 4715 33145 4771 33201
rect 4839 33145 4895 33201
rect 4963 33145 5019 33201
rect 4095 33021 4151 33077
rect 4219 33021 4275 33077
rect 4343 33021 4399 33077
rect 4467 33021 4523 33077
rect 4591 33021 4647 33077
rect 4715 33021 4771 33077
rect 4839 33021 4895 33077
rect 4963 33021 5019 33077
rect 4095 32897 4151 32953
rect 4219 32897 4275 32953
rect 4343 32897 4399 32953
rect 4467 32897 4523 32953
rect 4591 32897 4647 32953
rect 4715 32897 4771 32953
rect 4839 32897 4895 32953
rect 4963 32897 5019 32953
rect 4095 32773 4151 32829
rect 4219 32773 4275 32829
rect 4343 32773 4399 32829
rect 4467 32773 4523 32829
rect 4591 32773 4647 32829
rect 4715 32773 4771 32829
rect 4839 32773 4895 32829
rect 4963 32773 5019 32829
rect 4095 32649 4151 32705
rect 4219 32649 4275 32705
rect 4343 32649 4399 32705
rect 4467 32649 4523 32705
rect 4591 32649 4647 32705
rect 4715 32649 4771 32705
rect 4839 32649 4895 32705
rect 4963 32649 5019 32705
rect 4095 32525 4151 32581
rect 4219 32525 4275 32581
rect 4343 32525 4399 32581
rect 4467 32525 4523 32581
rect 4591 32525 4647 32581
rect 4715 32525 4771 32581
rect 4839 32525 4895 32581
rect 4963 32525 5019 32581
rect 4095 32401 4151 32457
rect 4219 32401 4275 32457
rect 4343 32401 4399 32457
rect 4467 32401 4523 32457
rect 4591 32401 4647 32457
rect 4715 32401 4771 32457
rect 4839 32401 4895 32457
rect 4963 32401 5019 32457
rect 4095 32277 4151 32333
rect 4219 32277 4275 32333
rect 4343 32277 4399 32333
rect 4467 32277 4523 32333
rect 4591 32277 4647 32333
rect 4715 32277 4771 32333
rect 4839 32277 4895 32333
rect 4963 32277 5019 32333
rect 4095 32153 4151 32209
rect 4219 32153 4275 32209
rect 4343 32153 4399 32209
rect 4467 32153 4523 32209
rect 4591 32153 4647 32209
rect 4715 32153 4771 32209
rect 4839 32153 4895 32209
rect 4963 32153 5019 32209
rect 4095 32029 4151 32085
rect 4219 32029 4275 32085
rect 4343 32029 4399 32085
rect 4467 32029 4523 32085
rect 4591 32029 4647 32085
rect 4715 32029 4771 32085
rect 4839 32029 4895 32085
rect 4963 32029 5019 32085
rect 4095 31905 4151 31961
rect 4219 31905 4275 31961
rect 4343 31905 4399 31961
rect 4467 31905 4523 31961
rect 4591 31905 4647 31961
rect 4715 31905 4771 31961
rect 4839 31905 4895 31961
rect 4963 31905 5019 31961
rect 4095 31781 4151 31837
rect 4219 31781 4275 31837
rect 4343 31781 4399 31837
rect 4467 31781 4523 31837
rect 4591 31781 4647 31837
rect 4715 31781 4771 31837
rect 4839 31781 4895 31837
rect 4963 31781 5019 31837
rect 4095 31657 4151 31713
rect 4219 31657 4275 31713
rect 4343 31657 4399 31713
rect 4467 31657 4523 31713
rect 4591 31657 4647 31713
rect 4715 31657 4771 31713
rect 4839 31657 4895 31713
rect 4963 31657 5019 31713
rect 4095 31533 4151 31589
rect 4219 31533 4275 31589
rect 4343 31533 4399 31589
rect 4467 31533 4523 31589
rect 4591 31533 4647 31589
rect 4715 31533 4771 31589
rect 4839 31533 4895 31589
rect 4963 31533 5019 31589
rect 4095 31409 4151 31465
rect 4219 31409 4275 31465
rect 4343 31409 4399 31465
rect 4467 31409 4523 31465
rect 4591 31409 4647 31465
rect 4715 31409 4771 31465
rect 4839 31409 4895 31465
rect 4963 31409 5019 31465
rect 4095 31285 4151 31341
rect 4219 31285 4275 31341
rect 4343 31285 4399 31341
rect 4467 31285 4523 31341
rect 4591 31285 4647 31341
rect 4715 31285 4771 31341
rect 4839 31285 4895 31341
rect 4963 31285 5019 31341
rect 3631 30157 3687 30159
rect 3631 30105 3633 30157
rect 3633 30105 3685 30157
rect 3685 30105 3687 30157
rect 3631 30103 3687 30105
rect 3755 30157 3811 30159
rect 3755 30105 3757 30157
rect 3757 30105 3809 30157
rect 3809 30105 3811 30157
rect 3755 30103 3811 30105
rect 3879 30157 3935 30159
rect 3879 30105 3881 30157
rect 3881 30105 3933 30157
rect 3933 30105 3935 30157
rect 3879 30103 3935 30105
rect 3631 30033 3687 30035
rect 3631 29981 3633 30033
rect 3633 29981 3685 30033
rect 3685 29981 3687 30033
rect 3631 29979 3687 29981
rect 3755 30033 3811 30035
rect 3755 29981 3757 30033
rect 3757 29981 3809 30033
rect 3809 29981 3811 30033
rect 3755 29979 3811 29981
rect 3879 30033 3935 30035
rect 3879 29981 3881 30033
rect 3881 29981 3933 30033
rect 3933 29981 3935 30033
rect 3879 29979 3935 29981
rect 3631 29909 3687 29911
rect 3631 29857 3633 29909
rect 3633 29857 3685 29909
rect 3685 29857 3687 29909
rect 3631 29855 3687 29857
rect 3755 29909 3811 29911
rect 3755 29857 3757 29909
rect 3757 29857 3809 29909
rect 3809 29857 3811 29909
rect 3755 29855 3811 29857
rect 3879 29909 3935 29911
rect 3879 29857 3881 29909
rect 3881 29857 3933 29909
rect 3933 29857 3935 29909
rect 3879 29855 3935 29857
rect 3631 29785 3687 29787
rect 3631 29733 3633 29785
rect 3633 29733 3685 29785
rect 3685 29733 3687 29785
rect 3631 29731 3687 29733
rect 3755 29785 3811 29787
rect 3755 29733 3757 29785
rect 3757 29733 3809 29785
rect 3809 29733 3811 29785
rect 3755 29731 3811 29733
rect 3879 29785 3935 29787
rect 3879 29733 3881 29785
rect 3881 29733 3933 29785
rect 3933 29733 3935 29785
rect 3879 29731 3935 29733
rect 3631 29661 3687 29663
rect 3631 29609 3633 29661
rect 3633 29609 3685 29661
rect 3685 29609 3687 29661
rect 3631 29607 3687 29609
rect 3755 29661 3811 29663
rect 3755 29609 3757 29661
rect 3757 29609 3809 29661
rect 3809 29609 3811 29661
rect 3755 29607 3811 29609
rect 3879 29661 3935 29663
rect 3879 29609 3881 29661
rect 3881 29609 3933 29661
rect 3933 29609 3935 29661
rect 3879 29607 3935 29609
rect 3631 29537 3687 29539
rect 3631 29485 3633 29537
rect 3633 29485 3685 29537
rect 3685 29485 3687 29537
rect 3631 29483 3687 29485
rect 3755 29537 3811 29539
rect 3755 29485 3757 29537
rect 3757 29485 3809 29537
rect 3809 29485 3811 29537
rect 3755 29483 3811 29485
rect 3879 29537 3935 29539
rect 3879 29485 3881 29537
rect 3881 29485 3933 29537
rect 3933 29485 3935 29537
rect 3879 29483 3935 29485
rect 3631 29413 3687 29415
rect 3631 29361 3633 29413
rect 3633 29361 3685 29413
rect 3685 29361 3687 29413
rect 3631 29359 3687 29361
rect 3755 29413 3811 29415
rect 3755 29361 3757 29413
rect 3757 29361 3809 29413
rect 3809 29361 3811 29413
rect 3755 29359 3811 29361
rect 3879 29413 3935 29415
rect 3879 29361 3881 29413
rect 3881 29361 3933 29413
rect 3933 29361 3935 29413
rect 3879 29359 3935 29361
rect 3631 29289 3687 29291
rect 3631 29237 3633 29289
rect 3633 29237 3685 29289
rect 3685 29237 3687 29289
rect 3631 29235 3687 29237
rect 3755 29289 3811 29291
rect 3755 29237 3757 29289
rect 3757 29237 3809 29289
rect 3809 29237 3811 29289
rect 3755 29235 3811 29237
rect 3879 29289 3935 29291
rect 3879 29237 3881 29289
rect 3881 29237 3933 29289
rect 3933 29237 3935 29289
rect 3879 29235 3935 29237
rect 3631 29165 3687 29167
rect 3631 29113 3633 29165
rect 3633 29113 3685 29165
rect 3685 29113 3687 29165
rect 3631 29111 3687 29113
rect 3755 29165 3811 29167
rect 3755 29113 3757 29165
rect 3757 29113 3809 29165
rect 3809 29113 3811 29165
rect 3755 29111 3811 29113
rect 3879 29165 3935 29167
rect 3879 29113 3881 29165
rect 3881 29113 3933 29165
rect 3933 29113 3935 29165
rect 3879 29111 3935 29113
rect 3631 29041 3687 29043
rect 3631 28989 3633 29041
rect 3633 28989 3685 29041
rect 3685 28989 3687 29041
rect 3631 28987 3687 28989
rect 3755 29041 3811 29043
rect 3755 28989 3757 29041
rect 3757 28989 3809 29041
rect 3809 28989 3811 29041
rect 3755 28987 3811 28989
rect 3879 29041 3935 29043
rect 3879 28989 3881 29041
rect 3881 28989 3933 29041
rect 3933 28989 3935 29041
rect 3879 28987 3935 28989
rect 3631 28917 3687 28919
rect 3631 28865 3633 28917
rect 3633 28865 3685 28917
rect 3685 28865 3687 28917
rect 3631 28863 3687 28865
rect 3755 28917 3811 28919
rect 3755 28865 3757 28917
rect 3757 28865 3809 28917
rect 3809 28865 3811 28917
rect 3755 28863 3811 28865
rect 3879 28917 3935 28919
rect 3879 28865 3881 28917
rect 3881 28865 3933 28917
rect 3933 28865 3935 28917
rect 3879 28863 3935 28865
rect 3631 28793 3687 28795
rect 3631 28741 3633 28793
rect 3633 28741 3685 28793
rect 3685 28741 3687 28793
rect 3631 28739 3687 28741
rect 3755 28793 3811 28795
rect 3755 28741 3757 28793
rect 3757 28741 3809 28793
rect 3809 28741 3811 28793
rect 3755 28739 3811 28741
rect 3879 28793 3935 28795
rect 3879 28741 3881 28793
rect 3881 28741 3933 28793
rect 3933 28741 3935 28793
rect 3879 28739 3935 28741
rect 3631 28669 3687 28671
rect 3631 28617 3633 28669
rect 3633 28617 3685 28669
rect 3685 28617 3687 28669
rect 3631 28615 3687 28617
rect 3755 28669 3811 28671
rect 3755 28617 3757 28669
rect 3757 28617 3809 28669
rect 3809 28617 3811 28669
rect 3755 28615 3811 28617
rect 3879 28669 3935 28671
rect 3879 28617 3881 28669
rect 3881 28617 3933 28669
rect 3933 28617 3935 28669
rect 3879 28615 3935 28617
rect 3631 28545 3687 28547
rect 3631 28493 3633 28545
rect 3633 28493 3685 28545
rect 3685 28493 3687 28545
rect 3631 28491 3687 28493
rect 3755 28545 3811 28547
rect 3755 28493 3757 28545
rect 3757 28493 3809 28545
rect 3809 28493 3811 28545
rect 3755 28491 3811 28493
rect 3879 28545 3935 28547
rect 3879 28493 3881 28545
rect 3881 28493 3933 28545
rect 3933 28493 3935 28545
rect 3879 28491 3935 28493
rect 3631 28421 3687 28423
rect 3631 28369 3633 28421
rect 3633 28369 3685 28421
rect 3685 28369 3687 28421
rect 3631 28367 3687 28369
rect 3755 28421 3811 28423
rect 3755 28369 3757 28421
rect 3757 28369 3809 28421
rect 3809 28369 3811 28421
rect 3755 28367 3811 28369
rect 3879 28421 3935 28423
rect 3879 28369 3881 28421
rect 3881 28369 3933 28421
rect 3933 28369 3935 28421
rect 3879 28367 3935 28369
rect 4095 25635 4151 25691
rect 4219 25635 4275 25691
rect 4343 25635 4399 25691
rect 4467 25635 4523 25691
rect 4591 25635 4647 25691
rect 4715 25635 4771 25691
rect 4839 25635 4895 25691
rect 4963 25635 5019 25691
rect 4095 25511 4151 25567
rect 4219 25511 4275 25567
rect 4343 25511 4399 25567
rect 4467 25511 4523 25567
rect 4591 25511 4647 25567
rect 4715 25511 4771 25567
rect 4839 25511 4895 25567
rect 4963 25511 5019 25567
rect 4095 25387 4151 25443
rect 4219 25387 4275 25443
rect 4343 25387 4399 25443
rect 4467 25387 4523 25443
rect 4591 25387 4647 25443
rect 4715 25387 4771 25443
rect 4839 25387 4895 25443
rect 4963 25387 5019 25443
rect 4095 25263 4151 25319
rect 4219 25263 4275 25319
rect 4343 25263 4399 25319
rect 4467 25263 4523 25319
rect 4591 25263 4647 25319
rect 4715 25263 4771 25319
rect 4839 25263 4895 25319
rect 4963 25263 5019 25319
rect 4095 25139 4151 25195
rect 4219 25139 4275 25195
rect 4343 25139 4399 25195
rect 4467 25139 4523 25195
rect 4591 25139 4647 25195
rect 4715 25139 4771 25195
rect 4839 25139 4895 25195
rect 4963 25139 5019 25195
rect 4095 25015 4151 25071
rect 4219 25015 4275 25071
rect 4343 25015 4399 25071
rect 4467 25015 4523 25071
rect 4591 25015 4647 25071
rect 4715 25015 4771 25071
rect 4839 25015 4895 25071
rect 4963 25015 5019 25071
rect 4095 24891 4151 24947
rect 4219 24891 4275 24947
rect 4343 24891 4399 24947
rect 4467 24891 4523 24947
rect 4591 24891 4647 24947
rect 4715 24891 4771 24947
rect 4839 24891 4895 24947
rect 4963 24891 5019 24947
rect 4095 24767 4151 24823
rect 4219 24767 4275 24823
rect 4343 24767 4399 24823
rect 4467 24767 4523 24823
rect 4591 24767 4647 24823
rect 4715 24767 4771 24823
rect 4839 24767 4895 24823
rect 4963 24767 5019 24823
rect 3631 24062 3687 24064
rect 3631 24010 3633 24062
rect 3633 24010 3685 24062
rect 3685 24010 3687 24062
rect 3631 24008 3687 24010
rect 3755 24062 3811 24064
rect 3755 24010 3757 24062
rect 3757 24010 3809 24062
rect 3809 24010 3811 24062
rect 3755 24008 3811 24010
rect 3879 24062 3935 24064
rect 3879 24010 3881 24062
rect 3881 24010 3933 24062
rect 3933 24010 3935 24062
rect 3879 24008 3935 24010
rect 3631 23938 3687 23940
rect 3631 23886 3633 23938
rect 3633 23886 3685 23938
rect 3685 23886 3687 23938
rect 3631 23884 3687 23886
rect 3755 23938 3811 23940
rect 3755 23886 3757 23938
rect 3757 23886 3809 23938
rect 3809 23886 3811 23938
rect 3755 23884 3811 23886
rect 3879 23938 3935 23940
rect 3879 23886 3881 23938
rect 3881 23886 3933 23938
rect 3933 23886 3935 23938
rect 3879 23884 3935 23886
rect 3631 23814 3687 23816
rect 3631 23762 3633 23814
rect 3633 23762 3685 23814
rect 3685 23762 3687 23814
rect 3631 23760 3687 23762
rect 3755 23814 3811 23816
rect 3755 23762 3757 23814
rect 3757 23762 3809 23814
rect 3809 23762 3811 23814
rect 3755 23760 3811 23762
rect 3879 23814 3935 23816
rect 3879 23762 3881 23814
rect 3881 23762 3933 23814
rect 3933 23762 3935 23814
rect 3879 23760 3935 23762
rect 3631 23690 3687 23692
rect 3631 23638 3633 23690
rect 3633 23638 3685 23690
rect 3685 23638 3687 23690
rect 3631 23636 3687 23638
rect 3755 23690 3811 23692
rect 3755 23638 3757 23690
rect 3757 23638 3809 23690
rect 3809 23638 3811 23690
rect 3755 23636 3811 23638
rect 3879 23690 3935 23692
rect 3879 23638 3881 23690
rect 3881 23638 3933 23690
rect 3933 23638 3935 23690
rect 3879 23636 3935 23638
rect 3631 23566 3687 23568
rect 3631 23514 3633 23566
rect 3633 23514 3685 23566
rect 3685 23514 3687 23566
rect 3631 23512 3687 23514
rect 3755 23566 3811 23568
rect 3755 23514 3757 23566
rect 3757 23514 3809 23566
rect 3809 23514 3811 23566
rect 3755 23512 3811 23514
rect 3879 23566 3935 23568
rect 3879 23514 3881 23566
rect 3881 23514 3933 23566
rect 3933 23514 3935 23566
rect 3879 23512 3935 23514
rect 3631 23442 3687 23444
rect 3631 23390 3633 23442
rect 3633 23390 3685 23442
rect 3685 23390 3687 23442
rect 3631 23388 3687 23390
rect 3755 23442 3811 23444
rect 3755 23390 3757 23442
rect 3757 23390 3809 23442
rect 3809 23390 3811 23442
rect 3755 23388 3811 23390
rect 3879 23442 3935 23444
rect 3879 23390 3881 23442
rect 3881 23390 3933 23442
rect 3933 23390 3935 23442
rect 3879 23388 3935 23390
rect 3631 23318 3687 23320
rect 3631 23266 3633 23318
rect 3633 23266 3685 23318
rect 3685 23266 3687 23318
rect 3631 23264 3687 23266
rect 3755 23318 3811 23320
rect 3755 23266 3757 23318
rect 3757 23266 3809 23318
rect 3809 23266 3811 23318
rect 3755 23264 3811 23266
rect 3879 23318 3935 23320
rect 3879 23266 3881 23318
rect 3881 23266 3933 23318
rect 3933 23266 3935 23318
rect 3879 23264 3935 23266
rect 3631 23194 3687 23196
rect 3631 23142 3633 23194
rect 3633 23142 3685 23194
rect 3685 23142 3687 23194
rect 3631 23140 3687 23142
rect 3755 23194 3811 23196
rect 3755 23142 3757 23194
rect 3757 23142 3809 23194
rect 3809 23142 3811 23194
rect 3755 23140 3811 23142
rect 3879 23194 3935 23196
rect 3879 23142 3881 23194
rect 3881 23142 3933 23194
rect 3933 23142 3935 23194
rect 3879 23140 3935 23142
rect 4095 22456 4151 22512
rect 4219 22456 4275 22512
rect 4343 22456 4399 22512
rect 4467 22456 4523 22512
rect 4591 22456 4647 22512
rect 4715 22456 4771 22512
rect 4839 22456 4895 22512
rect 4963 22456 5019 22512
rect 4095 22332 4151 22388
rect 4219 22332 4275 22388
rect 4343 22332 4399 22388
rect 4467 22332 4523 22388
rect 4591 22332 4647 22388
rect 4715 22332 4771 22388
rect 4839 22332 4895 22388
rect 4963 22332 5019 22388
rect 4095 22208 4151 22264
rect 4219 22208 4275 22264
rect 4343 22208 4399 22264
rect 4467 22208 4523 22264
rect 4591 22208 4647 22264
rect 4715 22208 4771 22264
rect 4839 22208 4895 22264
rect 4963 22208 5019 22264
rect 4095 22084 4151 22140
rect 4219 22084 4275 22140
rect 4343 22084 4399 22140
rect 4467 22084 4523 22140
rect 4591 22084 4647 22140
rect 4715 22084 4771 22140
rect 4839 22084 4895 22140
rect 4963 22084 5019 22140
rect 4095 21960 4151 22016
rect 4219 21960 4275 22016
rect 4343 21960 4399 22016
rect 4467 21960 4523 22016
rect 4591 21960 4647 22016
rect 4715 21960 4771 22016
rect 4839 21960 4895 22016
rect 4963 21960 5019 22016
rect 4095 21836 4151 21892
rect 4219 21836 4275 21892
rect 4343 21836 4399 21892
rect 4467 21836 4523 21892
rect 4591 21836 4647 21892
rect 4715 21836 4771 21892
rect 4839 21836 4895 21892
rect 4963 21836 5019 21892
rect 4095 21712 4151 21768
rect 4219 21712 4275 21768
rect 4343 21712 4399 21768
rect 4467 21712 4523 21768
rect 4591 21712 4647 21768
rect 4715 21712 4771 21768
rect 4839 21712 4895 21768
rect 4963 21712 5019 21768
rect 4095 21588 4151 21644
rect 4219 21588 4275 21644
rect 4343 21588 4399 21644
rect 4467 21588 4523 21644
rect 4591 21588 4647 21644
rect 4715 21588 4771 21644
rect 4839 21588 4895 21644
rect 4963 21588 5019 21644
rect 4095 21464 4151 21520
rect 4219 21464 4275 21520
rect 4343 21464 4399 21520
rect 4467 21464 4523 21520
rect 4591 21464 4647 21520
rect 4715 21464 4771 21520
rect 4839 21464 4895 21520
rect 4963 21464 5019 21520
rect 4095 21340 4151 21396
rect 4219 21340 4275 21396
rect 4343 21340 4399 21396
rect 4467 21340 4523 21396
rect 4591 21340 4647 21396
rect 4715 21340 4771 21396
rect 4839 21340 4895 21396
rect 4963 21340 5019 21396
rect 4095 21216 4151 21272
rect 4219 21216 4275 21272
rect 4343 21216 4399 21272
rect 4467 21216 4523 21272
rect 4591 21216 4647 21272
rect 4715 21216 4771 21272
rect 4839 21216 4895 21272
rect 4963 21216 5019 21272
rect 4095 21092 4151 21148
rect 4219 21092 4275 21148
rect 4343 21092 4399 21148
rect 4467 21092 4523 21148
rect 4591 21092 4647 21148
rect 4715 21092 4771 21148
rect 4839 21092 4895 21148
rect 4963 21092 5019 21148
rect 4095 20968 4151 21024
rect 4219 20968 4275 21024
rect 4343 20968 4399 21024
rect 4467 20968 4523 21024
rect 4591 20968 4647 21024
rect 4715 20968 4771 21024
rect 4839 20968 4895 21024
rect 4963 20968 5019 21024
rect 4095 20844 4151 20900
rect 4219 20844 4275 20900
rect 4343 20844 4399 20900
rect 4467 20844 4523 20900
rect 4591 20844 4647 20900
rect 4715 20844 4771 20900
rect 4839 20844 4895 20900
rect 4963 20844 5019 20900
rect 4095 20720 4151 20776
rect 4219 20720 4275 20776
rect 4343 20720 4399 20776
rect 4467 20720 4523 20776
rect 4591 20720 4647 20776
rect 4715 20720 4771 20776
rect 4839 20720 4895 20776
rect 4963 20720 5019 20776
rect 4095 20596 4151 20652
rect 4219 20596 4275 20652
rect 4343 20596 4399 20652
rect 4467 20596 4523 20652
rect 4591 20596 4647 20652
rect 4715 20596 4771 20652
rect 4839 20596 4895 20652
rect 4963 20596 5019 20652
rect 4095 20472 4151 20528
rect 4219 20472 4275 20528
rect 4343 20472 4399 20528
rect 4467 20472 4523 20528
rect 4591 20472 4647 20528
rect 4715 20472 4771 20528
rect 4839 20472 4895 20528
rect 4963 20472 5019 20528
rect 4095 20348 4151 20404
rect 4219 20348 4275 20404
rect 4343 20348 4399 20404
rect 4467 20348 4523 20404
rect 4591 20348 4647 20404
rect 4715 20348 4771 20404
rect 4839 20348 4895 20404
rect 4963 20348 5019 20404
rect 4095 20224 4151 20280
rect 4219 20224 4275 20280
rect 4343 20224 4399 20280
rect 4467 20224 4523 20280
rect 4591 20224 4647 20280
rect 4715 20224 4771 20280
rect 4839 20224 4895 20280
rect 4963 20224 5019 20280
rect 4095 20100 4151 20156
rect 4219 20100 4275 20156
rect 4343 20100 4399 20156
rect 4467 20100 4523 20156
rect 4591 20100 4647 20156
rect 4715 20100 4771 20156
rect 4839 20100 4895 20156
rect 4963 20100 5019 20156
rect 4095 19976 4151 20032
rect 4219 19976 4275 20032
rect 4343 19976 4399 20032
rect 4467 19976 4523 20032
rect 4591 19976 4647 20032
rect 4715 19976 4771 20032
rect 4839 19976 4895 20032
rect 4963 19976 5019 20032
rect 4095 19852 4151 19908
rect 4219 19852 4275 19908
rect 4343 19852 4399 19908
rect 4467 19852 4523 19908
rect 4591 19852 4647 19908
rect 4715 19852 4771 19908
rect 4839 19852 4895 19908
rect 4963 19852 5019 19908
rect 3631 19505 3687 19507
rect 3631 19453 3633 19505
rect 3633 19453 3685 19505
rect 3685 19453 3687 19505
rect 3631 19451 3687 19453
rect 3755 19505 3811 19507
rect 3755 19453 3757 19505
rect 3757 19453 3809 19505
rect 3809 19453 3811 19505
rect 3755 19451 3811 19453
rect 3879 19505 3935 19507
rect 3879 19453 3881 19505
rect 3881 19453 3933 19505
rect 3933 19453 3935 19505
rect 3879 19451 3935 19453
rect 3631 19381 3687 19383
rect 3631 19329 3633 19381
rect 3633 19329 3685 19381
rect 3685 19329 3687 19381
rect 3631 19327 3687 19329
rect 3755 19381 3811 19383
rect 3755 19329 3757 19381
rect 3757 19329 3809 19381
rect 3809 19329 3811 19381
rect 3755 19327 3811 19329
rect 3879 19381 3935 19383
rect 3879 19329 3881 19381
rect 3881 19329 3933 19381
rect 3933 19329 3935 19381
rect 3879 19327 3935 19329
rect 3631 19257 3687 19259
rect 3631 19205 3633 19257
rect 3633 19205 3685 19257
rect 3685 19205 3687 19257
rect 3631 19203 3687 19205
rect 3755 19257 3811 19259
rect 3755 19205 3757 19257
rect 3757 19205 3809 19257
rect 3809 19205 3811 19257
rect 3755 19203 3811 19205
rect 3879 19257 3935 19259
rect 3879 19205 3881 19257
rect 3881 19205 3933 19257
rect 3933 19205 3935 19257
rect 3879 19203 3935 19205
rect 3631 19133 3687 19135
rect 3631 19081 3633 19133
rect 3633 19081 3685 19133
rect 3685 19081 3687 19133
rect 3631 19079 3687 19081
rect 3755 19133 3811 19135
rect 3755 19081 3757 19133
rect 3757 19081 3809 19133
rect 3809 19081 3811 19133
rect 3755 19079 3811 19081
rect 3879 19133 3935 19135
rect 3879 19081 3881 19133
rect 3881 19081 3933 19133
rect 3933 19081 3935 19133
rect 3879 19079 3935 19081
rect 3631 19009 3687 19011
rect 3631 18957 3633 19009
rect 3633 18957 3685 19009
rect 3685 18957 3687 19009
rect 3631 18955 3687 18957
rect 3755 19009 3811 19011
rect 3755 18957 3757 19009
rect 3757 18957 3809 19009
rect 3809 18957 3811 19009
rect 3755 18955 3811 18957
rect 3879 19009 3935 19011
rect 3879 18957 3881 19009
rect 3881 18957 3933 19009
rect 3933 18957 3935 19009
rect 3879 18955 3935 18957
rect 3631 18885 3687 18887
rect 3631 18833 3633 18885
rect 3633 18833 3685 18885
rect 3685 18833 3687 18885
rect 3631 18831 3687 18833
rect 3755 18885 3811 18887
rect 3755 18833 3757 18885
rect 3757 18833 3809 18885
rect 3809 18833 3811 18885
rect 3755 18831 3811 18833
rect 3879 18885 3935 18887
rect 3879 18833 3881 18885
rect 3881 18833 3933 18885
rect 3933 18833 3935 18885
rect 3879 18831 3935 18833
rect 3631 18761 3687 18763
rect 3631 18709 3633 18761
rect 3633 18709 3685 18761
rect 3685 18709 3687 18761
rect 3631 18707 3687 18709
rect 3755 18761 3811 18763
rect 3755 18709 3757 18761
rect 3757 18709 3809 18761
rect 3809 18709 3811 18761
rect 3755 18707 3811 18709
rect 3879 18761 3935 18763
rect 3879 18709 3881 18761
rect 3881 18709 3933 18761
rect 3933 18709 3935 18761
rect 3879 18707 3935 18709
rect 3631 18637 3687 18639
rect 3631 18585 3633 18637
rect 3633 18585 3685 18637
rect 3685 18585 3687 18637
rect 3631 18583 3687 18585
rect 3755 18637 3811 18639
rect 3755 18585 3757 18637
rect 3757 18585 3809 18637
rect 3809 18585 3811 18637
rect 3755 18583 3811 18585
rect 3879 18637 3935 18639
rect 3879 18585 3881 18637
rect 3881 18585 3933 18637
rect 3933 18585 3935 18637
rect 3879 18583 3935 18585
rect 3631 18513 3687 18515
rect 3631 18461 3633 18513
rect 3633 18461 3685 18513
rect 3685 18461 3687 18513
rect 3631 18459 3687 18461
rect 3755 18513 3811 18515
rect 3755 18461 3757 18513
rect 3757 18461 3809 18513
rect 3809 18461 3811 18513
rect 3755 18459 3811 18461
rect 3879 18513 3935 18515
rect 3879 18461 3881 18513
rect 3881 18461 3933 18513
rect 3933 18461 3935 18513
rect 3879 18459 3935 18461
rect 3631 18389 3687 18391
rect 3631 18337 3633 18389
rect 3633 18337 3685 18389
rect 3685 18337 3687 18389
rect 3631 18335 3687 18337
rect 3755 18389 3811 18391
rect 3755 18337 3757 18389
rect 3757 18337 3809 18389
rect 3809 18337 3811 18389
rect 3755 18335 3811 18337
rect 3879 18389 3935 18391
rect 3879 18337 3881 18389
rect 3881 18337 3933 18389
rect 3933 18337 3935 18389
rect 3879 18335 3935 18337
rect 3631 18265 3687 18267
rect 3631 18213 3633 18265
rect 3633 18213 3685 18265
rect 3685 18213 3687 18265
rect 3631 18211 3687 18213
rect 3755 18265 3811 18267
rect 3755 18213 3757 18265
rect 3757 18213 3809 18265
rect 3809 18213 3811 18265
rect 3755 18211 3811 18213
rect 3879 18265 3935 18267
rect 3879 18213 3881 18265
rect 3881 18213 3933 18265
rect 3933 18213 3935 18265
rect 3879 18211 3935 18213
rect 3631 18141 3687 18143
rect 3631 18089 3633 18141
rect 3633 18089 3685 18141
rect 3685 18089 3687 18141
rect 3631 18087 3687 18089
rect 3755 18141 3811 18143
rect 3755 18089 3757 18141
rect 3757 18089 3809 18141
rect 3809 18089 3811 18141
rect 3755 18087 3811 18089
rect 3879 18141 3935 18143
rect 3879 18089 3881 18141
rect 3881 18089 3933 18141
rect 3933 18089 3935 18141
rect 3879 18087 3935 18089
rect 3631 18017 3687 18019
rect 3631 17965 3633 18017
rect 3633 17965 3685 18017
rect 3685 17965 3687 18017
rect 3631 17963 3687 17965
rect 3755 18017 3811 18019
rect 3755 17965 3757 18017
rect 3757 17965 3809 18017
rect 3809 17965 3811 18017
rect 3755 17963 3811 17965
rect 3879 18017 3935 18019
rect 3879 17965 3881 18017
rect 3881 17965 3933 18017
rect 3933 17965 3935 18017
rect 3879 17963 3935 17965
rect 3631 17893 3687 17895
rect 3631 17841 3633 17893
rect 3633 17841 3685 17893
rect 3685 17841 3687 17893
rect 3631 17839 3687 17841
rect 3755 17893 3811 17895
rect 3755 17841 3757 17893
rect 3757 17841 3809 17893
rect 3809 17841 3811 17893
rect 3755 17839 3811 17841
rect 3879 17893 3935 17895
rect 3879 17841 3881 17893
rect 3881 17841 3933 17893
rect 3933 17841 3935 17893
rect 3879 17839 3935 17841
rect 3631 17769 3687 17771
rect 3631 17717 3633 17769
rect 3633 17717 3685 17769
rect 3685 17717 3687 17769
rect 3631 17715 3687 17717
rect 3755 17769 3811 17771
rect 3755 17717 3757 17769
rect 3757 17717 3809 17769
rect 3809 17717 3811 17769
rect 3755 17715 3811 17717
rect 3879 17769 3935 17771
rect 3879 17717 3881 17769
rect 3881 17717 3933 17769
rect 3933 17717 3935 17769
rect 3879 17715 3935 17717
rect 3631 17645 3687 17647
rect 3631 17593 3633 17645
rect 3633 17593 3685 17645
rect 3685 17593 3687 17645
rect 3631 17591 3687 17593
rect 3755 17645 3811 17647
rect 3755 17593 3757 17645
rect 3757 17593 3809 17645
rect 3809 17593 3811 17645
rect 3755 17591 3811 17593
rect 3879 17645 3935 17647
rect 3879 17593 3881 17645
rect 3881 17593 3933 17645
rect 3933 17593 3935 17645
rect 3879 17591 3935 17593
rect 3631 17521 3687 17523
rect 3631 17469 3633 17521
rect 3633 17469 3685 17521
rect 3685 17469 3687 17521
rect 3631 17467 3687 17469
rect 3755 17521 3811 17523
rect 3755 17469 3757 17521
rect 3757 17469 3809 17521
rect 3809 17469 3811 17521
rect 3755 17467 3811 17469
rect 3879 17521 3935 17523
rect 3879 17469 3881 17521
rect 3881 17469 3933 17521
rect 3933 17469 3935 17521
rect 3879 17467 3935 17469
rect 3631 17397 3687 17399
rect 3631 17345 3633 17397
rect 3633 17345 3685 17397
rect 3685 17345 3687 17397
rect 3631 17343 3687 17345
rect 3755 17397 3811 17399
rect 3755 17345 3757 17397
rect 3757 17345 3809 17397
rect 3809 17345 3811 17397
rect 3755 17343 3811 17345
rect 3879 17397 3935 17399
rect 3879 17345 3881 17397
rect 3881 17345 3933 17397
rect 3933 17345 3935 17397
rect 3879 17343 3935 17345
rect 3631 17273 3687 17275
rect 3631 17221 3633 17273
rect 3633 17221 3685 17273
rect 3685 17221 3687 17273
rect 3631 17219 3687 17221
rect 3755 17273 3811 17275
rect 3755 17221 3757 17273
rect 3757 17221 3809 17273
rect 3809 17221 3811 17273
rect 3755 17219 3811 17221
rect 3879 17273 3935 17275
rect 3879 17221 3881 17273
rect 3881 17221 3933 17273
rect 3933 17221 3935 17273
rect 3879 17219 3935 17221
rect 3631 17149 3687 17151
rect 3631 17097 3633 17149
rect 3633 17097 3685 17149
rect 3685 17097 3687 17149
rect 3631 17095 3687 17097
rect 3755 17149 3811 17151
rect 3755 17097 3757 17149
rect 3757 17097 3809 17149
rect 3809 17097 3811 17149
rect 3755 17095 3811 17097
rect 3879 17149 3935 17151
rect 3879 17097 3881 17149
rect 3881 17097 3933 17149
rect 3933 17097 3935 17149
rect 3879 17095 3935 17097
rect 3631 17025 3687 17027
rect 3631 16973 3633 17025
rect 3633 16973 3685 17025
rect 3685 16973 3687 17025
rect 3631 16971 3687 16973
rect 3755 17025 3811 17027
rect 3755 16973 3757 17025
rect 3757 16973 3809 17025
rect 3809 16973 3811 17025
rect 3755 16971 3811 16973
rect 3879 17025 3935 17027
rect 3879 16973 3881 17025
rect 3881 16973 3933 17025
rect 3933 16973 3935 17025
rect 3879 16971 3935 16973
rect 3631 16901 3687 16903
rect 3631 16849 3633 16901
rect 3633 16849 3685 16901
rect 3685 16849 3687 16901
rect 3631 16847 3687 16849
rect 3755 16901 3811 16903
rect 3755 16849 3757 16901
rect 3757 16849 3809 16901
rect 3809 16849 3811 16901
rect 3755 16847 3811 16849
rect 3879 16901 3935 16903
rect 3879 16849 3881 16901
rect 3881 16849 3933 16901
rect 3933 16849 3935 16901
rect 3879 16847 3935 16849
rect 3631 16777 3687 16779
rect 3631 16725 3633 16777
rect 3633 16725 3685 16777
rect 3685 16725 3687 16777
rect 3631 16723 3687 16725
rect 3755 16777 3811 16779
rect 3755 16725 3757 16777
rect 3757 16725 3809 16777
rect 3809 16725 3811 16777
rect 3755 16723 3811 16725
rect 3879 16777 3935 16779
rect 3879 16725 3881 16777
rect 3881 16725 3933 16777
rect 3933 16725 3935 16777
rect 3879 16723 3935 16725
rect 3631 16653 3687 16655
rect 3631 16601 3633 16653
rect 3633 16601 3685 16653
rect 3685 16601 3687 16653
rect 3631 16599 3687 16601
rect 3755 16653 3811 16655
rect 3755 16601 3757 16653
rect 3757 16601 3809 16653
rect 3809 16601 3811 16653
rect 3755 16599 3811 16601
rect 3879 16653 3935 16655
rect 3879 16601 3881 16653
rect 3881 16601 3933 16653
rect 3933 16601 3935 16653
rect 3879 16599 3935 16601
rect 3631 16529 3687 16531
rect 3631 16477 3633 16529
rect 3633 16477 3685 16529
rect 3685 16477 3687 16529
rect 3631 16475 3687 16477
rect 3755 16529 3811 16531
rect 3755 16477 3757 16529
rect 3757 16477 3809 16529
rect 3809 16477 3811 16529
rect 3755 16475 3811 16477
rect 3879 16529 3935 16531
rect 3879 16477 3881 16529
rect 3881 16477 3933 16529
rect 3933 16477 3935 16529
rect 3879 16475 3935 16477
rect 3631 16405 3687 16407
rect 3631 16353 3633 16405
rect 3633 16353 3685 16405
rect 3685 16353 3687 16405
rect 3631 16351 3687 16353
rect 3755 16405 3811 16407
rect 3755 16353 3757 16405
rect 3757 16353 3809 16405
rect 3809 16353 3811 16405
rect 3755 16351 3811 16353
rect 3879 16405 3935 16407
rect 3879 16353 3881 16405
rect 3881 16353 3933 16405
rect 3933 16353 3935 16405
rect 3879 16351 3935 16353
rect 3631 16281 3687 16283
rect 3631 16229 3633 16281
rect 3633 16229 3685 16281
rect 3685 16229 3687 16281
rect 3631 16227 3687 16229
rect 3755 16281 3811 16283
rect 3755 16229 3757 16281
rect 3757 16229 3809 16281
rect 3809 16229 3811 16281
rect 3755 16227 3811 16229
rect 3879 16281 3935 16283
rect 3879 16229 3881 16281
rect 3881 16229 3933 16281
rect 3933 16229 3935 16281
rect 3879 16227 3935 16229
rect 4095 15886 4151 15942
rect 4219 15886 4275 15942
rect 4343 15886 4399 15942
rect 4467 15886 4523 15942
rect 4591 15886 4647 15942
rect 4715 15886 4771 15942
rect 4839 15886 4895 15942
rect 4963 15886 5019 15942
rect 4095 15762 4151 15818
rect 4219 15762 4275 15818
rect 4343 15762 4399 15818
rect 4467 15762 4523 15818
rect 4591 15762 4647 15818
rect 4715 15762 4771 15818
rect 4839 15762 4895 15818
rect 4963 15762 5019 15818
rect 4095 15638 4151 15694
rect 4219 15638 4275 15694
rect 4343 15638 4399 15694
rect 4467 15638 4523 15694
rect 4591 15638 4647 15694
rect 4715 15638 4771 15694
rect 4839 15638 4895 15694
rect 4963 15638 5019 15694
rect 4095 15514 4151 15570
rect 4219 15514 4275 15570
rect 4343 15514 4399 15570
rect 4467 15514 4523 15570
rect 4591 15514 4647 15570
rect 4715 15514 4771 15570
rect 4839 15514 4895 15570
rect 4963 15514 5019 15570
rect 4095 15390 4151 15446
rect 4219 15390 4275 15446
rect 4343 15390 4399 15446
rect 4467 15390 4523 15446
rect 4591 15390 4647 15446
rect 4715 15390 4771 15446
rect 4839 15390 4895 15446
rect 4963 15390 5019 15446
rect 4095 15266 4151 15322
rect 4219 15266 4275 15322
rect 4343 15266 4399 15322
rect 4467 15266 4523 15322
rect 4591 15266 4647 15322
rect 4715 15266 4771 15322
rect 4839 15266 4895 15322
rect 4963 15266 5019 15322
rect 4095 15142 4151 15198
rect 4219 15142 4275 15198
rect 4343 15142 4399 15198
rect 4467 15142 4523 15198
rect 4591 15142 4647 15198
rect 4715 15142 4771 15198
rect 4839 15142 4895 15198
rect 4963 15142 5019 15198
rect 4095 15018 4151 15074
rect 4219 15018 4275 15074
rect 4343 15018 4399 15074
rect 4467 15018 4523 15074
rect 4591 15018 4647 15074
rect 4715 15018 4771 15074
rect 4839 15018 4895 15074
rect 4963 15018 5019 15074
rect 4095 14894 4151 14950
rect 4219 14894 4275 14950
rect 4343 14894 4399 14950
rect 4467 14894 4523 14950
rect 4591 14894 4647 14950
rect 4715 14894 4771 14950
rect 4839 14894 4895 14950
rect 4963 14894 5019 14950
rect 4095 14770 4151 14826
rect 4219 14770 4275 14826
rect 4343 14770 4399 14826
rect 4467 14770 4523 14826
rect 4591 14770 4647 14826
rect 4715 14770 4771 14826
rect 4839 14770 4895 14826
rect 4963 14770 5019 14826
rect 4095 14646 4151 14702
rect 4219 14646 4275 14702
rect 4343 14646 4399 14702
rect 4467 14646 4523 14702
rect 4591 14646 4647 14702
rect 4715 14646 4771 14702
rect 4839 14646 4895 14702
rect 4963 14646 5019 14702
rect 4095 14522 4151 14578
rect 4219 14522 4275 14578
rect 4343 14522 4399 14578
rect 4467 14522 4523 14578
rect 4591 14522 4647 14578
rect 4715 14522 4771 14578
rect 4839 14522 4895 14578
rect 4963 14522 5019 14578
rect 4095 14398 4151 14454
rect 4219 14398 4275 14454
rect 4343 14398 4399 14454
rect 4467 14398 4523 14454
rect 4591 14398 4647 14454
rect 4715 14398 4771 14454
rect 4839 14398 4895 14454
rect 4963 14398 5019 14454
rect 4095 14274 4151 14330
rect 4219 14274 4275 14330
rect 4343 14274 4399 14330
rect 4467 14274 4523 14330
rect 4591 14274 4647 14330
rect 4715 14274 4771 14330
rect 4839 14274 4895 14330
rect 4963 14274 5019 14330
rect 4095 14150 4151 14206
rect 4219 14150 4275 14206
rect 4343 14150 4399 14206
rect 4467 14150 4523 14206
rect 4591 14150 4647 14206
rect 4715 14150 4771 14206
rect 4839 14150 4895 14206
rect 4963 14150 5019 14206
rect 4095 14026 4151 14082
rect 4219 14026 4275 14082
rect 4343 14026 4399 14082
rect 4467 14026 4523 14082
rect 4591 14026 4647 14082
rect 4715 14026 4771 14082
rect 4839 14026 4895 14082
rect 4963 14026 5019 14082
rect 4095 13902 4151 13958
rect 4219 13902 4275 13958
rect 4343 13902 4399 13958
rect 4467 13902 4523 13958
rect 4591 13902 4647 13958
rect 4715 13902 4771 13958
rect 4839 13902 4895 13958
rect 4963 13902 5019 13958
rect 3631 13226 3687 13228
rect 3631 13174 3633 13226
rect 3633 13174 3685 13226
rect 3685 13174 3687 13226
rect 3631 13172 3687 13174
rect 3755 13226 3811 13228
rect 3755 13174 3757 13226
rect 3757 13174 3809 13226
rect 3809 13174 3811 13226
rect 3755 13172 3811 13174
rect 3879 13226 3935 13228
rect 3879 13174 3881 13226
rect 3881 13174 3933 13226
rect 3933 13174 3935 13226
rect 3879 13172 3935 13174
rect 3631 13102 3687 13104
rect 3631 13050 3633 13102
rect 3633 13050 3685 13102
rect 3685 13050 3687 13102
rect 3631 13048 3687 13050
rect 3755 13102 3811 13104
rect 3755 13050 3757 13102
rect 3757 13050 3809 13102
rect 3809 13050 3811 13102
rect 3755 13048 3811 13050
rect 3879 13102 3935 13104
rect 3879 13050 3881 13102
rect 3881 13050 3933 13102
rect 3933 13050 3935 13102
rect 3879 13048 3935 13050
rect 3631 12978 3687 12980
rect 3631 12926 3633 12978
rect 3633 12926 3685 12978
rect 3685 12926 3687 12978
rect 3631 12924 3687 12926
rect 3755 12978 3811 12980
rect 3755 12926 3757 12978
rect 3757 12926 3809 12978
rect 3809 12926 3811 12978
rect 3755 12924 3811 12926
rect 3879 12978 3935 12980
rect 3879 12926 3881 12978
rect 3881 12926 3933 12978
rect 3933 12926 3935 12978
rect 3879 12924 3935 12926
rect 3631 12854 3687 12856
rect 3631 12802 3633 12854
rect 3633 12802 3685 12854
rect 3685 12802 3687 12854
rect 3631 12800 3687 12802
rect 3755 12854 3811 12856
rect 3755 12802 3757 12854
rect 3757 12802 3809 12854
rect 3809 12802 3811 12854
rect 3755 12800 3811 12802
rect 3879 12854 3935 12856
rect 3879 12802 3881 12854
rect 3881 12802 3933 12854
rect 3933 12802 3935 12854
rect 3879 12800 3935 12802
rect 3631 12730 3687 12732
rect 3631 12678 3633 12730
rect 3633 12678 3685 12730
rect 3685 12678 3687 12730
rect 3631 12676 3687 12678
rect 3755 12730 3811 12732
rect 3755 12678 3757 12730
rect 3757 12678 3809 12730
rect 3809 12678 3811 12730
rect 3755 12676 3811 12678
rect 3879 12730 3935 12732
rect 3879 12678 3881 12730
rect 3881 12678 3933 12730
rect 3933 12678 3935 12730
rect 3879 12676 3935 12678
rect 3631 12606 3687 12608
rect 3631 12554 3633 12606
rect 3633 12554 3685 12606
rect 3685 12554 3687 12606
rect 3631 12552 3687 12554
rect 3755 12606 3811 12608
rect 3755 12554 3757 12606
rect 3757 12554 3809 12606
rect 3809 12554 3811 12606
rect 3755 12552 3811 12554
rect 3879 12606 3935 12608
rect 3879 12554 3881 12606
rect 3881 12554 3933 12606
rect 3933 12554 3935 12606
rect 3879 12552 3935 12554
rect 3631 12482 3687 12484
rect 3631 12430 3633 12482
rect 3633 12430 3685 12482
rect 3685 12430 3687 12482
rect 3631 12428 3687 12430
rect 3755 12482 3811 12484
rect 3755 12430 3757 12482
rect 3757 12430 3809 12482
rect 3809 12430 3811 12482
rect 3755 12428 3811 12430
rect 3879 12482 3935 12484
rect 3879 12430 3881 12482
rect 3881 12430 3933 12482
rect 3933 12430 3935 12482
rect 3879 12428 3935 12430
rect 3631 12358 3687 12360
rect 3631 12306 3633 12358
rect 3633 12306 3685 12358
rect 3685 12306 3687 12358
rect 3631 12304 3687 12306
rect 3755 12358 3811 12360
rect 3755 12306 3757 12358
rect 3757 12306 3809 12358
rect 3809 12306 3811 12358
rect 3755 12304 3811 12306
rect 3879 12358 3935 12360
rect 3879 12306 3881 12358
rect 3881 12306 3933 12358
rect 3933 12306 3935 12358
rect 3879 12304 3935 12306
rect 3631 12234 3687 12236
rect 3631 12182 3633 12234
rect 3633 12182 3685 12234
rect 3685 12182 3687 12234
rect 3631 12180 3687 12182
rect 3755 12234 3811 12236
rect 3755 12182 3757 12234
rect 3757 12182 3809 12234
rect 3809 12182 3811 12234
rect 3755 12180 3811 12182
rect 3879 12234 3935 12236
rect 3879 12182 3881 12234
rect 3881 12182 3933 12234
rect 3933 12182 3935 12234
rect 3879 12180 3935 12182
rect 3631 12110 3687 12112
rect 3631 12058 3633 12110
rect 3633 12058 3685 12110
rect 3685 12058 3687 12110
rect 3631 12056 3687 12058
rect 3755 12110 3811 12112
rect 3755 12058 3757 12110
rect 3757 12058 3809 12110
rect 3809 12058 3811 12110
rect 3755 12056 3811 12058
rect 3879 12110 3935 12112
rect 3879 12058 3881 12110
rect 3881 12058 3933 12110
rect 3933 12058 3935 12110
rect 3879 12056 3935 12058
rect 4095 11236 4151 11292
rect 4219 11236 4275 11292
rect 4343 11236 4399 11292
rect 4467 11236 4523 11292
rect 4591 11236 4647 11292
rect 4715 11236 4771 11292
rect 4839 11236 4895 11292
rect 4963 11236 5019 11292
rect 4095 11112 4151 11168
rect 4219 11112 4275 11168
rect 4343 11112 4399 11168
rect 4467 11112 4523 11168
rect 4591 11112 4647 11168
rect 4715 11112 4771 11168
rect 4839 11112 4895 11168
rect 4963 11112 5019 11168
rect 4095 10988 4151 11044
rect 4219 10988 4275 11044
rect 4343 10988 4399 11044
rect 4467 10988 4523 11044
rect 4591 10988 4647 11044
rect 4715 10988 4771 11044
rect 4839 10988 4895 11044
rect 4963 10988 5019 11044
rect 4095 10864 4151 10920
rect 4219 10864 4275 10920
rect 4343 10864 4399 10920
rect 4467 10864 4523 10920
rect 4591 10864 4647 10920
rect 4715 10864 4771 10920
rect 4839 10864 4895 10920
rect 4963 10864 5019 10920
rect 4095 10740 4151 10796
rect 4219 10740 4275 10796
rect 4343 10740 4399 10796
rect 4467 10740 4523 10796
rect 4591 10740 4647 10796
rect 4715 10740 4771 10796
rect 4839 10740 4895 10796
rect 4963 10740 5019 10796
rect 4095 10616 4151 10672
rect 4219 10616 4275 10672
rect 4343 10616 4399 10672
rect 4467 10616 4523 10672
rect 4591 10616 4647 10672
rect 4715 10616 4771 10672
rect 4839 10616 4895 10672
rect 4963 10616 5019 10672
rect 4095 10492 4151 10548
rect 4219 10492 4275 10548
rect 4343 10492 4399 10548
rect 4467 10492 4523 10548
rect 4591 10492 4647 10548
rect 4715 10492 4771 10548
rect 4839 10492 4895 10548
rect 4963 10492 5019 10548
rect 4095 10368 4151 10424
rect 4219 10368 4275 10424
rect 4343 10368 4399 10424
rect 4467 10368 4523 10424
rect 4591 10368 4647 10424
rect 4715 10368 4771 10424
rect 4839 10368 4895 10424
rect 4963 10368 5019 10424
rect 4095 10244 4151 10300
rect 4219 10244 4275 10300
rect 4343 10244 4399 10300
rect 4467 10244 4523 10300
rect 4591 10244 4647 10300
rect 4715 10244 4771 10300
rect 4839 10244 4895 10300
rect 4963 10244 5019 10300
rect 4095 10120 4151 10176
rect 4219 10120 4275 10176
rect 4343 10120 4399 10176
rect 4467 10120 4523 10176
rect 4591 10120 4647 10176
rect 4715 10120 4771 10176
rect 4839 10120 4895 10176
rect 4963 10120 5019 10176
rect 4095 9996 4151 10052
rect 4219 9996 4275 10052
rect 4343 9996 4399 10052
rect 4467 9996 4523 10052
rect 4591 9996 4647 10052
rect 4715 9996 4771 10052
rect 4839 9996 4895 10052
rect 4963 9996 5019 10052
rect 3631 9390 3687 9392
rect 3631 9338 3633 9390
rect 3633 9338 3685 9390
rect 3685 9338 3687 9390
rect 3631 9336 3687 9338
rect 3755 9390 3811 9392
rect 3755 9338 3757 9390
rect 3757 9338 3809 9390
rect 3809 9338 3811 9390
rect 3755 9336 3811 9338
rect 3879 9390 3935 9392
rect 3879 9338 3881 9390
rect 3881 9338 3933 9390
rect 3933 9338 3935 9390
rect 3879 9336 3935 9338
rect 3631 9266 3687 9268
rect 3631 9214 3633 9266
rect 3633 9214 3685 9266
rect 3685 9214 3687 9266
rect 3631 9212 3687 9214
rect 3755 9266 3811 9268
rect 3755 9214 3757 9266
rect 3757 9214 3809 9266
rect 3809 9214 3811 9266
rect 3755 9212 3811 9214
rect 3879 9266 3935 9268
rect 3879 9214 3881 9266
rect 3881 9214 3933 9266
rect 3933 9214 3935 9266
rect 3879 9212 3935 9214
rect 3631 9142 3687 9144
rect 3631 9090 3633 9142
rect 3633 9090 3685 9142
rect 3685 9090 3687 9142
rect 3631 9088 3687 9090
rect 3755 9142 3811 9144
rect 3755 9090 3757 9142
rect 3757 9090 3809 9142
rect 3809 9090 3811 9142
rect 3755 9088 3811 9090
rect 3879 9142 3935 9144
rect 3879 9090 3881 9142
rect 3881 9090 3933 9142
rect 3933 9090 3935 9142
rect 3879 9088 3935 9090
rect 3631 9018 3687 9020
rect 3631 8966 3633 9018
rect 3633 8966 3685 9018
rect 3685 8966 3687 9018
rect 3631 8964 3687 8966
rect 3755 9018 3811 9020
rect 3755 8966 3757 9018
rect 3757 8966 3809 9018
rect 3809 8966 3811 9018
rect 3755 8964 3811 8966
rect 3879 9018 3935 9020
rect 3879 8966 3881 9018
rect 3881 8966 3933 9018
rect 3933 8966 3935 9018
rect 3879 8964 3935 8966
rect 3631 8894 3687 8896
rect 3631 8842 3633 8894
rect 3633 8842 3685 8894
rect 3685 8842 3687 8894
rect 3631 8840 3687 8842
rect 3755 8894 3811 8896
rect 3755 8842 3757 8894
rect 3757 8842 3809 8894
rect 3809 8842 3811 8894
rect 3755 8840 3811 8842
rect 3879 8894 3935 8896
rect 3879 8842 3881 8894
rect 3881 8842 3933 8894
rect 3933 8842 3935 8894
rect 3879 8840 3935 8842
rect 3631 8770 3687 8772
rect 3631 8718 3633 8770
rect 3633 8718 3685 8770
rect 3685 8718 3687 8770
rect 3631 8716 3687 8718
rect 3755 8770 3811 8772
rect 3755 8718 3757 8770
rect 3757 8718 3809 8770
rect 3809 8718 3811 8770
rect 3755 8716 3811 8718
rect 3879 8770 3935 8772
rect 3879 8718 3881 8770
rect 3881 8718 3933 8770
rect 3933 8718 3935 8770
rect 3879 8716 3935 8718
rect 3631 8646 3687 8648
rect 3631 8594 3633 8646
rect 3633 8594 3685 8646
rect 3685 8594 3687 8646
rect 3631 8592 3687 8594
rect 3755 8646 3811 8648
rect 3755 8594 3757 8646
rect 3757 8594 3809 8646
rect 3809 8594 3811 8646
rect 3755 8592 3811 8594
rect 3879 8646 3935 8648
rect 3879 8594 3881 8646
rect 3881 8594 3933 8646
rect 3933 8594 3935 8646
rect 3879 8592 3935 8594
rect 3631 8522 3687 8524
rect 3631 8470 3633 8522
rect 3633 8470 3685 8522
rect 3685 8470 3687 8522
rect 3631 8468 3687 8470
rect 3755 8522 3811 8524
rect 3755 8470 3757 8522
rect 3757 8470 3809 8522
rect 3809 8470 3811 8522
rect 3755 8468 3811 8470
rect 3879 8522 3935 8524
rect 3879 8470 3881 8522
rect 3881 8470 3933 8522
rect 3933 8470 3935 8522
rect 3879 8468 3935 8470
rect 3631 8398 3687 8400
rect 3631 8346 3633 8398
rect 3633 8346 3685 8398
rect 3685 8346 3687 8398
rect 3631 8344 3687 8346
rect 3755 8398 3811 8400
rect 3755 8346 3757 8398
rect 3757 8346 3809 8398
rect 3809 8346 3811 8398
rect 3755 8344 3811 8346
rect 3879 8398 3935 8400
rect 3879 8346 3881 8398
rect 3881 8346 3933 8398
rect 3933 8346 3935 8398
rect 3879 8344 3935 8346
rect 3631 8274 3687 8276
rect 3631 8222 3633 8274
rect 3633 8222 3685 8274
rect 3685 8222 3687 8274
rect 3631 8220 3687 8222
rect 3755 8274 3811 8276
rect 3755 8222 3757 8274
rect 3757 8222 3809 8274
rect 3809 8222 3811 8274
rect 3755 8220 3811 8222
rect 3879 8274 3935 8276
rect 3879 8222 3881 8274
rect 3881 8222 3933 8274
rect 3933 8222 3935 8274
rect 3879 8220 3935 8222
rect 3631 8150 3687 8152
rect 3631 8098 3633 8150
rect 3633 8098 3685 8150
rect 3685 8098 3687 8150
rect 3631 8096 3687 8098
rect 3755 8150 3811 8152
rect 3755 8098 3757 8150
rect 3757 8098 3809 8150
rect 3809 8098 3811 8150
rect 3755 8096 3811 8098
rect 3879 8150 3935 8152
rect 3879 8098 3881 8150
rect 3881 8098 3933 8150
rect 3933 8098 3935 8150
rect 3879 8096 3935 8098
rect 3631 8026 3687 8028
rect 3631 7974 3633 8026
rect 3633 7974 3685 8026
rect 3685 7974 3687 8026
rect 3631 7972 3687 7974
rect 3755 8026 3811 8028
rect 3755 7974 3757 8026
rect 3757 7974 3809 8026
rect 3809 7974 3811 8026
rect 3755 7972 3811 7974
rect 3879 8026 3935 8028
rect 3879 7974 3881 8026
rect 3881 7974 3933 8026
rect 3933 7974 3935 8026
rect 3879 7972 3935 7974
rect 3631 7902 3687 7904
rect 3631 7850 3633 7902
rect 3633 7850 3685 7902
rect 3685 7850 3687 7902
rect 3631 7848 3687 7850
rect 3755 7902 3811 7904
rect 3755 7850 3757 7902
rect 3757 7850 3809 7902
rect 3809 7850 3811 7902
rect 3755 7848 3811 7850
rect 3879 7902 3935 7904
rect 3879 7850 3881 7902
rect 3881 7850 3933 7902
rect 3933 7850 3935 7902
rect 3879 7848 3935 7850
rect 3631 7778 3687 7780
rect 3631 7726 3633 7778
rect 3633 7726 3685 7778
rect 3685 7726 3687 7778
rect 3631 7724 3687 7726
rect 3755 7778 3811 7780
rect 3755 7726 3757 7778
rect 3757 7726 3809 7778
rect 3809 7726 3811 7778
rect 3755 7724 3811 7726
rect 3879 7778 3935 7780
rect 3879 7726 3881 7778
rect 3881 7726 3933 7778
rect 3933 7726 3935 7778
rect 3879 7724 3935 7726
rect 3631 7654 3687 7656
rect 3631 7602 3633 7654
rect 3633 7602 3685 7654
rect 3685 7602 3687 7654
rect 3631 7600 3687 7602
rect 3755 7654 3811 7656
rect 3755 7602 3757 7654
rect 3757 7602 3809 7654
rect 3809 7602 3811 7654
rect 3755 7600 3811 7602
rect 3879 7654 3935 7656
rect 3879 7602 3881 7654
rect 3881 7602 3933 7654
rect 3933 7602 3935 7654
rect 3879 7600 3935 7602
rect 4095 7379 4151 7435
rect 4219 7379 4275 7435
rect 4343 7379 4399 7435
rect 4467 7379 4523 7435
rect 4591 7379 4647 7435
rect 4715 7379 4771 7435
rect 4839 7379 4895 7435
rect 4963 7379 5019 7435
rect 4095 7255 4151 7311
rect 4219 7255 4275 7311
rect 4343 7255 4399 7311
rect 4467 7255 4523 7311
rect 4591 7255 4647 7311
rect 4715 7255 4771 7311
rect 4839 7255 4895 7311
rect 4963 7255 5019 7311
rect 4095 7131 4151 7187
rect 4219 7131 4275 7187
rect 4343 7131 4399 7187
rect 4467 7131 4523 7187
rect 4591 7131 4647 7187
rect 4715 7131 4771 7187
rect 4839 7131 4895 7187
rect 4963 7131 5019 7187
rect 4095 7007 4151 7063
rect 4219 7007 4275 7063
rect 4343 7007 4399 7063
rect 4467 7007 4523 7063
rect 4591 7007 4647 7063
rect 4715 7007 4771 7063
rect 4839 7007 4895 7063
rect 4963 7007 5019 7063
rect 4095 6883 4151 6939
rect 4219 6883 4275 6939
rect 4343 6883 4399 6939
rect 4467 6883 4523 6939
rect 4591 6883 4647 6939
rect 4715 6883 4771 6939
rect 4839 6883 4895 6939
rect 4963 6883 5019 6939
rect 4095 6759 4151 6815
rect 4219 6759 4275 6815
rect 4343 6759 4399 6815
rect 4467 6759 4523 6815
rect 4591 6759 4647 6815
rect 4715 6759 4771 6815
rect 4839 6759 4895 6815
rect 4963 6759 5019 6815
rect 4095 6635 4151 6691
rect 4219 6635 4275 6691
rect 4343 6635 4399 6691
rect 4467 6635 4523 6691
rect 4591 6635 4647 6691
rect 4715 6635 4771 6691
rect 4839 6635 4895 6691
rect 4963 6635 5019 6691
rect 4095 6511 4151 6567
rect 4219 6511 4275 6567
rect 4343 6511 4399 6567
rect 4467 6511 4523 6567
rect 4591 6511 4647 6567
rect 4715 6511 4771 6567
rect 4839 6511 4895 6567
rect 4963 6511 5019 6567
rect 4095 6387 4151 6443
rect 4219 6387 4275 6443
rect 4343 6387 4399 6443
rect 4467 6387 4523 6443
rect 4591 6387 4647 6443
rect 4715 6387 4771 6443
rect 4839 6387 4895 6443
rect 4963 6387 5019 6443
rect 4095 6263 4151 6319
rect 4219 6263 4275 6319
rect 4343 6263 4399 6319
rect 4467 6263 4523 6319
rect 4591 6263 4647 6319
rect 4715 6263 4771 6319
rect 4839 6263 4895 6319
rect 4963 6263 5019 6319
rect 4095 6139 4151 6195
rect 4219 6139 4275 6195
rect 4343 6139 4399 6195
rect 4467 6139 4523 6195
rect 4591 6139 4647 6195
rect 4715 6139 4771 6195
rect 4839 6139 4895 6195
rect 4963 6139 5019 6195
rect 4095 6015 4151 6071
rect 4219 6015 4275 6071
rect 4343 6015 4399 6071
rect 4467 6015 4523 6071
rect 4591 6015 4647 6071
rect 4715 6015 4771 6071
rect 4839 6015 4895 6071
rect 4963 6015 5019 6071
rect 4095 5891 4151 5947
rect 4219 5891 4275 5947
rect 4343 5891 4399 5947
rect 4467 5891 4523 5947
rect 4591 5891 4647 5947
rect 4715 5891 4771 5947
rect 4839 5891 4895 5947
rect 4963 5891 5019 5947
rect 3631 5526 3687 5528
rect 3631 5474 3633 5526
rect 3633 5474 3685 5526
rect 3685 5474 3687 5526
rect 3631 5472 3687 5474
rect 3755 5526 3811 5528
rect 3755 5474 3757 5526
rect 3757 5474 3809 5526
rect 3809 5474 3811 5526
rect 3755 5472 3811 5474
rect 3879 5526 3935 5528
rect 3879 5474 3881 5526
rect 3881 5474 3933 5526
rect 3933 5474 3935 5526
rect 3879 5472 3935 5474
rect 3631 5402 3687 5404
rect 3631 5350 3633 5402
rect 3633 5350 3685 5402
rect 3685 5350 3687 5402
rect 3631 5348 3687 5350
rect 3755 5402 3811 5404
rect 3755 5350 3757 5402
rect 3757 5350 3809 5402
rect 3809 5350 3811 5402
rect 3755 5348 3811 5350
rect 3879 5402 3935 5404
rect 3879 5350 3881 5402
rect 3881 5350 3933 5402
rect 3933 5350 3935 5402
rect 3879 5348 3935 5350
rect 3631 5278 3687 5280
rect 3631 5226 3633 5278
rect 3633 5226 3685 5278
rect 3685 5226 3687 5278
rect 3631 5224 3687 5226
rect 3755 5278 3811 5280
rect 3755 5226 3757 5278
rect 3757 5226 3809 5278
rect 3809 5226 3811 5278
rect 3755 5224 3811 5226
rect 3879 5278 3935 5280
rect 3879 5226 3881 5278
rect 3881 5226 3933 5278
rect 3933 5226 3935 5278
rect 3879 5224 3935 5226
rect 3631 5154 3687 5156
rect 3631 5102 3633 5154
rect 3633 5102 3685 5154
rect 3685 5102 3687 5154
rect 3631 5100 3687 5102
rect 3755 5154 3811 5156
rect 3755 5102 3757 5154
rect 3757 5102 3809 5154
rect 3809 5102 3811 5154
rect 3755 5100 3811 5102
rect 3879 5154 3935 5156
rect 3879 5102 3881 5154
rect 3881 5102 3933 5154
rect 3933 5102 3935 5154
rect 3879 5100 3935 5102
rect 3631 5030 3687 5032
rect 3631 4978 3633 5030
rect 3633 4978 3685 5030
rect 3685 4978 3687 5030
rect 3631 4976 3687 4978
rect 3755 5030 3811 5032
rect 3755 4978 3757 5030
rect 3757 4978 3809 5030
rect 3809 4978 3811 5030
rect 3755 4976 3811 4978
rect 3879 5030 3935 5032
rect 3879 4978 3881 5030
rect 3881 4978 3933 5030
rect 3933 4978 3935 5030
rect 3879 4976 3935 4978
rect 3631 4906 3687 4908
rect 3631 4854 3633 4906
rect 3633 4854 3685 4906
rect 3685 4854 3687 4906
rect 3631 4852 3687 4854
rect 3755 4906 3811 4908
rect 3755 4854 3757 4906
rect 3757 4854 3809 4906
rect 3809 4854 3811 4906
rect 3755 4852 3811 4854
rect 3879 4906 3935 4908
rect 3879 4854 3881 4906
rect 3881 4854 3933 4906
rect 3933 4854 3935 4906
rect 3879 4852 3935 4854
rect 3631 4782 3687 4784
rect 3631 4730 3633 4782
rect 3633 4730 3685 4782
rect 3685 4730 3687 4782
rect 3631 4728 3687 4730
rect 3755 4782 3811 4784
rect 3755 4730 3757 4782
rect 3757 4730 3809 4782
rect 3809 4730 3811 4782
rect 3755 4728 3811 4730
rect 3879 4782 3935 4784
rect 3879 4730 3881 4782
rect 3881 4730 3933 4782
rect 3933 4730 3935 4782
rect 3879 4728 3935 4730
rect 3631 4658 3687 4660
rect 3631 4606 3633 4658
rect 3633 4606 3685 4658
rect 3685 4606 3687 4658
rect 3631 4604 3687 4606
rect 3755 4658 3811 4660
rect 3755 4606 3757 4658
rect 3757 4606 3809 4658
rect 3809 4606 3811 4658
rect 3755 4604 3811 4606
rect 3879 4658 3935 4660
rect 3879 4606 3881 4658
rect 3881 4606 3933 4658
rect 3933 4606 3935 4658
rect 3879 4604 3935 4606
rect 3631 4534 3687 4536
rect 3631 4482 3633 4534
rect 3633 4482 3685 4534
rect 3685 4482 3687 4534
rect 3631 4480 3687 4482
rect 3755 4534 3811 4536
rect 3755 4482 3757 4534
rect 3757 4482 3809 4534
rect 3809 4482 3811 4534
rect 3755 4480 3811 4482
rect 3879 4534 3935 4536
rect 3879 4482 3881 4534
rect 3881 4482 3933 4534
rect 3933 4482 3935 4534
rect 3879 4480 3935 4482
rect 3631 4410 3687 4412
rect 3631 4358 3633 4410
rect 3633 4358 3685 4410
rect 3685 4358 3687 4410
rect 3631 4356 3687 4358
rect 3755 4410 3811 4412
rect 3755 4358 3757 4410
rect 3757 4358 3809 4410
rect 3809 4358 3811 4410
rect 3755 4356 3811 4358
rect 3879 4410 3935 4412
rect 3879 4358 3881 4410
rect 3881 4358 3933 4410
rect 3933 4358 3935 4410
rect 3879 4356 3935 4358
rect 4095 3954 4151 4010
rect 4219 3954 4275 4010
rect 4343 3954 4399 4010
rect 4467 3954 4523 4010
rect 4591 3954 4647 4010
rect 4715 3954 4771 4010
rect 4839 3954 4895 4010
rect 4963 3954 5019 4010
rect 4095 3830 4151 3886
rect 4219 3830 4275 3886
rect 4343 3830 4399 3886
rect 4467 3830 4523 3886
rect 4591 3830 4647 3886
rect 4715 3830 4771 3886
rect 4839 3830 4895 3886
rect 4963 3830 5019 3886
rect 4095 3706 4151 3762
rect 4219 3706 4275 3762
rect 4343 3706 4399 3762
rect 4467 3706 4523 3762
rect 4591 3706 4647 3762
rect 4715 3706 4771 3762
rect 4839 3706 4895 3762
rect 4963 3706 5019 3762
rect 4095 3582 4151 3638
rect 4219 3582 4275 3638
rect 4343 3582 4399 3638
rect 4467 3582 4523 3638
rect 4591 3582 4647 3638
rect 4715 3582 4771 3638
rect 4839 3582 4895 3638
rect 4963 3582 5019 3638
rect 4095 3458 4151 3514
rect 4219 3458 4275 3514
rect 4343 3458 4399 3514
rect 4467 3458 4523 3514
rect 4591 3458 4647 3514
rect 4715 3458 4771 3514
rect 4839 3458 4895 3514
rect 4963 3458 5019 3514
rect 4095 3334 4151 3390
rect 4219 3334 4275 3390
rect 4343 3334 4399 3390
rect 4467 3334 4523 3390
rect 4591 3334 4647 3390
rect 4715 3334 4771 3390
rect 4839 3334 4895 3390
rect 4963 3334 5019 3390
rect 4095 3210 4151 3266
rect 4219 3210 4275 3266
rect 4343 3210 4399 3266
rect 4467 3210 4523 3266
rect 4591 3210 4647 3266
rect 4715 3210 4771 3266
rect 4839 3210 4895 3266
rect 4963 3210 5019 3266
rect 4095 3086 4151 3142
rect 4219 3086 4275 3142
rect 4343 3086 4399 3142
rect 4467 3086 4523 3142
rect 4591 3086 4647 3142
rect 4715 3086 4771 3142
rect 4839 3086 4895 3142
rect 4963 3086 5019 3142
<< metal3 >>
rect 3339 37083 6351 37145
rect 3339 37027 3631 37083
rect 3687 37027 3755 37083
rect 3811 37027 3879 37083
rect 3935 37027 6351 37083
rect 3339 36959 6351 37027
rect 3339 36903 3631 36959
rect 3687 36903 3755 36959
rect 3811 36903 3879 36959
rect 3935 36945 6351 36959
rect 3935 36903 4353 36945
rect 3339 36835 4353 36903
rect 3339 36779 3631 36835
rect 3687 36779 3755 36835
rect 3811 36779 3879 36835
rect 3935 36779 6350 36835
rect 3339 36711 6350 36779
rect 3339 36655 3631 36711
rect 3687 36655 3755 36711
rect 3811 36655 3879 36711
rect 3935 36655 6350 36711
rect 3339 36587 6350 36655
rect 3339 36531 3631 36587
rect 3687 36531 3755 36587
rect 3811 36531 3879 36587
rect 3935 36531 6350 36587
rect 3339 36463 6350 36531
rect 3339 36407 3631 36463
rect 3687 36407 3755 36463
rect 3811 36407 3879 36463
rect 3935 36407 6350 36463
rect 3339 36355 6350 36407
rect 3339 35929 6350 35944
rect 3339 35873 4095 35929
rect 4151 35873 4219 35929
rect 4275 35873 4343 35929
rect 4399 35873 4467 35929
rect 4523 35873 4591 35929
rect 4647 35873 4715 35929
rect 4771 35873 4839 35929
rect 4895 35873 4963 35929
rect 5019 35873 6350 35929
rect 3339 35805 6350 35873
rect 3339 35749 4095 35805
rect 4151 35749 4219 35805
rect 4275 35749 4343 35805
rect 4399 35749 4467 35805
rect 4523 35749 4591 35805
rect 4647 35749 4715 35805
rect 4771 35749 4839 35805
rect 4895 35749 4963 35805
rect 5019 35749 6350 35805
rect 3339 35681 6350 35749
rect 3339 35625 4095 35681
rect 4151 35625 4219 35681
rect 4275 35625 4343 35681
rect 4399 35625 4467 35681
rect 4523 35625 4591 35681
rect 4647 35625 4715 35681
rect 4771 35625 4839 35681
rect 4895 35625 4963 35681
rect 5019 35625 6350 35681
rect 3339 35557 6350 35625
rect 3339 35501 4095 35557
rect 4151 35501 4219 35557
rect 4275 35501 4343 35557
rect 4399 35501 4467 35557
rect 4523 35501 4591 35557
rect 4647 35501 4715 35557
rect 4771 35501 4839 35557
rect 4895 35501 4963 35557
rect 5019 35501 6350 35557
rect 3339 35433 6350 35501
rect 3339 35377 4095 35433
rect 4151 35377 4219 35433
rect 4275 35377 4343 35433
rect 4399 35377 4467 35433
rect 4523 35377 4591 35433
rect 4647 35377 4715 35433
rect 4771 35377 4839 35433
rect 4895 35377 4963 35433
rect 5019 35377 6350 35433
rect 3339 35309 6350 35377
rect 3339 35253 4095 35309
rect 4151 35253 4219 35309
rect 4275 35253 4343 35309
rect 4399 35253 4467 35309
rect 4523 35253 4591 35309
rect 4647 35253 4715 35309
rect 4771 35253 4839 35309
rect 4895 35253 4963 35309
rect 5019 35253 6350 35309
rect 3339 35185 6350 35253
rect 3339 35129 4095 35185
rect 4151 35129 4219 35185
rect 4275 35129 4343 35185
rect 4399 35129 4467 35185
rect 4523 35129 4591 35185
rect 4647 35129 4715 35185
rect 4771 35129 4839 35185
rect 4895 35129 4963 35185
rect 5019 35129 6350 35185
rect 3339 35061 6350 35129
rect 3339 35005 4095 35061
rect 4151 35005 4219 35061
rect 4275 35005 4343 35061
rect 4399 35005 4467 35061
rect 4523 35005 4591 35061
rect 4647 35005 4715 35061
rect 4771 35005 4839 35061
rect 4895 35005 4963 35061
rect 5019 35005 6350 35061
rect 3339 34937 6350 35005
rect 3339 34881 4095 34937
rect 4151 34881 4219 34937
rect 4275 34881 4343 34937
rect 4399 34881 4467 34937
rect 4523 34881 4591 34937
rect 4647 34881 4715 34937
rect 4771 34881 4839 34937
rect 4895 34881 4963 34937
rect 5019 34881 6350 34937
rect 3339 34813 6350 34881
rect 3339 34757 4095 34813
rect 4151 34757 4219 34813
rect 4275 34757 4343 34813
rect 4399 34757 4467 34813
rect 4523 34757 4591 34813
rect 4647 34757 4715 34813
rect 4771 34757 4839 34813
rect 4895 34757 4963 34813
rect 5019 34757 6350 34813
rect 3339 34689 6350 34757
rect 3339 34633 4095 34689
rect 4151 34633 4219 34689
rect 4275 34633 4343 34689
rect 4399 34633 4467 34689
rect 4523 34633 4591 34689
rect 4647 34633 4715 34689
rect 4771 34633 4839 34689
rect 4895 34633 4963 34689
rect 5019 34633 6350 34689
rect 3339 34565 6350 34633
rect 3339 34509 4095 34565
rect 4151 34509 4219 34565
rect 4275 34509 4343 34565
rect 4399 34509 4467 34565
rect 4523 34509 4591 34565
rect 4647 34509 4715 34565
rect 4771 34509 4839 34565
rect 4895 34509 4963 34565
rect 5019 34509 6350 34565
rect 3339 34441 6350 34509
rect 3339 34385 4095 34441
rect 4151 34385 4219 34441
rect 4275 34385 4343 34441
rect 4399 34385 4467 34441
rect 4523 34385 4591 34441
rect 4647 34385 4715 34441
rect 4771 34385 4839 34441
rect 4895 34385 4963 34441
rect 5019 34385 6350 34441
rect 3339 34317 6350 34385
rect 3339 34261 4095 34317
rect 4151 34261 4219 34317
rect 4275 34261 4343 34317
rect 4399 34261 4467 34317
rect 4523 34261 4591 34317
rect 4647 34261 4715 34317
rect 4771 34261 4839 34317
rect 4895 34261 4963 34317
rect 5019 34261 6350 34317
rect 3339 34193 6350 34261
rect 3339 34137 4095 34193
rect 4151 34137 4219 34193
rect 4275 34137 4343 34193
rect 4399 34137 4467 34193
rect 4523 34137 4591 34193
rect 4647 34137 4715 34193
rect 4771 34137 4839 34193
rect 4895 34137 4963 34193
rect 5019 34137 6350 34193
rect 3339 34134 6350 34137
rect 3339 34069 5045 34134
rect 3339 34013 4095 34069
rect 4151 34013 4219 34069
rect 4275 34013 4343 34069
rect 4399 34013 4467 34069
rect 4523 34013 4591 34069
rect 4647 34013 4715 34069
rect 4771 34013 4839 34069
rect 4895 34013 4963 34069
rect 5019 34013 5045 34069
rect 3339 33945 5045 34013
rect 3339 33889 4095 33945
rect 4151 33889 4219 33945
rect 4275 33889 4343 33945
rect 4399 33889 4467 33945
rect 4523 33889 4591 33945
rect 4647 33889 4715 33945
rect 4771 33889 4839 33945
rect 4895 33889 4963 33945
rect 5019 33889 5045 33945
rect 3339 33821 5045 33889
rect 3339 33765 4095 33821
rect 4151 33765 4219 33821
rect 4275 33765 4343 33821
rect 4399 33765 4467 33821
rect 4523 33765 4591 33821
rect 4647 33765 4715 33821
rect 4771 33765 4839 33821
rect 4895 33765 4963 33821
rect 5019 33765 5045 33821
rect 3339 33697 5045 33765
rect 3339 33641 4095 33697
rect 4151 33641 4219 33697
rect 4275 33641 4343 33697
rect 4399 33641 4467 33697
rect 4523 33641 4591 33697
rect 4647 33641 4715 33697
rect 4771 33641 4839 33697
rect 4895 33641 4963 33697
rect 5019 33641 5045 33697
rect 3339 33573 5045 33641
rect 3339 33517 4095 33573
rect 4151 33517 4219 33573
rect 4275 33517 4343 33573
rect 4399 33517 4467 33573
rect 4523 33517 4591 33573
rect 4647 33517 4715 33573
rect 4771 33517 4839 33573
rect 4895 33517 4963 33573
rect 5019 33517 5045 33573
rect 3339 33449 5045 33517
rect 3339 33393 4095 33449
rect 4151 33393 4219 33449
rect 4275 33393 4343 33449
rect 4399 33393 4467 33449
rect 4523 33393 4591 33449
rect 4647 33393 4715 33449
rect 4771 33393 4839 33449
rect 4895 33393 4963 33449
rect 5019 33393 5045 33449
rect 3339 33325 5045 33393
rect 3339 33269 4095 33325
rect 4151 33269 4219 33325
rect 4275 33269 4343 33325
rect 4399 33269 4467 33325
rect 4523 33269 4591 33325
rect 4647 33269 4715 33325
rect 4771 33269 4839 33325
rect 4895 33269 4963 33325
rect 5019 33269 5045 33325
rect 3339 33201 5045 33269
rect 3339 33145 4095 33201
rect 4151 33145 4219 33201
rect 4275 33145 4343 33201
rect 4399 33145 4467 33201
rect 4523 33145 4591 33201
rect 4647 33145 4715 33201
rect 4771 33145 4839 33201
rect 4895 33145 4963 33201
rect 5019 33145 5045 33201
rect 3339 33077 5045 33145
rect 3339 33021 4095 33077
rect 4151 33021 4219 33077
rect 4275 33021 4343 33077
rect 4399 33021 4467 33077
rect 4523 33021 4591 33077
rect 4647 33021 4715 33077
rect 4771 33021 4839 33077
rect 4895 33021 4963 33077
rect 5019 33021 5045 33077
rect 3339 32953 5045 33021
rect 3339 32897 4095 32953
rect 4151 32897 4219 32953
rect 4275 32897 4343 32953
rect 4399 32897 4467 32953
rect 4523 32897 4591 32953
rect 4647 32897 4715 32953
rect 4771 32897 4839 32953
rect 4895 32897 4963 32953
rect 5019 32897 5045 32953
rect 3339 32829 5045 32897
rect 3339 32773 4095 32829
rect 4151 32773 4219 32829
rect 4275 32773 4343 32829
rect 4399 32773 4467 32829
rect 4523 32773 4591 32829
rect 4647 32773 4715 32829
rect 4771 32773 4839 32829
rect 4895 32773 4963 32829
rect 5019 32773 5045 32829
rect 3339 32705 5045 32773
rect 3339 32649 4095 32705
rect 4151 32649 4219 32705
rect 4275 32649 4343 32705
rect 4399 32649 4467 32705
rect 4523 32649 4591 32705
rect 4647 32649 4715 32705
rect 4771 32649 4839 32705
rect 4895 32649 4963 32705
rect 5019 32649 5045 32705
rect 3339 32581 5045 32649
rect 3339 32525 4095 32581
rect 4151 32525 4219 32581
rect 4275 32525 4343 32581
rect 4399 32525 4467 32581
rect 4523 32525 4591 32581
rect 4647 32525 4715 32581
rect 4771 32525 4839 32581
rect 4895 32525 4963 32581
rect 5019 32525 5045 32581
rect 3339 32457 5045 32525
rect 3339 32401 4095 32457
rect 4151 32401 4219 32457
rect 4275 32401 4343 32457
rect 4399 32401 4467 32457
rect 4523 32401 4591 32457
rect 4647 32401 4715 32457
rect 4771 32401 4839 32457
rect 4895 32401 4963 32457
rect 5019 32401 5045 32457
rect 3339 32333 5045 32401
rect 3339 32277 4095 32333
rect 4151 32277 4219 32333
rect 4275 32277 4343 32333
rect 4399 32277 4467 32333
rect 4523 32277 4591 32333
rect 4647 32277 4715 32333
rect 4771 32277 4839 32333
rect 4895 32277 4963 32333
rect 5019 32277 5045 32333
rect 3339 32209 5045 32277
rect 3339 32153 4095 32209
rect 4151 32153 4219 32209
rect 4275 32153 4343 32209
rect 4399 32153 4467 32209
rect 4523 32153 4591 32209
rect 4647 32153 4715 32209
rect 4771 32153 4839 32209
rect 4895 32153 4963 32209
rect 5019 32153 5045 32209
rect 3339 32085 5045 32153
rect 3339 32029 4095 32085
rect 4151 32029 4219 32085
rect 4275 32029 4343 32085
rect 4399 32029 4467 32085
rect 4523 32029 4591 32085
rect 4647 32029 4715 32085
rect 4771 32029 4839 32085
rect 4895 32029 4963 32085
rect 5019 32029 5045 32085
rect 3339 31961 5045 32029
rect 3339 31905 4095 31961
rect 4151 31905 4219 31961
rect 4275 31905 4343 31961
rect 4399 31905 4467 31961
rect 4523 31905 4591 31961
rect 4647 31905 4715 31961
rect 4771 31905 4839 31961
rect 4895 31905 4963 31961
rect 5019 31905 5045 31961
rect 3339 31837 5045 31905
rect 3339 31781 4095 31837
rect 4151 31781 4219 31837
rect 4275 31781 4343 31837
rect 4399 31781 4467 31837
rect 4523 31781 4591 31837
rect 4647 31781 4715 31837
rect 4771 31781 4839 31837
rect 4895 31781 4963 31837
rect 5019 31781 5045 31837
rect 3339 31713 5045 31781
rect 3339 31657 4095 31713
rect 4151 31657 4219 31713
rect 4275 31657 4343 31713
rect 4399 31657 4467 31713
rect 4523 31657 4591 31713
rect 4647 31657 4715 31713
rect 4771 31657 4839 31713
rect 4895 31657 4963 31713
rect 5019 31657 5045 31713
rect 3339 31589 5045 31657
rect 3339 31533 4095 31589
rect 4151 31533 4219 31589
rect 4275 31533 4343 31589
rect 4399 31533 4467 31589
rect 4523 31533 4591 31589
rect 4647 31533 4715 31589
rect 4771 31533 4839 31589
rect 4895 31533 4963 31589
rect 5019 31533 5045 31589
rect 3339 31465 6632 31533
rect 3339 31409 4095 31465
rect 4151 31409 4219 31465
rect 4275 31409 4343 31465
rect 4399 31409 4467 31465
rect 4523 31409 4591 31465
rect 4647 31409 4715 31465
rect 4771 31409 4839 31465
rect 4895 31409 4963 31465
rect 5019 31409 6632 31465
rect 3339 31341 6632 31409
rect 3339 31285 4095 31341
rect 4151 31285 4219 31341
rect 4275 31285 4343 31341
rect 4399 31285 4467 31341
rect 4523 31285 4591 31341
rect 4647 31285 4715 31341
rect 4771 31285 4839 31341
rect 4895 31285 4963 31341
rect 5019 31285 6632 31341
rect 3339 31249 6632 31285
rect 3339 30159 6350 30235
rect 3339 30103 3631 30159
rect 3687 30103 3755 30159
rect 3811 30103 3879 30159
rect 3935 30103 6350 30159
rect 3339 30035 6350 30103
rect 3339 29979 3631 30035
rect 3687 29979 3755 30035
rect 3811 29979 3879 30035
rect 3935 29979 6350 30035
rect 3339 29911 6350 29979
rect 3339 29855 3631 29911
rect 3687 29855 3755 29911
rect 3811 29855 3879 29911
rect 3935 29855 6350 29911
rect 3339 29787 6350 29855
rect 3339 29731 3631 29787
rect 3687 29731 3755 29787
rect 3811 29731 3879 29787
rect 3935 29731 6350 29787
rect 3339 29663 6350 29731
rect 3339 29607 3631 29663
rect 3687 29607 3755 29663
rect 3811 29607 3879 29663
rect 3935 29607 6350 29663
rect 3339 29539 6350 29607
rect 3339 29483 3631 29539
rect 3687 29483 3755 29539
rect 3811 29483 3879 29539
rect 3935 29483 6350 29539
rect 3339 29415 6350 29483
rect 3339 29359 3631 29415
rect 3687 29359 3755 29415
rect 3811 29359 3879 29415
rect 3935 29359 6350 29415
rect 3339 29291 6350 29359
rect 3339 29235 3631 29291
rect 3687 29235 3755 29291
rect 3811 29235 3879 29291
rect 3935 29235 6350 29291
rect 3339 29167 6350 29235
rect 3339 29111 3631 29167
rect 3687 29111 3755 29167
rect 3811 29111 3879 29167
rect 3935 29111 6350 29167
rect 3339 29043 6350 29111
rect 3339 28987 3631 29043
rect 3687 28987 3755 29043
rect 3811 28987 3879 29043
rect 3935 28987 6350 29043
rect 3339 28919 6350 28987
rect 3339 28863 3631 28919
rect 3687 28863 3755 28919
rect 3811 28863 3879 28919
rect 3935 28863 6350 28919
rect 3339 28795 6350 28863
rect 3339 28739 3631 28795
rect 3687 28739 3755 28795
rect 3811 28739 3879 28795
rect 3935 28739 6350 28795
rect 3339 28671 6350 28739
rect 3339 28615 3631 28671
rect 3687 28615 3755 28671
rect 3811 28615 3879 28671
rect 3935 28615 6350 28671
rect 3339 28547 6350 28615
rect 3339 28491 3631 28547
rect 3687 28491 3755 28547
rect 3811 28491 3879 28547
rect 3935 28491 6350 28547
rect 3339 28423 6350 28491
rect 3339 28367 3631 28423
rect 3687 28367 3755 28423
rect 3811 28367 3879 28423
rect 3935 28367 6350 28423
rect 3339 28254 6350 28367
rect 3339 25691 5045 25757
rect 3339 25635 4095 25691
rect 4151 25635 4219 25691
rect 4275 25635 4343 25691
rect 4399 25635 4467 25691
rect 4523 25635 4591 25691
rect 4647 25635 4715 25691
rect 4771 25635 4839 25691
rect 4895 25635 4963 25691
rect 5019 25635 5045 25691
rect 3339 25567 5045 25635
rect 3339 25511 4095 25567
rect 4151 25511 4219 25567
rect 4275 25511 4343 25567
rect 4399 25511 4467 25567
rect 4523 25511 4591 25567
rect 4647 25511 4715 25567
rect 4771 25511 4839 25567
rect 4895 25511 4963 25567
rect 5019 25511 5045 25567
rect 3339 25443 5045 25511
rect 3339 25387 4095 25443
rect 4151 25387 4219 25443
rect 4275 25387 4343 25443
rect 4399 25387 4467 25443
rect 4523 25387 4591 25443
rect 4647 25387 4715 25443
rect 4771 25387 4839 25443
rect 4895 25387 4963 25443
rect 5019 25387 5045 25443
rect 3339 25319 5045 25387
rect 3339 25263 4095 25319
rect 4151 25263 4219 25319
rect 4275 25263 4343 25319
rect 4399 25263 4467 25319
rect 4523 25263 4591 25319
rect 4647 25263 4715 25319
rect 4771 25263 4839 25319
rect 4895 25263 4963 25319
rect 5019 25263 5045 25319
rect 3339 25199 5045 25263
rect 3339 25195 6350 25199
rect 3339 25139 4095 25195
rect 4151 25139 4219 25195
rect 4275 25139 4343 25195
rect 4399 25139 4467 25195
rect 4523 25139 4591 25195
rect 4647 25139 4715 25195
rect 4771 25139 4839 25195
rect 4895 25139 4963 25195
rect 5019 25139 6350 25195
rect 3339 25071 6350 25139
rect 3339 25015 4095 25071
rect 4151 25015 4219 25071
rect 4275 25015 4343 25071
rect 4399 25015 4467 25071
rect 4523 25015 4591 25071
rect 4647 25015 4715 25071
rect 4771 25015 4839 25071
rect 4895 25015 4963 25071
rect 5019 25015 6350 25071
rect 3339 24947 6350 25015
rect 3339 24891 4095 24947
rect 4151 24891 4219 24947
rect 4275 24891 4343 24947
rect 4399 24891 4467 24947
rect 4523 24891 4591 24947
rect 4647 24891 4715 24947
rect 4771 24891 4839 24947
rect 4895 24891 4963 24947
rect 5019 24891 6350 24947
rect 3339 24823 6350 24891
rect 3339 24767 4095 24823
rect 4151 24767 4219 24823
rect 4275 24767 4343 24823
rect 4399 24767 4467 24823
rect 4523 24767 4591 24823
rect 4647 24767 4715 24823
rect 4771 24767 4839 24823
rect 4895 24767 4963 24823
rect 5019 24767 6350 24823
rect 3339 24757 6350 24767
rect 3339 24064 6350 24101
rect 3339 24008 3631 24064
rect 3687 24008 3755 24064
rect 3811 24008 3879 24064
rect 3935 24008 6350 24064
rect 3339 23940 6350 24008
rect 3339 23884 3631 23940
rect 3687 23884 3755 23940
rect 3811 23884 3879 23940
rect 3935 23884 6350 23940
rect 3339 23816 6350 23884
rect 3339 23760 3631 23816
rect 3687 23760 3755 23816
rect 3811 23760 3879 23816
rect 3935 23760 6350 23816
rect 3339 23692 6350 23760
rect 3339 23636 3631 23692
rect 3687 23636 3755 23692
rect 3811 23636 3879 23692
rect 3935 23646 6350 23692
rect 3935 23636 4353 23646
rect 3339 23568 4353 23636
rect 3339 23512 3631 23568
rect 3687 23512 3755 23568
rect 3811 23512 3879 23568
rect 3935 23512 4353 23568
rect 3339 23444 4353 23512
rect 3339 23388 3631 23444
rect 3687 23388 3755 23444
rect 3811 23388 3879 23444
rect 3935 23388 4353 23444
rect 3339 23320 4353 23388
rect 3339 23264 3631 23320
rect 3687 23264 3755 23320
rect 3811 23264 3879 23320
rect 3935 23264 4353 23320
rect 3339 23196 4353 23264
rect 3339 23140 3631 23196
rect 3687 23140 3755 23196
rect 3811 23140 3879 23196
rect 3935 23140 4353 23196
rect 3339 23101 4353 23140
rect 3339 22512 6350 22558
rect 3339 22456 4095 22512
rect 4151 22456 4219 22512
rect 4275 22456 4343 22512
rect 4399 22456 4467 22512
rect 4523 22456 4591 22512
rect 4647 22456 4715 22512
rect 4771 22456 4839 22512
rect 4895 22456 4963 22512
rect 5019 22456 6350 22512
rect 3339 22388 6350 22456
rect 3339 22332 4095 22388
rect 4151 22332 4219 22388
rect 4275 22332 4343 22388
rect 4399 22332 4467 22388
rect 4523 22332 4591 22388
rect 4647 22332 4715 22388
rect 4771 22332 4839 22388
rect 4895 22332 4963 22388
rect 5019 22332 6350 22388
rect 3339 22264 6350 22332
rect 3339 22208 4095 22264
rect 4151 22208 4219 22264
rect 4275 22208 4343 22264
rect 4399 22208 4467 22264
rect 4523 22208 4591 22264
rect 4647 22208 4715 22264
rect 4771 22208 4839 22264
rect 4895 22208 4963 22264
rect 5019 22208 6350 22264
rect 3339 22140 6350 22208
rect 3339 22084 4095 22140
rect 4151 22084 4219 22140
rect 4275 22084 4343 22140
rect 4399 22084 4467 22140
rect 4523 22084 4591 22140
rect 4647 22084 4715 22140
rect 4771 22084 4839 22140
rect 4895 22084 4963 22140
rect 5019 22084 6350 22140
rect 3339 22016 6350 22084
rect 3339 21960 4095 22016
rect 4151 21960 4219 22016
rect 4275 21960 4343 22016
rect 4399 21960 4467 22016
rect 4523 21960 4591 22016
rect 4647 21960 4715 22016
rect 4771 21960 4839 22016
rect 4895 21960 4963 22016
rect 5019 21960 6350 22016
rect 3339 21892 6350 21960
rect 3339 21836 4095 21892
rect 4151 21836 4219 21892
rect 4275 21836 4343 21892
rect 4399 21836 4467 21892
rect 4523 21836 4591 21892
rect 4647 21836 4715 21892
rect 4771 21836 4839 21892
rect 4895 21836 4963 21892
rect 5019 21836 6350 21892
rect 3339 21768 6350 21836
rect 3339 21712 4095 21768
rect 4151 21712 4219 21768
rect 4275 21712 4343 21768
rect 4399 21712 4467 21768
rect 4523 21712 4591 21768
rect 4647 21712 4715 21768
rect 4771 21712 4839 21768
rect 4895 21712 4963 21768
rect 5019 21712 6350 21768
rect 3339 21644 6350 21712
rect 3339 21588 4095 21644
rect 4151 21588 4219 21644
rect 4275 21588 4343 21644
rect 4399 21588 4467 21644
rect 4523 21588 4591 21644
rect 4647 21588 4715 21644
rect 4771 21588 4839 21644
rect 4895 21588 4963 21644
rect 5019 21588 6350 21644
rect 3339 21520 6350 21588
rect 3339 21464 4095 21520
rect 4151 21464 4219 21520
rect 4275 21464 4343 21520
rect 4399 21464 4467 21520
rect 4523 21464 4591 21520
rect 4647 21464 4715 21520
rect 4771 21464 4839 21520
rect 4895 21464 4963 21520
rect 5019 21464 6350 21520
rect 3339 21396 6350 21464
rect 3339 21340 4095 21396
rect 4151 21340 4219 21396
rect 4275 21340 4343 21396
rect 4399 21340 4467 21396
rect 4523 21340 4591 21396
rect 4647 21340 4715 21396
rect 4771 21340 4839 21396
rect 4895 21340 4963 21396
rect 5019 21340 6350 21396
rect 3339 21272 6350 21340
rect 3339 21216 4095 21272
rect 4151 21216 4219 21272
rect 4275 21216 4343 21272
rect 4399 21216 4467 21272
rect 4523 21216 4591 21272
rect 4647 21216 4715 21272
rect 4771 21216 4839 21272
rect 4895 21216 4963 21272
rect 5019 21216 6350 21272
rect 3339 21148 6350 21216
rect 3339 21092 4095 21148
rect 4151 21092 4219 21148
rect 4275 21092 4343 21148
rect 4399 21092 4467 21148
rect 4523 21092 4591 21148
rect 4647 21092 4715 21148
rect 4771 21092 4839 21148
rect 4895 21092 4963 21148
rect 5019 21092 6350 21148
rect 3339 21024 6350 21092
rect 3339 20968 4095 21024
rect 4151 20968 4219 21024
rect 4275 20968 4343 21024
rect 4399 20968 4467 21024
rect 4523 20968 4591 21024
rect 4647 20968 4715 21024
rect 4771 20968 4839 21024
rect 4895 20968 4963 21024
rect 5019 20968 6350 21024
rect 3339 20900 6350 20968
rect 3339 20844 4095 20900
rect 4151 20844 4219 20900
rect 4275 20844 4343 20900
rect 4399 20844 4467 20900
rect 4523 20844 4591 20900
rect 4647 20844 4715 20900
rect 4771 20844 4839 20900
rect 4895 20844 4963 20900
rect 5019 20844 6350 20900
rect 3339 20776 6350 20844
rect 3339 20720 4095 20776
rect 4151 20720 4219 20776
rect 4275 20720 4343 20776
rect 4399 20720 4467 20776
rect 4523 20720 4591 20776
rect 4647 20720 4715 20776
rect 4771 20720 4839 20776
rect 4895 20720 4963 20776
rect 5019 20720 6350 20776
rect 3339 20652 6350 20720
rect 3339 20596 4095 20652
rect 4151 20596 4219 20652
rect 4275 20596 4343 20652
rect 4399 20596 4467 20652
rect 4523 20596 4591 20652
rect 4647 20596 4715 20652
rect 4771 20596 4839 20652
rect 4895 20596 4963 20652
rect 5019 20596 6350 20652
rect 3339 20528 6350 20596
rect 3339 20472 4095 20528
rect 4151 20472 4219 20528
rect 4275 20472 4343 20528
rect 4399 20472 4467 20528
rect 4523 20472 4591 20528
rect 4647 20472 4715 20528
rect 4771 20472 4839 20528
rect 4895 20472 4963 20528
rect 5019 20472 6350 20528
rect 3339 20404 6350 20472
rect 3339 20348 4095 20404
rect 4151 20348 4219 20404
rect 4275 20348 4343 20404
rect 4399 20348 4467 20404
rect 4523 20348 4591 20404
rect 4647 20348 4715 20404
rect 4771 20348 4839 20404
rect 4895 20348 4963 20404
rect 5019 20348 6350 20404
rect 3339 20280 6350 20348
rect 3339 20224 4095 20280
rect 4151 20224 4219 20280
rect 4275 20224 4343 20280
rect 4399 20224 4467 20280
rect 4523 20224 4591 20280
rect 4647 20224 4715 20280
rect 4771 20224 4839 20280
rect 4895 20224 4963 20280
rect 5019 20224 6350 20280
rect 3339 20156 6350 20224
rect 3339 20100 4095 20156
rect 4151 20100 4219 20156
rect 4275 20100 4343 20156
rect 4399 20100 4467 20156
rect 4523 20100 4591 20156
rect 4647 20100 4715 20156
rect 4771 20100 4839 20156
rect 4895 20100 4963 20156
rect 5019 20100 6350 20156
rect 3339 20032 6350 20100
rect 3339 19976 4095 20032
rect 4151 19976 4219 20032
rect 4275 19976 4343 20032
rect 4399 19976 4467 20032
rect 4523 19976 4591 20032
rect 4647 19976 4715 20032
rect 4771 19976 4839 20032
rect 4895 19976 4963 20032
rect 5019 19976 6350 20032
rect 3339 19908 6350 19976
rect 3339 19852 4095 19908
rect 4151 19852 4219 19908
rect 4275 19852 4343 19908
rect 4399 19852 4467 19908
rect 4523 19852 4591 19908
rect 4647 19852 4715 19908
rect 4771 19852 4839 19908
rect 4895 19852 4963 19908
rect 5019 19852 6350 19908
rect 3339 19835 6350 19852
rect 3339 19507 6350 19549
rect 3339 19451 3631 19507
rect 3687 19451 3755 19507
rect 3811 19451 3879 19507
rect 3935 19451 6350 19507
rect 3339 19383 6350 19451
rect 3339 19327 3631 19383
rect 3687 19327 3755 19383
rect 3811 19327 3879 19383
rect 3935 19327 6350 19383
rect 3339 19259 6350 19327
rect 3339 19203 3631 19259
rect 3687 19203 3755 19259
rect 3811 19203 3879 19259
rect 3935 19203 6350 19259
rect 3339 19135 6350 19203
rect 3339 19079 3631 19135
rect 3687 19079 3755 19135
rect 3811 19079 3879 19135
rect 3935 19079 6350 19135
rect 3339 19011 6350 19079
rect 3339 18955 3631 19011
rect 3687 18955 3755 19011
rect 3811 18955 3879 19011
rect 3935 18955 6350 19011
rect 3339 18887 6350 18955
rect 3339 18831 3631 18887
rect 3687 18831 3755 18887
rect 3811 18831 3879 18887
rect 3935 18831 6350 18887
rect 3339 18763 6350 18831
rect 3339 18707 3631 18763
rect 3687 18707 3755 18763
rect 3811 18707 3879 18763
rect 3935 18707 6350 18763
rect 3339 18639 6350 18707
rect 3339 18583 3631 18639
rect 3687 18583 3755 18639
rect 3811 18583 3879 18639
rect 3935 18583 6350 18639
rect 3339 18515 6350 18583
rect 3339 18459 3631 18515
rect 3687 18459 3755 18515
rect 3811 18459 3879 18515
rect 3935 18459 6350 18515
rect 3339 18391 6350 18459
rect 3339 18335 3631 18391
rect 3687 18335 3755 18391
rect 3811 18335 3879 18391
rect 3935 18335 6350 18391
rect 3339 18267 6350 18335
rect 3339 18211 3631 18267
rect 3687 18211 3755 18267
rect 3811 18211 3879 18267
rect 3935 18211 6350 18267
rect 3339 18143 6350 18211
rect 3339 18087 3631 18143
rect 3687 18087 3755 18143
rect 3811 18087 3879 18143
rect 3935 18087 6350 18143
rect 3339 18019 6350 18087
rect 3339 17963 3631 18019
rect 3687 17963 3755 18019
rect 3811 17963 3879 18019
rect 3935 17963 6350 18019
rect 3339 17895 6350 17963
rect 3339 17839 3631 17895
rect 3687 17839 3755 17895
rect 3811 17839 3879 17895
rect 3935 17839 6350 17895
rect 3339 17771 6350 17839
rect 3339 17715 3631 17771
rect 3687 17715 3755 17771
rect 3811 17715 3879 17771
rect 3935 17715 6350 17771
rect 3339 17647 6350 17715
rect 3339 17591 3631 17647
rect 3687 17591 3755 17647
rect 3811 17591 3879 17647
rect 3935 17591 6350 17647
rect 3339 17523 6350 17591
rect 3339 17467 3631 17523
rect 3687 17467 3755 17523
rect 3811 17467 3879 17523
rect 3935 17467 6350 17523
rect 3339 17399 6350 17467
rect 3339 17343 3631 17399
rect 3687 17343 3755 17399
rect 3811 17343 3879 17399
rect 3935 17343 6350 17399
rect 3339 17275 6350 17343
rect 3339 17219 3631 17275
rect 3687 17219 3755 17275
rect 3811 17219 3879 17275
rect 3935 17219 6350 17275
rect 3339 17151 6350 17219
rect 3339 17095 3631 17151
rect 3687 17095 3755 17151
rect 3811 17095 3879 17151
rect 3935 17095 6350 17151
rect 3339 17027 6350 17095
rect 3339 16971 3631 17027
rect 3687 16971 3755 17027
rect 3811 16971 3879 17027
rect 3935 16971 6350 17027
rect 3339 16903 6350 16971
rect 3339 16847 3631 16903
rect 3687 16847 3755 16903
rect 3811 16847 3879 16903
rect 3935 16847 6350 16903
rect 3339 16779 6350 16847
rect 3339 16723 3631 16779
rect 3687 16723 3755 16779
rect 3811 16723 3879 16779
rect 3935 16723 6350 16779
rect 3339 16655 6350 16723
rect 3339 16599 3631 16655
rect 3687 16599 3755 16655
rect 3811 16599 3879 16655
rect 3935 16599 6350 16655
rect 3339 16531 6350 16599
rect 3339 16475 3631 16531
rect 3687 16475 3755 16531
rect 3811 16475 3879 16531
rect 3935 16475 6350 16531
rect 3339 16407 6350 16475
rect 3339 16351 3631 16407
rect 3687 16351 3755 16407
rect 3811 16351 3879 16407
rect 3935 16351 6350 16407
rect 3339 16283 6350 16351
rect 3339 16227 3631 16283
rect 3687 16227 3755 16283
rect 3811 16227 3879 16283
rect 3935 16227 6350 16283
rect 3339 16147 6350 16227
rect 3339 15942 6350 15997
rect 3339 15886 4095 15942
rect 4151 15886 4219 15942
rect 4275 15886 4343 15942
rect 4399 15886 4467 15942
rect 4523 15886 4591 15942
rect 4647 15886 4715 15942
rect 4771 15886 4839 15942
rect 4895 15886 4963 15942
rect 5019 15886 6350 15942
rect 3339 15818 6350 15886
rect 3339 15762 4095 15818
rect 4151 15762 4219 15818
rect 4275 15762 4343 15818
rect 4399 15762 4467 15818
rect 4523 15762 4591 15818
rect 4647 15762 4715 15818
rect 4771 15762 4839 15818
rect 4895 15762 4963 15818
rect 5019 15762 6350 15818
rect 3339 15694 6350 15762
rect 3339 15638 4095 15694
rect 4151 15638 4219 15694
rect 4275 15638 4343 15694
rect 4399 15638 4467 15694
rect 4523 15638 4591 15694
rect 4647 15638 4715 15694
rect 4771 15638 4839 15694
rect 4895 15638 4963 15694
rect 5019 15638 6350 15694
rect 3339 15570 6350 15638
rect 3339 15514 4095 15570
rect 4151 15514 4219 15570
rect 4275 15514 4343 15570
rect 4399 15514 4467 15570
rect 4523 15514 4591 15570
rect 4647 15514 4715 15570
rect 4771 15514 4839 15570
rect 4895 15514 4963 15570
rect 5019 15514 6350 15570
rect 3339 15446 6350 15514
rect 3339 15390 4095 15446
rect 4151 15390 4219 15446
rect 4275 15390 4343 15446
rect 4399 15390 4467 15446
rect 4523 15390 4591 15446
rect 4647 15390 4715 15446
rect 4771 15390 4839 15446
rect 4895 15390 4963 15446
rect 5019 15390 6350 15446
rect 3339 15322 6350 15390
rect 3339 15266 4095 15322
rect 4151 15266 4219 15322
rect 4275 15266 4343 15322
rect 4399 15266 4467 15322
rect 4523 15266 4591 15322
rect 4647 15266 4715 15322
rect 4771 15266 4839 15322
rect 4895 15266 4963 15322
rect 5019 15280 6350 15322
rect 5019 15266 5045 15280
rect 3339 15198 5045 15266
rect 3339 15142 4095 15198
rect 4151 15142 4219 15198
rect 4275 15142 4343 15198
rect 4399 15142 4467 15198
rect 4523 15142 4591 15198
rect 4647 15142 4715 15198
rect 4771 15142 4839 15198
rect 4895 15142 4963 15198
rect 5019 15142 5045 15198
rect 3339 15074 5045 15142
rect 3339 15018 4095 15074
rect 4151 15018 4219 15074
rect 4275 15018 4343 15074
rect 4399 15018 4467 15074
rect 4523 15018 4591 15074
rect 4647 15018 4715 15074
rect 4771 15018 4839 15074
rect 4895 15018 4963 15074
rect 5019 15018 5045 15074
rect 3339 14950 5045 15018
rect 3339 14894 4095 14950
rect 4151 14894 4219 14950
rect 4275 14894 4343 14950
rect 4399 14894 4467 14950
rect 4523 14894 4591 14950
rect 4647 14894 4715 14950
rect 4771 14894 4839 14950
rect 4895 14894 4963 14950
rect 5019 14894 5045 14950
rect 3339 14826 5045 14894
rect 3339 14770 4095 14826
rect 4151 14770 4219 14826
rect 4275 14770 4343 14826
rect 4399 14770 4467 14826
rect 4523 14770 4591 14826
rect 4647 14770 4715 14826
rect 4771 14770 4839 14826
rect 4895 14770 4963 14826
rect 5019 14770 5045 14826
rect 3339 14702 5045 14770
rect 3339 14646 4095 14702
rect 4151 14646 4219 14702
rect 4275 14646 4343 14702
rect 4399 14646 4467 14702
rect 4523 14646 4591 14702
rect 4647 14646 4715 14702
rect 4771 14646 4839 14702
rect 4895 14646 4963 14702
rect 5019 14665 5045 14702
rect 5019 14646 6350 14665
rect 3339 14578 6350 14646
rect 3339 14522 4095 14578
rect 4151 14522 4219 14578
rect 4275 14522 4343 14578
rect 4399 14522 4467 14578
rect 4523 14522 4591 14578
rect 4647 14522 4715 14578
rect 4771 14522 4839 14578
rect 4895 14522 4963 14578
rect 5019 14522 6350 14578
rect 3339 14454 6350 14522
rect 3339 14398 4095 14454
rect 4151 14398 4219 14454
rect 4275 14398 4343 14454
rect 4399 14398 4467 14454
rect 4523 14398 4591 14454
rect 4647 14398 4715 14454
rect 4771 14398 4839 14454
rect 4895 14398 4963 14454
rect 5019 14398 6350 14454
rect 3339 14330 6350 14398
rect 3339 14274 4095 14330
rect 4151 14274 4219 14330
rect 4275 14274 4343 14330
rect 4399 14274 4467 14330
rect 4523 14274 4591 14330
rect 4647 14274 4715 14330
rect 4771 14274 4839 14330
rect 4895 14274 4963 14330
rect 5019 14274 6350 14330
rect 3339 14206 6350 14274
rect 3339 14150 4095 14206
rect 4151 14150 4219 14206
rect 4275 14150 4343 14206
rect 4399 14150 4467 14206
rect 4523 14150 4591 14206
rect 4647 14150 4715 14206
rect 4771 14150 4839 14206
rect 4895 14150 4963 14206
rect 5019 14150 6350 14206
rect 3339 14082 6350 14150
rect 3339 14026 4095 14082
rect 4151 14026 4219 14082
rect 4275 14026 4343 14082
rect 4399 14026 4467 14082
rect 4523 14026 4591 14082
rect 4647 14026 4715 14082
rect 4771 14026 4839 14082
rect 4895 14026 4963 14082
rect 5019 14026 6350 14082
rect 3339 13958 6350 14026
rect 3339 13902 4095 13958
rect 4151 13902 4219 13958
rect 4275 13902 4343 13958
rect 4399 13902 4467 13958
rect 4523 13902 4591 13958
rect 4647 13902 4715 13958
rect 4771 13902 4839 13958
rect 4895 13902 4963 13958
rect 5019 13902 6350 13958
rect 3339 13855 6350 13902
rect 3339 13228 6350 13312
rect 3339 13172 3631 13228
rect 3687 13172 3755 13228
rect 3811 13172 3879 13228
rect 3935 13172 6350 13228
rect 3339 13104 6350 13172
rect 3339 13048 3631 13104
rect 3687 13048 3755 13104
rect 3811 13048 3879 13104
rect 3935 13048 6350 13104
rect 3339 12980 6350 13048
rect 3339 12924 3631 12980
rect 3687 12924 3755 12980
rect 3811 12924 3879 12980
rect 3935 12924 6350 12980
rect 3339 12856 6350 12924
rect 3339 12800 3631 12856
rect 3687 12800 3755 12856
rect 3811 12800 3879 12856
rect 3935 12800 6350 12856
rect 3339 12732 6350 12800
rect 3339 12676 3631 12732
rect 3687 12676 3755 12732
rect 3811 12676 3879 12732
rect 3935 12676 6350 12732
rect 3339 12608 6350 12676
rect 3339 12552 3631 12608
rect 3687 12552 3755 12608
rect 3811 12552 3879 12608
rect 3935 12552 6350 12608
rect 3339 12484 6350 12552
rect 3339 12428 3631 12484
rect 3687 12428 3755 12484
rect 3811 12428 3879 12484
rect 3935 12428 6350 12484
rect 3339 12360 6350 12428
rect 3339 12304 3631 12360
rect 3687 12304 3755 12360
rect 3811 12304 3879 12360
rect 3935 12304 6350 12360
rect 3339 12236 6350 12304
rect 3339 12180 3631 12236
rect 3687 12180 3755 12236
rect 3811 12180 3879 12236
rect 3935 12180 6350 12236
rect 3339 12112 6350 12180
rect 3339 12056 3631 12112
rect 3687 12056 3755 12112
rect 3811 12056 3879 12112
rect 3935 12056 6350 12112
rect 3339 11995 6350 12056
rect 3339 11292 6350 11334
rect 3339 11236 4095 11292
rect 4151 11236 4219 11292
rect 4275 11236 4343 11292
rect 4399 11236 4467 11292
rect 4523 11236 4591 11292
rect 4647 11236 4715 11292
rect 4771 11236 4839 11292
rect 4895 11236 4963 11292
rect 5019 11236 6350 11292
rect 3339 11168 6350 11236
rect 3339 11112 4095 11168
rect 4151 11112 4219 11168
rect 4275 11112 4343 11168
rect 4399 11112 4467 11168
rect 4523 11112 4591 11168
rect 4647 11112 4715 11168
rect 4771 11112 4839 11168
rect 4895 11112 4963 11168
rect 5019 11112 6350 11168
rect 3339 11044 6350 11112
rect 3339 10988 4095 11044
rect 4151 10988 4219 11044
rect 4275 10988 4343 11044
rect 4399 10988 4467 11044
rect 4523 10988 4591 11044
rect 4647 10988 4715 11044
rect 4771 10988 4839 11044
rect 4895 10988 4963 11044
rect 5019 10988 6350 11044
rect 3339 10920 6350 10988
rect 3339 10864 4095 10920
rect 4151 10864 4219 10920
rect 4275 10864 4343 10920
rect 4399 10864 4467 10920
rect 4523 10864 4591 10920
rect 4647 10864 4715 10920
rect 4771 10864 4839 10920
rect 4895 10864 4963 10920
rect 5019 10864 6350 10920
rect 3339 10796 6350 10864
rect 3339 10740 4095 10796
rect 4151 10740 4219 10796
rect 4275 10740 4343 10796
rect 4399 10740 4467 10796
rect 4523 10740 4591 10796
rect 4647 10740 4715 10796
rect 4771 10740 4839 10796
rect 4895 10740 4963 10796
rect 5019 10740 6350 10796
rect 3339 10672 6350 10740
rect 3339 10616 4095 10672
rect 4151 10616 4219 10672
rect 4275 10616 4343 10672
rect 4399 10616 4467 10672
rect 4523 10616 4591 10672
rect 4647 10616 4715 10672
rect 4771 10616 4839 10672
rect 4895 10616 4963 10672
rect 5019 10616 6350 10672
rect 3339 10548 6350 10616
rect 3339 10492 4095 10548
rect 4151 10492 4219 10548
rect 4275 10492 4343 10548
rect 4399 10492 4467 10548
rect 4523 10492 4591 10548
rect 4647 10492 4715 10548
rect 4771 10492 4839 10548
rect 4895 10492 4963 10548
rect 5019 10492 6350 10548
rect 3339 10424 6350 10492
rect 3339 10368 4095 10424
rect 4151 10368 4219 10424
rect 4275 10368 4343 10424
rect 4399 10368 4467 10424
rect 4523 10368 4591 10424
rect 4647 10368 4715 10424
rect 4771 10368 4839 10424
rect 4895 10368 4963 10424
rect 5019 10368 6350 10424
rect 3339 10300 6350 10368
rect 3339 10244 4095 10300
rect 4151 10244 4219 10300
rect 4275 10244 4343 10300
rect 4399 10244 4467 10300
rect 4523 10244 4591 10300
rect 4647 10244 4715 10300
rect 4771 10244 4839 10300
rect 4895 10244 4963 10300
rect 5019 10244 6350 10300
rect 3339 10176 6350 10244
rect 3339 10120 4095 10176
rect 4151 10120 4219 10176
rect 4275 10120 4343 10176
rect 4399 10120 4467 10176
rect 4523 10120 4591 10176
rect 4647 10120 4715 10176
rect 4771 10120 4839 10176
rect 4895 10120 4963 10176
rect 5019 10120 6350 10176
rect 3339 10052 6350 10120
rect 3339 9996 4095 10052
rect 4151 9996 4219 10052
rect 4275 9996 4343 10052
rect 4399 9996 4467 10052
rect 4523 9996 4591 10052
rect 4647 9996 4715 10052
rect 4771 9996 4839 10052
rect 4895 9996 4963 10052
rect 5019 9996 6350 10052
rect 3339 9971 6350 9996
rect 3339 9392 6350 9415
rect 3339 9336 3631 9392
rect 3687 9336 3755 9392
rect 3811 9336 3879 9392
rect 3935 9336 6350 9392
rect 3339 9268 6350 9336
rect 3339 9212 3631 9268
rect 3687 9212 3755 9268
rect 3811 9212 3879 9268
rect 3935 9212 6350 9268
rect 3339 9144 6350 9212
rect 3339 9088 3631 9144
rect 3687 9088 3755 9144
rect 3811 9088 3879 9144
rect 3935 9088 6350 9144
rect 3339 9020 6350 9088
rect 3339 8964 3631 9020
rect 3687 8964 3755 9020
rect 3811 8964 3879 9020
rect 3935 8964 6350 9020
rect 3339 8896 6350 8964
rect 3339 8840 3631 8896
rect 3687 8840 3755 8896
rect 3811 8840 3879 8896
rect 3935 8840 6350 8896
rect 3339 8801 6350 8840
rect 3339 8772 4353 8801
rect 3339 8716 3631 8772
rect 3687 8716 3755 8772
rect 3811 8716 3879 8772
rect 3935 8716 4353 8772
rect 3339 8648 4353 8716
rect 3339 8592 3631 8648
rect 3687 8592 3755 8648
rect 3811 8592 3879 8648
rect 3935 8592 4353 8648
rect 3339 8524 4353 8592
rect 3339 8468 3631 8524
rect 3687 8468 3755 8524
rect 3811 8468 3879 8524
rect 3935 8468 4353 8524
rect 3339 8400 4353 8468
rect 3339 8344 3631 8400
rect 3687 8344 3755 8400
rect 3811 8344 3879 8400
rect 3935 8344 4353 8400
rect 3339 8276 4353 8344
rect 3339 8220 3631 8276
rect 3687 8220 3755 8276
rect 3811 8220 3879 8276
rect 3935 8220 4353 8276
rect 3339 8152 4353 8220
rect 3339 8096 3631 8152
rect 3687 8096 3755 8152
rect 3811 8096 3879 8152
rect 3935 8096 4353 8152
rect 3339 8028 4353 8096
rect 3339 7972 3631 8028
rect 3687 7972 3755 8028
rect 3811 7972 3879 8028
rect 3935 8018 4353 8028
rect 3935 7972 6350 8018
rect 3339 7904 6350 7972
rect 3339 7848 3631 7904
rect 3687 7848 3755 7904
rect 3811 7848 3879 7904
rect 3935 7848 6350 7904
rect 3339 7780 6350 7848
rect 3339 7724 3631 7780
rect 3687 7724 3755 7780
rect 3811 7724 3879 7780
rect 3935 7724 6350 7780
rect 3339 7656 6350 7724
rect 3339 7600 3631 7656
rect 3687 7600 3755 7656
rect 3811 7600 3879 7656
rect 3935 7600 6350 7656
rect 3339 7585 6350 7600
rect 3339 7435 6350 7448
rect 3339 7379 4095 7435
rect 4151 7379 4219 7435
rect 4275 7379 4343 7435
rect 4399 7379 4467 7435
rect 4523 7379 4591 7435
rect 4647 7379 4715 7435
rect 4771 7379 4839 7435
rect 4895 7379 4963 7435
rect 5019 7379 6350 7435
rect 3339 7311 6350 7379
rect 3339 7255 4095 7311
rect 4151 7255 4219 7311
rect 4275 7255 4343 7311
rect 4399 7255 4467 7311
rect 4523 7255 4591 7311
rect 4647 7255 4715 7311
rect 4771 7255 4839 7311
rect 4895 7255 4963 7311
rect 5019 7255 6350 7311
rect 3339 7187 6350 7255
rect 3339 7131 4095 7187
rect 4151 7131 4219 7187
rect 4275 7131 4343 7187
rect 4399 7131 4467 7187
rect 4523 7131 4591 7187
rect 4647 7131 4715 7187
rect 4771 7131 4839 7187
rect 4895 7131 4963 7187
rect 5019 7131 6350 7187
rect 3339 7063 6350 7131
rect 3339 7007 4095 7063
rect 4151 7007 4219 7063
rect 4275 7007 4343 7063
rect 4399 7007 4467 7063
rect 4523 7007 4591 7063
rect 4647 7007 4715 7063
rect 4771 7007 4839 7063
rect 4895 7007 4963 7063
rect 5019 7007 6350 7063
rect 3339 6992 6350 7007
rect 3339 6939 5051 6992
rect 3339 6883 4095 6939
rect 4151 6883 4219 6939
rect 4275 6883 4343 6939
rect 4399 6883 4467 6939
rect 4523 6883 4591 6939
rect 4647 6883 4715 6939
rect 4771 6883 4839 6939
rect 4895 6883 4963 6939
rect 5019 6883 5051 6939
rect 3339 6815 5051 6883
rect 3339 6759 4095 6815
rect 4151 6759 4219 6815
rect 4275 6759 4343 6815
rect 4399 6759 4467 6815
rect 4523 6759 4591 6815
rect 4647 6759 4715 6815
rect 4771 6759 4839 6815
rect 4895 6759 4963 6815
rect 5019 6759 5051 6815
rect 3339 6691 5051 6759
rect 3339 6635 4095 6691
rect 4151 6635 4219 6691
rect 4275 6635 4343 6691
rect 4399 6635 4467 6691
rect 4523 6635 4591 6691
rect 4647 6635 4715 6691
rect 4771 6635 4839 6691
rect 4895 6635 4963 6691
rect 5019 6635 5051 6691
rect 3339 6567 5051 6635
rect 3339 6511 4095 6567
rect 4151 6511 4219 6567
rect 4275 6511 4343 6567
rect 4399 6511 4467 6567
rect 4523 6511 4591 6567
rect 4647 6511 4715 6567
rect 4771 6511 4839 6567
rect 4895 6511 4963 6567
rect 5019 6511 5051 6567
rect 3339 6443 5051 6511
rect 3339 6387 4095 6443
rect 4151 6387 4219 6443
rect 4275 6387 4343 6443
rect 4399 6387 4467 6443
rect 4523 6387 4591 6443
rect 4647 6387 4715 6443
rect 4771 6387 4839 6443
rect 4895 6387 4963 6443
rect 5019 6387 5051 6443
rect 3339 6334 5051 6387
rect 3339 6319 6350 6334
rect 3339 6263 4095 6319
rect 4151 6263 4219 6319
rect 4275 6263 4343 6319
rect 4399 6263 4467 6319
rect 4523 6263 4591 6319
rect 4647 6263 4715 6319
rect 4771 6263 4839 6319
rect 4895 6263 4963 6319
rect 5019 6263 6350 6319
rect 3339 6195 6350 6263
rect 3339 6139 4095 6195
rect 4151 6139 4219 6195
rect 4275 6139 4343 6195
rect 4399 6139 4467 6195
rect 4523 6139 4591 6195
rect 4647 6139 4715 6195
rect 4771 6139 4839 6195
rect 4895 6139 4963 6195
rect 5019 6139 6350 6195
rect 3339 6071 6350 6139
rect 3339 6015 4095 6071
rect 4151 6015 4219 6071
rect 4275 6015 4343 6071
rect 4399 6015 4467 6071
rect 4523 6015 4591 6071
rect 4647 6015 4715 6071
rect 4771 6015 4839 6071
rect 4895 6015 4963 6071
rect 5019 6015 6350 6071
rect 3339 5947 6350 6015
rect 3339 5891 4095 5947
rect 4151 5891 4219 5947
rect 4275 5891 4343 5947
rect 4399 5891 4467 5947
rect 4523 5891 4591 5947
rect 4647 5891 4715 5947
rect 4771 5891 4839 5947
rect 4895 5891 4963 5947
rect 5019 5891 6350 5947
rect 3339 5879 6350 5891
rect 3339 5528 6350 5591
rect 3339 5472 3631 5528
rect 3687 5472 3755 5528
rect 3811 5472 3879 5528
rect 3935 5472 6350 5528
rect 3339 5404 6350 5472
rect 3339 5348 3631 5404
rect 3687 5348 3755 5404
rect 3811 5348 3879 5404
rect 3935 5348 6350 5404
rect 3339 5280 6350 5348
rect 3339 5224 3631 5280
rect 3687 5224 3755 5280
rect 3811 5224 3879 5280
rect 3935 5239 6350 5280
rect 3935 5224 4339 5239
rect 3339 5156 4339 5224
rect 3339 5100 3631 5156
rect 3687 5100 3755 5156
rect 3811 5100 3879 5156
rect 3935 5100 4339 5156
rect 3339 5032 4339 5100
rect 3339 4976 3631 5032
rect 3687 4976 3755 5032
rect 3811 4976 3879 5032
rect 3935 4976 4339 5032
rect 3339 4908 4339 4976
rect 3339 4852 3631 4908
rect 3687 4852 3755 4908
rect 3811 4852 3879 4908
rect 3935 4852 4339 4908
rect 3339 4784 4339 4852
rect 3339 4728 3631 4784
rect 3687 4728 3755 4784
rect 3811 4728 3879 4784
rect 3935 4728 4339 4784
rect 3339 4673 4339 4728
rect 3339 4660 6350 4673
rect 3339 4604 3631 4660
rect 3687 4604 3755 4660
rect 3811 4604 3879 4660
rect 3935 4604 6350 4660
rect 3339 4536 6350 4604
rect 3339 4480 3631 4536
rect 3687 4480 3755 4536
rect 3811 4480 3879 4536
rect 3935 4480 6350 4536
rect 3339 4412 6350 4480
rect 3339 4356 3631 4412
rect 3687 4356 3755 4412
rect 3811 4356 3879 4412
rect 3935 4356 6350 4412
rect 3339 4321 6350 4356
rect 3339 4010 6350 4051
rect 3339 3954 4095 4010
rect 4151 3954 4219 4010
rect 4275 3954 4343 4010
rect 4399 3954 4467 4010
rect 4523 3954 4591 4010
rect 4647 3954 4715 4010
rect 4771 3954 4839 4010
rect 4895 3954 4963 4010
rect 5019 3954 6350 4010
rect 3339 3886 6350 3954
rect 3339 3830 4095 3886
rect 4151 3830 4219 3886
rect 4275 3830 4343 3886
rect 4399 3830 4467 3886
rect 4523 3830 4591 3886
rect 4647 3830 4715 3886
rect 4771 3830 4839 3886
rect 4895 3830 4963 3886
rect 5019 3830 6350 3886
rect 3339 3762 6350 3830
rect 3339 3706 4095 3762
rect 4151 3706 4219 3762
rect 4275 3706 4343 3762
rect 4399 3706 4467 3762
rect 4523 3706 4591 3762
rect 4647 3706 4715 3762
rect 4771 3706 4839 3762
rect 4895 3706 4963 3762
rect 5019 3706 6350 3762
rect 3339 3638 6350 3706
rect 3339 3582 4095 3638
rect 4151 3582 4219 3638
rect 4275 3582 4343 3638
rect 4399 3582 4467 3638
rect 4523 3582 4591 3638
rect 4647 3582 4715 3638
rect 4771 3582 4839 3638
rect 4895 3582 4963 3638
rect 5019 3582 6350 3638
rect 3339 3514 6350 3582
rect 3339 3458 4095 3514
rect 4151 3458 4219 3514
rect 4275 3458 4343 3514
rect 4399 3458 4467 3514
rect 4523 3458 4591 3514
rect 4647 3458 4715 3514
rect 4771 3458 4839 3514
rect 4895 3458 4963 3514
rect 5019 3458 6350 3514
rect 3339 3390 6350 3458
rect 3339 3334 4095 3390
rect 4151 3334 4219 3390
rect 4275 3334 4343 3390
rect 4399 3334 4467 3390
rect 4523 3334 4591 3390
rect 4647 3334 4715 3390
rect 4771 3334 4839 3390
rect 4895 3334 4963 3390
rect 5019 3334 6350 3390
rect 3339 3266 6350 3334
rect 3339 3210 4095 3266
rect 4151 3210 4219 3266
rect 4275 3210 4343 3266
rect 4399 3210 4467 3266
rect 4523 3210 4591 3266
rect 4647 3210 4715 3266
rect 4771 3210 4839 3266
rect 4895 3210 4963 3266
rect 5019 3210 6350 3266
rect 3339 3142 6350 3210
rect 3339 3086 4095 3142
rect 4151 3086 4219 3142
rect 4275 3086 4343 3142
rect 4399 3086 4467 3142
rect 4523 3086 4591 3142
rect 4647 3086 4715 3142
rect 4771 3086 4839 3142
rect 4895 3086 4963 3142
rect 5019 3086 6350 3142
rect 3339 3051 6350 3086
use M2_M1431059054873_128x8m81  M2_M1431059054873_128x8m81_0
timestamp 1698431365
transform 1 0 3783 0 1 36745
box 0 0 1 1
use M2_M14310590548721_128x8m81  M2_M14310590548721_128x8m81_0
timestamp 1698431365
transform 1 0 3783 0 1 23602
box 0 0 1 1
use M2_M14310590548785_128x8m81  M2_M14310590548785_128x8m81_0
timestamp 1698431365
transform 1 0 3783 0 1 4942
box 0 0 1 1
use M2_M14310590548785_128x8m81  M2_M14310590548785_128x8m81_1
timestamp 1698431365
transform 1 0 3783 0 1 12642
box 0 0 1 1
use M2_M14310590548793_128x8m81  M2_M14310590548793_128x8m81_0
timestamp 1698431365
transform 1 0 3783 0 1 17867
box 0 0 1 1
use M2_M14310590548794_128x8m81  M2_M14310590548794_128x8m81_0
timestamp 1698431365
transform 1 0 3783 0 1 8496
box 0 0 1 1
use M2_M14310590548794_128x8m81  M2_M14310590548794_128x8m81_1
timestamp 1698431365
transform 1 0 3783 0 1 29263
box 0 0 1 1
use M3_M2431059054879_128x8m81  M3_M2431059054879_128x8m81_0
timestamp 1698431365
transform 1 0 3783 0 1 23602
box 0 0 1 1
use M3_M24310590548718_128x8m81  M3_M24310590548718_128x8m81_0
timestamp 1698431365
transform 1 0 3783 0 1 36745
box 0 0 1 1
use M3_M24310590548781_128x8m81  M3_M24310590548781_128x8m81_0
timestamp 1698431365
transform 1 0 4557 0 1 3548
box 0 0 1 1
use M3_M24310590548781_128x8m81  M3_M24310590548781_128x8m81_1
timestamp 1698431365
transform 1 0 4557 0 1 25229
box 0 0 1 1
use M3_M24310590548786_128x8m81  M3_M24310590548786_128x8m81_0
timestamp 1698431365
transform 1 0 4557 0 1 6663
box 0 0 1 1
use M3_M24310590548787_128x8m81  M3_M24310590548787_128x8m81_0
timestamp 1698431365
transform 1 0 4557 0 1 33607
box 0 0 1 1
use M3_M24310590548788_128x8m81  M3_M24310590548788_128x8m81_0
timestamp 1698431365
transform 1 0 3783 0 1 17867
box 0 0 1 1
use M3_M24310590548789_128x8m81  M3_M24310590548789_128x8m81_0
timestamp 1698431365
transform 1 0 3783 0 1 8496
box 0 0 1 1
use M3_M24310590548789_128x8m81  M3_M24310590548789_128x8m81_1
timestamp 1698431365
transform 1 0 3783 0 1 29263
box 0 0 1 1
use M3_M24310590548790_128x8m81  M3_M24310590548790_128x8m81_0
timestamp 1698431365
transform 1 0 4557 0 1 14922
box 0 0 1 1
use M3_M24310590548791_128x8m81  M3_M24310590548791_128x8m81_0
timestamp 1698431365
transform 1 0 3783 0 1 4942
box 0 0 1 1
use M3_M24310590548791_128x8m81  M3_M24310590548791_128x8m81_1
timestamp 1698431365
transform 1 0 3783 0 1 12642
box 0 0 1 1
use M3_M24310590548792_128x8m81  M3_M24310590548792_128x8m81_0
timestamp 1698431365
transform 1 0 4557 0 1 10644
box 0 0 1 1
use M3_M24310590548795_128x8m81  M3_M24310590548795_128x8m81_0
timestamp 1698431365
transform 1 0 4557 0 1 21182
box 0 0 1 1
<< properties >>
string GDS_END 1476260
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 1473616
<< end >>
