magic
tech gf180mcuB
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 352 4790 870
<< pwell >>
rect -86 -86 4790 352
<< mvnmos >>
rect 124 70 244 166
rect 348 70 468 166
rect 572 70 692 166
rect 796 70 916 166
rect 1020 70 1140 166
rect 1244 70 1364 166
rect 1468 70 1588 166
rect 1692 70 1812 166
rect 1916 70 2036 166
rect 2140 70 2260 166
rect 2364 70 2484 166
rect 2588 70 2708 166
rect 2812 70 2932 166
rect 3036 70 3156 166
rect 3260 70 3380 166
rect 3484 70 3604 166
rect 3708 70 3828 166
rect 3932 70 4052 166
rect 4156 70 4276 166
rect 4380 70 4500 166
<< mvpmos >>
rect 124 472 224 716
rect 348 472 448 716
rect 572 472 672 716
rect 796 472 896 716
rect 1020 472 1120 716
rect 1244 472 1344 716
rect 1468 472 1568 716
rect 1692 472 1792 716
rect 1916 472 2016 716
rect 2140 472 2240 716
rect 2364 472 2464 716
rect 2588 472 2688 716
rect 2812 472 2912 716
rect 3036 472 3136 716
rect 3260 472 3360 716
rect 3484 472 3584 716
rect 3708 472 3808 716
rect 3932 472 4032 716
rect 4156 472 4256 716
rect 4380 472 4480 716
<< mvndiff >>
rect 36 129 124 166
rect 36 83 49 129
rect 95 83 124 129
rect 36 70 124 83
rect 244 153 348 166
rect 244 107 273 153
rect 319 107 348 153
rect 244 70 348 107
rect 468 129 572 166
rect 468 83 497 129
rect 543 83 572 129
rect 468 70 572 83
rect 692 153 796 166
rect 692 107 721 153
rect 767 107 796 153
rect 692 70 796 107
rect 916 129 1020 166
rect 916 83 945 129
rect 991 83 1020 129
rect 916 70 1020 83
rect 1140 153 1244 166
rect 1140 107 1169 153
rect 1215 107 1244 153
rect 1140 70 1244 107
rect 1364 129 1468 166
rect 1364 83 1393 129
rect 1439 83 1468 129
rect 1364 70 1468 83
rect 1588 153 1692 166
rect 1588 107 1617 153
rect 1663 107 1692 153
rect 1588 70 1692 107
rect 1812 129 1916 166
rect 1812 83 1841 129
rect 1887 83 1916 129
rect 1812 70 1916 83
rect 2036 153 2140 166
rect 2036 107 2065 153
rect 2111 107 2140 153
rect 2036 70 2140 107
rect 2260 129 2364 166
rect 2260 83 2289 129
rect 2335 83 2364 129
rect 2260 70 2364 83
rect 2484 153 2588 166
rect 2484 107 2513 153
rect 2559 107 2588 153
rect 2484 70 2588 107
rect 2708 129 2812 166
rect 2708 83 2737 129
rect 2783 83 2812 129
rect 2708 70 2812 83
rect 2932 153 3036 166
rect 2932 107 2961 153
rect 3007 107 3036 153
rect 2932 70 3036 107
rect 3156 129 3260 166
rect 3156 83 3185 129
rect 3231 83 3260 129
rect 3156 70 3260 83
rect 3380 153 3484 166
rect 3380 107 3409 153
rect 3455 107 3484 153
rect 3380 70 3484 107
rect 3604 129 3708 166
rect 3604 83 3633 129
rect 3679 83 3708 129
rect 3604 70 3708 83
rect 3828 153 3932 166
rect 3828 107 3857 153
rect 3903 107 3932 153
rect 3828 70 3932 107
rect 4052 129 4156 166
rect 4052 83 4081 129
rect 4127 83 4156 129
rect 4052 70 4156 83
rect 4276 153 4380 166
rect 4276 107 4305 153
rect 4351 107 4380 153
rect 4276 70 4380 107
rect 4500 129 4588 166
rect 4500 83 4529 129
rect 4575 83 4588 129
rect 4500 70 4588 83
<< mvpdiff >>
rect 36 665 124 716
rect 36 525 49 665
rect 95 525 124 665
rect 36 472 124 525
rect 224 665 348 716
rect 224 525 273 665
rect 319 525 348 665
rect 224 472 348 525
rect 448 703 572 716
rect 448 657 477 703
rect 523 657 572 703
rect 448 472 572 657
rect 672 665 796 716
rect 672 525 701 665
rect 747 525 796 665
rect 672 472 796 525
rect 896 703 1020 716
rect 896 657 925 703
rect 971 657 1020 703
rect 896 472 1020 657
rect 1120 665 1244 716
rect 1120 525 1149 665
rect 1195 525 1244 665
rect 1120 472 1244 525
rect 1344 703 1468 716
rect 1344 657 1373 703
rect 1419 657 1468 703
rect 1344 472 1468 657
rect 1568 665 1692 716
rect 1568 525 1597 665
rect 1643 525 1692 665
rect 1568 472 1692 525
rect 1792 703 1916 716
rect 1792 657 1821 703
rect 1867 657 1916 703
rect 1792 472 1916 657
rect 2016 665 2140 716
rect 2016 525 2045 665
rect 2091 525 2140 665
rect 2016 472 2140 525
rect 2240 703 2364 716
rect 2240 657 2269 703
rect 2315 657 2364 703
rect 2240 472 2364 657
rect 2464 665 2588 716
rect 2464 525 2493 665
rect 2539 525 2588 665
rect 2464 472 2588 525
rect 2688 703 2812 716
rect 2688 657 2717 703
rect 2763 657 2812 703
rect 2688 472 2812 657
rect 2912 665 3036 716
rect 2912 525 2941 665
rect 2987 525 3036 665
rect 2912 472 3036 525
rect 3136 703 3260 716
rect 3136 657 3165 703
rect 3211 657 3260 703
rect 3136 472 3260 657
rect 3360 665 3484 716
rect 3360 525 3389 665
rect 3435 525 3484 665
rect 3360 472 3484 525
rect 3584 703 3708 716
rect 3584 657 3613 703
rect 3659 657 3708 703
rect 3584 472 3708 657
rect 3808 665 3932 716
rect 3808 525 3837 665
rect 3883 525 3932 665
rect 3808 472 3932 525
rect 4032 703 4156 716
rect 4032 657 4061 703
rect 4107 657 4156 703
rect 4032 472 4156 657
rect 4256 665 4380 716
rect 4256 525 4285 665
rect 4331 525 4380 665
rect 4256 472 4380 525
rect 4480 665 4568 716
rect 4480 525 4509 665
rect 4555 525 4568 665
rect 4480 472 4568 525
<< mvndiffc >>
rect 49 83 95 129
rect 273 107 319 153
rect 497 83 543 129
rect 721 107 767 153
rect 945 83 991 129
rect 1169 107 1215 153
rect 1393 83 1439 129
rect 1617 107 1663 153
rect 1841 83 1887 129
rect 2065 107 2111 153
rect 2289 83 2335 129
rect 2513 107 2559 153
rect 2737 83 2783 129
rect 2961 107 3007 153
rect 3185 83 3231 129
rect 3409 107 3455 153
rect 3633 83 3679 129
rect 3857 107 3903 153
rect 4081 83 4127 129
rect 4305 107 4351 153
rect 4529 83 4575 129
<< mvpdiffc >>
rect 49 525 95 665
rect 273 525 319 665
rect 477 657 523 703
rect 701 525 747 665
rect 925 657 971 703
rect 1149 525 1195 665
rect 1373 657 1419 703
rect 1597 525 1643 665
rect 1821 657 1867 703
rect 2045 525 2091 665
rect 2269 657 2315 703
rect 2493 525 2539 665
rect 2717 657 2763 703
rect 2941 525 2987 665
rect 3165 657 3211 703
rect 3389 525 3435 665
rect 3613 657 3659 703
rect 3837 525 3883 665
rect 4061 657 4107 703
rect 4285 525 4331 665
rect 4509 525 4555 665
<< polysilicon >>
rect 124 716 224 760
rect 348 716 448 760
rect 572 716 672 760
rect 796 716 896 760
rect 1020 716 1120 760
rect 1244 716 1344 760
rect 1468 716 1568 760
rect 1692 716 1792 760
rect 1916 716 2016 760
rect 2140 716 2240 760
rect 2364 716 2464 760
rect 2588 716 2688 760
rect 2812 716 2912 760
rect 3036 716 3136 760
rect 3260 716 3360 760
rect 3484 716 3584 760
rect 3708 716 3808 760
rect 3932 716 4032 760
rect 4156 716 4256 760
rect 4380 716 4480 760
rect 124 407 224 472
rect 348 407 448 472
rect 572 407 672 472
rect 796 407 896 472
rect 1020 407 1120 472
rect 1244 407 1344 472
rect 1468 407 1568 472
rect 1692 407 1792 472
rect 1916 407 2016 472
rect 2140 407 2240 472
rect 2364 407 2464 472
rect 2588 407 2688 472
rect 2812 407 2912 472
rect 3036 407 3136 472
rect 3260 407 3360 472
rect 3484 407 3584 472
rect 3708 407 3808 472
rect 3932 407 4032 472
rect 4156 407 4256 472
rect 4380 407 4480 472
rect 124 394 4480 407
rect 124 348 137 394
rect 1969 348 2515 394
rect 4441 348 4480 394
rect 124 335 4480 348
rect 124 166 244 335
rect 348 166 468 335
rect 572 166 692 335
rect 796 166 916 335
rect 1020 166 1140 335
rect 1244 166 1364 335
rect 1468 166 1588 335
rect 1692 166 1812 335
rect 1916 166 2036 335
rect 2140 166 2260 335
rect 2364 166 2484 335
rect 2588 166 2708 335
rect 2812 166 2932 335
rect 3036 166 3156 335
rect 3260 166 3380 335
rect 3484 166 3604 335
rect 3708 166 3828 335
rect 3932 166 4052 335
rect 4156 166 4276 335
rect 4380 288 4480 335
rect 4380 166 4500 288
rect 124 24 244 70
rect 348 24 468 70
rect 572 24 692 70
rect 796 24 916 70
rect 1020 24 1140 70
rect 1244 24 1364 70
rect 1468 24 1588 70
rect 1692 24 1812 70
rect 1916 24 2036 70
rect 2140 24 2260 70
rect 2364 24 2484 70
rect 2588 24 2708 70
rect 2812 24 2932 70
rect 3036 24 3156 70
rect 3260 24 3380 70
rect 3484 24 3604 70
rect 3708 24 3828 70
rect 3932 24 4052 70
rect 4156 24 4276 70
rect 4380 24 4500 70
<< polycontact >>
rect 137 348 1969 394
rect 2515 348 4441 394
<< metal1 >>
rect 0 724 4704 844
rect 49 665 95 724
rect 466 703 534 724
rect 49 506 95 525
rect 273 665 319 676
rect 466 657 477 703
rect 523 657 534 703
rect 914 703 982 724
rect 701 665 747 676
rect 319 525 701 611
rect 914 657 925 703
rect 971 657 982 703
rect 1362 703 1430 724
rect 1149 665 1195 676
rect 747 525 1149 611
rect 1362 657 1373 703
rect 1419 657 1430 703
rect 1810 703 1878 724
rect 1597 665 1643 676
rect 1195 525 1597 611
rect 1810 657 1821 703
rect 1867 657 1878 703
rect 2258 703 2326 724
rect 2034 665 2110 676
rect 2034 611 2045 665
rect 1643 525 2045 611
rect 2091 611 2110 665
rect 2258 657 2269 703
rect 2315 657 2326 703
rect 2706 703 2774 724
rect 2493 665 2539 676
rect 2091 525 2493 611
rect 2706 657 2717 703
rect 2763 657 2774 703
rect 3154 703 3222 724
rect 2941 665 2987 676
rect 2539 525 2941 611
rect 3154 657 3165 703
rect 3211 657 3222 703
rect 3602 703 3670 724
rect 3389 665 3435 676
rect 2987 525 3389 611
rect 3602 657 3613 703
rect 3659 657 3670 703
rect 4050 703 4118 724
rect 3837 665 3883 676
rect 3435 525 3837 611
rect 4050 657 4061 703
rect 4107 657 4118 703
rect 4285 665 4331 676
rect 3883 525 4285 611
rect 273 470 4331 525
rect 4509 665 4555 724
rect 4509 506 4555 525
rect 126 394 1980 424
rect 126 348 137 394
rect 1969 348 1980 394
rect 2206 301 2386 470
rect 2504 394 4480 424
rect 2504 348 2515 394
rect 4441 348 4480 394
rect 262 175 4362 301
rect 262 153 330 175
rect 49 129 95 140
rect 262 107 273 153
rect 319 107 330 153
rect 710 153 778 175
rect 49 60 95 83
rect 486 83 497 129
rect 543 83 554 129
rect 710 107 721 153
rect 767 107 778 153
rect 1158 153 1226 175
rect 486 60 554 83
rect 934 83 945 129
rect 991 83 1002 129
rect 1158 107 1169 153
rect 1215 107 1226 153
rect 1606 153 1674 175
rect 934 60 1002 83
rect 1382 83 1393 129
rect 1439 83 1450 129
rect 1606 107 1617 153
rect 1663 107 1674 153
rect 2054 153 2122 175
rect 1382 60 1450 83
rect 1830 83 1841 129
rect 1887 83 1898 129
rect 2054 107 2065 153
rect 2111 107 2122 153
rect 2502 153 2570 175
rect 1830 60 1898 83
rect 2278 83 2289 129
rect 2335 83 2346 129
rect 2502 107 2513 153
rect 2559 107 2570 153
rect 2950 153 3018 175
rect 2278 60 2346 83
rect 2726 83 2737 129
rect 2783 83 2794 129
rect 2950 107 2961 153
rect 3007 107 3018 153
rect 3398 153 3466 175
rect 2726 60 2794 83
rect 3174 83 3185 129
rect 3231 83 3242 129
rect 3398 107 3409 153
rect 3455 107 3466 153
rect 3846 153 3914 175
rect 3174 60 3242 83
rect 3622 83 3633 129
rect 3679 83 3690 129
rect 3846 107 3857 153
rect 3903 107 3914 153
rect 4294 153 4362 175
rect 3622 60 3690 83
rect 4070 83 4081 129
rect 4127 83 4138 129
rect 4294 107 4305 153
rect 4351 107 4362 153
rect 4070 60 4138 83
rect 4518 83 4529 129
rect 4575 83 4586 129
rect 4518 60 4586 83
rect 0 -60 4704 60
<< labels >>
flabel metal1 s 0 724 4704 844 0 FreeSans 600 0 0 0 VDD
port 3 nsew power bidirectional abutment
flabel metal1 s 49 129 95 140 0 FreeSans 600 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel metal1 s 4285 611 4331 676 0 FreeSans 600 0 0 0 ZN
port 2 nsew default output
flabel metal1 s 126 348 1980 424 0 FreeSans 600 0 0 0 I
port 1 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 4 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 2504 348 4480 424 1 I
port 1 nsew default input
rlabel metal1 s 3837 611 3883 676 1 ZN
port 2 nsew default output
rlabel metal1 s 3389 611 3435 676 1 ZN
port 2 nsew default output
rlabel metal1 s 2941 611 2987 676 1 ZN
port 2 nsew default output
rlabel metal1 s 2493 611 2539 676 1 ZN
port 2 nsew default output
rlabel metal1 s 2034 611 2110 676 1 ZN
port 2 nsew default output
rlabel metal1 s 1597 611 1643 676 1 ZN
port 2 nsew default output
rlabel metal1 s 1149 611 1195 676 1 ZN
port 2 nsew default output
rlabel metal1 s 701 611 747 676 1 ZN
port 2 nsew default output
rlabel metal1 s 273 611 319 676 1 ZN
port 2 nsew default output
rlabel metal1 s 273 470 4331 611 1 ZN
port 2 nsew default output
rlabel metal1 s 2206 301 2386 470 1 ZN
port 2 nsew default output
rlabel metal1 s 262 175 4362 301 1 ZN
port 2 nsew default output
rlabel metal1 s 4294 107 4362 175 1 ZN
port 2 nsew default output
rlabel metal1 s 3846 107 3914 175 1 ZN
port 2 nsew default output
rlabel metal1 s 3398 107 3466 175 1 ZN
port 2 nsew default output
rlabel metal1 s 2950 107 3018 175 1 ZN
port 2 nsew default output
rlabel metal1 s 2502 107 2570 175 1 ZN
port 2 nsew default output
rlabel metal1 s 2054 107 2122 175 1 ZN
port 2 nsew default output
rlabel metal1 s 1606 107 1674 175 1 ZN
port 2 nsew default output
rlabel metal1 s 1158 107 1226 175 1 ZN
port 2 nsew default output
rlabel metal1 s 710 107 778 175 1 ZN
port 2 nsew default output
rlabel metal1 s 262 107 330 175 1 ZN
port 2 nsew default output
rlabel metal1 s 4509 657 4555 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4050 657 4118 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3602 657 3670 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3154 657 3222 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2706 657 2774 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2258 657 2326 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1810 657 1878 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1362 657 1430 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 914 657 982 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 466 657 534 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 657 95 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4509 506 4555 657 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 506 95 657 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4518 60 4586 129 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 4070 60 4138 129 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3622 60 3690 129 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3174 60 3242 129 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2726 60 2794 129 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2278 60 2346 129 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1830 60 1898 129 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1382 60 1450 129 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 934 60 1002 129 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 486 60 554 129 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 129 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 4704 60 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4704 784
string GDS_END 857594
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 847270
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
