magic
tech gf180mcuB
magscale 1 10
timestamp 1698431365
<< metal2 >>
rect -400 12949 13200 13065
rect -400 12893 -254 12949
rect -198 12893 -130 12949
rect -74 12893 -6 12949
rect 50 12893 118 12949
rect 174 12893 242 12949
rect 298 12893 366 12949
rect 422 12893 490 12949
rect 546 12893 614 12949
rect 670 12893 738 12949
rect 794 12893 862 12949
rect 918 12893 986 12949
rect 1042 12893 1110 12949
rect 1166 12893 1234 12949
rect 1290 12893 1358 12949
rect 1414 12893 1482 12949
rect 1538 12893 1606 12949
rect 1662 12893 1730 12949
rect 1786 12893 1854 12949
rect 1910 12893 1978 12949
rect 2034 12893 2102 12949
rect 2158 12893 2226 12949
rect 2282 12893 2350 12949
rect 2406 12893 2474 12949
rect 2530 12893 2598 12949
rect 2654 12893 2722 12949
rect 2778 12893 2846 12949
rect 2902 12893 2970 12949
rect 3026 12893 3094 12949
rect 3150 12893 3218 12949
rect 3274 12893 3342 12949
rect 3398 12893 3466 12949
rect 3522 12893 3590 12949
rect 3646 12893 3714 12949
rect 3770 12893 3838 12949
rect 3894 12893 3962 12949
rect 4018 12893 4086 12949
rect 4142 12893 4210 12949
rect 4266 12893 4334 12949
rect 4390 12893 4458 12949
rect 4514 12893 4582 12949
rect 4638 12893 4706 12949
rect 4762 12893 4830 12949
rect 4886 12893 4954 12949
rect 5010 12893 5078 12949
rect 5134 12893 5202 12949
rect 5258 12893 5326 12949
rect 5382 12893 5450 12949
rect 5506 12893 5574 12949
rect 5630 12893 5698 12949
rect 5754 12893 5822 12949
rect 5878 12893 5946 12949
rect 6002 12893 6070 12949
rect 6126 12893 6194 12949
rect 6250 12893 6318 12949
rect 6374 12893 6442 12949
rect 6498 12893 6566 12949
rect 6622 12893 6690 12949
rect 6746 12893 6814 12949
rect 6870 12893 6938 12949
rect 6994 12893 7062 12949
rect 7118 12893 7186 12949
rect 7242 12893 7310 12949
rect 7366 12893 7434 12949
rect 7490 12893 7558 12949
rect 7614 12893 7682 12949
rect 7738 12893 7806 12949
rect 7862 12893 7930 12949
rect 7986 12893 8054 12949
rect 8110 12893 8178 12949
rect 8234 12893 8302 12949
rect 8358 12893 8426 12949
rect 8482 12893 8550 12949
rect 8606 12893 8674 12949
rect 8730 12893 8798 12949
rect 8854 12893 8922 12949
rect 8978 12893 9046 12949
rect 9102 12893 9170 12949
rect 9226 12893 9294 12949
rect 9350 12893 9418 12949
rect 9474 12893 9542 12949
rect 9598 12893 9666 12949
rect 9722 12893 9790 12949
rect 9846 12893 9914 12949
rect 9970 12893 10038 12949
rect 10094 12893 10162 12949
rect 10218 12893 10286 12949
rect 10342 12893 10410 12949
rect 10466 12893 10534 12949
rect 10590 12893 10658 12949
rect 10714 12893 10782 12949
rect 10838 12893 10906 12949
rect 10962 12893 11030 12949
rect 11086 12893 11154 12949
rect 11210 12893 11278 12949
rect 11334 12893 11402 12949
rect 11458 12893 11526 12949
rect 11582 12893 11650 12949
rect 11706 12893 11774 12949
rect 11830 12893 11898 12949
rect 11954 12893 12022 12949
rect 12078 12893 12146 12949
rect 12202 12893 12270 12949
rect 12326 12893 12394 12949
rect 12450 12893 12518 12949
rect 12574 12893 12642 12949
rect 12698 12893 12766 12949
rect 12822 12893 12890 12949
rect 12946 12893 13014 12949
rect 13070 12893 13200 12949
rect -400 12825 13200 12893
rect -400 12769 -254 12825
rect -198 12769 -130 12825
rect -74 12769 -6 12825
rect 50 12769 118 12825
rect 174 12769 242 12825
rect 298 12769 366 12825
rect 422 12769 490 12825
rect 546 12769 614 12825
rect 670 12769 738 12825
rect 794 12769 862 12825
rect 918 12769 986 12825
rect 1042 12769 1110 12825
rect 1166 12769 1234 12825
rect 1290 12769 1358 12825
rect 1414 12769 1482 12825
rect 1538 12769 1606 12825
rect 1662 12769 1730 12825
rect 1786 12769 1854 12825
rect 1910 12769 1978 12825
rect 2034 12769 2102 12825
rect 2158 12769 2226 12825
rect 2282 12769 2350 12825
rect 2406 12769 2474 12825
rect 2530 12769 2598 12825
rect 2654 12769 2722 12825
rect 2778 12769 2846 12825
rect 2902 12769 2970 12825
rect 3026 12769 3094 12825
rect 3150 12769 3218 12825
rect 3274 12769 3342 12825
rect 3398 12769 3466 12825
rect 3522 12769 3590 12825
rect 3646 12769 3714 12825
rect 3770 12769 3838 12825
rect 3894 12769 3962 12825
rect 4018 12769 4086 12825
rect 4142 12769 4210 12825
rect 4266 12769 4334 12825
rect 4390 12769 4458 12825
rect 4514 12769 4582 12825
rect 4638 12769 4706 12825
rect 4762 12769 4830 12825
rect 4886 12769 4954 12825
rect 5010 12769 5078 12825
rect 5134 12769 5202 12825
rect 5258 12769 5326 12825
rect 5382 12769 5450 12825
rect 5506 12769 5574 12825
rect 5630 12769 5698 12825
rect 5754 12769 5822 12825
rect 5878 12769 5946 12825
rect 6002 12769 6070 12825
rect 6126 12769 6194 12825
rect 6250 12769 6318 12825
rect 6374 12769 6442 12825
rect 6498 12769 6566 12825
rect 6622 12769 6690 12825
rect 6746 12769 6814 12825
rect 6870 12769 6938 12825
rect 6994 12769 7062 12825
rect 7118 12769 7186 12825
rect 7242 12769 7310 12825
rect 7366 12769 7434 12825
rect 7490 12769 7558 12825
rect 7614 12769 7682 12825
rect 7738 12769 7806 12825
rect 7862 12769 7930 12825
rect 7986 12769 8054 12825
rect 8110 12769 8178 12825
rect 8234 12769 8302 12825
rect 8358 12769 8426 12825
rect 8482 12769 8550 12825
rect 8606 12769 8674 12825
rect 8730 12769 8798 12825
rect 8854 12769 8922 12825
rect 8978 12769 9046 12825
rect 9102 12769 9170 12825
rect 9226 12769 9294 12825
rect 9350 12769 9418 12825
rect 9474 12769 9542 12825
rect 9598 12769 9666 12825
rect 9722 12769 9790 12825
rect 9846 12769 9914 12825
rect 9970 12769 10038 12825
rect 10094 12769 10162 12825
rect 10218 12769 10286 12825
rect 10342 12769 10410 12825
rect 10466 12769 10534 12825
rect 10590 12769 10658 12825
rect 10714 12769 10782 12825
rect 10838 12769 10906 12825
rect 10962 12769 11030 12825
rect 11086 12769 11154 12825
rect 11210 12769 11278 12825
rect 11334 12769 11402 12825
rect 11458 12769 11526 12825
rect 11582 12769 11650 12825
rect 11706 12769 11774 12825
rect 11830 12769 11898 12825
rect 11954 12769 12022 12825
rect 12078 12769 12146 12825
rect 12202 12769 12270 12825
rect 12326 12769 12394 12825
rect 12450 12769 12518 12825
rect 12574 12769 12642 12825
rect 12698 12769 12766 12825
rect 12822 12769 12890 12825
rect 12946 12769 13014 12825
rect 13070 12769 13200 12825
rect -400 12701 13200 12769
rect -400 12645 -254 12701
rect -198 12645 -130 12701
rect -74 12645 -6 12701
rect 50 12645 118 12701
rect 174 12645 242 12701
rect 298 12645 366 12701
rect 422 12645 490 12701
rect 546 12645 614 12701
rect 670 12645 738 12701
rect 794 12645 862 12701
rect 918 12645 986 12701
rect 1042 12645 1110 12701
rect 1166 12645 1234 12701
rect 1290 12645 1358 12701
rect 1414 12645 1482 12701
rect 1538 12645 1606 12701
rect 1662 12645 1730 12701
rect 1786 12645 1854 12701
rect 1910 12645 1978 12701
rect 2034 12645 2102 12701
rect 2158 12645 2226 12701
rect 2282 12645 2350 12701
rect 2406 12645 2474 12701
rect 2530 12645 2598 12701
rect 2654 12645 2722 12701
rect 2778 12645 2846 12701
rect 2902 12645 2970 12701
rect 3026 12645 3094 12701
rect 3150 12645 3218 12701
rect 3274 12645 3342 12701
rect 3398 12645 3466 12701
rect 3522 12645 3590 12701
rect 3646 12645 3714 12701
rect 3770 12645 3838 12701
rect 3894 12645 3962 12701
rect 4018 12645 4086 12701
rect 4142 12645 4210 12701
rect 4266 12645 4334 12701
rect 4390 12645 4458 12701
rect 4514 12645 4582 12701
rect 4638 12645 4706 12701
rect 4762 12645 4830 12701
rect 4886 12645 4954 12701
rect 5010 12645 5078 12701
rect 5134 12645 5202 12701
rect 5258 12645 5326 12701
rect 5382 12645 5450 12701
rect 5506 12645 5574 12701
rect 5630 12645 5698 12701
rect 5754 12645 5822 12701
rect 5878 12645 5946 12701
rect 6002 12645 6070 12701
rect 6126 12645 6194 12701
rect 6250 12645 6318 12701
rect 6374 12645 6442 12701
rect 6498 12645 6566 12701
rect 6622 12645 6690 12701
rect 6746 12645 6814 12701
rect 6870 12645 6938 12701
rect 6994 12645 7062 12701
rect 7118 12645 7186 12701
rect 7242 12645 7310 12701
rect 7366 12645 7434 12701
rect 7490 12645 7558 12701
rect 7614 12645 7682 12701
rect 7738 12645 7806 12701
rect 7862 12645 7930 12701
rect 7986 12645 8054 12701
rect 8110 12645 8178 12701
rect 8234 12645 8302 12701
rect 8358 12645 8426 12701
rect 8482 12645 8550 12701
rect 8606 12645 8674 12701
rect 8730 12645 8798 12701
rect 8854 12645 8922 12701
rect 8978 12645 9046 12701
rect 9102 12645 9170 12701
rect 9226 12645 9294 12701
rect 9350 12645 9418 12701
rect 9474 12645 9542 12701
rect 9598 12645 9666 12701
rect 9722 12645 9790 12701
rect 9846 12645 9914 12701
rect 9970 12645 10038 12701
rect 10094 12645 10162 12701
rect 10218 12645 10286 12701
rect 10342 12645 10410 12701
rect 10466 12645 10534 12701
rect 10590 12645 10658 12701
rect 10714 12645 10782 12701
rect 10838 12645 10906 12701
rect 10962 12645 11030 12701
rect 11086 12645 11154 12701
rect 11210 12645 11278 12701
rect 11334 12645 11402 12701
rect 11458 12645 11526 12701
rect 11582 12645 11650 12701
rect 11706 12645 11774 12701
rect 11830 12645 11898 12701
rect 11954 12645 12022 12701
rect 12078 12645 12146 12701
rect 12202 12645 12270 12701
rect 12326 12645 12394 12701
rect 12450 12645 12518 12701
rect 12574 12645 12642 12701
rect 12698 12645 12766 12701
rect 12822 12645 12890 12701
rect 12946 12645 13014 12701
rect 13070 12645 13200 12701
rect -400 12577 13200 12645
rect -400 12521 -254 12577
rect -198 12521 -130 12577
rect -74 12521 -6 12577
rect 50 12521 118 12577
rect 174 12521 242 12577
rect 298 12521 366 12577
rect 422 12521 490 12577
rect 546 12521 614 12577
rect 670 12521 738 12577
rect 794 12521 862 12577
rect 918 12521 986 12577
rect 1042 12521 1110 12577
rect 1166 12521 1234 12577
rect 1290 12521 1358 12577
rect 1414 12521 1482 12577
rect 1538 12521 1606 12577
rect 1662 12521 1730 12577
rect 1786 12521 1854 12577
rect 1910 12521 1978 12577
rect 2034 12521 2102 12577
rect 2158 12521 2226 12577
rect 2282 12521 2350 12577
rect 2406 12521 2474 12577
rect 2530 12521 2598 12577
rect 2654 12521 2722 12577
rect 2778 12521 2846 12577
rect 2902 12521 2970 12577
rect 3026 12521 3094 12577
rect 3150 12521 3218 12577
rect 3274 12521 3342 12577
rect 3398 12521 3466 12577
rect 3522 12521 3590 12577
rect 3646 12521 3714 12577
rect 3770 12521 3838 12577
rect 3894 12521 3962 12577
rect 4018 12521 4086 12577
rect 4142 12521 4210 12577
rect 4266 12521 4334 12577
rect 4390 12521 4458 12577
rect 4514 12521 4582 12577
rect 4638 12521 4706 12577
rect 4762 12521 4830 12577
rect 4886 12521 4954 12577
rect 5010 12521 5078 12577
rect 5134 12521 5202 12577
rect 5258 12521 5326 12577
rect 5382 12521 5450 12577
rect 5506 12521 5574 12577
rect 5630 12521 5698 12577
rect 5754 12521 5822 12577
rect 5878 12521 5946 12577
rect 6002 12521 6070 12577
rect 6126 12521 6194 12577
rect 6250 12521 6318 12577
rect 6374 12521 6442 12577
rect 6498 12521 6566 12577
rect 6622 12521 6690 12577
rect 6746 12521 6814 12577
rect 6870 12521 6938 12577
rect 6994 12521 7062 12577
rect 7118 12521 7186 12577
rect 7242 12521 7310 12577
rect 7366 12521 7434 12577
rect 7490 12521 7558 12577
rect 7614 12521 7682 12577
rect 7738 12521 7806 12577
rect 7862 12521 7930 12577
rect 7986 12521 8054 12577
rect 8110 12521 8178 12577
rect 8234 12521 8302 12577
rect 8358 12521 8426 12577
rect 8482 12521 8550 12577
rect 8606 12521 8674 12577
rect 8730 12521 8798 12577
rect 8854 12521 8922 12577
rect 8978 12521 9046 12577
rect 9102 12521 9170 12577
rect 9226 12521 9294 12577
rect 9350 12521 9418 12577
rect 9474 12521 9542 12577
rect 9598 12521 9666 12577
rect 9722 12521 9790 12577
rect 9846 12521 9914 12577
rect 9970 12521 10038 12577
rect 10094 12521 10162 12577
rect 10218 12521 10286 12577
rect 10342 12521 10410 12577
rect 10466 12521 10534 12577
rect 10590 12521 10658 12577
rect 10714 12521 10782 12577
rect 10838 12521 10906 12577
rect 10962 12521 11030 12577
rect 11086 12521 11154 12577
rect 11210 12521 11278 12577
rect 11334 12521 11402 12577
rect 11458 12521 11526 12577
rect 11582 12521 11650 12577
rect 11706 12521 11774 12577
rect 11830 12521 11898 12577
rect 11954 12521 12022 12577
rect 12078 12521 12146 12577
rect 12202 12521 12270 12577
rect 12326 12521 12394 12577
rect 12450 12521 12518 12577
rect 12574 12521 12642 12577
rect 12698 12521 12766 12577
rect 12822 12521 12890 12577
rect 12946 12521 13014 12577
rect 13070 12521 13200 12577
rect -400 12400 13200 12521
rect -400 12358 400 12400
rect -400 12302 -286 12358
rect -230 12302 -162 12358
rect -106 12302 -38 12358
rect 18 12302 86 12358
rect 142 12302 210 12358
rect 266 12302 400 12358
rect -400 12234 400 12302
rect -400 12178 -286 12234
rect -230 12178 -162 12234
rect -106 12178 -38 12234
rect 18 12178 86 12234
rect 142 12178 210 12234
rect 266 12178 400 12234
rect -400 12110 400 12178
rect -400 12054 -286 12110
rect -230 12054 -162 12110
rect -106 12054 -38 12110
rect 18 12054 86 12110
rect 142 12054 210 12110
rect 266 12054 400 12110
rect -400 11986 400 12054
rect -400 11930 -286 11986
rect -230 11930 -162 11986
rect -106 11930 -38 11986
rect 18 11930 86 11986
rect 142 11930 210 11986
rect 266 11930 400 11986
rect -400 11862 400 11930
rect -400 11806 -286 11862
rect -230 11806 -162 11862
rect -106 11806 -38 11862
rect 18 11806 86 11862
rect 142 11806 210 11862
rect 266 11806 400 11862
rect -400 11738 400 11806
rect -400 11682 -286 11738
rect -230 11682 -162 11738
rect -106 11682 -38 11738
rect 18 11682 86 11738
rect 142 11682 210 11738
rect 266 11682 400 11738
rect -400 11614 400 11682
rect -400 11558 -286 11614
rect -230 11558 -162 11614
rect -106 11558 -38 11614
rect 18 11558 86 11614
rect 142 11558 210 11614
rect 266 11558 400 11614
rect -400 11490 400 11558
rect -400 11434 -286 11490
rect -230 11434 -162 11490
rect -106 11434 -38 11490
rect 18 11434 86 11490
rect 142 11434 210 11490
rect 266 11434 400 11490
rect -400 11366 400 11434
rect -400 11310 -286 11366
rect -230 11310 -162 11366
rect -106 11310 -38 11366
rect 18 11310 86 11366
rect 142 11310 210 11366
rect 266 11310 400 11366
rect -400 11242 400 11310
rect -400 11186 -286 11242
rect -230 11186 -162 11242
rect -106 11186 -38 11242
rect 18 11186 86 11242
rect 142 11186 210 11242
rect 266 11186 400 11242
rect -400 11118 400 11186
rect -400 11062 -286 11118
rect -230 11062 -162 11118
rect -106 11062 -38 11118
rect 18 11062 86 11118
rect 142 11062 210 11118
rect 266 11062 400 11118
rect -400 10994 400 11062
rect -400 10938 -286 10994
rect -230 10938 -162 10994
rect -106 10938 -38 10994
rect 18 10938 86 10994
rect 142 10938 210 10994
rect 266 10938 400 10994
rect -400 10870 400 10938
rect -400 10814 -286 10870
rect -230 10814 -162 10870
rect -106 10814 -38 10870
rect 18 10814 86 10870
rect 142 10814 210 10870
rect 266 10814 400 10870
rect -400 10746 400 10814
rect -400 10690 -286 10746
rect -230 10690 -162 10746
rect -106 10690 -38 10746
rect 18 10690 86 10746
rect 142 10690 210 10746
rect 266 10690 400 10746
rect -400 10622 400 10690
rect -400 10566 -286 10622
rect -230 10566 -162 10622
rect -106 10566 -38 10622
rect 18 10566 86 10622
rect 142 10566 210 10622
rect 266 10566 400 10622
rect -400 10498 400 10566
rect -400 10442 -286 10498
rect -230 10442 -162 10498
rect -106 10442 -38 10498
rect 18 10442 86 10498
rect 142 10442 210 10498
rect 266 10442 400 10498
rect -400 10374 400 10442
rect -400 10318 -286 10374
rect -230 10318 -162 10374
rect -106 10318 -38 10374
rect 18 10318 86 10374
rect 142 10318 210 10374
rect 266 10318 400 10374
rect -400 10250 400 10318
rect -400 10194 -286 10250
rect -230 10194 -162 10250
rect -106 10194 -38 10250
rect 18 10194 86 10250
rect 142 10194 210 10250
rect 266 10194 400 10250
rect -400 10126 400 10194
rect -400 10070 -286 10126
rect -230 10070 -162 10126
rect -106 10070 -38 10126
rect 18 10070 86 10126
rect 142 10070 210 10126
rect 266 10070 400 10126
rect -400 10002 400 10070
rect -400 9946 -286 10002
rect -230 9946 -162 10002
rect -106 9946 -38 10002
rect 18 9946 86 10002
rect 142 9946 210 10002
rect 266 9946 400 10002
rect -400 9878 400 9946
rect -400 9822 -286 9878
rect -230 9822 -162 9878
rect -106 9822 -38 9878
rect 18 9822 86 9878
rect 142 9822 210 9878
rect 266 9822 400 9878
rect -400 9754 400 9822
rect -400 9698 -286 9754
rect -230 9698 -162 9754
rect -106 9698 -38 9754
rect 18 9698 86 9754
rect 142 9698 210 9754
rect 266 9698 400 9754
rect -400 9630 400 9698
rect -400 9574 -286 9630
rect -230 9574 -162 9630
rect -106 9574 -38 9630
rect 18 9574 86 9630
rect 142 9574 210 9630
rect 266 9574 400 9630
rect -400 9506 400 9574
rect -400 9450 -286 9506
rect -230 9450 -162 9506
rect -106 9450 -38 9506
rect 18 9450 86 9506
rect 142 9450 210 9506
rect 266 9450 400 9506
rect -400 9382 400 9450
rect -400 9326 -286 9382
rect -230 9326 -162 9382
rect -106 9326 -38 9382
rect 18 9326 86 9382
rect 142 9326 210 9382
rect 266 9326 400 9382
rect -400 9258 400 9326
rect -400 9202 -286 9258
rect -230 9202 -162 9258
rect -106 9202 -38 9258
rect 18 9202 86 9258
rect 142 9202 210 9258
rect 266 9202 400 9258
rect -400 9134 400 9202
rect -400 9078 -286 9134
rect -230 9078 -162 9134
rect -106 9078 -38 9134
rect 18 9078 86 9134
rect 142 9078 210 9134
rect 266 9078 400 9134
rect -400 9010 400 9078
rect -400 8954 -286 9010
rect -230 8954 -162 9010
rect -106 8954 -38 9010
rect 18 8954 86 9010
rect 142 8954 210 9010
rect 266 8954 400 9010
rect -400 8886 400 8954
rect -400 8830 -286 8886
rect -230 8830 -162 8886
rect -106 8830 -38 8886
rect 18 8830 86 8886
rect 142 8830 210 8886
rect 266 8830 400 8886
rect -400 8762 400 8830
rect -400 8706 -286 8762
rect -230 8706 -162 8762
rect -106 8706 -38 8762
rect 18 8706 86 8762
rect 142 8706 210 8762
rect 266 8706 400 8762
rect -400 8638 400 8706
rect -400 8582 -286 8638
rect -230 8582 -162 8638
rect -106 8582 -38 8638
rect 18 8582 86 8638
rect 142 8582 210 8638
rect 266 8582 400 8638
rect -400 8514 400 8582
rect -400 8458 -286 8514
rect -230 8458 -162 8514
rect -106 8458 -38 8514
rect 18 8458 86 8514
rect 142 8458 210 8514
rect 266 8458 400 8514
rect -400 8390 400 8458
rect -400 8334 -286 8390
rect -230 8334 -162 8390
rect -106 8334 -38 8390
rect 18 8334 86 8390
rect 142 8334 210 8390
rect 266 8334 400 8390
rect -400 8266 400 8334
rect -400 8210 -286 8266
rect -230 8210 -162 8266
rect -106 8210 -38 8266
rect 18 8210 86 8266
rect 142 8210 210 8266
rect 266 8210 400 8266
rect -400 8142 400 8210
rect -400 8086 -286 8142
rect -230 8086 -162 8142
rect -106 8086 -38 8142
rect 18 8086 86 8142
rect 142 8086 210 8142
rect 266 8086 400 8142
rect -400 8018 400 8086
rect -400 7962 -286 8018
rect -230 7962 -162 8018
rect -106 7962 -38 8018
rect 18 7962 86 8018
rect 142 7962 210 8018
rect 266 7962 400 8018
rect -400 7894 400 7962
rect -400 7838 -286 7894
rect -230 7838 -162 7894
rect -106 7838 -38 7894
rect 18 7838 86 7894
rect 142 7838 210 7894
rect 266 7838 400 7894
rect -400 7770 400 7838
rect -400 7714 -286 7770
rect -230 7714 -162 7770
rect -106 7714 -38 7770
rect 18 7714 86 7770
rect 142 7714 210 7770
rect 266 7714 400 7770
rect -400 7646 400 7714
rect -400 7590 -286 7646
rect -230 7590 -162 7646
rect -106 7590 -38 7646
rect 18 7590 86 7646
rect 142 7590 210 7646
rect 266 7590 400 7646
rect -400 7522 400 7590
rect -400 7466 -286 7522
rect -230 7466 -162 7522
rect -106 7466 -38 7522
rect 18 7466 86 7522
rect 142 7466 210 7522
rect 266 7466 400 7522
rect -400 7398 400 7466
rect -400 7342 -286 7398
rect -230 7342 -162 7398
rect -106 7342 -38 7398
rect 18 7342 86 7398
rect 142 7342 210 7398
rect 266 7342 400 7398
rect -400 7274 400 7342
rect -400 7218 -286 7274
rect -230 7218 -162 7274
rect -106 7218 -38 7274
rect 18 7218 86 7274
rect 142 7218 210 7274
rect 266 7218 400 7274
rect -400 7150 400 7218
rect -400 7094 -286 7150
rect -230 7094 -162 7150
rect -106 7094 -38 7150
rect 18 7094 86 7150
rect 142 7094 210 7150
rect 266 7094 400 7150
rect -400 7026 400 7094
rect -400 6970 -286 7026
rect -230 6970 -162 7026
rect -106 6970 -38 7026
rect 18 6970 86 7026
rect 142 6970 210 7026
rect 266 6970 400 7026
rect -400 6902 400 6970
rect -400 6846 -286 6902
rect -230 6846 -162 6902
rect -106 6846 -38 6902
rect 18 6846 86 6902
rect 142 6846 210 6902
rect 266 6846 400 6902
rect -400 6778 400 6846
rect -400 6722 -286 6778
rect -230 6722 -162 6778
rect -106 6722 -38 6778
rect 18 6722 86 6778
rect 142 6722 210 6778
rect 266 6722 400 6778
rect -400 6654 400 6722
rect -400 6598 -286 6654
rect -230 6598 -162 6654
rect -106 6598 -38 6654
rect 18 6598 86 6654
rect 142 6598 210 6654
rect 266 6598 400 6654
rect -400 6530 400 6598
rect -400 6474 -286 6530
rect -230 6474 -162 6530
rect -106 6474 -38 6530
rect 18 6474 86 6530
rect 142 6474 210 6530
rect 266 6474 400 6530
rect -400 6406 400 6474
rect -400 6350 -286 6406
rect -230 6350 -162 6406
rect -106 6350 -38 6406
rect 18 6350 86 6406
rect 142 6350 210 6406
rect 266 6350 400 6406
rect -400 6282 400 6350
rect -400 6226 -286 6282
rect -230 6226 -162 6282
rect -106 6226 -38 6282
rect 18 6226 86 6282
rect 142 6226 210 6282
rect 266 6226 400 6282
rect -400 6158 400 6226
rect -400 6102 -286 6158
rect -230 6102 -162 6158
rect -106 6102 -38 6158
rect 18 6102 86 6158
rect 142 6102 210 6158
rect 266 6102 400 6158
rect -400 6034 400 6102
rect -400 5978 -286 6034
rect -230 5978 -162 6034
rect -106 5978 -38 6034
rect 18 5978 86 6034
rect 142 5978 210 6034
rect 266 5978 400 6034
rect -400 5910 400 5978
rect -400 5854 -286 5910
rect -230 5854 -162 5910
rect -106 5854 -38 5910
rect 18 5854 86 5910
rect 142 5854 210 5910
rect 266 5854 400 5910
rect -400 5786 400 5854
rect -400 5730 -286 5786
rect -230 5730 -162 5786
rect -106 5730 -38 5786
rect 18 5730 86 5786
rect 142 5730 210 5786
rect 266 5730 400 5786
rect -400 5662 400 5730
rect -400 5606 -286 5662
rect -230 5606 -162 5662
rect -106 5606 -38 5662
rect 18 5606 86 5662
rect 142 5606 210 5662
rect 266 5606 400 5662
rect -400 5538 400 5606
rect -400 5482 -286 5538
rect -230 5482 -162 5538
rect -106 5482 -38 5538
rect 18 5482 86 5538
rect 142 5482 210 5538
rect 266 5482 400 5538
rect -400 5414 400 5482
rect -400 5358 -286 5414
rect -230 5358 -162 5414
rect -106 5358 -38 5414
rect 18 5358 86 5414
rect 142 5358 210 5414
rect 266 5358 400 5414
rect -400 5290 400 5358
rect -400 5234 -286 5290
rect -230 5234 -162 5290
rect -106 5234 -38 5290
rect 18 5234 86 5290
rect 142 5234 210 5290
rect 266 5234 400 5290
rect -400 5166 400 5234
rect -400 5110 -286 5166
rect -230 5110 -162 5166
rect -106 5110 -38 5166
rect 18 5110 86 5166
rect 142 5110 210 5166
rect 266 5110 400 5166
rect -400 5042 400 5110
rect -400 4986 -286 5042
rect -230 4986 -162 5042
rect -106 4986 -38 5042
rect 18 4986 86 5042
rect 142 4986 210 5042
rect 266 4986 400 5042
rect -400 4918 400 4986
rect -400 4862 -286 4918
rect -230 4862 -162 4918
rect -106 4862 -38 4918
rect 18 4862 86 4918
rect 142 4862 210 4918
rect 266 4862 400 4918
rect -400 4794 400 4862
rect -400 4738 -286 4794
rect -230 4738 -162 4794
rect -106 4738 -38 4794
rect 18 4738 86 4794
rect 142 4738 210 4794
rect 266 4738 400 4794
rect -400 4670 400 4738
rect -400 4614 -286 4670
rect -230 4614 -162 4670
rect -106 4614 -38 4670
rect 18 4614 86 4670
rect 142 4614 210 4670
rect 266 4614 400 4670
rect -400 4546 400 4614
rect -400 4490 -286 4546
rect -230 4490 -162 4546
rect -106 4490 -38 4546
rect 18 4490 86 4546
rect 142 4490 210 4546
rect 266 4490 400 4546
rect -400 4422 400 4490
rect -400 4366 -286 4422
rect -230 4366 -162 4422
rect -106 4366 -38 4422
rect 18 4366 86 4422
rect 142 4366 210 4422
rect 266 4366 400 4422
rect -400 4298 400 4366
rect -400 4242 -286 4298
rect -230 4242 -162 4298
rect -106 4242 -38 4298
rect 18 4242 86 4298
rect 142 4242 210 4298
rect 266 4242 400 4298
rect -400 4174 400 4242
rect -400 4118 -286 4174
rect -230 4118 -162 4174
rect -106 4118 -38 4174
rect 18 4118 86 4174
rect 142 4118 210 4174
rect 266 4118 400 4174
rect -400 4050 400 4118
rect -400 3994 -286 4050
rect -230 3994 -162 4050
rect -106 3994 -38 4050
rect 18 3994 86 4050
rect 142 3994 210 4050
rect 266 3994 400 4050
rect -400 3926 400 3994
rect -400 3870 -286 3926
rect -230 3870 -162 3926
rect -106 3870 -38 3926
rect 18 3870 86 3926
rect 142 3870 210 3926
rect 266 3870 400 3926
rect -400 3802 400 3870
rect -400 3746 -286 3802
rect -230 3746 -162 3802
rect -106 3746 -38 3802
rect 18 3746 86 3802
rect 142 3746 210 3802
rect 266 3746 400 3802
rect -400 3678 400 3746
rect -400 3622 -286 3678
rect -230 3622 -162 3678
rect -106 3622 -38 3678
rect 18 3622 86 3678
rect 142 3622 210 3678
rect 266 3622 400 3678
rect -400 3554 400 3622
rect -400 3498 -286 3554
rect -230 3498 -162 3554
rect -106 3498 -38 3554
rect 18 3498 86 3554
rect 142 3498 210 3554
rect 266 3498 400 3554
rect -400 3430 400 3498
rect -400 3374 -286 3430
rect -230 3374 -162 3430
rect -106 3374 -38 3430
rect 18 3374 86 3430
rect 142 3374 210 3430
rect 266 3374 400 3430
rect -400 3306 400 3374
rect -400 3250 -286 3306
rect -230 3250 -162 3306
rect -106 3250 -38 3306
rect 18 3250 86 3306
rect 142 3250 210 3306
rect 266 3250 400 3306
rect -400 3182 400 3250
rect -400 3126 -286 3182
rect -230 3126 -162 3182
rect -106 3126 -38 3182
rect 18 3126 86 3182
rect 142 3126 210 3182
rect 266 3126 400 3182
rect -400 3058 400 3126
rect -400 3002 -286 3058
rect -230 3002 -162 3058
rect -106 3002 -38 3058
rect 18 3002 86 3058
rect 142 3002 210 3058
rect 266 3002 400 3058
rect -400 2934 400 3002
rect -400 2878 -286 2934
rect -230 2878 -162 2934
rect -106 2878 -38 2934
rect 18 2878 86 2934
rect 142 2878 210 2934
rect 266 2878 400 2934
rect -400 2810 400 2878
rect -400 2754 -286 2810
rect -230 2754 -162 2810
rect -106 2754 -38 2810
rect 18 2754 86 2810
rect 142 2754 210 2810
rect 266 2754 400 2810
rect -400 2686 400 2754
rect -400 2630 -286 2686
rect -230 2630 -162 2686
rect -106 2630 -38 2686
rect 18 2630 86 2686
rect 142 2630 210 2686
rect 266 2630 400 2686
rect -400 2562 400 2630
rect -400 2506 -286 2562
rect -230 2506 -162 2562
rect -106 2506 -38 2562
rect 18 2506 86 2562
rect 142 2506 210 2562
rect 266 2506 400 2562
rect -400 2438 400 2506
rect -400 2382 -286 2438
rect -230 2382 -162 2438
rect -106 2382 -38 2438
rect 18 2382 86 2438
rect 142 2382 210 2438
rect 266 2382 400 2438
rect -400 2314 400 2382
rect -400 2258 -286 2314
rect -230 2258 -162 2314
rect -106 2258 -38 2314
rect 18 2258 86 2314
rect 142 2258 210 2314
rect 266 2258 400 2314
rect -400 2190 400 2258
rect -400 2134 -286 2190
rect -230 2134 -162 2190
rect -106 2134 -38 2190
rect 18 2134 86 2190
rect 142 2134 210 2190
rect 266 2134 400 2190
rect -400 2066 400 2134
rect -400 2010 -286 2066
rect -230 2010 -162 2066
rect -106 2010 -38 2066
rect 18 2010 86 2066
rect 142 2010 210 2066
rect 266 2010 400 2066
rect -400 1942 400 2010
rect -400 1886 -286 1942
rect -230 1886 -162 1942
rect -106 1886 -38 1942
rect 18 1886 86 1942
rect 142 1886 210 1942
rect 266 1886 400 1942
rect -400 1818 400 1886
rect -400 1762 -286 1818
rect -230 1762 -162 1818
rect -106 1762 -38 1818
rect 18 1762 86 1818
rect 142 1762 210 1818
rect 266 1762 400 1818
rect -400 1694 400 1762
rect -400 1638 -286 1694
rect -230 1638 -162 1694
rect -106 1638 -38 1694
rect 18 1638 86 1694
rect 142 1638 210 1694
rect 266 1638 400 1694
rect -400 1570 400 1638
rect -400 1514 -286 1570
rect -230 1514 -162 1570
rect -106 1514 -38 1570
rect 18 1514 86 1570
rect 142 1514 210 1570
rect 266 1514 400 1570
rect -400 1446 400 1514
rect -400 1390 -286 1446
rect -230 1390 -162 1446
rect -106 1390 -38 1446
rect 18 1390 86 1446
rect 142 1390 210 1446
rect 266 1390 400 1446
rect -400 1322 400 1390
rect -400 1266 -286 1322
rect -230 1266 -162 1322
rect -106 1266 -38 1322
rect 18 1266 86 1322
rect 142 1266 210 1322
rect 266 1266 400 1322
rect -400 1198 400 1266
rect -400 1142 -286 1198
rect -230 1142 -162 1198
rect -106 1142 -38 1198
rect 18 1142 86 1198
rect 142 1142 210 1198
rect 266 1142 400 1198
rect -400 1074 400 1142
rect -400 1018 -286 1074
rect -230 1018 -162 1074
rect -106 1018 -38 1074
rect 18 1018 86 1074
rect 142 1018 210 1074
rect 266 1018 400 1074
rect -400 950 400 1018
rect -400 894 -286 950
rect -230 894 -162 950
rect -106 894 -38 950
rect 18 894 86 950
rect 142 894 210 950
rect 266 894 400 950
rect -400 826 400 894
rect -400 770 -286 826
rect -230 770 -162 826
rect -106 770 -38 826
rect 18 770 86 826
rect 142 770 210 826
rect 266 770 400 826
rect -400 702 400 770
rect -400 646 -286 702
rect -230 646 -162 702
rect -106 646 -38 702
rect 18 646 86 702
rect 142 646 210 702
rect 266 646 400 702
rect -400 578 400 646
rect -400 522 -286 578
rect -230 522 -162 578
rect -106 522 -38 578
rect 18 522 86 578
rect 142 522 210 578
rect 266 522 400 578
rect -400 454 400 522
rect -400 398 -286 454
rect -230 398 -162 454
rect -106 398 -38 454
rect 18 398 86 454
rect 142 398 210 454
rect 266 400 400 454
rect 668 12310 1008 12400
rect 668 12254 741 12310
rect 797 12254 883 12310
rect 939 12254 1008 12310
rect 668 12168 1008 12254
rect 668 12112 741 12168
rect 797 12112 883 12168
rect 939 12112 1008 12168
rect 668 12026 1008 12112
rect 668 11970 741 12026
rect 797 11970 883 12026
rect 939 11970 1008 12026
rect 668 11884 1008 11970
rect 668 11828 741 11884
rect 797 11828 883 11884
rect 939 11828 1008 11884
rect 668 11742 1008 11828
rect 668 11686 741 11742
rect 797 11686 883 11742
rect 939 11686 1008 11742
rect 668 11600 1008 11686
rect 668 11544 741 11600
rect 797 11544 883 11600
rect 939 11544 1008 11600
rect 668 11458 1008 11544
rect 668 11402 741 11458
rect 797 11402 883 11458
rect 939 11402 1008 11458
rect 668 11316 1008 11402
rect 668 11260 741 11316
rect 797 11260 883 11316
rect 939 11260 1008 11316
rect 668 11174 1008 11260
rect 668 11118 741 11174
rect 797 11118 883 11174
rect 939 11118 1008 11174
rect 668 11032 1008 11118
rect 668 10976 741 11032
rect 797 10976 883 11032
rect 939 10976 1008 11032
rect 668 10890 1008 10976
rect 668 10834 741 10890
rect 797 10834 883 10890
rect 939 10834 1008 10890
rect 668 10748 1008 10834
rect 668 10692 741 10748
rect 797 10692 883 10748
rect 939 10692 1008 10748
rect 668 10606 1008 10692
rect 668 10550 741 10606
rect 797 10550 883 10606
rect 939 10550 1008 10606
rect 668 10464 1008 10550
rect 668 10408 741 10464
rect 797 10408 883 10464
rect 939 10408 1008 10464
rect 668 10322 1008 10408
rect 668 10266 741 10322
rect 797 10266 883 10322
rect 939 10266 1008 10322
rect 668 10180 1008 10266
rect 668 10124 741 10180
rect 797 10124 883 10180
rect 939 10124 1008 10180
rect 668 10038 1008 10124
rect 668 9982 741 10038
rect 797 9982 883 10038
rect 939 9982 1008 10038
rect 668 9896 1008 9982
rect 668 9840 741 9896
rect 797 9840 883 9896
rect 939 9840 1008 9896
rect 668 9754 1008 9840
rect 668 9698 741 9754
rect 797 9698 883 9754
rect 939 9698 1008 9754
rect 668 9612 1008 9698
rect 668 9556 741 9612
rect 797 9556 883 9612
rect 939 9556 1008 9612
rect 668 9470 1008 9556
rect 668 9414 741 9470
rect 797 9414 883 9470
rect 939 9414 1008 9470
rect 668 9328 1008 9414
rect 668 9272 741 9328
rect 797 9272 883 9328
rect 939 9272 1008 9328
rect 668 9186 1008 9272
rect 668 9130 741 9186
rect 797 9130 883 9186
rect 939 9130 1008 9186
rect 668 9044 1008 9130
rect 668 8988 741 9044
rect 797 8988 883 9044
rect 939 8988 1008 9044
rect 668 8902 1008 8988
rect 668 8846 741 8902
rect 797 8846 883 8902
rect 939 8846 1008 8902
rect 668 8760 1008 8846
rect 668 8704 741 8760
rect 797 8704 883 8760
rect 939 8704 1008 8760
rect 668 8618 1008 8704
rect 668 8562 741 8618
rect 797 8562 883 8618
rect 939 8562 1008 8618
rect 668 8476 1008 8562
rect 668 8420 741 8476
rect 797 8420 883 8476
rect 939 8420 1008 8476
rect 668 8334 1008 8420
rect 668 8278 741 8334
rect 797 8278 883 8334
rect 939 8278 1008 8334
rect 668 8192 1008 8278
rect 668 8136 741 8192
rect 797 8136 883 8192
rect 939 8136 1008 8192
rect 668 8050 1008 8136
rect 668 7994 741 8050
rect 797 7994 883 8050
rect 939 7994 1008 8050
rect 668 7908 1008 7994
rect 668 7852 741 7908
rect 797 7852 883 7908
rect 939 7852 1008 7908
rect 668 7766 1008 7852
rect 668 7710 741 7766
rect 797 7710 883 7766
rect 939 7710 1008 7766
rect 668 7624 1008 7710
rect 668 7568 741 7624
rect 797 7568 883 7624
rect 939 7568 1008 7624
rect 668 7482 1008 7568
rect 668 7426 741 7482
rect 797 7426 883 7482
rect 939 7426 1008 7482
rect 668 7340 1008 7426
rect 668 7284 741 7340
rect 797 7284 883 7340
rect 939 7284 1008 7340
rect 668 7198 1008 7284
rect 668 7142 741 7198
rect 797 7142 883 7198
rect 939 7142 1008 7198
rect 668 7056 1008 7142
rect 668 7000 741 7056
rect 797 7000 883 7056
rect 939 7000 1008 7056
rect 668 6914 1008 7000
rect 668 6858 741 6914
rect 797 6858 883 6914
rect 939 6858 1008 6914
rect 668 6772 1008 6858
rect 668 6716 741 6772
rect 797 6716 883 6772
rect 939 6716 1008 6772
rect 668 6630 1008 6716
rect 668 6574 741 6630
rect 797 6574 883 6630
rect 939 6574 1008 6630
rect 668 6488 1008 6574
rect 668 6432 741 6488
rect 797 6432 883 6488
rect 939 6432 1008 6488
rect 668 6346 1008 6432
rect 668 6290 741 6346
rect 797 6290 883 6346
rect 939 6290 1008 6346
rect 668 6204 1008 6290
rect 668 6148 741 6204
rect 797 6148 883 6204
rect 939 6148 1008 6204
rect 668 6062 1008 6148
rect 668 6006 741 6062
rect 797 6006 883 6062
rect 939 6006 1008 6062
rect 668 5920 1008 6006
rect 668 5864 741 5920
rect 797 5864 883 5920
rect 939 5864 1008 5920
rect 668 5778 1008 5864
rect 668 5722 741 5778
rect 797 5722 883 5778
rect 939 5722 1008 5778
rect 668 5636 1008 5722
rect 668 5580 741 5636
rect 797 5580 883 5636
rect 939 5580 1008 5636
rect 668 5494 1008 5580
rect 668 5438 741 5494
rect 797 5438 883 5494
rect 939 5438 1008 5494
rect 668 5352 1008 5438
rect 668 5296 741 5352
rect 797 5296 883 5352
rect 939 5296 1008 5352
rect 668 5210 1008 5296
rect 668 5154 741 5210
rect 797 5154 883 5210
rect 939 5154 1008 5210
rect 668 5068 1008 5154
rect 668 5012 741 5068
rect 797 5012 883 5068
rect 939 5012 1008 5068
rect 668 4926 1008 5012
rect 668 4870 741 4926
rect 797 4870 883 4926
rect 939 4870 1008 4926
rect 668 4784 1008 4870
rect 668 4728 741 4784
rect 797 4728 883 4784
rect 939 4728 1008 4784
rect 668 4642 1008 4728
rect 668 4586 741 4642
rect 797 4586 883 4642
rect 939 4586 1008 4642
rect 668 4500 1008 4586
rect 668 4444 741 4500
rect 797 4444 883 4500
rect 939 4444 1008 4500
rect 668 4358 1008 4444
rect 668 4302 741 4358
rect 797 4302 883 4358
rect 939 4302 1008 4358
rect 668 4216 1008 4302
rect 668 4160 741 4216
rect 797 4160 883 4216
rect 939 4160 1008 4216
rect 668 4074 1008 4160
rect 668 4018 741 4074
rect 797 4018 883 4074
rect 939 4018 1008 4074
rect 668 3932 1008 4018
rect 668 3876 741 3932
rect 797 3876 883 3932
rect 939 3876 1008 3932
rect 668 3790 1008 3876
rect 668 3734 741 3790
rect 797 3734 883 3790
rect 939 3734 1008 3790
rect 668 3648 1008 3734
rect 668 3592 741 3648
rect 797 3592 883 3648
rect 939 3592 1008 3648
rect 668 3506 1008 3592
rect 668 3450 741 3506
rect 797 3450 883 3506
rect 939 3450 1008 3506
rect 668 3364 1008 3450
rect 668 3308 741 3364
rect 797 3308 883 3364
rect 939 3308 1008 3364
rect 668 3222 1008 3308
rect 668 3166 741 3222
rect 797 3166 883 3222
rect 939 3166 1008 3222
rect 668 3080 1008 3166
rect 668 3024 741 3080
rect 797 3024 883 3080
rect 939 3024 1008 3080
rect 668 2938 1008 3024
rect 668 2882 741 2938
rect 797 2882 883 2938
rect 939 2882 1008 2938
rect 668 2796 1008 2882
rect 668 2740 741 2796
rect 797 2740 883 2796
rect 939 2740 1008 2796
rect 668 2654 1008 2740
rect 668 2598 741 2654
rect 797 2598 883 2654
rect 939 2598 1008 2654
rect 668 2512 1008 2598
rect 668 2456 741 2512
rect 797 2456 883 2512
rect 939 2456 1008 2512
rect 668 2370 1008 2456
rect 668 2314 741 2370
rect 797 2314 883 2370
rect 939 2314 1008 2370
rect 668 2228 1008 2314
rect 668 2172 741 2228
rect 797 2172 883 2228
rect 939 2172 1008 2228
rect 668 2086 1008 2172
rect 668 2030 741 2086
rect 797 2030 883 2086
rect 939 2030 1008 2086
rect 668 1944 1008 2030
rect 668 1888 741 1944
rect 797 1888 883 1944
rect 939 1888 1008 1944
rect 668 1802 1008 1888
rect 668 1746 741 1802
rect 797 1746 883 1802
rect 939 1746 1008 1802
rect 668 1660 1008 1746
rect 668 1604 741 1660
rect 797 1604 883 1660
rect 939 1604 1008 1660
rect 668 1518 1008 1604
rect 668 1462 741 1518
rect 797 1462 883 1518
rect 939 1462 1008 1518
rect 668 1376 1008 1462
rect 668 1320 741 1376
rect 797 1320 883 1376
rect 939 1320 1008 1376
rect 668 1234 1008 1320
rect 668 1178 741 1234
rect 797 1178 883 1234
rect 939 1178 1008 1234
rect 668 1092 1008 1178
rect 668 1036 741 1092
rect 797 1036 883 1092
rect 939 1036 1008 1092
rect 668 950 1008 1036
rect 668 894 741 950
rect 797 894 883 950
rect 939 894 1008 950
rect 668 808 1008 894
rect 668 752 741 808
rect 797 752 883 808
rect 939 752 1008 808
rect 668 666 1008 752
rect 668 610 741 666
rect 797 610 883 666
rect 939 610 1008 666
rect 668 524 1008 610
rect 668 468 741 524
rect 797 468 883 524
rect 939 468 1008 524
rect 668 400 1008 468
rect 1068 12310 1408 12400
rect 1068 12254 1142 12310
rect 1198 12254 1284 12310
rect 1340 12254 1408 12310
rect 1068 12168 1408 12254
rect 1068 12112 1142 12168
rect 1198 12112 1284 12168
rect 1340 12112 1408 12168
rect 1068 12026 1408 12112
rect 1068 11970 1142 12026
rect 1198 11970 1284 12026
rect 1340 11970 1408 12026
rect 1068 11884 1408 11970
rect 1068 11828 1142 11884
rect 1198 11828 1284 11884
rect 1340 11828 1408 11884
rect 1068 11742 1408 11828
rect 1068 11686 1142 11742
rect 1198 11686 1284 11742
rect 1340 11686 1408 11742
rect 1068 11600 1408 11686
rect 1068 11544 1142 11600
rect 1198 11544 1284 11600
rect 1340 11544 1408 11600
rect 1068 11458 1408 11544
rect 1068 11402 1142 11458
rect 1198 11402 1284 11458
rect 1340 11402 1408 11458
rect 1068 11316 1408 11402
rect 1068 11260 1142 11316
rect 1198 11260 1284 11316
rect 1340 11260 1408 11316
rect 1068 11174 1408 11260
rect 1068 11118 1142 11174
rect 1198 11118 1284 11174
rect 1340 11118 1408 11174
rect 1068 11032 1408 11118
rect 1068 10976 1142 11032
rect 1198 10976 1284 11032
rect 1340 10976 1408 11032
rect 1068 10890 1408 10976
rect 1068 10834 1142 10890
rect 1198 10834 1284 10890
rect 1340 10834 1408 10890
rect 1068 10748 1408 10834
rect 1068 10692 1142 10748
rect 1198 10692 1284 10748
rect 1340 10692 1408 10748
rect 1068 10606 1408 10692
rect 1068 10550 1142 10606
rect 1198 10550 1284 10606
rect 1340 10550 1408 10606
rect 1068 10464 1408 10550
rect 1068 10408 1142 10464
rect 1198 10408 1284 10464
rect 1340 10408 1408 10464
rect 1068 10322 1408 10408
rect 1068 10266 1142 10322
rect 1198 10266 1284 10322
rect 1340 10266 1408 10322
rect 1068 10180 1408 10266
rect 1068 10124 1142 10180
rect 1198 10124 1284 10180
rect 1340 10124 1408 10180
rect 1068 10038 1408 10124
rect 1068 9982 1142 10038
rect 1198 9982 1284 10038
rect 1340 9982 1408 10038
rect 1068 9896 1408 9982
rect 1068 9840 1142 9896
rect 1198 9840 1284 9896
rect 1340 9840 1408 9896
rect 1068 9754 1408 9840
rect 1068 9698 1142 9754
rect 1198 9698 1284 9754
rect 1340 9698 1408 9754
rect 1068 9612 1408 9698
rect 1068 9556 1142 9612
rect 1198 9556 1284 9612
rect 1340 9556 1408 9612
rect 1068 9470 1408 9556
rect 1068 9414 1142 9470
rect 1198 9414 1284 9470
rect 1340 9414 1408 9470
rect 1068 9328 1408 9414
rect 1068 9272 1142 9328
rect 1198 9272 1284 9328
rect 1340 9272 1408 9328
rect 1068 9186 1408 9272
rect 1068 9130 1142 9186
rect 1198 9130 1284 9186
rect 1340 9130 1408 9186
rect 1068 9044 1408 9130
rect 1068 8988 1142 9044
rect 1198 8988 1284 9044
rect 1340 8988 1408 9044
rect 1068 8902 1408 8988
rect 1068 8846 1142 8902
rect 1198 8846 1284 8902
rect 1340 8846 1408 8902
rect 1068 8760 1408 8846
rect 1068 8704 1142 8760
rect 1198 8704 1284 8760
rect 1340 8704 1408 8760
rect 1068 8618 1408 8704
rect 1068 8562 1142 8618
rect 1198 8562 1284 8618
rect 1340 8562 1408 8618
rect 1068 8476 1408 8562
rect 1068 8420 1142 8476
rect 1198 8420 1284 8476
rect 1340 8420 1408 8476
rect 1068 8334 1408 8420
rect 1068 8278 1142 8334
rect 1198 8278 1284 8334
rect 1340 8278 1408 8334
rect 1068 8192 1408 8278
rect 1068 8136 1142 8192
rect 1198 8136 1284 8192
rect 1340 8136 1408 8192
rect 1068 8050 1408 8136
rect 1068 7994 1142 8050
rect 1198 7994 1284 8050
rect 1340 7994 1408 8050
rect 1068 7908 1408 7994
rect 1068 7852 1142 7908
rect 1198 7852 1284 7908
rect 1340 7852 1408 7908
rect 1068 7766 1408 7852
rect 1068 7710 1142 7766
rect 1198 7710 1284 7766
rect 1340 7710 1408 7766
rect 1068 7624 1408 7710
rect 1068 7568 1142 7624
rect 1198 7568 1284 7624
rect 1340 7568 1408 7624
rect 1068 7482 1408 7568
rect 1068 7426 1142 7482
rect 1198 7426 1284 7482
rect 1340 7426 1408 7482
rect 1068 7340 1408 7426
rect 1068 7284 1142 7340
rect 1198 7284 1284 7340
rect 1340 7284 1408 7340
rect 1068 7198 1408 7284
rect 1068 7142 1142 7198
rect 1198 7142 1284 7198
rect 1340 7142 1408 7198
rect 1068 7056 1408 7142
rect 1068 7000 1142 7056
rect 1198 7000 1284 7056
rect 1340 7000 1408 7056
rect 1068 6914 1408 7000
rect 1068 6858 1142 6914
rect 1198 6858 1284 6914
rect 1340 6858 1408 6914
rect 1068 6772 1408 6858
rect 1068 6716 1142 6772
rect 1198 6716 1284 6772
rect 1340 6716 1408 6772
rect 1068 6630 1408 6716
rect 1068 6574 1142 6630
rect 1198 6574 1284 6630
rect 1340 6574 1408 6630
rect 1068 6488 1408 6574
rect 1068 6432 1142 6488
rect 1198 6432 1284 6488
rect 1340 6432 1408 6488
rect 1068 6346 1408 6432
rect 1068 6290 1142 6346
rect 1198 6290 1284 6346
rect 1340 6290 1408 6346
rect 1068 6204 1408 6290
rect 1068 6148 1142 6204
rect 1198 6148 1284 6204
rect 1340 6148 1408 6204
rect 1068 6062 1408 6148
rect 1068 6006 1142 6062
rect 1198 6006 1284 6062
rect 1340 6006 1408 6062
rect 1068 5920 1408 6006
rect 1068 5864 1142 5920
rect 1198 5864 1284 5920
rect 1340 5864 1408 5920
rect 1068 5778 1408 5864
rect 1068 5722 1142 5778
rect 1198 5722 1284 5778
rect 1340 5722 1408 5778
rect 1068 5636 1408 5722
rect 1068 5580 1142 5636
rect 1198 5580 1284 5636
rect 1340 5580 1408 5636
rect 1068 5494 1408 5580
rect 1068 5438 1142 5494
rect 1198 5438 1284 5494
rect 1340 5438 1408 5494
rect 1068 5352 1408 5438
rect 1068 5296 1142 5352
rect 1198 5296 1284 5352
rect 1340 5296 1408 5352
rect 1068 5210 1408 5296
rect 1068 5154 1142 5210
rect 1198 5154 1284 5210
rect 1340 5154 1408 5210
rect 1068 5068 1408 5154
rect 1068 5012 1142 5068
rect 1198 5012 1284 5068
rect 1340 5012 1408 5068
rect 1068 4926 1408 5012
rect 1068 4870 1142 4926
rect 1198 4870 1284 4926
rect 1340 4870 1408 4926
rect 1068 4784 1408 4870
rect 1068 4728 1142 4784
rect 1198 4728 1284 4784
rect 1340 4728 1408 4784
rect 1068 4642 1408 4728
rect 1068 4586 1142 4642
rect 1198 4586 1284 4642
rect 1340 4586 1408 4642
rect 1068 4500 1408 4586
rect 1068 4444 1142 4500
rect 1198 4444 1284 4500
rect 1340 4444 1408 4500
rect 1068 4358 1408 4444
rect 1068 4302 1142 4358
rect 1198 4302 1284 4358
rect 1340 4302 1408 4358
rect 1068 4216 1408 4302
rect 1068 4160 1142 4216
rect 1198 4160 1284 4216
rect 1340 4160 1408 4216
rect 1068 4074 1408 4160
rect 1068 4018 1142 4074
rect 1198 4018 1284 4074
rect 1340 4018 1408 4074
rect 1068 3932 1408 4018
rect 1068 3876 1142 3932
rect 1198 3876 1284 3932
rect 1340 3876 1408 3932
rect 1068 3790 1408 3876
rect 1068 3734 1142 3790
rect 1198 3734 1284 3790
rect 1340 3734 1408 3790
rect 1068 3648 1408 3734
rect 1068 3592 1142 3648
rect 1198 3592 1284 3648
rect 1340 3592 1408 3648
rect 1068 3506 1408 3592
rect 1068 3450 1142 3506
rect 1198 3450 1284 3506
rect 1340 3450 1408 3506
rect 1068 3364 1408 3450
rect 1068 3308 1142 3364
rect 1198 3308 1284 3364
rect 1340 3308 1408 3364
rect 1068 3222 1408 3308
rect 1068 3166 1142 3222
rect 1198 3166 1284 3222
rect 1340 3166 1408 3222
rect 1068 3080 1408 3166
rect 1068 3024 1142 3080
rect 1198 3024 1284 3080
rect 1340 3024 1408 3080
rect 1068 2938 1408 3024
rect 1068 2882 1142 2938
rect 1198 2882 1284 2938
rect 1340 2882 1408 2938
rect 1068 2796 1408 2882
rect 1068 2740 1142 2796
rect 1198 2740 1284 2796
rect 1340 2740 1408 2796
rect 1068 2654 1408 2740
rect 1068 2598 1142 2654
rect 1198 2598 1284 2654
rect 1340 2598 1408 2654
rect 1068 2512 1408 2598
rect 1068 2456 1142 2512
rect 1198 2456 1284 2512
rect 1340 2456 1408 2512
rect 1068 2370 1408 2456
rect 1068 2314 1142 2370
rect 1198 2314 1284 2370
rect 1340 2314 1408 2370
rect 1068 2228 1408 2314
rect 1068 2172 1142 2228
rect 1198 2172 1284 2228
rect 1340 2172 1408 2228
rect 1068 2086 1408 2172
rect 1068 2030 1142 2086
rect 1198 2030 1284 2086
rect 1340 2030 1408 2086
rect 1068 1944 1408 2030
rect 1068 1888 1142 1944
rect 1198 1888 1284 1944
rect 1340 1888 1408 1944
rect 1068 1802 1408 1888
rect 1068 1746 1142 1802
rect 1198 1746 1284 1802
rect 1340 1746 1408 1802
rect 1068 1660 1408 1746
rect 1068 1604 1142 1660
rect 1198 1604 1284 1660
rect 1340 1604 1408 1660
rect 1068 1518 1408 1604
rect 1068 1462 1142 1518
rect 1198 1462 1284 1518
rect 1340 1462 1408 1518
rect 1068 1376 1408 1462
rect 1068 1320 1142 1376
rect 1198 1320 1284 1376
rect 1340 1320 1408 1376
rect 1068 1234 1408 1320
rect 1068 1178 1142 1234
rect 1198 1178 1284 1234
rect 1340 1178 1408 1234
rect 1068 1092 1408 1178
rect 1068 1036 1142 1092
rect 1198 1036 1284 1092
rect 1340 1036 1408 1092
rect 1068 950 1408 1036
rect 1068 894 1142 950
rect 1198 894 1284 950
rect 1340 894 1408 950
rect 1068 808 1408 894
rect 1068 752 1142 808
rect 1198 752 1284 808
rect 1340 752 1408 808
rect 1068 666 1408 752
rect 1068 610 1142 666
rect 1198 610 1284 666
rect 1340 610 1408 666
rect 1068 524 1408 610
rect 1068 468 1142 524
rect 1198 468 1284 524
rect 1340 468 1408 524
rect 1068 400 1408 468
rect 1468 12310 1808 12400
rect 1468 12254 1542 12310
rect 1598 12254 1684 12310
rect 1740 12254 1808 12310
rect 1468 12168 1808 12254
rect 1468 12112 1542 12168
rect 1598 12112 1684 12168
rect 1740 12112 1808 12168
rect 1468 12026 1808 12112
rect 1468 11970 1542 12026
rect 1598 11970 1684 12026
rect 1740 11970 1808 12026
rect 1468 11884 1808 11970
rect 1468 11828 1542 11884
rect 1598 11828 1684 11884
rect 1740 11828 1808 11884
rect 1468 11742 1808 11828
rect 1468 11686 1542 11742
rect 1598 11686 1684 11742
rect 1740 11686 1808 11742
rect 1468 11600 1808 11686
rect 1468 11544 1542 11600
rect 1598 11544 1684 11600
rect 1740 11544 1808 11600
rect 1468 11458 1808 11544
rect 1468 11402 1542 11458
rect 1598 11402 1684 11458
rect 1740 11402 1808 11458
rect 1468 11316 1808 11402
rect 1468 11260 1542 11316
rect 1598 11260 1684 11316
rect 1740 11260 1808 11316
rect 1468 11174 1808 11260
rect 1468 11118 1542 11174
rect 1598 11118 1684 11174
rect 1740 11118 1808 11174
rect 1468 11032 1808 11118
rect 1468 10976 1542 11032
rect 1598 10976 1684 11032
rect 1740 10976 1808 11032
rect 1468 10890 1808 10976
rect 1468 10834 1542 10890
rect 1598 10834 1684 10890
rect 1740 10834 1808 10890
rect 1468 10748 1808 10834
rect 1468 10692 1542 10748
rect 1598 10692 1684 10748
rect 1740 10692 1808 10748
rect 1468 10606 1808 10692
rect 1468 10550 1542 10606
rect 1598 10550 1684 10606
rect 1740 10550 1808 10606
rect 1468 10464 1808 10550
rect 1468 10408 1542 10464
rect 1598 10408 1684 10464
rect 1740 10408 1808 10464
rect 1468 10322 1808 10408
rect 1468 10266 1542 10322
rect 1598 10266 1684 10322
rect 1740 10266 1808 10322
rect 1468 10180 1808 10266
rect 1468 10124 1542 10180
rect 1598 10124 1684 10180
rect 1740 10124 1808 10180
rect 1468 10038 1808 10124
rect 1468 9982 1542 10038
rect 1598 9982 1684 10038
rect 1740 9982 1808 10038
rect 1468 9896 1808 9982
rect 1468 9840 1542 9896
rect 1598 9840 1684 9896
rect 1740 9840 1808 9896
rect 1468 9754 1808 9840
rect 1468 9698 1542 9754
rect 1598 9698 1684 9754
rect 1740 9698 1808 9754
rect 1468 9612 1808 9698
rect 1468 9556 1542 9612
rect 1598 9556 1684 9612
rect 1740 9556 1808 9612
rect 1468 9470 1808 9556
rect 1468 9414 1542 9470
rect 1598 9414 1684 9470
rect 1740 9414 1808 9470
rect 1468 9328 1808 9414
rect 1468 9272 1542 9328
rect 1598 9272 1684 9328
rect 1740 9272 1808 9328
rect 1468 9186 1808 9272
rect 1468 9130 1542 9186
rect 1598 9130 1684 9186
rect 1740 9130 1808 9186
rect 1468 9044 1808 9130
rect 1468 8988 1542 9044
rect 1598 8988 1684 9044
rect 1740 8988 1808 9044
rect 1468 8902 1808 8988
rect 1468 8846 1542 8902
rect 1598 8846 1684 8902
rect 1740 8846 1808 8902
rect 1468 8760 1808 8846
rect 1468 8704 1542 8760
rect 1598 8704 1684 8760
rect 1740 8704 1808 8760
rect 1468 8618 1808 8704
rect 1468 8562 1542 8618
rect 1598 8562 1684 8618
rect 1740 8562 1808 8618
rect 1468 8476 1808 8562
rect 1468 8420 1542 8476
rect 1598 8420 1684 8476
rect 1740 8420 1808 8476
rect 1468 8334 1808 8420
rect 1468 8278 1542 8334
rect 1598 8278 1684 8334
rect 1740 8278 1808 8334
rect 1468 8192 1808 8278
rect 1468 8136 1542 8192
rect 1598 8136 1684 8192
rect 1740 8136 1808 8192
rect 1468 8050 1808 8136
rect 1468 7994 1542 8050
rect 1598 7994 1684 8050
rect 1740 7994 1808 8050
rect 1468 7908 1808 7994
rect 1468 7852 1542 7908
rect 1598 7852 1684 7908
rect 1740 7852 1808 7908
rect 1468 7766 1808 7852
rect 1468 7710 1542 7766
rect 1598 7710 1684 7766
rect 1740 7710 1808 7766
rect 1468 7624 1808 7710
rect 1468 7568 1542 7624
rect 1598 7568 1684 7624
rect 1740 7568 1808 7624
rect 1468 7482 1808 7568
rect 1468 7426 1542 7482
rect 1598 7426 1684 7482
rect 1740 7426 1808 7482
rect 1468 7340 1808 7426
rect 1468 7284 1542 7340
rect 1598 7284 1684 7340
rect 1740 7284 1808 7340
rect 1468 7198 1808 7284
rect 1468 7142 1542 7198
rect 1598 7142 1684 7198
rect 1740 7142 1808 7198
rect 1468 7056 1808 7142
rect 1468 7000 1542 7056
rect 1598 7000 1684 7056
rect 1740 7000 1808 7056
rect 1468 6914 1808 7000
rect 1468 6858 1542 6914
rect 1598 6858 1684 6914
rect 1740 6858 1808 6914
rect 1468 6772 1808 6858
rect 1468 6716 1542 6772
rect 1598 6716 1684 6772
rect 1740 6716 1808 6772
rect 1468 6630 1808 6716
rect 1468 6574 1542 6630
rect 1598 6574 1684 6630
rect 1740 6574 1808 6630
rect 1468 6488 1808 6574
rect 1468 6432 1542 6488
rect 1598 6432 1684 6488
rect 1740 6432 1808 6488
rect 1468 6346 1808 6432
rect 1468 6290 1542 6346
rect 1598 6290 1684 6346
rect 1740 6290 1808 6346
rect 1468 6204 1808 6290
rect 1468 6148 1542 6204
rect 1598 6148 1684 6204
rect 1740 6148 1808 6204
rect 1468 6062 1808 6148
rect 1468 6006 1542 6062
rect 1598 6006 1684 6062
rect 1740 6006 1808 6062
rect 1468 5920 1808 6006
rect 1468 5864 1542 5920
rect 1598 5864 1684 5920
rect 1740 5864 1808 5920
rect 1468 5778 1808 5864
rect 1468 5722 1542 5778
rect 1598 5722 1684 5778
rect 1740 5722 1808 5778
rect 1468 5636 1808 5722
rect 1468 5580 1542 5636
rect 1598 5580 1684 5636
rect 1740 5580 1808 5636
rect 1468 5494 1808 5580
rect 1468 5438 1542 5494
rect 1598 5438 1684 5494
rect 1740 5438 1808 5494
rect 1468 5352 1808 5438
rect 1468 5296 1542 5352
rect 1598 5296 1684 5352
rect 1740 5296 1808 5352
rect 1468 5210 1808 5296
rect 1468 5154 1542 5210
rect 1598 5154 1684 5210
rect 1740 5154 1808 5210
rect 1468 5068 1808 5154
rect 1468 5012 1542 5068
rect 1598 5012 1684 5068
rect 1740 5012 1808 5068
rect 1468 4926 1808 5012
rect 1468 4870 1542 4926
rect 1598 4870 1684 4926
rect 1740 4870 1808 4926
rect 1468 4784 1808 4870
rect 1468 4728 1542 4784
rect 1598 4728 1684 4784
rect 1740 4728 1808 4784
rect 1468 4642 1808 4728
rect 1468 4586 1542 4642
rect 1598 4586 1684 4642
rect 1740 4586 1808 4642
rect 1468 4500 1808 4586
rect 1468 4444 1542 4500
rect 1598 4444 1684 4500
rect 1740 4444 1808 4500
rect 1468 4358 1808 4444
rect 1468 4302 1542 4358
rect 1598 4302 1684 4358
rect 1740 4302 1808 4358
rect 1468 4216 1808 4302
rect 1468 4160 1542 4216
rect 1598 4160 1684 4216
rect 1740 4160 1808 4216
rect 1468 4074 1808 4160
rect 1468 4018 1542 4074
rect 1598 4018 1684 4074
rect 1740 4018 1808 4074
rect 1468 3932 1808 4018
rect 1468 3876 1542 3932
rect 1598 3876 1684 3932
rect 1740 3876 1808 3932
rect 1468 3790 1808 3876
rect 1468 3734 1542 3790
rect 1598 3734 1684 3790
rect 1740 3734 1808 3790
rect 1468 3648 1808 3734
rect 1468 3592 1542 3648
rect 1598 3592 1684 3648
rect 1740 3592 1808 3648
rect 1468 3506 1808 3592
rect 1468 3450 1542 3506
rect 1598 3450 1684 3506
rect 1740 3450 1808 3506
rect 1468 3364 1808 3450
rect 1468 3308 1542 3364
rect 1598 3308 1684 3364
rect 1740 3308 1808 3364
rect 1468 3222 1808 3308
rect 1468 3166 1542 3222
rect 1598 3166 1684 3222
rect 1740 3166 1808 3222
rect 1468 3080 1808 3166
rect 1468 3024 1542 3080
rect 1598 3024 1684 3080
rect 1740 3024 1808 3080
rect 1468 2938 1808 3024
rect 1468 2882 1542 2938
rect 1598 2882 1684 2938
rect 1740 2882 1808 2938
rect 1468 2796 1808 2882
rect 1468 2740 1542 2796
rect 1598 2740 1684 2796
rect 1740 2740 1808 2796
rect 1468 2654 1808 2740
rect 1468 2598 1542 2654
rect 1598 2598 1684 2654
rect 1740 2598 1808 2654
rect 1468 2512 1808 2598
rect 1468 2456 1542 2512
rect 1598 2456 1684 2512
rect 1740 2456 1808 2512
rect 1468 2370 1808 2456
rect 1468 2314 1542 2370
rect 1598 2314 1684 2370
rect 1740 2314 1808 2370
rect 1468 2228 1808 2314
rect 1468 2172 1542 2228
rect 1598 2172 1684 2228
rect 1740 2172 1808 2228
rect 1468 2086 1808 2172
rect 1468 2030 1542 2086
rect 1598 2030 1684 2086
rect 1740 2030 1808 2086
rect 1468 1944 1808 2030
rect 1468 1888 1542 1944
rect 1598 1888 1684 1944
rect 1740 1888 1808 1944
rect 1468 1802 1808 1888
rect 1468 1746 1542 1802
rect 1598 1746 1684 1802
rect 1740 1746 1808 1802
rect 1468 1660 1808 1746
rect 1468 1604 1542 1660
rect 1598 1604 1684 1660
rect 1740 1604 1808 1660
rect 1468 1518 1808 1604
rect 1468 1462 1542 1518
rect 1598 1462 1684 1518
rect 1740 1462 1808 1518
rect 1468 1376 1808 1462
rect 1468 1320 1542 1376
rect 1598 1320 1684 1376
rect 1740 1320 1808 1376
rect 1468 1234 1808 1320
rect 1468 1178 1542 1234
rect 1598 1178 1684 1234
rect 1740 1178 1808 1234
rect 1468 1092 1808 1178
rect 1468 1036 1542 1092
rect 1598 1036 1684 1092
rect 1740 1036 1808 1092
rect 1468 950 1808 1036
rect 1468 894 1542 950
rect 1598 894 1684 950
rect 1740 894 1808 950
rect 1468 808 1808 894
rect 1468 752 1542 808
rect 1598 752 1684 808
rect 1740 752 1808 808
rect 1468 666 1808 752
rect 1468 610 1542 666
rect 1598 610 1684 666
rect 1740 610 1808 666
rect 1468 524 1808 610
rect 1468 468 1542 524
rect 1598 468 1684 524
rect 1740 468 1808 524
rect 1468 400 1808 468
rect 1868 12310 2208 12400
rect 1868 12254 1939 12310
rect 1995 12254 2081 12310
rect 2137 12254 2208 12310
rect 1868 12168 2208 12254
rect 1868 12112 1939 12168
rect 1995 12112 2081 12168
rect 2137 12112 2208 12168
rect 1868 12026 2208 12112
rect 1868 11970 1939 12026
rect 1995 11970 2081 12026
rect 2137 11970 2208 12026
rect 1868 11884 2208 11970
rect 1868 11828 1939 11884
rect 1995 11828 2081 11884
rect 2137 11828 2208 11884
rect 1868 11742 2208 11828
rect 1868 11686 1939 11742
rect 1995 11686 2081 11742
rect 2137 11686 2208 11742
rect 1868 11600 2208 11686
rect 1868 11544 1939 11600
rect 1995 11544 2081 11600
rect 2137 11544 2208 11600
rect 1868 11458 2208 11544
rect 1868 11402 1939 11458
rect 1995 11402 2081 11458
rect 2137 11402 2208 11458
rect 1868 11316 2208 11402
rect 1868 11260 1939 11316
rect 1995 11260 2081 11316
rect 2137 11260 2208 11316
rect 1868 11174 2208 11260
rect 1868 11118 1939 11174
rect 1995 11118 2081 11174
rect 2137 11118 2208 11174
rect 1868 11032 2208 11118
rect 1868 10976 1939 11032
rect 1995 10976 2081 11032
rect 2137 10976 2208 11032
rect 1868 10890 2208 10976
rect 1868 10834 1939 10890
rect 1995 10834 2081 10890
rect 2137 10834 2208 10890
rect 1868 10748 2208 10834
rect 1868 10692 1939 10748
rect 1995 10692 2081 10748
rect 2137 10692 2208 10748
rect 1868 10606 2208 10692
rect 1868 10550 1939 10606
rect 1995 10550 2081 10606
rect 2137 10550 2208 10606
rect 1868 10464 2208 10550
rect 1868 10408 1939 10464
rect 1995 10408 2081 10464
rect 2137 10408 2208 10464
rect 1868 10322 2208 10408
rect 1868 10266 1939 10322
rect 1995 10266 2081 10322
rect 2137 10266 2208 10322
rect 1868 10180 2208 10266
rect 1868 10124 1939 10180
rect 1995 10124 2081 10180
rect 2137 10124 2208 10180
rect 1868 10038 2208 10124
rect 1868 9982 1939 10038
rect 1995 9982 2081 10038
rect 2137 9982 2208 10038
rect 1868 9896 2208 9982
rect 1868 9840 1939 9896
rect 1995 9840 2081 9896
rect 2137 9840 2208 9896
rect 1868 9754 2208 9840
rect 1868 9698 1939 9754
rect 1995 9698 2081 9754
rect 2137 9698 2208 9754
rect 1868 9612 2208 9698
rect 1868 9556 1939 9612
rect 1995 9556 2081 9612
rect 2137 9556 2208 9612
rect 1868 9470 2208 9556
rect 1868 9414 1939 9470
rect 1995 9414 2081 9470
rect 2137 9414 2208 9470
rect 1868 9328 2208 9414
rect 1868 9272 1939 9328
rect 1995 9272 2081 9328
rect 2137 9272 2208 9328
rect 1868 9186 2208 9272
rect 1868 9130 1939 9186
rect 1995 9130 2081 9186
rect 2137 9130 2208 9186
rect 1868 9044 2208 9130
rect 1868 8988 1939 9044
rect 1995 8988 2081 9044
rect 2137 8988 2208 9044
rect 1868 8902 2208 8988
rect 1868 8846 1939 8902
rect 1995 8846 2081 8902
rect 2137 8846 2208 8902
rect 1868 8760 2208 8846
rect 1868 8704 1939 8760
rect 1995 8704 2081 8760
rect 2137 8704 2208 8760
rect 1868 8618 2208 8704
rect 1868 8562 1939 8618
rect 1995 8562 2081 8618
rect 2137 8562 2208 8618
rect 1868 8476 2208 8562
rect 1868 8420 1939 8476
rect 1995 8420 2081 8476
rect 2137 8420 2208 8476
rect 1868 8334 2208 8420
rect 1868 8278 1939 8334
rect 1995 8278 2081 8334
rect 2137 8278 2208 8334
rect 1868 8192 2208 8278
rect 1868 8136 1939 8192
rect 1995 8136 2081 8192
rect 2137 8136 2208 8192
rect 1868 8050 2208 8136
rect 1868 7994 1939 8050
rect 1995 7994 2081 8050
rect 2137 7994 2208 8050
rect 1868 7908 2208 7994
rect 1868 7852 1939 7908
rect 1995 7852 2081 7908
rect 2137 7852 2208 7908
rect 1868 7766 2208 7852
rect 1868 7710 1939 7766
rect 1995 7710 2081 7766
rect 2137 7710 2208 7766
rect 1868 7624 2208 7710
rect 1868 7568 1939 7624
rect 1995 7568 2081 7624
rect 2137 7568 2208 7624
rect 1868 7482 2208 7568
rect 1868 7426 1939 7482
rect 1995 7426 2081 7482
rect 2137 7426 2208 7482
rect 1868 7340 2208 7426
rect 1868 7284 1939 7340
rect 1995 7284 2081 7340
rect 2137 7284 2208 7340
rect 1868 7198 2208 7284
rect 1868 7142 1939 7198
rect 1995 7142 2081 7198
rect 2137 7142 2208 7198
rect 1868 7056 2208 7142
rect 1868 7000 1939 7056
rect 1995 7000 2081 7056
rect 2137 7000 2208 7056
rect 1868 6914 2208 7000
rect 1868 6858 1939 6914
rect 1995 6858 2081 6914
rect 2137 6858 2208 6914
rect 1868 6772 2208 6858
rect 1868 6716 1939 6772
rect 1995 6716 2081 6772
rect 2137 6716 2208 6772
rect 1868 6630 2208 6716
rect 1868 6574 1939 6630
rect 1995 6574 2081 6630
rect 2137 6574 2208 6630
rect 1868 6488 2208 6574
rect 1868 6432 1939 6488
rect 1995 6432 2081 6488
rect 2137 6432 2208 6488
rect 1868 6346 2208 6432
rect 1868 6290 1939 6346
rect 1995 6290 2081 6346
rect 2137 6290 2208 6346
rect 1868 6204 2208 6290
rect 1868 6148 1939 6204
rect 1995 6148 2081 6204
rect 2137 6148 2208 6204
rect 1868 6062 2208 6148
rect 1868 6006 1939 6062
rect 1995 6006 2081 6062
rect 2137 6006 2208 6062
rect 1868 5920 2208 6006
rect 1868 5864 1939 5920
rect 1995 5864 2081 5920
rect 2137 5864 2208 5920
rect 1868 5778 2208 5864
rect 1868 5722 1939 5778
rect 1995 5722 2081 5778
rect 2137 5722 2208 5778
rect 1868 5636 2208 5722
rect 1868 5580 1939 5636
rect 1995 5580 2081 5636
rect 2137 5580 2208 5636
rect 1868 5494 2208 5580
rect 1868 5438 1939 5494
rect 1995 5438 2081 5494
rect 2137 5438 2208 5494
rect 1868 5352 2208 5438
rect 1868 5296 1939 5352
rect 1995 5296 2081 5352
rect 2137 5296 2208 5352
rect 1868 5210 2208 5296
rect 1868 5154 1939 5210
rect 1995 5154 2081 5210
rect 2137 5154 2208 5210
rect 1868 5068 2208 5154
rect 1868 5012 1939 5068
rect 1995 5012 2081 5068
rect 2137 5012 2208 5068
rect 1868 4926 2208 5012
rect 1868 4870 1939 4926
rect 1995 4870 2081 4926
rect 2137 4870 2208 4926
rect 1868 4784 2208 4870
rect 1868 4728 1939 4784
rect 1995 4728 2081 4784
rect 2137 4728 2208 4784
rect 1868 4642 2208 4728
rect 1868 4586 1939 4642
rect 1995 4586 2081 4642
rect 2137 4586 2208 4642
rect 1868 4500 2208 4586
rect 1868 4444 1939 4500
rect 1995 4444 2081 4500
rect 2137 4444 2208 4500
rect 1868 4358 2208 4444
rect 1868 4302 1939 4358
rect 1995 4302 2081 4358
rect 2137 4302 2208 4358
rect 1868 4216 2208 4302
rect 1868 4160 1939 4216
rect 1995 4160 2081 4216
rect 2137 4160 2208 4216
rect 1868 4074 2208 4160
rect 1868 4018 1939 4074
rect 1995 4018 2081 4074
rect 2137 4018 2208 4074
rect 1868 3932 2208 4018
rect 1868 3876 1939 3932
rect 1995 3876 2081 3932
rect 2137 3876 2208 3932
rect 1868 3790 2208 3876
rect 1868 3734 1939 3790
rect 1995 3734 2081 3790
rect 2137 3734 2208 3790
rect 1868 3648 2208 3734
rect 1868 3592 1939 3648
rect 1995 3592 2081 3648
rect 2137 3592 2208 3648
rect 1868 3506 2208 3592
rect 1868 3450 1939 3506
rect 1995 3450 2081 3506
rect 2137 3450 2208 3506
rect 1868 3364 2208 3450
rect 1868 3308 1939 3364
rect 1995 3308 2081 3364
rect 2137 3308 2208 3364
rect 1868 3222 2208 3308
rect 1868 3166 1939 3222
rect 1995 3166 2081 3222
rect 2137 3166 2208 3222
rect 1868 3080 2208 3166
rect 1868 3024 1939 3080
rect 1995 3024 2081 3080
rect 2137 3024 2208 3080
rect 1868 2938 2208 3024
rect 1868 2882 1939 2938
rect 1995 2882 2081 2938
rect 2137 2882 2208 2938
rect 1868 2796 2208 2882
rect 1868 2740 1939 2796
rect 1995 2740 2081 2796
rect 2137 2740 2208 2796
rect 1868 2654 2208 2740
rect 1868 2598 1939 2654
rect 1995 2598 2081 2654
rect 2137 2598 2208 2654
rect 1868 2512 2208 2598
rect 1868 2456 1939 2512
rect 1995 2456 2081 2512
rect 2137 2456 2208 2512
rect 1868 2370 2208 2456
rect 1868 2314 1939 2370
rect 1995 2314 2081 2370
rect 2137 2314 2208 2370
rect 1868 2228 2208 2314
rect 1868 2172 1939 2228
rect 1995 2172 2081 2228
rect 2137 2172 2208 2228
rect 1868 2086 2208 2172
rect 1868 2030 1939 2086
rect 1995 2030 2081 2086
rect 2137 2030 2208 2086
rect 1868 1944 2208 2030
rect 1868 1888 1939 1944
rect 1995 1888 2081 1944
rect 2137 1888 2208 1944
rect 1868 1802 2208 1888
rect 1868 1746 1939 1802
rect 1995 1746 2081 1802
rect 2137 1746 2208 1802
rect 1868 1660 2208 1746
rect 1868 1604 1939 1660
rect 1995 1604 2081 1660
rect 2137 1604 2208 1660
rect 1868 1518 2208 1604
rect 1868 1462 1939 1518
rect 1995 1462 2081 1518
rect 2137 1462 2208 1518
rect 1868 1376 2208 1462
rect 1868 1320 1939 1376
rect 1995 1320 2081 1376
rect 2137 1320 2208 1376
rect 1868 1234 2208 1320
rect 1868 1178 1939 1234
rect 1995 1178 2081 1234
rect 2137 1178 2208 1234
rect 1868 1092 2208 1178
rect 1868 1036 1939 1092
rect 1995 1036 2081 1092
rect 2137 1036 2208 1092
rect 1868 950 2208 1036
rect 1868 894 1939 950
rect 1995 894 2081 950
rect 2137 894 2208 950
rect 1868 808 2208 894
rect 1868 752 1939 808
rect 1995 752 2081 808
rect 2137 752 2208 808
rect 1868 666 2208 752
rect 1868 610 1939 666
rect 1995 610 2081 666
rect 2137 610 2208 666
rect 1868 524 2208 610
rect 1868 468 1939 524
rect 1995 468 2081 524
rect 2137 468 2208 524
rect 1868 400 2208 468
rect 2268 12310 2608 12400
rect 2268 12254 2336 12310
rect 2392 12254 2478 12310
rect 2534 12254 2608 12310
rect 2268 12168 2608 12254
rect 2268 12112 2336 12168
rect 2392 12112 2478 12168
rect 2534 12112 2608 12168
rect 2268 12026 2608 12112
rect 2268 11970 2336 12026
rect 2392 11970 2478 12026
rect 2534 11970 2608 12026
rect 2268 11884 2608 11970
rect 2268 11828 2336 11884
rect 2392 11828 2478 11884
rect 2534 11828 2608 11884
rect 2268 11742 2608 11828
rect 2268 11686 2336 11742
rect 2392 11686 2478 11742
rect 2534 11686 2608 11742
rect 2268 11600 2608 11686
rect 2268 11544 2336 11600
rect 2392 11544 2478 11600
rect 2534 11544 2608 11600
rect 2268 11458 2608 11544
rect 2268 11402 2336 11458
rect 2392 11402 2478 11458
rect 2534 11402 2608 11458
rect 2268 11316 2608 11402
rect 2268 11260 2336 11316
rect 2392 11260 2478 11316
rect 2534 11260 2608 11316
rect 2268 11174 2608 11260
rect 2268 11118 2336 11174
rect 2392 11118 2478 11174
rect 2534 11118 2608 11174
rect 2268 11032 2608 11118
rect 2268 10976 2336 11032
rect 2392 10976 2478 11032
rect 2534 10976 2608 11032
rect 2268 10890 2608 10976
rect 2268 10834 2336 10890
rect 2392 10834 2478 10890
rect 2534 10834 2608 10890
rect 2268 10748 2608 10834
rect 2268 10692 2336 10748
rect 2392 10692 2478 10748
rect 2534 10692 2608 10748
rect 2268 10606 2608 10692
rect 2268 10550 2336 10606
rect 2392 10550 2478 10606
rect 2534 10550 2608 10606
rect 2268 10464 2608 10550
rect 2268 10408 2336 10464
rect 2392 10408 2478 10464
rect 2534 10408 2608 10464
rect 2268 10322 2608 10408
rect 2268 10266 2336 10322
rect 2392 10266 2478 10322
rect 2534 10266 2608 10322
rect 2268 10180 2608 10266
rect 2268 10124 2336 10180
rect 2392 10124 2478 10180
rect 2534 10124 2608 10180
rect 2268 10038 2608 10124
rect 2268 9982 2336 10038
rect 2392 9982 2478 10038
rect 2534 9982 2608 10038
rect 2268 9896 2608 9982
rect 2268 9840 2336 9896
rect 2392 9840 2478 9896
rect 2534 9840 2608 9896
rect 2268 9754 2608 9840
rect 2268 9698 2336 9754
rect 2392 9698 2478 9754
rect 2534 9698 2608 9754
rect 2268 9612 2608 9698
rect 2268 9556 2336 9612
rect 2392 9556 2478 9612
rect 2534 9556 2608 9612
rect 2268 9470 2608 9556
rect 2268 9414 2336 9470
rect 2392 9414 2478 9470
rect 2534 9414 2608 9470
rect 2268 9328 2608 9414
rect 2268 9272 2336 9328
rect 2392 9272 2478 9328
rect 2534 9272 2608 9328
rect 2268 9186 2608 9272
rect 2268 9130 2336 9186
rect 2392 9130 2478 9186
rect 2534 9130 2608 9186
rect 2268 9044 2608 9130
rect 2268 8988 2336 9044
rect 2392 8988 2478 9044
rect 2534 8988 2608 9044
rect 2268 8902 2608 8988
rect 2268 8846 2336 8902
rect 2392 8846 2478 8902
rect 2534 8846 2608 8902
rect 2268 8760 2608 8846
rect 2268 8704 2336 8760
rect 2392 8704 2478 8760
rect 2534 8704 2608 8760
rect 2268 8618 2608 8704
rect 2268 8562 2336 8618
rect 2392 8562 2478 8618
rect 2534 8562 2608 8618
rect 2268 8476 2608 8562
rect 2268 8420 2336 8476
rect 2392 8420 2478 8476
rect 2534 8420 2608 8476
rect 2268 8334 2608 8420
rect 2268 8278 2336 8334
rect 2392 8278 2478 8334
rect 2534 8278 2608 8334
rect 2268 8192 2608 8278
rect 2268 8136 2336 8192
rect 2392 8136 2478 8192
rect 2534 8136 2608 8192
rect 2268 8050 2608 8136
rect 2268 7994 2336 8050
rect 2392 7994 2478 8050
rect 2534 7994 2608 8050
rect 2268 7908 2608 7994
rect 2268 7852 2336 7908
rect 2392 7852 2478 7908
rect 2534 7852 2608 7908
rect 2268 7766 2608 7852
rect 2268 7710 2336 7766
rect 2392 7710 2478 7766
rect 2534 7710 2608 7766
rect 2268 7624 2608 7710
rect 2268 7568 2336 7624
rect 2392 7568 2478 7624
rect 2534 7568 2608 7624
rect 2268 7482 2608 7568
rect 2268 7426 2336 7482
rect 2392 7426 2478 7482
rect 2534 7426 2608 7482
rect 2268 7340 2608 7426
rect 2268 7284 2336 7340
rect 2392 7284 2478 7340
rect 2534 7284 2608 7340
rect 2268 7198 2608 7284
rect 2268 7142 2336 7198
rect 2392 7142 2478 7198
rect 2534 7142 2608 7198
rect 2268 7056 2608 7142
rect 2268 7000 2336 7056
rect 2392 7000 2478 7056
rect 2534 7000 2608 7056
rect 2268 6914 2608 7000
rect 2268 6858 2336 6914
rect 2392 6858 2478 6914
rect 2534 6858 2608 6914
rect 2268 6772 2608 6858
rect 2268 6716 2336 6772
rect 2392 6716 2478 6772
rect 2534 6716 2608 6772
rect 2268 6630 2608 6716
rect 2268 6574 2336 6630
rect 2392 6574 2478 6630
rect 2534 6574 2608 6630
rect 2268 6488 2608 6574
rect 2268 6432 2336 6488
rect 2392 6432 2478 6488
rect 2534 6432 2608 6488
rect 2268 6346 2608 6432
rect 2268 6290 2336 6346
rect 2392 6290 2478 6346
rect 2534 6290 2608 6346
rect 2268 6204 2608 6290
rect 2268 6148 2336 6204
rect 2392 6148 2478 6204
rect 2534 6148 2608 6204
rect 2268 6062 2608 6148
rect 2268 6006 2336 6062
rect 2392 6006 2478 6062
rect 2534 6006 2608 6062
rect 2268 5920 2608 6006
rect 2268 5864 2336 5920
rect 2392 5864 2478 5920
rect 2534 5864 2608 5920
rect 2268 5778 2608 5864
rect 2268 5722 2336 5778
rect 2392 5722 2478 5778
rect 2534 5722 2608 5778
rect 2268 5636 2608 5722
rect 2268 5580 2336 5636
rect 2392 5580 2478 5636
rect 2534 5580 2608 5636
rect 2268 5494 2608 5580
rect 2268 5438 2336 5494
rect 2392 5438 2478 5494
rect 2534 5438 2608 5494
rect 2268 5352 2608 5438
rect 2268 5296 2336 5352
rect 2392 5296 2478 5352
rect 2534 5296 2608 5352
rect 2268 5210 2608 5296
rect 2268 5154 2336 5210
rect 2392 5154 2478 5210
rect 2534 5154 2608 5210
rect 2268 5068 2608 5154
rect 2268 5012 2336 5068
rect 2392 5012 2478 5068
rect 2534 5012 2608 5068
rect 2268 4926 2608 5012
rect 2268 4870 2336 4926
rect 2392 4870 2478 4926
rect 2534 4870 2608 4926
rect 2268 4784 2608 4870
rect 2268 4728 2336 4784
rect 2392 4728 2478 4784
rect 2534 4728 2608 4784
rect 2268 4642 2608 4728
rect 2268 4586 2336 4642
rect 2392 4586 2478 4642
rect 2534 4586 2608 4642
rect 2268 4500 2608 4586
rect 2268 4444 2336 4500
rect 2392 4444 2478 4500
rect 2534 4444 2608 4500
rect 2268 4358 2608 4444
rect 2268 4302 2336 4358
rect 2392 4302 2478 4358
rect 2534 4302 2608 4358
rect 2268 4216 2608 4302
rect 2268 4160 2336 4216
rect 2392 4160 2478 4216
rect 2534 4160 2608 4216
rect 2268 4074 2608 4160
rect 2268 4018 2336 4074
rect 2392 4018 2478 4074
rect 2534 4018 2608 4074
rect 2268 3932 2608 4018
rect 2268 3876 2336 3932
rect 2392 3876 2478 3932
rect 2534 3876 2608 3932
rect 2268 3790 2608 3876
rect 2268 3734 2336 3790
rect 2392 3734 2478 3790
rect 2534 3734 2608 3790
rect 2268 3648 2608 3734
rect 2268 3592 2336 3648
rect 2392 3592 2478 3648
rect 2534 3592 2608 3648
rect 2268 3506 2608 3592
rect 2268 3450 2336 3506
rect 2392 3450 2478 3506
rect 2534 3450 2608 3506
rect 2268 3364 2608 3450
rect 2268 3308 2336 3364
rect 2392 3308 2478 3364
rect 2534 3308 2608 3364
rect 2268 3222 2608 3308
rect 2268 3166 2336 3222
rect 2392 3166 2478 3222
rect 2534 3166 2608 3222
rect 2268 3080 2608 3166
rect 2268 3024 2336 3080
rect 2392 3024 2478 3080
rect 2534 3024 2608 3080
rect 2268 2938 2608 3024
rect 2268 2882 2336 2938
rect 2392 2882 2478 2938
rect 2534 2882 2608 2938
rect 2268 2796 2608 2882
rect 2268 2740 2336 2796
rect 2392 2740 2478 2796
rect 2534 2740 2608 2796
rect 2268 2654 2608 2740
rect 2268 2598 2336 2654
rect 2392 2598 2478 2654
rect 2534 2598 2608 2654
rect 2268 2512 2608 2598
rect 2268 2456 2336 2512
rect 2392 2456 2478 2512
rect 2534 2456 2608 2512
rect 2268 2370 2608 2456
rect 2268 2314 2336 2370
rect 2392 2314 2478 2370
rect 2534 2314 2608 2370
rect 2268 2228 2608 2314
rect 2268 2172 2336 2228
rect 2392 2172 2478 2228
rect 2534 2172 2608 2228
rect 2268 2086 2608 2172
rect 2268 2030 2336 2086
rect 2392 2030 2478 2086
rect 2534 2030 2608 2086
rect 2268 1944 2608 2030
rect 2268 1888 2336 1944
rect 2392 1888 2478 1944
rect 2534 1888 2608 1944
rect 2268 1802 2608 1888
rect 2268 1746 2336 1802
rect 2392 1746 2478 1802
rect 2534 1746 2608 1802
rect 2268 1660 2608 1746
rect 2268 1604 2336 1660
rect 2392 1604 2478 1660
rect 2534 1604 2608 1660
rect 2268 1518 2608 1604
rect 2268 1462 2336 1518
rect 2392 1462 2478 1518
rect 2534 1462 2608 1518
rect 2268 1376 2608 1462
rect 2268 1320 2336 1376
rect 2392 1320 2478 1376
rect 2534 1320 2608 1376
rect 2268 1234 2608 1320
rect 2268 1178 2336 1234
rect 2392 1178 2478 1234
rect 2534 1178 2608 1234
rect 2268 1092 2608 1178
rect 2268 1036 2336 1092
rect 2392 1036 2478 1092
rect 2534 1036 2608 1092
rect 2268 950 2608 1036
rect 2268 894 2336 950
rect 2392 894 2478 950
rect 2534 894 2608 950
rect 2268 808 2608 894
rect 2268 752 2336 808
rect 2392 752 2478 808
rect 2534 752 2608 808
rect 2268 666 2608 752
rect 2268 610 2336 666
rect 2392 610 2478 666
rect 2534 610 2608 666
rect 2268 524 2608 610
rect 2268 468 2336 524
rect 2392 468 2478 524
rect 2534 468 2608 524
rect 2268 400 2608 468
rect 2668 12310 3008 12400
rect 2668 12254 2740 12310
rect 2796 12254 2882 12310
rect 2938 12254 3008 12310
rect 2668 12168 3008 12254
rect 2668 12112 2740 12168
rect 2796 12112 2882 12168
rect 2938 12112 3008 12168
rect 2668 12026 3008 12112
rect 2668 11970 2740 12026
rect 2796 11970 2882 12026
rect 2938 11970 3008 12026
rect 2668 11884 3008 11970
rect 2668 11828 2740 11884
rect 2796 11828 2882 11884
rect 2938 11828 3008 11884
rect 2668 11742 3008 11828
rect 2668 11686 2740 11742
rect 2796 11686 2882 11742
rect 2938 11686 3008 11742
rect 2668 11600 3008 11686
rect 2668 11544 2740 11600
rect 2796 11544 2882 11600
rect 2938 11544 3008 11600
rect 2668 11458 3008 11544
rect 2668 11402 2740 11458
rect 2796 11402 2882 11458
rect 2938 11402 3008 11458
rect 2668 11316 3008 11402
rect 2668 11260 2740 11316
rect 2796 11260 2882 11316
rect 2938 11260 3008 11316
rect 2668 11174 3008 11260
rect 2668 11118 2740 11174
rect 2796 11118 2882 11174
rect 2938 11118 3008 11174
rect 2668 11032 3008 11118
rect 2668 10976 2740 11032
rect 2796 10976 2882 11032
rect 2938 10976 3008 11032
rect 2668 10890 3008 10976
rect 2668 10834 2740 10890
rect 2796 10834 2882 10890
rect 2938 10834 3008 10890
rect 2668 10748 3008 10834
rect 2668 10692 2740 10748
rect 2796 10692 2882 10748
rect 2938 10692 3008 10748
rect 2668 10606 3008 10692
rect 2668 10550 2740 10606
rect 2796 10550 2882 10606
rect 2938 10550 3008 10606
rect 2668 10464 3008 10550
rect 2668 10408 2740 10464
rect 2796 10408 2882 10464
rect 2938 10408 3008 10464
rect 2668 10322 3008 10408
rect 2668 10266 2740 10322
rect 2796 10266 2882 10322
rect 2938 10266 3008 10322
rect 2668 10180 3008 10266
rect 2668 10124 2740 10180
rect 2796 10124 2882 10180
rect 2938 10124 3008 10180
rect 2668 10038 3008 10124
rect 2668 9982 2740 10038
rect 2796 9982 2882 10038
rect 2938 9982 3008 10038
rect 2668 9896 3008 9982
rect 2668 9840 2740 9896
rect 2796 9840 2882 9896
rect 2938 9840 3008 9896
rect 2668 9754 3008 9840
rect 2668 9698 2740 9754
rect 2796 9698 2882 9754
rect 2938 9698 3008 9754
rect 2668 9612 3008 9698
rect 2668 9556 2740 9612
rect 2796 9556 2882 9612
rect 2938 9556 3008 9612
rect 2668 9470 3008 9556
rect 2668 9414 2740 9470
rect 2796 9414 2882 9470
rect 2938 9414 3008 9470
rect 2668 9328 3008 9414
rect 2668 9272 2740 9328
rect 2796 9272 2882 9328
rect 2938 9272 3008 9328
rect 2668 9186 3008 9272
rect 2668 9130 2740 9186
rect 2796 9130 2882 9186
rect 2938 9130 3008 9186
rect 2668 9044 3008 9130
rect 2668 8988 2740 9044
rect 2796 8988 2882 9044
rect 2938 8988 3008 9044
rect 2668 8902 3008 8988
rect 2668 8846 2740 8902
rect 2796 8846 2882 8902
rect 2938 8846 3008 8902
rect 2668 8760 3008 8846
rect 2668 8704 2740 8760
rect 2796 8704 2882 8760
rect 2938 8704 3008 8760
rect 2668 8618 3008 8704
rect 2668 8562 2740 8618
rect 2796 8562 2882 8618
rect 2938 8562 3008 8618
rect 2668 8476 3008 8562
rect 2668 8420 2740 8476
rect 2796 8420 2882 8476
rect 2938 8420 3008 8476
rect 2668 8334 3008 8420
rect 2668 8278 2740 8334
rect 2796 8278 2882 8334
rect 2938 8278 3008 8334
rect 2668 8192 3008 8278
rect 2668 8136 2740 8192
rect 2796 8136 2882 8192
rect 2938 8136 3008 8192
rect 2668 8050 3008 8136
rect 2668 7994 2740 8050
rect 2796 7994 2882 8050
rect 2938 7994 3008 8050
rect 2668 7908 3008 7994
rect 2668 7852 2740 7908
rect 2796 7852 2882 7908
rect 2938 7852 3008 7908
rect 2668 7766 3008 7852
rect 2668 7710 2740 7766
rect 2796 7710 2882 7766
rect 2938 7710 3008 7766
rect 2668 7624 3008 7710
rect 2668 7568 2740 7624
rect 2796 7568 2882 7624
rect 2938 7568 3008 7624
rect 2668 7482 3008 7568
rect 2668 7426 2740 7482
rect 2796 7426 2882 7482
rect 2938 7426 3008 7482
rect 2668 7340 3008 7426
rect 2668 7284 2740 7340
rect 2796 7284 2882 7340
rect 2938 7284 3008 7340
rect 2668 7198 3008 7284
rect 2668 7142 2740 7198
rect 2796 7142 2882 7198
rect 2938 7142 3008 7198
rect 2668 7056 3008 7142
rect 2668 7000 2740 7056
rect 2796 7000 2882 7056
rect 2938 7000 3008 7056
rect 2668 6914 3008 7000
rect 2668 6858 2740 6914
rect 2796 6858 2882 6914
rect 2938 6858 3008 6914
rect 2668 6772 3008 6858
rect 2668 6716 2740 6772
rect 2796 6716 2882 6772
rect 2938 6716 3008 6772
rect 2668 6630 3008 6716
rect 2668 6574 2740 6630
rect 2796 6574 2882 6630
rect 2938 6574 3008 6630
rect 2668 6488 3008 6574
rect 2668 6432 2740 6488
rect 2796 6432 2882 6488
rect 2938 6432 3008 6488
rect 2668 6346 3008 6432
rect 2668 6290 2740 6346
rect 2796 6290 2882 6346
rect 2938 6290 3008 6346
rect 2668 6204 3008 6290
rect 2668 6148 2740 6204
rect 2796 6148 2882 6204
rect 2938 6148 3008 6204
rect 2668 6062 3008 6148
rect 2668 6006 2740 6062
rect 2796 6006 2882 6062
rect 2938 6006 3008 6062
rect 2668 5920 3008 6006
rect 2668 5864 2740 5920
rect 2796 5864 2882 5920
rect 2938 5864 3008 5920
rect 2668 5778 3008 5864
rect 2668 5722 2740 5778
rect 2796 5722 2882 5778
rect 2938 5722 3008 5778
rect 2668 5636 3008 5722
rect 2668 5580 2740 5636
rect 2796 5580 2882 5636
rect 2938 5580 3008 5636
rect 2668 5494 3008 5580
rect 2668 5438 2740 5494
rect 2796 5438 2882 5494
rect 2938 5438 3008 5494
rect 2668 5352 3008 5438
rect 2668 5296 2740 5352
rect 2796 5296 2882 5352
rect 2938 5296 3008 5352
rect 2668 5210 3008 5296
rect 2668 5154 2740 5210
rect 2796 5154 2882 5210
rect 2938 5154 3008 5210
rect 2668 5068 3008 5154
rect 2668 5012 2740 5068
rect 2796 5012 2882 5068
rect 2938 5012 3008 5068
rect 2668 4926 3008 5012
rect 2668 4870 2740 4926
rect 2796 4870 2882 4926
rect 2938 4870 3008 4926
rect 2668 4784 3008 4870
rect 2668 4728 2740 4784
rect 2796 4728 2882 4784
rect 2938 4728 3008 4784
rect 2668 4642 3008 4728
rect 2668 4586 2740 4642
rect 2796 4586 2882 4642
rect 2938 4586 3008 4642
rect 2668 4500 3008 4586
rect 2668 4444 2740 4500
rect 2796 4444 2882 4500
rect 2938 4444 3008 4500
rect 2668 4358 3008 4444
rect 2668 4302 2740 4358
rect 2796 4302 2882 4358
rect 2938 4302 3008 4358
rect 2668 4216 3008 4302
rect 2668 4160 2740 4216
rect 2796 4160 2882 4216
rect 2938 4160 3008 4216
rect 2668 4074 3008 4160
rect 2668 4018 2740 4074
rect 2796 4018 2882 4074
rect 2938 4018 3008 4074
rect 2668 3932 3008 4018
rect 2668 3876 2740 3932
rect 2796 3876 2882 3932
rect 2938 3876 3008 3932
rect 2668 3790 3008 3876
rect 2668 3734 2740 3790
rect 2796 3734 2882 3790
rect 2938 3734 3008 3790
rect 2668 3648 3008 3734
rect 2668 3592 2740 3648
rect 2796 3592 2882 3648
rect 2938 3592 3008 3648
rect 2668 3506 3008 3592
rect 2668 3450 2740 3506
rect 2796 3450 2882 3506
rect 2938 3450 3008 3506
rect 2668 3364 3008 3450
rect 2668 3308 2740 3364
rect 2796 3308 2882 3364
rect 2938 3308 3008 3364
rect 2668 3222 3008 3308
rect 2668 3166 2740 3222
rect 2796 3166 2882 3222
rect 2938 3166 3008 3222
rect 2668 3080 3008 3166
rect 2668 3024 2740 3080
rect 2796 3024 2882 3080
rect 2938 3024 3008 3080
rect 2668 2938 3008 3024
rect 2668 2882 2740 2938
rect 2796 2882 2882 2938
rect 2938 2882 3008 2938
rect 2668 2796 3008 2882
rect 2668 2740 2740 2796
rect 2796 2740 2882 2796
rect 2938 2740 3008 2796
rect 2668 2654 3008 2740
rect 2668 2598 2740 2654
rect 2796 2598 2882 2654
rect 2938 2598 3008 2654
rect 2668 2512 3008 2598
rect 2668 2456 2740 2512
rect 2796 2456 2882 2512
rect 2938 2456 3008 2512
rect 2668 2370 3008 2456
rect 2668 2314 2740 2370
rect 2796 2314 2882 2370
rect 2938 2314 3008 2370
rect 2668 2228 3008 2314
rect 2668 2172 2740 2228
rect 2796 2172 2882 2228
rect 2938 2172 3008 2228
rect 2668 2086 3008 2172
rect 2668 2030 2740 2086
rect 2796 2030 2882 2086
rect 2938 2030 3008 2086
rect 2668 1944 3008 2030
rect 2668 1888 2740 1944
rect 2796 1888 2882 1944
rect 2938 1888 3008 1944
rect 2668 1802 3008 1888
rect 2668 1746 2740 1802
rect 2796 1746 2882 1802
rect 2938 1746 3008 1802
rect 2668 1660 3008 1746
rect 2668 1604 2740 1660
rect 2796 1604 2882 1660
rect 2938 1604 3008 1660
rect 2668 1518 3008 1604
rect 2668 1462 2740 1518
rect 2796 1462 2882 1518
rect 2938 1462 3008 1518
rect 2668 1376 3008 1462
rect 2668 1320 2740 1376
rect 2796 1320 2882 1376
rect 2938 1320 3008 1376
rect 2668 1234 3008 1320
rect 2668 1178 2740 1234
rect 2796 1178 2882 1234
rect 2938 1178 3008 1234
rect 2668 1092 3008 1178
rect 2668 1036 2740 1092
rect 2796 1036 2882 1092
rect 2938 1036 3008 1092
rect 2668 950 3008 1036
rect 2668 894 2740 950
rect 2796 894 2882 950
rect 2938 894 3008 950
rect 2668 808 3008 894
rect 2668 752 2740 808
rect 2796 752 2882 808
rect 2938 752 3008 808
rect 2668 666 3008 752
rect 2668 610 2740 666
rect 2796 610 2882 666
rect 2938 610 3008 666
rect 2668 524 3008 610
rect 2668 468 2740 524
rect 2796 468 2882 524
rect 2938 468 3008 524
rect 2668 400 3008 468
rect 3068 12310 3408 12400
rect 3068 12254 3136 12310
rect 3192 12254 3278 12310
rect 3334 12254 3408 12310
rect 3068 12168 3408 12254
rect 3068 12112 3136 12168
rect 3192 12112 3278 12168
rect 3334 12112 3408 12168
rect 3068 12026 3408 12112
rect 3068 11970 3136 12026
rect 3192 11970 3278 12026
rect 3334 11970 3408 12026
rect 3068 11884 3408 11970
rect 3068 11828 3136 11884
rect 3192 11828 3278 11884
rect 3334 11828 3408 11884
rect 3068 11742 3408 11828
rect 3068 11686 3136 11742
rect 3192 11686 3278 11742
rect 3334 11686 3408 11742
rect 3068 11600 3408 11686
rect 3068 11544 3136 11600
rect 3192 11544 3278 11600
rect 3334 11544 3408 11600
rect 3068 11458 3408 11544
rect 3068 11402 3136 11458
rect 3192 11402 3278 11458
rect 3334 11402 3408 11458
rect 3068 11316 3408 11402
rect 3068 11260 3136 11316
rect 3192 11260 3278 11316
rect 3334 11260 3408 11316
rect 3068 11174 3408 11260
rect 3068 11118 3136 11174
rect 3192 11118 3278 11174
rect 3334 11118 3408 11174
rect 3068 11032 3408 11118
rect 3068 10976 3136 11032
rect 3192 10976 3278 11032
rect 3334 10976 3408 11032
rect 3068 10890 3408 10976
rect 3068 10834 3136 10890
rect 3192 10834 3278 10890
rect 3334 10834 3408 10890
rect 3068 10748 3408 10834
rect 3068 10692 3136 10748
rect 3192 10692 3278 10748
rect 3334 10692 3408 10748
rect 3068 10606 3408 10692
rect 3068 10550 3136 10606
rect 3192 10550 3278 10606
rect 3334 10550 3408 10606
rect 3068 10464 3408 10550
rect 3068 10408 3136 10464
rect 3192 10408 3278 10464
rect 3334 10408 3408 10464
rect 3068 10322 3408 10408
rect 3068 10266 3136 10322
rect 3192 10266 3278 10322
rect 3334 10266 3408 10322
rect 3068 10180 3408 10266
rect 3068 10124 3136 10180
rect 3192 10124 3278 10180
rect 3334 10124 3408 10180
rect 3068 10038 3408 10124
rect 3068 9982 3136 10038
rect 3192 9982 3278 10038
rect 3334 9982 3408 10038
rect 3068 9896 3408 9982
rect 3068 9840 3136 9896
rect 3192 9840 3278 9896
rect 3334 9840 3408 9896
rect 3068 9754 3408 9840
rect 3068 9698 3136 9754
rect 3192 9698 3278 9754
rect 3334 9698 3408 9754
rect 3068 9612 3408 9698
rect 3068 9556 3136 9612
rect 3192 9556 3278 9612
rect 3334 9556 3408 9612
rect 3068 9470 3408 9556
rect 3068 9414 3136 9470
rect 3192 9414 3278 9470
rect 3334 9414 3408 9470
rect 3068 9328 3408 9414
rect 3068 9272 3136 9328
rect 3192 9272 3278 9328
rect 3334 9272 3408 9328
rect 3068 9186 3408 9272
rect 3068 9130 3136 9186
rect 3192 9130 3278 9186
rect 3334 9130 3408 9186
rect 3068 9044 3408 9130
rect 3068 8988 3136 9044
rect 3192 8988 3278 9044
rect 3334 8988 3408 9044
rect 3068 8902 3408 8988
rect 3068 8846 3136 8902
rect 3192 8846 3278 8902
rect 3334 8846 3408 8902
rect 3068 8760 3408 8846
rect 3068 8704 3136 8760
rect 3192 8704 3278 8760
rect 3334 8704 3408 8760
rect 3068 8618 3408 8704
rect 3068 8562 3136 8618
rect 3192 8562 3278 8618
rect 3334 8562 3408 8618
rect 3068 8476 3408 8562
rect 3068 8420 3136 8476
rect 3192 8420 3278 8476
rect 3334 8420 3408 8476
rect 3068 8334 3408 8420
rect 3068 8278 3136 8334
rect 3192 8278 3278 8334
rect 3334 8278 3408 8334
rect 3068 8192 3408 8278
rect 3068 8136 3136 8192
rect 3192 8136 3278 8192
rect 3334 8136 3408 8192
rect 3068 8050 3408 8136
rect 3068 7994 3136 8050
rect 3192 7994 3278 8050
rect 3334 7994 3408 8050
rect 3068 7908 3408 7994
rect 3068 7852 3136 7908
rect 3192 7852 3278 7908
rect 3334 7852 3408 7908
rect 3068 7766 3408 7852
rect 3068 7710 3136 7766
rect 3192 7710 3278 7766
rect 3334 7710 3408 7766
rect 3068 7624 3408 7710
rect 3068 7568 3136 7624
rect 3192 7568 3278 7624
rect 3334 7568 3408 7624
rect 3068 7482 3408 7568
rect 3068 7426 3136 7482
rect 3192 7426 3278 7482
rect 3334 7426 3408 7482
rect 3068 7340 3408 7426
rect 3068 7284 3136 7340
rect 3192 7284 3278 7340
rect 3334 7284 3408 7340
rect 3068 7198 3408 7284
rect 3068 7142 3136 7198
rect 3192 7142 3278 7198
rect 3334 7142 3408 7198
rect 3068 7056 3408 7142
rect 3068 7000 3136 7056
rect 3192 7000 3278 7056
rect 3334 7000 3408 7056
rect 3068 6914 3408 7000
rect 3068 6858 3136 6914
rect 3192 6858 3278 6914
rect 3334 6858 3408 6914
rect 3068 6772 3408 6858
rect 3068 6716 3136 6772
rect 3192 6716 3278 6772
rect 3334 6716 3408 6772
rect 3068 6630 3408 6716
rect 3068 6574 3136 6630
rect 3192 6574 3278 6630
rect 3334 6574 3408 6630
rect 3068 6488 3408 6574
rect 3068 6432 3136 6488
rect 3192 6432 3278 6488
rect 3334 6432 3408 6488
rect 3068 6346 3408 6432
rect 3068 6290 3136 6346
rect 3192 6290 3278 6346
rect 3334 6290 3408 6346
rect 3068 6204 3408 6290
rect 3068 6148 3136 6204
rect 3192 6148 3278 6204
rect 3334 6148 3408 6204
rect 3068 6062 3408 6148
rect 3068 6006 3136 6062
rect 3192 6006 3278 6062
rect 3334 6006 3408 6062
rect 3068 5920 3408 6006
rect 3068 5864 3136 5920
rect 3192 5864 3278 5920
rect 3334 5864 3408 5920
rect 3068 5778 3408 5864
rect 3068 5722 3136 5778
rect 3192 5722 3278 5778
rect 3334 5722 3408 5778
rect 3068 5636 3408 5722
rect 3068 5580 3136 5636
rect 3192 5580 3278 5636
rect 3334 5580 3408 5636
rect 3068 5494 3408 5580
rect 3068 5438 3136 5494
rect 3192 5438 3278 5494
rect 3334 5438 3408 5494
rect 3068 5352 3408 5438
rect 3068 5296 3136 5352
rect 3192 5296 3278 5352
rect 3334 5296 3408 5352
rect 3068 5210 3408 5296
rect 3068 5154 3136 5210
rect 3192 5154 3278 5210
rect 3334 5154 3408 5210
rect 3068 5068 3408 5154
rect 3068 5012 3136 5068
rect 3192 5012 3278 5068
rect 3334 5012 3408 5068
rect 3068 4926 3408 5012
rect 3068 4870 3136 4926
rect 3192 4870 3278 4926
rect 3334 4870 3408 4926
rect 3068 4784 3408 4870
rect 3068 4728 3136 4784
rect 3192 4728 3278 4784
rect 3334 4728 3408 4784
rect 3068 4642 3408 4728
rect 3068 4586 3136 4642
rect 3192 4586 3278 4642
rect 3334 4586 3408 4642
rect 3068 4500 3408 4586
rect 3068 4444 3136 4500
rect 3192 4444 3278 4500
rect 3334 4444 3408 4500
rect 3068 4358 3408 4444
rect 3068 4302 3136 4358
rect 3192 4302 3278 4358
rect 3334 4302 3408 4358
rect 3068 4216 3408 4302
rect 3068 4160 3136 4216
rect 3192 4160 3278 4216
rect 3334 4160 3408 4216
rect 3068 4074 3408 4160
rect 3068 4018 3136 4074
rect 3192 4018 3278 4074
rect 3334 4018 3408 4074
rect 3068 3932 3408 4018
rect 3068 3876 3136 3932
rect 3192 3876 3278 3932
rect 3334 3876 3408 3932
rect 3068 3790 3408 3876
rect 3068 3734 3136 3790
rect 3192 3734 3278 3790
rect 3334 3734 3408 3790
rect 3068 3648 3408 3734
rect 3068 3592 3136 3648
rect 3192 3592 3278 3648
rect 3334 3592 3408 3648
rect 3068 3506 3408 3592
rect 3068 3450 3136 3506
rect 3192 3450 3278 3506
rect 3334 3450 3408 3506
rect 3068 3364 3408 3450
rect 3068 3308 3136 3364
rect 3192 3308 3278 3364
rect 3334 3308 3408 3364
rect 3068 3222 3408 3308
rect 3068 3166 3136 3222
rect 3192 3166 3278 3222
rect 3334 3166 3408 3222
rect 3068 3080 3408 3166
rect 3068 3024 3136 3080
rect 3192 3024 3278 3080
rect 3334 3024 3408 3080
rect 3068 2938 3408 3024
rect 3068 2882 3136 2938
rect 3192 2882 3278 2938
rect 3334 2882 3408 2938
rect 3068 2796 3408 2882
rect 3068 2740 3136 2796
rect 3192 2740 3278 2796
rect 3334 2740 3408 2796
rect 3068 2654 3408 2740
rect 3068 2598 3136 2654
rect 3192 2598 3278 2654
rect 3334 2598 3408 2654
rect 3068 2512 3408 2598
rect 3068 2456 3136 2512
rect 3192 2456 3278 2512
rect 3334 2456 3408 2512
rect 3068 2370 3408 2456
rect 3068 2314 3136 2370
rect 3192 2314 3278 2370
rect 3334 2314 3408 2370
rect 3068 2228 3408 2314
rect 3068 2172 3136 2228
rect 3192 2172 3278 2228
rect 3334 2172 3408 2228
rect 3068 2086 3408 2172
rect 3068 2030 3136 2086
rect 3192 2030 3278 2086
rect 3334 2030 3408 2086
rect 3068 1944 3408 2030
rect 3068 1888 3136 1944
rect 3192 1888 3278 1944
rect 3334 1888 3408 1944
rect 3068 1802 3408 1888
rect 3068 1746 3136 1802
rect 3192 1746 3278 1802
rect 3334 1746 3408 1802
rect 3068 1660 3408 1746
rect 3068 1604 3136 1660
rect 3192 1604 3278 1660
rect 3334 1604 3408 1660
rect 3068 1518 3408 1604
rect 3068 1462 3136 1518
rect 3192 1462 3278 1518
rect 3334 1462 3408 1518
rect 3068 1376 3408 1462
rect 3068 1320 3136 1376
rect 3192 1320 3278 1376
rect 3334 1320 3408 1376
rect 3068 1234 3408 1320
rect 3068 1178 3136 1234
rect 3192 1178 3278 1234
rect 3334 1178 3408 1234
rect 3068 1092 3408 1178
rect 3068 1036 3136 1092
rect 3192 1036 3278 1092
rect 3334 1036 3408 1092
rect 3068 950 3408 1036
rect 3068 894 3136 950
rect 3192 894 3278 950
rect 3334 894 3408 950
rect 3068 808 3408 894
rect 3068 752 3136 808
rect 3192 752 3278 808
rect 3334 752 3408 808
rect 3068 666 3408 752
rect 3068 610 3136 666
rect 3192 610 3278 666
rect 3334 610 3408 666
rect 3068 524 3408 610
rect 3068 468 3136 524
rect 3192 468 3278 524
rect 3334 468 3408 524
rect 3068 400 3408 468
rect 3468 12310 3808 12400
rect 3468 12254 3536 12310
rect 3592 12254 3678 12310
rect 3734 12254 3808 12310
rect 3468 12168 3808 12254
rect 3468 12112 3536 12168
rect 3592 12112 3678 12168
rect 3734 12112 3808 12168
rect 3468 12026 3808 12112
rect 3468 11970 3536 12026
rect 3592 11970 3678 12026
rect 3734 11970 3808 12026
rect 3468 11884 3808 11970
rect 3468 11828 3536 11884
rect 3592 11828 3678 11884
rect 3734 11828 3808 11884
rect 3468 11742 3808 11828
rect 3468 11686 3536 11742
rect 3592 11686 3678 11742
rect 3734 11686 3808 11742
rect 3468 11600 3808 11686
rect 3468 11544 3536 11600
rect 3592 11544 3678 11600
rect 3734 11544 3808 11600
rect 3468 11458 3808 11544
rect 3468 11402 3536 11458
rect 3592 11402 3678 11458
rect 3734 11402 3808 11458
rect 3468 11316 3808 11402
rect 3468 11260 3536 11316
rect 3592 11260 3678 11316
rect 3734 11260 3808 11316
rect 3468 11174 3808 11260
rect 3468 11118 3536 11174
rect 3592 11118 3678 11174
rect 3734 11118 3808 11174
rect 3468 11032 3808 11118
rect 3468 10976 3536 11032
rect 3592 10976 3678 11032
rect 3734 10976 3808 11032
rect 3468 10890 3808 10976
rect 3468 10834 3536 10890
rect 3592 10834 3678 10890
rect 3734 10834 3808 10890
rect 3468 10748 3808 10834
rect 3468 10692 3536 10748
rect 3592 10692 3678 10748
rect 3734 10692 3808 10748
rect 3468 10606 3808 10692
rect 3468 10550 3536 10606
rect 3592 10550 3678 10606
rect 3734 10550 3808 10606
rect 3468 10464 3808 10550
rect 3468 10408 3536 10464
rect 3592 10408 3678 10464
rect 3734 10408 3808 10464
rect 3468 10322 3808 10408
rect 3468 10266 3536 10322
rect 3592 10266 3678 10322
rect 3734 10266 3808 10322
rect 3468 10180 3808 10266
rect 3468 10124 3536 10180
rect 3592 10124 3678 10180
rect 3734 10124 3808 10180
rect 3468 10038 3808 10124
rect 3468 9982 3536 10038
rect 3592 9982 3678 10038
rect 3734 9982 3808 10038
rect 3468 9896 3808 9982
rect 3468 9840 3536 9896
rect 3592 9840 3678 9896
rect 3734 9840 3808 9896
rect 3468 9754 3808 9840
rect 3468 9698 3536 9754
rect 3592 9698 3678 9754
rect 3734 9698 3808 9754
rect 3468 9612 3808 9698
rect 3468 9556 3536 9612
rect 3592 9556 3678 9612
rect 3734 9556 3808 9612
rect 3468 9470 3808 9556
rect 3468 9414 3536 9470
rect 3592 9414 3678 9470
rect 3734 9414 3808 9470
rect 3468 9328 3808 9414
rect 3468 9272 3536 9328
rect 3592 9272 3678 9328
rect 3734 9272 3808 9328
rect 3468 9186 3808 9272
rect 3468 9130 3536 9186
rect 3592 9130 3678 9186
rect 3734 9130 3808 9186
rect 3468 9044 3808 9130
rect 3468 8988 3536 9044
rect 3592 8988 3678 9044
rect 3734 8988 3808 9044
rect 3468 8902 3808 8988
rect 3468 8846 3536 8902
rect 3592 8846 3678 8902
rect 3734 8846 3808 8902
rect 3468 8760 3808 8846
rect 3468 8704 3536 8760
rect 3592 8704 3678 8760
rect 3734 8704 3808 8760
rect 3468 8618 3808 8704
rect 3468 8562 3536 8618
rect 3592 8562 3678 8618
rect 3734 8562 3808 8618
rect 3468 8476 3808 8562
rect 3468 8420 3536 8476
rect 3592 8420 3678 8476
rect 3734 8420 3808 8476
rect 3468 8334 3808 8420
rect 3468 8278 3536 8334
rect 3592 8278 3678 8334
rect 3734 8278 3808 8334
rect 3468 8192 3808 8278
rect 3468 8136 3536 8192
rect 3592 8136 3678 8192
rect 3734 8136 3808 8192
rect 3468 8050 3808 8136
rect 3468 7994 3536 8050
rect 3592 7994 3678 8050
rect 3734 7994 3808 8050
rect 3468 7908 3808 7994
rect 3468 7852 3536 7908
rect 3592 7852 3678 7908
rect 3734 7852 3808 7908
rect 3468 7766 3808 7852
rect 3468 7710 3536 7766
rect 3592 7710 3678 7766
rect 3734 7710 3808 7766
rect 3468 7624 3808 7710
rect 3468 7568 3536 7624
rect 3592 7568 3678 7624
rect 3734 7568 3808 7624
rect 3468 7482 3808 7568
rect 3468 7426 3536 7482
rect 3592 7426 3678 7482
rect 3734 7426 3808 7482
rect 3468 7340 3808 7426
rect 3468 7284 3536 7340
rect 3592 7284 3678 7340
rect 3734 7284 3808 7340
rect 3468 7198 3808 7284
rect 3468 7142 3536 7198
rect 3592 7142 3678 7198
rect 3734 7142 3808 7198
rect 3468 7056 3808 7142
rect 3468 7000 3536 7056
rect 3592 7000 3678 7056
rect 3734 7000 3808 7056
rect 3468 6914 3808 7000
rect 3468 6858 3536 6914
rect 3592 6858 3678 6914
rect 3734 6858 3808 6914
rect 3468 6772 3808 6858
rect 3468 6716 3536 6772
rect 3592 6716 3678 6772
rect 3734 6716 3808 6772
rect 3468 6630 3808 6716
rect 3468 6574 3536 6630
rect 3592 6574 3678 6630
rect 3734 6574 3808 6630
rect 3468 6488 3808 6574
rect 3468 6432 3536 6488
rect 3592 6432 3678 6488
rect 3734 6432 3808 6488
rect 3468 6346 3808 6432
rect 3468 6290 3536 6346
rect 3592 6290 3678 6346
rect 3734 6290 3808 6346
rect 3468 6204 3808 6290
rect 3468 6148 3536 6204
rect 3592 6148 3678 6204
rect 3734 6148 3808 6204
rect 3468 6062 3808 6148
rect 3468 6006 3536 6062
rect 3592 6006 3678 6062
rect 3734 6006 3808 6062
rect 3468 5920 3808 6006
rect 3468 5864 3536 5920
rect 3592 5864 3678 5920
rect 3734 5864 3808 5920
rect 3468 5778 3808 5864
rect 3468 5722 3536 5778
rect 3592 5722 3678 5778
rect 3734 5722 3808 5778
rect 3468 5636 3808 5722
rect 3468 5580 3536 5636
rect 3592 5580 3678 5636
rect 3734 5580 3808 5636
rect 3468 5494 3808 5580
rect 3468 5438 3536 5494
rect 3592 5438 3678 5494
rect 3734 5438 3808 5494
rect 3468 5352 3808 5438
rect 3468 5296 3536 5352
rect 3592 5296 3678 5352
rect 3734 5296 3808 5352
rect 3468 5210 3808 5296
rect 3468 5154 3536 5210
rect 3592 5154 3678 5210
rect 3734 5154 3808 5210
rect 3468 5068 3808 5154
rect 3468 5012 3536 5068
rect 3592 5012 3678 5068
rect 3734 5012 3808 5068
rect 3468 4926 3808 5012
rect 3468 4870 3536 4926
rect 3592 4870 3678 4926
rect 3734 4870 3808 4926
rect 3468 4784 3808 4870
rect 3468 4728 3536 4784
rect 3592 4728 3678 4784
rect 3734 4728 3808 4784
rect 3468 4642 3808 4728
rect 3468 4586 3536 4642
rect 3592 4586 3678 4642
rect 3734 4586 3808 4642
rect 3468 4500 3808 4586
rect 3468 4444 3536 4500
rect 3592 4444 3678 4500
rect 3734 4444 3808 4500
rect 3468 4358 3808 4444
rect 3468 4302 3536 4358
rect 3592 4302 3678 4358
rect 3734 4302 3808 4358
rect 3468 4216 3808 4302
rect 3468 4160 3536 4216
rect 3592 4160 3678 4216
rect 3734 4160 3808 4216
rect 3468 4074 3808 4160
rect 3468 4018 3536 4074
rect 3592 4018 3678 4074
rect 3734 4018 3808 4074
rect 3468 3932 3808 4018
rect 3468 3876 3536 3932
rect 3592 3876 3678 3932
rect 3734 3876 3808 3932
rect 3468 3790 3808 3876
rect 3468 3734 3536 3790
rect 3592 3734 3678 3790
rect 3734 3734 3808 3790
rect 3468 3648 3808 3734
rect 3468 3592 3536 3648
rect 3592 3592 3678 3648
rect 3734 3592 3808 3648
rect 3468 3506 3808 3592
rect 3468 3450 3536 3506
rect 3592 3450 3678 3506
rect 3734 3450 3808 3506
rect 3468 3364 3808 3450
rect 3468 3308 3536 3364
rect 3592 3308 3678 3364
rect 3734 3308 3808 3364
rect 3468 3222 3808 3308
rect 3468 3166 3536 3222
rect 3592 3166 3678 3222
rect 3734 3166 3808 3222
rect 3468 3080 3808 3166
rect 3468 3024 3536 3080
rect 3592 3024 3678 3080
rect 3734 3024 3808 3080
rect 3468 2938 3808 3024
rect 3468 2882 3536 2938
rect 3592 2882 3678 2938
rect 3734 2882 3808 2938
rect 3468 2796 3808 2882
rect 3468 2740 3536 2796
rect 3592 2740 3678 2796
rect 3734 2740 3808 2796
rect 3468 2654 3808 2740
rect 3468 2598 3536 2654
rect 3592 2598 3678 2654
rect 3734 2598 3808 2654
rect 3468 2512 3808 2598
rect 3468 2456 3536 2512
rect 3592 2456 3678 2512
rect 3734 2456 3808 2512
rect 3468 2370 3808 2456
rect 3468 2314 3536 2370
rect 3592 2314 3678 2370
rect 3734 2314 3808 2370
rect 3468 2228 3808 2314
rect 3468 2172 3536 2228
rect 3592 2172 3678 2228
rect 3734 2172 3808 2228
rect 3468 2086 3808 2172
rect 3468 2030 3536 2086
rect 3592 2030 3678 2086
rect 3734 2030 3808 2086
rect 3468 1944 3808 2030
rect 3468 1888 3536 1944
rect 3592 1888 3678 1944
rect 3734 1888 3808 1944
rect 3468 1802 3808 1888
rect 3468 1746 3536 1802
rect 3592 1746 3678 1802
rect 3734 1746 3808 1802
rect 3468 1660 3808 1746
rect 3468 1604 3536 1660
rect 3592 1604 3678 1660
rect 3734 1604 3808 1660
rect 3468 1518 3808 1604
rect 3468 1462 3536 1518
rect 3592 1462 3678 1518
rect 3734 1462 3808 1518
rect 3468 1376 3808 1462
rect 3468 1320 3536 1376
rect 3592 1320 3678 1376
rect 3734 1320 3808 1376
rect 3468 1234 3808 1320
rect 3468 1178 3536 1234
rect 3592 1178 3678 1234
rect 3734 1178 3808 1234
rect 3468 1092 3808 1178
rect 3468 1036 3536 1092
rect 3592 1036 3678 1092
rect 3734 1036 3808 1092
rect 3468 950 3808 1036
rect 3468 894 3536 950
rect 3592 894 3678 950
rect 3734 894 3808 950
rect 3468 808 3808 894
rect 3468 752 3536 808
rect 3592 752 3678 808
rect 3734 752 3808 808
rect 3468 666 3808 752
rect 3468 610 3536 666
rect 3592 610 3678 666
rect 3734 610 3808 666
rect 3468 524 3808 610
rect 3468 468 3536 524
rect 3592 468 3678 524
rect 3734 468 3808 524
rect 3468 400 3808 468
rect 3868 12310 4208 12400
rect 3868 12254 3933 12310
rect 3989 12254 4075 12310
rect 4131 12254 4208 12310
rect 3868 12168 4208 12254
rect 3868 12112 3933 12168
rect 3989 12112 4075 12168
rect 4131 12112 4208 12168
rect 3868 12026 4208 12112
rect 3868 11970 3933 12026
rect 3989 11970 4075 12026
rect 4131 11970 4208 12026
rect 3868 11884 4208 11970
rect 3868 11828 3933 11884
rect 3989 11828 4075 11884
rect 4131 11828 4208 11884
rect 3868 11742 4208 11828
rect 3868 11686 3933 11742
rect 3989 11686 4075 11742
rect 4131 11686 4208 11742
rect 3868 11600 4208 11686
rect 3868 11544 3933 11600
rect 3989 11544 4075 11600
rect 4131 11544 4208 11600
rect 3868 11458 4208 11544
rect 3868 11402 3933 11458
rect 3989 11402 4075 11458
rect 4131 11402 4208 11458
rect 3868 11316 4208 11402
rect 3868 11260 3933 11316
rect 3989 11260 4075 11316
rect 4131 11260 4208 11316
rect 3868 11174 4208 11260
rect 3868 11118 3933 11174
rect 3989 11118 4075 11174
rect 4131 11118 4208 11174
rect 3868 11032 4208 11118
rect 3868 10976 3933 11032
rect 3989 10976 4075 11032
rect 4131 10976 4208 11032
rect 3868 10890 4208 10976
rect 3868 10834 3933 10890
rect 3989 10834 4075 10890
rect 4131 10834 4208 10890
rect 3868 10748 4208 10834
rect 3868 10692 3933 10748
rect 3989 10692 4075 10748
rect 4131 10692 4208 10748
rect 3868 10606 4208 10692
rect 3868 10550 3933 10606
rect 3989 10550 4075 10606
rect 4131 10550 4208 10606
rect 3868 10464 4208 10550
rect 3868 10408 3933 10464
rect 3989 10408 4075 10464
rect 4131 10408 4208 10464
rect 3868 10322 4208 10408
rect 3868 10266 3933 10322
rect 3989 10266 4075 10322
rect 4131 10266 4208 10322
rect 3868 10180 4208 10266
rect 3868 10124 3933 10180
rect 3989 10124 4075 10180
rect 4131 10124 4208 10180
rect 3868 10038 4208 10124
rect 3868 9982 3933 10038
rect 3989 9982 4075 10038
rect 4131 9982 4208 10038
rect 3868 9896 4208 9982
rect 3868 9840 3933 9896
rect 3989 9840 4075 9896
rect 4131 9840 4208 9896
rect 3868 9754 4208 9840
rect 3868 9698 3933 9754
rect 3989 9698 4075 9754
rect 4131 9698 4208 9754
rect 3868 9612 4208 9698
rect 3868 9556 3933 9612
rect 3989 9556 4075 9612
rect 4131 9556 4208 9612
rect 3868 9470 4208 9556
rect 3868 9414 3933 9470
rect 3989 9414 4075 9470
rect 4131 9414 4208 9470
rect 3868 9328 4208 9414
rect 3868 9272 3933 9328
rect 3989 9272 4075 9328
rect 4131 9272 4208 9328
rect 3868 9186 4208 9272
rect 3868 9130 3933 9186
rect 3989 9130 4075 9186
rect 4131 9130 4208 9186
rect 3868 9044 4208 9130
rect 3868 8988 3933 9044
rect 3989 8988 4075 9044
rect 4131 8988 4208 9044
rect 3868 8902 4208 8988
rect 3868 8846 3933 8902
rect 3989 8846 4075 8902
rect 4131 8846 4208 8902
rect 3868 8760 4208 8846
rect 3868 8704 3933 8760
rect 3989 8704 4075 8760
rect 4131 8704 4208 8760
rect 3868 8618 4208 8704
rect 3868 8562 3933 8618
rect 3989 8562 4075 8618
rect 4131 8562 4208 8618
rect 3868 8476 4208 8562
rect 3868 8420 3933 8476
rect 3989 8420 4075 8476
rect 4131 8420 4208 8476
rect 3868 8334 4208 8420
rect 3868 8278 3933 8334
rect 3989 8278 4075 8334
rect 4131 8278 4208 8334
rect 3868 8192 4208 8278
rect 3868 8136 3933 8192
rect 3989 8136 4075 8192
rect 4131 8136 4208 8192
rect 3868 8050 4208 8136
rect 3868 7994 3933 8050
rect 3989 7994 4075 8050
rect 4131 7994 4208 8050
rect 3868 7908 4208 7994
rect 3868 7852 3933 7908
rect 3989 7852 4075 7908
rect 4131 7852 4208 7908
rect 3868 7766 4208 7852
rect 3868 7710 3933 7766
rect 3989 7710 4075 7766
rect 4131 7710 4208 7766
rect 3868 7624 4208 7710
rect 3868 7568 3933 7624
rect 3989 7568 4075 7624
rect 4131 7568 4208 7624
rect 3868 7482 4208 7568
rect 3868 7426 3933 7482
rect 3989 7426 4075 7482
rect 4131 7426 4208 7482
rect 3868 7340 4208 7426
rect 3868 7284 3933 7340
rect 3989 7284 4075 7340
rect 4131 7284 4208 7340
rect 3868 7198 4208 7284
rect 3868 7142 3933 7198
rect 3989 7142 4075 7198
rect 4131 7142 4208 7198
rect 3868 7056 4208 7142
rect 3868 7000 3933 7056
rect 3989 7000 4075 7056
rect 4131 7000 4208 7056
rect 3868 6914 4208 7000
rect 3868 6858 3933 6914
rect 3989 6858 4075 6914
rect 4131 6858 4208 6914
rect 3868 6772 4208 6858
rect 3868 6716 3933 6772
rect 3989 6716 4075 6772
rect 4131 6716 4208 6772
rect 3868 6630 4208 6716
rect 3868 6574 3933 6630
rect 3989 6574 4075 6630
rect 4131 6574 4208 6630
rect 3868 6488 4208 6574
rect 3868 6432 3933 6488
rect 3989 6432 4075 6488
rect 4131 6432 4208 6488
rect 3868 6346 4208 6432
rect 3868 6290 3933 6346
rect 3989 6290 4075 6346
rect 4131 6290 4208 6346
rect 3868 6204 4208 6290
rect 3868 6148 3933 6204
rect 3989 6148 4075 6204
rect 4131 6148 4208 6204
rect 3868 6062 4208 6148
rect 3868 6006 3933 6062
rect 3989 6006 4075 6062
rect 4131 6006 4208 6062
rect 3868 5920 4208 6006
rect 3868 5864 3933 5920
rect 3989 5864 4075 5920
rect 4131 5864 4208 5920
rect 3868 5778 4208 5864
rect 3868 5722 3933 5778
rect 3989 5722 4075 5778
rect 4131 5722 4208 5778
rect 3868 5636 4208 5722
rect 3868 5580 3933 5636
rect 3989 5580 4075 5636
rect 4131 5580 4208 5636
rect 3868 5494 4208 5580
rect 3868 5438 3933 5494
rect 3989 5438 4075 5494
rect 4131 5438 4208 5494
rect 3868 5352 4208 5438
rect 3868 5296 3933 5352
rect 3989 5296 4075 5352
rect 4131 5296 4208 5352
rect 3868 5210 4208 5296
rect 3868 5154 3933 5210
rect 3989 5154 4075 5210
rect 4131 5154 4208 5210
rect 3868 5068 4208 5154
rect 3868 5012 3933 5068
rect 3989 5012 4075 5068
rect 4131 5012 4208 5068
rect 3868 4926 4208 5012
rect 3868 4870 3933 4926
rect 3989 4870 4075 4926
rect 4131 4870 4208 4926
rect 3868 4784 4208 4870
rect 3868 4728 3933 4784
rect 3989 4728 4075 4784
rect 4131 4728 4208 4784
rect 3868 4642 4208 4728
rect 3868 4586 3933 4642
rect 3989 4586 4075 4642
rect 4131 4586 4208 4642
rect 3868 4500 4208 4586
rect 3868 4444 3933 4500
rect 3989 4444 4075 4500
rect 4131 4444 4208 4500
rect 3868 4358 4208 4444
rect 3868 4302 3933 4358
rect 3989 4302 4075 4358
rect 4131 4302 4208 4358
rect 3868 4216 4208 4302
rect 3868 4160 3933 4216
rect 3989 4160 4075 4216
rect 4131 4160 4208 4216
rect 3868 4074 4208 4160
rect 3868 4018 3933 4074
rect 3989 4018 4075 4074
rect 4131 4018 4208 4074
rect 3868 3932 4208 4018
rect 3868 3876 3933 3932
rect 3989 3876 4075 3932
rect 4131 3876 4208 3932
rect 3868 3790 4208 3876
rect 3868 3734 3933 3790
rect 3989 3734 4075 3790
rect 4131 3734 4208 3790
rect 3868 3648 4208 3734
rect 3868 3592 3933 3648
rect 3989 3592 4075 3648
rect 4131 3592 4208 3648
rect 3868 3506 4208 3592
rect 3868 3450 3933 3506
rect 3989 3450 4075 3506
rect 4131 3450 4208 3506
rect 3868 3364 4208 3450
rect 3868 3308 3933 3364
rect 3989 3308 4075 3364
rect 4131 3308 4208 3364
rect 3868 3222 4208 3308
rect 3868 3166 3933 3222
rect 3989 3166 4075 3222
rect 4131 3166 4208 3222
rect 3868 3080 4208 3166
rect 3868 3024 3933 3080
rect 3989 3024 4075 3080
rect 4131 3024 4208 3080
rect 3868 2938 4208 3024
rect 3868 2882 3933 2938
rect 3989 2882 4075 2938
rect 4131 2882 4208 2938
rect 3868 2796 4208 2882
rect 3868 2740 3933 2796
rect 3989 2740 4075 2796
rect 4131 2740 4208 2796
rect 3868 2654 4208 2740
rect 3868 2598 3933 2654
rect 3989 2598 4075 2654
rect 4131 2598 4208 2654
rect 3868 2512 4208 2598
rect 3868 2456 3933 2512
rect 3989 2456 4075 2512
rect 4131 2456 4208 2512
rect 3868 2370 4208 2456
rect 3868 2314 3933 2370
rect 3989 2314 4075 2370
rect 4131 2314 4208 2370
rect 3868 2228 4208 2314
rect 3868 2172 3933 2228
rect 3989 2172 4075 2228
rect 4131 2172 4208 2228
rect 3868 2086 4208 2172
rect 3868 2030 3933 2086
rect 3989 2030 4075 2086
rect 4131 2030 4208 2086
rect 3868 1944 4208 2030
rect 3868 1888 3933 1944
rect 3989 1888 4075 1944
rect 4131 1888 4208 1944
rect 3868 1802 4208 1888
rect 3868 1746 3933 1802
rect 3989 1746 4075 1802
rect 4131 1746 4208 1802
rect 3868 1660 4208 1746
rect 3868 1604 3933 1660
rect 3989 1604 4075 1660
rect 4131 1604 4208 1660
rect 3868 1518 4208 1604
rect 3868 1462 3933 1518
rect 3989 1462 4075 1518
rect 4131 1462 4208 1518
rect 3868 1376 4208 1462
rect 3868 1320 3933 1376
rect 3989 1320 4075 1376
rect 4131 1320 4208 1376
rect 3868 1234 4208 1320
rect 3868 1178 3933 1234
rect 3989 1178 4075 1234
rect 4131 1178 4208 1234
rect 3868 1092 4208 1178
rect 3868 1036 3933 1092
rect 3989 1036 4075 1092
rect 4131 1036 4208 1092
rect 3868 950 4208 1036
rect 3868 894 3933 950
rect 3989 894 4075 950
rect 4131 894 4208 950
rect 3868 808 4208 894
rect 3868 752 3933 808
rect 3989 752 4075 808
rect 4131 752 4208 808
rect 3868 666 4208 752
rect 3868 610 3933 666
rect 3989 610 4075 666
rect 4131 610 4208 666
rect 3868 524 4208 610
rect 3868 468 3933 524
rect 3989 468 4075 524
rect 4131 468 4208 524
rect 3868 400 4208 468
rect 4268 12310 4608 12400
rect 4268 12254 4338 12310
rect 4394 12254 4480 12310
rect 4536 12254 4608 12310
rect 4268 12168 4608 12254
rect 4268 12112 4338 12168
rect 4394 12112 4480 12168
rect 4536 12112 4608 12168
rect 4268 12026 4608 12112
rect 4268 11970 4338 12026
rect 4394 11970 4480 12026
rect 4536 11970 4608 12026
rect 4268 11884 4608 11970
rect 4268 11828 4338 11884
rect 4394 11828 4480 11884
rect 4536 11828 4608 11884
rect 4268 11742 4608 11828
rect 4268 11686 4338 11742
rect 4394 11686 4480 11742
rect 4536 11686 4608 11742
rect 4268 11600 4608 11686
rect 4268 11544 4338 11600
rect 4394 11544 4480 11600
rect 4536 11544 4608 11600
rect 4268 11458 4608 11544
rect 4268 11402 4338 11458
rect 4394 11402 4480 11458
rect 4536 11402 4608 11458
rect 4268 11316 4608 11402
rect 4268 11260 4338 11316
rect 4394 11260 4480 11316
rect 4536 11260 4608 11316
rect 4268 11174 4608 11260
rect 4268 11118 4338 11174
rect 4394 11118 4480 11174
rect 4536 11118 4608 11174
rect 4268 11032 4608 11118
rect 4268 10976 4338 11032
rect 4394 10976 4480 11032
rect 4536 10976 4608 11032
rect 4268 10890 4608 10976
rect 4268 10834 4338 10890
rect 4394 10834 4480 10890
rect 4536 10834 4608 10890
rect 4268 10748 4608 10834
rect 4268 10692 4338 10748
rect 4394 10692 4480 10748
rect 4536 10692 4608 10748
rect 4268 10606 4608 10692
rect 4268 10550 4338 10606
rect 4394 10550 4480 10606
rect 4536 10550 4608 10606
rect 4268 10464 4608 10550
rect 4268 10408 4338 10464
rect 4394 10408 4480 10464
rect 4536 10408 4608 10464
rect 4268 10322 4608 10408
rect 4268 10266 4338 10322
rect 4394 10266 4480 10322
rect 4536 10266 4608 10322
rect 4268 10180 4608 10266
rect 4268 10124 4338 10180
rect 4394 10124 4480 10180
rect 4536 10124 4608 10180
rect 4268 10038 4608 10124
rect 4268 9982 4338 10038
rect 4394 9982 4480 10038
rect 4536 9982 4608 10038
rect 4268 9896 4608 9982
rect 4268 9840 4338 9896
rect 4394 9840 4480 9896
rect 4536 9840 4608 9896
rect 4268 9754 4608 9840
rect 4268 9698 4338 9754
rect 4394 9698 4480 9754
rect 4536 9698 4608 9754
rect 4268 9612 4608 9698
rect 4268 9556 4338 9612
rect 4394 9556 4480 9612
rect 4536 9556 4608 9612
rect 4268 9470 4608 9556
rect 4268 9414 4338 9470
rect 4394 9414 4480 9470
rect 4536 9414 4608 9470
rect 4268 9328 4608 9414
rect 4268 9272 4338 9328
rect 4394 9272 4480 9328
rect 4536 9272 4608 9328
rect 4268 9186 4608 9272
rect 4268 9130 4338 9186
rect 4394 9130 4480 9186
rect 4536 9130 4608 9186
rect 4268 9044 4608 9130
rect 4268 8988 4338 9044
rect 4394 8988 4480 9044
rect 4536 8988 4608 9044
rect 4268 8902 4608 8988
rect 4268 8846 4338 8902
rect 4394 8846 4480 8902
rect 4536 8846 4608 8902
rect 4268 8760 4608 8846
rect 4268 8704 4338 8760
rect 4394 8704 4480 8760
rect 4536 8704 4608 8760
rect 4268 8618 4608 8704
rect 4268 8562 4338 8618
rect 4394 8562 4480 8618
rect 4536 8562 4608 8618
rect 4268 8476 4608 8562
rect 4268 8420 4338 8476
rect 4394 8420 4480 8476
rect 4536 8420 4608 8476
rect 4268 8334 4608 8420
rect 4268 8278 4338 8334
rect 4394 8278 4480 8334
rect 4536 8278 4608 8334
rect 4268 8192 4608 8278
rect 4268 8136 4338 8192
rect 4394 8136 4480 8192
rect 4536 8136 4608 8192
rect 4268 8050 4608 8136
rect 4268 7994 4338 8050
rect 4394 7994 4480 8050
rect 4536 7994 4608 8050
rect 4268 7908 4608 7994
rect 4268 7852 4338 7908
rect 4394 7852 4480 7908
rect 4536 7852 4608 7908
rect 4268 7766 4608 7852
rect 4268 7710 4338 7766
rect 4394 7710 4480 7766
rect 4536 7710 4608 7766
rect 4268 7624 4608 7710
rect 4268 7568 4338 7624
rect 4394 7568 4480 7624
rect 4536 7568 4608 7624
rect 4268 7482 4608 7568
rect 4268 7426 4338 7482
rect 4394 7426 4480 7482
rect 4536 7426 4608 7482
rect 4268 7340 4608 7426
rect 4268 7284 4338 7340
rect 4394 7284 4480 7340
rect 4536 7284 4608 7340
rect 4268 7198 4608 7284
rect 4268 7142 4338 7198
rect 4394 7142 4480 7198
rect 4536 7142 4608 7198
rect 4268 7056 4608 7142
rect 4268 7000 4338 7056
rect 4394 7000 4480 7056
rect 4536 7000 4608 7056
rect 4268 6914 4608 7000
rect 4268 6858 4338 6914
rect 4394 6858 4480 6914
rect 4536 6858 4608 6914
rect 4268 6772 4608 6858
rect 4268 6716 4338 6772
rect 4394 6716 4480 6772
rect 4536 6716 4608 6772
rect 4268 6630 4608 6716
rect 4268 6574 4338 6630
rect 4394 6574 4480 6630
rect 4536 6574 4608 6630
rect 4268 6488 4608 6574
rect 4268 6432 4338 6488
rect 4394 6432 4480 6488
rect 4536 6432 4608 6488
rect 4268 6346 4608 6432
rect 4268 6290 4338 6346
rect 4394 6290 4480 6346
rect 4536 6290 4608 6346
rect 4268 6204 4608 6290
rect 4268 6148 4338 6204
rect 4394 6148 4480 6204
rect 4536 6148 4608 6204
rect 4268 6062 4608 6148
rect 4268 6006 4338 6062
rect 4394 6006 4480 6062
rect 4536 6006 4608 6062
rect 4268 5920 4608 6006
rect 4268 5864 4338 5920
rect 4394 5864 4480 5920
rect 4536 5864 4608 5920
rect 4268 5778 4608 5864
rect 4268 5722 4338 5778
rect 4394 5722 4480 5778
rect 4536 5722 4608 5778
rect 4268 5636 4608 5722
rect 4268 5580 4338 5636
rect 4394 5580 4480 5636
rect 4536 5580 4608 5636
rect 4268 5494 4608 5580
rect 4268 5438 4338 5494
rect 4394 5438 4480 5494
rect 4536 5438 4608 5494
rect 4268 5352 4608 5438
rect 4268 5296 4338 5352
rect 4394 5296 4480 5352
rect 4536 5296 4608 5352
rect 4268 5210 4608 5296
rect 4268 5154 4338 5210
rect 4394 5154 4480 5210
rect 4536 5154 4608 5210
rect 4268 5068 4608 5154
rect 4268 5012 4338 5068
rect 4394 5012 4480 5068
rect 4536 5012 4608 5068
rect 4268 4926 4608 5012
rect 4268 4870 4338 4926
rect 4394 4870 4480 4926
rect 4536 4870 4608 4926
rect 4268 4784 4608 4870
rect 4268 4728 4338 4784
rect 4394 4728 4480 4784
rect 4536 4728 4608 4784
rect 4268 4642 4608 4728
rect 4268 4586 4338 4642
rect 4394 4586 4480 4642
rect 4536 4586 4608 4642
rect 4268 4500 4608 4586
rect 4268 4444 4338 4500
rect 4394 4444 4480 4500
rect 4536 4444 4608 4500
rect 4268 4358 4608 4444
rect 4268 4302 4338 4358
rect 4394 4302 4480 4358
rect 4536 4302 4608 4358
rect 4268 4216 4608 4302
rect 4268 4160 4338 4216
rect 4394 4160 4480 4216
rect 4536 4160 4608 4216
rect 4268 4074 4608 4160
rect 4268 4018 4338 4074
rect 4394 4018 4480 4074
rect 4536 4018 4608 4074
rect 4268 3932 4608 4018
rect 4268 3876 4338 3932
rect 4394 3876 4480 3932
rect 4536 3876 4608 3932
rect 4268 3790 4608 3876
rect 4268 3734 4338 3790
rect 4394 3734 4480 3790
rect 4536 3734 4608 3790
rect 4268 3648 4608 3734
rect 4268 3592 4338 3648
rect 4394 3592 4480 3648
rect 4536 3592 4608 3648
rect 4268 3506 4608 3592
rect 4268 3450 4338 3506
rect 4394 3450 4480 3506
rect 4536 3450 4608 3506
rect 4268 3364 4608 3450
rect 4268 3308 4338 3364
rect 4394 3308 4480 3364
rect 4536 3308 4608 3364
rect 4268 3222 4608 3308
rect 4268 3166 4338 3222
rect 4394 3166 4480 3222
rect 4536 3166 4608 3222
rect 4268 3080 4608 3166
rect 4268 3024 4338 3080
rect 4394 3024 4480 3080
rect 4536 3024 4608 3080
rect 4268 2938 4608 3024
rect 4268 2882 4338 2938
rect 4394 2882 4480 2938
rect 4536 2882 4608 2938
rect 4268 2796 4608 2882
rect 4268 2740 4338 2796
rect 4394 2740 4480 2796
rect 4536 2740 4608 2796
rect 4268 2654 4608 2740
rect 4268 2598 4338 2654
rect 4394 2598 4480 2654
rect 4536 2598 4608 2654
rect 4268 2512 4608 2598
rect 4268 2456 4338 2512
rect 4394 2456 4480 2512
rect 4536 2456 4608 2512
rect 4268 2370 4608 2456
rect 4268 2314 4338 2370
rect 4394 2314 4480 2370
rect 4536 2314 4608 2370
rect 4268 2228 4608 2314
rect 4268 2172 4338 2228
rect 4394 2172 4480 2228
rect 4536 2172 4608 2228
rect 4268 2086 4608 2172
rect 4268 2030 4338 2086
rect 4394 2030 4480 2086
rect 4536 2030 4608 2086
rect 4268 1944 4608 2030
rect 4268 1888 4338 1944
rect 4394 1888 4480 1944
rect 4536 1888 4608 1944
rect 4268 1802 4608 1888
rect 4268 1746 4338 1802
rect 4394 1746 4480 1802
rect 4536 1746 4608 1802
rect 4268 1660 4608 1746
rect 4268 1604 4338 1660
rect 4394 1604 4480 1660
rect 4536 1604 4608 1660
rect 4268 1518 4608 1604
rect 4268 1462 4338 1518
rect 4394 1462 4480 1518
rect 4536 1462 4608 1518
rect 4268 1376 4608 1462
rect 4268 1320 4338 1376
rect 4394 1320 4480 1376
rect 4536 1320 4608 1376
rect 4268 1234 4608 1320
rect 4268 1178 4338 1234
rect 4394 1178 4480 1234
rect 4536 1178 4608 1234
rect 4268 1092 4608 1178
rect 4268 1036 4338 1092
rect 4394 1036 4480 1092
rect 4536 1036 4608 1092
rect 4268 950 4608 1036
rect 4268 894 4338 950
rect 4394 894 4480 950
rect 4536 894 4608 950
rect 4268 808 4608 894
rect 4268 752 4338 808
rect 4394 752 4480 808
rect 4536 752 4608 808
rect 4268 666 4608 752
rect 4268 610 4338 666
rect 4394 610 4480 666
rect 4536 610 4608 666
rect 4268 524 4608 610
rect 4268 468 4338 524
rect 4394 468 4480 524
rect 4536 468 4608 524
rect 4268 400 4608 468
rect 4668 12310 5008 12400
rect 4668 12254 4738 12310
rect 4794 12254 4880 12310
rect 4936 12254 5008 12310
rect 4668 12168 5008 12254
rect 4668 12112 4738 12168
rect 4794 12112 4880 12168
rect 4936 12112 5008 12168
rect 4668 12026 5008 12112
rect 4668 11970 4738 12026
rect 4794 11970 4880 12026
rect 4936 11970 5008 12026
rect 4668 11884 5008 11970
rect 4668 11828 4738 11884
rect 4794 11828 4880 11884
rect 4936 11828 5008 11884
rect 4668 11742 5008 11828
rect 4668 11686 4738 11742
rect 4794 11686 4880 11742
rect 4936 11686 5008 11742
rect 4668 11600 5008 11686
rect 4668 11544 4738 11600
rect 4794 11544 4880 11600
rect 4936 11544 5008 11600
rect 4668 11458 5008 11544
rect 4668 11402 4738 11458
rect 4794 11402 4880 11458
rect 4936 11402 5008 11458
rect 4668 11316 5008 11402
rect 4668 11260 4738 11316
rect 4794 11260 4880 11316
rect 4936 11260 5008 11316
rect 4668 11174 5008 11260
rect 4668 11118 4738 11174
rect 4794 11118 4880 11174
rect 4936 11118 5008 11174
rect 4668 11032 5008 11118
rect 4668 10976 4738 11032
rect 4794 10976 4880 11032
rect 4936 10976 5008 11032
rect 4668 10890 5008 10976
rect 4668 10834 4738 10890
rect 4794 10834 4880 10890
rect 4936 10834 5008 10890
rect 4668 10748 5008 10834
rect 4668 10692 4738 10748
rect 4794 10692 4880 10748
rect 4936 10692 5008 10748
rect 4668 10606 5008 10692
rect 4668 10550 4738 10606
rect 4794 10550 4880 10606
rect 4936 10550 5008 10606
rect 4668 10464 5008 10550
rect 4668 10408 4738 10464
rect 4794 10408 4880 10464
rect 4936 10408 5008 10464
rect 4668 10322 5008 10408
rect 4668 10266 4738 10322
rect 4794 10266 4880 10322
rect 4936 10266 5008 10322
rect 4668 10180 5008 10266
rect 4668 10124 4738 10180
rect 4794 10124 4880 10180
rect 4936 10124 5008 10180
rect 4668 10038 5008 10124
rect 4668 9982 4738 10038
rect 4794 9982 4880 10038
rect 4936 9982 5008 10038
rect 4668 9896 5008 9982
rect 4668 9840 4738 9896
rect 4794 9840 4880 9896
rect 4936 9840 5008 9896
rect 4668 9754 5008 9840
rect 4668 9698 4738 9754
rect 4794 9698 4880 9754
rect 4936 9698 5008 9754
rect 4668 9612 5008 9698
rect 4668 9556 4738 9612
rect 4794 9556 4880 9612
rect 4936 9556 5008 9612
rect 4668 9470 5008 9556
rect 4668 9414 4738 9470
rect 4794 9414 4880 9470
rect 4936 9414 5008 9470
rect 4668 9328 5008 9414
rect 4668 9272 4738 9328
rect 4794 9272 4880 9328
rect 4936 9272 5008 9328
rect 4668 9186 5008 9272
rect 4668 9130 4738 9186
rect 4794 9130 4880 9186
rect 4936 9130 5008 9186
rect 4668 9044 5008 9130
rect 4668 8988 4738 9044
rect 4794 8988 4880 9044
rect 4936 8988 5008 9044
rect 4668 8902 5008 8988
rect 4668 8846 4738 8902
rect 4794 8846 4880 8902
rect 4936 8846 5008 8902
rect 4668 8760 5008 8846
rect 4668 8704 4738 8760
rect 4794 8704 4880 8760
rect 4936 8704 5008 8760
rect 4668 8618 5008 8704
rect 4668 8562 4738 8618
rect 4794 8562 4880 8618
rect 4936 8562 5008 8618
rect 4668 8476 5008 8562
rect 4668 8420 4738 8476
rect 4794 8420 4880 8476
rect 4936 8420 5008 8476
rect 4668 8334 5008 8420
rect 4668 8278 4738 8334
rect 4794 8278 4880 8334
rect 4936 8278 5008 8334
rect 4668 8192 5008 8278
rect 4668 8136 4738 8192
rect 4794 8136 4880 8192
rect 4936 8136 5008 8192
rect 4668 8050 5008 8136
rect 4668 7994 4738 8050
rect 4794 7994 4880 8050
rect 4936 7994 5008 8050
rect 4668 7908 5008 7994
rect 4668 7852 4738 7908
rect 4794 7852 4880 7908
rect 4936 7852 5008 7908
rect 4668 7766 5008 7852
rect 4668 7710 4738 7766
rect 4794 7710 4880 7766
rect 4936 7710 5008 7766
rect 4668 7624 5008 7710
rect 4668 7568 4738 7624
rect 4794 7568 4880 7624
rect 4936 7568 5008 7624
rect 4668 7482 5008 7568
rect 4668 7426 4738 7482
rect 4794 7426 4880 7482
rect 4936 7426 5008 7482
rect 4668 7340 5008 7426
rect 4668 7284 4738 7340
rect 4794 7284 4880 7340
rect 4936 7284 5008 7340
rect 4668 7198 5008 7284
rect 4668 7142 4738 7198
rect 4794 7142 4880 7198
rect 4936 7142 5008 7198
rect 4668 7056 5008 7142
rect 4668 7000 4738 7056
rect 4794 7000 4880 7056
rect 4936 7000 5008 7056
rect 4668 6914 5008 7000
rect 4668 6858 4738 6914
rect 4794 6858 4880 6914
rect 4936 6858 5008 6914
rect 4668 6772 5008 6858
rect 4668 6716 4738 6772
rect 4794 6716 4880 6772
rect 4936 6716 5008 6772
rect 4668 6630 5008 6716
rect 4668 6574 4738 6630
rect 4794 6574 4880 6630
rect 4936 6574 5008 6630
rect 4668 6488 5008 6574
rect 4668 6432 4738 6488
rect 4794 6432 4880 6488
rect 4936 6432 5008 6488
rect 4668 6346 5008 6432
rect 4668 6290 4738 6346
rect 4794 6290 4880 6346
rect 4936 6290 5008 6346
rect 4668 6204 5008 6290
rect 4668 6148 4738 6204
rect 4794 6148 4880 6204
rect 4936 6148 5008 6204
rect 4668 6062 5008 6148
rect 4668 6006 4738 6062
rect 4794 6006 4880 6062
rect 4936 6006 5008 6062
rect 4668 5920 5008 6006
rect 4668 5864 4738 5920
rect 4794 5864 4880 5920
rect 4936 5864 5008 5920
rect 4668 5778 5008 5864
rect 4668 5722 4738 5778
rect 4794 5722 4880 5778
rect 4936 5722 5008 5778
rect 4668 5636 5008 5722
rect 4668 5580 4738 5636
rect 4794 5580 4880 5636
rect 4936 5580 5008 5636
rect 4668 5494 5008 5580
rect 4668 5438 4738 5494
rect 4794 5438 4880 5494
rect 4936 5438 5008 5494
rect 4668 5352 5008 5438
rect 4668 5296 4738 5352
rect 4794 5296 4880 5352
rect 4936 5296 5008 5352
rect 4668 5210 5008 5296
rect 4668 5154 4738 5210
rect 4794 5154 4880 5210
rect 4936 5154 5008 5210
rect 4668 5068 5008 5154
rect 4668 5012 4738 5068
rect 4794 5012 4880 5068
rect 4936 5012 5008 5068
rect 4668 4926 5008 5012
rect 4668 4870 4738 4926
rect 4794 4870 4880 4926
rect 4936 4870 5008 4926
rect 4668 4784 5008 4870
rect 4668 4728 4738 4784
rect 4794 4728 4880 4784
rect 4936 4728 5008 4784
rect 4668 4642 5008 4728
rect 4668 4586 4738 4642
rect 4794 4586 4880 4642
rect 4936 4586 5008 4642
rect 4668 4500 5008 4586
rect 4668 4444 4738 4500
rect 4794 4444 4880 4500
rect 4936 4444 5008 4500
rect 4668 4358 5008 4444
rect 4668 4302 4738 4358
rect 4794 4302 4880 4358
rect 4936 4302 5008 4358
rect 4668 4216 5008 4302
rect 4668 4160 4738 4216
rect 4794 4160 4880 4216
rect 4936 4160 5008 4216
rect 4668 4074 5008 4160
rect 4668 4018 4738 4074
rect 4794 4018 4880 4074
rect 4936 4018 5008 4074
rect 4668 3932 5008 4018
rect 4668 3876 4738 3932
rect 4794 3876 4880 3932
rect 4936 3876 5008 3932
rect 4668 3790 5008 3876
rect 4668 3734 4738 3790
rect 4794 3734 4880 3790
rect 4936 3734 5008 3790
rect 4668 3648 5008 3734
rect 4668 3592 4738 3648
rect 4794 3592 4880 3648
rect 4936 3592 5008 3648
rect 4668 3506 5008 3592
rect 4668 3450 4738 3506
rect 4794 3450 4880 3506
rect 4936 3450 5008 3506
rect 4668 3364 5008 3450
rect 4668 3308 4738 3364
rect 4794 3308 4880 3364
rect 4936 3308 5008 3364
rect 4668 3222 5008 3308
rect 4668 3166 4738 3222
rect 4794 3166 4880 3222
rect 4936 3166 5008 3222
rect 4668 3080 5008 3166
rect 4668 3024 4738 3080
rect 4794 3024 4880 3080
rect 4936 3024 5008 3080
rect 4668 2938 5008 3024
rect 4668 2882 4738 2938
rect 4794 2882 4880 2938
rect 4936 2882 5008 2938
rect 4668 2796 5008 2882
rect 4668 2740 4738 2796
rect 4794 2740 4880 2796
rect 4936 2740 5008 2796
rect 4668 2654 5008 2740
rect 4668 2598 4738 2654
rect 4794 2598 4880 2654
rect 4936 2598 5008 2654
rect 4668 2512 5008 2598
rect 4668 2456 4738 2512
rect 4794 2456 4880 2512
rect 4936 2456 5008 2512
rect 4668 2370 5008 2456
rect 4668 2314 4738 2370
rect 4794 2314 4880 2370
rect 4936 2314 5008 2370
rect 4668 2228 5008 2314
rect 4668 2172 4738 2228
rect 4794 2172 4880 2228
rect 4936 2172 5008 2228
rect 4668 2086 5008 2172
rect 4668 2030 4738 2086
rect 4794 2030 4880 2086
rect 4936 2030 5008 2086
rect 4668 1944 5008 2030
rect 4668 1888 4738 1944
rect 4794 1888 4880 1944
rect 4936 1888 5008 1944
rect 4668 1802 5008 1888
rect 4668 1746 4738 1802
rect 4794 1746 4880 1802
rect 4936 1746 5008 1802
rect 4668 1660 5008 1746
rect 4668 1604 4738 1660
rect 4794 1604 4880 1660
rect 4936 1604 5008 1660
rect 4668 1518 5008 1604
rect 4668 1462 4738 1518
rect 4794 1462 4880 1518
rect 4936 1462 5008 1518
rect 4668 1376 5008 1462
rect 4668 1320 4738 1376
rect 4794 1320 4880 1376
rect 4936 1320 5008 1376
rect 4668 1234 5008 1320
rect 4668 1178 4738 1234
rect 4794 1178 4880 1234
rect 4936 1178 5008 1234
rect 4668 1092 5008 1178
rect 4668 1036 4738 1092
rect 4794 1036 4880 1092
rect 4936 1036 5008 1092
rect 4668 950 5008 1036
rect 4668 894 4738 950
rect 4794 894 4880 950
rect 4936 894 5008 950
rect 4668 808 5008 894
rect 4668 752 4738 808
rect 4794 752 4880 808
rect 4936 752 5008 808
rect 4668 666 5008 752
rect 4668 610 4738 666
rect 4794 610 4880 666
rect 4936 610 5008 666
rect 4668 524 5008 610
rect 4668 468 4738 524
rect 4794 468 4880 524
rect 4936 468 5008 524
rect 4668 400 5008 468
rect 5068 12310 5408 12400
rect 5068 12254 5143 12310
rect 5199 12254 5285 12310
rect 5341 12254 5408 12310
rect 5068 12168 5408 12254
rect 5068 12112 5143 12168
rect 5199 12112 5285 12168
rect 5341 12112 5408 12168
rect 5068 12026 5408 12112
rect 5068 11970 5143 12026
rect 5199 11970 5285 12026
rect 5341 11970 5408 12026
rect 5068 11884 5408 11970
rect 5068 11828 5143 11884
rect 5199 11828 5285 11884
rect 5341 11828 5408 11884
rect 5068 11742 5408 11828
rect 5068 11686 5143 11742
rect 5199 11686 5285 11742
rect 5341 11686 5408 11742
rect 5068 11600 5408 11686
rect 5068 11544 5143 11600
rect 5199 11544 5285 11600
rect 5341 11544 5408 11600
rect 5068 11458 5408 11544
rect 5068 11402 5143 11458
rect 5199 11402 5285 11458
rect 5341 11402 5408 11458
rect 5068 11316 5408 11402
rect 5068 11260 5143 11316
rect 5199 11260 5285 11316
rect 5341 11260 5408 11316
rect 5068 11174 5408 11260
rect 5068 11118 5143 11174
rect 5199 11118 5285 11174
rect 5341 11118 5408 11174
rect 5068 11032 5408 11118
rect 5068 10976 5143 11032
rect 5199 10976 5285 11032
rect 5341 10976 5408 11032
rect 5068 10890 5408 10976
rect 5068 10834 5143 10890
rect 5199 10834 5285 10890
rect 5341 10834 5408 10890
rect 5068 10748 5408 10834
rect 5068 10692 5143 10748
rect 5199 10692 5285 10748
rect 5341 10692 5408 10748
rect 5068 10606 5408 10692
rect 5068 10550 5143 10606
rect 5199 10550 5285 10606
rect 5341 10550 5408 10606
rect 5068 10464 5408 10550
rect 5068 10408 5143 10464
rect 5199 10408 5285 10464
rect 5341 10408 5408 10464
rect 5068 10322 5408 10408
rect 5068 10266 5143 10322
rect 5199 10266 5285 10322
rect 5341 10266 5408 10322
rect 5068 10180 5408 10266
rect 5068 10124 5143 10180
rect 5199 10124 5285 10180
rect 5341 10124 5408 10180
rect 5068 10038 5408 10124
rect 5068 9982 5143 10038
rect 5199 9982 5285 10038
rect 5341 9982 5408 10038
rect 5068 9896 5408 9982
rect 5068 9840 5143 9896
rect 5199 9840 5285 9896
rect 5341 9840 5408 9896
rect 5068 9754 5408 9840
rect 5068 9698 5143 9754
rect 5199 9698 5285 9754
rect 5341 9698 5408 9754
rect 5068 9612 5408 9698
rect 5068 9556 5143 9612
rect 5199 9556 5285 9612
rect 5341 9556 5408 9612
rect 5068 9470 5408 9556
rect 5068 9414 5143 9470
rect 5199 9414 5285 9470
rect 5341 9414 5408 9470
rect 5068 9328 5408 9414
rect 5068 9272 5143 9328
rect 5199 9272 5285 9328
rect 5341 9272 5408 9328
rect 5068 9186 5408 9272
rect 5068 9130 5143 9186
rect 5199 9130 5285 9186
rect 5341 9130 5408 9186
rect 5068 9044 5408 9130
rect 5068 8988 5143 9044
rect 5199 8988 5285 9044
rect 5341 8988 5408 9044
rect 5068 8902 5408 8988
rect 5068 8846 5143 8902
rect 5199 8846 5285 8902
rect 5341 8846 5408 8902
rect 5068 8760 5408 8846
rect 5068 8704 5143 8760
rect 5199 8704 5285 8760
rect 5341 8704 5408 8760
rect 5068 8618 5408 8704
rect 5068 8562 5143 8618
rect 5199 8562 5285 8618
rect 5341 8562 5408 8618
rect 5068 8476 5408 8562
rect 5068 8420 5143 8476
rect 5199 8420 5285 8476
rect 5341 8420 5408 8476
rect 5068 8334 5408 8420
rect 5068 8278 5143 8334
rect 5199 8278 5285 8334
rect 5341 8278 5408 8334
rect 5068 8192 5408 8278
rect 5068 8136 5143 8192
rect 5199 8136 5285 8192
rect 5341 8136 5408 8192
rect 5068 8050 5408 8136
rect 5068 7994 5143 8050
rect 5199 7994 5285 8050
rect 5341 7994 5408 8050
rect 5068 7908 5408 7994
rect 5068 7852 5143 7908
rect 5199 7852 5285 7908
rect 5341 7852 5408 7908
rect 5068 7766 5408 7852
rect 5068 7710 5143 7766
rect 5199 7710 5285 7766
rect 5341 7710 5408 7766
rect 5068 7624 5408 7710
rect 5068 7568 5143 7624
rect 5199 7568 5285 7624
rect 5341 7568 5408 7624
rect 5068 7482 5408 7568
rect 5068 7426 5143 7482
rect 5199 7426 5285 7482
rect 5341 7426 5408 7482
rect 5068 7340 5408 7426
rect 5068 7284 5143 7340
rect 5199 7284 5285 7340
rect 5341 7284 5408 7340
rect 5068 7198 5408 7284
rect 5068 7142 5143 7198
rect 5199 7142 5285 7198
rect 5341 7142 5408 7198
rect 5068 7056 5408 7142
rect 5068 7000 5143 7056
rect 5199 7000 5285 7056
rect 5341 7000 5408 7056
rect 5068 6914 5408 7000
rect 5068 6858 5143 6914
rect 5199 6858 5285 6914
rect 5341 6858 5408 6914
rect 5068 6772 5408 6858
rect 5068 6716 5143 6772
rect 5199 6716 5285 6772
rect 5341 6716 5408 6772
rect 5068 6630 5408 6716
rect 5068 6574 5143 6630
rect 5199 6574 5285 6630
rect 5341 6574 5408 6630
rect 5068 6488 5408 6574
rect 5068 6432 5143 6488
rect 5199 6432 5285 6488
rect 5341 6432 5408 6488
rect 5068 6346 5408 6432
rect 5068 6290 5143 6346
rect 5199 6290 5285 6346
rect 5341 6290 5408 6346
rect 5068 6204 5408 6290
rect 5068 6148 5143 6204
rect 5199 6148 5285 6204
rect 5341 6148 5408 6204
rect 5068 6062 5408 6148
rect 5068 6006 5143 6062
rect 5199 6006 5285 6062
rect 5341 6006 5408 6062
rect 5068 5920 5408 6006
rect 5068 5864 5143 5920
rect 5199 5864 5285 5920
rect 5341 5864 5408 5920
rect 5068 5778 5408 5864
rect 5068 5722 5143 5778
rect 5199 5722 5285 5778
rect 5341 5722 5408 5778
rect 5068 5636 5408 5722
rect 5068 5580 5143 5636
rect 5199 5580 5285 5636
rect 5341 5580 5408 5636
rect 5068 5494 5408 5580
rect 5068 5438 5143 5494
rect 5199 5438 5285 5494
rect 5341 5438 5408 5494
rect 5068 5352 5408 5438
rect 5068 5296 5143 5352
rect 5199 5296 5285 5352
rect 5341 5296 5408 5352
rect 5068 5210 5408 5296
rect 5068 5154 5143 5210
rect 5199 5154 5285 5210
rect 5341 5154 5408 5210
rect 5068 5068 5408 5154
rect 5068 5012 5143 5068
rect 5199 5012 5285 5068
rect 5341 5012 5408 5068
rect 5068 4926 5408 5012
rect 5068 4870 5143 4926
rect 5199 4870 5285 4926
rect 5341 4870 5408 4926
rect 5068 4784 5408 4870
rect 5068 4728 5143 4784
rect 5199 4728 5285 4784
rect 5341 4728 5408 4784
rect 5068 4642 5408 4728
rect 5068 4586 5143 4642
rect 5199 4586 5285 4642
rect 5341 4586 5408 4642
rect 5068 4500 5408 4586
rect 5068 4444 5143 4500
rect 5199 4444 5285 4500
rect 5341 4444 5408 4500
rect 5068 4358 5408 4444
rect 5068 4302 5143 4358
rect 5199 4302 5285 4358
rect 5341 4302 5408 4358
rect 5068 4216 5408 4302
rect 5068 4160 5143 4216
rect 5199 4160 5285 4216
rect 5341 4160 5408 4216
rect 5068 4074 5408 4160
rect 5068 4018 5143 4074
rect 5199 4018 5285 4074
rect 5341 4018 5408 4074
rect 5068 3932 5408 4018
rect 5068 3876 5143 3932
rect 5199 3876 5285 3932
rect 5341 3876 5408 3932
rect 5068 3790 5408 3876
rect 5068 3734 5143 3790
rect 5199 3734 5285 3790
rect 5341 3734 5408 3790
rect 5068 3648 5408 3734
rect 5068 3592 5143 3648
rect 5199 3592 5285 3648
rect 5341 3592 5408 3648
rect 5068 3506 5408 3592
rect 5068 3450 5143 3506
rect 5199 3450 5285 3506
rect 5341 3450 5408 3506
rect 5068 3364 5408 3450
rect 5068 3308 5143 3364
rect 5199 3308 5285 3364
rect 5341 3308 5408 3364
rect 5068 3222 5408 3308
rect 5068 3166 5143 3222
rect 5199 3166 5285 3222
rect 5341 3166 5408 3222
rect 5068 3080 5408 3166
rect 5068 3024 5143 3080
rect 5199 3024 5285 3080
rect 5341 3024 5408 3080
rect 5068 2938 5408 3024
rect 5068 2882 5143 2938
rect 5199 2882 5285 2938
rect 5341 2882 5408 2938
rect 5068 2796 5408 2882
rect 5068 2740 5143 2796
rect 5199 2740 5285 2796
rect 5341 2740 5408 2796
rect 5068 2654 5408 2740
rect 5068 2598 5143 2654
rect 5199 2598 5285 2654
rect 5341 2598 5408 2654
rect 5068 2512 5408 2598
rect 5068 2456 5143 2512
rect 5199 2456 5285 2512
rect 5341 2456 5408 2512
rect 5068 2370 5408 2456
rect 5068 2314 5143 2370
rect 5199 2314 5285 2370
rect 5341 2314 5408 2370
rect 5068 2228 5408 2314
rect 5068 2172 5143 2228
rect 5199 2172 5285 2228
rect 5341 2172 5408 2228
rect 5068 2086 5408 2172
rect 5068 2030 5143 2086
rect 5199 2030 5285 2086
rect 5341 2030 5408 2086
rect 5068 1944 5408 2030
rect 5068 1888 5143 1944
rect 5199 1888 5285 1944
rect 5341 1888 5408 1944
rect 5068 1802 5408 1888
rect 5068 1746 5143 1802
rect 5199 1746 5285 1802
rect 5341 1746 5408 1802
rect 5068 1660 5408 1746
rect 5068 1604 5143 1660
rect 5199 1604 5285 1660
rect 5341 1604 5408 1660
rect 5068 1518 5408 1604
rect 5068 1462 5143 1518
rect 5199 1462 5285 1518
rect 5341 1462 5408 1518
rect 5068 1376 5408 1462
rect 5068 1320 5143 1376
rect 5199 1320 5285 1376
rect 5341 1320 5408 1376
rect 5068 1234 5408 1320
rect 5068 1178 5143 1234
rect 5199 1178 5285 1234
rect 5341 1178 5408 1234
rect 5068 1092 5408 1178
rect 5068 1036 5143 1092
rect 5199 1036 5285 1092
rect 5341 1036 5408 1092
rect 5068 950 5408 1036
rect 5068 894 5143 950
rect 5199 894 5285 950
rect 5341 894 5408 950
rect 5068 808 5408 894
rect 5068 752 5143 808
rect 5199 752 5285 808
rect 5341 752 5408 808
rect 5068 666 5408 752
rect 5068 610 5143 666
rect 5199 610 5285 666
rect 5341 610 5408 666
rect 5068 524 5408 610
rect 5068 468 5143 524
rect 5199 468 5285 524
rect 5341 468 5408 524
rect 5068 400 5408 468
rect 5468 12310 5808 12400
rect 5468 12254 5540 12310
rect 5596 12254 5682 12310
rect 5738 12254 5808 12310
rect 5468 12168 5808 12254
rect 5468 12112 5540 12168
rect 5596 12112 5682 12168
rect 5738 12112 5808 12168
rect 5468 12026 5808 12112
rect 5468 11970 5540 12026
rect 5596 11970 5682 12026
rect 5738 11970 5808 12026
rect 5468 11884 5808 11970
rect 5468 11828 5540 11884
rect 5596 11828 5682 11884
rect 5738 11828 5808 11884
rect 5468 11742 5808 11828
rect 5468 11686 5540 11742
rect 5596 11686 5682 11742
rect 5738 11686 5808 11742
rect 5468 11600 5808 11686
rect 5468 11544 5540 11600
rect 5596 11544 5682 11600
rect 5738 11544 5808 11600
rect 5468 11458 5808 11544
rect 5468 11402 5540 11458
rect 5596 11402 5682 11458
rect 5738 11402 5808 11458
rect 5468 11316 5808 11402
rect 5468 11260 5540 11316
rect 5596 11260 5682 11316
rect 5738 11260 5808 11316
rect 5468 11174 5808 11260
rect 5468 11118 5540 11174
rect 5596 11118 5682 11174
rect 5738 11118 5808 11174
rect 5468 11032 5808 11118
rect 5468 10976 5540 11032
rect 5596 10976 5682 11032
rect 5738 10976 5808 11032
rect 5468 10890 5808 10976
rect 5468 10834 5540 10890
rect 5596 10834 5682 10890
rect 5738 10834 5808 10890
rect 5468 10748 5808 10834
rect 5468 10692 5540 10748
rect 5596 10692 5682 10748
rect 5738 10692 5808 10748
rect 5468 10606 5808 10692
rect 5468 10550 5540 10606
rect 5596 10550 5682 10606
rect 5738 10550 5808 10606
rect 5468 10464 5808 10550
rect 5468 10408 5540 10464
rect 5596 10408 5682 10464
rect 5738 10408 5808 10464
rect 5468 10322 5808 10408
rect 5468 10266 5540 10322
rect 5596 10266 5682 10322
rect 5738 10266 5808 10322
rect 5468 10180 5808 10266
rect 5468 10124 5540 10180
rect 5596 10124 5682 10180
rect 5738 10124 5808 10180
rect 5468 10038 5808 10124
rect 5468 9982 5540 10038
rect 5596 9982 5682 10038
rect 5738 9982 5808 10038
rect 5468 9896 5808 9982
rect 5468 9840 5540 9896
rect 5596 9840 5682 9896
rect 5738 9840 5808 9896
rect 5468 9754 5808 9840
rect 5468 9698 5540 9754
rect 5596 9698 5682 9754
rect 5738 9698 5808 9754
rect 5468 9612 5808 9698
rect 5468 9556 5540 9612
rect 5596 9556 5682 9612
rect 5738 9556 5808 9612
rect 5468 9470 5808 9556
rect 5468 9414 5540 9470
rect 5596 9414 5682 9470
rect 5738 9414 5808 9470
rect 5468 9328 5808 9414
rect 5468 9272 5540 9328
rect 5596 9272 5682 9328
rect 5738 9272 5808 9328
rect 5468 9186 5808 9272
rect 5468 9130 5540 9186
rect 5596 9130 5682 9186
rect 5738 9130 5808 9186
rect 5468 9044 5808 9130
rect 5468 8988 5540 9044
rect 5596 8988 5682 9044
rect 5738 8988 5808 9044
rect 5468 8902 5808 8988
rect 5468 8846 5540 8902
rect 5596 8846 5682 8902
rect 5738 8846 5808 8902
rect 5468 8760 5808 8846
rect 5468 8704 5540 8760
rect 5596 8704 5682 8760
rect 5738 8704 5808 8760
rect 5468 8618 5808 8704
rect 5468 8562 5540 8618
rect 5596 8562 5682 8618
rect 5738 8562 5808 8618
rect 5468 8476 5808 8562
rect 5468 8420 5540 8476
rect 5596 8420 5682 8476
rect 5738 8420 5808 8476
rect 5468 8334 5808 8420
rect 5468 8278 5540 8334
rect 5596 8278 5682 8334
rect 5738 8278 5808 8334
rect 5468 8192 5808 8278
rect 5468 8136 5540 8192
rect 5596 8136 5682 8192
rect 5738 8136 5808 8192
rect 5468 8050 5808 8136
rect 5468 7994 5540 8050
rect 5596 7994 5682 8050
rect 5738 7994 5808 8050
rect 5468 7908 5808 7994
rect 5468 7852 5540 7908
rect 5596 7852 5682 7908
rect 5738 7852 5808 7908
rect 5468 7766 5808 7852
rect 5468 7710 5540 7766
rect 5596 7710 5682 7766
rect 5738 7710 5808 7766
rect 5468 7624 5808 7710
rect 5468 7568 5540 7624
rect 5596 7568 5682 7624
rect 5738 7568 5808 7624
rect 5468 7482 5808 7568
rect 5468 7426 5540 7482
rect 5596 7426 5682 7482
rect 5738 7426 5808 7482
rect 5468 7340 5808 7426
rect 5468 7284 5540 7340
rect 5596 7284 5682 7340
rect 5738 7284 5808 7340
rect 5468 7198 5808 7284
rect 5468 7142 5540 7198
rect 5596 7142 5682 7198
rect 5738 7142 5808 7198
rect 5468 7056 5808 7142
rect 5468 7000 5540 7056
rect 5596 7000 5682 7056
rect 5738 7000 5808 7056
rect 5468 6914 5808 7000
rect 5468 6858 5540 6914
rect 5596 6858 5682 6914
rect 5738 6858 5808 6914
rect 5468 6772 5808 6858
rect 5468 6716 5540 6772
rect 5596 6716 5682 6772
rect 5738 6716 5808 6772
rect 5468 6630 5808 6716
rect 5468 6574 5540 6630
rect 5596 6574 5682 6630
rect 5738 6574 5808 6630
rect 5468 6488 5808 6574
rect 5468 6432 5540 6488
rect 5596 6432 5682 6488
rect 5738 6432 5808 6488
rect 5468 6346 5808 6432
rect 5468 6290 5540 6346
rect 5596 6290 5682 6346
rect 5738 6290 5808 6346
rect 5468 6204 5808 6290
rect 5468 6148 5540 6204
rect 5596 6148 5682 6204
rect 5738 6148 5808 6204
rect 5468 6062 5808 6148
rect 5468 6006 5540 6062
rect 5596 6006 5682 6062
rect 5738 6006 5808 6062
rect 5468 5920 5808 6006
rect 5468 5864 5540 5920
rect 5596 5864 5682 5920
rect 5738 5864 5808 5920
rect 5468 5778 5808 5864
rect 5468 5722 5540 5778
rect 5596 5722 5682 5778
rect 5738 5722 5808 5778
rect 5468 5636 5808 5722
rect 5468 5580 5540 5636
rect 5596 5580 5682 5636
rect 5738 5580 5808 5636
rect 5468 5494 5808 5580
rect 5468 5438 5540 5494
rect 5596 5438 5682 5494
rect 5738 5438 5808 5494
rect 5468 5352 5808 5438
rect 5468 5296 5540 5352
rect 5596 5296 5682 5352
rect 5738 5296 5808 5352
rect 5468 5210 5808 5296
rect 5468 5154 5540 5210
rect 5596 5154 5682 5210
rect 5738 5154 5808 5210
rect 5468 5068 5808 5154
rect 5468 5012 5540 5068
rect 5596 5012 5682 5068
rect 5738 5012 5808 5068
rect 5468 4926 5808 5012
rect 5468 4870 5540 4926
rect 5596 4870 5682 4926
rect 5738 4870 5808 4926
rect 5468 4784 5808 4870
rect 5468 4728 5540 4784
rect 5596 4728 5682 4784
rect 5738 4728 5808 4784
rect 5468 4642 5808 4728
rect 5468 4586 5540 4642
rect 5596 4586 5682 4642
rect 5738 4586 5808 4642
rect 5468 4500 5808 4586
rect 5468 4444 5540 4500
rect 5596 4444 5682 4500
rect 5738 4444 5808 4500
rect 5468 4358 5808 4444
rect 5468 4302 5540 4358
rect 5596 4302 5682 4358
rect 5738 4302 5808 4358
rect 5468 4216 5808 4302
rect 5468 4160 5540 4216
rect 5596 4160 5682 4216
rect 5738 4160 5808 4216
rect 5468 4074 5808 4160
rect 5468 4018 5540 4074
rect 5596 4018 5682 4074
rect 5738 4018 5808 4074
rect 5468 3932 5808 4018
rect 5468 3876 5540 3932
rect 5596 3876 5682 3932
rect 5738 3876 5808 3932
rect 5468 3790 5808 3876
rect 5468 3734 5540 3790
rect 5596 3734 5682 3790
rect 5738 3734 5808 3790
rect 5468 3648 5808 3734
rect 5468 3592 5540 3648
rect 5596 3592 5682 3648
rect 5738 3592 5808 3648
rect 5468 3506 5808 3592
rect 5468 3450 5540 3506
rect 5596 3450 5682 3506
rect 5738 3450 5808 3506
rect 5468 3364 5808 3450
rect 5468 3308 5540 3364
rect 5596 3308 5682 3364
rect 5738 3308 5808 3364
rect 5468 3222 5808 3308
rect 5468 3166 5540 3222
rect 5596 3166 5682 3222
rect 5738 3166 5808 3222
rect 5468 3080 5808 3166
rect 5468 3024 5540 3080
rect 5596 3024 5682 3080
rect 5738 3024 5808 3080
rect 5468 2938 5808 3024
rect 5468 2882 5540 2938
rect 5596 2882 5682 2938
rect 5738 2882 5808 2938
rect 5468 2796 5808 2882
rect 5468 2740 5540 2796
rect 5596 2740 5682 2796
rect 5738 2740 5808 2796
rect 5468 2654 5808 2740
rect 5468 2598 5540 2654
rect 5596 2598 5682 2654
rect 5738 2598 5808 2654
rect 5468 2512 5808 2598
rect 5468 2456 5540 2512
rect 5596 2456 5682 2512
rect 5738 2456 5808 2512
rect 5468 2370 5808 2456
rect 5468 2314 5540 2370
rect 5596 2314 5682 2370
rect 5738 2314 5808 2370
rect 5468 2228 5808 2314
rect 5468 2172 5540 2228
rect 5596 2172 5682 2228
rect 5738 2172 5808 2228
rect 5468 2086 5808 2172
rect 5468 2030 5540 2086
rect 5596 2030 5682 2086
rect 5738 2030 5808 2086
rect 5468 1944 5808 2030
rect 5468 1888 5540 1944
rect 5596 1888 5682 1944
rect 5738 1888 5808 1944
rect 5468 1802 5808 1888
rect 5468 1746 5540 1802
rect 5596 1746 5682 1802
rect 5738 1746 5808 1802
rect 5468 1660 5808 1746
rect 5468 1604 5540 1660
rect 5596 1604 5682 1660
rect 5738 1604 5808 1660
rect 5468 1518 5808 1604
rect 5468 1462 5540 1518
rect 5596 1462 5682 1518
rect 5738 1462 5808 1518
rect 5468 1376 5808 1462
rect 5468 1320 5540 1376
rect 5596 1320 5682 1376
rect 5738 1320 5808 1376
rect 5468 1234 5808 1320
rect 5468 1178 5540 1234
rect 5596 1178 5682 1234
rect 5738 1178 5808 1234
rect 5468 1092 5808 1178
rect 5468 1036 5540 1092
rect 5596 1036 5682 1092
rect 5738 1036 5808 1092
rect 5468 950 5808 1036
rect 5468 894 5540 950
rect 5596 894 5682 950
rect 5738 894 5808 950
rect 5468 808 5808 894
rect 5468 752 5540 808
rect 5596 752 5682 808
rect 5738 752 5808 808
rect 5468 666 5808 752
rect 5468 610 5540 666
rect 5596 610 5682 666
rect 5738 610 5808 666
rect 5468 524 5808 610
rect 5468 468 5540 524
rect 5596 468 5682 524
rect 5738 468 5808 524
rect 5468 400 5808 468
rect 5868 12310 6208 12400
rect 5868 12254 5937 12310
rect 5993 12254 6079 12310
rect 6135 12254 6208 12310
rect 5868 12168 6208 12254
rect 5868 12112 5937 12168
rect 5993 12112 6079 12168
rect 6135 12112 6208 12168
rect 5868 12026 6208 12112
rect 5868 11970 5937 12026
rect 5993 11970 6079 12026
rect 6135 11970 6208 12026
rect 5868 11884 6208 11970
rect 5868 11828 5937 11884
rect 5993 11828 6079 11884
rect 6135 11828 6208 11884
rect 5868 11742 6208 11828
rect 5868 11686 5937 11742
rect 5993 11686 6079 11742
rect 6135 11686 6208 11742
rect 5868 11600 6208 11686
rect 5868 11544 5937 11600
rect 5993 11544 6079 11600
rect 6135 11544 6208 11600
rect 5868 11458 6208 11544
rect 5868 11402 5937 11458
rect 5993 11402 6079 11458
rect 6135 11402 6208 11458
rect 5868 11316 6208 11402
rect 5868 11260 5937 11316
rect 5993 11260 6079 11316
rect 6135 11260 6208 11316
rect 5868 11174 6208 11260
rect 5868 11118 5937 11174
rect 5993 11118 6079 11174
rect 6135 11118 6208 11174
rect 5868 11032 6208 11118
rect 5868 10976 5937 11032
rect 5993 10976 6079 11032
rect 6135 10976 6208 11032
rect 5868 10890 6208 10976
rect 5868 10834 5937 10890
rect 5993 10834 6079 10890
rect 6135 10834 6208 10890
rect 5868 10748 6208 10834
rect 5868 10692 5937 10748
rect 5993 10692 6079 10748
rect 6135 10692 6208 10748
rect 5868 10606 6208 10692
rect 5868 10550 5937 10606
rect 5993 10550 6079 10606
rect 6135 10550 6208 10606
rect 5868 10464 6208 10550
rect 5868 10408 5937 10464
rect 5993 10408 6079 10464
rect 6135 10408 6208 10464
rect 5868 10322 6208 10408
rect 5868 10266 5937 10322
rect 5993 10266 6079 10322
rect 6135 10266 6208 10322
rect 5868 10180 6208 10266
rect 5868 10124 5937 10180
rect 5993 10124 6079 10180
rect 6135 10124 6208 10180
rect 5868 10038 6208 10124
rect 5868 9982 5937 10038
rect 5993 9982 6079 10038
rect 6135 9982 6208 10038
rect 5868 9896 6208 9982
rect 5868 9840 5937 9896
rect 5993 9840 6079 9896
rect 6135 9840 6208 9896
rect 5868 9754 6208 9840
rect 5868 9698 5937 9754
rect 5993 9698 6079 9754
rect 6135 9698 6208 9754
rect 5868 9612 6208 9698
rect 5868 9556 5937 9612
rect 5993 9556 6079 9612
rect 6135 9556 6208 9612
rect 5868 9470 6208 9556
rect 5868 9414 5937 9470
rect 5993 9414 6079 9470
rect 6135 9414 6208 9470
rect 5868 9328 6208 9414
rect 5868 9272 5937 9328
rect 5993 9272 6079 9328
rect 6135 9272 6208 9328
rect 5868 9186 6208 9272
rect 5868 9130 5937 9186
rect 5993 9130 6079 9186
rect 6135 9130 6208 9186
rect 5868 9044 6208 9130
rect 5868 8988 5937 9044
rect 5993 8988 6079 9044
rect 6135 8988 6208 9044
rect 5868 8902 6208 8988
rect 5868 8846 5937 8902
rect 5993 8846 6079 8902
rect 6135 8846 6208 8902
rect 5868 8760 6208 8846
rect 5868 8704 5937 8760
rect 5993 8704 6079 8760
rect 6135 8704 6208 8760
rect 5868 8618 6208 8704
rect 5868 8562 5937 8618
rect 5993 8562 6079 8618
rect 6135 8562 6208 8618
rect 5868 8476 6208 8562
rect 5868 8420 5937 8476
rect 5993 8420 6079 8476
rect 6135 8420 6208 8476
rect 5868 8334 6208 8420
rect 5868 8278 5937 8334
rect 5993 8278 6079 8334
rect 6135 8278 6208 8334
rect 5868 8192 6208 8278
rect 5868 8136 5937 8192
rect 5993 8136 6079 8192
rect 6135 8136 6208 8192
rect 5868 8050 6208 8136
rect 5868 7994 5937 8050
rect 5993 7994 6079 8050
rect 6135 7994 6208 8050
rect 5868 7908 6208 7994
rect 5868 7852 5937 7908
rect 5993 7852 6079 7908
rect 6135 7852 6208 7908
rect 5868 7766 6208 7852
rect 5868 7710 5937 7766
rect 5993 7710 6079 7766
rect 6135 7710 6208 7766
rect 5868 7624 6208 7710
rect 5868 7568 5937 7624
rect 5993 7568 6079 7624
rect 6135 7568 6208 7624
rect 5868 7482 6208 7568
rect 5868 7426 5937 7482
rect 5993 7426 6079 7482
rect 6135 7426 6208 7482
rect 5868 7340 6208 7426
rect 5868 7284 5937 7340
rect 5993 7284 6079 7340
rect 6135 7284 6208 7340
rect 5868 7198 6208 7284
rect 5868 7142 5937 7198
rect 5993 7142 6079 7198
rect 6135 7142 6208 7198
rect 5868 7056 6208 7142
rect 5868 7000 5937 7056
rect 5993 7000 6079 7056
rect 6135 7000 6208 7056
rect 5868 6914 6208 7000
rect 5868 6858 5937 6914
rect 5993 6858 6079 6914
rect 6135 6858 6208 6914
rect 5868 6772 6208 6858
rect 5868 6716 5937 6772
rect 5993 6716 6079 6772
rect 6135 6716 6208 6772
rect 5868 6630 6208 6716
rect 5868 6574 5937 6630
rect 5993 6574 6079 6630
rect 6135 6574 6208 6630
rect 5868 6488 6208 6574
rect 5868 6432 5937 6488
rect 5993 6432 6079 6488
rect 6135 6432 6208 6488
rect 5868 6346 6208 6432
rect 5868 6290 5937 6346
rect 5993 6290 6079 6346
rect 6135 6290 6208 6346
rect 5868 6204 6208 6290
rect 5868 6148 5937 6204
rect 5993 6148 6079 6204
rect 6135 6148 6208 6204
rect 5868 6062 6208 6148
rect 5868 6006 5937 6062
rect 5993 6006 6079 6062
rect 6135 6006 6208 6062
rect 5868 5920 6208 6006
rect 5868 5864 5937 5920
rect 5993 5864 6079 5920
rect 6135 5864 6208 5920
rect 5868 5778 6208 5864
rect 5868 5722 5937 5778
rect 5993 5722 6079 5778
rect 6135 5722 6208 5778
rect 5868 5636 6208 5722
rect 5868 5580 5937 5636
rect 5993 5580 6079 5636
rect 6135 5580 6208 5636
rect 5868 5494 6208 5580
rect 5868 5438 5937 5494
rect 5993 5438 6079 5494
rect 6135 5438 6208 5494
rect 5868 5352 6208 5438
rect 5868 5296 5937 5352
rect 5993 5296 6079 5352
rect 6135 5296 6208 5352
rect 5868 5210 6208 5296
rect 5868 5154 5937 5210
rect 5993 5154 6079 5210
rect 6135 5154 6208 5210
rect 5868 5068 6208 5154
rect 5868 5012 5937 5068
rect 5993 5012 6079 5068
rect 6135 5012 6208 5068
rect 5868 4926 6208 5012
rect 5868 4870 5937 4926
rect 5993 4870 6079 4926
rect 6135 4870 6208 4926
rect 5868 4784 6208 4870
rect 5868 4728 5937 4784
rect 5993 4728 6079 4784
rect 6135 4728 6208 4784
rect 5868 4642 6208 4728
rect 5868 4586 5937 4642
rect 5993 4586 6079 4642
rect 6135 4586 6208 4642
rect 5868 4500 6208 4586
rect 5868 4444 5937 4500
rect 5993 4444 6079 4500
rect 6135 4444 6208 4500
rect 5868 4358 6208 4444
rect 5868 4302 5937 4358
rect 5993 4302 6079 4358
rect 6135 4302 6208 4358
rect 5868 4216 6208 4302
rect 5868 4160 5937 4216
rect 5993 4160 6079 4216
rect 6135 4160 6208 4216
rect 5868 4074 6208 4160
rect 5868 4018 5937 4074
rect 5993 4018 6079 4074
rect 6135 4018 6208 4074
rect 5868 3932 6208 4018
rect 5868 3876 5937 3932
rect 5993 3876 6079 3932
rect 6135 3876 6208 3932
rect 5868 3790 6208 3876
rect 5868 3734 5937 3790
rect 5993 3734 6079 3790
rect 6135 3734 6208 3790
rect 5868 3648 6208 3734
rect 5868 3592 5937 3648
rect 5993 3592 6079 3648
rect 6135 3592 6208 3648
rect 5868 3506 6208 3592
rect 5868 3450 5937 3506
rect 5993 3450 6079 3506
rect 6135 3450 6208 3506
rect 5868 3364 6208 3450
rect 5868 3308 5937 3364
rect 5993 3308 6079 3364
rect 6135 3308 6208 3364
rect 5868 3222 6208 3308
rect 5868 3166 5937 3222
rect 5993 3166 6079 3222
rect 6135 3166 6208 3222
rect 5868 3080 6208 3166
rect 5868 3024 5937 3080
rect 5993 3024 6079 3080
rect 6135 3024 6208 3080
rect 5868 2938 6208 3024
rect 5868 2882 5937 2938
rect 5993 2882 6079 2938
rect 6135 2882 6208 2938
rect 5868 2796 6208 2882
rect 5868 2740 5937 2796
rect 5993 2740 6079 2796
rect 6135 2740 6208 2796
rect 5868 2654 6208 2740
rect 5868 2598 5937 2654
rect 5993 2598 6079 2654
rect 6135 2598 6208 2654
rect 5868 2512 6208 2598
rect 5868 2456 5937 2512
rect 5993 2456 6079 2512
rect 6135 2456 6208 2512
rect 5868 2370 6208 2456
rect 5868 2314 5937 2370
rect 5993 2314 6079 2370
rect 6135 2314 6208 2370
rect 5868 2228 6208 2314
rect 5868 2172 5937 2228
rect 5993 2172 6079 2228
rect 6135 2172 6208 2228
rect 5868 2086 6208 2172
rect 5868 2030 5937 2086
rect 5993 2030 6079 2086
rect 6135 2030 6208 2086
rect 5868 1944 6208 2030
rect 5868 1888 5937 1944
rect 5993 1888 6079 1944
rect 6135 1888 6208 1944
rect 5868 1802 6208 1888
rect 5868 1746 5937 1802
rect 5993 1746 6079 1802
rect 6135 1746 6208 1802
rect 5868 1660 6208 1746
rect 5868 1604 5937 1660
rect 5993 1604 6079 1660
rect 6135 1604 6208 1660
rect 5868 1518 6208 1604
rect 5868 1462 5937 1518
rect 5993 1462 6079 1518
rect 6135 1462 6208 1518
rect 5868 1376 6208 1462
rect 5868 1320 5937 1376
rect 5993 1320 6079 1376
rect 6135 1320 6208 1376
rect 5868 1234 6208 1320
rect 5868 1178 5937 1234
rect 5993 1178 6079 1234
rect 6135 1178 6208 1234
rect 5868 1092 6208 1178
rect 5868 1036 5937 1092
rect 5993 1036 6079 1092
rect 6135 1036 6208 1092
rect 5868 950 6208 1036
rect 5868 894 5937 950
rect 5993 894 6079 950
rect 6135 894 6208 950
rect 5868 808 6208 894
rect 5868 752 5937 808
rect 5993 752 6079 808
rect 6135 752 6208 808
rect 5868 666 6208 752
rect 5868 610 5937 666
rect 5993 610 6079 666
rect 6135 610 6208 666
rect 5868 524 6208 610
rect 5868 468 5937 524
rect 5993 468 6079 524
rect 6135 468 6208 524
rect 5868 400 6208 468
rect 6268 12310 6608 12400
rect 6268 12254 6340 12310
rect 6396 12254 6482 12310
rect 6538 12254 6608 12310
rect 6268 12168 6608 12254
rect 6268 12112 6340 12168
rect 6396 12112 6482 12168
rect 6538 12112 6608 12168
rect 6268 12026 6608 12112
rect 6268 11970 6340 12026
rect 6396 11970 6482 12026
rect 6538 11970 6608 12026
rect 6268 11884 6608 11970
rect 6268 11828 6340 11884
rect 6396 11828 6482 11884
rect 6538 11828 6608 11884
rect 6268 11742 6608 11828
rect 6268 11686 6340 11742
rect 6396 11686 6482 11742
rect 6538 11686 6608 11742
rect 6268 11600 6608 11686
rect 6268 11544 6340 11600
rect 6396 11544 6482 11600
rect 6538 11544 6608 11600
rect 6268 11458 6608 11544
rect 6268 11402 6340 11458
rect 6396 11402 6482 11458
rect 6538 11402 6608 11458
rect 6268 11316 6608 11402
rect 6268 11260 6340 11316
rect 6396 11260 6482 11316
rect 6538 11260 6608 11316
rect 6268 11174 6608 11260
rect 6268 11118 6340 11174
rect 6396 11118 6482 11174
rect 6538 11118 6608 11174
rect 6268 11032 6608 11118
rect 6268 10976 6340 11032
rect 6396 10976 6482 11032
rect 6538 10976 6608 11032
rect 6268 10890 6608 10976
rect 6268 10834 6340 10890
rect 6396 10834 6482 10890
rect 6538 10834 6608 10890
rect 6268 10748 6608 10834
rect 6268 10692 6340 10748
rect 6396 10692 6482 10748
rect 6538 10692 6608 10748
rect 6268 10606 6608 10692
rect 6268 10550 6340 10606
rect 6396 10550 6482 10606
rect 6538 10550 6608 10606
rect 6268 10464 6608 10550
rect 6268 10408 6340 10464
rect 6396 10408 6482 10464
rect 6538 10408 6608 10464
rect 6268 10322 6608 10408
rect 6268 10266 6340 10322
rect 6396 10266 6482 10322
rect 6538 10266 6608 10322
rect 6268 10180 6608 10266
rect 6268 10124 6340 10180
rect 6396 10124 6482 10180
rect 6538 10124 6608 10180
rect 6268 10038 6608 10124
rect 6268 9982 6340 10038
rect 6396 9982 6482 10038
rect 6538 9982 6608 10038
rect 6268 9896 6608 9982
rect 6268 9840 6340 9896
rect 6396 9840 6482 9896
rect 6538 9840 6608 9896
rect 6268 9754 6608 9840
rect 6268 9698 6340 9754
rect 6396 9698 6482 9754
rect 6538 9698 6608 9754
rect 6268 9612 6608 9698
rect 6268 9556 6340 9612
rect 6396 9556 6482 9612
rect 6538 9556 6608 9612
rect 6268 9470 6608 9556
rect 6268 9414 6340 9470
rect 6396 9414 6482 9470
rect 6538 9414 6608 9470
rect 6268 9328 6608 9414
rect 6268 9272 6340 9328
rect 6396 9272 6482 9328
rect 6538 9272 6608 9328
rect 6268 9186 6608 9272
rect 6268 9130 6340 9186
rect 6396 9130 6482 9186
rect 6538 9130 6608 9186
rect 6268 9044 6608 9130
rect 6268 8988 6340 9044
rect 6396 8988 6482 9044
rect 6538 8988 6608 9044
rect 6268 8902 6608 8988
rect 6268 8846 6340 8902
rect 6396 8846 6482 8902
rect 6538 8846 6608 8902
rect 6268 8760 6608 8846
rect 6268 8704 6340 8760
rect 6396 8704 6482 8760
rect 6538 8704 6608 8760
rect 6268 8618 6608 8704
rect 6268 8562 6340 8618
rect 6396 8562 6482 8618
rect 6538 8562 6608 8618
rect 6268 8476 6608 8562
rect 6268 8420 6340 8476
rect 6396 8420 6482 8476
rect 6538 8420 6608 8476
rect 6268 8334 6608 8420
rect 6268 8278 6340 8334
rect 6396 8278 6482 8334
rect 6538 8278 6608 8334
rect 6268 8192 6608 8278
rect 6268 8136 6340 8192
rect 6396 8136 6482 8192
rect 6538 8136 6608 8192
rect 6268 8050 6608 8136
rect 6268 7994 6340 8050
rect 6396 7994 6482 8050
rect 6538 7994 6608 8050
rect 6268 7908 6608 7994
rect 6268 7852 6340 7908
rect 6396 7852 6482 7908
rect 6538 7852 6608 7908
rect 6268 7766 6608 7852
rect 6268 7710 6340 7766
rect 6396 7710 6482 7766
rect 6538 7710 6608 7766
rect 6268 7624 6608 7710
rect 6268 7568 6340 7624
rect 6396 7568 6482 7624
rect 6538 7568 6608 7624
rect 6268 7482 6608 7568
rect 6268 7426 6340 7482
rect 6396 7426 6482 7482
rect 6538 7426 6608 7482
rect 6268 7340 6608 7426
rect 6268 7284 6340 7340
rect 6396 7284 6482 7340
rect 6538 7284 6608 7340
rect 6268 7198 6608 7284
rect 6268 7142 6340 7198
rect 6396 7142 6482 7198
rect 6538 7142 6608 7198
rect 6268 7056 6608 7142
rect 6268 7000 6340 7056
rect 6396 7000 6482 7056
rect 6538 7000 6608 7056
rect 6268 6914 6608 7000
rect 6268 6858 6340 6914
rect 6396 6858 6482 6914
rect 6538 6858 6608 6914
rect 6268 6772 6608 6858
rect 6268 6716 6340 6772
rect 6396 6716 6482 6772
rect 6538 6716 6608 6772
rect 6268 6630 6608 6716
rect 6268 6574 6340 6630
rect 6396 6574 6482 6630
rect 6538 6574 6608 6630
rect 6268 6488 6608 6574
rect 6268 6432 6340 6488
rect 6396 6432 6482 6488
rect 6538 6432 6608 6488
rect 6268 6346 6608 6432
rect 6268 6290 6340 6346
rect 6396 6290 6482 6346
rect 6538 6290 6608 6346
rect 6268 6204 6608 6290
rect 6268 6148 6340 6204
rect 6396 6148 6482 6204
rect 6538 6148 6608 6204
rect 6268 6062 6608 6148
rect 6268 6006 6340 6062
rect 6396 6006 6482 6062
rect 6538 6006 6608 6062
rect 6268 5920 6608 6006
rect 6268 5864 6340 5920
rect 6396 5864 6482 5920
rect 6538 5864 6608 5920
rect 6268 5778 6608 5864
rect 6268 5722 6340 5778
rect 6396 5722 6482 5778
rect 6538 5722 6608 5778
rect 6268 5636 6608 5722
rect 6268 5580 6340 5636
rect 6396 5580 6482 5636
rect 6538 5580 6608 5636
rect 6268 5494 6608 5580
rect 6268 5438 6340 5494
rect 6396 5438 6482 5494
rect 6538 5438 6608 5494
rect 6268 5352 6608 5438
rect 6268 5296 6340 5352
rect 6396 5296 6482 5352
rect 6538 5296 6608 5352
rect 6268 5210 6608 5296
rect 6268 5154 6340 5210
rect 6396 5154 6482 5210
rect 6538 5154 6608 5210
rect 6268 5068 6608 5154
rect 6268 5012 6340 5068
rect 6396 5012 6482 5068
rect 6538 5012 6608 5068
rect 6268 4926 6608 5012
rect 6268 4870 6340 4926
rect 6396 4870 6482 4926
rect 6538 4870 6608 4926
rect 6268 4784 6608 4870
rect 6268 4728 6340 4784
rect 6396 4728 6482 4784
rect 6538 4728 6608 4784
rect 6268 4642 6608 4728
rect 6268 4586 6340 4642
rect 6396 4586 6482 4642
rect 6538 4586 6608 4642
rect 6268 4500 6608 4586
rect 6268 4444 6340 4500
rect 6396 4444 6482 4500
rect 6538 4444 6608 4500
rect 6268 4358 6608 4444
rect 6268 4302 6340 4358
rect 6396 4302 6482 4358
rect 6538 4302 6608 4358
rect 6268 4216 6608 4302
rect 6268 4160 6340 4216
rect 6396 4160 6482 4216
rect 6538 4160 6608 4216
rect 6268 4074 6608 4160
rect 6268 4018 6340 4074
rect 6396 4018 6482 4074
rect 6538 4018 6608 4074
rect 6268 3932 6608 4018
rect 6268 3876 6340 3932
rect 6396 3876 6482 3932
rect 6538 3876 6608 3932
rect 6268 3790 6608 3876
rect 6268 3734 6340 3790
rect 6396 3734 6482 3790
rect 6538 3734 6608 3790
rect 6268 3648 6608 3734
rect 6268 3592 6340 3648
rect 6396 3592 6482 3648
rect 6538 3592 6608 3648
rect 6268 3506 6608 3592
rect 6268 3450 6340 3506
rect 6396 3450 6482 3506
rect 6538 3450 6608 3506
rect 6268 3364 6608 3450
rect 6268 3308 6340 3364
rect 6396 3308 6482 3364
rect 6538 3308 6608 3364
rect 6268 3222 6608 3308
rect 6268 3166 6340 3222
rect 6396 3166 6482 3222
rect 6538 3166 6608 3222
rect 6268 3080 6608 3166
rect 6268 3024 6340 3080
rect 6396 3024 6482 3080
rect 6538 3024 6608 3080
rect 6268 2938 6608 3024
rect 6268 2882 6340 2938
rect 6396 2882 6482 2938
rect 6538 2882 6608 2938
rect 6268 2796 6608 2882
rect 6268 2740 6340 2796
rect 6396 2740 6482 2796
rect 6538 2740 6608 2796
rect 6268 2654 6608 2740
rect 6268 2598 6340 2654
rect 6396 2598 6482 2654
rect 6538 2598 6608 2654
rect 6268 2512 6608 2598
rect 6268 2456 6340 2512
rect 6396 2456 6482 2512
rect 6538 2456 6608 2512
rect 6268 2370 6608 2456
rect 6268 2314 6340 2370
rect 6396 2314 6482 2370
rect 6538 2314 6608 2370
rect 6268 2228 6608 2314
rect 6268 2172 6340 2228
rect 6396 2172 6482 2228
rect 6538 2172 6608 2228
rect 6268 2086 6608 2172
rect 6268 2030 6340 2086
rect 6396 2030 6482 2086
rect 6538 2030 6608 2086
rect 6268 1944 6608 2030
rect 6268 1888 6340 1944
rect 6396 1888 6482 1944
rect 6538 1888 6608 1944
rect 6268 1802 6608 1888
rect 6268 1746 6340 1802
rect 6396 1746 6482 1802
rect 6538 1746 6608 1802
rect 6268 1660 6608 1746
rect 6268 1604 6340 1660
rect 6396 1604 6482 1660
rect 6538 1604 6608 1660
rect 6268 1518 6608 1604
rect 6268 1462 6340 1518
rect 6396 1462 6482 1518
rect 6538 1462 6608 1518
rect 6268 1376 6608 1462
rect 6268 1320 6340 1376
rect 6396 1320 6482 1376
rect 6538 1320 6608 1376
rect 6268 1234 6608 1320
rect 6268 1178 6340 1234
rect 6396 1178 6482 1234
rect 6538 1178 6608 1234
rect 6268 1092 6608 1178
rect 6268 1036 6340 1092
rect 6396 1036 6482 1092
rect 6538 1036 6608 1092
rect 6268 950 6608 1036
rect 6268 894 6340 950
rect 6396 894 6482 950
rect 6538 894 6608 950
rect 6268 808 6608 894
rect 6268 752 6340 808
rect 6396 752 6482 808
rect 6538 752 6608 808
rect 6268 666 6608 752
rect 6268 610 6340 666
rect 6396 610 6482 666
rect 6538 610 6608 666
rect 6268 524 6608 610
rect 6268 468 6340 524
rect 6396 468 6482 524
rect 6538 468 6608 524
rect 6268 400 6608 468
rect 6668 12310 7008 12400
rect 6668 12254 6742 12310
rect 6798 12254 6884 12310
rect 6940 12254 7008 12310
rect 6668 12168 7008 12254
rect 6668 12112 6742 12168
rect 6798 12112 6884 12168
rect 6940 12112 7008 12168
rect 6668 12026 7008 12112
rect 6668 11970 6742 12026
rect 6798 11970 6884 12026
rect 6940 11970 7008 12026
rect 6668 11884 7008 11970
rect 6668 11828 6742 11884
rect 6798 11828 6884 11884
rect 6940 11828 7008 11884
rect 6668 11742 7008 11828
rect 6668 11686 6742 11742
rect 6798 11686 6884 11742
rect 6940 11686 7008 11742
rect 6668 11600 7008 11686
rect 6668 11544 6742 11600
rect 6798 11544 6884 11600
rect 6940 11544 7008 11600
rect 6668 11458 7008 11544
rect 6668 11402 6742 11458
rect 6798 11402 6884 11458
rect 6940 11402 7008 11458
rect 6668 11316 7008 11402
rect 6668 11260 6742 11316
rect 6798 11260 6884 11316
rect 6940 11260 7008 11316
rect 6668 11174 7008 11260
rect 6668 11118 6742 11174
rect 6798 11118 6884 11174
rect 6940 11118 7008 11174
rect 6668 11032 7008 11118
rect 6668 10976 6742 11032
rect 6798 10976 6884 11032
rect 6940 10976 7008 11032
rect 6668 10890 7008 10976
rect 6668 10834 6742 10890
rect 6798 10834 6884 10890
rect 6940 10834 7008 10890
rect 6668 10748 7008 10834
rect 6668 10692 6742 10748
rect 6798 10692 6884 10748
rect 6940 10692 7008 10748
rect 6668 10606 7008 10692
rect 6668 10550 6742 10606
rect 6798 10550 6884 10606
rect 6940 10550 7008 10606
rect 6668 10464 7008 10550
rect 6668 10408 6742 10464
rect 6798 10408 6884 10464
rect 6940 10408 7008 10464
rect 6668 10322 7008 10408
rect 6668 10266 6742 10322
rect 6798 10266 6884 10322
rect 6940 10266 7008 10322
rect 6668 10180 7008 10266
rect 6668 10124 6742 10180
rect 6798 10124 6884 10180
rect 6940 10124 7008 10180
rect 6668 10038 7008 10124
rect 6668 9982 6742 10038
rect 6798 9982 6884 10038
rect 6940 9982 7008 10038
rect 6668 9896 7008 9982
rect 6668 9840 6742 9896
rect 6798 9840 6884 9896
rect 6940 9840 7008 9896
rect 6668 9754 7008 9840
rect 6668 9698 6742 9754
rect 6798 9698 6884 9754
rect 6940 9698 7008 9754
rect 6668 9612 7008 9698
rect 6668 9556 6742 9612
rect 6798 9556 6884 9612
rect 6940 9556 7008 9612
rect 6668 9470 7008 9556
rect 6668 9414 6742 9470
rect 6798 9414 6884 9470
rect 6940 9414 7008 9470
rect 6668 9328 7008 9414
rect 6668 9272 6742 9328
rect 6798 9272 6884 9328
rect 6940 9272 7008 9328
rect 6668 9186 7008 9272
rect 6668 9130 6742 9186
rect 6798 9130 6884 9186
rect 6940 9130 7008 9186
rect 6668 9044 7008 9130
rect 6668 8988 6742 9044
rect 6798 8988 6884 9044
rect 6940 8988 7008 9044
rect 6668 8902 7008 8988
rect 6668 8846 6742 8902
rect 6798 8846 6884 8902
rect 6940 8846 7008 8902
rect 6668 8760 7008 8846
rect 6668 8704 6742 8760
rect 6798 8704 6884 8760
rect 6940 8704 7008 8760
rect 6668 8618 7008 8704
rect 6668 8562 6742 8618
rect 6798 8562 6884 8618
rect 6940 8562 7008 8618
rect 6668 8476 7008 8562
rect 6668 8420 6742 8476
rect 6798 8420 6884 8476
rect 6940 8420 7008 8476
rect 6668 8334 7008 8420
rect 6668 8278 6742 8334
rect 6798 8278 6884 8334
rect 6940 8278 7008 8334
rect 6668 8192 7008 8278
rect 6668 8136 6742 8192
rect 6798 8136 6884 8192
rect 6940 8136 7008 8192
rect 6668 8050 7008 8136
rect 6668 7994 6742 8050
rect 6798 7994 6884 8050
rect 6940 7994 7008 8050
rect 6668 7908 7008 7994
rect 6668 7852 6742 7908
rect 6798 7852 6884 7908
rect 6940 7852 7008 7908
rect 6668 7766 7008 7852
rect 6668 7710 6742 7766
rect 6798 7710 6884 7766
rect 6940 7710 7008 7766
rect 6668 7624 7008 7710
rect 6668 7568 6742 7624
rect 6798 7568 6884 7624
rect 6940 7568 7008 7624
rect 6668 7482 7008 7568
rect 6668 7426 6742 7482
rect 6798 7426 6884 7482
rect 6940 7426 7008 7482
rect 6668 7340 7008 7426
rect 6668 7284 6742 7340
rect 6798 7284 6884 7340
rect 6940 7284 7008 7340
rect 6668 7198 7008 7284
rect 6668 7142 6742 7198
rect 6798 7142 6884 7198
rect 6940 7142 7008 7198
rect 6668 7056 7008 7142
rect 6668 7000 6742 7056
rect 6798 7000 6884 7056
rect 6940 7000 7008 7056
rect 6668 6914 7008 7000
rect 6668 6858 6742 6914
rect 6798 6858 6884 6914
rect 6940 6858 7008 6914
rect 6668 6772 7008 6858
rect 6668 6716 6742 6772
rect 6798 6716 6884 6772
rect 6940 6716 7008 6772
rect 6668 6630 7008 6716
rect 6668 6574 6742 6630
rect 6798 6574 6884 6630
rect 6940 6574 7008 6630
rect 6668 6488 7008 6574
rect 6668 6432 6742 6488
rect 6798 6432 6884 6488
rect 6940 6432 7008 6488
rect 6668 6346 7008 6432
rect 6668 6290 6742 6346
rect 6798 6290 6884 6346
rect 6940 6290 7008 6346
rect 6668 6204 7008 6290
rect 6668 6148 6742 6204
rect 6798 6148 6884 6204
rect 6940 6148 7008 6204
rect 6668 6062 7008 6148
rect 6668 6006 6742 6062
rect 6798 6006 6884 6062
rect 6940 6006 7008 6062
rect 6668 5920 7008 6006
rect 6668 5864 6742 5920
rect 6798 5864 6884 5920
rect 6940 5864 7008 5920
rect 6668 5778 7008 5864
rect 6668 5722 6742 5778
rect 6798 5722 6884 5778
rect 6940 5722 7008 5778
rect 6668 5636 7008 5722
rect 6668 5580 6742 5636
rect 6798 5580 6884 5636
rect 6940 5580 7008 5636
rect 6668 5494 7008 5580
rect 6668 5438 6742 5494
rect 6798 5438 6884 5494
rect 6940 5438 7008 5494
rect 6668 5352 7008 5438
rect 6668 5296 6742 5352
rect 6798 5296 6884 5352
rect 6940 5296 7008 5352
rect 6668 5210 7008 5296
rect 6668 5154 6742 5210
rect 6798 5154 6884 5210
rect 6940 5154 7008 5210
rect 6668 5068 7008 5154
rect 6668 5012 6742 5068
rect 6798 5012 6884 5068
rect 6940 5012 7008 5068
rect 6668 4926 7008 5012
rect 6668 4870 6742 4926
rect 6798 4870 6884 4926
rect 6940 4870 7008 4926
rect 6668 4784 7008 4870
rect 6668 4728 6742 4784
rect 6798 4728 6884 4784
rect 6940 4728 7008 4784
rect 6668 4642 7008 4728
rect 6668 4586 6742 4642
rect 6798 4586 6884 4642
rect 6940 4586 7008 4642
rect 6668 4500 7008 4586
rect 6668 4444 6742 4500
rect 6798 4444 6884 4500
rect 6940 4444 7008 4500
rect 6668 4358 7008 4444
rect 6668 4302 6742 4358
rect 6798 4302 6884 4358
rect 6940 4302 7008 4358
rect 6668 4216 7008 4302
rect 6668 4160 6742 4216
rect 6798 4160 6884 4216
rect 6940 4160 7008 4216
rect 6668 4074 7008 4160
rect 6668 4018 6742 4074
rect 6798 4018 6884 4074
rect 6940 4018 7008 4074
rect 6668 3932 7008 4018
rect 6668 3876 6742 3932
rect 6798 3876 6884 3932
rect 6940 3876 7008 3932
rect 6668 3790 7008 3876
rect 6668 3734 6742 3790
rect 6798 3734 6884 3790
rect 6940 3734 7008 3790
rect 6668 3648 7008 3734
rect 6668 3592 6742 3648
rect 6798 3592 6884 3648
rect 6940 3592 7008 3648
rect 6668 3506 7008 3592
rect 6668 3450 6742 3506
rect 6798 3450 6884 3506
rect 6940 3450 7008 3506
rect 6668 3364 7008 3450
rect 6668 3308 6742 3364
rect 6798 3308 6884 3364
rect 6940 3308 7008 3364
rect 6668 3222 7008 3308
rect 6668 3166 6742 3222
rect 6798 3166 6884 3222
rect 6940 3166 7008 3222
rect 6668 3080 7008 3166
rect 6668 3024 6742 3080
rect 6798 3024 6884 3080
rect 6940 3024 7008 3080
rect 6668 2938 7008 3024
rect 6668 2882 6742 2938
rect 6798 2882 6884 2938
rect 6940 2882 7008 2938
rect 6668 2796 7008 2882
rect 6668 2740 6742 2796
rect 6798 2740 6884 2796
rect 6940 2740 7008 2796
rect 6668 2654 7008 2740
rect 6668 2598 6742 2654
rect 6798 2598 6884 2654
rect 6940 2598 7008 2654
rect 6668 2512 7008 2598
rect 6668 2456 6742 2512
rect 6798 2456 6884 2512
rect 6940 2456 7008 2512
rect 6668 2370 7008 2456
rect 6668 2314 6742 2370
rect 6798 2314 6884 2370
rect 6940 2314 7008 2370
rect 6668 2228 7008 2314
rect 6668 2172 6742 2228
rect 6798 2172 6884 2228
rect 6940 2172 7008 2228
rect 6668 2086 7008 2172
rect 6668 2030 6742 2086
rect 6798 2030 6884 2086
rect 6940 2030 7008 2086
rect 6668 1944 7008 2030
rect 6668 1888 6742 1944
rect 6798 1888 6884 1944
rect 6940 1888 7008 1944
rect 6668 1802 7008 1888
rect 6668 1746 6742 1802
rect 6798 1746 6884 1802
rect 6940 1746 7008 1802
rect 6668 1660 7008 1746
rect 6668 1604 6742 1660
rect 6798 1604 6884 1660
rect 6940 1604 7008 1660
rect 6668 1518 7008 1604
rect 6668 1462 6742 1518
rect 6798 1462 6884 1518
rect 6940 1462 7008 1518
rect 6668 1376 7008 1462
rect 6668 1320 6742 1376
rect 6798 1320 6884 1376
rect 6940 1320 7008 1376
rect 6668 1234 7008 1320
rect 6668 1178 6742 1234
rect 6798 1178 6884 1234
rect 6940 1178 7008 1234
rect 6668 1092 7008 1178
rect 6668 1036 6742 1092
rect 6798 1036 6884 1092
rect 6940 1036 7008 1092
rect 6668 950 7008 1036
rect 6668 894 6742 950
rect 6798 894 6884 950
rect 6940 894 7008 950
rect 6668 808 7008 894
rect 6668 752 6742 808
rect 6798 752 6884 808
rect 6940 752 7008 808
rect 6668 666 7008 752
rect 6668 610 6742 666
rect 6798 610 6884 666
rect 6940 610 7008 666
rect 6668 524 7008 610
rect 6668 468 6742 524
rect 6798 468 6884 524
rect 6940 468 7008 524
rect 6668 400 7008 468
rect 7068 12310 7408 12400
rect 7068 12254 7145 12310
rect 7201 12254 7287 12310
rect 7343 12254 7408 12310
rect 7068 12168 7408 12254
rect 7068 12112 7145 12168
rect 7201 12112 7287 12168
rect 7343 12112 7408 12168
rect 7068 12026 7408 12112
rect 7068 11970 7145 12026
rect 7201 11970 7287 12026
rect 7343 11970 7408 12026
rect 7068 11884 7408 11970
rect 7068 11828 7145 11884
rect 7201 11828 7287 11884
rect 7343 11828 7408 11884
rect 7068 11742 7408 11828
rect 7068 11686 7145 11742
rect 7201 11686 7287 11742
rect 7343 11686 7408 11742
rect 7068 11600 7408 11686
rect 7068 11544 7145 11600
rect 7201 11544 7287 11600
rect 7343 11544 7408 11600
rect 7068 11458 7408 11544
rect 7068 11402 7145 11458
rect 7201 11402 7287 11458
rect 7343 11402 7408 11458
rect 7068 11316 7408 11402
rect 7068 11260 7145 11316
rect 7201 11260 7287 11316
rect 7343 11260 7408 11316
rect 7068 11174 7408 11260
rect 7068 11118 7145 11174
rect 7201 11118 7287 11174
rect 7343 11118 7408 11174
rect 7068 11032 7408 11118
rect 7068 10976 7145 11032
rect 7201 10976 7287 11032
rect 7343 10976 7408 11032
rect 7068 10890 7408 10976
rect 7068 10834 7145 10890
rect 7201 10834 7287 10890
rect 7343 10834 7408 10890
rect 7068 10748 7408 10834
rect 7068 10692 7145 10748
rect 7201 10692 7287 10748
rect 7343 10692 7408 10748
rect 7068 10606 7408 10692
rect 7068 10550 7145 10606
rect 7201 10550 7287 10606
rect 7343 10550 7408 10606
rect 7068 10464 7408 10550
rect 7068 10408 7145 10464
rect 7201 10408 7287 10464
rect 7343 10408 7408 10464
rect 7068 10322 7408 10408
rect 7068 10266 7145 10322
rect 7201 10266 7287 10322
rect 7343 10266 7408 10322
rect 7068 10180 7408 10266
rect 7068 10124 7145 10180
rect 7201 10124 7287 10180
rect 7343 10124 7408 10180
rect 7068 10038 7408 10124
rect 7068 9982 7145 10038
rect 7201 9982 7287 10038
rect 7343 9982 7408 10038
rect 7068 9896 7408 9982
rect 7068 9840 7145 9896
rect 7201 9840 7287 9896
rect 7343 9840 7408 9896
rect 7068 9754 7408 9840
rect 7068 9698 7145 9754
rect 7201 9698 7287 9754
rect 7343 9698 7408 9754
rect 7068 9612 7408 9698
rect 7068 9556 7145 9612
rect 7201 9556 7287 9612
rect 7343 9556 7408 9612
rect 7068 9470 7408 9556
rect 7068 9414 7145 9470
rect 7201 9414 7287 9470
rect 7343 9414 7408 9470
rect 7068 9328 7408 9414
rect 7068 9272 7145 9328
rect 7201 9272 7287 9328
rect 7343 9272 7408 9328
rect 7068 9186 7408 9272
rect 7068 9130 7145 9186
rect 7201 9130 7287 9186
rect 7343 9130 7408 9186
rect 7068 9044 7408 9130
rect 7068 8988 7145 9044
rect 7201 8988 7287 9044
rect 7343 8988 7408 9044
rect 7068 8902 7408 8988
rect 7068 8846 7145 8902
rect 7201 8846 7287 8902
rect 7343 8846 7408 8902
rect 7068 8760 7408 8846
rect 7068 8704 7145 8760
rect 7201 8704 7287 8760
rect 7343 8704 7408 8760
rect 7068 8618 7408 8704
rect 7068 8562 7145 8618
rect 7201 8562 7287 8618
rect 7343 8562 7408 8618
rect 7068 8476 7408 8562
rect 7068 8420 7145 8476
rect 7201 8420 7287 8476
rect 7343 8420 7408 8476
rect 7068 8334 7408 8420
rect 7068 8278 7145 8334
rect 7201 8278 7287 8334
rect 7343 8278 7408 8334
rect 7068 8192 7408 8278
rect 7068 8136 7145 8192
rect 7201 8136 7287 8192
rect 7343 8136 7408 8192
rect 7068 8050 7408 8136
rect 7068 7994 7145 8050
rect 7201 7994 7287 8050
rect 7343 7994 7408 8050
rect 7068 7908 7408 7994
rect 7068 7852 7145 7908
rect 7201 7852 7287 7908
rect 7343 7852 7408 7908
rect 7068 7766 7408 7852
rect 7068 7710 7145 7766
rect 7201 7710 7287 7766
rect 7343 7710 7408 7766
rect 7068 7624 7408 7710
rect 7068 7568 7145 7624
rect 7201 7568 7287 7624
rect 7343 7568 7408 7624
rect 7068 7482 7408 7568
rect 7068 7426 7145 7482
rect 7201 7426 7287 7482
rect 7343 7426 7408 7482
rect 7068 7340 7408 7426
rect 7068 7284 7145 7340
rect 7201 7284 7287 7340
rect 7343 7284 7408 7340
rect 7068 7198 7408 7284
rect 7068 7142 7145 7198
rect 7201 7142 7287 7198
rect 7343 7142 7408 7198
rect 7068 7056 7408 7142
rect 7068 7000 7145 7056
rect 7201 7000 7287 7056
rect 7343 7000 7408 7056
rect 7068 6914 7408 7000
rect 7068 6858 7145 6914
rect 7201 6858 7287 6914
rect 7343 6858 7408 6914
rect 7068 6772 7408 6858
rect 7068 6716 7145 6772
rect 7201 6716 7287 6772
rect 7343 6716 7408 6772
rect 7068 6630 7408 6716
rect 7068 6574 7145 6630
rect 7201 6574 7287 6630
rect 7343 6574 7408 6630
rect 7068 6488 7408 6574
rect 7068 6432 7145 6488
rect 7201 6432 7287 6488
rect 7343 6432 7408 6488
rect 7068 6346 7408 6432
rect 7068 6290 7145 6346
rect 7201 6290 7287 6346
rect 7343 6290 7408 6346
rect 7068 6204 7408 6290
rect 7068 6148 7145 6204
rect 7201 6148 7287 6204
rect 7343 6148 7408 6204
rect 7068 6062 7408 6148
rect 7068 6006 7145 6062
rect 7201 6006 7287 6062
rect 7343 6006 7408 6062
rect 7068 5920 7408 6006
rect 7068 5864 7145 5920
rect 7201 5864 7287 5920
rect 7343 5864 7408 5920
rect 7068 5778 7408 5864
rect 7068 5722 7145 5778
rect 7201 5722 7287 5778
rect 7343 5722 7408 5778
rect 7068 5636 7408 5722
rect 7068 5580 7145 5636
rect 7201 5580 7287 5636
rect 7343 5580 7408 5636
rect 7068 5494 7408 5580
rect 7068 5438 7145 5494
rect 7201 5438 7287 5494
rect 7343 5438 7408 5494
rect 7068 5352 7408 5438
rect 7068 5296 7145 5352
rect 7201 5296 7287 5352
rect 7343 5296 7408 5352
rect 7068 5210 7408 5296
rect 7068 5154 7145 5210
rect 7201 5154 7287 5210
rect 7343 5154 7408 5210
rect 7068 5068 7408 5154
rect 7068 5012 7145 5068
rect 7201 5012 7287 5068
rect 7343 5012 7408 5068
rect 7068 4926 7408 5012
rect 7068 4870 7145 4926
rect 7201 4870 7287 4926
rect 7343 4870 7408 4926
rect 7068 4784 7408 4870
rect 7068 4728 7145 4784
rect 7201 4728 7287 4784
rect 7343 4728 7408 4784
rect 7068 4642 7408 4728
rect 7068 4586 7145 4642
rect 7201 4586 7287 4642
rect 7343 4586 7408 4642
rect 7068 4500 7408 4586
rect 7068 4444 7145 4500
rect 7201 4444 7287 4500
rect 7343 4444 7408 4500
rect 7068 4358 7408 4444
rect 7068 4302 7145 4358
rect 7201 4302 7287 4358
rect 7343 4302 7408 4358
rect 7068 4216 7408 4302
rect 7068 4160 7145 4216
rect 7201 4160 7287 4216
rect 7343 4160 7408 4216
rect 7068 4074 7408 4160
rect 7068 4018 7145 4074
rect 7201 4018 7287 4074
rect 7343 4018 7408 4074
rect 7068 3932 7408 4018
rect 7068 3876 7145 3932
rect 7201 3876 7287 3932
rect 7343 3876 7408 3932
rect 7068 3790 7408 3876
rect 7068 3734 7145 3790
rect 7201 3734 7287 3790
rect 7343 3734 7408 3790
rect 7068 3648 7408 3734
rect 7068 3592 7145 3648
rect 7201 3592 7287 3648
rect 7343 3592 7408 3648
rect 7068 3506 7408 3592
rect 7068 3450 7145 3506
rect 7201 3450 7287 3506
rect 7343 3450 7408 3506
rect 7068 3364 7408 3450
rect 7068 3308 7145 3364
rect 7201 3308 7287 3364
rect 7343 3308 7408 3364
rect 7068 3222 7408 3308
rect 7068 3166 7145 3222
rect 7201 3166 7287 3222
rect 7343 3166 7408 3222
rect 7068 3080 7408 3166
rect 7068 3024 7145 3080
rect 7201 3024 7287 3080
rect 7343 3024 7408 3080
rect 7068 2938 7408 3024
rect 7068 2882 7145 2938
rect 7201 2882 7287 2938
rect 7343 2882 7408 2938
rect 7068 2796 7408 2882
rect 7068 2740 7145 2796
rect 7201 2740 7287 2796
rect 7343 2740 7408 2796
rect 7068 2654 7408 2740
rect 7068 2598 7145 2654
rect 7201 2598 7287 2654
rect 7343 2598 7408 2654
rect 7068 2512 7408 2598
rect 7068 2456 7145 2512
rect 7201 2456 7287 2512
rect 7343 2456 7408 2512
rect 7068 2370 7408 2456
rect 7068 2314 7145 2370
rect 7201 2314 7287 2370
rect 7343 2314 7408 2370
rect 7068 2228 7408 2314
rect 7068 2172 7145 2228
rect 7201 2172 7287 2228
rect 7343 2172 7408 2228
rect 7068 2086 7408 2172
rect 7068 2030 7145 2086
rect 7201 2030 7287 2086
rect 7343 2030 7408 2086
rect 7068 1944 7408 2030
rect 7068 1888 7145 1944
rect 7201 1888 7287 1944
rect 7343 1888 7408 1944
rect 7068 1802 7408 1888
rect 7068 1746 7145 1802
rect 7201 1746 7287 1802
rect 7343 1746 7408 1802
rect 7068 1660 7408 1746
rect 7068 1604 7145 1660
rect 7201 1604 7287 1660
rect 7343 1604 7408 1660
rect 7068 1518 7408 1604
rect 7068 1462 7145 1518
rect 7201 1462 7287 1518
rect 7343 1462 7408 1518
rect 7068 1376 7408 1462
rect 7068 1320 7145 1376
rect 7201 1320 7287 1376
rect 7343 1320 7408 1376
rect 7068 1234 7408 1320
rect 7068 1178 7145 1234
rect 7201 1178 7287 1234
rect 7343 1178 7408 1234
rect 7068 1092 7408 1178
rect 7068 1036 7145 1092
rect 7201 1036 7287 1092
rect 7343 1036 7408 1092
rect 7068 950 7408 1036
rect 7068 894 7145 950
rect 7201 894 7287 950
rect 7343 894 7408 950
rect 7068 808 7408 894
rect 7068 752 7145 808
rect 7201 752 7287 808
rect 7343 752 7408 808
rect 7068 666 7408 752
rect 7068 610 7145 666
rect 7201 610 7287 666
rect 7343 610 7408 666
rect 7068 524 7408 610
rect 7068 468 7145 524
rect 7201 468 7287 524
rect 7343 468 7408 524
rect 7068 400 7408 468
rect 7468 12310 7808 12400
rect 7468 12254 7539 12310
rect 7595 12254 7681 12310
rect 7737 12254 7808 12310
rect 7468 12168 7808 12254
rect 7468 12112 7539 12168
rect 7595 12112 7681 12168
rect 7737 12112 7808 12168
rect 7468 12026 7808 12112
rect 7468 11970 7539 12026
rect 7595 11970 7681 12026
rect 7737 11970 7808 12026
rect 7468 11884 7808 11970
rect 7468 11828 7539 11884
rect 7595 11828 7681 11884
rect 7737 11828 7808 11884
rect 7468 11742 7808 11828
rect 7468 11686 7539 11742
rect 7595 11686 7681 11742
rect 7737 11686 7808 11742
rect 7468 11600 7808 11686
rect 7468 11544 7539 11600
rect 7595 11544 7681 11600
rect 7737 11544 7808 11600
rect 7468 11458 7808 11544
rect 7468 11402 7539 11458
rect 7595 11402 7681 11458
rect 7737 11402 7808 11458
rect 7468 11316 7808 11402
rect 7468 11260 7539 11316
rect 7595 11260 7681 11316
rect 7737 11260 7808 11316
rect 7468 11174 7808 11260
rect 7468 11118 7539 11174
rect 7595 11118 7681 11174
rect 7737 11118 7808 11174
rect 7468 11032 7808 11118
rect 7468 10976 7539 11032
rect 7595 10976 7681 11032
rect 7737 10976 7808 11032
rect 7468 10890 7808 10976
rect 7468 10834 7539 10890
rect 7595 10834 7681 10890
rect 7737 10834 7808 10890
rect 7468 10748 7808 10834
rect 7468 10692 7539 10748
rect 7595 10692 7681 10748
rect 7737 10692 7808 10748
rect 7468 10606 7808 10692
rect 7468 10550 7539 10606
rect 7595 10550 7681 10606
rect 7737 10550 7808 10606
rect 7468 10464 7808 10550
rect 7468 10408 7539 10464
rect 7595 10408 7681 10464
rect 7737 10408 7808 10464
rect 7468 10322 7808 10408
rect 7468 10266 7539 10322
rect 7595 10266 7681 10322
rect 7737 10266 7808 10322
rect 7468 10180 7808 10266
rect 7468 10124 7539 10180
rect 7595 10124 7681 10180
rect 7737 10124 7808 10180
rect 7468 10038 7808 10124
rect 7468 9982 7539 10038
rect 7595 9982 7681 10038
rect 7737 9982 7808 10038
rect 7468 9896 7808 9982
rect 7468 9840 7539 9896
rect 7595 9840 7681 9896
rect 7737 9840 7808 9896
rect 7468 9754 7808 9840
rect 7468 9698 7539 9754
rect 7595 9698 7681 9754
rect 7737 9698 7808 9754
rect 7468 9612 7808 9698
rect 7468 9556 7539 9612
rect 7595 9556 7681 9612
rect 7737 9556 7808 9612
rect 7468 9470 7808 9556
rect 7468 9414 7539 9470
rect 7595 9414 7681 9470
rect 7737 9414 7808 9470
rect 7468 9328 7808 9414
rect 7468 9272 7539 9328
rect 7595 9272 7681 9328
rect 7737 9272 7808 9328
rect 7468 9186 7808 9272
rect 7468 9130 7539 9186
rect 7595 9130 7681 9186
rect 7737 9130 7808 9186
rect 7468 9044 7808 9130
rect 7468 8988 7539 9044
rect 7595 8988 7681 9044
rect 7737 8988 7808 9044
rect 7468 8902 7808 8988
rect 7468 8846 7539 8902
rect 7595 8846 7681 8902
rect 7737 8846 7808 8902
rect 7468 8760 7808 8846
rect 7468 8704 7539 8760
rect 7595 8704 7681 8760
rect 7737 8704 7808 8760
rect 7468 8618 7808 8704
rect 7468 8562 7539 8618
rect 7595 8562 7681 8618
rect 7737 8562 7808 8618
rect 7468 8476 7808 8562
rect 7468 8420 7539 8476
rect 7595 8420 7681 8476
rect 7737 8420 7808 8476
rect 7468 8334 7808 8420
rect 7468 8278 7539 8334
rect 7595 8278 7681 8334
rect 7737 8278 7808 8334
rect 7468 8192 7808 8278
rect 7468 8136 7539 8192
rect 7595 8136 7681 8192
rect 7737 8136 7808 8192
rect 7468 8050 7808 8136
rect 7468 7994 7539 8050
rect 7595 7994 7681 8050
rect 7737 7994 7808 8050
rect 7468 7908 7808 7994
rect 7468 7852 7539 7908
rect 7595 7852 7681 7908
rect 7737 7852 7808 7908
rect 7468 7766 7808 7852
rect 7468 7710 7539 7766
rect 7595 7710 7681 7766
rect 7737 7710 7808 7766
rect 7468 7624 7808 7710
rect 7468 7568 7539 7624
rect 7595 7568 7681 7624
rect 7737 7568 7808 7624
rect 7468 7482 7808 7568
rect 7468 7426 7539 7482
rect 7595 7426 7681 7482
rect 7737 7426 7808 7482
rect 7468 7340 7808 7426
rect 7468 7284 7539 7340
rect 7595 7284 7681 7340
rect 7737 7284 7808 7340
rect 7468 7198 7808 7284
rect 7468 7142 7539 7198
rect 7595 7142 7681 7198
rect 7737 7142 7808 7198
rect 7468 7056 7808 7142
rect 7468 7000 7539 7056
rect 7595 7000 7681 7056
rect 7737 7000 7808 7056
rect 7468 6914 7808 7000
rect 7468 6858 7539 6914
rect 7595 6858 7681 6914
rect 7737 6858 7808 6914
rect 7468 6772 7808 6858
rect 7468 6716 7539 6772
rect 7595 6716 7681 6772
rect 7737 6716 7808 6772
rect 7468 6630 7808 6716
rect 7468 6574 7539 6630
rect 7595 6574 7681 6630
rect 7737 6574 7808 6630
rect 7468 6488 7808 6574
rect 7468 6432 7539 6488
rect 7595 6432 7681 6488
rect 7737 6432 7808 6488
rect 7468 6346 7808 6432
rect 7468 6290 7539 6346
rect 7595 6290 7681 6346
rect 7737 6290 7808 6346
rect 7468 6204 7808 6290
rect 7468 6148 7539 6204
rect 7595 6148 7681 6204
rect 7737 6148 7808 6204
rect 7468 6062 7808 6148
rect 7468 6006 7539 6062
rect 7595 6006 7681 6062
rect 7737 6006 7808 6062
rect 7468 5920 7808 6006
rect 7468 5864 7539 5920
rect 7595 5864 7681 5920
rect 7737 5864 7808 5920
rect 7468 5778 7808 5864
rect 7468 5722 7539 5778
rect 7595 5722 7681 5778
rect 7737 5722 7808 5778
rect 7468 5636 7808 5722
rect 7468 5580 7539 5636
rect 7595 5580 7681 5636
rect 7737 5580 7808 5636
rect 7468 5494 7808 5580
rect 7468 5438 7539 5494
rect 7595 5438 7681 5494
rect 7737 5438 7808 5494
rect 7468 5352 7808 5438
rect 7468 5296 7539 5352
rect 7595 5296 7681 5352
rect 7737 5296 7808 5352
rect 7468 5210 7808 5296
rect 7468 5154 7539 5210
rect 7595 5154 7681 5210
rect 7737 5154 7808 5210
rect 7468 5068 7808 5154
rect 7468 5012 7539 5068
rect 7595 5012 7681 5068
rect 7737 5012 7808 5068
rect 7468 4926 7808 5012
rect 7468 4870 7539 4926
rect 7595 4870 7681 4926
rect 7737 4870 7808 4926
rect 7468 4784 7808 4870
rect 7468 4728 7539 4784
rect 7595 4728 7681 4784
rect 7737 4728 7808 4784
rect 7468 4642 7808 4728
rect 7468 4586 7539 4642
rect 7595 4586 7681 4642
rect 7737 4586 7808 4642
rect 7468 4500 7808 4586
rect 7468 4444 7539 4500
rect 7595 4444 7681 4500
rect 7737 4444 7808 4500
rect 7468 4358 7808 4444
rect 7468 4302 7539 4358
rect 7595 4302 7681 4358
rect 7737 4302 7808 4358
rect 7468 4216 7808 4302
rect 7468 4160 7539 4216
rect 7595 4160 7681 4216
rect 7737 4160 7808 4216
rect 7468 4074 7808 4160
rect 7468 4018 7539 4074
rect 7595 4018 7681 4074
rect 7737 4018 7808 4074
rect 7468 3932 7808 4018
rect 7468 3876 7539 3932
rect 7595 3876 7681 3932
rect 7737 3876 7808 3932
rect 7468 3790 7808 3876
rect 7468 3734 7539 3790
rect 7595 3734 7681 3790
rect 7737 3734 7808 3790
rect 7468 3648 7808 3734
rect 7468 3592 7539 3648
rect 7595 3592 7681 3648
rect 7737 3592 7808 3648
rect 7468 3506 7808 3592
rect 7468 3450 7539 3506
rect 7595 3450 7681 3506
rect 7737 3450 7808 3506
rect 7468 3364 7808 3450
rect 7468 3308 7539 3364
rect 7595 3308 7681 3364
rect 7737 3308 7808 3364
rect 7468 3222 7808 3308
rect 7468 3166 7539 3222
rect 7595 3166 7681 3222
rect 7737 3166 7808 3222
rect 7468 3080 7808 3166
rect 7468 3024 7539 3080
rect 7595 3024 7681 3080
rect 7737 3024 7808 3080
rect 7468 2938 7808 3024
rect 7468 2882 7539 2938
rect 7595 2882 7681 2938
rect 7737 2882 7808 2938
rect 7468 2796 7808 2882
rect 7468 2740 7539 2796
rect 7595 2740 7681 2796
rect 7737 2740 7808 2796
rect 7468 2654 7808 2740
rect 7468 2598 7539 2654
rect 7595 2598 7681 2654
rect 7737 2598 7808 2654
rect 7468 2512 7808 2598
rect 7468 2456 7539 2512
rect 7595 2456 7681 2512
rect 7737 2456 7808 2512
rect 7468 2370 7808 2456
rect 7468 2314 7539 2370
rect 7595 2314 7681 2370
rect 7737 2314 7808 2370
rect 7468 2228 7808 2314
rect 7468 2172 7539 2228
rect 7595 2172 7681 2228
rect 7737 2172 7808 2228
rect 7468 2086 7808 2172
rect 7468 2030 7539 2086
rect 7595 2030 7681 2086
rect 7737 2030 7808 2086
rect 7468 1944 7808 2030
rect 7468 1888 7539 1944
rect 7595 1888 7681 1944
rect 7737 1888 7808 1944
rect 7468 1802 7808 1888
rect 7468 1746 7539 1802
rect 7595 1746 7681 1802
rect 7737 1746 7808 1802
rect 7468 1660 7808 1746
rect 7468 1604 7539 1660
rect 7595 1604 7681 1660
rect 7737 1604 7808 1660
rect 7468 1518 7808 1604
rect 7468 1462 7539 1518
rect 7595 1462 7681 1518
rect 7737 1462 7808 1518
rect 7468 1376 7808 1462
rect 7468 1320 7539 1376
rect 7595 1320 7681 1376
rect 7737 1320 7808 1376
rect 7468 1234 7808 1320
rect 7468 1178 7539 1234
rect 7595 1178 7681 1234
rect 7737 1178 7808 1234
rect 7468 1092 7808 1178
rect 7468 1036 7539 1092
rect 7595 1036 7681 1092
rect 7737 1036 7808 1092
rect 7468 950 7808 1036
rect 7468 894 7539 950
rect 7595 894 7681 950
rect 7737 894 7808 950
rect 7468 808 7808 894
rect 7468 752 7539 808
rect 7595 752 7681 808
rect 7737 752 7808 808
rect 7468 666 7808 752
rect 7468 610 7539 666
rect 7595 610 7681 666
rect 7737 610 7808 666
rect 7468 524 7808 610
rect 7468 468 7539 524
rect 7595 468 7681 524
rect 7737 468 7808 524
rect 7468 400 7808 468
rect 7868 12310 8208 12400
rect 7868 12254 7940 12310
rect 7996 12254 8082 12310
rect 8138 12254 8208 12310
rect 7868 12168 8208 12254
rect 7868 12112 7940 12168
rect 7996 12112 8082 12168
rect 8138 12112 8208 12168
rect 7868 12026 8208 12112
rect 7868 11970 7940 12026
rect 7996 11970 8082 12026
rect 8138 11970 8208 12026
rect 7868 11884 8208 11970
rect 7868 11828 7940 11884
rect 7996 11828 8082 11884
rect 8138 11828 8208 11884
rect 7868 11742 8208 11828
rect 7868 11686 7940 11742
rect 7996 11686 8082 11742
rect 8138 11686 8208 11742
rect 7868 11600 8208 11686
rect 7868 11544 7940 11600
rect 7996 11544 8082 11600
rect 8138 11544 8208 11600
rect 7868 11458 8208 11544
rect 7868 11402 7940 11458
rect 7996 11402 8082 11458
rect 8138 11402 8208 11458
rect 7868 11316 8208 11402
rect 7868 11260 7940 11316
rect 7996 11260 8082 11316
rect 8138 11260 8208 11316
rect 7868 11174 8208 11260
rect 7868 11118 7940 11174
rect 7996 11118 8082 11174
rect 8138 11118 8208 11174
rect 7868 11032 8208 11118
rect 7868 10976 7940 11032
rect 7996 10976 8082 11032
rect 8138 10976 8208 11032
rect 7868 10890 8208 10976
rect 7868 10834 7940 10890
rect 7996 10834 8082 10890
rect 8138 10834 8208 10890
rect 7868 10748 8208 10834
rect 7868 10692 7940 10748
rect 7996 10692 8082 10748
rect 8138 10692 8208 10748
rect 7868 10606 8208 10692
rect 7868 10550 7940 10606
rect 7996 10550 8082 10606
rect 8138 10550 8208 10606
rect 7868 10464 8208 10550
rect 7868 10408 7940 10464
rect 7996 10408 8082 10464
rect 8138 10408 8208 10464
rect 7868 10322 8208 10408
rect 7868 10266 7940 10322
rect 7996 10266 8082 10322
rect 8138 10266 8208 10322
rect 7868 10180 8208 10266
rect 7868 10124 7940 10180
rect 7996 10124 8082 10180
rect 8138 10124 8208 10180
rect 7868 10038 8208 10124
rect 7868 9982 7940 10038
rect 7996 9982 8082 10038
rect 8138 9982 8208 10038
rect 7868 9896 8208 9982
rect 7868 9840 7940 9896
rect 7996 9840 8082 9896
rect 8138 9840 8208 9896
rect 7868 9754 8208 9840
rect 7868 9698 7940 9754
rect 7996 9698 8082 9754
rect 8138 9698 8208 9754
rect 7868 9612 8208 9698
rect 7868 9556 7940 9612
rect 7996 9556 8082 9612
rect 8138 9556 8208 9612
rect 7868 9470 8208 9556
rect 7868 9414 7940 9470
rect 7996 9414 8082 9470
rect 8138 9414 8208 9470
rect 7868 9328 8208 9414
rect 7868 9272 7940 9328
rect 7996 9272 8082 9328
rect 8138 9272 8208 9328
rect 7868 9186 8208 9272
rect 7868 9130 7940 9186
rect 7996 9130 8082 9186
rect 8138 9130 8208 9186
rect 7868 9044 8208 9130
rect 7868 8988 7940 9044
rect 7996 8988 8082 9044
rect 8138 8988 8208 9044
rect 7868 8902 8208 8988
rect 7868 8846 7940 8902
rect 7996 8846 8082 8902
rect 8138 8846 8208 8902
rect 7868 8760 8208 8846
rect 7868 8704 7940 8760
rect 7996 8704 8082 8760
rect 8138 8704 8208 8760
rect 7868 8618 8208 8704
rect 7868 8562 7940 8618
rect 7996 8562 8082 8618
rect 8138 8562 8208 8618
rect 7868 8476 8208 8562
rect 7868 8420 7940 8476
rect 7996 8420 8082 8476
rect 8138 8420 8208 8476
rect 7868 8334 8208 8420
rect 7868 8278 7940 8334
rect 7996 8278 8082 8334
rect 8138 8278 8208 8334
rect 7868 8192 8208 8278
rect 7868 8136 7940 8192
rect 7996 8136 8082 8192
rect 8138 8136 8208 8192
rect 7868 8050 8208 8136
rect 7868 7994 7940 8050
rect 7996 7994 8082 8050
rect 8138 7994 8208 8050
rect 7868 7908 8208 7994
rect 7868 7852 7940 7908
rect 7996 7852 8082 7908
rect 8138 7852 8208 7908
rect 7868 7766 8208 7852
rect 7868 7710 7940 7766
rect 7996 7710 8082 7766
rect 8138 7710 8208 7766
rect 7868 7624 8208 7710
rect 7868 7568 7940 7624
rect 7996 7568 8082 7624
rect 8138 7568 8208 7624
rect 7868 7482 8208 7568
rect 7868 7426 7940 7482
rect 7996 7426 8082 7482
rect 8138 7426 8208 7482
rect 7868 7340 8208 7426
rect 7868 7284 7940 7340
rect 7996 7284 8082 7340
rect 8138 7284 8208 7340
rect 7868 7198 8208 7284
rect 7868 7142 7940 7198
rect 7996 7142 8082 7198
rect 8138 7142 8208 7198
rect 7868 7056 8208 7142
rect 7868 7000 7940 7056
rect 7996 7000 8082 7056
rect 8138 7000 8208 7056
rect 7868 6914 8208 7000
rect 7868 6858 7940 6914
rect 7996 6858 8082 6914
rect 8138 6858 8208 6914
rect 7868 6772 8208 6858
rect 7868 6716 7940 6772
rect 7996 6716 8082 6772
rect 8138 6716 8208 6772
rect 7868 6630 8208 6716
rect 7868 6574 7940 6630
rect 7996 6574 8082 6630
rect 8138 6574 8208 6630
rect 7868 6488 8208 6574
rect 7868 6432 7940 6488
rect 7996 6432 8082 6488
rect 8138 6432 8208 6488
rect 7868 6346 8208 6432
rect 7868 6290 7940 6346
rect 7996 6290 8082 6346
rect 8138 6290 8208 6346
rect 7868 6204 8208 6290
rect 7868 6148 7940 6204
rect 7996 6148 8082 6204
rect 8138 6148 8208 6204
rect 7868 6062 8208 6148
rect 7868 6006 7940 6062
rect 7996 6006 8082 6062
rect 8138 6006 8208 6062
rect 7868 5920 8208 6006
rect 7868 5864 7940 5920
rect 7996 5864 8082 5920
rect 8138 5864 8208 5920
rect 7868 5778 8208 5864
rect 7868 5722 7940 5778
rect 7996 5722 8082 5778
rect 8138 5722 8208 5778
rect 7868 5636 8208 5722
rect 7868 5580 7940 5636
rect 7996 5580 8082 5636
rect 8138 5580 8208 5636
rect 7868 5494 8208 5580
rect 7868 5438 7940 5494
rect 7996 5438 8082 5494
rect 8138 5438 8208 5494
rect 7868 5352 8208 5438
rect 7868 5296 7940 5352
rect 7996 5296 8082 5352
rect 8138 5296 8208 5352
rect 7868 5210 8208 5296
rect 7868 5154 7940 5210
rect 7996 5154 8082 5210
rect 8138 5154 8208 5210
rect 7868 5068 8208 5154
rect 7868 5012 7940 5068
rect 7996 5012 8082 5068
rect 8138 5012 8208 5068
rect 7868 4926 8208 5012
rect 7868 4870 7940 4926
rect 7996 4870 8082 4926
rect 8138 4870 8208 4926
rect 7868 4784 8208 4870
rect 7868 4728 7940 4784
rect 7996 4728 8082 4784
rect 8138 4728 8208 4784
rect 7868 4642 8208 4728
rect 7868 4586 7940 4642
rect 7996 4586 8082 4642
rect 8138 4586 8208 4642
rect 7868 4500 8208 4586
rect 7868 4444 7940 4500
rect 7996 4444 8082 4500
rect 8138 4444 8208 4500
rect 7868 4358 8208 4444
rect 7868 4302 7940 4358
rect 7996 4302 8082 4358
rect 8138 4302 8208 4358
rect 7868 4216 8208 4302
rect 7868 4160 7940 4216
rect 7996 4160 8082 4216
rect 8138 4160 8208 4216
rect 7868 4074 8208 4160
rect 7868 4018 7940 4074
rect 7996 4018 8082 4074
rect 8138 4018 8208 4074
rect 7868 3932 8208 4018
rect 7868 3876 7940 3932
rect 7996 3876 8082 3932
rect 8138 3876 8208 3932
rect 7868 3790 8208 3876
rect 7868 3734 7940 3790
rect 7996 3734 8082 3790
rect 8138 3734 8208 3790
rect 7868 3648 8208 3734
rect 7868 3592 7940 3648
rect 7996 3592 8082 3648
rect 8138 3592 8208 3648
rect 7868 3506 8208 3592
rect 7868 3450 7940 3506
rect 7996 3450 8082 3506
rect 8138 3450 8208 3506
rect 7868 3364 8208 3450
rect 7868 3308 7940 3364
rect 7996 3308 8082 3364
rect 8138 3308 8208 3364
rect 7868 3222 8208 3308
rect 7868 3166 7940 3222
rect 7996 3166 8082 3222
rect 8138 3166 8208 3222
rect 7868 3080 8208 3166
rect 7868 3024 7940 3080
rect 7996 3024 8082 3080
rect 8138 3024 8208 3080
rect 7868 2938 8208 3024
rect 7868 2882 7940 2938
rect 7996 2882 8082 2938
rect 8138 2882 8208 2938
rect 7868 2796 8208 2882
rect 7868 2740 7940 2796
rect 7996 2740 8082 2796
rect 8138 2740 8208 2796
rect 7868 2654 8208 2740
rect 7868 2598 7940 2654
rect 7996 2598 8082 2654
rect 8138 2598 8208 2654
rect 7868 2512 8208 2598
rect 7868 2456 7940 2512
rect 7996 2456 8082 2512
rect 8138 2456 8208 2512
rect 7868 2370 8208 2456
rect 7868 2314 7940 2370
rect 7996 2314 8082 2370
rect 8138 2314 8208 2370
rect 7868 2228 8208 2314
rect 7868 2172 7940 2228
rect 7996 2172 8082 2228
rect 8138 2172 8208 2228
rect 7868 2086 8208 2172
rect 7868 2030 7940 2086
rect 7996 2030 8082 2086
rect 8138 2030 8208 2086
rect 7868 1944 8208 2030
rect 7868 1888 7940 1944
rect 7996 1888 8082 1944
rect 8138 1888 8208 1944
rect 7868 1802 8208 1888
rect 7868 1746 7940 1802
rect 7996 1746 8082 1802
rect 8138 1746 8208 1802
rect 7868 1660 8208 1746
rect 7868 1604 7940 1660
rect 7996 1604 8082 1660
rect 8138 1604 8208 1660
rect 7868 1518 8208 1604
rect 7868 1462 7940 1518
rect 7996 1462 8082 1518
rect 8138 1462 8208 1518
rect 7868 1376 8208 1462
rect 7868 1320 7940 1376
rect 7996 1320 8082 1376
rect 8138 1320 8208 1376
rect 7868 1234 8208 1320
rect 7868 1178 7940 1234
rect 7996 1178 8082 1234
rect 8138 1178 8208 1234
rect 7868 1092 8208 1178
rect 7868 1036 7940 1092
rect 7996 1036 8082 1092
rect 8138 1036 8208 1092
rect 7868 950 8208 1036
rect 7868 894 7940 950
rect 7996 894 8082 950
rect 8138 894 8208 950
rect 7868 808 8208 894
rect 7868 752 7940 808
rect 7996 752 8082 808
rect 8138 752 8208 808
rect 7868 666 8208 752
rect 7868 610 7940 666
rect 7996 610 8082 666
rect 8138 610 8208 666
rect 7868 524 8208 610
rect 7868 468 7940 524
rect 7996 468 8082 524
rect 8138 468 8208 524
rect 7868 400 8208 468
rect 8268 12310 8608 12400
rect 8268 12254 8340 12310
rect 8396 12254 8482 12310
rect 8538 12254 8608 12310
rect 8268 12168 8608 12254
rect 8268 12112 8340 12168
rect 8396 12112 8482 12168
rect 8538 12112 8608 12168
rect 8268 12026 8608 12112
rect 8268 11970 8340 12026
rect 8396 11970 8482 12026
rect 8538 11970 8608 12026
rect 8268 11884 8608 11970
rect 8268 11828 8340 11884
rect 8396 11828 8482 11884
rect 8538 11828 8608 11884
rect 8268 11742 8608 11828
rect 8268 11686 8340 11742
rect 8396 11686 8482 11742
rect 8538 11686 8608 11742
rect 8268 11600 8608 11686
rect 8268 11544 8340 11600
rect 8396 11544 8482 11600
rect 8538 11544 8608 11600
rect 8268 11458 8608 11544
rect 8268 11402 8340 11458
rect 8396 11402 8482 11458
rect 8538 11402 8608 11458
rect 8268 11316 8608 11402
rect 8268 11260 8340 11316
rect 8396 11260 8482 11316
rect 8538 11260 8608 11316
rect 8268 11174 8608 11260
rect 8268 11118 8340 11174
rect 8396 11118 8482 11174
rect 8538 11118 8608 11174
rect 8268 11032 8608 11118
rect 8268 10976 8340 11032
rect 8396 10976 8482 11032
rect 8538 10976 8608 11032
rect 8268 10890 8608 10976
rect 8268 10834 8340 10890
rect 8396 10834 8482 10890
rect 8538 10834 8608 10890
rect 8268 10748 8608 10834
rect 8268 10692 8340 10748
rect 8396 10692 8482 10748
rect 8538 10692 8608 10748
rect 8268 10606 8608 10692
rect 8268 10550 8340 10606
rect 8396 10550 8482 10606
rect 8538 10550 8608 10606
rect 8268 10464 8608 10550
rect 8268 10408 8340 10464
rect 8396 10408 8482 10464
rect 8538 10408 8608 10464
rect 8268 10322 8608 10408
rect 8268 10266 8340 10322
rect 8396 10266 8482 10322
rect 8538 10266 8608 10322
rect 8268 10180 8608 10266
rect 8268 10124 8340 10180
rect 8396 10124 8482 10180
rect 8538 10124 8608 10180
rect 8268 10038 8608 10124
rect 8268 9982 8340 10038
rect 8396 9982 8482 10038
rect 8538 9982 8608 10038
rect 8268 9896 8608 9982
rect 8268 9840 8340 9896
rect 8396 9840 8482 9896
rect 8538 9840 8608 9896
rect 8268 9754 8608 9840
rect 8268 9698 8340 9754
rect 8396 9698 8482 9754
rect 8538 9698 8608 9754
rect 8268 9612 8608 9698
rect 8268 9556 8340 9612
rect 8396 9556 8482 9612
rect 8538 9556 8608 9612
rect 8268 9470 8608 9556
rect 8268 9414 8340 9470
rect 8396 9414 8482 9470
rect 8538 9414 8608 9470
rect 8268 9328 8608 9414
rect 8268 9272 8340 9328
rect 8396 9272 8482 9328
rect 8538 9272 8608 9328
rect 8268 9186 8608 9272
rect 8268 9130 8340 9186
rect 8396 9130 8482 9186
rect 8538 9130 8608 9186
rect 8268 9044 8608 9130
rect 8268 8988 8340 9044
rect 8396 8988 8482 9044
rect 8538 8988 8608 9044
rect 8268 8902 8608 8988
rect 8268 8846 8340 8902
rect 8396 8846 8482 8902
rect 8538 8846 8608 8902
rect 8268 8760 8608 8846
rect 8268 8704 8340 8760
rect 8396 8704 8482 8760
rect 8538 8704 8608 8760
rect 8268 8618 8608 8704
rect 8268 8562 8340 8618
rect 8396 8562 8482 8618
rect 8538 8562 8608 8618
rect 8268 8476 8608 8562
rect 8268 8420 8340 8476
rect 8396 8420 8482 8476
rect 8538 8420 8608 8476
rect 8268 8334 8608 8420
rect 8268 8278 8340 8334
rect 8396 8278 8482 8334
rect 8538 8278 8608 8334
rect 8268 8192 8608 8278
rect 8268 8136 8340 8192
rect 8396 8136 8482 8192
rect 8538 8136 8608 8192
rect 8268 8050 8608 8136
rect 8268 7994 8340 8050
rect 8396 7994 8482 8050
rect 8538 7994 8608 8050
rect 8268 7908 8608 7994
rect 8268 7852 8340 7908
rect 8396 7852 8482 7908
rect 8538 7852 8608 7908
rect 8268 7766 8608 7852
rect 8268 7710 8340 7766
rect 8396 7710 8482 7766
rect 8538 7710 8608 7766
rect 8268 7624 8608 7710
rect 8268 7568 8340 7624
rect 8396 7568 8482 7624
rect 8538 7568 8608 7624
rect 8268 7482 8608 7568
rect 8268 7426 8340 7482
rect 8396 7426 8482 7482
rect 8538 7426 8608 7482
rect 8268 7340 8608 7426
rect 8268 7284 8340 7340
rect 8396 7284 8482 7340
rect 8538 7284 8608 7340
rect 8268 7198 8608 7284
rect 8268 7142 8340 7198
rect 8396 7142 8482 7198
rect 8538 7142 8608 7198
rect 8268 7056 8608 7142
rect 8268 7000 8340 7056
rect 8396 7000 8482 7056
rect 8538 7000 8608 7056
rect 8268 6914 8608 7000
rect 8268 6858 8340 6914
rect 8396 6858 8482 6914
rect 8538 6858 8608 6914
rect 8268 6772 8608 6858
rect 8268 6716 8340 6772
rect 8396 6716 8482 6772
rect 8538 6716 8608 6772
rect 8268 6630 8608 6716
rect 8268 6574 8340 6630
rect 8396 6574 8482 6630
rect 8538 6574 8608 6630
rect 8268 6488 8608 6574
rect 8268 6432 8340 6488
rect 8396 6432 8482 6488
rect 8538 6432 8608 6488
rect 8268 6346 8608 6432
rect 8268 6290 8340 6346
rect 8396 6290 8482 6346
rect 8538 6290 8608 6346
rect 8268 6204 8608 6290
rect 8268 6148 8340 6204
rect 8396 6148 8482 6204
rect 8538 6148 8608 6204
rect 8268 6062 8608 6148
rect 8268 6006 8340 6062
rect 8396 6006 8482 6062
rect 8538 6006 8608 6062
rect 8268 5920 8608 6006
rect 8268 5864 8340 5920
rect 8396 5864 8482 5920
rect 8538 5864 8608 5920
rect 8268 5778 8608 5864
rect 8268 5722 8340 5778
rect 8396 5722 8482 5778
rect 8538 5722 8608 5778
rect 8268 5636 8608 5722
rect 8268 5580 8340 5636
rect 8396 5580 8482 5636
rect 8538 5580 8608 5636
rect 8268 5494 8608 5580
rect 8268 5438 8340 5494
rect 8396 5438 8482 5494
rect 8538 5438 8608 5494
rect 8268 5352 8608 5438
rect 8268 5296 8340 5352
rect 8396 5296 8482 5352
rect 8538 5296 8608 5352
rect 8268 5210 8608 5296
rect 8268 5154 8340 5210
rect 8396 5154 8482 5210
rect 8538 5154 8608 5210
rect 8268 5068 8608 5154
rect 8268 5012 8340 5068
rect 8396 5012 8482 5068
rect 8538 5012 8608 5068
rect 8268 4926 8608 5012
rect 8268 4870 8340 4926
rect 8396 4870 8482 4926
rect 8538 4870 8608 4926
rect 8268 4784 8608 4870
rect 8268 4728 8340 4784
rect 8396 4728 8482 4784
rect 8538 4728 8608 4784
rect 8268 4642 8608 4728
rect 8268 4586 8340 4642
rect 8396 4586 8482 4642
rect 8538 4586 8608 4642
rect 8268 4500 8608 4586
rect 8268 4444 8340 4500
rect 8396 4444 8482 4500
rect 8538 4444 8608 4500
rect 8268 4358 8608 4444
rect 8268 4302 8340 4358
rect 8396 4302 8482 4358
rect 8538 4302 8608 4358
rect 8268 4216 8608 4302
rect 8268 4160 8340 4216
rect 8396 4160 8482 4216
rect 8538 4160 8608 4216
rect 8268 4074 8608 4160
rect 8268 4018 8340 4074
rect 8396 4018 8482 4074
rect 8538 4018 8608 4074
rect 8268 3932 8608 4018
rect 8268 3876 8340 3932
rect 8396 3876 8482 3932
rect 8538 3876 8608 3932
rect 8268 3790 8608 3876
rect 8268 3734 8340 3790
rect 8396 3734 8482 3790
rect 8538 3734 8608 3790
rect 8268 3648 8608 3734
rect 8268 3592 8340 3648
rect 8396 3592 8482 3648
rect 8538 3592 8608 3648
rect 8268 3506 8608 3592
rect 8268 3450 8340 3506
rect 8396 3450 8482 3506
rect 8538 3450 8608 3506
rect 8268 3364 8608 3450
rect 8268 3308 8340 3364
rect 8396 3308 8482 3364
rect 8538 3308 8608 3364
rect 8268 3222 8608 3308
rect 8268 3166 8340 3222
rect 8396 3166 8482 3222
rect 8538 3166 8608 3222
rect 8268 3080 8608 3166
rect 8268 3024 8340 3080
rect 8396 3024 8482 3080
rect 8538 3024 8608 3080
rect 8268 2938 8608 3024
rect 8268 2882 8340 2938
rect 8396 2882 8482 2938
rect 8538 2882 8608 2938
rect 8268 2796 8608 2882
rect 8268 2740 8340 2796
rect 8396 2740 8482 2796
rect 8538 2740 8608 2796
rect 8268 2654 8608 2740
rect 8268 2598 8340 2654
rect 8396 2598 8482 2654
rect 8538 2598 8608 2654
rect 8268 2512 8608 2598
rect 8268 2456 8340 2512
rect 8396 2456 8482 2512
rect 8538 2456 8608 2512
rect 8268 2370 8608 2456
rect 8268 2314 8340 2370
rect 8396 2314 8482 2370
rect 8538 2314 8608 2370
rect 8268 2228 8608 2314
rect 8268 2172 8340 2228
rect 8396 2172 8482 2228
rect 8538 2172 8608 2228
rect 8268 2086 8608 2172
rect 8268 2030 8340 2086
rect 8396 2030 8482 2086
rect 8538 2030 8608 2086
rect 8268 1944 8608 2030
rect 8268 1888 8340 1944
rect 8396 1888 8482 1944
rect 8538 1888 8608 1944
rect 8268 1802 8608 1888
rect 8268 1746 8340 1802
rect 8396 1746 8482 1802
rect 8538 1746 8608 1802
rect 8268 1660 8608 1746
rect 8268 1604 8340 1660
rect 8396 1604 8482 1660
rect 8538 1604 8608 1660
rect 8268 1518 8608 1604
rect 8268 1462 8340 1518
rect 8396 1462 8482 1518
rect 8538 1462 8608 1518
rect 8268 1376 8608 1462
rect 8268 1320 8340 1376
rect 8396 1320 8482 1376
rect 8538 1320 8608 1376
rect 8268 1234 8608 1320
rect 8268 1178 8340 1234
rect 8396 1178 8482 1234
rect 8538 1178 8608 1234
rect 8268 1092 8608 1178
rect 8268 1036 8340 1092
rect 8396 1036 8482 1092
rect 8538 1036 8608 1092
rect 8268 950 8608 1036
rect 8268 894 8340 950
rect 8396 894 8482 950
rect 8538 894 8608 950
rect 8268 808 8608 894
rect 8268 752 8340 808
rect 8396 752 8482 808
rect 8538 752 8608 808
rect 8268 666 8608 752
rect 8268 610 8340 666
rect 8396 610 8482 666
rect 8538 610 8608 666
rect 8268 524 8608 610
rect 8268 468 8340 524
rect 8396 468 8482 524
rect 8538 468 8608 524
rect 8268 400 8608 468
rect 8668 12310 9008 12400
rect 8668 12254 8737 12310
rect 8793 12254 8879 12310
rect 8935 12254 9008 12310
rect 8668 12168 9008 12254
rect 8668 12112 8737 12168
rect 8793 12112 8879 12168
rect 8935 12112 9008 12168
rect 8668 12026 9008 12112
rect 8668 11970 8737 12026
rect 8793 11970 8879 12026
rect 8935 11970 9008 12026
rect 8668 11884 9008 11970
rect 8668 11828 8737 11884
rect 8793 11828 8879 11884
rect 8935 11828 9008 11884
rect 8668 11742 9008 11828
rect 8668 11686 8737 11742
rect 8793 11686 8879 11742
rect 8935 11686 9008 11742
rect 8668 11600 9008 11686
rect 8668 11544 8737 11600
rect 8793 11544 8879 11600
rect 8935 11544 9008 11600
rect 8668 11458 9008 11544
rect 8668 11402 8737 11458
rect 8793 11402 8879 11458
rect 8935 11402 9008 11458
rect 8668 11316 9008 11402
rect 8668 11260 8737 11316
rect 8793 11260 8879 11316
rect 8935 11260 9008 11316
rect 8668 11174 9008 11260
rect 8668 11118 8737 11174
rect 8793 11118 8879 11174
rect 8935 11118 9008 11174
rect 8668 11032 9008 11118
rect 8668 10976 8737 11032
rect 8793 10976 8879 11032
rect 8935 10976 9008 11032
rect 8668 10890 9008 10976
rect 8668 10834 8737 10890
rect 8793 10834 8879 10890
rect 8935 10834 9008 10890
rect 8668 10748 9008 10834
rect 8668 10692 8737 10748
rect 8793 10692 8879 10748
rect 8935 10692 9008 10748
rect 8668 10606 9008 10692
rect 8668 10550 8737 10606
rect 8793 10550 8879 10606
rect 8935 10550 9008 10606
rect 8668 10464 9008 10550
rect 8668 10408 8737 10464
rect 8793 10408 8879 10464
rect 8935 10408 9008 10464
rect 8668 10322 9008 10408
rect 8668 10266 8737 10322
rect 8793 10266 8879 10322
rect 8935 10266 9008 10322
rect 8668 10180 9008 10266
rect 8668 10124 8737 10180
rect 8793 10124 8879 10180
rect 8935 10124 9008 10180
rect 8668 10038 9008 10124
rect 8668 9982 8737 10038
rect 8793 9982 8879 10038
rect 8935 9982 9008 10038
rect 8668 9896 9008 9982
rect 8668 9840 8737 9896
rect 8793 9840 8879 9896
rect 8935 9840 9008 9896
rect 8668 9754 9008 9840
rect 8668 9698 8737 9754
rect 8793 9698 8879 9754
rect 8935 9698 9008 9754
rect 8668 9612 9008 9698
rect 8668 9556 8737 9612
rect 8793 9556 8879 9612
rect 8935 9556 9008 9612
rect 8668 9470 9008 9556
rect 8668 9414 8737 9470
rect 8793 9414 8879 9470
rect 8935 9414 9008 9470
rect 8668 9328 9008 9414
rect 8668 9272 8737 9328
rect 8793 9272 8879 9328
rect 8935 9272 9008 9328
rect 8668 9186 9008 9272
rect 8668 9130 8737 9186
rect 8793 9130 8879 9186
rect 8935 9130 9008 9186
rect 8668 9044 9008 9130
rect 8668 8988 8737 9044
rect 8793 8988 8879 9044
rect 8935 8988 9008 9044
rect 8668 8902 9008 8988
rect 8668 8846 8737 8902
rect 8793 8846 8879 8902
rect 8935 8846 9008 8902
rect 8668 8760 9008 8846
rect 8668 8704 8737 8760
rect 8793 8704 8879 8760
rect 8935 8704 9008 8760
rect 8668 8618 9008 8704
rect 8668 8562 8737 8618
rect 8793 8562 8879 8618
rect 8935 8562 9008 8618
rect 8668 8476 9008 8562
rect 8668 8420 8737 8476
rect 8793 8420 8879 8476
rect 8935 8420 9008 8476
rect 8668 8334 9008 8420
rect 8668 8278 8737 8334
rect 8793 8278 8879 8334
rect 8935 8278 9008 8334
rect 8668 8192 9008 8278
rect 8668 8136 8737 8192
rect 8793 8136 8879 8192
rect 8935 8136 9008 8192
rect 8668 8050 9008 8136
rect 8668 7994 8737 8050
rect 8793 7994 8879 8050
rect 8935 7994 9008 8050
rect 8668 7908 9008 7994
rect 8668 7852 8737 7908
rect 8793 7852 8879 7908
rect 8935 7852 9008 7908
rect 8668 7766 9008 7852
rect 8668 7710 8737 7766
rect 8793 7710 8879 7766
rect 8935 7710 9008 7766
rect 8668 7624 9008 7710
rect 8668 7568 8737 7624
rect 8793 7568 8879 7624
rect 8935 7568 9008 7624
rect 8668 7482 9008 7568
rect 8668 7426 8737 7482
rect 8793 7426 8879 7482
rect 8935 7426 9008 7482
rect 8668 7340 9008 7426
rect 8668 7284 8737 7340
rect 8793 7284 8879 7340
rect 8935 7284 9008 7340
rect 8668 7198 9008 7284
rect 8668 7142 8737 7198
rect 8793 7142 8879 7198
rect 8935 7142 9008 7198
rect 8668 7056 9008 7142
rect 8668 7000 8737 7056
rect 8793 7000 8879 7056
rect 8935 7000 9008 7056
rect 8668 6914 9008 7000
rect 8668 6858 8737 6914
rect 8793 6858 8879 6914
rect 8935 6858 9008 6914
rect 8668 6772 9008 6858
rect 8668 6716 8737 6772
rect 8793 6716 8879 6772
rect 8935 6716 9008 6772
rect 8668 6630 9008 6716
rect 8668 6574 8737 6630
rect 8793 6574 8879 6630
rect 8935 6574 9008 6630
rect 8668 6488 9008 6574
rect 8668 6432 8737 6488
rect 8793 6432 8879 6488
rect 8935 6432 9008 6488
rect 8668 6346 9008 6432
rect 8668 6290 8737 6346
rect 8793 6290 8879 6346
rect 8935 6290 9008 6346
rect 8668 6204 9008 6290
rect 8668 6148 8737 6204
rect 8793 6148 8879 6204
rect 8935 6148 9008 6204
rect 8668 6062 9008 6148
rect 8668 6006 8737 6062
rect 8793 6006 8879 6062
rect 8935 6006 9008 6062
rect 8668 5920 9008 6006
rect 8668 5864 8737 5920
rect 8793 5864 8879 5920
rect 8935 5864 9008 5920
rect 8668 5778 9008 5864
rect 8668 5722 8737 5778
rect 8793 5722 8879 5778
rect 8935 5722 9008 5778
rect 8668 5636 9008 5722
rect 8668 5580 8737 5636
rect 8793 5580 8879 5636
rect 8935 5580 9008 5636
rect 8668 5494 9008 5580
rect 8668 5438 8737 5494
rect 8793 5438 8879 5494
rect 8935 5438 9008 5494
rect 8668 5352 9008 5438
rect 8668 5296 8737 5352
rect 8793 5296 8879 5352
rect 8935 5296 9008 5352
rect 8668 5210 9008 5296
rect 8668 5154 8737 5210
rect 8793 5154 8879 5210
rect 8935 5154 9008 5210
rect 8668 5068 9008 5154
rect 8668 5012 8737 5068
rect 8793 5012 8879 5068
rect 8935 5012 9008 5068
rect 8668 4926 9008 5012
rect 8668 4870 8737 4926
rect 8793 4870 8879 4926
rect 8935 4870 9008 4926
rect 8668 4784 9008 4870
rect 8668 4728 8737 4784
rect 8793 4728 8879 4784
rect 8935 4728 9008 4784
rect 8668 4642 9008 4728
rect 8668 4586 8737 4642
rect 8793 4586 8879 4642
rect 8935 4586 9008 4642
rect 8668 4500 9008 4586
rect 8668 4444 8737 4500
rect 8793 4444 8879 4500
rect 8935 4444 9008 4500
rect 8668 4358 9008 4444
rect 8668 4302 8737 4358
rect 8793 4302 8879 4358
rect 8935 4302 9008 4358
rect 8668 4216 9008 4302
rect 8668 4160 8737 4216
rect 8793 4160 8879 4216
rect 8935 4160 9008 4216
rect 8668 4074 9008 4160
rect 8668 4018 8737 4074
rect 8793 4018 8879 4074
rect 8935 4018 9008 4074
rect 8668 3932 9008 4018
rect 8668 3876 8737 3932
rect 8793 3876 8879 3932
rect 8935 3876 9008 3932
rect 8668 3790 9008 3876
rect 8668 3734 8737 3790
rect 8793 3734 8879 3790
rect 8935 3734 9008 3790
rect 8668 3648 9008 3734
rect 8668 3592 8737 3648
rect 8793 3592 8879 3648
rect 8935 3592 9008 3648
rect 8668 3506 9008 3592
rect 8668 3450 8737 3506
rect 8793 3450 8879 3506
rect 8935 3450 9008 3506
rect 8668 3364 9008 3450
rect 8668 3308 8737 3364
rect 8793 3308 8879 3364
rect 8935 3308 9008 3364
rect 8668 3222 9008 3308
rect 8668 3166 8737 3222
rect 8793 3166 8879 3222
rect 8935 3166 9008 3222
rect 8668 3080 9008 3166
rect 8668 3024 8737 3080
rect 8793 3024 8879 3080
rect 8935 3024 9008 3080
rect 8668 2938 9008 3024
rect 8668 2882 8737 2938
rect 8793 2882 8879 2938
rect 8935 2882 9008 2938
rect 8668 2796 9008 2882
rect 8668 2740 8737 2796
rect 8793 2740 8879 2796
rect 8935 2740 9008 2796
rect 8668 2654 9008 2740
rect 8668 2598 8737 2654
rect 8793 2598 8879 2654
rect 8935 2598 9008 2654
rect 8668 2512 9008 2598
rect 8668 2456 8737 2512
rect 8793 2456 8879 2512
rect 8935 2456 9008 2512
rect 8668 2370 9008 2456
rect 8668 2314 8737 2370
rect 8793 2314 8879 2370
rect 8935 2314 9008 2370
rect 8668 2228 9008 2314
rect 8668 2172 8737 2228
rect 8793 2172 8879 2228
rect 8935 2172 9008 2228
rect 8668 2086 9008 2172
rect 8668 2030 8737 2086
rect 8793 2030 8879 2086
rect 8935 2030 9008 2086
rect 8668 1944 9008 2030
rect 8668 1888 8737 1944
rect 8793 1888 8879 1944
rect 8935 1888 9008 1944
rect 8668 1802 9008 1888
rect 8668 1746 8737 1802
rect 8793 1746 8879 1802
rect 8935 1746 9008 1802
rect 8668 1660 9008 1746
rect 8668 1604 8737 1660
rect 8793 1604 8879 1660
rect 8935 1604 9008 1660
rect 8668 1518 9008 1604
rect 8668 1462 8737 1518
rect 8793 1462 8879 1518
rect 8935 1462 9008 1518
rect 8668 1376 9008 1462
rect 8668 1320 8737 1376
rect 8793 1320 8879 1376
rect 8935 1320 9008 1376
rect 8668 1234 9008 1320
rect 8668 1178 8737 1234
rect 8793 1178 8879 1234
rect 8935 1178 9008 1234
rect 8668 1092 9008 1178
rect 8668 1036 8737 1092
rect 8793 1036 8879 1092
rect 8935 1036 9008 1092
rect 8668 950 9008 1036
rect 8668 894 8737 950
rect 8793 894 8879 950
rect 8935 894 9008 950
rect 8668 808 9008 894
rect 8668 752 8737 808
rect 8793 752 8879 808
rect 8935 752 9008 808
rect 8668 666 9008 752
rect 8668 610 8737 666
rect 8793 610 8879 666
rect 8935 610 9008 666
rect 8668 524 9008 610
rect 8668 468 8737 524
rect 8793 468 8879 524
rect 8935 468 9008 524
rect 8668 400 9008 468
rect 9068 12310 9408 12400
rect 9068 12254 9134 12310
rect 9190 12254 9276 12310
rect 9332 12254 9408 12310
rect 9068 12168 9408 12254
rect 9068 12112 9134 12168
rect 9190 12112 9276 12168
rect 9332 12112 9408 12168
rect 9068 12026 9408 12112
rect 9068 11970 9134 12026
rect 9190 11970 9276 12026
rect 9332 11970 9408 12026
rect 9068 11884 9408 11970
rect 9068 11828 9134 11884
rect 9190 11828 9276 11884
rect 9332 11828 9408 11884
rect 9068 11742 9408 11828
rect 9068 11686 9134 11742
rect 9190 11686 9276 11742
rect 9332 11686 9408 11742
rect 9068 11600 9408 11686
rect 9068 11544 9134 11600
rect 9190 11544 9276 11600
rect 9332 11544 9408 11600
rect 9068 11458 9408 11544
rect 9068 11402 9134 11458
rect 9190 11402 9276 11458
rect 9332 11402 9408 11458
rect 9068 11316 9408 11402
rect 9068 11260 9134 11316
rect 9190 11260 9276 11316
rect 9332 11260 9408 11316
rect 9068 11174 9408 11260
rect 9068 11118 9134 11174
rect 9190 11118 9276 11174
rect 9332 11118 9408 11174
rect 9068 11032 9408 11118
rect 9068 10976 9134 11032
rect 9190 10976 9276 11032
rect 9332 10976 9408 11032
rect 9068 10890 9408 10976
rect 9068 10834 9134 10890
rect 9190 10834 9276 10890
rect 9332 10834 9408 10890
rect 9068 10748 9408 10834
rect 9068 10692 9134 10748
rect 9190 10692 9276 10748
rect 9332 10692 9408 10748
rect 9068 10606 9408 10692
rect 9068 10550 9134 10606
rect 9190 10550 9276 10606
rect 9332 10550 9408 10606
rect 9068 10464 9408 10550
rect 9068 10408 9134 10464
rect 9190 10408 9276 10464
rect 9332 10408 9408 10464
rect 9068 10322 9408 10408
rect 9068 10266 9134 10322
rect 9190 10266 9276 10322
rect 9332 10266 9408 10322
rect 9068 10180 9408 10266
rect 9068 10124 9134 10180
rect 9190 10124 9276 10180
rect 9332 10124 9408 10180
rect 9068 10038 9408 10124
rect 9068 9982 9134 10038
rect 9190 9982 9276 10038
rect 9332 9982 9408 10038
rect 9068 9896 9408 9982
rect 9068 9840 9134 9896
rect 9190 9840 9276 9896
rect 9332 9840 9408 9896
rect 9068 9754 9408 9840
rect 9068 9698 9134 9754
rect 9190 9698 9276 9754
rect 9332 9698 9408 9754
rect 9068 9612 9408 9698
rect 9068 9556 9134 9612
rect 9190 9556 9276 9612
rect 9332 9556 9408 9612
rect 9068 9470 9408 9556
rect 9068 9414 9134 9470
rect 9190 9414 9276 9470
rect 9332 9414 9408 9470
rect 9068 9328 9408 9414
rect 9068 9272 9134 9328
rect 9190 9272 9276 9328
rect 9332 9272 9408 9328
rect 9068 9186 9408 9272
rect 9068 9130 9134 9186
rect 9190 9130 9276 9186
rect 9332 9130 9408 9186
rect 9068 9044 9408 9130
rect 9068 8988 9134 9044
rect 9190 8988 9276 9044
rect 9332 8988 9408 9044
rect 9068 8902 9408 8988
rect 9068 8846 9134 8902
rect 9190 8846 9276 8902
rect 9332 8846 9408 8902
rect 9068 8760 9408 8846
rect 9068 8704 9134 8760
rect 9190 8704 9276 8760
rect 9332 8704 9408 8760
rect 9068 8618 9408 8704
rect 9068 8562 9134 8618
rect 9190 8562 9276 8618
rect 9332 8562 9408 8618
rect 9068 8476 9408 8562
rect 9068 8420 9134 8476
rect 9190 8420 9276 8476
rect 9332 8420 9408 8476
rect 9068 8334 9408 8420
rect 9068 8278 9134 8334
rect 9190 8278 9276 8334
rect 9332 8278 9408 8334
rect 9068 8192 9408 8278
rect 9068 8136 9134 8192
rect 9190 8136 9276 8192
rect 9332 8136 9408 8192
rect 9068 8050 9408 8136
rect 9068 7994 9134 8050
rect 9190 7994 9276 8050
rect 9332 7994 9408 8050
rect 9068 7908 9408 7994
rect 9068 7852 9134 7908
rect 9190 7852 9276 7908
rect 9332 7852 9408 7908
rect 9068 7766 9408 7852
rect 9068 7710 9134 7766
rect 9190 7710 9276 7766
rect 9332 7710 9408 7766
rect 9068 7624 9408 7710
rect 9068 7568 9134 7624
rect 9190 7568 9276 7624
rect 9332 7568 9408 7624
rect 9068 7482 9408 7568
rect 9068 7426 9134 7482
rect 9190 7426 9276 7482
rect 9332 7426 9408 7482
rect 9068 7340 9408 7426
rect 9068 7284 9134 7340
rect 9190 7284 9276 7340
rect 9332 7284 9408 7340
rect 9068 7198 9408 7284
rect 9068 7142 9134 7198
rect 9190 7142 9276 7198
rect 9332 7142 9408 7198
rect 9068 7056 9408 7142
rect 9068 7000 9134 7056
rect 9190 7000 9276 7056
rect 9332 7000 9408 7056
rect 9068 6914 9408 7000
rect 9068 6858 9134 6914
rect 9190 6858 9276 6914
rect 9332 6858 9408 6914
rect 9068 6772 9408 6858
rect 9068 6716 9134 6772
rect 9190 6716 9276 6772
rect 9332 6716 9408 6772
rect 9068 6630 9408 6716
rect 9068 6574 9134 6630
rect 9190 6574 9276 6630
rect 9332 6574 9408 6630
rect 9068 6488 9408 6574
rect 9068 6432 9134 6488
rect 9190 6432 9276 6488
rect 9332 6432 9408 6488
rect 9068 6346 9408 6432
rect 9068 6290 9134 6346
rect 9190 6290 9276 6346
rect 9332 6290 9408 6346
rect 9068 6204 9408 6290
rect 9068 6148 9134 6204
rect 9190 6148 9276 6204
rect 9332 6148 9408 6204
rect 9068 6062 9408 6148
rect 9068 6006 9134 6062
rect 9190 6006 9276 6062
rect 9332 6006 9408 6062
rect 9068 5920 9408 6006
rect 9068 5864 9134 5920
rect 9190 5864 9276 5920
rect 9332 5864 9408 5920
rect 9068 5778 9408 5864
rect 9068 5722 9134 5778
rect 9190 5722 9276 5778
rect 9332 5722 9408 5778
rect 9068 5636 9408 5722
rect 9068 5580 9134 5636
rect 9190 5580 9276 5636
rect 9332 5580 9408 5636
rect 9068 5494 9408 5580
rect 9068 5438 9134 5494
rect 9190 5438 9276 5494
rect 9332 5438 9408 5494
rect 9068 5352 9408 5438
rect 9068 5296 9134 5352
rect 9190 5296 9276 5352
rect 9332 5296 9408 5352
rect 9068 5210 9408 5296
rect 9068 5154 9134 5210
rect 9190 5154 9276 5210
rect 9332 5154 9408 5210
rect 9068 5068 9408 5154
rect 9068 5012 9134 5068
rect 9190 5012 9276 5068
rect 9332 5012 9408 5068
rect 9068 4926 9408 5012
rect 9068 4870 9134 4926
rect 9190 4870 9276 4926
rect 9332 4870 9408 4926
rect 9068 4784 9408 4870
rect 9068 4728 9134 4784
rect 9190 4728 9276 4784
rect 9332 4728 9408 4784
rect 9068 4642 9408 4728
rect 9068 4586 9134 4642
rect 9190 4586 9276 4642
rect 9332 4586 9408 4642
rect 9068 4500 9408 4586
rect 9068 4444 9134 4500
rect 9190 4444 9276 4500
rect 9332 4444 9408 4500
rect 9068 4358 9408 4444
rect 9068 4302 9134 4358
rect 9190 4302 9276 4358
rect 9332 4302 9408 4358
rect 9068 4216 9408 4302
rect 9068 4160 9134 4216
rect 9190 4160 9276 4216
rect 9332 4160 9408 4216
rect 9068 4074 9408 4160
rect 9068 4018 9134 4074
rect 9190 4018 9276 4074
rect 9332 4018 9408 4074
rect 9068 3932 9408 4018
rect 9068 3876 9134 3932
rect 9190 3876 9276 3932
rect 9332 3876 9408 3932
rect 9068 3790 9408 3876
rect 9068 3734 9134 3790
rect 9190 3734 9276 3790
rect 9332 3734 9408 3790
rect 9068 3648 9408 3734
rect 9068 3592 9134 3648
rect 9190 3592 9276 3648
rect 9332 3592 9408 3648
rect 9068 3506 9408 3592
rect 9068 3450 9134 3506
rect 9190 3450 9276 3506
rect 9332 3450 9408 3506
rect 9068 3364 9408 3450
rect 9068 3308 9134 3364
rect 9190 3308 9276 3364
rect 9332 3308 9408 3364
rect 9068 3222 9408 3308
rect 9068 3166 9134 3222
rect 9190 3166 9276 3222
rect 9332 3166 9408 3222
rect 9068 3080 9408 3166
rect 9068 3024 9134 3080
rect 9190 3024 9276 3080
rect 9332 3024 9408 3080
rect 9068 2938 9408 3024
rect 9068 2882 9134 2938
rect 9190 2882 9276 2938
rect 9332 2882 9408 2938
rect 9068 2796 9408 2882
rect 9068 2740 9134 2796
rect 9190 2740 9276 2796
rect 9332 2740 9408 2796
rect 9068 2654 9408 2740
rect 9068 2598 9134 2654
rect 9190 2598 9276 2654
rect 9332 2598 9408 2654
rect 9068 2512 9408 2598
rect 9068 2456 9134 2512
rect 9190 2456 9276 2512
rect 9332 2456 9408 2512
rect 9068 2370 9408 2456
rect 9068 2314 9134 2370
rect 9190 2314 9276 2370
rect 9332 2314 9408 2370
rect 9068 2228 9408 2314
rect 9068 2172 9134 2228
rect 9190 2172 9276 2228
rect 9332 2172 9408 2228
rect 9068 2086 9408 2172
rect 9068 2030 9134 2086
rect 9190 2030 9276 2086
rect 9332 2030 9408 2086
rect 9068 1944 9408 2030
rect 9068 1888 9134 1944
rect 9190 1888 9276 1944
rect 9332 1888 9408 1944
rect 9068 1802 9408 1888
rect 9068 1746 9134 1802
rect 9190 1746 9276 1802
rect 9332 1746 9408 1802
rect 9068 1660 9408 1746
rect 9068 1604 9134 1660
rect 9190 1604 9276 1660
rect 9332 1604 9408 1660
rect 9068 1518 9408 1604
rect 9068 1462 9134 1518
rect 9190 1462 9276 1518
rect 9332 1462 9408 1518
rect 9068 1376 9408 1462
rect 9068 1320 9134 1376
rect 9190 1320 9276 1376
rect 9332 1320 9408 1376
rect 9068 1234 9408 1320
rect 9068 1178 9134 1234
rect 9190 1178 9276 1234
rect 9332 1178 9408 1234
rect 9068 1092 9408 1178
rect 9068 1036 9134 1092
rect 9190 1036 9276 1092
rect 9332 1036 9408 1092
rect 9068 950 9408 1036
rect 9068 894 9134 950
rect 9190 894 9276 950
rect 9332 894 9408 950
rect 9068 808 9408 894
rect 9068 752 9134 808
rect 9190 752 9276 808
rect 9332 752 9408 808
rect 9068 666 9408 752
rect 9068 610 9134 666
rect 9190 610 9276 666
rect 9332 610 9408 666
rect 9068 524 9408 610
rect 9068 468 9134 524
rect 9190 468 9276 524
rect 9332 468 9408 524
rect 9068 400 9408 468
rect 9468 12310 9808 12400
rect 9468 12254 9538 12310
rect 9594 12254 9680 12310
rect 9736 12254 9808 12310
rect 9468 12168 9808 12254
rect 9468 12112 9538 12168
rect 9594 12112 9680 12168
rect 9736 12112 9808 12168
rect 9468 12026 9808 12112
rect 9468 11970 9538 12026
rect 9594 11970 9680 12026
rect 9736 11970 9808 12026
rect 9468 11884 9808 11970
rect 9468 11828 9538 11884
rect 9594 11828 9680 11884
rect 9736 11828 9808 11884
rect 9468 11742 9808 11828
rect 9468 11686 9538 11742
rect 9594 11686 9680 11742
rect 9736 11686 9808 11742
rect 9468 11600 9808 11686
rect 9468 11544 9538 11600
rect 9594 11544 9680 11600
rect 9736 11544 9808 11600
rect 9468 11458 9808 11544
rect 9468 11402 9538 11458
rect 9594 11402 9680 11458
rect 9736 11402 9808 11458
rect 9468 11316 9808 11402
rect 9468 11260 9538 11316
rect 9594 11260 9680 11316
rect 9736 11260 9808 11316
rect 9468 11174 9808 11260
rect 9468 11118 9538 11174
rect 9594 11118 9680 11174
rect 9736 11118 9808 11174
rect 9468 11032 9808 11118
rect 9468 10976 9538 11032
rect 9594 10976 9680 11032
rect 9736 10976 9808 11032
rect 9468 10890 9808 10976
rect 9468 10834 9538 10890
rect 9594 10834 9680 10890
rect 9736 10834 9808 10890
rect 9468 10748 9808 10834
rect 9468 10692 9538 10748
rect 9594 10692 9680 10748
rect 9736 10692 9808 10748
rect 9468 10606 9808 10692
rect 9468 10550 9538 10606
rect 9594 10550 9680 10606
rect 9736 10550 9808 10606
rect 9468 10464 9808 10550
rect 9468 10408 9538 10464
rect 9594 10408 9680 10464
rect 9736 10408 9808 10464
rect 9468 10322 9808 10408
rect 9468 10266 9538 10322
rect 9594 10266 9680 10322
rect 9736 10266 9808 10322
rect 9468 10180 9808 10266
rect 9468 10124 9538 10180
rect 9594 10124 9680 10180
rect 9736 10124 9808 10180
rect 9468 10038 9808 10124
rect 9468 9982 9538 10038
rect 9594 9982 9680 10038
rect 9736 9982 9808 10038
rect 9468 9896 9808 9982
rect 9468 9840 9538 9896
rect 9594 9840 9680 9896
rect 9736 9840 9808 9896
rect 9468 9754 9808 9840
rect 9468 9698 9538 9754
rect 9594 9698 9680 9754
rect 9736 9698 9808 9754
rect 9468 9612 9808 9698
rect 9468 9556 9538 9612
rect 9594 9556 9680 9612
rect 9736 9556 9808 9612
rect 9468 9470 9808 9556
rect 9468 9414 9538 9470
rect 9594 9414 9680 9470
rect 9736 9414 9808 9470
rect 9468 9328 9808 9414
rect 9468 9272 9538 9328
rect 9594 9272 9680 9328
rect 9736 9272 9808 9328
rect 9468 9186 9808 9272
rect 9468 9130 9538 9186
rect 9594 9130 9680 9186
rect 9736 9130 9808 9186
rect 9468 9044 9808 9130
rect 9468 8988 9538 9044
rect 9594 8988 9680 9044
rect 9736 8988 9808 9044
rect 9468 8902 9808 8988
rect 9468 8846 9538 8902
rect 9594 8846 9680 8902
rect 9736 8846 9808 8902
rect 9468 8760 9808 8846
rect 9468 8704 9538 8760
rect 9594 8704 9680 8760
rect 9736 8704 9808 8760
rect 9468 8618 9808 8704
rect 9468 8562 9538 8618
rect 9594 8562 9680 8618
rect 9736 8562 9808 8618
rect 9468 8476 9808 8562
rect 9468 8420 9538 8476
rect 9594 8420 9680 8476
rect 9736 8420 9808 8476
rect 9468 8334 9808 8420
rect 9468 8278 9538 8334
rect 9594 8278 9680 8334
rect 9736 8278 9808 8334
rect 9468 8192 9808 8278
rect 9468 8136 9538 8192
rect 9594 8136 9680 8192
rect 9736 8136 9808 8192
rect 9468 8050 9808 8136
rect 9468 7994 9538 8050
rect 9594 7994 9680 8050
rect 9736 7994 9808 8050
rect 9468 7908 9808 7994
rect 9468 7852 9538 7908
rect 9594 7852 9680 7908
rect 9736 7852 9808 7908
rect 9468 7766 9808 7852
rect 9468 7710 9538 7766
rect 9594 7710 9680 7766
rect 9736 7710 9808 7766
rect 9468 7624 9808 7710
rect 9468 7568 9538 7624
rect 9594 7568 9680 7624
rect 9736 7568 9808 7624
rect 9468 7482 9808 7568
rect 9468 7426 9538 7482
rect 9594 7426 9680 7482
rect 9736 7426 9808 7482
rect 9468 7340 9808 7426
rect 9468 7284 9538 7340
rect 9594 7284 9680 7340
rect 9736 7284 9808 7340
rect 9468 7198 9808 7284
rect 9468 7142 9538 7198
rect 9594 7142 9680 7198
rect 9736 7142 9808 7198
rect 9468 7056 9808 7142
rect 9468 7000 9538 7056
rect 9594 7000 9680 7056
rect 9736 7000 9808 7056
rect 9468 6914 9808 7000
rect 9468 6858 9538 6914
rect 9594 6858 9680 6914
rect 9736 6858 9808 6914
rect 9468 6772 9808 6858
rect 9468 6716 9538 6772
rect 9594 6716 9680 6772
rect 9736 6716 9808 6772
rect 9468 6630 9808 6716
rect 9468 6574 9538 6630
rect 9594 6574 9680 6630
rect 9736 6574 9808 6630
rect 9468 6488 9808 6574
rect 9468 6432 9538 6488
rect 9594 6432 9680 6488
rect 9736 6432 9808 6488
rect 9468 6346 9808 6432
rect 9468 6290 9538 6346
rect 9594 6290 9680 6346
rect 9736 6290 9808 6346
rect 9468 6204 9808 6290
rect 9468 6148 9538 6204
rect 9594 6148 9680 6204
rect 9736 6148 9808 6204
rect 9468 6062 9808 6148
rect 9468 6006 9538 6062
rect 9594 6006 9680 6062
rect 9736 6006 9808 6062
rect 9468 5920 9808 6006
rect 9468 5864 9538 5920
rect 9594 5864 9680 5920
rect 9736 5864 9808 5920
rect 9468 5778 9808 5864
rect 9468 5722 9538 5778
rect 9594 5722 9680 5778
rect 9736 5722 9808 5778
rect 9468 5636 9808 5722
rect 9468 5580 9538 5636
rect 9594 5580 9680 5636
rect 9736 5580 9808 5636
rect 9468 5494 9808 5580
rect 9468 5438 9538 5494
rect 9594 5438 9680 5494
rect 9736 5438 9808 5494
rect 9468 5352 9808 5438
rect 9468 5296 9538 5352
rect 9594 5296 9680 5352
rect 9736 5296 9808 5352
rect 9468 5210 9808 5296
rect 9468 5154 9538 5210
rect 9594 5154 9680 5210
rect 9736 5154 9808 5210
rect 9468 5068 9808 5154
rect 9468 5012 9538 5068
rect 9594 5012 9680 5068
rect 9736 5012 9808 5068
rect 9468 4926 9808 5012
rect 9468 4870 9538 4926
rect 9594 4870 9680 4926
rect 9736 4870 9808 4926
rect 9468 4784 9808 4870
rect 9468 4728 9538 4784
rect 9594 4728 9680 4784
rect 9736 4728 9808 4784
rect 9468 4642 9808 4728
rect 9468 4586 9538 4642
rect 9594 4586 9680 4642
rect 9736 4586 9808 4642
rect 9468 4500 9808 4586
rect 9468 4444 9538 4500
rect 9594 4444 9680 4500
rect 9736 4444 9808 4500
rect 9468 4358 9808 4444
rect 9468 4302 9538 4358
rect 9594 4302 9680 4358
rect 9736 4302 9808 4358
rect 9468 4216 9808 4302
rect 9468 4160 9538 4216
rect 9594 4160 9680 4216
rect 9736 4160 9808 4216
rect 9468 4074 9808 4160
rect 9468 4018 9538 4074
rect 9594 4018 9680 4074
rect 9736 4018 9808 4074
rect 9468 3932 9808 4018
rect 9468 3876 9538 3932
rect 9594 3876 9680 3932
rect 9736 3876 9808 3932
rect 9468 3790 9808 3876
rect 9468 3734 9538 3790
rect 9594 3734 9680 3790
rect 9736 3734 9808 3790
rect 9468 3648 9808 3734
rect 9468 3592 9538 3648
rect 9594 3592 9680 3648
rect 9736 3592 9808 3648
rect 9468 3506 9808 3592
rect 9468 3450 9538 3506
rect 9594 3450 9680 3506
rect 9736 3450 9808 3506
rect 9468 3364 9808 3450
rect 9468 3308 9538 3364
rect 9594 3308 9680 3364
rect 9736 3308 9808 3364
rect 9468 3222 9808 3308
rect 9468 3166 9538 3222
rect 9594 3166 9680 3222
rect 9736 3166 9808 3222
rect 9468 3080 9808 3166
rect 9468 3024 9538 3080
rect 9594 3024 9680 3080
rect 9736 3024 9808 3080
rect 9468 2938 9808 3024
rect 9468 2882 9538 2938
rect 9594 2882 9680 2938
rect 9736 2882 9808 2938
rect 9468 2796 9808 2882
rect 9468 2740 9538 2796
rect 9594 2740 9680 2796
rect 9736 2740 9808 2796
rect 9468 2654 9808 2740
rect 9468 2598 9538 2654
rect 9594 2598 9680 2654
rect 9736 2598 9808 2654
rect 9468 2512 9808 2598
rect 9468 2456 9538 2512
rect 9594 2456 9680 2512
rect 9736 2456 9808 2512
rect 9468 2370 9808 2456
rect 9468 2314 9538 2370
rect 9594 2314 9680 2370
rect 9736 2314 9808 2370
rect 9468 2228 9808 2314
rect 9468 2172 9538 2228
rect 9594 2172 9680 2228
rect 9736 2172 9808 2228
rect 9468 2086 9808 2172
rect 9468 2030 9538 2086
rect 9594 2030 9680 2086
rect 9736 2030 9808 2086
rect 9468 1944 9808 2030
rect 9468 1888 9538 1944
rect 9594 1888 9680 1944
rect 9736 1888 9808 1944
rect 9468 1802 9808 1888
rect 9468 1746 9538 1802
rect 9594 1746 9680 1802
rect 9736 1746 9808 1802
rect 9468 1660 9808 1746
rect 9468 1604 9538 1660
rect 9594 1604 9680 1660
rect 9736 1604 9808 1660
rect 9468 1518 9808 1604
rect 9468 1462 9538 1518
rect 9594 1462 9680 1518
rect 9736 1462 9808 1518
rect 9468 1376 9808 1462
rect 9468 1320 9538 1376
rect 9594 1320 9680 1376
rect 9736 1320 9808 1376
rect 9468 1234 9808 1320
rect 9468 1178 9538 1234
rect 9594 1178 9680 1234
rect 9736 1178 9808 1234
rect 9468 1092 9808 1178
rect 9468 1036 9538 1092
rect 9594 1036 9680 1092
rect 9736 1036 9808 1092
rect 9468 950 9808 1036
rect 9468 894 9538 950
rect 9594 894 9680 950
rect 9736 894 9808 950
rect 9468 808 9808 894
rect 9468 752 9538 808
rect 9594 752 9680 808
rect 9736 752 9808 808
rect 9468 666 9808 752
rect 9468 610 9538 666
rect 9594 610 9680 666
rect 9736 610 9808 666
rect 9468 524 9808 610
rect 9468 468 9538 524
rect 9594 468 9680 524
rect 9736 468 9808 524
rect 9468 400 9808 468
rect 9868 12310 10208 12400
rect 9868 12254 9934 12310
rect 9990 12254 10076 12310
rect 10132 12254 10208 12310
rect 9868 12168 10208 12254
rect 9868 12112 9934 12168
rect 9990 12112 10076 12168
rect 10132 12112 10208 12168
rect 9868 12026 10208 12112
rect 9868 11970 9934 12026
rect 9990 11970 10076 12026
rect 10132 11970 10208 12026
rect 9868 11884 10208 11970
rect 9868 11828 9934 11884
rect 9990 11828 10076 11884
rect 10132 11828 10208 11884
rect 9868 11742 10208 11828
rect 9868 11686 9934 11742
rect 9990 11686 10076 11742
rect 10132 11686 10208 11742
rect 9868 11600 10208 11686
rect 9868 11544 9934 11600
rect 9990 11544 10076 11600
rect 10132 11544 10208 11600
rect 9868 11458 10208 11544
rect 9868 11402 9934 11458
rect 9990 11402 10076 11458
rect 10132 11402 10208 11458
rect 9868 11316 10208 11402
rect 9868 11260 9934 11316
rect 9990 11260 10076 11316
rect 10132 11260 10208 11316
rect 9868 11174 10208 11260
rect 9868 11118 9934 11174
rect 9990 11118 10076 11174
rect 10132 11118 10208 11174
rect 9868 11032 10208 11118
rect 9868 10976 9934 11032
rect 9990 10976 10076 11032
rect 10132 10976 10208 11032
rect 9868 10890 10208 10976
rect 9868 10834 9934 10890
rect 9990 10834 10076 10890
rect 10132 10834 10208 10890
rect 9868 10748 10208 10834
rect 9868 10692 9934 10748
rect 9990 10692 10076 10748
rect 10132 10692 10208 10748
rect 9868 10606 10208 10692
rect 9868 10550 9934 10606
rect 9990 10550 10076 10606
rect 10132 10550 10208 10606
rect 9868 10464 10208 10550
rect 9868 10408 9934 10464
rect 9990 10408 10076 10464
rect 10132 10408 10208 10464
rect 9868 10322 10208 10408
rect 9868 10266 9934 10322
rect 9990 10266 10076 10322
rect 10132 10266 10208 10322
rect 9868 10180 10208 10266
rect 9868 10124 9934 10180
rect 9990 10124 10076 10180
rect 10132 10124 10208 10180
rect 9868 10038 10208 10124
rect 9868 9982 9934 10038
rect 9990 9982 10076 10038
rect 10132 9982 10208 10038
rect 9868 9896 10208 9982
rect 9868 9840 9934 9896
rect 9990 9840 10076 9896
rect 10132 9840 10208 9896
rect 9868 9754 10208 9840
rect 9868 9698 9934 9754
rect 9990 9698 10076 9754
rect 10132 9698 10208 9754
rect 9868 9612 10208 9698
rect 9868 9556 9934 9612
rect 9990 9556 10076 9612
rect 10132 9556 10208 9612
rect 9868 9470 10208 9556
rect 9868 9414 9934 9470
rect 9990 9414 10076 9470
rect 10132 9414 10208 9470
rect 9868 9328 10208 9414
rect 9868 9272 9934 9328
rect 9990 9272 10076 9328
rect 10132 9272 10208 9328
rect 9868 9186 10208 9272
rect 9868 9130 9934 9186
rect 9990 9130 10076 9186
rect 10132 9130 10208 9186
rect 9868 9044 10208 9130
rect 9868 8988 9934 9044
rect 9990 8988 10076 9044
rect 10132 8988 10208 9044
rect 9868 8902 10208 8988
rect 9868 8846 9934 8902
rect 9990 8846 10076 8902
rect 10132 8846 10208 8902
rect 9868 8760 10208 8846
rect 9868 8704 9934 8760
rect 9990 8704 10076 8760
rect 10132 8704 10208 8760
rect 9868 8618 10208 8704
rect 9868 8562 9934 8618
rect 9990 8562 10076 8618
rect 10132 8562 10208 8618
rect 9868 8476 10208 8562
rect 9868 8420 9934 8476
rect 9990 8420 10076 8476
rect 10132 8420 10208 8476
rect 9868 8334 10208 8420
rect 9868 8278 9934 8334
rect 9990 8278 10076 8334
rect 10132 8278 10208 8334
rect 9868 8192 10208 8278
rect 9868 8136 9934 8192
rect 9990 8136 10076 8192
rect 10132 8136 10208 8192
rect 9868 8050 10208 8136
rect 9868 7994 9934 8050
rect 9990 7994 10076 8050
rect 10132 7994 10208 8050
rect 9868 7908 10208 7994
rect 9868 7852 9934 7908
rect 9990 7852 10076 7908
rect 10132 7852 10208 7908
rect 9868 7766 10208 7852
rect 9868 7710 9934 7766
rect 9990 7710 10076 7766
rect 10132 7710 10208 7766
rect 9868 7624 10208 7710
rect 9868 7568 9934 7624
rect 9990 7568 10076 7624
rect 10132 7568 10208 7624
rect 9868 7482 10208 7568
rect 9868 7426 9934 7482
rect 9990 7426 10076 7482
rect 10132 7426 10208 7482
rect 9868 7340 10208 7426
rect 9868 7284 9934 7340
rect 9990 7284 10076 7340
rect 10132 7284 10208 7340
rect 9868 7198 10208 7284
rect 9868 7142 9934 7198
rect 9990 7142 10076 7198
rect 10132 7142 10208 7198
rect 9868 7056 10208 7142
rect 9868 7000 9934 7056
rect 9990 7000 10076 7056
rect 10132 7000 10208 7056
rect 9868 6914 10208 7000
rect 9868 6858 9934 6914
rect 9990 6858 10076 6914
rect 10132 6858 10208 6914
rect 9868 6772 10208 6858
rect 9868 6716 9934 6772
rect 9990 6716 10076 6772
rect 10132 6716 10208 6772
rect 9868 6630 10208 6716
rect 9868 6574 9934 6630
rect 9990 6574 10076 6630
rect 10132 6574 10208 6630
rect 9868 6488 10208 6574
rect 9868 6432 9934 6488
rect 9990 6432 10076 6488
rect 10132 6432 10208 6488
rect 9868 6346 10208 6432
rect 9868 6290 9934 6346
rect 9990 6290 10076 6346
rect 10132 6290 10208 6346
rect 9868 6204 10208 6290
rect 9868 6148 9934 6204
rect 9990 6148 10076 6204
rect 10132 6148 10208 6204
rect 9868 6062 10208 6148
rect 9868 6006 9934 6062
rect 9990 6006 10076 6062
rect 10132 6006 10208 6062
rect 9868 5920 10208 6006
rect 9868 5864 9934 5920
rect 9990 5864 10076 5920
rect 10132 5864 10208 5920
rect 9868 5778 10208 5864
rect 9868 5722 9934 5778
rect 9990 5722 10076 5778
rect 10132 5722 10208 5778
rect 9868 5636 10208 5722
rect 9868 5580 9934 5636
rect 9990 5580 10076 5636
rect 10132 5580 10208 5636
rect 9868 5494 10208 5580
rect 9868 5438 9934 5494
rect 9990 5438 10076 5494
rect 10132 5438 10208 5494
rect 9868 5352 10208 5438
rect 9868 5296 9934 5352
rect 9990 5296 10076 5352
rect 10132 5296 10208 5352
rect 9868 5210 10208 5296
rect 9868 5154 9934 5210
rect 9990 5154 10076 5210
rect 10132 5154 10208 5210
rect 9868 5068 10208 5154
rect 9868 5012 9934 5068
rect 9990 5012 10076 5068
rect 10132 5012 10208 5068
rect 9868 4926 10208 5012
rect 9868 4870 9934 4926
rect 9990 4870 10076 4926
rect 10132 4870 10208 4926
rect 9868 4784 10208 4870
rect 9868 4728 9934 4784
rect 9990 4728 10076 4784
rect 10132 4728 10208 4784
rect 9868 4642 10208 4728
rect 9868 4586 9934 4642
rect 9990 4586 10076 4642
rect 10132 4586 10208 4642
rect 9868 4500 10208 4586
rect 9868 4444 9934 4500
rect 9990 4444 10076 4500
rect 10132 4444 10208 4500
rect 9868 4358 10208 4444
rect 9868 4302 9934 4358
rect 9990 4302 10076 4358
rect 10132 4302 10208 4358
rect 9868 4216 10208 4302
rect 9868 4160 9934 4216
rect 9990 4160 10076 4216
rect 10132 4160 10208 4216
rect 9868 4074 10208 4160
rect 9868 4018 9934 4074
rect 9990 4018 10076 4074
rect 10132 4018 10208 4074
rect 9868 3932 10208 4018
rect 9868 3876 9934 3932
rect 9990 3876 10076 3932
rect 10132 3876 10208 3932
rect 9868 3790 10208 3876
rect 9868 3734 9934 3790
rect 9990 3734 10076 3790
rect 10132 3734 10208 3790
rect 9868 3648 10208 3734
rect 9868 3592 9934 3648
rect 9990 3592 10076 3648
rect 10132 3592 10208 3648
rect 9868 3506 10208 3592
rect 9868 3450 9934 3506
rect 9990 3450 10076 3506
rect 10132 3450 10208 3506
rect 9868 3364 10208 3450
rect 9868 3308 9934 3364
rect 9990 3308 10076 3364
rect 10132 3308 10208 3364
rect 9868 3222 10208 3308
rect 9868 3166 9934 3222
rect 9990 3166 10076 3222
rect 10132 3166 10208 3222
rect 9868 3080 10208 3166
rect 9868 3024 9934 3080
rect 9990 3024 10076 3080
rect 10132 3024 10208 3080
rect 9868 2938 10208 3024
rect 9868 2882 9934 2938
rect 9990 2882 10076 2938
rect 10132 2882 10208 2938
rect 9868 2796 10208 2882
rect 9868 2740 9934 2796
rect 9990 2740 10076 2796
rect 10132 2740 10208 2796
rect 9868 2654 10208 2740
rect 9868 2598 9934 2654
rect 9990 2598 10076 2654
rect 10132 2598 10208 2654
rect 9868 2512 10208 2598
rect 9868 2456 9934 2512
rect 9990 2456 10076 2512
rect 10132 2456 10208 2512
rect 9868 2370 10208 2456
rect 9868 2314 9934 2370
rect 9990 2314 10076 2370
rect 10132 2314 10208 2370
rect 9868 2228 10208 2314
rect 9868 2172 9934 2228
rect 9990 2172 10076 2228
rect 10132 2172 10208 2228
rect 9868 2086 10208 2172
rect 9868 2030 9934 2086
rect 9990 2030 10076 2086
rect 10132 2030 10208 2086
rect 9868 1944 10208 2030
rect 9868 1888 9934 1944
rect 9990 1888 10076 1944
rect 10132 1888 10208 1944
rect 9868 1802 10208 1888
rect 9868 1746 9934 1802
rect 9990 1746 10076 1802
rect 10132 1746 10208 1802
rect 9868 1660 10208 1746
rect 9868 1604 9934 1660
rect 9990 1604 10076 1660
rect 10132 1604 10208 1660
rect 9868 1518 10208 1604
rect 9868 1462 9934 1518
rect 9990 1462 10076 1518
rect 10132 1462 10208 1518
rect 9868 1376 10208 1462
rect 9868 1320 9934 1376
rect 9990 1320 10076 1376
rect 10132 1320 10208 1376
rect 9868 1234 10208 1320
rect 9868 1178 9934 1234
rect 9990 1178 10076 1234
rect 10132 1178 10208 1234
rect 9868 1092 10208 1178
rect 9868 1036 9934 1092
rect 9990 1036 10076 1092
rect 10132 1036 10208 1092
rect 9868 950 10208 1036
rect 9868 894 9934 950
rect 9990 894 10076 950
rect 10132 894 10208 950
rect 9868 808 10208 894
rect 9868 752 9934 808
rect 9990 752 10076 808
rect 10132 752 10208 808
rect 9868 666 10208 752
rect 9868 610 9934 666
rect 9990 610 10076 666
rect 10132 610 10208 666
rect 9868 524 10208 610
rect 9868 468 9934 524
rect 9990 468 10076 524
rect 10132 468 10208 524
rect 9868 400 10208 468
rect 10268 12310 10608 12400
rect 10268 12254 10334 12310
rect 10390 12254 10476 12310
rect 10532 12254 10608 12310
rect 10268 12168 10608 12254
rect 10268 12112 10334 12168
rect 10390 12112 10476 12168
rect 10532 12112 10608 12168
rect 10268 12026 10608 12112
rect 10268 11970 10334 12026
rect 10390 11970 10476 12026
rect 10532 11970 10608 12026
rect 10268 11884 10608 11970
rect 10268 11828 10334 11884
rect 10390 11828 10476 11884
rect 10532 11828 10608 11884
rect 10268 11742 10608 11828
rect 10268 11686 10334 11742
rect 10390 11686 10476 11742
rect 10532 11686 10608 11742
rect 10268 11600 10608 11686
rect 10268 11544 10334 11600
rect 10390 11544 10476 11600
rect 10532 11544 10608 11600
rect 10268 11458 10608 11544
rect 10268 11402 10334 11458
rect 10390 11402 10476 11458
rect 10532 11402 10608 11458
rect 10268 11316 10608 11402
rect 10268 11260 10334 11316
rect 10390 11260 10476 11316
rect 10532 11260 10608 11316
rect 10268 11174 10608 11260
rect 10268 11118 10334 11174
rect 10390 11118 10476 11174
rect 10532 11118 10608 11174
rect 10268 11032 10608 11118
rect 10268 10976 10334 11032
rect 10390 10976 10476 11032
rect 10532 10976 10608 11032
rect 10268 10890 10608 10976
rect 10268 10834 10334 10890
rect 10390 10834 10476 10890
rect 10532 10834 10608 10890
rect 10268 10748 10608 10834
rect 10268 10692 10334 10748
rect 10390 10692 10476 10748
rect 10532 10692 10608 10748
rect 10268 10606 10608 10692
rect 10268 10550 10334 10606
rect 10390 10550 10476 10606
rect 10532 10550 10608 10606
rect 10268 10464 10608 10550
rect 10268 10408 10334 10464
rect 10390 10408 10476 10464
rect 10532 10408 10608 10464
rect 10268 10322 10608 10408
rect 10268 10266 10334 10322
rect 10390 10266 10476 10322
rect 10532 10266 10608 10322
rect 10268 10180 10608 10266
rect 10268 10124 10334 10180
rect 10390 10124 10476 10180
rect 10532 10124 10608 10180
rect 10268 10038 10608 10124
rect 10268 9982 10334 10038
rect 10390 9982 10476 10038
rect 10532 9982 10608 10038
rect 10268 9896 10608 9982
rect 10268 9840 10334 9896
rect 10390 9840 10476 9896
rect 10532 9840 10608 9896
rect 10268 9754 10608 9840
rect 10268 9698 10334 9754
rect 10390 9698 10476 9754
rect 10532 9698 10608 9754
rect 10268 9612 10608 9698
rect 10268 9556 10334 9612
rect 10390 9556 10476 9612
rect 10532 9556 10608 9612
rect 10268 9470 10608 9556
rect 10268 9414 10334 9470
rect 10390 9414 10476 9470
rect 10532 9414 10608 9470
rect 10268 9328 10608 9414
rect 10268 9272 10334 9328
rect 10390 9272 10476 9328
rect 10532 9272 10608 9328
rect 10268 9186 10608 9272
rect 10268 9130 10334 9186
rect 10390 9130 10476 9186
rect 10532 9130 10608 9186
rect 10268 9044 10608 9130
rect 10268 8988 10334 9044
rect 10390 8988 10476 9044
rect 10532 8988 10608 9044
rect 10268 8902 10608 8988
rect 10268 8846 10334 8902
rect 10390 8846 10476 8902
rect 10532 8846 10608 8902
rect 10268 8760 10608 8846
rect 10268 8704 10334 8760
rect 10390 8704 10476 8760
rect 10532 8704 10608 8760
rect 10268 8618 10608 8704
rect 10268 8562 10334 8618
rect 10390 8562 10476 8618
rect 10532 8562 10608 8618
rect 10268 8476 10608 8562
rect 10268 8420 10334 8476
rect 10390 8420 10476 8476
rect 10532 8420 10608 8476
rect 10268 8334 10608 8420
rect 10268 8278 10334 8334
rect 10390 8278 10476 8334
rect 10532 8278 10608 8334
rect 10268 8192 10608 8278
rect 10268 8136 10334 8192
rect 10390 8136 10476 8192
rect 10532 8136 10608 8192
rect 10268 8050 10608 8136
rect 10268 7994 10334 8050
rect 10390 7994 10476 8050
rect 10532 7994 10608 8050
rect 10268 7908 10608 7994
rect 10268 7852 10334 7908
rect 10390 7852 10476 7908
rect 10532 7852 10608 7908
rect 10268 7766 10608 7852
rect 10268 7710 10334 7766
rect 10390 7710 10476 7766
rect 10532 7710 10608 7766
rect 10268 7624 10608 7710
rect 10268 7568 10334 7624
rect 10390 7568 10476 7624
rect 10532 7568 10608 7624
rect 10268 7482 10608 7568
rect 10268 7426 10334 7482
rect 10390 7426 10476 7482
rect 10532 7426 10608 7482
rect 10268 7340 10608 7426
rect 10268 7284 10334 7340
rect 10390 7284 10476 7340
rect 10532 7284 10608 7340
rect 10268 7198 10608 7284
rect 10268 7142 10334 7198
rect 10390 7142 10476 7198
rect 10532 7142 10608 7198
rect 10268 7056 10608 7142
rect 10268 7000 10334 7056
rect 10390 7000 10476 7056
rect 10532 7000 10608 7056
rect 10268 6914 10608 7000
rect 10268 6858 10334 6914
rect 10390 6858 10476 6914
rect 10532 6858 10608 6914
rect 10268 6772 10608 6858
rect 10268 6716 10334 6772
rect 10390 6716 10476 6772
rect 10532 6716 10608 6772
rect 10268 6630 10608 6716
rect 10268 6574 10334 6630
rect 10390 6574 10476 6630
rect 10532 6574 10608 6630
rect 10268 6488 10608 6574
rect 10268 6432 10334 6488
rect 10390 6432 10476 6488
rect 10532 6432 10608 6488
rect 10268 6346 10608 6432
rect 10268 6290 10334 6346
rect 10390 6290 10476 6346
rect 10532 6290 10608 6346
rect 10268 6204 10608 6290
rect 10268 6148 10334 6204
rect 10390 6148 10476 6204
rect 10532 6148 10608 6204
rect 10268 6062 10608 6148
rect 10268 6006 10334 6062
rect 10390 6006 10476 6062
rect 10532 6006 10608 6062
rect 10268 5920 10608 6006
rect 10268 5864 10334 5920
rect 10390 5864 10476 5920
rect 10532 5864 10608 5920
rect 10268 5778 10608 5864
rect 10268 5722 10334 5778
rect 10390 5722 10476 5778
rect 10532 5722 10608 5778
rect 10268 5636 10608 5722
rect 10268 5580 10334 5636
rect 10390 5580 10476 5636
rect 10532 5580 10608 5636
rect 10268 5494 10608 5580
rect 10268 5438 10334 5494
rect 10390 5438 10476 5494
rect 10532 5438 10608 5494
rect 10268 5352 10608 5438
rect 10268 5296 10334 5352
rect 10390 5296 10476 5352
rect 10532 5296 10608 5352
rect 10268 5210 10608 5296
rect 10268 5154 10334 5210
rect 10390 5154 10476 5210
rect 10532 5154 10608 5210
rect 10268 5068 10608 5154
rect 10268 5012 10334 5068
rect 10390 5012 10476 5068
rect 10532 5012 10608 5068
rect 10268 4926 10608 5012
rect 10268 4870 10334 4926
rect 10390 4870 10476 4926
rect 10532 4870 10608 4926
rect 10268 4784 10608 4870
rect 10268 4728 10334 4784
rect 10390 4728 10476 4784
rect 10532 4728 10608 4784
rect 10268 4642 10608 4728
rect 10268 4586 10334 4642
rect 10390 4586 10476 4642
rect 10532 4586 10608 4642
rect 10268 4500 10608 4586
rect 10268 4444 10334 4500
rect 10390 4444 10476 4500
rect 10532 4444 10608 4500
rect 10268 4358 10608 4444
rect 10268 4302 10334 4358
rect 10390 4302 10476 4358
rect 10532 4302 10608 4358
rect 10268 4216 10608 4302
rect 10268 4160 10334 4216
rect 10390 4160 10476 4216
rect 10532 4160 10608 4216
rect 10268 4074 10608 4160
rect 10268 4018 10334 4074
rect 10390 4018 10476 4074
rect 10532 4018 10608 4074
rect 10268 3932 10608 4018
rect 10268 3876 10334 3932
rect 10390 3876 10476 3932
rect 10532 3876 10608 3932
rect 10268 3790 10608 3876
rect 10268 3734 10334 3790
rect 10390 3734 10476 3790
rect 10532 3734 10608 3790
rect 10268 3648 10608 3734
rect 10268 3592 10334 3648
rect 10390 3592 10476 3648
rect 10532 3592 10608 3648
rect 10268 3506 10608 3592
rect 10268 3450 10334 3506
rect 10390 3450 10476 3506
rect 10532 3450 10608 3506
rect 10268 3364 10608 3450
rect 10268 3308 10334 3364
rect 10390 3308 10476 3364
rect 10532 3308 10608 3364
rect 10268 3222 10608 3308
rect 10268 3166 10334 3222
rect 10390 3166 10476 3222
rect 10532 3166 10608 3222
rect 10268 3080 10608 3166
rect 10268 3024 10334 3080
rect 10390 3024 10476 3080
rect 10532 3024 10608 3080
rect 10268 2938 10608 3024
rect 10268 2882 10334 2938
rect 10390 2882 10476 2938
rect 10532 2882 10608 2938
rect 10268 2796 10608 2882
rect 10268 2740 10334 2796
rect 10390 2740 10476 2796
rect 10532 2740 10608 2796
rect 10268 2654 10608 2740
rect 10268 2598 10334 2654
rect 10390 2598 10476 2654
rect 10532 2598 10608 2654
rect 10268 2512 10608 2598
rect 10268 2456 10334 2512
rect 10390 2456 10476 2512
rect 10532 2456 10608 2512
rect 10268 2370 10608 2456
rect 10268 2314 10334 2370
rect 10390 2314 10476 2370
rect 10532 2314 10608 2370
rect 10268 2228 10608 2314
rect 10268 2172 10334 2228
rect 10390 2172 10476 2228
rect 10532 2172 10608 2228
rect 10268 2086 10608 2172
rect 10268 2030 10334 2086
rect 10390 2030 10476 2086
rect 10532 2030 10608 2086
rect 10268 1944 10608 2030
rect 10268 1888 10334 1944
rect 10390 1888 10476 1944
rect 10532 1888 10608 1944
rect 10268 1802 10608 1888
rect 10268 1746 10334 1802
rect 10390 1746 10476 1802
rect 10532 1746 10608 1802
rect 10268 1660 10608 1746
rect 10268 1604 10334 1660
rect 10390 1604 10476 1660
rect 10532 1604 10608 1660
rect 10268 1518 10608 1604
rect 10268 1462 10334 1518
rect 10390 1462 10476 1518
rect 10532 1462 10608 1518
rect 10268 1376 10608 1462
rect 10268 1320 10334 1376
rect 10390 1320 10476 1376
rect 10532 1320 10608 1376
rect 10268 1234 10608 1320
rect 10268 1178 10334 1234
rect 10390 1178 10476 1234
rect 10532 1178 10608 1234
rect 10268 1092 10608 1178
rect 10268 1036 10334 1092
rect 10390 1036 10476 1092
rect 10532 1036 10608 1092
rect 10268 950 10608 1036
rect 10268 894 10334 950
rect 10390 894 10476 950
rect 10532 894 10608 950
rect 10268 808 10608 894
rect 10268 752 10334 808
rect 10390 752 10476 808
rect 10532 752 10608 808
rect 10268 666 10608 752
rect 10268 610 10334 666
rect 10390 610 10476 666
rect 10532 610 10608 666
rect 10268 524 10608 610
rect 10268 468 10334 524
rect 10390 468 10476 524
rect 10532 468 10608 524
rect 10268 400 10608 468
rect 10668 12310 11008 12400
rect 10668 12254 10731 12310
rect 10787 12254 10873 12310
rect 10929 12254 11008 12310
rect 10668 12168 11008 12254
rect 10668 12112 10731 12168
rect 10787 12112 10873 12168
rect 10929 12112 11008 12168
rect 10668 12026 11008 12112
rect 10668 11970 10731 12026
rect 10787 11970 10873 12026
rect 10929 11970 11008 12026
rect 10668 11884 11008 11970
rect 10668 11828 10731 11884
rect 10787 11828 10873 11884
rect 10929 11828 11008 11884
rect 10668 11742 11008 11828
rect 10668 11686 10731 11742
rect 10787 11686 10873 11742
rect 10929 11686 11008 11742
rect 10668 11600 11008 11686
rect 10668 11544 10731 11600
rect 10787 11544 10873 11600
rect 10929 11544 11008 11600
rect 10668 11458 11008 11544
rect 10668 11402 10731 11458
rect 10787 11402 10873 11458
rect 10929 11402 11008 11458
rect 10668 11316 11008 11402
rect 10668 11260 10731 11316
rect 10787 11260 10873 11316
rect 10929 11260 11008 11316
rect 10668 11174 11008 11260
rect 10668 11118 10731 11174
rect 10787 11118 10873 11174
rect 10929 11118 11008 11174
rect 10668 11032 11008 11118
rect 10668 10976 10731 11032
rect 10787 10976 10873 11032
rect 10929 10976 11008 11032
rect 10668 10890 11008 10976
rect 10668 10834 10731 10890
rect 10787 10834 10873 10890
rect 10929 10834 11008 10890
rect 10668 10748 11008 10834
rect 10668 10692 10731 10748
rect 10787 10692 10873 10748
rect 10929 10692 11008 10748
rect 10668 10606 11008 10692
rect 10668 10550 10731 10606
rect 10787 10550 10873 10606
rect 10929 10550 11008 10606
rect 10668 10464 11008 10550
rect 10668 10408 10731 10464
rect 10787 10408 10873 10464
rect 10929 10408 11008 10464
rect 10668 10322 11008 10408
rect 10668 10266 10731 10322
rect 10787 10266 10873 10322
rect 10929 10266 11008 10322
rect 10668 10180 11008 10266
rect 10668 10124 10731 10180
rect 10787 10124 10873 10180
rect 10929 10124 11008 10180
rect 10668 10038 11008 10124
rect 10668 9982 10731 10038
rect 10787 9982 10873 10038
rect 10929 9982 11008 10038
rect 10668 9896 11008 9982
rect 10668 9840 10731 9896
rect 10787 9840 10873 9896
rect 10929 9840 11008 9896
rect 10668 9754 11008 9840
rect 10668 9698 10731 9754
rect 10787 9698 10873 9754
rect 10929 9698 11008 9754
rect 10668 9612 11008 9698
rect 10668 9556 10731 9612
rect 10787 9556 10873 9612
rect 10929 9556 11008 9612
rect 10668 9470 11008 9556
rect 10668 9414 10731 9470
rect 10787 9414 10873 9470
rect 10929 9414 11008 9470
rect 10668 9328 11008 9414
rect 10668 9272 10731 9328
rect 10787 9272 10873 9328
rect 10929 9272 11008 9328
rect 10668 9186 11008 9272
rect 10668 9130 10731 9186
rect 10787 9130 10873 9186
rect 10929 9130 11008 9186
rect 10668 9044 11008 9130
rect 10668 8988 10731 9044
rect 10787 8988 10873 9044
rect 10929 8988 11008 9044
rect 10668 8902 11008 8988
rect 10668 8846 10731 8902
rect 10787 8846 10873 8902
rect 10929 8846 11008 8902
rect 10668 8760 11008 8846
rect 10668 8704 10731 8760
rect 10787 8704 10873 8760
rect 10929 8704 11008 8760
rect 10668 8618 11008 8704
rect 10668 8562 10731 8618
rect 10787 8562 10873 8618
rect 10929 8562 11008 8618
rect 10668 8476 11008 8562
rect 10668 8420 10731 8476
rect 10787 8420 10873 8476
rect 10929 8420 11008 8476
rect 10668 8334 11008 8420
rect 10668 8278 10731 8334
rect 10787 8278 10873 8334
rect 10929 8278 11008 8334
rect 10668 8192 11008 8278
rect 10668 8136 10731 8192
rect 10787 8136 10873 8192
rect 10929 8136 11008 8192
rect 10668 8050 11008 8136
rect 10668 7994 10731 8050
rect 10787 7994 10873 8050
rect 10929 7994 11008 8050
rect 10668 7908 11008 7994
rect 10668 7852 10731 7908
rect 10787 7852 10873 7908
rect 10929 7852 11008 7908
rect 10668 7766 11008 7852
rect 10668 7710 10731 7766
rect 10787 7710 10873 7766
rect 10929 7710 11008 7766
rect 10668 7624 11008 7710
rect 10668 7568 10731 7624
rect 10787 7568 10873 7624
rect 10929 7568 11008 7624
rect 10668 7482 11008 7568
rect 10668 7426 10731 7482
rect 10787 7426 10873 7482
rect 10929 7426 11008 7482
rect 10668 7340 11008 7426
rect 10668 7284 10731 7340
rect 10787 7284 10873 7340
rect 10929 7284 11008 7340
rect 10668 7198 11008 7284
rect 10668 7142 10731 7198
rect 10787 7142 10873 7198
rect 10929 7142 11008 7198
rect 10668 7056 11008 7142
rect 10668 7000 10731 7056
rect 10787 7000 10873 7056
rect 10929 7000 11008 7056
rect 10668 6914 11008 7000
rect 10668 6858 10731 6914
rect 10787 6858 10873 6914
rect 10929 6858 11008 6914
rect 10668 6772 11008 6858
rect 10668 6716 10731 6772
rect 10787 6716 10873 6772
rect 10929 6716 11008 6772
rect 10668 6630 11008 6716
rect 10668 6574 10731 6630
rect 10787 6574 10873 6630
rect 10929 6574 11008 6630
rect 10668 6488 11008 6574
rect 10668 6432 10731 6488
rect 10787 6432 10873 6488
rect 10929 6432 11008 6488
rect 10668 6346 11008 6432
rect 10668 6290 10731 6346
rect 10787 6290 10873 6346
rect 10929 6290 11008 6346
rect 10668 6204 11008 6290
rect 10668 6148 10731 6204
rect 10787 6148 10873 6204
rect 10929 6148 11008 6204
rect 10668 6062 11008 6148
rect 10668 6006 10731 6062
rect 10787 6006 10873 6062
rect 10929 6006 11008 6062
rect 10668 5920 11008 6006
rect 10668 5864 10731 5920
rect 10787 5864 10873 5920
rect 10929 5864 11008 5920
rect 10668 5778 11008 5864
rect 10668 5722 10731 5778
rect 10787 5722 10873 5778
rect 10929 5722 11008 5778
rect 10668 5636 11008 5722
rect 10668 5580 10731 5636
rect 10787 5580 10873 5636
rect 10929 5580 11008 5636
rect 10668 5494 11008 5580
rect 10668 5438 10731 5494
rect 10787 5438 10873 5494
rect 10929 5438 11008 5494
rect 10668 5352 11008 5438
rect 10668 5296 10731 5352
rect 10787 5296 10873 5352
rect 10929 5296 11008 5352
rect 10668 5210 11008 5296
rect 10668 5154 10731 5210
rect 10787 5154 10873 5210
rect 10929 5154 11008 5210
rect 10668 5068 11008 5154
rect 10668 5012 10731 5068
rect 10787 5012 10873 5068
rect 10929 5012 11008 5068
rect 10668 4926 11008 5012
rect 10668 4870 10731 4926
rect 10787 4870 10873 4926
rect 10929 4870 11008 4926
rect 10668 4784 11008 4870
rect 10668 4728 10731 4784
rect 10787 4728 10873 4784
rect 10929 4728 11008 4784
rect 10668 4642 11008 4728
rect 10668 4586 10731 4642
rect 10787 4586 10873 4642
rect 10929 4586 11008 4642
rect 10668 4500 11008 4586
rect 10668 4444 10731 4500
rect 10787 4444 10873 4500
rect 10929 4444 11008 4500
rect 10668 4358 11008 4444
rect 10668 4302 10731 4358
rect 10787 4302 10873 4358
rect 10929 4302 11008 4358
rect 10668 4216 11008 4302
rect 10668 4160 10731 4216
rect 10787 4160 10873 4216
rect 10929 4160 11008 4216
rect 10668 4074 11008 4160
rect 10668 4018 10731 4074
rect 10787 4018 10873 4074
rect 10929 4018 11008 4074
rect 10668 3932 11008 4018
rect 10668 3876 10731 3932
rect 10787 3876 10873 3932
rect 10929 3876 11008 3932
rect 10668 3790 11008 3876
rect 10668 3734 10731 3790
rect 10787 3734 10873 3790
rect 10929 3734 11008 3790
rect 10668 3648 11008 3734
rect 10668 3592 10731 3648
rect 10787 3592 10873 3648
rect 10929 3592 11008 3648
rect 10668 3506 11008 3592
rect 10668 3450 10731 3506
rect 10787 3450 10873 3506
rect 10929 3450 11008 3506
rect 10668 3364 11008 3450
rect 10668 3308 10731 3364
rect 10787 3308 10873 3364
rect 10929 3308 11008 3364
rect 10668 3222 11008 3308
rect 10668 3166 10731 3222
rect 10787 3166 10873 3222
rect 10929 3166 11008 3222
rect 10668 3080 11008 3166
rect 10668 3024 10731 3080
rect 10787 3024 10873 3080
rect 10929 3024 11008 3080
rect 10668 2938 11008 3024
rect 10668 2882 10731 2938
rect 10787 2882 10873 2938
rect 10929 2882 11008 2938
rect 10668 2796 11008 2882
rect 10668 2740 10731 2796
rect 10787 2740 10873 2796
rect 10929 2740 11008 2796
rect 10668 2654 11008 2740
rect 10668 2598 10731 2654
rect 10787 2598 10873 2654
rect 10929 2598 11008 2654
rect 10668 2512 11008 2598
rect 10668 2456 10731 2512
rect 10787 2456 10873 2512
rect 10929 2456 11008 2512
rect 10668 2370 11008 2456
rect 10668 2314 10731 2370
rect 10787 2314 10873 2370
rect 10929 2314 11008 2370
rect 10668 2228 11008 2314
rect 10668 2172 10731 2228
rect 10787 2172 10873 2228
rect 10929 2172 11008 2228
rect 10668 2086 11008 2172
rect 10668 2030 10731 2086
rect 10787 2030 10873 2086
rect 10929 2030 11008 2086
rect 10668 1944 11008 2030
rect 10668 1888 10731 1944
rect 10787 1888 10873 1944
rect 10929 1888 11008 1944
rect 10668 1802 11008 1888
rect 10668 1746 10731 1802
rect 10787 1746 10873 1802
rect 10929 1746 11008 1802
rect 10668 1660 11008 1746
rect 10668 1604 10731 1660
rect 10787 1604 10873 1660
rect 10929 1604 11008 1660
rect 10668 1518 11008 1604
rect 10668 1462 10731 1518
rect 10787 1462 10873 1518
rect 10929 1462 11008 1518
rect 10668 1376 11008 1462
rect 10668 1320 10731 1376
rect 10787 1320 10873 1376
rect 10929 1320 11008 1376
rect 10668 1234 11008 1320
rect 10668 1178 10731 1234
rect 10787 1178 10873 1234
rect 10929 1178 11008 1234
rect 10668 1092 11008 1178
rect 10668 1036 10731 1092
rect 10787 1036 10873 1092
rect 10929 1036 11008 1092
rect 10668 950 11008 1036
rect 10668 894 10731 950
rect 10787 894 10873 950
rect 10929 894 11008 950
rect 10668 808 11008 894
rect 10668 752 10731 808
rect 10787 752 10873 808
rect 10929 752 11008 808
rect 10668 666 11008 752
rect 10668 610 10731 666
rect 10787 610 10873 666
rect 10929 610 11008 666
rect 10668 524 11008 610
rect 10668 468 10731 524
rect 10787 468 10873 524
rect 10929 468 11008 524
rect 10668 400 11008 468
rect 11068 12310 11408 12400
rect 11068 12254 11136 12310
rect 11192 12254 11278 12310
rect 11334 12254 11408 12310
rect 11068 12168 11408 12254
rect 11068 12112 11136 12168
rect 11192 12112 11278 12168
rect 11334 12112 11408 12168
rect 11068 12026 11408 12112
rect 11068 11970 11136 12026
rect 11192 11970 11278 12026
rect 11334 11970 11408 12026
rect 11068 11884 11408 11970
rect 11068 11828 11136 11884
rect 11192 11828 11278 11884
rect 11334 11828 11408 11884
rect 11068 11742 11408 11828
rect 11068 11686 11136 11742
rect 11192 11686 11278 11742
rect 11334 11686 11408 11742
rect 11068 11600 11408 11686
rect 11068 11544 11136 11600
rect 11192 11544 11278 11600
rect 11334 11544 11408 11600
rect 11068 11458 11408 11544
rect 11068 11402 11136 11458
rect 11192 11402 11278 11458
rect 11334 11402 11408 11458
rect 11068 11316 11408 11402
rect 11068 11260 11136 11316
rect 11192 11260 11278 11316
rect 11334 11260 11408 11316
rect 11068 11174 11408 11260
rect 11068 11118 11136 11174
rect 11192 11118 11278 11174
rect 11334 11118 11408 11174
rect 11068 11032 11408 11118
rect 11068 10976 11136 11032
rect 11192 10976 11278 11032
rect 11334 10976 11408 11032
rect 11068 10890 11408 10976
rect 11068 10834 11136 10890
rect 11192 10834 11278 10890
rect 11334 10834 11408 10890
rect 11068 10748 11408 10834
rect 11068 10692 11136 10748
rect 11192 10692 11278 10748
rect 11334 10692 11408 10748
rect 11068 10606 11408 10692
rect 11068 10550 11136 10606
rect 11192 10550 11278 10606
rect 11334 10550 11408 10606
rect 11068 10464 11408 10550
rect 11068 10408 11136 10464
rect 11192 10408 11278 10464
rect 11334 10408 11408 10464
rect 11068 10322 11408 10408
rect 11068 10266 11136 10322
rect 11192 10266 11278 10322
rect 11334 10266 11408 10322
rect 11068 10180 11408 10266
rect 11068 10124 11136 10180
rect 11192 10124 11278 10180
rect 11334 10124 11408 10180
rect 11068 10038 11408 10124
rect 11068 9982 11136 10038
rect 11192 9982 11278 10038
rect 11334 9982 11408 10038
rect 11068 9896 11408 9982
rect 11068 9840 11136 9896
rect 11192 9840 11278 9896
rect 11334 9840 11408 9896
rect 11068 9754 11408 9840
rect 11068 9698 11136 9754
rect 11192 9698 11278 9754
rect 11334 9698 11408 9754
rect 11068 9612 11408 9698
rect 11068 9556 11136 9612
rect 11192 9556 11278 9612
rect 11334 9556 11408 9612
rect 11068 9470 11408 9556
rect 11068 9414 11136 9470
rect 11192 9414 11278 9470
rect 11334 9414 11408 9470
rect 11068 9328 11408 9414
rect 11068 9272 11136 9328
rect 11192 9272 11278 9328
rect 11334 9272 11408 9328
rect 11068 9186 11408 9272
rect 11068 9130 11136 9186
rect 11192 9130 11278 9186
rect 11334 9130 11408 9186
rect 11068 9044 11408 9130
rect 11068 8988 11136 9044
rect 11192 8988 11278 9044
rect 11334 8988 11408 9044
rect 11068 8902 11408 8988
rect 11068 8846 11136 8902
rect 11192 8846 11278 8902
rect 11334 8846 11408 8902
rect 11068 8760 11408 8846
rect 11068 8704 11136 8760
rect 11192 8704 11278 8760
rect 11334 8704 11408 8760
rect 11068 8618 11408 8704
rect 11068 8562 11136 8618
rect 11192 8562 11278 8618
rect 11334 8562 11408 8618
rect 11068 8476 11408 8562
rect 11068 8420 11136 8476
rect 11192 8420 11278 8476
rect 11334 8420 11408 8476
rect 11068 8334 11408 8420
rect 11068 8278 11136 8334
rect 11192 8278 11278 8334
rect 11334 8278 11408 8334
rect 11068 8192 11408 8278
rect 11068 8136 11136 8192
rect 11192 8136 11278 8192
rect 11334 8136 11408 8192
rect 11068 8050 11408 8136
rect 11068 7994 11136 8050
rect 11192 7994 11278 8050
rect 11334 7994 11408 8050
rect 11068 7908 11408 7994
rect 11068 7852 11136 7908
rect 11192 7852 11278 7908
rect 11334 7852 11408 7908
rect 11068 7766 11408 7852
rect 11068 7710 11136 7766
rect 11192 7710 11278 7766
rect 11334 7710 11408 7766
rect 11068 7624 11408 7710
rect 11068 7568 11136 7624
rect 11192 7568 11278 7624
rect 11334 7568 11408 7624
rect 11068 7482 11408 7568
rect 11068 7426 11136 7482
rect 11192 7426 11278 7482
rect 11334 7426 11408 7482
rect 11068 7340 11408 7426
rect 11068 7284 11136 7340
rect 11192 7284 11278 7340
rect 11334 7284 11408 7340
rect 11068 7198 11408 7284
rect 11068 7142 11136 7198
rect 11192 7142 11278 7198
rect 11334 7142 11408 7198
rect 11068 7056 11408 7142
rect 11068 7000 11136 7056
rect 11192 7000 11278 7056
rect 11334 7000 11408 7056
rect 11068 6914 11408 7000
rect 11068 6858 11136 6914
rect 11192 6858 11278 6914
rect 11334 6858 11408 6914
rect 11068 6772 11408 6858
rect 11068 6716 11136 6772
rect 11192 6716 11278 6772
rect 11334 6716 11408 6772
rect 11068 6630 11408 6716
rect 11068 6574 11136 6630
rect 11192 6574 11278 6630
rect 11334 6574 11408 6630
rect 11068 6488 11408 6574
rect 11068 6432 11136 6488
rect 11192 6432 11278 6488
rect 11334 6432 11408 6488
rect 11068 6346 11408 6432
rect 11068 6290 11136 6346
rect 11192 6290 11278 6346
rect 11334 6290 11408 6346
rect 11068 6204 11408 6290
rect 11068 6148 11136 6204
rect 11192 6148 11278 6204
rect 11334 6148 11408 6204
rect 11068 6062 11408 6148
rect 11068 6006 11136 6062
rect 11192 6006 11278 6062
rect 11334 6006 11408 6062
rect 11068 5920 11408 6006
rect 11068 5864 11136 5920
rect 11192 5864 11278 5920
rect 11334 5864 11408 5920
rect 11068 5778 11408 5864
rect 11068 5722 11136 5778
rect 11192 5722 11278 5778
rect 11334 5722 11408 5778
rect 11068 5636 11408 5722
rect 11068 5580 11136 5636
rect 11192 5580 11278 5636
rect 11334 5580 11408 5636
rect 11068 5494 11408 5580
rect 11068 5438 11136 5494
rect 11192 5438 11278 5494
rect 11334 5438 11408 5494
rect 11068 5352 11408 5438
rect 11068 5296 11136 5352
rect 11192 5296 11278 5352
rect 11334 5296 11408 5352
rect 11068 5210 11408 5296
rect 11068 5154 11136 5210
rect 11192 5154 11278 5210
rect 11334 5154 11408 5210
rect 11068 5068 11408 5154
rect 11068 5012 11136 5068
rect 11192 5012 11278 5068
rect 11334 5012 11408 5068
rect 11068 4926 11408 5012
rect 11068 4870 11136 4926
rect 11192 4870 11278 4926
rect 11334 4870 11408 4926
rect 11068 4784 11408 4870
rect 11068 4728 11136 4784
rect 11192 4728 11278 4784
rect 11334 4728 11408 4784
rect 11068 4642 11408 4728
rect 11068 4586 11136 4642
rect 11192 4586 11278 4642
rect 11334 4586 11408 4642
rect 11068 4500 11408 4586
rect 11068 4444 11136 4500
rect 11192 4444 11278 4500
rect 11334 4444 11408 4500
rect 11068 4358 11408 4444
rect 11068 4302 11136 4358
rect 11192 4302 11278 4358
rect 11334 4302 11408 4358
rect 11068 4216 11408 4302
rect 11068 4160 11136 4216
rect 11192 4160 11278 4216
rect 11334 4160 11408 4216
rect 11068 4074 11408 4160
rect 11068 4018 11136 4074
rect 11192 4018 11278 4074
rect 11334 4018 11408 4074
rect 11068 3932 11408 4018
rect 11068 3876 11136 3932
rect 11192 3876 11278 3932
rect 11334 3876 11408 3932
rect 11068 3790 11408 3876
rect 11068 3734 11136 3790
rect 11192 3734 11278 3790
rect 11334 3734 11408 3790
rect 11068 3648 11408 3734
rect 11068 3592 11136 3648
rect 11192 3592 11278 3648
rect 11334 3592 11408 3648
rect 11068 3506 11408 3592
rect 11068 3450 11136 3506
rect 11192 3450 11278 3506
rect 11334 3450 11408 3506
rect 11068 3364 11408 3450
rect 11068 3308 11136 3364
rect 11192 3308 11278 3364
rect 11334 3308 11408 3364
rect 11068 3222 11408 3308
rect 11068 3166 11136 3222
rect 11192 3166 11278 3222
rect 11334 3166 11408 3222
rect 11068 3080 11408 3166
rect 11068 3024 11136 3080
rect 11192 3024 11278 3080
rect 11334 3024 11408 3080
rect 11068 2938 11408 3024
rect 11068 2882 11136 2938
rect 11192 2882 11278 2938
rect 11334 2882 11408 2938
rect 11068 2796 11408 2882
rect 11068 2740 11136 2796
rect 11192 2740 11278 2796
rect 11334 2740 11408 2796
rect 11068 2654 11408 2740
rect 11068 2598 11136 2654
rect 11192 2598 11278 2654
rect 11334 2598 11408 2654
rect 11068 2512 11408 2598
rect 11068 2456 11136 2512
rect 11192 2456 11278 2512
rect 11334 2456 11408 2512
rect 11068 2370 11408 2456
rect 11068 2314 11136 2370
rect 11192 2314 11278 2370
rect 11334 2314 11408 2370
rect 11068 2228 11408 2314
rect 11068 2172 11136 2228
rect 11192 2172 11278 2228
rect 11334 2172 11408 2228
rect 11068 2086 11408 2172
rect 11068 2030 11136 2086
rect 11192 2030 11278 2086
rect 11334 2030 11408 2086
rect 11068 1944 11408 2030
rect 11068 1888 11136 1944
rect 11192 1888 11278 1944
rect 11334 1888 11408 1944
rect 11068 1802 11408 1888
rect 11068 1746 11136 1802
rect 11192 1746 11278 1802
rect 11334 1746 11408 1802
rect 11068 1660 11408 1746
rect 11068 1604 11136 1660
rect 11192 1604 11278 1660
rect 11334 1604 11408 1660
rect 11068 1518 11408 1604
rect 11068 1462 11136 1518
rect 11192 1462 11278 1518
rect 11334 1462 11408 1518
rect 11068 1376 11408 1462
rect 11068 1320 11136 1376
rect 11192 1320 11278 1376
rect 11334 1320 11408 1376
rect 11068 1234 11408 1320
rect 11068 1178 11136 1234
rect 11192 1178 11278 1234
rect 11334 1178 11408 1234
rect 11068 1092 11408 1178
rect 11068 1036 11136 1092
rect 11192 1036 11278 1092
rect 11334 1036 11408 1092
rect 11068 950 11408 1036
rect 11068 894 11136 950
rect 11192 894 11278 950
rect 11334 894 11408 950
rect 11068 808 11408 894
rect 11068 752 11136 808
rect 11192 752 11278 808
rect 11334 752 11408 808
rect 11068 666 11408 752
rect 11068 610 11136 666
rect 11192 610 11278 666
rect 11334 610 11408 666
rect 11068 524 11408 610
rect 11068 468 11136 524
rect 11192 468 11278 524
rect 11334 468 11408 524
rect 11068 400 11408 468
rect 11468 12310 11808 12400
rect 11468 12254 11536 12310
rect 11592 12254 11678 12310
rect 11734 12254 11808 12310
rect 11468 12168 11808 12254
rect 11468 12112 11536 12168
rect 11592 12112 11678 12168
rect 11734 12112 11808 12168
rect 11468 12026 11808 12112
rect 11468 11970 11536 12026
rect 11592 11970 11678 12026
rect 11734 11970 11808 12026
rect 11468 11884 11808 11970
rect 11468 11828 11536 11884
rect 11592 11828 11678 11884
rect 11734 11828 11808 11884
rect 11468 11742 11808 11828
rect 11468 11686 11536 11742
rect 11592 11686 11678 11742
rect 11734 11686 11808 11742
rect 11468 11600 11808 11686
rect 11468 11544 11536 11600
rect 11592 11544 11678 11600
rect 11734 11544 11808 11600
rect 11468 11458 11808 11544
rect 11468 11402 11536 11458
rect 11592 11402 11678 11458
rect 11734 11402 11808 11458
rect 11468 11316 11808 11402
rect 11468 11260 11536 11316
rect 11592 11260 11678 11316
rect 11734 11260 11808 11316
rect 11468 11174 11808 11260
rect 11468 11118 11536 11174
rect 11592 11118 11678 11174
rect 11734 11118 11808 11174
rect 11468 11032 11808 11118
rect 11468 10976 11536 11032
rect 11592 10976 11678 11032
rect 11734 10976 11808 11032
rect 11468 10890 11808 10976
rect 11468 10834 11536 10890
rect 11592 10834 11678 10890
rect 11734 10834 11808 10890
rect 11468 10748 11808 10834
rect 11468 10692 11536 10748
rect 11592 10692 11678 10748
rect 11734 10692 11808 10748
rect 11468 10606 11808 10692
rect 11468 10550 11536 10606
rect 11592 10550 11678 10606
rect 11734 10550 11808 10606
rect 11468 10464 11808 10550
rect 11468 10408 11536 10464
rect 11592 10408 11678 10464
rect 11734 10408 11808 10464
rect 11468 10322 11808 10408
rect 11468 10266 11536 10322
rect 11592 10266 11678 10322
rect 11734 10266 11808 10322
rect 11468 10180 11808 10266
rect 11468 10124 11536 10180
rect 11592 10124 11678 10180
rect 11734 10124 11808 10180
rect 11468 10038 11808 10124
rect 11468 9982 11536 10038
rect 11592 9982 11678 10038
rect 11734 9982 11808 10038
rect 11468 9896 11808 9982
rect 11468 9840 11536 9896
rect 11592 9840 11678 9896
rect 11734 9840 11808 9896
rect 11468 9754 11808 9840
rect 11468 9698 11536 9754
rect 11592 9698 11678 9754
rect 11734 9698 11808 9754
rect 11468 9612 11808 9698
rect 11468 9556 11536 9612
rect 11592 9556 11678 9612
rect 11734 9556 11808 9612
rect 11468 9470 11808 9556
rect 11468 9414 11536 9470
rect 11592 9414 11678 9470
rect 11734 9414 11808 9470
rect 11468 9328 11808 9414
rect 11468 9272 11536 9328
rect 11592 9272 11678 9328
rect 11734 9272 11808 9328
rect 11468 9186 11808 9272
rect 11468 9130 11536 9186
rect 11592 9130 11678 9186
rect 11734 9130 11808 9186
rect 11468 9044 11808 9130
rect 11468 8988 11536 9044
rect 11592 8988 11678 9044
rect 11734 8988 11808 9044
rect 11468 8902 11808 8988
rect 11468 8846 11536 8902
rect 11592 8846 11678 8902
rect 11734 8846 11808 8902
rect 11468 8760 11808 8846
rect 11468 8704 11536 8760
rect 11592 8704 11678 8760
rect 11734 8704 11808 8760
rect 11468 8618 11808 8704
rect 11468 8562 11536 8618
rect 11592 8562 11678 8618
rect 11734 8562 11808 8618
rect 11468 8476 11808 8562
rect 11468 8420 11536 8476
rect 11592 8420 11678 8476
rect 11734 8420 11808 8476
rect 11468 8334 11808 8420
rect 11468 8278 11536 8334
rect 11592 8278 11678 8334
rect 11734 8278 11808 8334
rect 11468 8192 11808 8278
rect 11468 8136 11536 8192
rect 11592 8136 11678 8192
rect 11734 8136 11808 8192
rect 11468 8050 11808 8136
rect 11468 7994 11536 8050
rect 11592 7994 11678 8050
rect 11734 7994 11808 8050
rect 11468 7908 11808 7994
rect 11468 7852 11536 7908
rect 11592 7852 11678 7908
rect 11734 7852 11808 7908
rect 11468 7766 11808 7852
rect 11468 7710 11536 7766
rect 11592 7710 11678 7766
rect 11734 7710 11808 7766
rect 11468 7624 11808 7710
rect 11468 7568 11536 7624
rect 11592 7568 11678 7624
rect 11734 7568 11808 7624
rect 11468 7482 11808 7568
rect 11468 7426 11536 7482
rect 11592 7426 11678 7482
rect 11734 7426 11808 7482
rect 11468 7340 11808 7426
rect 11468 7284 11536 7340
rect 11592 7284 11678 7340
rect 11734 7284 11808 7340
rect 11468 7198 11808 7284
rect 11468 7142 11536 7198
rect 11592 7142 11678 7198
rect 11734 7142 11808 7198
rect 11468 7056 11808 7142
rect 11468 7000 11536 7056
rect 11592 7000 11678 7056
rect 11734 7000 11808 7056
rect 11468 6914 11808 7000
rect 11468 6858 11536 6914
rect 11592 6858 11678 6914
rect 11734 6858 11808 6914
rect 11468 6772 11808 6858
rect 11468 6716 11536 6772
rect 11592 6716 11678 6772
rect 11734 6716 11808 6772
rect 11468 6630 11808 6716
rect 11468 6574 11536 6630
rect 11592 6574 11678 6630
rect 11734 6574 11808 6630
rect 11468 6488 11808 6574
rect 11468 6432 11536 6488
rect 11592 6432 11678 6488
rect 11734 6432 11808 6488
rect 11468 6346 11808 6432
rect 11468 6290 11536 6346
rect 11592 6290 11678 6346
rect 11734 6290 11808 6346
rect 11468 6204 11808 6290
rect 11468 6148 11536 6204
rect 11592 6148 11678 6204
rect 11734 6148 11808 6204
rect 11468 6062 11808 6148
rect 11468 6006 11536 6062
rect 11592 6006 11678 6062
rect 11734 6006 11808 6062
rect 11468 5920 11808 6006
rect 11468 5864 11536 5920
rect 11592 5864 11678 5920
rect 11734 5864 11808 5920
rect 11468 5778 11808 5864
rect 11468 5722 11536 5778
rect 11592 5722 11678 5778
rect 11734 5722 11808 5778
rect 11468 5636 11808 5722
rect 11468 5580 11536 5636
rect 11592 5580 11678 5636
rect 11734 5580 11808 5636
rect 11468 5494 11808 5580
rect 11468 5438 11536 5494
rect 11592 5438 11678 5494
rect 11734 5438 11808 5494
rect 11468 5352 11808 5438
rect 11468 5296 11536 5352
rect 11592 5296 11678 5352
rect 11734 5296 11808 5352
rect 11468 5210 11808 5296
rect 11468 5154 11536 5210
rect 11592 5154 11678 5210
rect 11734 5154 11808 5210
rect 11468 5068 11808 5154
rect 11468 5012 11536 5068
rect 11592 5012 11678 5068
rect 11734 5012 11808 5068
rect 11468 4926 11808 5012
rect 11468 4870 11536 4926
rect 11592 4870 11678 4926
rect 11734 4870 11808 4926
rect 11468 4784 11808 4870
rect 11468 4728 11536 4784
rect 11592 4728 11678 4784
rect 11734 4728 11808 4784
rect 11468 4642 11808 4728
rect 11468 4586 11536 4642
rect 11592 4586 11678 4642
rect 11734 4586 11808 4642
rect 11468 4500 11808 4586
rect 11468 4444 11536 4500
rect 11592 4444 11678 4500
rect 11734 4444 11808 4500
rect 11468 4358 11808 4444
rect 11468 4302 11536 4358
rect 11592 4302 11678 4358
rect 11734 4302 11808 4358
rect 11468 4216 11808 4302
rect 11468 4160 11536 4216
rect 11592 4160 11678 4216
rect 11734 4160 11808 4216
rect 11468 4074 11808 4160
rect 11468 4018 11536 4074
rect 11592 4018 11678 4074
rect 11734 4018 11808 4074
rect 11468 3932 11808 4018
rect 11468 3876 11536 3932
rect 11592 3876 11678 3932
rect 11734 3876 11808 3932
rect 11468 3790 11808 3876
rect 11468 3734 11536 3790
rect 11592 3734 11678 3790
rect 11734 3734 11808 3790
rect 11468 3648 11808 3734
rect 11468 3592 11536 3648
rect 11592 3592 11678 3648
rect 11734 3592 11808 3648
rect 11468 3506 11808 3592
rect 11468 3450 11536 3506
rect 11592 3450 11678 3506
rect 11734 3450 11808 3506
rect 11468 3364 11808 3450
rect 11468 3308 11536 3364
rect 11592 3308 11678 3364
rect 11734 3308 11808 3364
rect 11468 3222 11808 3308
rect 11468 3166 11536 3222
rect 11592 3166 11678 3222
rect 11734 3166 11808 3222
rect 11468 3080 11808 3166
rect 11468 3024 11536 3080
rect 11592 3024 11678 3080
rect 11734 3024 11808 3080
rect 11468 2938 11808 3024
rect 11468 2882 11536 2938
rect 11592 2882 11678 2938
rect 11734 2882 11808 2938
rect 11468 2796 11808 2882
rect 11468 2740 11536 2796
rect 11592 2740 11678 2796
rect 11734 2740 11808 2796
rect 11468 2654 11808 2740
rect 11468 2598 11536 2654
rect 11592 2598 11678 2654
rect 11734 2598 11808 2654
rect 11468 2512 11808 2598
rect 11468 2456 11536 2512
rect 11592 2456 11678 2512
rect 11734 2456 11808 2512
rect 11468 2370 11808 2456
rect 11468 2314 11536 2370
rect 11592 2314 11678 2370
rect 11734 2314 11808 2370
rect 11468 2228 11808 2314
rect 11468 2172 11536 2228
rect 11592 2172 11678 2228
rect 11734 2172 11808 2228
rect 11468 2086 11808 2172
rect 11468 2030 11536 2086
rect 11592 2030 11678 2086
rect 11734 2030 11808 2086
rect 11468 1944 11808 2030
rect 11468 1888 11536 1944
rect 11592 1888 11678 1944
rect 11734 1888 11808 1944
rect 11468 1802 11808 1888
rect 11468 1746 11536 1802
rect 11592 1746 11678 1802
rect 11734 1746 11808 1802
rect 11468 1660 11808 1746
rect 11468 1604 11536 1660
rect 11592 1604 11678 1660
rect 11734 1604 11808 1660
rect 11468 1518 11808 1604
rect 11468 1462 11536 1518
rect 11592 1462 11678 1518
rect 11734 1462 11808 1518
rect 11468 1376 11808 1462
rect 11468 1320 11536 1376
rect 11592 1320 11678 1376
rect 11734 1320 11808 1376
rect 11468 1234 11808 1320
rect 11468 1178 11536 1234
rect 11592 1178 11678 1234
rect 11734 1178 11808 1234
rect 11468 1092 11808 1178
rect 11468 1036 11536 1092
rect 11592 1036 11678 1092
rect 11734 1036 11808 1092
rect 11468 950 11808 1036
rect 11468 894 11536 950
rect 11592 894 11678 950
rect 11734 894 11808 950
rect 11468 808 11808 894
rect 11468 752 11536 808
rect 11592 752 11678 808
rect 11734 752 11808 808
rect 11468 666 11808 752
rect 11468 610 11536 666
rect 11592 610 11678 666
rect 11734 610 11808 666
rect 11468 524 11808 610
rect 11468 468 11536 524
rect 11592 468 11678 524
rect 11734 468 11808 524
rect 11468 400 11808 468
rect 11868 12310 12208 12400
rect 11868 12254 11941 12310
rect 11997 12254 12083 12310
rect 12139 12254 12208 12310
rect 11868 12168 12208 12254
rect 11868 12112 11941 12168
rect 11997 12112 12083 12168
rect 12139 12112 12208 12168
rect 11868 12026 12208 12112
rect 11868 11970 11941 12026
rect 11997 11970 12083 12026
rect 12139 11970 12208 12026
rect 11868 11884 12208 11970
rect 11868 11828 11941 11884
rect 11997 11828 12083 11884
rect 12139 11828 12208 11884
rect 11868 11742 12208 11828
rect 11868 11686 11941 11742
rect 11997 11686 12083 11742
rect 12139 11686 12208 11742
rect 11868 11600 12208 11686
rect 11868 11544 11941 11600
rect 11997 11544 12083 11600
rect 12139 11544 12208 11600
rect 11868 11458 12208 11544
rect 11868 11402 11941 11458
rect 11997 11402 12083 11458
rect 12139 11402 12208 11458
rect 11868 11316 12208 11402
rect 11868 11260 11941 11316
rect 11997 11260 12083 11316
rect 12139 11260 12208 11316
rect 11868 11174 12208 11260
rect 11868 11118 11941 11174
rect 11997 11118 12083 11174
rect 12139 11118 12208 11174
rect 11868 11032 12208 11118
rect 11868 10976 11941 11032
rect 11997 10976 12083 11032
rect 12139 10976 12208 11032
rect 11868 10890 12208 10976
rect 11868 10834 11941 10890
rect 11997 10834 12083 10890
rect 12139 10834 12208 10890
rect 11868 10748 12208 10834
rect 11868 10692 11941 10748
rect 11997 10692 12083 10748
rect 12139 10692 12208 10748
rect 11868 10606 12208 10692
rect 11868 10550 11941 10606
rect 11997 10550 12083 10606
rect 12139 10550 12208 10606
rect 11868 10464 12208 10550
rect 11868 10408 11941 10464
rect 11997 10408 12083 10464
rect 12139 10408 12208 10464
rect 11868 10322 12208 10408
rect 11868 10266 11941 10322
rect 11997 10266 12083 10322
rect 12139 10266 12208 10322
rect 11868 10180 12208 10266
rect 11868 10124 11941 10180
rect 11997 10124 12083 10180
rect 12139 10124 12208 10180
rect 11868 10038 12208 10124
rect 11868 9982 11941 10038
rect 11997 9982 12083 10038
rect 12139 9982 12208 10038
rect 11868 9896 12208 9982
rect 11868 9840 11941 9896
rect 11997 9840 12083 9896
rect 12139 9840 12208 9896
rect 11868 9754 12208 9840
rect 11868 9698 11941 9754
rect 11997 9698 12083 9754
rect 12139 9698 12208 9754
rect 11868 9612 12208 9698
rect 11868 9556 11941 9612
rect 11997 9556 12083 9612
rect 12139 9556 12208 9612
rect 11868 9470 12208 9556
rect 11868 9414 11941 9470
rect 11997 9414 12083 9470
rect 12139 9414 12208 9470
rect 11868 9328 12208 9414
rect 11868 9272 11941 9328
rect 11997 9272 12083 9328
rect 12139 9272 12208 9328
rect 11868 9186 12208 9272
rect 11868 9130 11941 9186
rect 11997 9130 12083 9186
rect 12139 9130 12208 9186
rect 11868 9044 12208 9130
rect 11868 8988 11941 9044
rect 11997 8988 12083 9044
rect 12139 8988 12208 9044
rect 11868 8902 12208 8988
rect 11868 8846 11941 8902
rect 11997 8846 12083 8902
rect 12139 8846 12208 8902
rect 11868 8760 12208 8846
rect 11868 8704 11941 8760
rect 11997 8704 12083 8760
rect 12139 8704 12208 8760
rect 11868 8618 12208 8704
rect 11868 8562 11941 8618
rect 11997 8562 12083 8618
rect 12139 8562 12208 8618
rect 11868 8476 12208 8562
rect 11868 8420 11941 8476
rect 11997 8420 12083 8476
rect 12139 8420 12208 8476
rect 11868 8334 12208 8420
rect 11868 8278 11941 8334
rect 11997 8278 12083 8334
rect 12139 8278 12208 8334
rect 11868 8192 12208 8278
rect 11868 8136 11941 8192
rect 11997 8136 12083 8192
rect 12139 8136 12208 8192
rect 11868 8050 12208 8136
rect 11868 7994 11941 8050
rect 11997 7994 12083 8050
rect 12139 7994 12208 8050
rect 11868 7908 12208 7994
rect 11868 7852 11941 7908
rect 11997 7852 12083 7908
rect 12139 7852 12208 7908
rect 11868 7766 12208 7852
rect 11868 7710 11941 7766
rect 11997 7710 12083 7766
rect 12139 7710 12208 7766
rect 11868 7624 12208 7710
rect 11868 7568 11941 7624
rect 11997 7568 12083 7624
rect 12139 7568 12208 7624
rect 11868 7482 12208 7568
rect 11868 7426 11941 7482
rect 11997 7426 12083 7482
rect 12139 7426 12208 7482
rect 11868 7340 12208 7426
rect 11868 7284 11941 7340
rect 11997 7284 12083 7340
rect 12139 7284 12208 7340
rect 11868 7198 12208 7284
rect 11868 7142 11941 7198
rect 11997 7142 12083 7198
rect 12139 7142 12208 7198
rect 11868 7056 12208 7142
rect 11868 7000 11941 7056
rect 11997 7000 12083 7056
rect 12139 7000 12208 7056
rect 11868 6914 12208 7000
rect 11868 6858 11941 6914
rect 11997 6858 12083 6914
rect 12139 6858 12208 6914
rect 11868 6772 12208 6858
rect 11868 6716 11941 6772
rect 11997 6716 12083 6772
rect 12139 6716 12208 6772
rect 11868 6630 12208 6716
rect 11868 6574 11941 6630
rect 11997 6574 12083 6630
rect 12139 6574 12208 6630
rect 11868 6488 12208 6574
rect 11868 6432 11941 6488
rect 11997 6432 12083 6488
rect 12139 6432 12208 6488
rect 11868 6346 12208 6432
rect 11868 6290 11941 6346
rect 11997 6290 12083 6346
rect 12139 6290 12208 6346
rect 11868 6204 12208 6290
rect 11868 6148 11941 6204
rect 11997 6148 12083 6204
rect 12139 6148 12208 6204
rect 11868 6062 12208 6148
rect 11868 6006 11941 6062
rect 11997 6006 12083 6062
rect 12139 6006 12208 6062
rect 11868 5920 12208 6006
rect 11868 5864 11941 5920
rect 11997 5864 12083 5920
rect 12139 5864 12208 5920
rect 11868 5778 12208 5864
rect 11868 5722 11941 5778
rect 11997 5722 12083 5778
rect 12139 5722 12208 5778
rect 11868 5636 12208 5722
rect 11868 5580 11941 5636
rect 11997 5580 12083 5636
rect 12139 5580 12208 5636
rect 11868 5494 12208 5580
rect 11868 5438 11941 5494
rect 11997 5438 12083 5494
rect 12139 5438 12208 5494
rect 11868 5352 12208 5438
rect 11868 5296 11941 5352
rect 11997 5296 12083 5352
rect 12139 5296 12208 5352
rect 11868 5210 12208 5296
rect 11868 5154 11941 5210
rect 11997 5154 12083 5210
rect 12139 5154 12208 5210
rect 11868 5068 12208 5154
rect 11868 5012 11941 5068
rect 11997 5012 12083 5068
rect 12139 5012 12208 5068
rect 11868 4926 12208 5012
rect 11868 4870 11941 4926
rect 11997 4870 12083 4926
rect 12139 4870 12208 4926
rect 11868 4784 12208 4870
rect 11868 4728 11941 4784
rect 11997 4728 12083 4784
rect 12139 4728 12208 4784
rect 11868 4642 12208 4728
rect 11868 4586 11941 4642
rect 11997 4586 12083 4642
rect 12139 4586 12208 4642
rect 11868 4500 12208 4586
rect 11868 4444 11941 4500
rect 11997 4444 12083 4500
rect 12139 4444 12208 4500
rect 11868 4358 12208 4444
rect 11868 4302 11941 4358
rect 11997 4302 12083 4358
rect 12139 4302 12208 4358
rect 11868 4216 12208 4302
rect 11868 4160 11941 4216
rect 11997 4160 12083 4216
rect 12139 4160 12208 4216
rect 11868 4074 12208 4160
rect 11868 4018 11941 4074
rect 11997 4018 12083 4074
rect 12139 4018 12208 4074
rect 11868 3932 12208 4018
rect 11868 3876 11941 3932
rect 11997 3876 12083 3932
rect 12139 3876 12208 3932
rect 11868 3790 12208 3876
rect 11868 3734 11941 3790
rect 11997 3734 12083 3790
rect 12139 3734 12208 3790
rect 11868 3648 12208 3734
rect 11868 3592 11941 3648
rect 11997 3592 12083 3648
rect 12139 3592 12208 3648
rect 11868 3506 12208 3592
rect 11868 3450 11941 3506
rect 11997 3450 12083 3506
rect 12139 3450 12208 3506
rect 11868 3364 12208 3450
rect 11868 3308 11941 3364
rect 11997 3308 12083 3364
rect 12139 3308 12208 3364
rect 11868 3222 12208 3308
rect 11868 3166 11941 3222
rect 11997 3166 12083 3222
rect 12139 3166 12208 3222
rect 11868 3080 12208 3166
rect 11868 3024 11941 3080
rect 11997 3024 12083 3080
rect 12139 3024 12208 3080
rect 11868 2938 12208 3024
rect 11868 2882 11941 2938
rect 11997 2882 12083 2938
rect 12139 2882 12208 2938
rect 11868 2796 12208 2882
rect 11868 2740 11941 2796
rect 11997 2740 12083 2796
rect 12139 2740 12208 2796
rect 11868 2654 12208 2740
rect 11868 2598 11941 2654
rect 11997 2598 12083 2654
rect 12139 2598 12208 2654
rect 11868 2512 12208 2598
rect 11868 2456 11941 2512
rect 11997 2456 12083 2512
rect 12139 2456 12208 2512
rect 11868 2370 12208 2456
rect 11868 2314 11941 2370
rect 11997 2314 12083 2370
rect 12139 2314 12208 2370
rect 11868 2228 12208 2314
rect 11868 2172 11941 2228
rect 11997 2172 12083 2228
rect 12139 2172 12208 2228
rect 11868 2086 12208 2172
rect 11868 2030 11941 2086
rect 11997 2030 12083 2086
rect 12139 2030 12208 2086
rect 11868 1944 12208 2030
rect 11868 1888 11941 1944
rect 11997 1888 12083 1944
rect 12139 1888 12208 1944
rect 11868 1802 12208 1888
rect 11868 1746 11941 1802
rect 11997 1746 12083 1802
rect 12139 1746 12208 1802
rect 11868 1660 12208 1746
rect 11868 1604 11941 1660
rect 11997 1604 12083 1660
rect 12139 1604 12208 1660
rect 11868 1518 12208 1604
rect 11868 1462 11941 1518
rect 11997 1462 12083 1518
rect 12139 1462 12208 1518
rect 11868 1376 12208 1462
rect 11868 1320 11941 1376
rect 11997 1320 12083 1376
rect 12139 1320 12208 1376
rect 11868 1234 12208 1320
rect 11868 1178 11941 1234
rect 11997 1178 12083 1234
rect 12139 1178 12208 1234
rect 11868 1092 12208 1178
rect 11868 1036 11941 1092
rect 11997 1036 12083 1092
rect 12139 1036 12208 1092
rect 11868 950 12208 1036
rect 11868 894 11941 950
rect 11997 894 12083 950
rect 12139 894 12208 950
rect 11868 808 12208 894
rect 11868 752 11941 808
rect 11997 752 12083 808
rect 12139 752 12208 808
rect 11868 666 12208 752
rect 11868 610 11941 666
rect 11997 610 12083 666
rect 12139 610 12208 666
rect 11868 524 12208 610
rect 11868 468 11941 524
rect 11997 468 12083 524
rect 12139 468 12208 524
rect 11868 400 12208 468
rect 12400 12358 13200 12400
rect 12400 12302 12526 12358
rect 12582 12302 12650 12358
rect 12706 12302 12774 12358
rect 12830 12302 12898 12358
rect 12954 12302 13022 12358
rect 13078 12302 13200 12358
rect 12400 12234 13200 12302
rect 12400 12178 12526 12234
rect 12582 12178 12650 12234
rect 12706 12178 12774 12234
rect 12830 12178 12898 12234
rect 12954 12178 13022 12234
rect 13078 12178 13200 12234
rect 12400 12110 13200 12178
rect 12400 12054 12526 12110
rect 12582 12054 12650 12110
rect 12706 12054 12774 12110
rect 12830 12054 12898 12110
rect 12954 12054 13022 12110
rect 13078 12054 13200 12110
rect 12400 11986 13200 12054
rect 12400 11930 12526 11986
rect 12582 11930 12650 11986
rect 12706 11930 12774 11986
rect 12830 11930 12898 11986
rect 12954 11930 13022 11986
rect 13078 11930 13200 11986
rect 12400 11862 13200 11930
rect 12400 11806 12526 11862
rect 12582 11806 12650 11862
rect 12706 11806 12774 11862
rect 12830 11806 12898 11862
rect 12954 11806 13022 11862
rect 13078 11806 13200 11862
rect 12400 11738 13200 11806
rect 12400 11682 12526 11738
rect 12582 11682 12650 11738
rect 12706 11682 12774 11738
rect 12830 11682 12898 11738
rect 12954 11682 13022 11738
rect 13078 11682 13200 11738
rect 12400 11614 13200 11682
rect 12400 11558 12526 11614
rect 12582 11558 12650 11614
rect 12706 11558 12774 11614
rect 12830 11558 12898 11614
rect 12954 11558 13022 11614
rect 13078 11558 13200 11614
rect 12400 11490 13200 11558
rect 12400 11434 12526 11490
rect 12582 11434 12650 11490
rect 12706 11434 12774 11490
rect 12830 11434 12898 11490
rect 12954 11434 13022 11490
rect 13078 11434 13200 11490
rect 12400 11366 13200 11434
rect 12400 11310 12526 11366
rect 12582 11310 12650 11366
rect 12706 11310 12774 11366
rect 12830 11310 12898 11366
rect 12954 11310 13022 11366
rect 13078 11310 13200 11366
rect 12400 11242 13200 11310
rect 12400 11186 12526 11242
rect 12582 11186 12650 11242
rect 12706 11186 12774 11242
rect 12830 11186 12898 11242
rect 12954 11186 13022 11242
rect 13078 11186 13200 11242
rect 12400 11118 13200 11186
rect 12400 11062 12526 11118
rect 12582 11062 12650 11118
rect 12706 11062 12774 11118
rect 12830 11062 12898 11118
rect 12954 11062 13022 11118
rect 13078 11062 13200 11118
rect 12400 10994 13200 11062
rect 12400 10938 12526 10994
rect 12582 10938 12650 10994
rect 12706 10938 12774 10994
rect 12830 10938 12898 10994
rect 12954 10938 13022 10994
rect 13078 10938 13200 10994
rect 12400 10870 13200 10938
rect 12400 10814 12526 10870
rect 12582 10814 12650 10870
rect 12706 10814 12774 10870
rect 12830 10814 12898 10870
rect 12954 10814 13022 10870
rect 13078 10814 13200 10870
rect 12400 10746 13200 10814
rect 12400 10690 12526 10746
rect 12582 10690 12650 10746
rect 12706 10690 12774 10746
rect 12830 10690 12898 10746
rect 12954 10690 13022 10746
rect 13078 10690 13200 10746
rect 12400 10622 13200 10690
rect 12400 10566 12526 10622
rect 12582 10566 12650 10622
rect 12706 10566 12774 10622
rect 12830 10566 12898 10622
rect 12954 10566 13022 10622
rect 13078 10566 13200 10622
rect 12400 10498 13200 10566
rect 12400 10442 12526 10498
rect 12582 10442 12650 10498
rect 12706 10442 12774 10498
rect 12830 10442 12898 10498
rect 12954 10442 13022 10498
rect 13078 10442 13200 10498
rect 12400 10374 13200 10442
rect 12400 10318 12526 10374
rect 12582 10318 12650 10374
rect 12706 10318 12774 10374
rect 12830 10318 12898 10374
rect 12954 10318 13022 10374
rect 13078 10318 13200 10374
rect 12400 10250 13200 10318
rect 12400 10194 12526 10250
rect 12582 10194 12650 10250
rect 12706 10194 12774 10250
rect 12830 10194 12898 10250
rect 12954 10194 13022 10250
rect 13078 10194 13200 10250
rect 12400 10126 13200 10194
rect 12400 10070 12526 10126
rect 12582 10070 12650 10126
rect 12706 10070 12774 10126
rect 12830 10070 12898 10126
rect 12954 10070 13022 10126
rect 13078 10070 13200 10126
rect 12400 10002 13200 10070
rect 12400 9946 12526 10002
rect 12582 9946 12650 10002
rect 12706 9946 12774 10002
rect 12830 9946 12898 10002
rect 12954 9946 13022 10002
rect 13078 9946 13200 10002
rect 12400 9878 13200 9946
rect 12400 9822 12526 9878
rect 12582 9822 12650 9878
rect 12706 9822 12774 9878
rect 12830 9822 12898 9878
rect 12954 9822 13022 9878
rect 13078 9822 13200 9878
rect 12400 9754 13200 9822
rect 12400 9698 12526 9754
rect 12582 9698 12650 9754
rect 12706 9698 12774 9754
rect 12830 9698 12898 9754
rect 12954 9698 13022 9754
rect 13078 9698 13200 9754
rect 12400 9630 13200 9698
rect 12400 9574 12526 9630
rect 12582 9574 12650 9630
rect 12706 9574 12774 9630
rect 12830 9574 12898 9630
rect 12954 9574 13022 9630
rect 13078 9574 13200 9630
rect 12400 9506 13200 9574
rect 12400 9450 12526 9506
rect 12582 9450 12650 9506
rect 12706 9450 12774 9506
rect 12830 9450 12898 9506
rect 12954 9450 13022 9506
rect 13078 9450 13200 9506
rect 12400 9382 13200 9450
rect 12400 9326 12526 9382
rect 12582 9326 12650 9382
rect 12706 9326 12774 9382
rect 12830 9326 12898 9382
rect 12954 9326 13022 9382
rect 13078 9326 13200 9382
rect 12400 9258 13200 9326
rect 12400 9202 12526 9258
rect 12582 9202 12650 9258
rect 12706 9202 12774 9258
rect 12830 9202 12898 9258
rect 12954 9202 13022 9258
rect 13078 9202 13200 9258
rect 12400 9134 13200 9202
rect 12400 9078 12526 9134
rect 12582 9078 12650 9134
rect 12706 9078 12774 9134
rect 12830 9078 12898 9134
rect 12954 9078 13022 9134
rect 13078 9078 13200 9134
rect 12400 9010 13200 9078
rect 12400 8954 12526 9010
rect 12582 8954 12650 9010
rect 12706 8954 12774 9010
rect 12830 8954 12898 9010
rect 12954 8954 13022 9010
rect 13078 8954 13200 9010
rect 12400 8886 13200 8954
rect 12400 8830 12526 8886
rect 12582 8830 12650 8886
rect 12706 8830 12774 8886
rect 12830 8830 12898 8886
rect 12954 8830 13022 8886
rect 13078 8830 13200 8886
rect 12400 8762 13200 8830
rect 12400 8706 12526 8762
rect 12582 8706 12650 8762
rect 12706 8706 12774 8762
rect 12830 8706 12898 8762
rect 12954 8706 13022 8762
rect 13078 8706 13200 8762
rect 12400 8638 13200 8706
rect 12400 8582 12526 8638
rect 12582 8582 12650 8638
rect 12706 8582 12774 8638
rect 12830 8582 12898 8638
rect 12954 8582 13022 8638
rect 13078 8582 13200 8638
rect 12400 8514 13200 8582
rect 12400 8458 12526 8514
rect 12582 8458 12650 8514
rect 12706 8458 12774 8514
rect 12830 8458 12898 8514
rect 12954 8458 13022 8514
rect 13078 8458 13200 8514
rect 12400 8390 13200 8458
rect 12400 8334 12526 8390
rect 12582 8334 12650 8390
rect 12706 8334 12774 8390
rect 12830 8334 12898 8390
rect 12954 8334 13022 8390
rect 13078 8334 13200 8390
rect 12400 8266 13200 8334
rect 12400 8210 12526 8266
rect 12582 8210 12650 8266
rect 12706 8210 12774 8266
rect 12830 8210 12898 8266
rect 12954 8210 13022 8266
rect 13078 8210 13200 8266
rect 12400 8142 13200 8210
rect 12400 8086 12526 8142
rect 12582 8086 12650 8142
rect 12706 8086 12774 8142
rect 12830 8086 12898 8142
rect 12954 8086 13022 8142
rect 13078 8086 13200 8142
rect 12400 8018 13200 8086
rect 12400 7962 12526 8018
rect 12582 7962 12650 8018
rect 12706 7962 12774 8018
rect 12830 7962 12898 8018
rect 12954 7962 13022 8018
rect 13078 7962 13200 8018
rect 12400 7894 13200 7962
rect 12400 7838 12526 7894
rect 12582 7838 12650 7894
rect 12706 7838 12774 7894
rect 12830 7838 12898 7894
rect 12954 7838 13022 7894
rect 13078 7838 13200 7894
rect 12400 7770 13200 7838
rect 12400 7714 12526 7770
rect 12582 7714 12650 7770
rect 12706 7714 12774 7770
rect 12830 7714 12898 7770
rect 12954 7714 13022 7770
rect 13078 7714 13200 7770
rect 12400 7646 13200 7714
rect 12400 7590 12526 7646
rect 12582 7590 12650 7646
rect 12706 7590 12774 7646
rect 12830 7590 12898 7646
rect 12954 7590 13022 7646
rect 13078 7590 13200 7646
rect 12400 7522 13200 7590
rect 12400 7466 12526 7522
rect 12582 7466 12650 7522
rect 12706 7466 12774 7522
rect 12830 7466 12898 7522
rect 12954 7466 13022 7522
rect 13078 7466 13200 7522
rect 12400 7398 13200 7466
rect 12400 7342 12526 7398
rect 12582 7342 12650 7398
rect 12706 7342 12774 7398
rect 12830 7342 12898 7398
rect 12954 7342 13022 7398
rect 13078 7342 13200 7398
rect 12400 7274 13200 7342
rect 12400 7218 12526 7274
rect 12582 7218 12650 7274
rect 12706 7218 12774 7274
rect 12830 7218 12898 7274
rect 12954 7218 13022 7274
rect 13078 7218 13200 7274
rect 12400 7150 13200 7218
rect 12400 7094 12526 7150
rect 12582 7094 12650 7150
rect 12706 7094 12774 7150
rect 12830 7094 12898 7150
rect 12954 7094 13022 7150
rect 13078 7094 13200 7150
rect 12400 7026 13200 7094
rect 12400 6970 12526 7026
rect 12582 6970 12650 7026
rect 12706 6970 12774 7026
rect 12830 6970 12898 7026
rect 12954 6970 13022 7026
rect 13078 6970 13200 7026
rect 12400 6902 13200 6970
rect 12400 6846 12526 6902
rect 12582 6846 12650 6902
rect 12706 6846 12774 6902
rect 12830 6846 12898 6902
rect 12954 6846 13022 6902
rect 13078 6846 13200 6902
rect 12400 6778 13200 6846
rect 12400 6722 12526 6778
rect 12582 6722 12650 6778
rect 12706 6722 12774 6778
rect 12830 6722 12898 6778
rect 12954 6722 13022 6778
rect 13078 6722 13200 6778
rect 12400 6654 13200 6722
rect 12400 6598 12526 6654
rect 12582 6598 12650 6654
rect 12706 6598 12774 6654
rect 12830 6598 12898 6654
rect 12954 6598 13022 6654
rect 13078 6598 13200 6654
rect 12400 6530 13200 6598
rect 12400 6474 12526 6530
rect 12582 6474 12650 6530
rect 12706 6474 12774 6530
rect 12830 6474 12898 6530
rect 12954 6474 13022 6530
rect 13078 6474 13200 6530
rect 12400 6406 13200 6474
rect 12400 6350 12526 6406
rect 12582 6350 12650 6406
rect 12706 6350 12774 6406
rect 12830 6350 12898 6406
rect 12954 6350 13022 6406
rect 13078 6350 13200 6406
rect 12400 6282 13200 6350
rect 12400 6226 12526 6282
rect 12582 6226 12650 6282
rect 12706 6226 12774 6282
rect 12830 6226 12898 6282
rect 12954 6226 13022 6282
rect 13078 6226 13200 6282
rect 12400 6158 13200 6226
rect 12400 6102 12526 6158
rect 12582 6102 12650 6158
rect 12706 6102 12774 6158
rect 12830 6102 12898 6158
rect 12954 6102 13022 6158
rect 13078 6102 13200 6158
rect 12400 6034 13200 6102
rect 12400 5978 12526 6034
rect 12582 5978 12650 6034
rect 12706 5978 12774 6034
rect 12830 5978 12898 6034
rect 12954 5978 13022 6034
rect 13078 5978 13200 6034
rect 12400 5910 13200 5978
rect 12400 5854 12526 5910
rect 12582 5854 12650 5910
rect 12706 5854 12774 5910
rect 12830 5854 12898 5910
rect 12954 5854 13022 5910
rect 13078 5854 13200 5910
rect 12400 5786 13200 5854
rect 12400 5730 12526 5786
rect 12582 5730 12650 5786
rect 12706 5730 12774 5786
rect 12830 5730 12898 5786
rect 12954 5730 13022 5786
rect 13078 5730 13200 5786
rect 12400 5662 13200 5730
rect 12400 5606 12526 5662
rect 12582 5606 12650 5662
rect 12706 5606 12774 5662
rect 12830 5606 12898 5662
rect 12954 5606 13022 5662
rect 13078 5606 13200 5662
rect 12400 5538 13200 5606
rect 12400 5482 12526 5538
rect 12582 5482 12650 5538
rect 12706 5482 12774 5538
rect 12830 5482 12898 5538
rect 12954 5482 13022 5538
rect 13078 5482 13200 5538
rect 12400 5414 13200 5482
rect 12400 5358 12526 5414
rect 12582 5358 12650 5414
rect 12706 5358 12774 5414
rect 12830 5358 12898 5414
rect 12954 5358 13022 5414
rect 13078 5358 13200 5414
rect 12400 5290 13200 5358
rect 12400 5234 12526 5290
rect 12582 5234 12650 5290
rect 12706 5234 12774 5290
rect 12830 5234 12898 5290
rect 12954 5234 13022 5290
rect 13078 5234 13200 5290
rect 12400 5166 13200 5234
rect 12400 5110 12526 5166
rect 12582 5110 12650 5166
rect 12706 5110 12774 5166
rect 12830 5110 12898 5166
rect 12954 5110 13022 5166
rect 13078 5110 13200 5166
rect 12400 5042 13200 5110
rect 12400 4986 12526 5042
rect 12582 4986 12650 5042
rect 12706 4986 12774 5042
rect 12830 4986 12898 5042
rect 12954 4986 13022 5042
rect 13078 4986 13200 5042
rect 12400 4918 13200 4986
rect 12400 4862 12526 4918
rect 12582 4862 12650 4918
rect 12706 4862 12774 4918
rect 12830 4862 12898 4918
rect 12954 4862 13022 4918
rect 13078 4862 13200 4918
rect 12400 4794 13200 4862
rect 12400 4738 12526 4794
rect 12582 4738 12650 4794
rect 12706 4738 12774 4794
rect 12830 4738 12898 4794
rect 12954 4738 13022 4794
rect 13078 4738 13200 4794
rect 12400 4670 13200 4738
rect 12400 4614 12526 4670
rect 12582 4614 12650 4670
rect 12706 4614 12774 4670
rect 12830 4614 12898 4670
rect 12954 4614 13022 4670
rect 13078 4614 13200 4670
rect 12400 4546 13200 4614
rect 12400 4490 12526 4546
rect 12582 4490 12650 4546
rect 12706 4490 12774 4546
rect 12830 4490 12898 4546
rect 12954 4490 13022 4546
rect 13078 4490 13200 4546
rect 12400 4422 13200 4490
rect 12400 4366 12526 4422
rect 12582 4366 12650 4422
rect 12706 4366 12774 4422
rect 12830 4366 12898 4422
rect 12954 4366 13022 4422
rect 13078 4366 13200 4422
rect 12400 4298 13200 4366
rect 12400 4242 12526 4298
rect 12582 4242 12650 4298
rect 12706 4242 12774 4298
rect 12830 4242 12898 4298
rect 12954 4242 13022 4298
rect 13078 4242 13200 4298
rect 12400 4174 13200 4242
rect 12400 4118 12526 4174
rect 12582 4118 12650 4174
rect 12706 4118 12774 4174
rect 12830 4118 12898 4174
rect 12954 4118 13022 4174
rect 13078 4118 13200 4174
rect 12400 4050 13200 4118
rect 12400 3994 12526 4050
rect 12582 3994 12650 4050
rect 12706 3994 12774 4050
rect 12830 3994 12898 4050
rect 12954 3994 13022 4050
rect 13078 3994 13200 4050
rect 12400 3926 13200 3994
rect 12400 3870 12526 3926
rect 12582 3870 12650 3926
rect 12706 3870 12774 3926
rect 12830 3870 12898 3926
rect 12954 3870 13022 3926
rect 13078 3870 13200 3926
rect 12400 3802 13200 3870
rect 12400 3746 12526 3802
rect 12582 3746 12650 3802
rect 12706 3746 12774 3802
rect 12830 3746 12898 3802
rect 12954 3746 13022 3802
rect 13078 3746 13200 3802
rect 12400 3678 13200 3746
rect 12400 3622 12526 3678
rect 12582 3622 12650 3678
rect 12706 3622 12774 3678
rect 12830 3622 12898 3678
rect 12954 3622 13022 3678
rect 13078 3622 13200 3678
rect 12400 3554 13200 3622
rect 12400 3498 12526 3554
rect 12582 3498 12650 3554
rect 12706 3498 12774 3554
rect 12830 3498 12898 3554
rect 12954 3498 13022 3554
rect 13078 3498 13200 3554
rect 12400 3430 13200 3498
rect 12400 3374 12526 3430
rect 12582 3374 12650 3430
rect 12706 3374 12774 3430
rect 12830 3374 12898 3430
rect 12954 3374 13022 3430
rect 13078 3374 13200 3430
rect 12400 3306 13200 3374
rect 12400 3250 12526 3306
rect 12582 3250 12650 3306
rect 12706 3250 12774 3306
rect 12830 3250 12898 3306
rect 12954 3250 13022 3306
rect 13078 3250 13200 3306
rect 12400 3182 13200 3250
rect 12400 3126 12526 3182
rect 12582 3126 12650 3182
rect 12706 3126 12774 3182
rect 12830 3126 12898 3182
rect 12954 3126 13022 3182
rect 13078 3126 13200 3182
rect 12400 3058 13200 3126
rect 12400 3002 12526 3058
rect 12582 3002 12650 3058
rect 12706 3002 12774 3058
rect 12830 3002 12898 3058
rect 12954 3002 13022 3058
rect 13078 3002 13200 3058
rect 12400 2934 13200 3002
rect 12400 2878 12526 2934
rect 12582 2878 12650 2934
rect 12706 2878 12774 2934
rect 12830 2878 12898 2934
rect 12954 2878 13022 2934
rect 13078 2878 13200 2934
rect 12400 2810 13200 2878
rect 12400 2754 12526 2810
rect 12582 2754 12650 2810
rect 12706 2754 12774 2810
rect 12830 2754 12898 2810
rect 12954 2754 13022 2810
rect 13078 2754 13200 2810
rect 12400 2686 13200 2754
rect 12400 2630 12526 2686
rect 12582 2630 12650 2686
rect 12706 2630 12774 2686
rect 12830 2630 12898 2686
rect 12954 2630 13022 2686
rect 13078 2630 13200 2686
rect 12400 2562 13200 2630
rect 12400 2506 12526 2562
rect 12582 2506 12650 2562
rect 12706 2506 12774 2562
rect 12830 2506 12898 2562
rect 12954 2506 13022 2562
rect 13078 2506 13200 2562
rect 12400 2438 13200 2506
rect 12400 2382 12526 2438
rect 12582 2382 12650 2438
rect 12706 2382 12774 2438
rect 12830 2382 12898 2438
rect 12954 2382 13022 2438
rect 13078 2382 13200 2438
rect 12400 2314 13200 2382
rect 12400 2258 12526 2314
rect 12582 2258 12650 2314
rect 12706 2258 12774 2314
rect 12830 2258 12898 2314
rect 12954 2258 13022 2314
rect 13078 2258 13200 2314
rect 12400 2190 13200 2258
rect 12400 2134 12526 2190
rect 12582 2134 12650 2190
rect 12706 2134 12774 2190
rect 12830 2134 12898 2190
rect 12954 2134 13022 2190
rect 13078 2134 13200 2190
rect 12400 2066 13200 2134
rect 12400 2010 12526 2066
rect 12582 2010 12650 2066
rect 12706 2010 12774 2066
rect 12830 2010 12898 2066
rect 12954 2010 13022 2066
rect 13078 2010 13200 2066
rect 12400 1942 13200 2010
rect 12400 1886 12526 1942
rect 12582 1886 12650 1942
rect 12706 1886 12774 1942
rect 12830 1886 12898 1942
rect 12954 1886 13022 1942
rect 13078 1886 13200 1942
rect 12400 1818 13200 1886
rect 12400 1762 12526 1818
rect 12582 1762 12650 1818
rect 12706 1762 12774 1818
rect 12830 1762 12898 1818
rect 12954 1762 13022 1818
rect 13078 1762 13200 1818
rect 12400 1694 13200 1762
rect 12400 1638 12526 1694
rect 12582 1638 12650 1694
rect 12706 1638 12774 1694
rect 12830 1638 12898 1694
rect 12954 1638 13022 1694
rect 13078 1638 13200 1694
rect 12400 1570 13200 1638
rect 12400 1514 12526 1570
rect 12582 1514 12650 1570
rect 12706 1514 12774 1570
rect 12830 1514 12898 1570
rect 12954 1514 13022 1570
rect 13078 1514 13200 1570
rect 12400 1446 13200 1514
rect 12400 1390 12526 1446
rect 12582 1390 12650 1446
rect 12706 1390 12774 1446
rect 12830 1390 12898 1446
rect 12954 1390 13022 1446
rect 13078 1390 13200 1446
rect 12400 1322 13200 1390
rect 12400 1266 12526 1322
rect 12582 1266 12650 1322
rect 12706 1266 12774 1322
rect 12830 1266 12898 1322
rect 12954 1266 13022 1322
rect 13078 1266 13200 1322
rect 12400 1198 13200 1266
rect 12400 1142 12526 1198
rect 12582 1142 12650 1198
rect 12706 1142 12774 1198
rect 12830 1142 12898 1198
rect 12954 1142 13022 1198
rect 13078 1142 13200 1198
rect 12400 1074 13200 1142
rect 12400 1018 12526 1074
rect 12582 1018 12650 1074
rect 12706 1018 12774 1074
rect 12830 1018 12898 1074
rect 12954 1018 13022 1074
rect 13078 1018 13200 1074
rect 12400 950 13200 1018
rect 12400 894 12526 950
rect 12582 894 12650 950
rect 12706 894 12774 950
rect 12830 894 12898 950
rect 12954 894 13022 950
rect 13078 894 13200 950
rect 12400 826 13200 894
rect 12400 770 12526 826
rect 12582 770 12650 826
rect 12706 770 12774 826
rect 12830 770 12898 826
rect 12954 770 13022 826
rect 13078 770 13200 826
rect 12400 702 13200 770
rect 12400 646 12526 702
rect 12582 646 12650 702
rect 12706 646 12774 702
rect 12830 646 12898 702
rect 12954 646 13022 702
rect 13078 646 13200 702
rect 12400 578 13200 646
rect 12400 522 12526 578
rect 12582 522 12650 578
rect 12706 522 12774 578
rect 12830 522 12898 578
rect 12954 522 13022 578
rect 13078 522 13200 578
rect 12400 454 13200 522
rect 12400 400 12526 454
rect 266 398 12526 400
rect 12582 398 12650 454
rect 12706 398 12774 454
rect 12830 398 12898 454
rect 12954 398 13022 454
rect 13078 398 13200 454
rect -400 330 13200 398
rect -400 274 -286 330
rect -230 274 -162 330
rect -106 274 -38 330
rect 18 274 86 330
rect 142 274 210 330
rect 266 302 12526 330
rect 266 274 415 302
rect -400 246 415 274
rect 471 246 557 302
rect 613 246 699 302
rect 755 246 841 302
rect 897 246 983 302
rect 1039 246 1125 302
rect 1181 246 1267 302
rect 1323 246 1409 302
rect 1465 246 1551 302
rect 1607 246 1693 302
rect 1749 246 1835 302
rect 1891 246 1977 302
rect 2033 246 2119 302
rect 2175 246 2261 302
rect 2317 246 2403 302
rect 2459 246 2545 302
rect 2601 246 2687 302
rect 2743 246 2829 302
rect 2885 246 2971 302
rect 3027 246 3113 302
rect 3169 246 3255 302
rect 3311 246 3397 302
rect 3453 246 3539 302
rect 3595 246 3681 302
rect 3737 246 3823 302
rect 3879 246 3965 302
rect 4021 246 4107 302
rect 4163 246 4249 302
rect 4305 246 4391 302
rect 4447 246 4533 302
rect 4589 246 4675 302
rect 4731 246 4817 302
rect 4873 246 4959 302
rect 5015 246 5101 302
rect 5157 246 5243 302
rect 5299 246 5385 302
rect 5441 246 5527 302
rect 5583 246 5669 302
rect 5725 246 5811 302
rect 5867 246 5953 302
rect 6009 246 6095 302
rect 6151 246 6237 302
rect 6293 246 6379 302
rect 6435 246 6521 302
rect 6577 246 6663 302
rect 6719 246 6805 302
rect 6861 246 6947 302
rect 7003 246 7089 302
rect 7145 246 7231 302
rect 7287 246 7373 302
rect 7429 246 7515 302
rect 7571 246 7657 302
rect 7713 246 7799 302
rect 7855 246 7941 302
rect 7997 246 8083 302
rect 8139 246 8225 302
rect 8281 246 8367 302
rect 8423 246 8509 302
rect 8565 246 8651 302
rect 8707 246 8793 302
rect 8849 246 8935 302
rect 8991 246 9077 302
rect 9133 246 9219 302
rect 9275 246 9361 302
rect 9417 246 9503 302
rect 9559 246 9645 302
rect 9701 246 9787 302
rect 9843 246 9929 302
rect 9985 246 10071 302
rect 10127 246 10213 302
rect 10269 246 10355 302
rect 10411 246 10497 302
rect 10553 246 10639 302
rect 10695 246 10781 302
rect 10837 246 10923 302
rect 10979 246 11065 302
rect 11121 246 11207 302
rect 11263 246 11349 302
rect 11405 246 11491 302
rect 11547 246 11633 302
rect 11689 246 11775 302
rect 11831 246 11917 302
rect 11973 246 12059 302
rect 12115 246 12201 302
rect 12257 246 12343 302
rect 12399 274 12526 302
rect 12582 274 12650 330
rect 12706 274 12774 330
rect 12830 274 12898 330
rect 12954 274 13022 330
rect 13078 274 13200 330
rect 12399 246 13200 274
rect -400 206 13200 246
rect -400 150 -286 206
rect -230 150 -162 206
rect -106 150 -38 206
rect 18 150 86 206
rect 142 150 210 206
rect 266 160 12526 206
rect 266 150 415 160
rect -400 104 415 150
rect 471 104 557 160
rect 613 104 699 160
rect 755 104 841 160
rect 897 104 983 160
rect 1039 104 1125 160
rect 1181 104 1267 160
rect 1323 104 1409 160
rect 1465 104 1551 160
rect 1607 104 1693 160
rect 1749 104 1835 160
rect 1891 104 1977 160
rect 2033 104 2119 160
rect 2175 104 2261 160
rect 2317 104 2403 160
rect 2459 104 2545 160
rect 2601 104 2687 160
rect 2743 104 2829 160
rect 2885 104 2971 160
rect 3027 104 3113 160
rect 3169 104 3255 160
rect 3311 104 3397 160
rect 3453 104 3539 160
rect 3595 104 3681 160
rect 3737 104 3823 160
rect 3879 104 3965 160
rect 4021 104 4107 160
rect 4163 104 4249 160
rect 4305 104 4391 160
rect 4447 104 4533 160
rect 4589 104 4675 160
rect 4731 104 4817 160
rect 4873 104 4959 160
rect 5015 104 5101 160
rect 5157 104 5243 160
rect 5299 104 5385 160
rect 5441 104 5527 160
rect 5583 104 5669 160
rect 5725 104 5811 160
rect 5867 104 5953 160
rect 6009 104 6095 160
rect 6151 104 6237 160
rect 6293 104 6379 160
rect 6435 104 6521 160
rect 6577 104 6663 160
rect 6719 104 6805 160
rect 6861 104 6947 160
rect 7003 104 7089 160
rect 7145 104 7231 160
rect 7287 104 7373 160
rect 7429 104 7515 160
rect 7571 104 7657 160
rect 7713 104 7799 160
rect 7855 104 7941 160
rect 7997 104 8083 160
rect 8139 104 8225 160
rect 8281 104 8367 160
rect 8423 104 8509 160
rect 8565 104 8651 160
rect 8707 104 8793 160
rect 8849 104 8935 160
rect 8991 104 9077 160
rect 9133 104 9219 160
rect 9275 104 9361 160
rect 9417 104 9503 160
rect 9559 104 9645 160
rect 9701 104 9787 160
rect 9843 104 9929 160
rect 9985 104 10071 160
rect 10127 104 10213 160
rect 10269 104 10355 160
rect 10411 104 10497 160
rect 10553 104 10639 160
rect 10695 104 10781 160
rect 10837 104 10923 160
rect 10979 104 11065 160
rect 11121 104 11207 160
rect 11263 104 11349 160
rect 11405 104 11491 160
rect 11547 104 11633 160
rect 11689 104 11775 160
rect 11831 104 11917 160
rect 11973 104 12059 160
rect 12115 104 12201 160
rect 12257 104 12343 160
rect 12399 150 12526 160
rect 12582 150 12650 206
rect 12706 150 12774 206
rect 12830 150 12898 206
rect 12954 150 13022 206
rect 13078 150 13200 206
rect 12399 104 13200 150
rect -400 0 13200 104
<< via2 >>
rect -254 12893 -198 12949
rect -130 12893 -74 12949
rect -6 12893 50 12949
rect 118 12893 174 12949
rect 242 12893 298 12949
rect 366 12893 422 12949
rect 490 12893 546 12949
rect 614 12893 670 12949
rect 738 12893 794 12949
rect 862 12893 918 12949
rect 986 12893 1042 12949
rect 1110 12893 1166 12949
rect 1234 12893 1290 12949
rect 1358 12893 1414 12949
rect 1482 12893 1538 12949
rect 1606 12893 1662 12949
rect 1730 12893 1786 12949
rect 1854 12893 1910 12949
rect 1978 12893 2034 12949
rect 2102 12893 2158 12949
rect 2226 12893 2282 12949
rect 2350 12893 2406 12949
rect 2474 12893 2530 12949
rect 2598 12893 2654 12949
rect 2722 12893 2778 12949
rect 2846 12893 2902 12949
rect 2970 12893 3026 12949
rect 3094 12893 3150 12949
rect 3218 12893 3274 12949
rect 3342 12893 3398 12949
rect 3466 12893 3522 12949
rect 3590 12893 3646 12949
rect 3714 12893 3770 12949
rect 3838 12893 3894 12949
rect 3962 12893 4018 12949
rect 4086 12893 4142 12949
rect 4210 12893 4266 12949
rect 4334 12893 4390 12949
rect 4458 12893 4514 12949
rect 4582 12893 4638 12949
rect 4706 12893 4762 12949
rect 4830 12893 4886 12949
rect 4954 12893 5010 12949
rect 5078 12893 5134 12949
rect 5202 12893 5258 12949
rect 5326 12893 5382 12949
rect 5450 12893 5506 12949
rect 5574 12893 5630 12949
rect 5698 12893 5754 12949
rect 5822 12893 5878 12949
rect 5946 12893 6002 12949
rect 6070 12893 6126 12949
rect 6194 12893 6250 12949
rect 6318 12893 6374 12949
rect 6442 12893 6498 12949
rect 6566 12893 6622 12949
rect 6690 12893 6746 12949
rect 6814 12893 6870 12949
rect 6938 12893 6994 12949
rect 7062 12893 7118 12949
rect 7186 12893 7242 12949
rect 7310 12893 7366 12949
rect 7434 12893 7490 12949
rect 7558 12893 7614 12949
rect 7682 12893 7738 12949
rect 7806 12893 7862 12949
rect 7930 12893 7986 12949
rect 8054 12893 8110 12949
rect 8178 12893 8234 12949
rect 8302 12893 8358 12949
rect 8426 12893 8482 12949
rect 8550 12893 8606 12949
rect 8674 12893 8730 12949
rect 8798 12893 8854 12949
rect 8922 12893 8978 12949
rect 9046 12893 9102 12949
rect 9170 12893 9226 12949
rect 9294 12893 9350 12949
rect 9418 12893 9474 12949
rect 9542 12893 9598 12949
rect 9666 12893 9722 12949
rect 9790 12893 9846 12949
rect 9914 12893 9970 12949
rect 10038 12893 10094 12949
rect 10162 12893 10218 12949
rect 10286 12893 10342 12949
rect 10410 12893 10466 12949
rect 10534 12893 10590 12949
rect 10658 12893 10714 12949
rect 10782 12893 10838 12949
rect 10906 12893 10962 12949
rect 11030 12893 11086 12949
rect 11154 12893 11210 12949
rect 11278 12893 11334 12949
rect 11402 12893 11458 12949
rect 11526 12893 11582 12949
rect 11650 12893 11706 12949
rect 11774 12893 11830 12949
rect 11898 12893 11954 12949
rect 12022 12893 12078 12949
rect 12146 12893 12202 12949
rect 12270 12893 12326 12949
rect 12394 12893 12450 12949
rect 12518 12893 12574 12949
rect 12642 12893 12698 12949
rect 12766 12893 12822 12949
rect 12890 12893 12946 12949
rect 13014 12893 13070 12949
rect -254 12769 -198 12825
rect -130 12769 -74 12825
rect -6 12769 50 12825
rect 118 12769 174 12825
rect 242 12769 298 12825
rect 366 12769 422 12825
rect 490 12769 546 12825
rect 614 12769 670 12825
rect 738 12769 794 12825
rect 862 12769 918 12825
rect 986 12769 1042 12825
rect 1110 12769 1166 12825
rect 1234 12769 1290 12825
rect 1358 12769 1414 12825
rect 1482 12769 1538 12825
rect 1606 12769 1662 12825
rect 1730 12769 1786 12825
rect 1854 12769 1910 12825
rect 1978 12769 2034 12825
rect 2102 12769 2158 12825
rect 2226 12769 2282 12825
rect 2350 12769 2406 12825
rect 2474 12769 2530 12825
rect 2598 12769 2654 12825
rect 2722 12769 2778 12825
rect 2846 12769 2902 12825
rect 2970 12769 3026 12825
rect 3094 12769 3150 12825
rect 3218 12769 3274 12825
rect 3342 12769 3398 12825
rect 3466 12769 3522 12825
rect 3590 12769 3646 12825
rect 3714 12769 3770 12825
rect 3838 12769 3894 12825
rect 3962 12769 4018 12825
rect 4086 12769 4142 12825
rect 4210 12769 4266 12825
rect 4334 12769 4390 12825
rect 4458 12769 4514 12825
rect 4582 12769 4638 12825
rect 4706 12769 4762 12825
rect 4830 12769 4886 12825
rect 4954 12769 5010 12825
rect 5078 12769 5134 12825
rect 5202 12769 5258 12825
rect 5326 12769 5382 12825
rect 5450 12769 5506 12825
rect 5574 12769 5630 12825
rect 5698 12769 5754 12825
rect 5822 12769 5878 12825
rect 5946 12769 6002 12825
rect 6070 12769 6126 12825
rect 6194 12769 6250 12825
rect 6318 12769 6374 12825
rect 6442 12769 6498 12825
rect 6566 12769 6622 12825
rect 6690 12769 6746 12825
rect 6814 12769 6870 12825
rect 6938 12769 6994 12825
rect 7062 12769 7118 12825
rect 7186 12769 7242 12825
rect 7310 12769 7366 12825
rect 7434 12769 7490 12825
rect 7558 12769 7614 12825
rect 7682 12769 7738 12825
rect 7806 12769 7862 12825
rect 7930 12769 7986 12825
rect 8054 12769 8110 12825
rect 8178 12769 8234 12825
rect 8302 12769 8358 12825
rect 8426 12769 8482 12825
rect 8550 12769 8606 12825
rect 8674 12769 8730 12825
rect 8798 12769 8854 12825
rect 8922 12769 8978 12825
rect 9046 12769 9102 12825
rect 9170 12769 9226 12825
rect 9294 12769 9350 12825
rect 9418 12769 9474 12825
rect 9542 12769 9598 12825
rect 9666 12769 9722 12825
rect 9790 12769 9846 12825
rect 9914 12769 9970 12825
rect 10038 12769 10094 12825
rect 10162 12769 10218 12825
rect 10286 12769 10342 12825
rect 10410 12769 10466 12825
rect 10534 12769 10590 12825
rect 10658 12769 10714 12825
rect 10782 12769 10838 12825
rect 10906 12769 10962 12825
rect 11030 12769 11086 12825
rect 11154 12769 11210 12825
rect 11278 12769 11334 12825
rect 11402 12769 11458 12825
rect 11526 12769 11582 12825
rect 11650 12769 11706 12825
rect 11774 12769 11830 12825
rect 11898 12769 11954 12825
rect 12022 12769 12078 12825
rect 12146 12769 12202 12825
rect 12270 12769 12326 12825
rect 12394 12769 12450 12825
rect 12518 12769 12574 12825
rect 12642 12769 12698 12825
rect 12766 12769 12822 12825
rect 12890 12769 12946 12825
rect 13014 12769 13070 12825
rect -254 12645 -198 12701
rect -130 12645 -74 12701
rect -6 12645 50 12701
rect 118 12645 174 12701
rect 242 12645 298 12701
rect 366 12645 422 12701
rect 490 12645 546 12701
rect 614 12645 670 12701
rect 738 12645 794 12701
rect 862 12645 918 12701
rect 986 12645 1042 12701
rect 1110 12645 1166 12701
rect 1234 12645 1290 12701
rect 1358 12645 1414 12701
rect 1482 12645 1538 12701
rect 1606 12645 1662 12701
rect 1730 12645 1786 12701
rect 1854 12645 1910 12701
rect 1978 12645 2034 12701
rect 2102 12645 2158 12701
rect 2226 12645 2282 12701
rect 2350 12645 2406 12701
rect 2474 12645 2530 12701
rect 2598 12645 2654 12701
rect 2722 12645 2778 12701
rect 2846 12645 2902 12701
rect 2970 12645 3026 12701
rect 3094 12645 3150 12701
rect 3218 12645 3274 12701
rect 3342 12645 3398 12701
rect 3466 12645 3522 12701
rect 3590 12645 3646 12701
rect 3714 12645 3770 12701
rect 3838 12645 3894 12701
rect 3962 12645 4018 12701
rect 4086 12645 4142 12701
rect 4210 12645 4266 12701
rect 4334 12645 4390 12701
rect 4458 12645 4514 12701
rect 4582 12645 4638 12701
rect 4706 12645 4762 12701
rect 4830 12645 4886 12701
rect 4954 12645 5010 12701
rect 5078 12645 5134 12701
rect 5202 12645 5258 12701
rect 5326 12645 5382 12701
rect 5450 12645 5506 12701
rect 5574 12645 5630 12701
rect 5698 12645 5754 12701
rect 5822 12645 5878 12701
rect 5946 12645 6002 12701
rect 6070 12645 6126 12701
rect 6194 12645 6250 12701
rect 6318 12645 6374 12701
rect 6442 12645 6498 12701
rect 6566 12645 6622 12701
rect 6690 12645 6746 12701
rect 6814 12645 6870 12701
rect 6938 12645 6994 12701
rect 7062 12645 7118 12701
rect 7186 12645 7242 12701
rect 7310 12645 7366 12701
rect 7434 12645 7490 12701
rect 7558 12645 7614 12701
rect 7682 12645 7738 12701
rect 7806 12645 7862 12701
rect 7930 12645 7986 12701
rect 8054 12645 8110 12701
rect 8178 12645 8234 12701
rect 8302 12645 8358 12701
rect 8426 12645 8482 12701
rect 8550 12645 8606 12701
rect 8674 12645 8730 12701
rect 8798 12645 8854 12701
rect 8922 12645 8978 12701
rect 9046 12645 9102 12701
rect 9170 12645 9226 12701
rect 9294 12645 9350 12701
rect 9418 12645 9474 12701
rect 9542 12645 9598 12701
rect 9666 12645 9722 12701
rect 9790 12645 9846 12701
rect 9914 12645 9970 12701
rect 10038 12645 10094 12701
rect 10162 12645 10218 12701
rect 10286 12645 10342 12701
rect 10410 12645 10466 12701
rect 10534 12645 10590 12701
rect 10658 12645 10714 12701
rect 10782 12645 10838 12701
rect 10906 12645 10962 12701
rect 11030 12645 11086 12701
rect 11154 12645 11210 12701
rect 11278 12645 11334 12701
rect 11402 12645 11458 12701
rect 11526 12645 11582 12701
rect 11650 12645 11706 12701
rect 11774 12645 11830 12701
rect 11898 12645 11954 12701
rect 12022 12645 12078 12701
rect 12146 12645 12202 12701
rect 12270 12645 12326 12701
rect 12394 12645 12450 12701
rect 12518 12645 12574 12701
rect 12642 12645 12698 12701
rect 12766 12645 12822 12701
rect 12890 12645 12946 12701
rect 13014 12645 13070 12701
rect -254 12521 -198 12577
rect -130 12521 -74 12577
rect -6 12521 50 12577
rect 118 12521 174 12577
rect 242 12521 298 12577
rect 366 12521 422 12577
rect 490 12521 546 12577
rect 614 12521 670 12577
rect 738 12521 794 12577
rect 862 12521 918 12577
rect 986 12521 1042 12577
rect 1110 12521 1166 12577
rect 1234 12521 1290 12577
rect 1358 12521 1414 12577
rect 1482 12521 1538 12577
rect 1606 12521 1662 12577
rect 1730 12521 1786 12577
rect 1854 12521 1910 12577
rect 1978 12521 2034 12577
rect 2102 12521 2158 12577
rect 2226 12521 2282 12577
rect 2350 12521 2406 12577
rect 2474 12521 2530 12577
rect 2598 12521 2654 12577
rect 2722 12521 2778 12577
rect 2846 12521 2902 12577
rect 2970 12521 3026 12577
rect 3094 12521 3150 12577
rect 3218 12521 3274 12577
rect 3342 12521 3398 12577
rect 3466 12521 3522 12577
rect 3590 12521 3646 12577
rect 3714 12521 3770 12577
rect 3838 12521 3894 12577
rect 3962 12521 4018 12577
rect 4086 12521 4142 12577
rect 4210 12521 4266 12577
rect 4334 12521 4390 12577
rect 4458 12521 4514 12577
rect 4582 12521 4638 12577
rect 4706 12521 4762 12577
rect 4830 12521 4886 12577
rect 4954 12521 5010 12577
rect 5078 12521 5134 12577
rect 5202 12521 5258 12577
rect 5326 12521 5382 12577
rect 5450 12521 5506 12577
rect 5574 12521 5630 12577
rect 5698 12521 5754 12577
rect 5822 12521 5878 12577
rect 5946 12521 6002 12577
rect 6070 12521 6126 12577
rect 6194 12521 6250 12577
rect 6318 12521 6374 12577
rect 6442 12521 6498 12577
rect 6566 12521 6622 12577
rect 6690 12521 6746 12577
rect 6814 12521 6870 12577
rect 6938 12521 6994 12577
rect 7062 12521 7118 12577
rect 7186 12521 7242 12577
rect 7310 12521 7366 12577
rect 7434 12521 7490 12577
rect 7558 12521 7614 12577
rect 7682 12521 7738 12577
rect 7806 12521 7862 12577
rect 7930 12521 7986 12577
rect 8054 12521 8110 12577
rect 8178 12521 8234 12577
rect 8302 12521 8358 12577
rect 8426 12521 8482 12577
rect 8550 12521 8606 12577
rect 8674 12521 8730 12577
rect 8798 12521 8854 12577
rect 8922 12521 8978 12577
rect 9046 12521 9102 12577
rect 9170 12521 9226 12577
rect 9294 12521 9350 12577
rect 9418 12521 9474 12577
rect 9542 12521 9598 12577
rect 9666 12521 9722 12577
rect 9790 12521 9846 12577
rect 9914 12521 9970 12577
rect 10038 12521 10094 12577
rect 10162 12521 10218 12577
rect 10286 12521 10342 12577
rect 10410 12521 10466 12577
rect 10534 12521 10590 12577
rect 10658 12521 10714 12577
rect 10782 12521 10838 12577
rect 10906 12521 10962 12577
rect 11030 12521 11086 12577
rect 11154 12521 11210 12577
rect 11278 12521 11334 12577
rect 11402 12521 11458 12577
rect 11526 12521 11582 12577
rect 11650 12521 11706 12577
rect 11774 12521 11830 12577
rect 11898 12521 11954 12577
rect 12022 12521 12078 12577
rect 12146 12521 12202 12577
rect 12270 12521 12326 12577
rect 12394 12521 12450 12577
rect 12518 12521 12574 12577
rect 12642 12521 12698 12577
rect 12766 12521 12822 12577
rect 12890 12521 12946 12577
rect 13014 12521 13070 12577
rect -286 12302 -230 12358
rect -162 12302 -106 12358
rect -38 12302 18 12358
rect 86 12302 142 12358
rect 210 12302 266 12358
rect -286 12178 -230 12234
rect -162 12178 -106 12234
rect -38 12178 18 12234
rect 86 12178 142 12234
rect 210 12178 266 12234
rect -286 12054 -230 12110
rect -162 12054 -106 12110
rect -38 12054 18 12110
rect 86 12054 142 12110
rect 210 12054 266 12110
rect -286 11930 -230 11986
rect -162 11930 -106 11986
rect -38 11930 18 11986
rect 86 11930 142 11986
rect 210 11930 266 11986
rect -286 11806 -230 11862
rect -162 11806 -106 11862
rect -38 11806 18 11862
rect 86 11806 142 11862
rect 210 11806 266 11862
rect -286 11682 -230 11738
rect -162 11682 -106 11738
rect -38 11682 18 11738
rect 86 11682 142 11738
rect 210 11682 266 11738
rect -286 11558 -230 11614
rect -162 11558 -106 11614
rect -38 11558 18 11614
rect 86 11558 142 11614
rect 210 11558 266 11614
rect -286 11434 -230 11490
rect -162 11434 -106 11490
rect -38 11434 18 11490
rect 86 11434 142 11490
rect 210 11434 266 11490
rect -286 11310 -230 11366
rect -162 11310 -106 11366
rect -38 11310 18 11366
rect 86 11310 142 11366
rect 210 11310 266 11366
rect -286 11186 -230 11242
rect -162 11186 -106 11242
rect -38 11186 18 11242
rect 86 11186 142 11242
rect 210 11186 266 11242
rect -286 11062 -230 11118
rect -162 11062 -106 11118
rect -38 11062 18 11118
rect 86 11062 142 11118
rect 210 11062 266 11118
rect -286 10938 -230 10994
rect -162 10938 -106 10994
rect -38 10938 18 10994
rect 86 10938 142 10994
rect 210 10938 266 10994
rect -286 10814 -230 10870
rect -162 10814 -106 10870
rect -38 10814 18 10870
rect 86 10814 142 10870
rect 210 10814 266 10870
rect -286 10690 -230 10746
rect -162 10690 -106 10746
rect -38 10690 18 10746
rect 86 10690 142 10746
rect 210 10690 266 10746
rect -286 10566 -230 10622
rect -162 10566 -106 10622
rect -38 10566 18 10622
rect 86 10566 142 10622
rect 210 10566 266 10622
rect -286 10442 -230 10498
rect -162 10442 -106 10498
rect -38 10442 18 10498
rect 86 10442 142 10498
rect 210 10442 266 10498
rect -286 10318 -230 10374
rect -162 10318 -106 10374
rect -38 10318 18 10374
rect 86 10318 142 10374
rect 210 10318 266 10374
rect -286 10194 -230 10250
rect -162 10194 -106 10250
rect -38 10194 18 10250
rect 86 10194 142 10250
rect 210 10194 266 10250
rect -286 10070 -230 10126
rect -162 10070 -106 10126
rect -38 10070 18 10126
rect 86 10070 142 10126
rect 210 10070 266 10126
rect -286 9946 -230 10002
rect -162 9946 -106 10002
rect -38 9946 18 10002
rect 86 9946 142 10002
rect 210 9946 266 10002
rect -286 9822 -230 9878
rect -162 9822 -106 9878
rect -38 9822 18 9878
rect 86 9822 142 9878
rect 210 9822 266 9878
rect -286 9698 -230 9754
rect -162 9698 -106 9754
rect -38 9698 18 9754
rect 86 9698 142 9754
rect 210 9698 266 9754
rect -286 9574 -230 9630
rect -162 9574 -106 9630
rect -38 9574 18 9630
rect 86 9574 142 9630
rect 210 9574 266 9630
rect -286 9450 -230 9506
rect -162 9450 -106 9506
rect -38 9450 18 9506
rect 86 9450 142 9506
rect 210 9450 266 9506
rect -286 9326 -230 9382
rect -162 9326 -106 9382
rect -38 9326 18 9382
rect 86 9326 142 9382
rect 210 9326 266 9382
rect -286 9202 -230 9258
rect -162 9202 -106 9258
rect -38 9202 18 9258
rect 86 9202 142 9258
rect 210 9202 266 9258
rect -286 9078 -230 9134
rect -162 9078 -106 9134
rect -38 9078 18 9134
rect 86 9078 142 9134
rect 210 9078 266 9134
rect -286 8954 -230 9010
rect -162 8954 -106 9010
rect -38 8954 18 9010
rect 86 8954 142 9010
rect 210 8954 266 9010
rect -286 8830 -230 8886
rect -162 8830 -106 8886
rect -38 8830 18 8886
rect 86 8830 142 8886
rect 210 8830 266 8886
rect -286 8706 -230 8762
rect -162 8706 -106 8762
rect -38 8706 18 8762
rect 86 8706 142 8762
rect 210 8706 266 8762
rect -286 8582 -230 8638
rect -162 8582 -106 8638
rect -38 8582 18 8638
rect 86 8582 142 8638
rect 210 8582 266 8638
rect -286 8458 -230 8514
rect -162 8458 -106 8514
rect -38 8458 18 8514
rect 86 8458 142 8514
rect 210 8458 266 8514
rect -286 8334 -230 8390
rect -162 8334 -106 8390
rect -38 8334 18 8390
rect 86 8334 142 8390
rect 210 8334 266 8390
rect -286 8210 -230 8266
rect -162 8210 -106 8266
rect -38 8210 18 8266
rect 86 8210 142 8266
rect 210 8210 266 8266
rect -286 8086 -230 8142
rect -162 8086 -106 8142
rect -38 8086 18 8142
rect 86 8086 142 8142
rect 210 8086 266 8142
rect -286 7962 -230 8018
rect -162 7962 -106 8018
rect -38 7962 18 8018
rect 86 7962 142 8018
rect 210 7962 266 8018
rect -286 7838 -230 7894
rect -162 7838 -106 7894
rect -38 7838 18 7894
rect 86 7838 142 7894
rect 210 7838 266 7894
rect -286 7714 -230 7770
rect -162 7714 -106 7770
rect -38 7714 18 7770
rect 86 7714 142 7770
rect 210 7714 266 7770
rect -286 7590 -230 7646
rect -162 7590 -106 7646
rect -38 7590 18 7646
rect 86 7590 142 7646
rect 210 7590 266 7646
rect -286 7466 -230 7522
rect -162 7466 -106 7522
rect -38 7466 18 7522
rect 86 7466 142 7522
rect 210 7466 266 7522
rect -286 7342 -230 7398
rect -162 7342 -106 7398
rect -38 7342 18 7398
rect 86 7342 142 7398
rect 210 7342 266 7398
rect -286 7218 -230 7274
rect -162 7218 -106 7274
rect -38 7218 18 7274
rect 86 7218 142 7274
rect 210 7218 266 7274
rect -286 7094 -230 7150
rect -162 7094 -106 7150
rect -38 7094 18 7150
rect 86 7094 142 7150
rect 210 7094 266 7150
rect -286 6970 -230 7026
rect -162 6970 -106 7026
rect -38 6970 18 7026
rect 86 6970 142 7026
rect 210 6970 266 7026
rect -286 6846 -230 6902
rect -162 6846 -106 6902
rect -38 6846 18 6902
rect 86 6846 142 6902
rect 210 6846 266 6902
rect -286 6722 -230 6778
rect -162 6722 -106 6778
rect -38 6722 18 6778
rect 86 6722 142 6778
rect 210 6722 266 6778
rect -286 6598 -230 6654
rect -162 6598 -106 6654
rect -38 6598 18 6654
rect 86 6598 142 6654
rect 210 6598 266 6654
rect -286 6474 -230 6530
rect -162 6474 -106 6530
rect -38 6474 18 6530
rect 86 6474 142 6530
rect 210 6474 266 6530
rect -286 6350 -230 6406
rect -162 6350 -106 6406
rect -38 6350 18 6406
rect 86 6350 142 6406
rect 210 6350 266 6406
rect -286 6226 -230 6282
rect -162 6226 -106 6282
rect -38 6226 18 6282
rect 86 6226 142 6282
rect 210 6226 266 6282
rect -286 6102 -230 6158
rect -162 6102 -106 6158
rect -38 6102 18 6158
rect 86 6102 142 6158
rect 210 6102 266 6158
rect -286 5978 -230 6034
rect -162 5978 -106 6034
rect -38 5978 18 6034
rect 86 5978 142 6034
rect 210 5978 266 6034
rect -286 5854 -230 5910
rect -162 5854 -106 5910
rect -38 5854 18 5910
rect 86 5854 142 5910
rect 210 5854 266 5910
rect -286 5730 -230 5786
rect -162 5730 -106 5786
rect -38 5730 18 5786
rect 86 5730 142 5786
rect 210 5730 266 5786
rect -286 5606 -230 5662
rect -162 5606 -106 5662
rect -38 5606 18 5662
rect 86 5606 142 5662
rect 210 5606 266 5662
rect -286 5482 -230 5538
rect -162 5482 -106 5538
rect -38 5482 18 5538
rect 86 5482 142 5538
rect 210 5482 266 5538
rect -286 5358 -230 5414
rect -162 5358 -106 5414
rect -38 5358 18 5414
rect 86 5358 142 5414
rect 210 5358 266 5414
rect -286 5234 -230 5290
rect -162 5234 -106 5290
rect -38 5234 18 5290
rect 86 5234 142 5290
rect 210 5234 266 5290
rect -286 5110 -230 5166
rect -162 5110 -106 5166
rect -38 5110 18 5166
rect 86 5110 142 5166
rect 210 5110 266 5166
rect -286 4986 -230 5042
rect -162 4986 -106 5042
rect -38 4986 18 5042
rect 86 4986 142 5042
rect 210 4986 266 5042
rect -286 4862 -230 4918
rect -162 4862 -106 4918
rect -38 4862 18 4918
rect 86 4862 142 4918
rect 210 4862 266 4918
rect -286 4738 -230 4794
rect -162 4738 -106 4794
rect -38 4738 18 4794
rect 86 4738 142 4794
rect 210 4738 266 4794
rect -286 4614 -230 4670
rect -162 4614 -106 4670
rect -38 4614 18 4670
rect 86 4614 142 4670
rect 210 4614 266 4670
rect -286 4490 -230 4546
rect -162 4490 -106 4546
rect -38 4490 18 4546
rect 86 4490 142 4546
rect 210 4490 266 4546
rect -286 4366 -230 4422
rect -162 4366 -106 4422
rect -38 4366 18 4422
rect 86 4366 142 4422
rect 210 4366 266 4422
rect -286 4242 -230 4298
rect -162 4242 -106 4298
rect -38 4242 18 4298
rect 86 4242 142 4298
rect 210 4242 266 4298
rect -286 4118 -230 4174
rect -162 4118 -106 4174
rect -38 4118 18 4174
rect 86 4118 142 4174
rect 210 4118 266 4174
rect -286 3994 -230 4050
rect -162 3994 -106 4050
rect -38 3994 18 4050
rect 86 3994 142 4050
rect 210 3994 266 4050
rect -286 3870 -230 3926
rect -162 3870 -106 3926
rect -38 3870 18 3926
rect 86 3870 142 3926
rect 210 3870 266 3926
rect -286 3746 -230 3802
rect -162 3746 -106 3802
rect -38 3746 18 3802
rect 86 3746 142 3802
rect 210 3746 266 3802
rect -286 3622 -230 3678
rect -162 3622 -106 3678
rect -38 3622 18 3678
rect 86 3622 142 3678
rect 210 3622 266 3678
rect -286 3498 -230 3554
rect -162 3498 -106 3554
rect -38 3498 18 3554
rect 86 3498 142 3554
rect 210 3498 266 3554
rect -286 3374 -230 3430
rect -162 3374 -106 3430
rect -38 3374 18 3430
rect 86 3374 142 3430
rect 210 3374 266 3430
rect -286 3250 -230 3306
rect -162 3250 -106 3306
rect -38 3250 18 3306
rect 86 3250 142 3306
rect 210 3250 266 3306
rect -286 3126 -230 3182
rect -162 3126 -106 3182
rect -38 3126 18 3182
rect 86 3126 142 3182
rect 210 3126 266 3182
rect -286 3002 -230 3058
rect -162 3002 -106 3058
rect -38 3002 18 3058
rect 86 3002 142 3058
rect 210 3002 266 3058
rect -286 2878 -230 2934
rect -162 2878 -106 2934
rect -38 2878 18 2934
rect 86 2878 142 2934
rect 210 2878 266 2934
rect -286 2754 -230 2810
rect -162 2754 -106 2810
rect -38 2754 18 2810
rect 86 2754 142 2810
rect 210 2754 266 2810
rect -286 2630 -230 2686
rect -162 2630 -106 2686
rect -38 2630 18 2686
rect 86 2630 142 2686
rect 210 2630 266 2686
rect -286 2506 -230 2562
rect -162 2506 -106 2562
rect -38 2506 18 2562
rect 86 2506 142 2562
rect 210 2506 266 2562
rect -286 2382 -230 2438
rect -162 2382 -106 2438
rect -38 2382 18 2438
rect 86 2382 142 2438
rect 210 2382 266 2438
rect -286 2258 -230 2314
rect -162 2258 -106 2314
rect -38 2258 18 2314
rect 86 2258 142 2314
rect 210 2258 266 2314
rect -286 2134 -230 2190
rect -162 2134 -106 2190
rect -38 2134 18 2190
rect 86 2134 142 2190
rect 210 2134 266 2190
rect -286 2010 -230 2066
rect -162 2010 -106 2066
rect -38 2010 18 2066
rect 86 2010 142 2066
rect 210 2010 266 2066
rect -286 1886 -230 1942
rect -162 1886 -106 1942
rect -38 1886 18 1942
rect 86 1886 142 1942
rect 210 1886 266 1942
rect -286 1762 -230 1818
rect -162 1762 -106 1818
rect -38 1762 18 1818
rect 86 1762 142 1818
rect 210 1762 266 1818
rect -286 1638 -230 1694
rect -162 1638 -106 1694
rect -38 1638 18 1694
rect 86 1638 142 1694
rect 210 1638 266 1694
rect -286 1514 -230 1570
rect -162 1514 -106 1570
rect -38 1514 18 1570
rect 86 1514 142 1570
rect 210 1514 266 1570
rect -286 1390 -230 1446
rect -162 1390 -106 1446
rect -38 1390 18 1446
rect 86 1390 142 1446
rect 210 1390 266 1446
rect -286 1266 -230 1322
rect -162 1266 -106 1322
rect -38 1266 18 1322
rect 86 1266 142 1322
rect 210 1266 266 1322
rect -286 1142 -230 1198
rect -162 1142 -106 1198
rect -38 1142 18 1198
rect 86 1142 142 1198
rect 210 1142 266 1198
rect -286 1018 -230 1074
rect -162 1018 -106 1074
rect -38 1018 18 1074
rect 86 1018 142 1074
rect 210 1018 266 1074
rect -286 894 -230 950
rect -162 894 -106 950
rect -38 894 18 950
rect 86 894 142 950
rect 210 894 266 950
rect -286 770 -230 826
rect -162 770 -106 826
rect -38 770 18 826
rect 86 770 142 826
rect 210 770 266 826
rect -286 646 -230 702
rect -162 646 -106 702
rect -38 646 18 702
rect 86 646 142 702
rect 210 646 266 702
rect -286 522 -230 578
rect -162 522 -106 578
rect -38 522 18 578
rect 86 522 142 578
rect 210 522 266 578
rect -286 398 -230 454
rect -162 398 -106 454
rect -38 398 18 454
rect 86 398 142 454
rect 210 398 266 454
rect 741 12254 797 12310
rect 883 12254 939 12310
rect 741 12112 797 12168
rect 883 12112 939 12168
rect 741 11970 797 12026
rect 883 11970 939 12026
rect 741 11828 797 11884
rect 883 11828 939 11884
rect 741 11686 797 11742
rect 883 11686 939 11742
rect 741 11544 797 11600
rect 883 11544 939 11600
rect 741 11402 797 11458
rect 883 11402 939 11458
rect 741 11260 797 11316
rect 883 11260 939 11316
rect 741 11118 797 11174
rect 883 11118 939 11174
rect 741 10976 797 11032
rect 883 10976 939 11032
rect 741 10834 797 10890
rect 883 10834 939 10890
rect 741 10692 797 10748
rect 883 10692 939 10748
rect 741 10550 797 10606
rect 883 10550 939 10606
rect 741 10408 797 10464
rect 883 10408 939 10464
rect 741 10266 797 10322
rect 883 10266 939 10322
rect 741 10124 797 10180
rect 883 10124 939 10180
rect 741 9982 797 10038
rect 883 9982 939 10038
rect 741 9840 797 9896
rect 883 9840 939 9896
rect 741 9698 797 9754
rect 883 9698 939 9754
rect 741 9556 797 9612
rect 883 9556 939 9612
rect 741 9414 797 9470
rect 883 9414 939 9470
rect 741 9272 797 9328
rect 883 9272 939 9328
rect 741 9130 797 9186
rect 883 9130 939 9186
rect 741 8988 797 9044
rect 883 8988 939 9044
rect 741 8846 797 8902
rect 883 8846 939 8902
rect 741 8704 797 8760
rect 883 8704 939 8760
rect 741 8562 797 8618
rect 883 8562 939 8618
rect 741 8420 797 8476
rect 883 8420 939 8476
rect 741 8278 797 8334
rect 883 8278 939 8334
rect 741 8136 797 8192
rect 883 8136 939 8192
rect 741 7994 797 8050
rect 883 7994 939 8050
rect 741 7852 797 7908
rect 883 7852 939 7908
rect 741 7710 797 7766
rect 883 7710 939 7766
rect 741 7568 797 7624
rect 883 7568 939 7624
rect 741 7426 797 7482
rect 883 7426 939 7482
rect 741 7284 797 7340
rect 883 7284 939 7340
rect 741 7142 797 7198
rect 883 7142 939 7198
rect 741 7000 797 7056
rect 883 7000 939 7056
rect 741 6858 797 6914
rect 883 6858 939 6914
rect 741 6716 797 6772
rect 883 6716 939 6772
rect 741 6574 797 6630
rect 883 6574 939 6630
rect 741 6432 797 6488
rect 883 6432 939 6488
rect 741 6290 797 6346
rect 883 6290 939 6346
rect 741 6148 797 6204
rect 883 6148 939 6204
rect 741 6006 797 6062
rect 883 6006 939 6062
rect 741 5864 797 5920
rect 883 5864 939 5920
rect 741 5722 797 5778
rect 883 5722 939 5778
rect 741 5580 797 5636
rect 883 5580 939 5636
rect 741 5438 797 5494
rect 883 5438 939 5494
rect 741 5296 797 5352
rect 883 5296 939 5352
rect 741 5154 797 5210
rect 883 5154 939 5210
rect 741 5012 797 5068
rect 883 5012 939 5068
rect 741 4870 797 4926
rect 883 4870 939 4926
rect 741 4728 797 4784
rect 883 4728 939 4784
rect 741 4586 797 4642
rect 883 4586 939 4642
rect 741 4444 797 4500
rect 883 4444 939 4500
rect 741 4302 797 4358
rect 883 4302 939 4358
rect 741 4160 797 4216
rect 883 4160 939 4216
rect 741 4018 797 4074
rect 883 4018 939 4074
rect 741 3876 797 3932
rect 883 3876 939 3932
rect 741 3734 797 3790
rect 883 3734 939 3790
rect 741 3592 797 3648
rect 883 3592 939 3648
rect 741 3450 797 3506
rect 883 3450 939 3506
rect 741 3308 797 3364
rect 883 3308 939 3364
rect 741 3166 797 3222
rect 883 3166 939 3222
rect 741 3024 797 3080
rect 883 3024 939 3080
rect 741 2882 797 2938
rect 883 2882 939 2938
rect 741 2740 797 2796
rect 883 2740 939 2796
rect 741 2598 797 2654
rect 883 2598 939 2654
rect 741 2456 797 2512
rect 883 2456 939 2512
rect 741 2314 797 2370
rect 883 2314 939 2370
rect 741 2172 797 2228
rect 883 2172 939 2228
rect 741 2030 797 2086
rect 883 2030 939 2086
rect 741 1888 797 1944
rect 883 1888 939 1944
rect 741 1746 797 1802
rect 883 1746 939 1802
rect 741 1604 797 1660
rect 883 1604 939 1660
rect 741 1462 797 1518
rect 883 1462 939 1518
rect 741 1320 797 1376
rect 883 1320 939 1376
rect 741 1178 797 1234
rect 883 1178 939 1234
rect 741 1036 797 1092
rect 883 1036 939 1092
rect 741 894 797 950
rect 883 894 939 950
rect 741 752 797 808
rect 883 752 939 808
rect 741 610 797 666
rect 883 610 939 666
rect 741 468 797 524
rect 883 468 939 524
rect 1142 12254 1198 12310
rect 1284 12254 1340 12310
rect 1142 12112 1198 12168
rect 1284 12112 1340 12168
rect 1142 11970 1198 12026
rect 1284 11970 1340 12026
rect 1142 11828 1198 11884
rect 1284 11828 1340 11884
rect 1142 11686 1198 11742
rect 1284 11686 1340 11742
rect 1142 11544 1198 11600
rect 1284 11544 1340 11600
rect 1142 11402 1198 11458
rect 1284 11402 1340 11458
rect 1142 11260 1198 11316
rect 1284 11260 1340 11316
rect 1142 11118 1198 11174
rect 1284 11118 1340 11174
rect 1142 10976 1198 11032
rect 1284 10976 1340 11032
rect 1142 10834 1198 10890
rect 1284 10834 1340 10890
rect 1142 10692 1198 10748
rect 1284 10692 1340 10748
rect 1142 10550 1198 10606
rect 1284 10550 1340 10606
rect 1142 10408 1198 10464
rect 1284 10408 1340 10464
rect 1142 10266 1198 10322
rect 1284 10266 1340 10322
rect 1142 10124 1198 10180
rect 1284 10124 1340 10180
rect 1142 9982 1198 10038
rect 1284 9982 1340 10038
rect 1142 9840 1198 9896
rect 1284 9840 1340 9896
rect 1142 9698 1198 9754
rect 1284 9698 1340 9754
rect 1142 9556 1198 9612
rect 1284 9556 1340 9612
rect 1142 9414 1198 9470
rect 1284 9414 1340 9470
rect 1142 9272 1198 9328
rect 1284 9272 1340 9328
rect 1142 9130 1198 9186
rect 1284 9130 1340 9186
rect 1142 8988 1198 9044
rect 1284 8988 1340 9044
rect 1142 8846 1198 8902
rect 1284 8846 1340 8902
rect 1142 8704 1198 8760
rect 1284 8704 1340 8760
rect 1142 8562 1198 8618
rect 1284 8562 1340 8618
rect 1142 8420 1198 8476
rect 1284 8420 1340 8476
rect 1142 8278 1198 8334
rect 1284 8278 1340 8334
rect 1142 8136 1198 8192
rect 1284 8136 1340 8192
rect 1142 7994 1198 8050
rect 1284 7994 1340 8050
rect 1142 7852 1198 7908
rect 1284 7852 1340 7908
rect 1142 7710 1198 7766
rect 1284 7710 1340 7766
rect 1142 7568 1198 7624
rect 1284 7568 1340 7624
rect 1142 7426 1198 7482
rect 1284 7426 1340 7482
rect 1142 7284 1198 7340
rect 1284 7284 1340 7340
rect 1142 7142 1198 7198
rect 1284 7142 1340 7198
rect 1142 7000 1198 7056
rect 1284 7000 1340 7056
rect 1142 6858 1198 6914
rect 1284 6858 1340 6914
rect 1142 6716 1198 6772
rect 1284 6716 1340 6772
rect 1142 6574 1198 6630
rect 1284 6574 1340 6630
rect 1142 6432 1198 6488
rect 1284 6432 1340 6488
rect 1142 6290 1198 6346
rect 1284 6290 1340 6346
rect 1142 6148 1198 6204
rect 1284 6148 1340 6204
rect 1142 6006 1198 6062
rect 1284 6006 1340 6062
rect 1142 5864 1198 5920
rect 1284 5864 1340 5920
rect 1142 5722 1198 5778
rect 1284 5722 1340 5778
rect 1142 5580 1198 5636
rect 1284 5580 1340 5636
rect 1142 5438 1198 5494
rect 1284 5438 1340 5494
rect 1142 5296 1198 5352
rect 1284 5296 1340 5352
rect 1142 5154 1198 5210
rect 1284 5154 1340 5210
rect 1142 5012 1198 5068
rect 1284 5012 1340 5068
rect 1142 4870 1198 4926
rect 1284 4870 1340 4926
rect 1142 4728 1198 4784
rect 1284 4728 1340 4784
rect 1142 4586 1198 4642
rect 1284 4586 1340 4642
rect 1142 4444 1198 4500
rect 1284 4444 1340 4500
rect 1142 4302 1198 4358
rect 1284 4302 1340 4358
rect 1142 4160 1198 4216
rect 1284 4160 1340 4216
rect 1142 4018 1198 4074
rect 1284 4018 1340 4074
rect 1142 3876 1198 3932
rect 1284 3876 1340 3932
rect 1142 3734 1198 3790
rect 1284 3734 1340 3790
rect 1142 3592 1198 3648
rect 1284 3592 1340 3648
rect 1142 3450 1198 3506
rect 1284 3450 1340 3506
rect 1142 3308 1198 3364
rect 1284 3308 1340 3364
rect 1142 3166 1198 3222
rect 1284 3166 1340 3222
rect 1142 3024 1198 3080
rect 1284 3024 1340 3080
rect 1142 2882 1198 2938
rect 1284 2882 1340 2938
rect 1142 2740 1198 2796
rect 1284 2740 1340 2796
rect 1142 2598 1198 2654
rect 1284 2598 1340 2654
rect 1142 2456 1198 2512
rect 1284 2456 1340 2512
rect 1142 2314 1198 2370
rect 1284 2314 1340 2370
rect 1142 2172 1198 2228
rect 1284 2172 1340 2228
rect 1142 2030 1198 2086
rect 1284 2030 1340 2086
rect 1142 1888 1198 1944
rect 1284 1888 1340 1944
rect 1142 1746 1198 1802
rect 1284 1746 1340 1802
rect 1142 1604 1198 1660
rect 1284 1604 1340 1660
rect 1142 1462 1198 1518
rect 1284 1462 1340 1518
rect 1142 1320 1198 1376
rect 1284 1320 1340 1376
rect 1142 1178 1198 1234
rect 1284 1178 1340 1234
rect 1142 1036 1198 1092
rect 1284 1036 1340 1092
rect 1142 894 1198 950
rect 1284 894 1340 950
rect 1142 752 1198 808
rect 1284 752 1340 808
rect 1142 610 1198 666
rect 1284 610 1340 666
rect 1142 468 1198 524
rect 1284 468 1340 524
rect 1542 12254 1598 12310
rect 1684 12254 1740 12310
rect 1542 12112 1598 12168
rect 1684 12112 1740 12168
rect 1542 11970 1598 12026
rect 1684 11970 1740 12026
rect 1542 11828 1598 11884
rect 1684 11828 1740 11884
rect 1542 11686 1598 11742
rect 1684 11686 1740 11742
rect 1542 11544 1598 11600
rect 1684 11544 1740 11600
rect 1542 11402 1598 11458
rect 1684 11402 1740 11458
rect 1542 11260 1598 11316
rect 1684 11260 1740 11316
rect 1542 11118 1598 11174
rect 1684 11118 1740 11174
rect 1542 10976 1598 11032
rect 1684 10976 1740 11032
rect 1542 10834 1598 10890
rect 1684 10834 1740 10890
rect 1542 10692 1598 10748
rect 1684 10692 1740 10748
rect 1542 10550 1598 10606
rect 1684 10550 1740 10606
rect 1542 10408 1598 10464
rect 1684 10408 1740 10464
rect 1542 10266 1598 10322
rect 1684 10266 1740 10322
rect 1542 10124 1598 10180
rect 1684 10124 1740 10180
rect 1542 9982 1598 10038
rect 1684 9982 1740 10038
rect 1542 9840 1598 9896
rect 1684 9840 1740 9896
rect 1542 9698 1598 9754
rect 1684 9698 1740 9754
rect 1542 9556 1598 9612
rect 1684 9556 1740 9612
rect 1542 9414 1598 9470
rect 1684 9414 1740 9470
rect 1542 9272 1598 9328
rect 1684 9272 1740 9328
rect 1542 9130 1598 9186
rect 1684 9130 1740 9186
rect 1542 8988 1598 9044
rect 1684 8988 1740 9044
rect 1542 8846 1598 8902
rect 1684 8846 1740 8902
rect 1542 8704 1598 8760
rect 1684 8704 1740 8760
rect 1542 8562 1598 8618
rect 1684 8562 1740 8618
rect 1542 8420 1598 8476
rect 1684 8420 1740 8476
rect 1542 8278 1598 8334
rect 1684 8278 1740 8334
rect 1542 8136 1598 8192
rect 1684 8136 1740 8192
rect 1542 7994 1598 8050
rect 1684 7994 1740 8050
rect 1542 7852 1598 7908
rect 1684 7852 1740 7908
rect 1542 7710 1598 7766
rect 1684 7710 1740 7766
rect 1542 7568 1598 7624
rect 1684 7568 1740 7624
rect 1542 7426 1598 7482
rect 1684 7426 1740 7482
rect 1542 7284 1598 7340
rect 1684 7284 1740 7340
rect 1542 7142 1598 7198
rect 1684 7142 1740 7198
rect 1542 7000 1598 7056
rect 1684 7000 1740 7056
rect 1542 6858 1598 6914
rect 1684 6858 1740 6914
rect 1542 6716 1598 6772
rect 1684 6716 1740 6772
rect 1542 6574 1598 6630
rect 1684 6574 1740 6630
rect 1542 6432 1598 6488
rect 1684 6432 1740 6488
rect 1542 6290 1598 6346
rect 1684 6290 1740 6346
rect 1542 6148 1598 6204
rect 1684 6148 1740 6204
rect 1542 6006 1598 6062
rect 1684 6006 1740 6062
rect 1542 5864 1598 5920
rect 1684 5864 1740 5920
rect 1542 5722 1598 5778
rect 1684 5722 1740 5778
rect 1542 5580 1598 5636
rect 1684 5580 1740 5636
rect 1542 5438 1598 5494
rect 1684 5438 1740 5494
rect 1542 5296 1598 5352
rect 1684 5296 1740 5352
rect 1542 5154 1598 5210
rect 1684 5154 1740 5210
rect 1542 5012 1598 5068
rect 1684 5012 1740 5068
rect 1542 4870 1598 4926
rect 1684 4870 1740 4926
rect 1542 4728 1598 4784
rect 1684 4728 1740 4784
rect 1542 4586 1598 4642
rect 1684 4586 1740 4642
rect 1542 4444 1598 4500
rect 1684 4444 1740 4500
rect 1542 4302 1598 4358
rect 1684 4302 1740 4358
rect 1542 4160 1598 4216
rect 1684 4160 1740 4216
rect 1542 4018 1598 4074
rect 1684 4018 1740 4074
rect 1542 3876 1598 3932
rect 1684 3876 1740 3932
rect 1542 3734 1598 3790
rect 1684 3734 1740 3790
rect 1542 3592 1598 3648
rect 1684 3592 1740 3648
rect 1542 3450 1598 3506
rect 1684 3450 1740 3506
rect 1542 3308 1598 3364
rect 1684 3308 1740 3364
rect 1542 3166 1598 3222
rect 1684 3166 1740 3222
rect 1542 3024 1598 3080
rect 1684 3024 1740 3080
rect 1542 2882 1598 2938
rect 1684 2882 1740 2938
rect 1542 2740 1598 2796
rect 1684 2740 1740 2796
rect 1542 2598 1598 2654
rect 1684 2598 1740 2654
rect 1542 2456 1598 2512
rect 1684 2456 1740 2512
rect 1542 2314 1598 2370
rect 1684 2314 1740 2370
rect 1542 2172 1598 2228
rect 1684 2172 1740 2228
rect 1542 2030 1598 2086
rect 1684 2030 1740 2086
rect 1542 1888 1598 1944
rect 1684 1888 1740 1944
rect 1542 1746 1598 1802
rect 1684 1746 1740 1802
rect 1542 1604 1598 1660
rect 1684 1604 1740 1660
rect 1542 1462 1598 1518
rect 1684 1462 1740 1518
rect 1542 1320 1598 1376
rect 1684 1320 1740 1376
rect 1542 1178 1598 1234
rect 1684 1178 1740 1234
rect 1542 1036 1598 1092
rect 1684 1036 1740 1092
rect 1542 894 1598 950
rect 1684 894 1740 950
rect 1542 752 1598 808
rect 1684 752 1740 808
rect 1542 610 1598 666
rect 1684 610 1740 666
rect 1542 468 1598 524
rect 1684 468 1740 524
rect 1939 12254 1995 12310
rect 2081 12254 2137 12310
rect 1939 12112 1995 12168
rect 2081 12112 2137 12168
rect 1939 11970 1995 12026
rect 2081 11970 2137 12026
rect 1939 11828 1995 11884
rect 2081 11828 2137 11884
rect 1939 11686 1995 11742
rect 2081 11686 2137 11742
rect 1939 11544 1995 11600
rect 2081 11544 2137 11600
rect 1939 11402 1995 11458
rect 2081 11402 2137 11458
rect 1939 11260 1995 11316
rect 2081 11260 2137 11316
rect 1939 11118 1995 11174
rect 2081 11118 2137 11174
rect 1939 10976 1995 11032
rect 2081 10976 2137 11032
rect 1939 10834 1995 10890
rect 2081 10834 2137 10890
rect 1939 10692 1995 10748
rect 2081 10692 2137 10748
rect 1939 10550 1995 10606
rect 2081 10550 2137 10606
rect 1939 10408 1995 10464
rect 2081 10408 2137 10464
rect 1939 10266 1995 10322
rect 2081 10266 2137 10322
rect 1939 10124 1995 10180
rect 2081 10124 2137 10180
rect 1939 9982 1995 10038
rect 2081 9982 2137 10038
rect 1939 9840 1995 9896
rect 2081 9840 2137 9896
rect 1939 9698 1995 9754
rect 2081 9698 2137 9754
rect 1939 9556 1995 9612
rect 2081 9556 2137 9612
rect 1939 9414 1995 9470
rect 2081 9414 2137 9470
rect 1939 9272 1995 9328
rect 2081 9272 2137 9328
rect 1939 9130 1995 9186
rect 2081 9130 2137 9186
rect 1939 8988 1995 9044
rect 2081 8988 2137 9044
rect 1939 8846 1995 8902
rect 2081 8846 2137 8902
rect 1939 8704 1995 8760
rect 2081 8704 2137 8760
rect 1939 8562 1995 8618
rect 2081 8562 2137 8618
rect 1939 8420 1995 8476
rect 2081 8420 2137 8476
rect 1939 8278 1995 8334
rect 2081 8278 2137 8334
rect 1939 8136 1995 8192
rect 2081 8136 2137 8192
rect 1939 7994 1995 8050
rect 2081 7994 2137 8050
rect 1939 7852 1995 7908
rect 2081 7852 2137 7908
rect 1939 7710 1995 7766
rect 2081 7710 2137 7766
rect 1939 7568 1995 7624
rect 2081 7568 2137 7624
rect 1939 7426 1995 7482
rect 2081 7426 2137 7482
rect 1939 7284 1995 7340
rect 2081 7284 2137 7340
rect 1939 7142 1995 7198
rect 2081 7142 2137 7198
rect 1939 7000 1995 7056
rect 2081 7000 2137 7056
rect 1939 6858 1995 6914
rect 2081 6858 2137 6914
rect 1939 6716 1995 6772
rect 2081 6716 2137 6772
rect 1939 6574 1995 6630
rect 2081 6574 2137 6630
rect 1939 6432 1995 6488
rect 2081 6432 2137 6488
rect 1939 6290 1995 6346
rect 2081 6290 2137 6346
rect 1939 6148 1995 6204
rect 2081 6148 2137 6204
rect 1939 6006 1995 6062
rect 2081 6006 2137 6062
rect 1939 5864 1995 5920
rect 2081 5864 2137 5920
rect 1939 5722 1995 5778
rect 2081 5722 2137 5778
rect 1939 5580 1995 5636
rect 2081 5580 2137 5636
rect 1939 5438 1995 5494
rect 2081 5438 2137 5494
rect 1939 5296 1995 5352
rect 2081 5296 2137 5352
rect 1939 5154 1995 5210
rect 2081 5154 2137 5210
rect 1939 5012 1995 5068
rect 2081 5012 2137 5068
rect 1939 4870 1995 4926
rect 2081 4870 2137 4926
rect 1939 4728 1995 4784
rect 2081 4728 2137 4784
rect 1939 4586 1995 4642
rect 2081 4586 2137 4642
rect 1939 4444 1995 4500
rect 2081 4444 2137 4500
rect 1939 4302 1995 4358
rect 2081 4302 2137 4358
rect 1939 4160 1995 4216
rect 2081 4160 2137 4216
rect 1939 4018 1995 4074
rect 2081 4018 2137 4074
rect 1939 3876 1995 3932
rect 2081 3876 2137 3932
rect 1939 3734 1995 3790
rect 2081 3734 2137 3790
rect 1939 3592 1995 3648
rect 2081 3592 2137 3648
rect 1939 3450 1995 3506
rect 2081 3450 2137 3506
rect 1939 3308 1995 3364
rect 2081 3308 2137 3364
rect 1939 3166 1995 3222
rect 2081 3166 2137 3222
rect 1939 3024 1995 3080
rect 2081 3024 2137 3080
rect 1939 2882 1995 2938
rect 2081 2882 2137 2938
rect 1939 2740 1995 2796
rect 2081 2740 2137 2796
rect 1939 2598 1995 2654
rect 2081 2598 2137 2654
rect 1939 2456 1995 2512
rect 2081 2456 2137 2512
rect 1939 2314 1995 2370
rect 2081 2314 2137 2370
rect 1939 2172 1995 2228
rect 2081 2172 2137 2228
rect 1939 2030 1995 2086
rect 2081 2030 2137 2086
rect 1939 1888 1995 1944
rect 2081 1888 2137 1944
rect 1939 1746 1995 1802
rect 2081 1746 2137 1802
rect 1939 1604 1995 1660
rect 2081 1604 2137 1660
rect 1939 1462 1995 1518
rect 2081 1462 2137 1518
rect 1939 1320 1995 1376
rect 2081 1320 2137 1376
rect 1939 1178 1995 1234
rect 2081 1178 2137 1234
rect 1939 1036 1995 1092
rect 2081 1036 2137 1092
rect 1939 894 1995 950
rect 2081 894 2137 950
rect 1939 752 1995 808
rect 2081 752 2137 808
rect 1939 610 1995 666
rect 2081 610 2137 666
rect 1939 468 1995 524
rect 2081 468 2137 524
rect 2336 12254 2392 12310
rect 2478 12254 2534 12310
rect 2336 12112 2392 12168
rect 2478 12112 2534 12168
rect 2336 11970 2392 12026
rect 2478 11970 2534 12026
rect 2336 11828 2392 11884
rect 2478 11828 2534 11884
rect 2336 11686 2392 11742
rect 2478 11686 2534 11742
rect 2336 11544 2392 11600
rect 2478 11544 2534 11600
rect 2336 11402 2392 11458
rect 2478 11402 2534 11458
rect 2336 11260 2392 11316
rect 2478 11260 2534 11316
rect 2336 11118 2392 11174
rect 2478 11118 2534 11174
rect 2336 10976 2392 11032
rect 2478 10976 2534 11032
rect 2336 10834 2392 10890
rect 2478 10834 2534 10890
rect 2336 10692 2392 10748
rect 2478 10692 2534 10748
rect 2336 10550 2392 10606
rect 2478 10550 2534 10606
rect 2336 10408 2392 10464
rect 2478 10408 2534 10464
rect 2336 10266 2392 10322
rect 2478 10266 2534 10322
rect 2336 10124 2392 10180
rect 2478 10124 2534 10180
rect 2336 9982 2392 10038
rect 2478 9982 2534 10038
rect 2336 9840 2392 9896
rect 2478 9840 2534 9896
rect 2336 9698 2392 9754
rect 2478 9698 2534 9754
rect 2336 9556 2392 9612
rect 2478 9556 2534 9612
rect 2336 9414 2392 9470
rect 2478 9414 2534 9470
rect 2336 9272 2392 9328
rect 2478 9272 2534 9328
rect 2336 9130 2392 9186
rect 2478 9130 2534 9186
rect 2336 8988 2392 9044
rect 2478 8988 2534 9044
rect 2336 8846 2392 8902
rect 2478 8846 2534 8902
rect 2336 8704 2392 8760
rect 2478 8704 2534 8760
rect 2336 8562 2392 8618
rect 2478 8562 2534 8618
rect 2336 8420 2392 8476
rect 2478 8420 2534 8476
rect 2336 8278 2392 8334
rect 2478 8278 2534 8334
rect 2336 8136 2392 8192
rect 2478 8136 2534 8192
rect 2336 7994 2392 8050
rect 2478 7994 2534 8050
rect 2336 7852 2392 7908
rect 2478 7852 2534 7908
rect 2336 7710 2392 7766
rect 2478 7710 2534 7766
rect 2336 7568 2392 7624
rect 2478 7568 2534 7624
rect 2336 7426 2392 7482
rect 2478 7426 2534 7482
rect 2336 7284 2392 7340
rect 2478 7284 2534 7340
rect 2336 7142 2392 7198
rect 2478 7142 2534 7198
rect 2336 7000 2392 7056
rect 2478 7000 2534 7056
rect 2336 6858 2392 6914
rect 2478 6858 2534 6914
rect 2336 6716 2392 6772
rect 2478 6716 2534 6772
rect 2336 6574 2392 6630
rect 2478 6574 2534 6630
rect 2336 6432 2392 6488
rect 2478 6432 2534 6488
rect 2336 6290 2392 6346
rect 2478 6290 2534 6346
rect 2336 6148 2392 6204
rect 2478 6148 2534 6204
rect 2336 6006 2392 6062
rect 2478 6006 2534 6062
rect 2336 5864 2392 5920
rect 2478 5864 2534 5920
rect 2336 5722 2392 5778
rect 2478 5722 2534 5778
rect 2336 5580 2392 5636
rect 2478 5580 2534 5636
rect 2336 5438 2392 5494
rect 2478 5438 2534 5494
rect 2336 5296 2392 5352
rect 2478 5296 2534 5352
rect 2336 5154 2392 5210
rect 2478 5154 2534 5210
rect 2336 5012 2392 5068
rect 2478 5012 2534 5068
rect 2336 4870 2392 4926
rect 2478 4870 2534 4926
rect 2336 4728 2392 4784
rect 2478 4728 2534 4784
rect 2336 4586 2392 4642
rect 2478 4586 2534 4642
rect 2336 4444 2392 4500
rect 2478 4444 2534 4500
rect 2336 4302 2392 4358
rect 2478 4302 2534 4358
rect 2336 4160 2392 4216
rect 2478 4160 2534 4216
rect 2336 4018 2392 4074
rect 2478 4018 2534 4074
rect 2336 3876 2392 3932
rect 2478 3876 2534 3932
rect 2336 3734 2392 3790
rect 2478 3734 2534 3790
rect 2336 3592 2392 3648
rect 2478 3592 2534 3648
rect 2336 3450 2392 3506
rect 2478 3450 2534 3506
rect 2336 3308 2392 3364
rect 2478 3308 2534 3364
rect 2336 3166 2392 3222
rect 2478 3166 2534 3222
rect 2336 3024 2392 3080
rect 2478 3024 2534 3080
rect 2336 2882 2392 2938
rect 2478 2882 2534 2938
rect 2336 2740 2392 2796
rect 2478 2740 2534 2796
rect 2336 2598 2392 2654
rect 2478 2598 2534 2654
rect 2336 2456 2392 2512
rect 2478 2456 2534 2512
rect 2336 2314 2392 2370
rect 2478 2314 2534 2370
rect 2336 2172 2392 2228
rect 2478 2172 2534 2228
rect 2336 2030 2392 2086
rect 2478 2030 2534 2086
rect 2336 1888 2392 1944
rect 2478 1888 2534 1944
rect 2336 1746 2392 1802
rect 2478 1746 2534 1802
rect 2336 1604 2392 1660
rect 2478 1604 2534 1660
rect 2336 1462 2392 1518
rect 2478 1462 2534 1518
rect 2336 1320 2392 1376
rect 2478 1320 2534 1376
rect 2336 1178 2392 1234
rect 2478 1178 2534 1234
rect 2336 1036 2392 1092
rect 2478 1036 2534 1092
rect 2336 894 2392 950
rect 2478 894 2534 950
rect 2336 752 2392 808
rect 2478 752 2534 808
rect 2336 610 2392 666
rect 2478 610 2534 666
rect 2336 468 2392 524
rect 2478 468 2534 524
rect 2740 12254 2796 12310
rect 2882 12254 2938 12310
rect 2740 12112 2796 12168
rect 2882 12112 2938 12168
rect 2740 11970 2796 12026
rect 2882 11970 2938 12026
rect 2740 11828 2796 11884
rect 2882 11828 2938 11884
rect 2740 11686 2796 11742
rect 2882 11686 2938 11742
rect 2740 11544 2796 11600
rect 2882 11544 2938 11600
rect 2740 11402 2796 11458
rect 2882 11402 2938 11458
rect 2740 11260 2796 11316
rect 2882 11260 2938 11316
rect 2740 11118 2796 11174
rect 2882 11118 2938 11174
rect 2740 10976 2796 11032
rect 2882 10976 2938 11032
rect 2740 10834 2796 10890
rect 2882 10834 2938 10890
rect 2740 10692 2796 10748
rect 2882 10692 2938 10748
rect 2740 10550 2796 10606
rect 2882 10550 2938 10606
rect 2740 10408 2796 10464
rect 2882 10408 2938 10464
rect 2740 10266 2796 10322
rect 2882 10266 2938 10322
rect 2740 10124 2796 10180
rect 2882 10124 2938 10180
rect 2740 9982 2796 10038
rect 2882 9982 2938 10038
rect 2740 9840 2796 9896
rect 2882 9840 2938 9896
rect 2740 9698 2796 9754
rect 2882 9698 2938 9754
rect 2740 9556 2796 9612
rect 2882 9556 2938 9612
rect 2740 9414 2796 9470
rect 2882 9414 2938 9470
rect 2740 9272 2796 9328
rect 2882 9272 2938 9328
rect 2740 9130 2796 9186
rect 2882 9130 2938 9186
rect 2740 8988 2796 9044
rect 2882 8988 2938 9044
rect 2740 8846 2796 8902
rect 2882 8846 2938 8902
rect 2740 8704 2796 8760
rect 2882 8704 2938 8760
rect 2740 8562 2796 8618
rect 2882 8562 2938 8618
rect 2740 8420 2796 8476
rect 2882 8420 2938 8476
rect 2740 8278 2796 8334
rect 2882 8278 2938 8334
rect 2740 8136 2796 8192
rect 2882 8136 2938 8192
rect 2740 7994 2796 8050
rect 2882 7994 2938 8050
rect 2740 7852 2796 7908
rect 2882 7852 2938 7908
rect 2740 7710 2796 7766
rect 2882 7710 2938 7766
rect 2740 7568 2796 7624
rect 2882 7568 2938 7624
rect 2740 7426 2796 7482
rect 2882 7426 2938 7482
rect 2740 7284 2796 7340
rect 2882 7284 2938 7340
rect 2740 7142 2796 7198
rect 2882 7142 2938 7198
rect 2740 7000 2796 7056
rect 2882 7000 2938 7056
rect 2740 6858 2796 6914
rect 2882 6858 2938 6914
rect 2740 6716 2796 6772
rect 2882 6716 2938 6772
rect 2740 6574 2796 6630
rect 2882 6574 2938 6630
rect 2740 6432 2796 6488
rect 2882 6432 2938 6488
rect 2740 6290 2796 6346
rect 2882 6290 2938 6346
rect 2740 6148 2796 6204
rect 2882 6148 2938 6204
rect 2740 6006 2796 6062
rect 2882 6006 2938 6062
rect 2740 5864 2796 5920
rect 2882 5864 2938 5920
rect 2740 5722 2796 5778
rect 2882 5722 2938 5778
rect 2740 5580 2796 5636
rect 2882 5580 2938 5636
rect 2740 5438 2796 5494
rect 2882 5438 2938 5494
rect 2740 5296 2796 5352
rect 2882 5296 2938 5352
rect 2740 5154 2796 5210
rect 2882 5154 2938 5210
rect 2740 5012 2796 5068
rect 2882 5012 2938 5068
rect 2740 4870 2796 4926
rect 2882 4870 2938 4926
rect 2740 4728 2796 4784
rect 2882 4728 2938 4784
rect 2740 4586 2796 4642
rect 2882 4586 2938 4642
rect 2740 4444 2796 4500
rect 2882 4444 2938 4500
rect 2740 4302 2796 4358
rect 2882 4302 2938 4358
rect 2740 4160 2796 4216
rect 2882 4160 2938 4216
rect 2740 4018 2796 4074
rect 2882 4018 2938 4074
rect 2740 3876 2796 3932
rect 2882 3876 2938 3932
rect 2740 3734 2796 3790
rect 2882 3734 2938 3790
rect 2740 3592 2796 3648
rect 2882 3592 2938 3648
rect 2740 3450 2796 3506
rect 2882 3450 2938 3506
rect 2740 3308 2796 3364
rect 2882 3308 2938 3364
rect 2740 3166 2796 3222
rect 2882 3166 2938 3222
rect 2740 3024 2796 3080
rect 2882 3024 2938 3080
rect 2740 2882 2796 2938
rect 2882 2882 2938 2938
rect 2740 2740 2796 2796
rect 2882 2740 2938 2796
rect 2740 2598 2796 2654
rect 2882 2598 2938 2654
rect 2740 2456 2796 2512
rect 2882 2456 2938 2512
rect 2740 2314 2796 2370
rect 2882 2314 2938 2370
rect 2740 2172 2796 2228
rect 2882 2172 2938 2228
rect 2740 2030 2796 2086
rect 2882 2030 2938 2086
rect 2740 1888 2796 1944
rect 2882 1888 2938 1944
rect 2740 1746 2796 1802
rect 2882 1746 2938 1802
rect 2740 1604 2796 1660
rect 2882 1604 2938 1660
rect 2740 1462 2796 1518
rect 2882 1462 2938 1518
rect 2740 1320 2796 1376
rect 2882 1320 2938 1376
rect 2740 1178 2796 1234
rect 2882 1178 2938 1234
rect 2740 1036 2796 1092
rect 2882 1036 2938 1092
rect 2740 894 2796 950
rect 2882 894 2938 950
rect 2740 752 2796 808
rect 2882 752 2938 808
rect 2740 610 2796 666
rect 2882 610 2938 666
rect 2740 468 2796 524
rect 2882 468 2938 524
rect 3136 12254 3192 12310
rect 3278 12254 3334 12310
rect 3136 12112 3192 12168
rect 3278 12112 3334 12168
rect 3136 11970 3192 12026
rect 3278 11970 3334 12026
rect 3136 11828 3192 11884
rect 3278 11828 3334 11884
rect 3136 11686 3192 11742
rect 3278 11686 3334 11742
rect 3136 11544 3192 11600
rect 3278 11544 3334 11600
rect 3136 11402 3192 11458
rect 3278 11402 3334 11458
rect 3136 11260 3192 11316
rect 3278 11260 3334 11316
rect 3136 11118 3192 11174
rect 3278 11118 3334 11174
rect 3136 10976 3192 11032
rect 3278 10976 3334 11032
rect 3136 10834 3192 10890
rect 3278 10834 3334 10890
rect 3136 10692 3192 10748
rect 3278 10692 3334 10748
rect 3136 10550 3192 10606
rect 3278 10550 3334 10606
rect 3136 10408 3192 10464
rect 3278 10408 3334 10464
rect 3136 10266 3192 10322
rect 3278 10266 3334 10322
rect 3136 10124 3192 10180
rect 3278 10124 3334 10180
rect 3136 9982 3192 10038
rect 3278 9982 3334 10038
rect 3136 9840 3192 9896
rect 3278 9840 3334 9896
rect 3136 9698 3192 9754
rect 3278 9698 3334 9754
rect 3136 9556 3192 9612
rect 3278 9556 3334 9612
rect 3136 9414 3192 9470
rect 3278 9414 3334 9470
rect 3136 9272 3192 9328
rect 3278 9272 3334 9328
rect 3136 9130 3192 9186
rect 3278 9130 3334 9186
rect 3136 8988 3192 9044
rect 3278 8988 3334 9044
rect 3136 8846 3192 8902
rect 3278 8846 3334 8902
rect 3136 8704 3192 8760
rect 3278 8704 3334 8760
rect 3136 8562 3192 8618
rect 3278 8562 3334 8618
rect 3136 8420 3192 8476
rect 3278 8420 3334 8476
rect 3136 8278 3192 8334
rect 3278 8278 3334 8334
rect 3136 8136 3192 8192
rect 3278 8136 3334 8192
rect 3136 7994 3192 8050
rect 3278 7994 3334 8050
rect 3136 7852 3192 7908
rect 3278 7852 3334 7908
rect 3136 7710 3192 7766
rect 3278 7710 3334 7766
rect 3136 7568 3192 7624
rect 3278 7568 3334 7624
rect 3136 7426 3192 7482
rect 3278 7426 3334 7482
rect 3136 7284 3192 7340
rect 3278 7284 3334 7340
rect 3136 7142 3192 7198
rect 3278 7142 3334 7198
rect 3136 7000 3192 7056
rect 3278 7000 3334 7056
rect 3136 6858 3192 6914
rect 3278 6858 3334 6914
rect 3136 6716 3192 6772
rect 3278 6716 3334 6772
rect 3136 6574 3192 6630
rect 3278 6574 3334 6630
rect 3136 6432 3192 6488
rect 3278 6432 3334 6488
rect 3136 6290 3192 6346
rect 3278 6290 3334 6346
rect 3136 6148 3192 6204
rect 3278 6148 3334 6204
rect 3136 6006 3192 6062
rect 3278 6006 3334 6062
rect 3136 5864 3192 5920
rect 3278 5864 3334 5920
rect 3136 5722 3192 5778
rect 3278 5722 3334 5778
rect 3136 5580 3192 5636
rect 3278 5580 3334 5636
rect 3136 5438 3192 5494
rect 3278 5438 3334 5494
rect 3136 5296 3192 5352
rect 3278 5296 3334 5352
rect 3136 5154 3192 5210
rect 3278 5154 3334 5210
rect 3136 5012 3192 5068
rect 3278 5012 3334 5068
rect 3136 4870 3192 4926
rect 3278 4870 3334 4926
rect 3136 4728 3192 4784
rect 3278 4728 3334 4784
rect 3136 4586 3192 4642
rect 3278 4586 3334 4642
rect 3136 4444 3192 4500
rect 3278 4444 3334 4500
rect 3136 4302 3192 4358
rect 3278 4302 3334 4358
rect 3136 4160 3192 4216
rect 3278 4160 3334 4216
rect 3136 4018 3192 4074
rect 3278 4018 3334 4074
rect 3136 3876 3192 3932
rect 3278 3876 3334 3932
rect 3136 3734 3192 3790
rect 3278 3734 3334 3790
rect 3136 3592 3192 3648
rect 3278 3592 3334 3648
rect 3136 3450 3192 3506
rect 3278 3450 3334 3506
rect 3136 3308 3192 3364
rect 3278 3308 3334 3364
rect 3136 3166 3192 3222
rect 3278 3166 3334 3222
rect 3136 3024 3192 3080
rect 3278 3024 3334 3080
rect 3136 2882 3192 2938
rect 3278 2882 3334 2938
rect 3136 2740 3192 2796
rect 3278 2740 3334 2796
rect 3136 2598 3192 2654
rect 3278 2598 3334 2654
rect 3136 2456 3192 2512
rect 3278 2456 3334 2512
rect 3136 2314 3192 2370
rect 3278 2314 3334 2370
rect 3136 2172 3192 2228
rect 3278 2172 3334 2228
rect 3136 2030 3192 2086
rect 3278 2030 3334 2086
rect 3136 1888 3192 1944
rect 3278 1888 3334 1944
rect 3136 1746 3192 1802
rect 3278 1746 3334 1802
rect 3136 1604 3192 1660
rect 3278 1604 3334 1660
rect 3136 1462 3192 1518
rect 3278 1462 3334 1518
rect 3136 1320 3192 1376
rect 3278 1320 3334 1376
rect 3136 1178 3192 1234
rect 3278 1178 3334 1234
rect 3136 1036 3192 1092
rect 3278 1036 3334 1092
rect 3136 894 3192 950
rect 3278 894 3334 950
rect 3136 752 3192 808
rect 3278 752 3334 808
rect 3136 610 3192 666
rect 3278 610 3334 666
rect 3136 468 3192 524
rect 3278 468 3334 524
rect 3536 12254 3592 12310
rect 3678 12254 3734 12310
rect 3536 12112 3592 12168
rect 3678 12112 3734 12168
rect 3536 11970 3592 12026
rect 3678 11970 3734 12026
rect 3536 11828 3592 11884
rect 3678 11828 3734 11884
rect 3536 11686 3592 11742
rect 3678 11686 3734 11742
rect 3536 11544 3592 11600
rect 3678 11544 3734 11600
rect 3536 11402 3592 11458
rect 3678 11402 3734 11458
rect 3536 11260 3592 11316
rect 3678 11260 3734 11316
rect 3536 11118 3592 11174
rect 3678 11118 3734 11174
rect 3536 10976 3592 11032
rect 3678 10976 3734 11032
rect 3536 10834 3592 10890
rect 3678 10834 3734 10890
rect 3536 10692 3592 10748
rect 3678 10692 3734 10748
rect 3536 10550 3592 10606
rect 3678 10550 3734 10606
rect 3536 10408 3592 10464
rect 3678 10408 3734 10464
rect 3536 10266 3592 10322
rect 3678 10266 3734 10322
rect 3536 10124 3592 10180
rect 3678 10124 3734 10180
rect 3536 9982 3592 10038
rect 3678 9982 3734 10038
rect 3536 9840 3592 9896
rect 3678 9840 3734 9896
rect 3536 9698 3592 9754
rect 3678 9698 3734 9754
rect 3536 9556 3592 9612
rect 3678 9556 3734 9612
rect 3536 9414 3592 9470
rect 3678 9414 3734 9470
rect 3536 9272 3592 9328
rect 3678 9272 3734 9328
rect 3536 9130 3592 9186
rect 3678 9130 3734 9186
rect 3536 8988 3592 9044
rect 3678 8988 3734 9044
rect 3536 8846 3592 8902
rect 3678 8846 3734 8902
rect 3536 8704 3592 8760
rect 3678 8704 3734 8760
rect 3536 8562 3592 8618
rect 3678 8562 3734 8618
rect 3536 8420 3592 8476
rect 3678 8420 3734 8476
rect 3536 8278 3592 8334
rect 3678 8278 3734 8334
rect 3536 8136 3592 8192
rect 3678 8136 3734 8192
rect 3536 7994 3592 8050
rect 3678 7994 3734 8050
rect 3536 7852 3592 7908
rect 3678 7852 3734 7908
rect 3536 7710 3592 7766
rect 3678 7710 3734 7766
rect 3536 7568 3592 7624
rect 3678 7568 3734 7624
rect 3536 7426 3592 7482
rect 3678 7426 3734 7482
rect 3536 7284 3592 7340
rect 3678 7284 3734 7340
rect 3536 7142 3592 7198
rect 3678 7142 3734 7198
rect 3536 7000 3592 7056
rect 3678 7000 3734 7056
rect 3536 6858 3592 6914
rect 3678 6858 3734 6914
rect 3536 6716 3592 6772
rect 3678 6716 3734 6772
rect 3536 6574 3592 6630
rect 3678 6574 3734 6630
rect 3536 6432 3592 6488
rect 3678 6432 3734 6488
rect 3536 6290 3592 6346
rect 3678 6290 3734 6346
rect 3536 6148 3592 6204
rect 3678 6148 3734 6204
rect 3536 6006 3592 6062
rect 3678 6006 3734 6062
rect 3536 5864 3592 5920
rect 3678 5864 3734 5920
rect 3536 5722 3592 5778
rect 3678 5722 3734 5778
rect 3536 5580 3592 5636
rect 3678 5580 3734 5636
rect 3536 5438 3592 5494
rect 3678 5438 3734 5494
rect 3536 5296 3592 5352
rect 3678 5296 3734 5352
rect 3536 5154 3592 5210
rect 3678 5154 3734 5210
rect 3536 5012 3592 5068
rect 3678 5012 3734 5068
rect 3536 4870 3592 4926
rect 3678 4870 3734 4926
rect 3536 4728 3592 4784
rect 3678 4728 3734 4784
rect 3536 4586 3592 4642
rect 3678 4586 3734 4642
rect 3536 4444 3592 4500
rect 3678 4444 3734 4500
rect 3536 4302 3592 4358
rect 3678 4302 3734 4358
rect 3536 4160 3592 4216
rect 3678 4160 3734 4216
rect 3536 4018 3592 4074
rect 3678 4018 3734 4074
rect 3536 3876 3592 3932
rect 3678 3876 3734 3932
rect 3536 3734 3592 3790
rect 3678 3734 3734 3790
rect 3536 3592 3592 3648
rect 3678 3592 3734 3648
rect 3536 3450 3592 3506
rect 3678 3450 3734 3506
rect 3536 3308 3592 3364
rect 3678 3308 3734 3364
rect 3536 3166 3592 3222
rect 3678 3166 3734 3222
rect 3536 3024 3592 3080
rect 3678 3024 3734 3080
rect 3536 2882 3592 2938
rect 3678 2882 3734 2938
rect 3536 2740 3592 2796
rect 3678 2740 3734 2796
rect 3536 2598 3592 2654
rect 3678 2598 3734 2654
rect 3536 2456 3592 2512
rect 3678 2456 3734 2512
rect 3536 2314 3592 2370
rect 3678 2314 3734 2370
rect 3536 2172 3592 2228
rect 3678 2172 3734 2228
rect 3536 2030 3592 2086
rect 3678 2030 3734 2086
rect 3536 1888 3592 1944
rect 3678 1888 3734 1944
rect 3536 1746 3592 1802
rect 3678 1746 3734 1802
rect 3536 1604 3592 1660
rect 3678 1604 3734 1660
rect 3536 1462 3592 1518
rect 3678 1462 3734 1518
rect 3536 1320 3592 1376
rect 3678 1320 3734 1376
rect 3536 1178 3592 1234
rect 3678 1178 3734 1234
rect 3536 1036 3592 1092
rect 3678 1036 3734 1092
rect 3536 894 3592 950
rect 3678 894 3734 950
rect 3536 752 3592 808
rect 3678 752 3734 808
rect 3536 610 3592 666
rect 3678 610 3734 666
rect 3536 468 3592 524
rect 3678 468 3734 524
rect 3933 12254 3989 12310
rect 4075 12254 4131 12310
rect 3933 12112 3989 12168
rect 4075 12112 4131 12168
rect 3933 11970 3989 12026
rect 4075 11970 4131 12026
rect 3933 11828 3989 11884
rect 4075 11828 4131 11884
rect 3933 11686 3989 11742
rect 4075 11686 4131 11742
rect 3933 11544 3989 11600
rect 4075 11544 4131 11600
rect 3933 11402 3989 11458
rect 4075 11402 4131 11458
rect 3933 11260 3989 11316
rect 4075 11260 4131 11316
rect 3933 11118 3989 11174
rect 4075 11118 4131 11174
rect 3933 10976 3989 11032
rect 4075 10976 4131 11032
rect 3933 10834 3989 10890
rect 4075 10834 4131 10890
rect 3933 10692 3989 10748
rect 4075 10692 4131 10748
rect 3933 10550 3989 10606
rect 4075 10550 4131 10606
rect 3933 10408 3989 10464
rect 4075 10408 4131 10464
rect 3933 10266 3989 10322
rect 4075 10266 4131 10322
rect 3933 10124 3989 10180
rect 4075 10124 4131 10180
rect 3933 9982 3989 10038
rect 4075 9982 4131 10038
rect 3933 9840 3989 9896
rect 4075 9840 4131 9896
rect 3933 9698 3989 9754
rect 4075 9698 4131 9754
rect 3933 9556 3989 9612
rect 4075 9556 4131 9612
rect 3933 9414 3989 9470
rect 4075 9414 4131 9470
rect 3933 9272 3989 9328
rect 4075 9272 4131 9328
rect 3933 9130 3989 9186
rect 4075 9130 4131 9186
rect 3933 8988 3989 9044
rect 4075 8988 4131 9044
rect 3933 8846 3989 8902
rect 4075 8846 4131 8902
rect 3933 8704 3989 8760
rect 4075 8704 4131 8760
rect 3933 8562 3989 8618
rect 4075 8562 4131 8618
rect 3933 8420 3989 8476
rect 4075 8420 4131 8476
rect 3933 8278 3989 8334
rect 4075 8278 4131 8334
rect 3933 8136 3989 8192
rect 4075 8136 4131 8192
rect 3933 7994 3989 8050
rect 4075 7994 4131 8050
rect 3933 7852 3989 7908
rect 4075 7852 4131 7908
rect 3933 7710 3989 7766
rect 4075 7710 4131 7766
rect 3933 7568 3989 7624
rect 4075 7568 4131 7624
rect 3933 7426 3989 7482
rect 4075 7426 4131 7482
rect 3933 7284 3989 7340
rect 4075 7284 4131 7340
rect 3933 7142 3989 7198
rect 4075 7142 4131 7198
rect 3933 7000 3989 7056
rect 4075 7000 4131 7056
rect 3933 6858 3989 6914
rect 4075 6858 4131 6914
rect 3933 6716 3989 6772
rect 4075 6716 4131 6772
rect 3933 6574 3989 6630
rect 4075 6574 4131 6630
rect 3933 6432 3989 6488
rect 4075 6432 4131 6488
rect 3933 6290 3989 6346
rect 4075 6290 4131 6346
rect 3933 6148 3989 6204
rect 4075 6148 4131 6204
rect 3933 6006 3989 6062
rect 4075 6006 4131 6062
rect 3933 5864 3989 5920
rect 4075 5864 4131 5920
rect 3933 5722 3989 5778
rect 4075 5722 4131 5778
rect 3933 5580 3989 5636
rect 4075 5580 4131 5636
rect 3933 5438 3989 5494
rect 4075 5438 4131 5494
rect 3933 5296 3989 5352
rect 4075 5296 4131 5352
rect 3933 5154 3989 5210
rect 4075 5154 4131 5210
rect 3933 5012 3989 5068
rect 4075 5012 4131 5068
rect 3933 4870 3989 4926
rect 4075 4870 4131 4926
rect 3933 4728 3989 4784
rect 4075 4728 4131 4784
rect 3933 4586 3989 4642
rect 4075 4586 4131 4642
rect 3933 4444 3989 4500
rect 4075 4444 4131 4500
rect 3933 4302 3989 4358
rect 4075 4302 4131 4358
rect 3933 4160 3989 4216
rect 4075 4160 4131 4216
rect 3933 4018 3989 4074
rect 4075 4018 4131 4074
rect 3933 3876 3989 3932
rect 4075 3876 4131 3932
rect 3933 3734 3989 3790
rect 4075 3734 4131 3790
rect 3933 3592 3989 3648
rect 4075 3592 4131 3648
rect 3933 3450 3989 3506
rect 4075 3450 4131 3506
rect 3933 3308 3989 3364
rect 4075 3308 4131 3364
rect 3933 3166 3989 3222
rect 4075 3166 4131 3222
rect 3933 3024 3989 3080
rect 4075 3024 4131 3080
rect 3933 2882 3989 2938
rect 4075 2882 4131 2938
rect 3933 2740 3989 2796
rect 4075 2740 4131 2796
rect 3933 2598 3989 2654
rect 4075 2598 4131 2654
rect 3933 2456 3989 2512
rect 4075 2456 4131 2512
rect 3933 2314 3989 2370
rect 4075 2314 4131 2370
rect 3933 2172 3989 2228
rect 4075 2172 4131 2228
rect 3933 2030 3989 2086
rect 4075 2030 4131 2086
rect 3933 1888 3989 1944
rect 4075 1888 4131 1944
rect 3933 1746 3989 1802
rect 4075 1746 4131 1802
rect 3933 1604 3989 1660
rect 4075 1604 4131 1660
rect 3933 1462 3989 1518
rect 4075 1462 4131 1518
rect 3933 1320 3989 1376
rect 4075 1320 4131 1376
rect 3933 1178 3989 1234
rect 4075 1178 4131 1234
rect 3933 1036 3989 1092
rect 4075 1036 4131 1092
rect 3933 894 3989 950
rect 4075 894 4131 950
rect 3933 752 3989 808
rect 4075 752 4131 808
rect 3933 610 3989 666
rect 4075 610 4131 666
rect 3933 468 3989 524
rect 4075 468 4131 524
rect 4338 12254 4394 12310
rect 4480 12254 4536 12310
rect 4338 12112 4394 12168
rect 4480 12112 4536 12168
rect 4338 11970 4394 12026
rect 4480 11970 4536 12026
rect 4338 11828 4394 11884
rect 4480 11828 4536 11884
rect 4338 11686 4394 11742
rect 4480 11686 4536 11742
rect 4338 11544 4394 11600
rect 4480 11544 4536 11600
rect 4338 11402 4394 11458
rect 4480 11402 4536 11458
rect 4338 11260 4394 11316
rect 4480 11260 4536 11316
rect 4338 11118 4394 11174
rect 4480 11118 4536 11174
rect 4338 10976 4394 11032
rect 4480 10976 4536 11032
rect 4338 10834 4394 10890
rect 4480 10834 4536 10890
rect 4338 10692 4394 10748
rect 4480 10692 4536 10748
rect 4338 10550 4394 10606
rect 4480 10550 4536 10606
rect 4338 10408 4394 10464
rect 4480 10408 4536 10464
rect 4338 10266 4394 10322
rect 4480 10266 4536 10322
rect 4338 10124 4394 10180
rect 4480 10124 4536 10180
rect 4338 9982 4394 10038
rect 4480 9982 4536 10038
rect 4338 9840 4394 9896
rect 4480 9840 4536 9896
rect 4338 9698 4394 9754
rect 4480 9698 4536 9754
rect 4338 9556 4394 9612
rect 4480 9556 4536 9612
rect 4338 9414 4394 9470
rect 4480 9414 4536 9470
rect 4338 9272 4394 9328
rect 4480 9272 4536 9328
rect 4338 9130 4394 9186
rect 4480 9130 4536 9186
rect 4338 8988 4394 9044
rect 4480 8988 4536 9044
rect 4338 8846 4394 8902
rect 4480 8846 4536 8902
rect 4338 8704 4394 8760
rect 4480 8704 4536 8760
rect 4338 8562 4394 8618
rect 4480 8562 4536 8618
rect 4338 8420 4394 8476
rect 4480 8420 4536 8476
rect 4338 8278 4394 8334
rect 4480 8278 4536 8334
rect 4338 8136 4394 8192
rect 4480 8136 4536 8192
rect 4338 7994 4394 8050
rect 4480 7994 4536 8050
rect 4338 7852 4394 7908
rect 4480 7852 4536 7908
rect 4338 7710 4394 7766
rect 4480 7710 4536 7766
rect 4338 7568 4394 7624
rect 4480 7568 4536 7624
rect 4338 7426 4394 7482
rect 4480 7426 4536 7482
rect 4338 7284 4394 7340
rect 4480 7284 4536 7340
rect 4338 7142 4394 7198
rect 4480 7142 4536 7198
rect 4338 7000 4394 7056
rect 4480 7000 4536 7056
rect 4338 6858 4394 6914
rect 4480 6858 4536 6914
rect 4338 6716 4394 6772
rect 4480 6716 4536 6772
rect 4338 6574 4394 6630
rect 4480 6574 4536 6630
rect 4338 6432 4394 6488
rect 4480 6432 4536 6488
rect 4338 6290 4394 6346
rect 4480 6290 4536 6346
rect 4338 6148 4394 6204
rect 4480 6148 4536 6204
rect 4338 6006 4394 6062
rect 4480 6006 4536 6062
rect 4338 5864 4394 5920
rect 4480 5864 4536 5920
rect 4338 5722 4394 5778
rect 4480 5722 4536 5778
rect 4338 5580 4394 5636
rect 4480 5580 4536 5636
rect 4338 5438 4394 5494
rect 4480 5438 4536 5494
rect 4338 5296 4394 5352
rect 4480 5296 4536 5352
rect 4338 5154 4394 5210
rect 4480 5154 4536 5210
rect 4338 5012 4394 5068
rect 4480 5012 4536 5068
rect 4338 4870 4394 4926
rect 4480 4870 4536 4926
rect 4338 4728 4394 4784
rect 4480 4728 4536 4784
rect 4338 4586 4394 4642
rect 4480 4586 4536 4642
rect 4338 4444 4394 4500
rect 4480 4444 4536 4500
rect 4338 4302 4394 4358
rect 4480 4302 4536 4358
rect 4338 4160 4394 4216
rect 4480 4160 4536 4216
rect 4338 4018 4394 4074
rect 4480 4018 4536 4074
rect 4338 3876 4394 3932
rect 4480 3876 4536 3932
rect 4338 3734 4394 3790
rect 4480 3734 4536 3790
rect 4338 3592 4394 3648
rect 4480 3592 4536 3648
rect 4338 3450 4394 3506
rect 4480 3450 4536 3506
rect 4338 3308 4394 3364
rect 4480 3308 4536 3364
rect 4338 3166 4394 3222
rect 4480 3166 4536 3222
rect 4338 3024 4394 3080
rect 4480 3024 4536 3080
rect 4338 2882 4394 2938
rect 4480 2882 4536 2938
rect 4338 2740 4394 2796
rect 4480 2740 4536 2796
rect 4338 2598 4394 2654
rect 4480 2598 4536 2654
rect 4338 2456 4394 2512
rect 4480 2456 4536 2512
rect 4338 2314 4394 2370
rect 4480 2314 4536 2370
rect 4338 2172 4394 2228
rect 4480 2172 4536 2228
rect 4338 2030 4394 2086
rect 4480 2030 4536 2086
rect 4338 1888 4394 1944
rect 4480 1888 4536 1944
rect 4338 1746 4394 1802
rect 4480 1746 4536 1802
rect 4338 1604 4394 1660
rect 4480 1604 4536 1660
rect 4338 1462 4394 1518
rect 4480 1462 4536 1518
rect 4338 1320 4394 1376
rect 4480 1320 4536 1376
rect 4338 1178 4394 1234
rect 4480 1178 4536 1234
rect 4338 1036 4394 1092
rect 4480 1036 4536 1092
rect 4338 894 4394 950
rect 4480 894 4536 950
rect 4338 752 4394 808
rect 4480 752 4536 808
rect 4338 610 4394 666
rect 4480 610 4536 666
rect 4338 468 4394 524
rect 4480 468 4536 524
rect 4738 12254 4794 12310
rect 4880 12254 4936 12310
rect 4738 12112 4794 12168
rect 4880 12112 4936 12168
rect 4738 11970 4794 12026
rect 4880 11970 4936 12026
rect 4738 11828 4794 11884
rect 4880 11828 4936 11884
rect 4738 11686 4794 11742
rect 4880 11686 4936 11742
rect 4738 11544 4794 11600
rect 4880 11544 4936 11600
rect 4738 11402 4794 11458
rect 4880 11402 4936 11458
rect 4738 11260 4794 11316
rect 4880 11260 4936 11316
rect 4738 11118 4794 11174
rect 4880 11118 4936 11174
rect 4738 10976 4794 11032
rect 4880 10976 4936 11032
rect 4738 10834 4794 10890
rect 4880 10834 4936 10890
rect 4738 10692 4794 10748
rect 4880 10692 4936 10748
rect 4738 10550 4794 10606
rect 4880 10550 4936 10606
rect 4738 10408 4794 10464
rect 4880 10408 4936 10464
rect 4738 10266 4794 10322
rect 4880 10266 4936 10322
rect 4738 10124 4794 10180
rect 4880 10124 4936 10180
rect 4738 9982 4794 10038
rect 4880 9982 4936 10038
rect 4738 9840 4794 9896
rect 4880 9840 4936 9896
rect 4738 9698 4794 9754
rect 4880 9698 4936 9754
rect 4738 9556 4794 9612
rect 4880 9556 4936 9612
rect 4738 9414 4794 9470
rect 4880 9414 4936 9470
rect 4738 9272 4794 9328
rect 4880 9272 4936 9328
rect 4738 9130 4794 9186
rect 4880 9130 4936 9186
rect 4738 8988 4794 9044
rect 4880 8988 4936 9044
rect 4738 8846 4794 8902
rect 4880 8846 4936 8902
rect 4738 8704 4794 8760
rect 4880 8704 4936 8760
rect 4738 8562 4794 8618
rect 4880 8562 4936 8618
rect 4738 8420 4794 8476
rect 4880 8420 4936 8476
rect 4738 8278 4794 8334
rect 4880 8278 4936 8334
rect 4738 8136 4794 8192
rect 4880 8136 4936 8192
rect 4738 7994 4794 8050
rect 4880 7994 4936 8050
rect 4738 7852 4794 7908
rect 4880 7852 4936 7908
rect 4738 7710 4794 7766
rect 4880 7710 4936 7766
rect 4738 7568 4794 7624
rect 4880 7568 4936 7624
rect 4738 7426 4794 7482
rect 4880 7426 4936 7482
rect 4738 7284 4794 7340
rect 4880 7284 4936 7340
rect 4738 7142 4794 7198
rect 4880 7142 4936 7198
rect 4738 7000 4794 7056
rect 4880 7000 4936 7056
rect 4738 6858 4794 6914
rect 4880 6858 4936 6914
rect 4738 6716 4794 6772
rect 4880 6716 4936 6772
rect 4738 6574 4794 6630
rect 4880 6574 4936 6630
rect 4738 6432 4794 6488
rect 4880 6432 4936 6488
rect 4738 6290 4794 6346
rect 4880 6290 4936 6346
rect 4738 6148 4794 6204
rect 4880 6148 4936 6204
rect 4738 6006 4794 6062
rect 4880 6006 4936 6062
rect 4738 5864 4794 5920
rect 4880 5864 4936 5920
rect 4738 5722 4794 5778
rect 4880 5722 4936 5778
rect 4738 5580 4794 5636
rect 4880 5580 4936 5636
rect 4738 5438 4794 5494
rect 4880 5438 4936 5494
rect 4738 5296 4794 5352
rect 4880 5296 4936 5352
rect 4738 5154 4794 5210
rect 4880 5154 4936 5210
rect 4738 5012 4794 5068
rect 4880 5012 4936 5068
rect 4738 4870 4794 4926
rect 4880 4870 4936 4926
rect 4738 4728 4794 4784
rect 4880 4728 4936 4784
rect 4738 4586 4794 4642
rect 4880 4586 4936 4642
rect 4738 4444 4794 4500
rect 4880 4444 4936 4500
rect 4738 4302 4794 4358
rect 4880 4302 4936 4358
rect 4738 4160 4794 4216
rect 4880 4160 4936 4216
rect 4738 4018 4794 4074
rect 4880 4018 4936 4074
rect 4738 3876 4794 3932
rect 4880 3876 4936 3932
rect 4738 3734 4794 3790
rect 4880 3734 4936 3790
rect 4738 3592 4794 3648
rect 4880 3592 4936 3648
rect 4738 3450 4794 3506
rect 4880 3450 4936 3506
rect 4738 3308 4794 3364
rect 4880 3308 4936 3364
rect 4738 3166 4794 3222
rect 4880 3166 4936 3222
rect 4738 3024 4794 3080
rect 4880 3024 4936 3080
rect 4738 2882 4794 2938
rect 4880 2882 4936 2938
rect 4738 2740 4794 2796
rect 4880 2740 4936 2796
rect 4738 2598 4794 2654
rect 4880 2598 4936 2654
rect 4738 2456 4794 2512
rect 4880 2456 4936 2512
rect 4738 2314 4794 2370
rect 4880 2314 4936 2370
rect 4738 2172 4794 2228
rect 4880 2172 4936 2228
rect 4738 2030 4794 2086
rect 4880 2030 4936 2086
rect 4738 1888 4794 1944
rect 4880 1888 4936 1944
rect 4738 1746 4794 1802
rect 4880 1746 4936 1802
rect 4738 1604 4794 1660
rect 4880 1604 4936 1660
rect 4738 1462 4794 1518
rect 4880 1462 4936 1518
rect 4738 1320 4794 1376
rect 4880 1320 4936 1376
rect 4738 1178 4794 1234
rect 4880 1178 4936 1234
rect 4738 1036 4794 1092
rect 4880 1036 4936 1092
rect 4738 894 4794 950
rect 4880 894 4936 950
rect 4738 752 4794 808
rect 4880 752 4936 808
rect 4738 610 4794 666
rect 4880 610 4936 666
rect 4738 468 4794 524
rect 4880 468 4936 524
rect 5143 12254 5199 12310
rect 5285 12254 5341 12310
rect 5143 12112 5199 12168
rect 5285 12112 5341 12168
rect 5143 11970 5199 12026
rect 5285 11970 5341 12026
rect 5143 11828 5199 11884
rect 5285 11828 5341 11884
rect 5143 11686 5199 11742
rect 5285 11686 5341 11742
rect 5143 11544 5199 11600
rect 5285 11544 5341 11600
rect 5143 11402 5199 11458
rect 5285 11402 5341 11458
rect 5143 11260 5199 11316
rect 5285 11260 5341 11316
rect 5143 11118 5199 11174
rect 5285 11118 5341 11174
rect 5143 10976 5199 11032
rect 5285 10976 5341 11032
rect 5143 10834 5199 10890
rect 5285 10834 5341 10890
rect 5143 10692 5199 10748
rect 5285 10692 5341 10748
rect 5143 10550 5199 10606
rect 5285 10550 5341 10606
rect 5143 10408 5199 10464
rect 5285 10408 5341 10464
rect 5143 10266 5199 10322
rect 5285 10266 5341 10322
rect 5143 10124 5199 10180
rect 5285 10124 5341 10180
rect 5143 9982 5199 10038
rect 5285 9982 5341 10038
rect 5143 9840 5199 9896
rect 5285 9840 5341 9896
rect 5143 9698 5199 9754
rect 5285 9698 5341 9754
rect 5143 9556 5199 9612
rect 5285 9556 5341 9612
rect 5143 9414 5199 9470
rect 5285 9414 5341 9470
rect 5143 9272 5199 9328
rect 5285 9272 5341 9328
rect 5143 9130 5199 9186
rect 5285 9130 5341 9186
rect 5143 8988 5199 9044
rect 5285 8988 5341 9044
rect 5143 8846 5199 8902
rect 5285 8846 5341 8902
rect 5143 8704 5199 8760
rect 5285 8704 5341 8760
rect 5143 8562 5199 8618
rect 5285 8562 5341 8618
rect 5143 8420 5199 8476
rect 5285 8420 5341 8476
rect 5143 8278 5199 8334
rect 5285 8278 5341 8334
rect 5143 8136 5199 8192
rect 5285 8136 5341 8192
rect 5143 7994 5199 8050
rect 5285 7994 5341 8050
rect 5143 7852 5199 7908
rect 5285 7852 5341 7908
rect 5143 7710 5199 7766
rect 5285 7710 5341 7766
rect 5143 7568 5199 7624
rect 5285 7568 5341 7624
rect 5143 7426 5199 7482
rect 5285 7426 5341 7482
rect 5143 7284 5199 7340
rect 5285 7284 5341 7340
rect 5143 7142 5199 7198
rect 5285 7142 5341 7198
rect 5143 7000 5199 7056
rect 5285 7000 5341 7056
rect 5143 6858 5199 6914
rect 5285 6858 5341 6914
rect 5143 6716 5199 6772
rect 5285 6716 5341 6772
rect 5143 6574 5199 6630
rect 5285 6574 5341 6630
rect 5143 6432 5199 6488
rect 5285 6432 5341 6488
rect 5143 6290 5199 6346
rect 5285 6290 5341 6346
rect 5143 6148 5199 6204
rect 5285 6148 5341 6204
rect 5143 6006 5199 6062
rect 5285 6006 5341 6062
rect 5143 5864 5199 5920
rect 5285 5864 5341 5920
rect 5143 5722 5199 5778
rect 5285 5722 5341 5778
rect 5143 5580 5199 5636
rect 5285 5580 5341 5636
rect 5143 5438 5199 5494
rect 5285 5438 5341 5494
rect 5143 5296 5199 5352
rect 5285 5296 5341 5352
rect 5143 5154 5199 5210
rect 5285 5154 5341 5210
rect 5143 5012 5199 5068
rect 5285 5012 5341 5068
rect 5143 4870 5199 4926
rect 5285 4870 5341 4926
rect 5143 4728 5199 4784
rect 5285 4728 5341 4784
rect 5143 4586 5199 4642
rect 5285 4586 5341 4642
rect 5143 4444 5199 4500
rect 5285 4444 5341 4500
rect 5143 4302 5199 4358
rect 5285 4302 5341 4358
rect 5143 4160 5199 4216
rect 5285 4160 5341 4216
rect 5143 4018 5199 4074
rect 5285 4018 5341 4074
rect 5143 3876 5199 3932
rect 5285 3876 5341 3932
rect 5143 3734 5199 3790
rect 5285 3734 5341 3790
rect 5143 3592 5199 3648
rect 5285 3592 5341 3648
rect 5143 3450 5199 3506
rect 5285 3450 5341 3506
rect 5143 3308 5199 3364
rect 5285 3308 5341 3364
rect 5143 3166 5199 3222
rect 5285 3166 5341 3222
rect 5143 3024 5199 3080
rect 5285 3024 5341 3080
rect 5143 2882 5199 2938
rect 5285 2882 5341 2938
rect 5143 2740 5199 2796
rect 5285 2740 5341 2796
rect 5143 2598 5199 2654
rect 5285 2598 5341 2654
rect 5143 2456 5199 2512
rect 5285 2456 5341 2512
rect 5143 2314 5199 2370
rect 5285 2314 5341 2370
rect 5143 2172 5199 2228
rect 5285 2172 5341 2228
rect 5143 2030 5199 2086
rect 5285 2030 5341 2086
rect 5143 1888 5199 1944
rect 5285 1888 5341 1944
rect 5143 1746 5199 1802
rect 5285 1746 5341 1802
rect 5143 1604 5199 1660
rect 5285 1604 5341 1660
rect 5143 1462 5199 1518
rect 5285 1462 5341 1518
rect 5143 1320 5199 1376
rect 5285 1320 5341 1376
rect 5143 1178 5199 1234
rect 5285 1178 5341 1234
rect 5143 1036 5199 1092
rect 5285 1036 5341 1092
rect 5143 894 5199 950
rect 5285 894 5341 950
rect 5143 752 5199 808
rect 5285 752 5341 808
rect 5143 610 5199 666
rect 5285 610 5341 666
rect 5143 468 5199 524
rect 5285 468 5341 524
rect 5540 12254 5596 12310
rect 5682 12254 5738 12310
rect 5540 12112 5596 12168
rect 5682 12112 5738 12168
rect 5540 11970 5596 12026
rect 5682 11970 5738 12026
rect 5540 11828 5596 11884
rect 5682 11828 5738 11884
rect 5540 11686 5596 11742
rect 5682 11686 5738 11742
rect 5540 11544 5596 11600
rect 5682 11544 5738 11600
rect 5540 11402 5596 11458
rect 5682 11402 5738 11458
rect 5540 11260 5596 11316
rect 5682 11260 5738 11316
rect 5540 11118 5596 11174
rect 5682 11118 5738 11174
rect 5540 10976 5596 11032
rect 5682 10976 5738 11032
rect 5540 10834 5596 10890
rect 5682 10834 5738 10890
rect 5540 10692 5596 10748
rect 5682 10692 5738 10748
rect 5540 10550 5596 10606
rect 5682 10550 5738 10606
rect 5540 10408 5596 10464
rect 5682 10408 5738 10464
rect 5540 10266 5596 10322
rect 5682 10266 5738 10322
rect 5540 10124 5596 10180
rect 5682 10124 5738 10180
rect 5540 9982 5596 10038
rect 5682 9982 5738 10038
rect 5540 9840 5596 9896
rect 5682 9840 5738 9896
rect 5540 9698 5596 9754
rect 5682 9698 5738 9754
rect 5540 9556 5596 9612
rect 5682 9556 5738 9612
rect 5540 9414 5596 9470
rect 5682 9414 5738 9470
rect 5540 9272 5596 9328
rect 5682 9272 5738 9328
rect 5540 9130 5596 9186
rect 5682 9130 5738 9186
rect 5540 8988 5596 9044
rect 5682 8988 5738 9044
rect 5540 8846 5596 8902
rect 5682 8846 5738 8902
rect 5540 8704 5596 8760
rect 5682 8704 5738 8760
rect 5540 8562 5596 8618
rect 5682 8562 5738 8618
rect 5540 8420 5596 8476
rect 5682 8420 5738 8476
rect 5540 8278 5596 8334
rect 5682 8278 5738 8334
rect 5540 8136 5596 8192
rect 5682 8136 5738 8192
rect 5540 7994 5596 8050
rect 5682 7994 5738 8050
rect 5540 7852 5596 7908
rect 5682 7852 5738 7908
rect 5540 7710 5596 7766
rect 5682 7710 5738 7766
rect 5540 7568 5596 7624
rect 5682 7568 5738 7624
rect 5540 7426 5596 7482
rect 5682 7426 5738 7482
rect 5540 7284 5596 7340
rect 5682 7284 5738 7340
rect 5540 7142 5596 7198
rect 5682 7142 5738 7198
rect 5540 7000 5596 7056
rect 5682 7000 5738 7056
rect 5540 6858 5596 6914
rect 5682 6858 5738 6914
rect 5540 6716 5596 6772
rect 5682 6716 5738 6772
rect 5540 6574 5596 6630
rect 5682 6574 5738 6630
rect 5540 6432 5596 6488
rect 5682 6432 5738 6488
rect 5540 6290 5596 6346
rect 5682 6290 5738 6346
rect 5540 6148 5596 6204
rect 5682 6148 5738 6204
rect 5540 6006 5596 6062
rect 5682 6006 5738 6062
rect 5540 5864 5596 5920
rect 5682 5864 5738 5920
rect 5540 5722 5596 5778
rect 5682 5722 5738 5778
rect 5540 5580 5596 5636
rect 5682 5580 5738 5636
rect 5540 5438 5596 5494
rect 5682 5438 5738 5494
rect 5540 5296 5596 5352
rect 5682 5296 5738 5352
rect 5540 5154 5596 5210
rect 5682 5154 5738 5210
rect 5540 5012 5596 5068
rect 5682 5012 5738 5068
rect 5540 4870 5596 4926
rect 5682 4870 5738 4926
rect 5540 4728 5596 4784
rect 5682 4728 5738 4784
rect 5540 4586 5596 4642
rect 5682 4586 5738 4642
rect 5540 4444 5596 4500
rect 5682 4444 5738 4500
rect 5540 4302 5596 4358
rect 5682 4302 5738 4358
rect 5540 4160 5596 4216
rect 5682 4160 5738 4216
rect 5540 4018 5596 4074
rect 5682 4018 5738 4074
rect 5540 3876 5596 3932
rect 5682 3876 5738 3932
rect 5540 3734 5596 3790
rect 5682 3734 5738 3790
rect 5540 3592 5596 3648
rect 5682 3592 5738 3648
rect 5540 3450 5596 3506
rect 5682 3450 5738 3506
rect 5540 3308 5596 3364
rect 5682 3308 5738 3364
rect 5540 3166 5596 3222
rect 5682 3166 5738 3222
rect 5540 3024 5596 3080
rect 5682 3024 5738 3080
rect 5540 2882 5596 2938
rect 5682 2882 5738 2938
rect 5540 2740 5596 2796
rect 5682 2740 5738 2796
rect 5540 2598 5596 2654
rect 5682 2598 5738 2654
rect 5540 2456 5596 2512
rect 5682 2456 5738 2512
rect 5540 2314 5596 2370
rect 5682 2314 5738 2370
rect 5540 2172 5596 2228
rect 5682 2172 5738 2228
rect 5540 2030 5596 2086
rect 5682 2030 5738 2086
rect 5540 1888 5596 1944
rect 5682 1888 5738 1944
rect 5540 1746 5596 1802
rect 5682 1746 5738 1802
rect 5540 1604 5596 1660
rect 5682 1604 5738 1660
rect 5540 1462 5596 1518
rect 5682 1462 5738 1518
rect 5540 1320 5596 1376
rect 5682 1320 5738 1376
rect 5540 1178 5596 1234
rect 5682 1178 5738 1234
rect 5540 1036 5596 1092
rect 5682 1036 5738 1092
rect 5540 894 5596 950
rect 5682 894 5738 950
rect 5540 752 5596 808
rect 5682 752 5738 808
rect 5540 610 5596 666
rect 5682 610 5738 666
rect 5540 468 5596 524
rect 5682 468 5738 524
rect 5937 12254 5993 12310
rect 6079 12254 6135 12310
rect 5937 12112 5993 12168
rect 6079 12112 6135 12168
rect 5937 11970 5993 12026
rect 6079 11970 6135 12026
rect 5937 11828 5993 11884
rect 6079 11828 6135 11884
rect 5937 11686 5993 11742
rect 6079 11686 6135 11742
rect 5937 11544 5993 11600
rect 6079 11544 6135 11600
rect 5937 11402 5993 11458
rect 6079 11402 6135 11458
rect 5937 11260 5993 11316
rect 6079 11260 6135 11316
rect 5937 11118 5993 11174
rect 6079 11118 6135 11174
rect 5937 10976 5993 11032
rect 6079 10976 6135 11032
rect 5937 10834 5993 10890
rect 6079 10834 6135 10890
rect 5937 10692 5993 10748
rect 6079 10692 6135 10748
rect 5937 10550 5993 10606
rect 6079 10550 6135 10606
rect 5937 10408 5993 10464
rect 6079 10408 6135 10464
rect 5937 10266 5993 10322
rect 6079 10266 6135 10322
rect 5937 10124 5993 10180
rect 6079 10124 6135 10180
rect 5937 9982 5993 10038
rect 6079 9982 6135 10038
rect 5937 9840 5993 9896
rect 6079 9840 6135 9896
rect 5937 9698 5993 9754
rect 6079 9698 6135 9754
rect 5937 9556 5993 9612
rect 6079 9556 6135 9612
rect 5937 9414 5993 9470
rect 6079 9414 6135 9470
rect 5937 9272 5993 9328
rect 6079 9272 6135 9328
rect 5937 9130 5993 9186
rect 6079 9130 6135 9186
rect 5937 8988 5993 9044
rect 6079 8988 6135 9044
rect 5937 8846 5993 8902
rect 6079 8846 6135 8902
rect 5937 8704 5993 8760
rect 6079 8704 6135 8760
rect 5937 8562 5993 8618
rect 6079 8562 6135 8618
rect 5937 8420 5993 8476
rect 6079 8420 6135 8476
rect 5937 8278 5993 8334
rect 6079 8278 6135 8334
rect 5937 8136 5993 8192
rect 6079 8136 6135 8192
rect 5937 7994 5993 8050
rect 6079 7994 6135 8050
rect 5937 7852 5993 7908
rect 6079 7852 6135 7908
rect 5937 7710 5993 7766
rect 6079 7710 6135 7766
rect 5937 7568 5993 7624
rect 6079 7568 6135 7624
rect 5937 7426 5993 7482
rect 6079 7426 6135 7482
rect 5937 7284 5993 7340
rect 6079 7284 6135 7340
rect 5937 7142 5993 7198
rect 6079 7142 6135 7198
rect 5937 7000 5993 7056
rect 6079 7000 6135 7056
rect 5937 6858 5993 6914
rect 6079 6858 6135 6914
rect 5937 6716 5993 6772
rect 6079 6716 6135 6772
rect 5937 6574 5993 6630
rect 6079 6574 6135 6630
rect 5937 6432 5993 6488
rect 6079 6432 6135 6488
rect 5937 6290 5993 6346
rect 6079 6290 6135 6346
rect 5937 6148 5993 6204
rect 6079 6148 6135 6204
rect 5937 6006 5993 6062
rect 6079 6006 6135 6062
rect 5937 5864 5993 5920
rect 6079 5864 6135 5920
rect 5937 5722 5993 5778
rect 6079 5722 6135 5778
rect 5937 5580 5993 5636
rect 6079 5580 6135 5636
rect 5937 5438 5993 5494
rect 6079 5438 6135 5494
rect 5937 5296 5993 5352
rect 6079 5296 6135 5352
rect 5937 5154 5993 5210
rect 6079 5154 6135 5210
rect 5937 5012 5993 5068
rect 6079 5012 6135 5068
rect 5937 4870 5993 4926
rect 6079 4870 6135 4926
rect 5937 4728 5993 4784
rect 6079 4728 6135 4784
rect 5937 4586 5993 4642
rect 6079 4586 6135 4642
rect 5937 4444 5993 4500
rect 6079 4444 6135 4500
rect 5937 4302 5993 4358
rect 6079 4302 6135 4358
rect 5937 4160 5993 4216
rect 6079 4160 6135 4216
rect 5937 4018 5993 4074
rect 6079 4018 6135 4074
rect 5937 3876 5993 3932
rect 6079 3876 6135 3932
rect 5937 3734 5993 3790
rect 6079 3734 6135 3790
rect 5937 3592 5993 3648
rect 6079 3592 6135 3648
rect 5937 3450 5993 3506
rect 6079 3450 6135 3506
rect 5937 3308 5993 3364
rect 6079 3308 6135 3364
rect 5937 3166 5993 3222
rect 6079 3166 6135 3222
rect 5937 3024 5993 3080
rect 6079 3024 6135 3080
rect 5937 2882 5993 2938
rect 6079 2882 6135 2938
rect 5937 2740 5993 2796
rect 6079 2740 6135 2796
rect 5937 2598 5993 2654
rect 6079 2598 6135 2654
rect 5937 2456 5993 2512
rect 6079 2456 6135 2512
rect 5937 2314 5993 2370
rect 6079 2314 6135 2370
rect 5937 2172 5993 2228
rect 6079 2172 6135 2228
rect 5937 2030 5993 2086
rect 6079 2030 6135 2086
rect 5937 1888 5993 1944
rect 6079 1888 6135 1944
rect 5937 1746 5993 1802
rect 6079 1746 6135 1802
rect 5937 1604 5993 1660
rect 6079 1604 6135 1660
rect 5937 1462 5993 1518
rect 6079 1462 6135 1518
rect 5937 1320 5993 1376
rect 6079 1320 6135 1376
rect 5937 1178 5993 1234
rect 6079 1178 6135 1234
rect 5937 1036 5993 1092
rect 6079 1036 6135 1092
rect 5937 894 5993 950
rect 6079 894 6135 950
rect 5937 752 5993 808
rect 6079 752 6135 808
rect 5937 610 5993 666
rect 6079 610 6135 666
rect 5937 468 5993 524
rect 6079 468 6135 524
rect 6340 12254 6396 12310
rect 6482 12254 6538 12310
rect 6340 12112 6396 12168
rect 6482 12112 6538 12168
rect 6340 11970 6396 12026
rect 6482 11970 6538 12026
rect 6340 11828 6396 11884
rect 6482 11828 6538 11884
rect 6340 11686 6396 11742
rect 6482 11686 6538 11742
rect 6340 11544 6396 11600
rect 6482 11544 6538 11600
rect 6340 11402 6396 11458
rect 6482 11402 6538 11458
rect 6340 11260 6396 11316
rect 6482 11260 6538 11316
rect 6340 11118 6396 11174
rect 6482 11118 6538 11174
rect 6340 10976 6396 11032
rect 6482 10976 6538 11032
rect 6340 10834 6396 10890
rect 6482 10834 6538 10890
rect 6340 10692 6396 10748
rect 6482 10692 6538 10748
rect 6340 10550 6396 10606
rect 6482 10550 6538 10606
rect 6340 10408 6396 10464
rect 6482 10408 6538 10464
rect 6340 10266 6396 10322
rect 6482 10266 6538 10322
rect 6340 10124 6396 10180
rect 6482 10124 6538 10180
rect 6340 9982 6396 10038
rect 6482 9982 6538 10038
rect 6340 9840 6396 9896
rect 6482 9840 6538 9896
rect 6340 9698 6396 9754
rect 6482 9698 6538 9754
rect 6340 9556 6396 9612
rect 6482 9556 6538 9612
rect 6340 9414 6396 9470
rect 6482 9414 6538 9470
rect 6340 9272 6396 9328
rect 6482 9272 6538 9328
rect 6340 9130 6396 9186
rect 6482 9130 6538 9186
rect 6340 8988 6396 9044
rect 6482 8988 6538 9044
rect 6340 8846 6396 8902
rect 6482 8846 6538 8902
rect 6340 8704 6396 8760
rect 6482 8704 6538 8760
rect 6340 8562 6396 8618
rect 6482 8562 6538 8618
rect 6340 8420 6396 8476
rect 6482 8420 6538 8476
rect 6340 8278 6396 8334
rect 6482 8278 6538 8334
rect 6340 8136 6396 8192
rect 6482 8136 6538 8192
rect 6340 7994 6396 8050
rect 6482 7994 6538 8050
rect 6340 7852 6396 7908
rect 6482 7852 6538 7908
rect 6340 7710 6396 7766
rect 6482 7710 6538 7766
rect 6340 7568 6396 7624
rect 6482 7568 6538 7624
rect 6340 7426 6396 7482
rect 6482 7426 6538 7482
rect 6340 7284 6396 7340
rect 6482 7284 6538 7340
rect 6340 7142 6396 7198
rect 6482 7142 6538 7198
rect 6340 7000 6396 7056
rect 6482 7000 6538 7056
rect 6340 6858 6396 6914
rect 6482 6858 6538 6914
rect 6340 6716 6396 6772
rect 6482 6716 6538 6772
rect 6340 6574 6396 6630
rect 6482 6574 6538 6630
rect 6340 6432 6396 6488
rect 6482 6432 6538 6488
rect 6340 6290 6396 6346
rect 6482 6290 6538 6346
rect 6340 6148 6396 6204
rect 6482 6148 6538 6204
rect 6340 6006 6396 6062
rect 6482 6006 6538 6062
rect 6340 5864 6396 5920
rect 6482 5864 6538 5920
rect 6340 5722 6396 5778
rect 6482 5722 6538 5778
rect 6340 5580 6396 5636
rect 6482 5580 6538 5636
rect 6340 5438 6396 5494
rect 6482 5438 6538 5494
rect 6340 5296 6396 5352
rect 6482 5296 6538 5352
rect 6340 5154 6396 5210
rect 6482 5154 6538 5210
rect 6340 5012 6396 5068
rect 6482 5012 6538 5068
rect 6340 4870 6396 4926
rect 6482 4870 6538 4926
rect 6340 4728 6396 4784
rect 6482 4728 6538 4784
rect 6340 4586 6396 4642
rect 6482 4586 6538 4642
rect 6340 4444 6396 4500
rect 6482 4444 6538 4500
rect 6340 4302 6396 4358
rect 6482 4302 6538 4358
rect 6340 4160 6396 4216
rect 6482 4160 6538 4216
rect 6340 4018 6396 4074
rect 6482 4018 6538 4074
rect 6340 3876 6396 3932
rect 6482 3876 6538 3932
rect 6340 3734 6396 3790
rect 6482 3734 6538 3790
rect 6340 3592 6396 3648
rect 6482 3592 6538 3648
rect 6340 3450 6396 3506
rect 6482 3450 6538 3506
rect 6340 3308 6396 3364
rect 6482 3308 6538 3364
rect 6340 3166 6396 3222
rect 6482 3166 6538 3222
rect 6340 3024 6396 3080
rect 6482 3024 6538 3080
rect 6340 2882 6396 2938
rect 6482 2882 6538 2938
rect 6340 2740 6396 2796
rect 6482 2740 6538 2796
rect 6340 2598 6396 2654
rect 6482 2598 6538 2654
rect 6340 2456 6396 2512
rect 6482 2456 6538 2512
rect 6340 2314 6396 2370
rect 6482 2314 6538 2370
rect 6340 2172 6396 2228
rect 6482 2172 6538 2228
rect 6340 2030 6396 2086
rect 6482 2030 6538 2086
rect 6340 1888 6396 1944
rect 6482 1888 6538 1944
rect 6340 1746 6396 1802
rect 6482 1746 6538 1802
rect 6340 1604 6396 1660
rect 6482 1604 6538 1660
rect 6340 1462 6396 1518
rect 6482 1462 6538 1518
rect 6340 1320 6396 1376
rect 6482 1320 6538 1376
rect 6340 1178 6396 1234
rect 6482 1178 6538 1234
rect 6340 1036 6396 1092
rect 6482 1036 6538 1092
rect 6340 894 6396 950
rect 6482 894 6538 950
rect 6340 752 6396 808
rect 6482 752 6538 808
rect 6340 610 6396 666
rect 6482 610 6538 666
rect 6340 468 6396 524
rect 6482 468 6538 524
rect 6742 12254 6798 12310
rect 6884 12254 6940 12310
rect 6742 12112 6798 12168
rect 6884 12112 6940 12168
rect 6742 11970 6798 12026
rect 6884 11970 6940 12026
rect 6742 11828 6798 11884
rect 6884 11828 6940 11884
rect 6742 11686 6798 11742
rect 6884 11686 6940 11742
rect 6742 11544 6798 11600
rect 6884 11544 6940 11600
rect 6742 11402 6798 11458
rect 6884 11402 6940 11458
rect 6742 11260 6798 11316
rect 6884 11260 6940 11316
rect 6742 11118 6798 11174
rect 6884 11118 6940 11174
rect 6742 10976 6798 11032
rect 6884 10976 6940 11032
rect 6742 10834 6798 10890
rect 6884 10834 6940 10890
rect 6742 10692 6798 10748
rect 6884 10692 6940 10748
rect 6742 10550 6798 10606
rect 6884 10550 6940 10606
rect 6742 10408 6798 10464
rect 6884 10408 6940 10464
rect 6742 10266 6798 10322
rect 6884 10266 6940 10322
rect 6742 10124 6798 10180
rect 6884 10124 6940 10180
rect 6742 9982 6798 10038
rect 6884 9982 6940 10038
rect 6742 9840 6798 9896
rect 6884 9840 6940 9896
rect 6742 9698 6798 9754
rect 6884 9698 6940 9754
rect 6742 9556 6798 9612
rect 6884 9556 6940 9612
rect 6742 9414 6798 9470
rect 6884 9414 6940 9470
rect 6742 9272 6798 9328
rect 6884 9272 6940 9328
rect 6742 9130 6798 9186
rect 6884 9130 6940 9186
rect 6742 8988 6798 9044
rect 6884 8988 6940 9044
rect 6742 8846 6798 8902
rect 6884 8846 6940 8902
rect 6742 8704 6798 8760
rect 6884 8704 6940 8760
rect 6742 8562 6798 8618
rect 6884 8562 6940 8618
rect 6742 8420 6798 8476
rect 6884 8420 6940 8476
rect 6742 8278 6798 8334
rect 6884 8278 6940 8334
rect 6742 8136 6798 8192
rect 6884 8136 6940 8192
rect 6742 7994 6798 8050
rect 6884 7994 6940 8050
rect 6742 7852 6798 7908
rect 6884 7852 6940 7908
rect 6742 7710 6798 7766
rect 6884 7710 6940 7766
rect 6742 7568 6798 7624
rect 6884 7568 6940 7624
rect 6742 7426 6798 7482
rect 6884 7426 6940 7482
rect 6742 7284 6798 7340
rect 6884 7284 6940 7340
rect 6742 7142 6798 7198
rect 6884 7142 6940 7198
rect 6742 7000 6798 7056
rect 6884 7000 6940 7056
rect 6742 6858 6798 6914
rect 6884 6858 6940 6914
rect 6742 6716 6798 6772
rect 6884 6716 6940 6772
rect 6742 6574 6798 6630
rect 6884 6574 6940 6630
rect 6742 6432 6798 6488
rect 6884 6432 6940 6488
rect 6742 6290 6798 6346
rect 6884 6290 6940 6346
rect 6742 6148 6798 6204
rect 6884 6148 6940 6204
rect 6742 6006 6798 6062
rect 6884 6006 6940 6062
rect 6742 5864 6798 5920
rect 6884 5864 6940 5920
rect 6742 5722 6798 5778
rect 6884 5722 6940 5778
rect 6742 5580 6798 5636
rect 6884 5580 6940 5636
rect 6742 5438 6798 5494
rect 6884 5438 6940 5494
rect 6742 5296 6798 5352
rect 6884 5296 6940 5352
rect 6742 5154 6798 5210
rect 6884 5154 6940 5210
rect 6742 5012 6798 5068
rect 6884 5012 6940 5068
rect 6742 4870 6798 4926
rect 6884 4870 6940 4926
rect 6742 4728 6798 4784
rect 6884 4728 6940 4784
rect 6742 4586 6798 4642
rect 6884 4586 6940 4642
rect 6742 4444 6798 4500
rect 6884 4444 6940 4500
rect 6742 4302 6798 4358
rect 6884 4302 6940 4358
rect 6742 4160 6798 4216
rect 6884 4160 6940 4216
rect 6742 4018 6798 4074
rect 6884 4018 6940 4074
rect 6742 3876 6798 3932
rect 6884 3876 6940 3932
rect 6742 3734 6798 3790
rect 6884 3734 6940 3790
rect 6742 3592 6798 3648
rect 6884 3592 6940 3648
rect 6742 3450 6798 3506
rect 6884 3450 6940 3506
rect 6742 3308 6798 3364
rect 6884 3308 6940 3364
rect 6742 3166 6798 3222
rect 6884 3166 6940 3222
rect 6742 3024 6798 3080
rect 6884 3024 6940 3080
rect 6742 2882 6798 2938
rect 6884 2882 6940 2938
rect 6742 2740 6798 2796
rect 6884 2740 6940 2796
rect 6742 2598 6798 2654
rect 6884 2598 6940 2654
rect 6742 2456 6798 2512
rect 6884 2456 6940 2512
rect 6742 2314 6798 2370
rect 6884 2314 6940 2370
rect 6742 2172 6798 2228
rect 6884 2172 6940 2228
rect 6742 2030 6798 2086
rect 6884 2030 6940 2086
rect 6742 1888 6798 1944
rect 6884 1888 6940 1944
rect 6742 1746 6798 1802
rect 6884 1746 6940 1802
rect 6742 1604 6798 1660
rect 6884 1604 6940 1660
rect 6742 1462 6798 1518
rect 6884 1462 6940 1518
rect 6742 1320 6798 1376
rect 6884 1320 6940 1376
rect 6742 1178 6798 1234
rect 6884 1178 6940 1234
rect 6742 1036 6798 1092
rect 6884 1036 6940 1092
rect 6742 894 6798 950
rect 6884 894 6940 950
rect 6742 752 6798 808
rect 6884 752 6940 808
rect 6742 610 6798 666
rect 6884 610 6940 666
rect 6742 468 6798 524
rect 6884 468 6940 524
rect 7145 12254 7201 12310
rect 7287 12254 7343 12310
rect 7145 12112 7201 12168
rect 7287 12112 7343 12168
rect 7145 11970 7201 12026
rect 7287 11970 7343 12026
rect 7145 11828 7201 11884
rect 7287 11828 7343 11884
rect 7145 11686 7201 11742
rect 7287 11686 7343 11742
rect 7145 11544 7201 11600
rect 7287 11544 7343 11600
rect 7145 11402 7201 11458
rect 7287 11402 7343 11458
rect 7145 11260 7201 11316
rect 7287 11260 7343 11316
rect 7145 11118 7201 11174
rect 7287 11118 7343 11174
rect 7145 10976 7201 11032
rect 7287 10976 7343 11032
rect 7145 10834 7201 10890
rect 7287 10834 7343 10890
rect 7145 10692 7201 10748
rect 7287 10692 7343 10748
rect 7145 10550 7201 10606
rect 7287 10550 7343 10606
rect 7145 10408 7201 10464
rect 7287 10408 7343 10464
rect 7145 10266 7201 10322
rect 7287 10266 7343 10322
rect 7145 10124 7201 10180
rect 7287 10124 7343 10180
rect 7145 9982 7201 10038
rect 7287 9982 7343 10038
rect 7145 9840 7201 9896
rect 7287 9840 7343 9896
rect 7145 9698 7201 9754
rect 7287 9698 7343 9754
rect 7145 9556 7201 9612
rect 7287 9556 7343 9612
rect 7145 9414 7201 9470
rect 7287 9414 7343 9470
rect 7145 9272 7201 9328
rect 7287 9272 7343 9328
rect 7145 9130 7201 9186
rect 7287 9130 7343 9186
rect 7145 8988 7201 9044
rect 7287 8988 7343 9044
rect 7145 8846 7201 8902
rect 7287 8846 7343 8902
rect 7145 8704 7201 8760
rect 7287 8704 7343 8760
rect 7145 8562 7201 8618
rect 7287 8562 7343 8618
rect 7145 8420 7201 8476
rect 7287 8420 7343 8476
rect 7145 8278 7201 8334
rect 7287 8278 7343 8334
rect 7145 8136 7201 8192
rect 7287 8136 7343 8192
rect 7145 7994 7201 8050
rect 7287 7994 7343 8050
rect 7145 7852 7201 7908
rect 7287 7852 7343 7908
rect 7145 7710 7201 7766
rect 7287 7710 7343 7766
rect 7145 7568 7201 7624
rect 7287 7568 7343 7624
rect 7145 7426 7201 7482
rect 7287 7426 7343 7482
rect 7145 7284 7201 7340
rect 7287 7284 7343 7340
rect 7145 7142 7201 7198
rect 7287 7142 7343 7198
rect 7145 7000 7201 7056
rect 7287 7000 7343 7056
rect 7145 6858 7201 6914
rect 7287 6858 7343 6914
rect 7145 6716 7201 6772
rect 7287 6716 7343 6772
rect 7145 6574 7201 6630
rect 7287 6574 7343 6630
rect 7145 6432 7201 6488
rect 7287 6432 7343 6488
rect 7145 6290 7201 6346
rect 7287 6290 7343 6346
rect 7145 6148 7201 6204
rect 7287 6148 7343 6204
rect 7145 6006 7201 6062
rect 7287 6006 7343 6062
rect 7145 5864 7201 5920
rect 7287 5864 7343 5920
rect 7145 5722 7201 5778
rect 7287 5722 7343 5778
rect 7145 5580 7201 5636
rect 7287 5580 7343 5636
rect 7145 5438 7201 5494
rect 7287 5438 7343 5494
rect 7145 5296 7201 5352
rect 7287 5296 7343 5352
rect 7145 5154 7201 5210
rect 7287 5154 7343 5210
rect 7145 5012 7201 5068
rect 7287 5012 7343 5068
rect 7145 4870 7201 4926
rect 7287 4870 7343 4926
rect 7145 4728 7201 4784
rect 7287 4728 7343 4784
rect 7145 4586 7201 4642
rect 7287 4586 7343 4642
rect 7145 4444 7201 4500
rect 7287 4444 7343 4500
rect 7145 4302 7201 4358
rect 7287 4302 7343 4358
rect 7145 4160 7201 4216
rect 7287 4160 7343 4216
rect 7145 4018 7201 4074
rect 7287 4018 7343 4074
rect 7145 3876 7201 3932
rect 7287 3876 7343 3932
rect 7145 3734 7201 3790
rect 7287 3734 7343 3790
rect 7145 3592 7201 3648
rect 7287 3592 7343 3648
rect 7145 3450 7201 3506
rect 7287 3450 7343 3506
rect 7145 3308 7201 3364
rect 7287 3308 7343 3364
rect 7145 3166 7201 3222
rect 7287 3166 7343 3222
rect 7145 3024 7201 3080
rect 7287 3024 7343 3080
rect 7145 2882 7201 2938
rect 7287 2882 7343 2938
rect 7145 2740 7201 2796
rect 7287 2740 7343 2796
rect 7145 2598 7201 2654
rect 7287 2598 7343 2654
rect 7145 2456 7201 2512
rect 7287 2456 7343 2512
rect 7145 2314 7201 2370
rect 7287 2314 7343 2370
rect 7145 2172 7201 2228
rect 7287 2172 7343 2228
rect 7145 2030 7201 2086
rect 7287 2030 7343 2086
rect 7145 1888 7201 1944
rect 7287 1888 7343 1944
rect 7145 1746 7201 1802
rect 7287 1746 7343 1802
rect 7145 1604 7201 1660
rect 7287 1604 7343 1660
rect 7145 1462 7201 1518
rect 7287 1462 7343 1518
rect 7145 1320 7201 1376
rect 7287 1320 7343 1376
rect 7145 1178 7201 1234
rect 7287 1178 7343 1234
rect 7145 1036 7201 1092
rect 7287 1036 7343 1092
rect 7145 894 7201 950
rect 7287 894 7343 950
rect 7145 752 7201 808
rect 7287 752 7343 808
rect 7145 610 7201 666
rect 7287 610 7343 666
rect 7145 468 7201 524
rect 7287 468 7343 524
rect 7539 12254 7595 12310
rect 7681 12254 7737 12310
rect 7539 12112 7595 12168
rect 7681 12112 7737 12168
rect 7539 11970 7595 12026
rect 7681 11970 7737 12026
rect 7539 11828 7595 11884
rect 7681 11828 7737 11884
rect 7539 11686 7595 11742
rect 7681 11686 7737 11742
rect 7539 11544 7595 11600
rect 7681 11544 7737 11600
rect 7539 11402 7595 11458
rect 7681 11402 7737 11458
rect 7539 11260 7595 11316
rect 7681 11260 7737 11316
rect 7539 11118 7595 11174
rect 7681 11118 7737 11174
rect 7539 10976 7595 11032
rect 7681 10976 7737 11032
rect 7539 10834 7595 10890
rect 7681 10834 7737 10890
rect 7539 10692 7595 10748
rect 7681 10692 7737 10748
rect 7539 10550 7595 10606
rect 7681 10550 7737 10606
rect 7539 10408 7595 10464
rect 7681 10408 7737 10464
rect 7539 10266 7595 10322
rect 7681 10266 7737 10322
rect 7539 10124 7595 10180
rect 7681 10124 7737 10180
rect 7539 9982 7595 10038
rect 7681 9982 7737 10038
rect 7539 9840 7595 9896
rect 7681 9840 7737 9896
rect 7539 9698 7595 9754
rect 7681 9698 7737 9754
rect 7539 9556 7595 9612
rect 7681 9556 7737 9612
rect 7539 9414 7595 9470
rect 7681 9414 7737 9470
rect 7539 9272 7595 9328
rect 7681 9272 7737 9328
rect 7539 9130 7595 9186
rect 7681 9130 7737 9186
rect 7539 8988 7595 9044
rect 7681 8988 7737 9044
rect 7539 8846 7595 8902
rect 7681 8846 7737 8902
rect 7539 8704 7595 8760
rect 7681 8704 7737 8760
rect 7539 8562 7595 8618
rect 7681 8562 7737 8618
rect 7539 8420 7595 8476
rect 7681 8420 7737 8476
rect 7539 8278 7595 8334
rect 7681 8278 7737 8334
rect 7539 8136 7595 8192
rect 7681 8136 7737 8192
rect 7539 7994 7595 8050
rect 7681 7994 7737 8050
rect 7539 7852 7595 7908
rect 7681 7852 7737 7908
rect 7539 7710 7595 7766
rect 7681 7710 7737 7766
rect 7539 7568 7595 7624
rect 7681 7568 7737 7624
rect 7539 7426 7595 7482
rect 7681 7426 7737 7482
rect 7539 7284 7595 7340
rect 7681 7284 7737 7340
rect 7539 7142 7595 7198
rect 7681 7142 7737 7198
rect 7539 7000 7595 7056
rect 7681 7000 7737 7056
rect 7539 6858 7595 6914
rect 7681 6858 7737 6914
rect 7539 6716 7595 6772
rect 7681 6716 7737 6772
rect 7539 6574 7595 6630
rect 7681 6574 7737 6630
rect 7539 6432 7595 6488
rect 7681 6432 7737 6488
rect 7539 6290 7595 6346
rect 7681 6290 7737 6346
rect 7539 6148 7595 6204
rect 7681 6148 7737 6204
rect 7539 6006 7595 6062
rect 7681 6006 7737 6062
rect 7539 5864 7595 5920
rect 7681 5864 7737 5920
rect 7539 5722 7595 5778
rect 7681 5722 7737 5778
rect 7539 5580 7595 5636
rect 7681 5580 7737 5636
rect 7539 5438 7595 5494
rect 7681 5438 7737 5494
rect 7539 5296 7595 5352
rect 7681 5296 7737 5352
rect 7539 5154 7595 5210
rect 7681 5154 7737 5210
rect 7539 5012 7595 5068
rect 7681 5012 7737 5068
rect 7539 4870 7595 4926
rect 7681 4870 7737 4926
rect 7539 4728 7595 4784
rect 7681 4728 7737 4784
rect 7539 4586 7595 4642
rect 7681 4586 7737 4642
rect 7539 4444 7595 4500
rect 7681 4444 7737 4500
rect 7539 4302 7595 4358
rect 7681 4302 7737 4358
rect 7539 4160 7595 4216
rect 7681 4160 7737 4216
rect 7539 4018 7595 4074
rect 7681 4018 7737 4074
rect 7539 3876 7595 3932
rect 7681 3876 7737 3932
rect 7539 3734 7595 3790
rect 7681 3734 7737 3790
rect 7539 3592 7595 3648
rect 7681 3592 7737 3648
rect 7539 3450 7595 3506
rect 7681 3450 7737 3506
rect 7539 3308 7595 3364
rect 7681 3308 7737 3364
rect 7539 3166 7595 3222
rect 7681 3166 7737 3222
rect 7539 3024 7595 3080
rect 7681 3024 7737 3080
rect 7539 2882 7595 2938
rect 7681 2882 7737 2938
rect 7539 2740 7595 2796
rect 7681 2740 7737 2796
rect 7539 2598 7595 2654
rect 7681 2598 7737 2654
rect 7539 2456 7595 2512
rect 7681 2456 7737 2512
rect 7539 2314 7595 2370
rect 7681 2314 7737 2370
rect 7539 2172 7595 2228
rect 7681 2172 7737 2228
rect 7539 2030 7595 2086
rect 7681 2030 7737 2086
rect 7539 1888 7595 1944
rect 7681 1888 7737 1944
rect 7539 1746 7595 1802
rect 7681 1746 7737 1802
rect 7539 1604 7595 1660
rect 7681 1604 7737 1660
rect 7539 1462 7595 1518
rect 7681 1462 7737 1518
rect 7539 1320 7595 1376
rect 7681 1320 7737 1376
rect 7539 1178 7595 1234
rect 7681 1178 7737 1234
rect 7539 1036 7595 1092
rect 7681 1036 7737 1092
rect 7539 894 7595 950
rect 7681 894 7737 950
rect 7539 752 7595 808
rect 7681 752 7737 808
rect 7539 610 7595 666
rect 7681 610 7737 666
rect 7539 468 7595 524
rect 7681 468 7737 524
rect 7940 12254 7996 12310
rect 8082 12254 8138 12310
rect 7940 12112 7996 12168
rect 8082 12112 8138 12168
rect 7940 11970 7996 12026
rect 8082 11970 8138 12026
rect 7940 11828 7996 11884
rect 8082 11828 8138 11884
rect 7940 11686 7996 11742
rect 8082 11686 8138 11742
rect 7940 11544 7996 11600
rect 8082 11544 8138 11600
rect 7940 11402 7996 11458
rect 8082 11402 8138 11458
rect 7940 11260 7996 11316
rect 8082 11260 8138 11316
rect 7940 11118 7996 11174
rect 8082 11118 8138 11174
rect 7940 10976 7996 11032
rect 8082 10976 8138 11032
rect 7940 10834 7996 10890
rect 8082 10834 8138 10890
rect 7940 10692 7996 10748
rect 8082 10692 8138 10748
rect 7940 10550 7996 10606
rect 8082 10550 8138 10606
rect 7940 10408 7996 10464
rect 8082 10408 8138 10464
rect 7940 10266 7996 10322
rect 8082 10266 8138 10322
rect 7940 10124 7996 10180
rect 8082 10124 8138 10180
rect 7940 9982 7996 10038
rect 8082 9982 8138 10038
rect 7940 9840 7996 9896
rect 8082 9840 8138 9896
rect 7940 9698 7996 9754
rect 8082 9698 8138 9754
rect 7940 9556 7996 9612
rect 8082 9556 8138 9612
rect 7940 9414 7996 9470
rect 8082 9414 8138 9470
rect 7940 9272 7996 9328
rect 8082 9272 8138 9328
rect 7940 9130 7996 9186
rect 8082 9130 8138 9186
rect 7940 8988 7996 9044
rect 8082 8988 8138 9044
rect 7940 8846 7996 8902
rect 8082 8846 8138 8902
rect 7940 8704 7996 8760
rect 8082 8704 8138 8760
rect 7940 8562 7996 8618
rect 8082 8562 8138 8618
rect 7940 8420 7996 8476
rect 8082 8420 8138 8476
rect 7940 8278 7996 8334
rect 8082 8278 8138 8334
rect 7940 8136 7996 8192
rect 8082 8136 8138 8192
rect 7940 7994 7996 8050
rect 8082 7994 8138 8050
rect 7940 7852 7996 7908
rect 8082 7852 8138 7908
rect 7940 7710 7996 7766
rect 8082 7710 8138 7766
rect 7940 7568 7996 7624
rect 8082 7568 8138 7624
rect 7940 7426 7996 7482
rect 8082 7426 8138 7482
rect 7940 7284 7996 7340
rect 8082 7284 8138 7340
rect 7940 7142 7996 7198
rect 8082 7142 8138 7198
rect 7940 7000 7996 7056
rect 8082 7000 8138 7056
rect 7940 6858 7996 6914
rect 8082 6858 8138 6914
rect 7940 6716 7996 6772
rect 8082 6716 8138 6772
rect 7940 6574 7996 6630
rect 8082 6574 8138 6630
rect 7940 6432 7996 6488
rect 8082 6432 8138 6488
rect 7940 6290 7996 6346
rect 8082 6290 8138 6346
rect 7940 6148 7996 6204
rect 8082 6148 8138 6204
rect 7940 6006 7996 6062
rect 8082 6006 8138 6062
rect 7940 5864 7996 5920
rect 8082 5864 8138 5920
rect 7940 5722 7996 5778
rect 8082 5722 8138 5778
rect 7940 5580 7996 5636
rect 8082 5580 8138 5636
rect 7940 5438 7996 5494
rect 8082 5438 8138 5494
rect 7940 5296 7996 5352
rect 8082 5296 8138 5352
rect 7940 5154 7996 5210
rect 8082 5154 8138 5210
rect 7940 5012 7996 5068
rect 8082 5012 8138 5068
rect 7940 4870 7996 4926
rect 8082 4870 8138 4926
rect 7940 4728 7996 4784
rect 8082 4728 8138 4784
rect 7940 4586 7996 4642
rect 8082 4586 8138 4642
rect 7940 4444 7996 4500
rect 8082 4444 8138 4500
rect 7940 4302 7996 4358
rect 8082 4302 8138 4358
rect 7940 4160 7996 4216
rect 8082 4160 8138 4216
rect 7940 4018 7996 4074
rect 8082 4018 8138 4074
rect 7940 3876 7996 3932
rect 8082 3876 8138 3932
rect 7940 3734 7996 3790
rect 8082 3734 8138 3790
rect 7940 3592 7996 3648
rect 8082 3592 8138 3648
rect 7940 3450 7996 3506
rect 8082 3450 8138 3506
rect 7940 3308 7996 3364
rect 8082 3308 8138 3364
rect 7940 3166 7996 3222
rect 8082 3166 8138 3222
rect 7940 3024 7996 3080
rect 8082 3024 8138 3080
rect 7940 2882 7996 2938
rect 8082 2882 8138 2938
rect 7940 2740 7996 2796
rect 8082 2740 8138 2796
rect 7940 2598 7996 2654
rect 8082 2598 8138 2654
rect 7940 2456 7996 2512
rect 8082 2456 8138 2512
rect 7940 2314 7996 2370
rect 8082 2314 8138 2370
rect 7940 2172 7996 2228
rect 8082 2172 8138 2228
rect 7940 2030 7996 2086
rect 8082 2030 8138 2086
rect 7940 1888 7996 1944
rect 8082 1888 8138 1944
rect 7940 1746 7996 1802
rect 8082 1746 8138 1802
rect 7940 1604 7996 1660
rect 8082 1604 8138 1660
rect 7940 1462 7996 1518
rect 8082 1462 8138 1518
rect 7940 1320 7996 1376
rect 8082 1320 8138 1376
rect 7940 1178 7996 1234
rect 8082 1178 8138 1234
rect 7940 1036 7996 1092
rect 8082 1036 8138 1092
rect 7940 894 7996 950
rect 8082 894 8138 950
rect 7940 752 7996 808
rect 8082 752 8138 808
rect 7940 610 7996 666
rect 8082 610 8138 666
rect 7940 468 7996 524
rect 8082 468 8138 524
rect 8340 12254 8396 12310
rect 8482 12254 8538 12310
rect 8340 12112 8396 12168
rect 8482 12112 8538 12168
rect 8340 11970 8396 12026
rect 8482 11970 8538 12026
rect 8340 11828 8396 11884
rect 8482 11828 8538 11884
rect 8340 11686 8396 11742
rect 8482 11686 8538 11742
rect 8340 11544 8396 11600
rect 8482 11544 8538 11600
rect 8340 11402 8396 11458
rect 8482 11402 8538 11458
rect 8340 11260 8396 11316
rect 8482 11260 8538 11316
rect 8340 11118 8396 11174
rect 8482 11118 8538 11174
rect 8340 10976 8396 11032
rect 8482 10976 8538 11032
rect 8340 10834 8396 10890
rect 8482 10834 8538 10890
rect 8340 10692 8396 10748
rect 8482 10692 8538 10748
rect 8340 10550 8396 10606
rect 8482 10550 8538 10606
rect 8340 10408 8396 10464
rect 8482 10408 8538 10464
rect 8340 10266 8396 10322
rect 8482 10266 8538 10322
rect 8340 10124 8396 10180
rect 8482 10124 8538 10180
rect 8340 9982 8396 10038
rect 8482 9982 8538 10038
rect 8340 9840 8396 9896
rect 8482 9840 8538 9896
rect 8340 9698 8396 9754
rect 8482 9698 8538 9754
rect 8340 9556 8396 9612
rect 8482 9556 8538 9612
rect 8340 9414 8396 9470
rect 8482 9414 8538 9470
rect 8340 9272 8396 9328
rect 8482 9272 8538 9328
rect 8340 9130 8396 9186
rect 8482 9130 8538 9186
rect 8340 8988 8396 9044
rect 8482 8988 8538 9044
rect 8340 8846 8396 8902
rect 8482 8846 8538 8902
rect 8340 8704 8396 8760
rect 8482 8704 8538 8760
rect 8340 8562 8396 8618
rect 8482 8562 8538 8618
rect 8340 8420 8396 8476
rect 8482 8420 8538 8476
rect 8340 8278 8396 8334
rect 8482 8278 8538 8334
rect 8340 8136 8396 8192
rect 8482 8136 8538 8192
rect 8340 7994 8396 8050
rect 8482 7994 8538 8050
rect 8340 7852 8396 7908
rect 8482 7852 8538 7908
rect 8340 7710 8396 7766
rect 8482 7710 8538 7766
rect 8340 7568 8396 7624
rect 8482 7568 8538 7624
rect 8340 7426 8396 7482
rect 8482 7426 8538 7482
rect 8340 7284 8396 7340
rect 8482 7284 8538 7340
rect 8340 7142 8396 7198
rect 8482 7142 8538 7198
rect 8340 7000 8396 7056
rect 8482 7000 8538 7056
rect 8340 6858 8396 6914
rect 8482 6858 8538 6914
rect 8340 6716 8396 6772
rect 8482 6716 8538 6772
rect 8340 6574 8396 6630
rect 8482 6574 8538 6630
rect 8340 6432 8396 6488
rect 8482 6432 8538 6488
rect 8340 6290 8396 6346
rect 8482 6290 8538 6346
rect 8340 6148 8396 6204
rect 8482 6148 8538 6204
rect 8340 6006 8396 6062
rect 8482 6006 8538 6062
rect 8340 5864 8396 5920
rect 8482 5864 8538 5920
rect 8340 5722 8396 5778
rect 8482 5722 8538 5778
rect 8340 5580 8396 5636
rect 8482 5580 8538 5636
rect 8340 5438 8396 5494
rect 8482 5438 8538 5494
rect 8340 5296 8396 5352
rect 8482 5296 8538 5352
rect 8340 5154 8396 5210
rect 8482 5154 8538 5210
rect 8340 5012 8396 5068
rect 8482 5012 8538 5068
rect 8340 4870 8396 4926
rect 8482 4870 8538 4926
rect 8340 4728 8396 4784
rect 8482 4728 8538 4784
rect 8340 4586 8396 4642
rect 8482 4586 8538 4642
rect 8340 4444 8396 4500
rect 8482 4444 8538 4500
rect 8340 4302 8396 4358
rect 8482 4302 8538 4358
rect 8340 4160 8396 4216
rect 8482 4160 8538 4216
rect 8340 4018 8396 4074
rect 8482 4018 8538 4074
rect 8340 3876 8396 3932
rect 8482 3876 8538 3932
rect 8340 3734 8396 3790
rect 8482 3734 8538 3790
rect 8340 3592 8396 3648
rect 8482 3592 8538 3648
rect 8340 3450 8396 3506
rect 8482 3450 8538 3506
rect 8340 3308 8396 3364
rect 8482 3308 8538 3364
rect 8340 3166 8396 3222
rect 8482 3166 8538 3222
rect 8340 3024 8396 3080
rect 8482 3024 8538 3080
rect 8340 2882 8396 2938
rect 8482 2882 8538 2938
rect 8340 2740 8396 2796
rect 8482 2740 8538 2796
rect 8340 2598 8396 2654
rect 8482 2598 8538 2654
rect 8340 2456 8396 2512
rect 8482 2456 8538 2512
rect 8340 2314 8396 2370
rect 8482 2314 8538 2370
rect 8340 2172 8396 2228
rect 8482 2172 8538 2228
rect 8340 2030 8396 2086
rect 8482 2030 8538 2086
rect 8340 1888 8396 1944
rect 8482 1888 8538 1944
rect 8340 1746 8396 1802
rect 8482 1746 8538 1802
rect 8340 1604 8396 1660
rect 8482 1604 8538 1660
rect 8340 1462 8396 1518
rect 8482 1462 8538 1518
rect 8340 1320 8396 1376
rect 8482 1320 8538 1376
rect 8340 1178 8396 1234
rect 8482 1178 8538 1234
rect 8340 1036 8396 1092
rect 8482 1036 8538 1092
rect 8340 894 8396 950
rect 8482 894 8538 950
rect 8340 752 8396 808
rect 8482 752 8538 808
rect 8340 610 8396 666
rect 8482 610 8538 666
rect 8340 468 8396 524
rect 8482 468 8538 524
rect 8737 12254 8793 12310
rect 8879 12254 8935 12310
rect 8737 12112 8793 12168
rect 8879 12112 8935 12168
rect 8737 11970 8793 12026
rect 8879 11970 8935 12026
rect 8737 11828 8793 11884
rect 8879 11828 8935 11884
rect 8737 11686 8793 11742
rect 8879 11686 8935 11742
rect 8737 11544 8793 11600
rect 8879 11544 8935 11600
rect 8737 11402 8793 11458
rect 8879 11402 8935 11458
rect 8737 11260 8793 11316
rect 8879 11260 8935 11316
rect 8737 11118 8793 11174
rect 8879 11118 8935 11174
rect 8737 10976 8793 11032
rect 8879 10976 8935 11032
rect 8737 10834 8793 10890
rect 8879 10834 8935 10890
rect 8737 10692 8793 10748
rect 8879 10692 8935 10748
rect 8737 10550 8793 10606
rect 8879 10550 8935 10606
rect 8737 10408 8793 10464
rect 8879 10408 8935 10464
rect 8737 10266 8793 10322
rect 8879 10266 8935 10322
rect 8737 10124 8793 10180
rect 8879 10124 8935 10180
rect 8737 9982 8793 10038
rect 8879 9982 8935 10038
rect 8737 9840 8793 9896
rect 8879 9840 8935 9896
rect 8737 9698 8793 9754
rect 8879 9698 8935 9754
rect 8737 9556 8793 9612
rect 8879 9556 8935 9612
rect 8737 9414 8793 9470
rect 8879 9414 8935 9470
rect 8737 9272 8793 9328
rect 8879 9272 8935 9328
rect 8737 9130 8793 9186
rect 8879 9130 8935 9186
rect 8737 8988 8793 9044
rect 8879 8988 8935 9044
rect 8737 8846 8793 8902
rect 8879 8846 8935 8902
rect 8737 8704 8793 8760
rect 8879 8704 8935 8760
rect 8737 8562 8793 8618
rect 8879 8562 8935 8618
rect 8737 8420 8793 8476
rect 8879 8420 8935 8476
rect 8737 8278 8793 8334
rect 8879 8278 8935 8334
rect 8737 8136 8793 8192
rect 8879 8136 8935 8192
rect 8737 7994 8793 8050
rect 8879 7994 8935 8050
rect 8737 7852 8793 7908
rect 8879 7852 8935 7908
rect 8737 7710 8793 7766
rect 8879 7710 8935 7766
rect 8737 7568 8793 7624
rect 8879 7568 8935 7624
rect 8737 7426 8793 7482
rect 8879 7426 8935 7482
rect 8737 7284 8793 7340
rect 8879 7284 8935 7340
rect 8737 7142 8793 7198
rect 8879 7142 8935 7198
rect 8737 7000 8793 7056
rect 8879 7000 8935 7056
rect 8737 6858 8793 6914
rect 8879 6858 8935 6914
rect 8737 6716 8793 6772
rect 8879 6716 8935 6772
rect 8737 6574 8793 6630
rect 8879 6574 8935 6630
rect 8737 6432 8793 6488
rect 8879 6432 8935 6488
rect 8737 6290 8793 6346
rect 8879 6290 8935 6346
rect 8737 6148 8793 6204
rect 8879 6148 8935 6204
rect 8737 6006 8793 6062
rect 8879 6006 8935 6062
rect 8737 5864 8793 5920
rect 8879 5864 8935 5920
rect 8737 5722 8793 5778
rect 8879 5722 8935 5778
rect 8737 5580 8793 5636
rect 8879 5580 8935 5636
rect 8737 5438 8793 5494
rect 8879 5438 8935 5494
rect 8737 5296 8793 5352
rect 8879 5296 8935 5352
rect 8737 5154 8793 5210
rect 8879 5154 8935 5210
rect 8737 5012 8793 5068
rect 8879 5012 8935 5068
rect 8737 4870 8793 4926
rect 8879 4870 8935 4926
rect 8737 4728 8793 4784
rect 8879 4728 8935 4784
rect 8737 4586 8793 4642
rect 8879 4586 8935 4642
rect 8737 4444 8793 4500
rect 8879 4444 8935 4500
rect 8737 4302 8793 4358
rect 8879 4302 8935 4358
rect 8737 4160 8793 4216
rect 8879 4160 8935 4216
rect 8737 4018 8793 4074
rect 8879 4018 8935 4074
rect 8737 3876 8793 3932
rect 8879 3876 8935 3932
rect 8737 3734 8793 3790
rect 8879 3734 8935 3790
rect 8737 3592 8793 3648
rect 8879 3592 8935 3648
rect 8737 3450 8793 3506
rect 8879 3450 8935 3506
rect 8737 3308 8793 3364
rect 8879 3308 8935 3364
rect 8737 3166 8793 3222
rect 8879 3166 8935 3222
rect 8737 3024 8793 3080
rect 8879 3024 8935 3080
rect 8737 2882 8793 2938
rect 8879 2882 8935 2938
rect 8737 2740 8793 2796
rect 8879 2740 8935 2796
rect 8737 2598 8793 2654
rect 8879 2598 8935 2654
rect 8737 2456 8793 2512
rect 8879 2456 8935 2512
rect 8737 2314 8793 2370
rect 8879 2314 8935 2370
rect 8737 2172 8793 2228
rect 8879 2172 8935 2228
rect 8737 2030 8793 2086
rect 8879 2030 8935 2086
rect 8737 1888 8793 1944
rect 8879 1888 8935 1944
rect 8737 1746 8793 1802
rect 8879 1746 8935 1802
rect 8737 1604 8793 1660
rect 8879 1604 8935 1660
rect 8737 1462 8793 1518
rect 8879 1462 8935 1518
rect 8737 1320 8793 1376
rect 8879 1320 8935 1376
rect 8737 1178 8793 1234
rect 8879 1178 8935 1234
rect 8737 1036 8793 1092
rect 8879 1036 8935 1092
rect 8737 894 8793 950
rect 8879 894 8935 950
rect 8737 752 8793 808
rect 8879 752 8935 808
rect 8737 610 8793 666
rect 8879 610 8935 666
rect 8737 468 8793 524
rect 8879 468 8935 524
rect 9134 12254 9190 12310
rect 9276 12254 9332 12310
rect 9134 12112 9190 12168
rect 9276 12112 9332 12168
rect 9134 11970 9190 12026
rect 9276 11970 9332 12026
rect 9134 11828 9190 11884
rect 9276 11828 9332 11884
rect 9134 11686 9190 11742
rect 9276 11686 9332 11742
rect 9134 11544 9190 11600
rect 9276 11544 9332 11600
rect 9134 11402 9190 11458
rect 9276 11402 9332 11458
rect 9134 11260 9190 11316
rect 9276 11260 9332 11316
rect 9134 11118 9190 11174
rect 9276 11118 9332 11174
rect 9134 10976 9190 11032
rect 9276 10976 9332 11032
rect 9134 10834 9190 10890
rect 9276 10834 9332 10890
rect 9134 10692 9190 10748
rect 9276 10692 9332 10748
rect 9134 10550 9190 10606
rect 9276 10550 9332 10606
rect 9134 10408 9190 10464
rect 9276 10408 9332 10464
rect 9134 10266 9190 10322
rect 9276 10266 9332 10322
rect 9134 10124 9190 10180
rect 9276 10124 9332 10180
rect 9134 9982 9190 10038
rect 9276 9982 9332 10038
rect 9134 9840 9190 9896
rect 9276 9840 9332 9896
rect 9134 9698 9190 9754
rect 9276 9698 9332 9754
rect 9134 9556 9190 9612
rect 9276 9556 9332 9612
rect 9134 9414 9190 9470
rect 9276 9414 9332 9470
rect 9134 9272 9190 9328
rect 9276 9272 9332 9328
rect 9134 9130 9190 9186
rect 9276 9130 9332 9186
rect 9134 8988 9190 9044
rect 9276 8988 9332 9044
rect 9134 8846 9190 8902
rect 9276 8846 9332 8902
rect 9134 8704 9190 8760
rect 9276 8704 9332 8760
rect 9134 8562 9190 8618
rect 9276 8562 9332 8618
rect 9134 8420 9190 8476
rect 9276 8420 9332 8476
rect 9134 8278 9190 8334
rect 9276 8278 9332 8334
rect 9134 8136 9190 8192
rect 9276 8136 9332 8192
rect 9134 7994 9190 8050
rect 9276 7994 9332 8050
rect 9134 7852 9190 7908
rect 9276 7852 9332 7908
rect 9134 7710 9190 7766
rect 9276 7710 9332 7766
rect 9134 7568 9190 7624
rect 9276 7568 9332 7624
rect 9134 7426 9190 7482
rect 9276 7426 9332 7482
rect 9134 7284 9190 7340
rect 9276 7284 9332 7340
rect 9134 7142 9190 7198
rect 9276 7142 9332 7198
rect 9134 7000 9190 7056
rect 9276 7000 9332 7056
rect 9134 6858 9190 6914
rect 9276 6858 9332 6914
rect 9134 6716 9190 6772
rect 9276 6716 9332 6772
rect 9134 6574 9190 6630
rect 9276 6574 9332 6630
rect 9134 6432 9190 6488
rect 9276 6432 9332 6488
rect 9134 6290 9190 6346
rect 9276 6290 9332 6346
rect 9134 6148 9190 6204
rect 9276 6148 9332 6204
rect 9134 6006 9190 6062
rect 9276 6006 9332 6062
rect 9134 5864 9190 5920
rect 9276 5864 9332 5920
rect 9134 5722 9190 5778
rect 9276 5722 9332 5778
rect 9134 5580 9190 5636
rect 9276 5580 9332 5636
rect 9134 5438 9190 5494
rect 9276 5438 9332 5494
rect 9134 5296 9190 5352
rect 9276 5296 9332 5352
rect 9134 5154 9190 5210
rect 9276 5154 9332 5210
rect 9134 5012 9190 5068
rect 9276 5012 9332 5068
rect 9134 4870 9190 4926
rect 9276 4870 9332 4926
rect 9134 4728 9190 4784
rect 9276 4728 9332 4784
rect 9134 4586 9190 4642
rect 9276 4586 9332 4642
rect 9134 4444 9190 4500
rect 9276 4444 9332 4500
rect 9134 4302 9190 4358
rect 9276 4302 9332 4358
rect 9134 4160 9190 4216
rect 9276 4160 9332 4216
rect 9134 4018 9190 4074
rect 9276 4018 9332 4074
rect 9134 3876 9190 3932
rect 9276 3876 9332 3932
rect 9134 3734 9190 3790
rect 9276 3734 9332 3790
rect 9134 3592 9190 3648
rect 9276 3592 9332 3648
rect 9134 3450 9190 3506
rect 9276 3450 9332 3506
rect 9134 3308 9190 3364
rect 9276 3308 9332 3364
rect 9134 3166 9190 3222
rect 9276 3166 9332 3222
rect 9134 3024 9190 3080
rect 9276 3024 9332 3080
rect 9134 2882 9190 2938
rect 9276 2882 9332 2938
rect 9134 2740 9190 2796
rect 9276 2740 9332 2796
rect 9134 2598 9190 2654
rect 9276 2598 9332 2654
rect 9134 2456 9190 2512
rect 9276 2456 9332 2512
rect 9134 2314 9190 2370
rect 9276 2314 9332 2370
rect 9134 2172 9190 2228
rect 9276 2172 9332 2228
rect 9134 2030 9190 2086
rect 9276 2030 9332 2086
rect 9134 1888 9190 1944
rect 9276 1888 9332 1944
rect 9134 1746 9190 1802
rect 9276 1746 9332 1802
rect 9134 1604 9190 1660
rect 9276 1604 9332 1660
rect 9134 1462 9190 1518
rect 9276 1462 9332 1518
rect 9134 1320 9190 1376
rect 9276 1320 9332 1376
rect 9134 1178 9190 1234
rect 9276 1178 9332 1234
rect 9134 1036 9190 1092
rect 9276 1036 9332 1092
rect 9134 894 9190 950
rect 9276 894 9332 950
rect 9134 752 9190 808
rect 9276 752 9332 808
rect 9134 610 9190 666
rect 9276 610 9332 666
rect 9134 468 9190 524
rect 9276 468 9332 524
rect 9538 12254 9594 12310
rect 9680 12254 9736 12310
rect 9538 12112 9594 12168
rect 9680 12112 9736 12168
rect 9538 11970 9594 12026
rect 9680 11970 9736 12026
rect 9538 11828 9594 11884
rect 9680 11828 9736 11884
rect 9538 11686 9594 11742
rect 9680 11686 9736 11742
rect 9538 11544 9594 11600
rect 9680 11544 9736 11600
rect 9538 11402 9594 11458
rect 9680 11402 9736 11458
rect 9538 11260 9594 11316
rect 9680 11260 9736 11316
rect 9538 11118 9594 11174
rect 9680 11118 9736 11174
rect 9538 10976 9594 11032
rect 9680 10976 9736 11032
rect 9538 10834 9594 10890
rect 9680 10834 9736 10890
rect 9538 10692 9594 10748
rect 9680 10692 9736 10748
rect 9538 10550 9594 10606
rect 9680 10550 9736 10606
rect 9538 10408 9594 10464
rect 9680 10408 9736 10464
rect 9538 10266 9594 10322
rect 9680 10266 9736 10322
rect 9538 10124 9594 10180
rect 9680 10124 9736 10180
rect 9538 9982 9594 10038
rect 9680 9982 9736 10038
rect 9538 9840 9594 9896
rect 9680 9840 9736 9896
rect 9538 9698 9594 9754
rect 9680 9698 9736 9754
rect 9538 9556 9594 9612
rect 9680 9556 9736 9612
rect 9538 9414 9594 9470
rect 9680 9414 9736 9470
rect 9538 9272 9594 9328
rect 9680 9272 9736 9328
rect 9538 9130 9594 9186
rect 9680 9130 9736 9186
rect 9538 8988 9594 9044
rect 9680 8988 9736 9044
rect 9538 8846 9594 8902
rect 9680 8846 9736 8902
rect 9538 8704 9594 8760
rect 9680 8704 9736 8760
rect 9538 8562 9594 8618
rect 9680 8562 9736 8618
rect 9538 8420 9594 8476
rect 9680 8420 9736 8476
rect 9538 8278 9594 8334
rect 9680 8278 9736 8334
rect 9538 8136 9594 8192
rect 9680 8136 9736 8192
rect 9538 7994 9594 8050
rect 9680 7994 9736 8050
rect 9538 7852 9594 7908
rect 9680 7852 9736 7908
rect 9538 7710 9594 7766
rect 9680 7710 9736 7766
rect 9538 7568 9594 7624
rect 9680 7568 9736 7624
rect 9538 7426 9594 7482
rect 9680 7426 9736 7482
rect 9538 7284 9594 7340
rect 9680 7284 9736 7340
rect 9538 7142 9594 7198
rect 9680 7142 9736 7198
rect 9538 7000 9594 7056
rect 9680 7000 9736 7056
rect 9538 6858 9594 6914
rect 9680 6858 9736 6914
rect 9538 6716 9594 6772
rect 9680 6716 9736 6772
rect 9538 6574 9594 6630
rect 9680 6574 9736 6630
rect 9538 6432 9594 6488
rect 9680 6432 9736 6488
rect 9538 6290 9594 6346
rect 9680 6290 9736 6346
rect 9538 6148 9594 6204
rect 9680 6148 9736 6204
rect 9538 6006 9594 6062
rect 9680 6006 9736 6062
rect 9538 5864 9594 5920
rect 9680 5864 9736 5920
rect 9538 5722 9594 5778
rect 9680 5722 9736 5778
rect 9538 5580 9594 5636
rect 9680 5580 9736 5636
rect 9538 5438 9594 5494
rect 9680 5438 9736 5494
rect 9538 5296 9594 5352
rect 9680 5296 9736 5352
rect 9538 5154 9594 5210
rect 9680 5154 9736 5210
rect 9538 5012 9594 5068
rect 9680 5012 9736 5068
rect 9538 4870 9594 4926
rect 9680 4870 9736 4926
rect 9538 4728 9594 4784
rect 9680 4728 9736 4784
rect 9538 4586 9594 4642
rect 9680 4586 9736 4642
rect 9538 4444 9594 4500
rect 9680 4444 9736 4500
rect 9538 4302 9594 4358
rect 9680 4302 9736 4358
rect 9538 4160 9594 4216
rect 9680 4160 9736 4216
rect 9538 4018 9594 4074
rect 9680 4018 9736 4074
rect 9538 3876 9594 3932
rect 9680 3876 9736 3932
rect 9538 3734 9594 3790
rect 9680 3734 9736 3790
rect 9538 3592 9594 3648
rect 9680 3592 9736 3648
rect 9538 3450 9594 3506
rect 9680 3450 9736 3506
rect 9538 3308 9594 3364
rect 9680 3308 9736 3364
rect 9538 3166 9594 3222
rect 9680 3166 9736 3222
rect 9538 3024 9594 3080
rect 9680 3024 9736 3080
rect 9538 2882 9594 2938
rect 9680 2882 9736 2938
rect 9538 2740 9594 2796
rect 9680 2740 9736 2796
rect 9538 2598 9594 2654
rect 9680 2598 9736 2654
rect 9538 2456 9594 2512
rect 9680 2456 9736 2512
rect 9538 2314 9594 2370
rect 9680 2314 9736 2370
rect 9538 2172 9594 2228
rect 9680 2172 9736 2228
rect 9538 2030 9594 2086
rect 9680 2030 9736 2086
rect 9538 1888 9594 1944
rect 9680 1888 9736 1944
rect 9538 1746 9594 1802
rect 9680 1746 9736 1802
rect 9538 1604 9594 1660
rect 9680 1604 9736 1660
rect 9538 1462 9594 1518
rect 9680 1462 9736 1518
rect 9538 1320 9594 1376
rect 9680 1320 9736 1376
rect 9538 1178 9594 1234
rect 9680 1178 9736 1234
rect 9538 1036 9594 1092
rect 9680 1036 9736 1092
rect 9538 894 9594 950
rect 9680 894 9736 950
rect 9538 752 9594 808
rect 9680 752 9736 808
rect 9538 610 9594 666
rect 9680 610 9736 666
rect 9538 468 9594 524
rect 9680 468 9736 524
rect 9934 12254 9990 12310
rect 10076 12254 10132 12310
rect 9934 12112 9990 12168
rect 10076 12112 10132 12168
rect 9934 11970 9990 12026
rect 10076 11970 10132 12026
rect 9934 11828 9990 11884
rect 10076 11828 10132 11884
rect 9934 11686 9990 11742
rect 10076 11686 10132 11742
rect 9934 11544 9990 11600
rect 10076 11544 10132 11600
rect 9934 11402 9990 11458
rect 10076 11402 10132 11458
rect 9934 11260 9990 11316
rect 10076 11260 10132 11316
rect 9934 11118 9990 11174
rect 10076 11118 10132 11174
rect 9934 10976 9990 11032
rect 10076 10976 10132 11032
rect 9934 10834 9990 10890
rect 10076 10834 10132 10890
rect 9934 10692 9990 10748
rect 10076 10692 10132 10748
rect 9934 10550 9990 10606
rect 10076 10550 10132 10606
rect 9934 10408 9990 10464
rect 10076 10408 10132 10464
rect 9934 10266 9990 10322
rect 10076 10266 10132 10322
rect 9934 10124 9990 10180
rect 10076 10124 10132 10180
rect 9934 9982 9990 10038
rect 10076 9982 10132 10038
rect 9934 9840 9990 9896
rect 10076 9840 10132 9896
rect 9934 9698 9990 9754
rect 10076 9698 10132 9754
rect 9934 9556 9990 9612
rect 10076 9556 10132 9612
rect 9934 9414 9990 9470
rect 10076 9414 10132 9470
rect 9934 9272 9990 9328
rect 10076 9272 10132 9328
rect 9934 9130 9990 9186
rect 10076 9130 10132 9186
rect 9934 8988 9990 9044
rect 10076 8988 10132 9044
rect 9934 8846 9990 8902
rect 10076 8846 10132 8902
rect 9934 8704 9990 8760
rect 10076 8704 10132 8760
rect 9934 8562 9990 8618
rect 10076 8562 10132 8618
rect 9934 8420 9990 8476
rect 10076 8420 10132 8476
rect 9934 8278 9990 8334
rect 10076 8278 10132 8334
rect 9934 8136 9990 8192
rect 10076 8136 10132 8192
rect 9934 7994 9990 8050
rect 10076 7994 10132 8050
rect 9934 7852 9990 7908
rect 10076 7852 10132 7908
rect 9934 7710 9990 7766
rect 10076 7710 10132 7766
rect 9934 7568 9990 7624
rect 10076 7568 10132 7624
rect 9934 7426 9990 7482
rect 10076 7426 10132 7482
rect 9934 7284 9990 7340
rect 10076 7284 10132 7340
rect 9934 7142 9990 7198
rect 10076 7142 10132 7198
rect 9934 7000 9990 7056
rect 10076 7000 10132 7056
rect 9934 6858 9990 6914
rect 10076 6858 10132 6914
rect 9934 6716 9990 6772
rect 10076 6716 10132 6772
rect 9934 6574 9990 6630
rect 10076 6574 10132 6630
rect 9934 6432 9990 6488
rect 10076 6432 10132 6488
rect 9934 6290 9990 6346
rect 10076 6290 10132 6346
rect 9934 6148 9990 6204
rect 10076 6148 10132 6204
rect 9934 6006 9990 6062
rect 10076 6006 10132 6062
rect 9934 5864 9990 5920
rect 10076 5864 10132 5920
rect 9934 5722 9990 5778
rect 10076 5722 10132 5778
rect 9934 5580 9990 5636
rect 10076 5580 10132 5636
rect 9934 5438 9990 5494
rect 10076 5438 10132 5494
rect 9934 5296 9990 5352
rect 10076 5296 10132 5352
rect 9934 5154 9990 5210
rect 10076 5154 10132 5210
rect 9934 5012 9990 5068
rect 10076 5012 10132 5068
rect 9934 4870 9990 4926
rect 10076 4870 10132 4926
rect 9934 4728 9990 4784
rect 10076 4728 10132 4784
rect 9934 4586 9990 4642
rect 10076 4586 10132 4642
rect 9934 4444 9990 4500
rect 10076 4444 10132 4500
rect 9934 4302 9990 4358
rect 10076 4302 10132 4358
rect 9934 4160 9990 4216
rect 10076 4160 10132 4216
rect 9934 4018 9990 4074
rect 10076 4018 10132 4074
rect 9934 3876 9990 3932
rect 10076 3876 10132 3932
rect 9934 3734 9990 3790
rect 10076 3734 10132 3790
rect 9934 3592 9990 3648
rect 10076 3592 10132 3648
rect 9934 3450 9990 3506
rect 10076 3450 10132 3506
rect 9934 3308 9990 3364
rect 10076 3308 10132 3364
rect 9934 3166 9990 3222
rect 10076 3166 10132 3222
rect 9934 3024 9990 3080
rect 10076 3024 10132 3080
rect 9934 2882 9990 2938
rect 10076 2882 10132 2938
rect 9934 2740 9990 2796
rect 10076 2740 10132 2796
rect 9934 2598 9990 2654
rect 10076 2598 10132 2654
rect 9934 2456 9990 2512
rect 10076 2456 10132 2512
rect 9934 2314 9990 2370
rect 10076 2314 10132 2370
rect 9934 2172 9990 2228
rect 10076 2172 10132 2228
rect 9934 2030 9990 2086
rect 10076 2030 10132 2086
rect 9934 1888 9990 1944
rect 10076 1888 10132 1944
rect 9934 1746 9990 1802
rect 10076 1746 10132 1802
rect 9934 1604 9990 1660
rect 10076 1604 10132 1660
rect 9934 1462 9990 1518
rect 10076 1462 10132 1518
rect 9934 1320 9990 1376
rect 10076 1320 10132 1376
rect 9934 1178 9990 1234
rect 10076 1178 10132 1234
rect 9934 1036 9990 1092
rect 10076 1036 10132 1092
rect 9934 894 9990 950
rect 10076 894 10132 950
rect 9934 752 9990 808
rect 10076 752 10132 808
rect 9934 610 9990 666
rect 10076 610 10132 666
rect 9934 468 9990 524
rect 10076 468 10132 524
rect 10334 12254 10390 12310
rect 10476 12254 10532 12310
rect 10334 12112 10390 12168
rect 10476 12112 10532 12168
rect 10334 11970 10390 12026
rect 10476 11970 10532 12026
rect 10334 11828 10390 11884
rect 10476 11828 10532 11884
rect 10334 11686 10390 11742
rect 10476 11686 10532 11742
rect 10334 11544 10390 11600
rect 10476 11544 10532 11600
rect 10334 11402 10390 11458
rect 10476 11402 10532 11458
rect 10334 11260 10390 11316
rect 10476 11260 10532 11316
rect 10334 11118 10390 11174
rect 10476 11118 10532 11174
rect 10334 10976 10390 11032
rect 10476 10976 10532 11032
rect 10334 10834 10390 10890
rect 10476 10834 10532 10890
rect 10334 10692 10390 10748
rect 10476 10692 10532 10748
rect 10334 10550 10390 10606
rect 10476 10550 10532 10606
rect 10334 10408 10390 10464
rect 10476 10408 10532 10464
rect 10334 10266 10390 10322
rect 10476 10266 10532 10322
rect 10334 10124 10390 10180
rect 10476 10124 10532 10180
rect 10334 9982 10390 10038
rect 10476 9982 10532 10038
rect 10334 9840 10390 9896
rect 10476 9840 10532 9896
rect 10334 9698 10390 9754
rect 10476 9698 10532 9754
rect 10334 9556 10390 9612
rect 10476 9556 10532 9612
rect 10334 9414 10390 9470
rect 10476 9414 10532 9470
rect 10334 9272 10390 9328
rect 10476 9272 10532 9328
rect 10334 9130 10390 9186
rect 10476 9130 10532 9186
rect 10334 8988 10390 9044
rect 10476 8988 10532 9044
rect 10334 8846 10390 8902
rect 10476 8846 10532 8902
rect 10334 8704 10390 8760
rect 10476 8704 10532 8760
rect 10334 8562 10390 8618
rect 10476 8562 10532 8618
rect 10334 8420 10390 8476
rect 10476 8420 10532 8476
rect 10334 8278 10390 8334
rect 10476 8278 10532 8334
rect 10334 8136 10390 8192
rect 10476 8136 10532 8192
rect 10334 7994 10390 8050
rect 10476 7994 10532 8050
rect 10334 7852 10390 7908
rect 10476 7852 10532 7908
rect 10334 7710 10390 7766
rect 10476 7710 10532 7766
rect 10334 7568 10390 7624
rect 10476 7568 10532 7624
rect 10334 7426 10390 7482
rect 10476 7426 10532 7482
rect 10334 7284 10390 7340
rect 10476 7284 10532 7340
rect 10334 7142 10390 7198
rect 10476 7142 10532 7198
rect 10334 7000 10390 7056
rect 10476 7000 10532 7056
rect 10334 6858 10390 6914
rect 10476 6858 10532 6914
rect 10334 6716 10390 6772
rect 10476 6716 10532 6772
rect 10334 6574 10390 6630
rect 10476 6574 10532 6630
rect 10334 6432 10390 6488
rect 10476 6432 10532 6488
rect 10334 6290 10390 6346
rect 10476 6290 10532 6346
rect 10334 6148 10390 6204
rect 10476 6148 10532 6204
rect 10334 6006 10390 6062
rect 10476 6006 10532 6062
rect 10334 5864 10390 5920
rect 10476 5864 10532 5920
rect 10334 5722 10390 5778
rect 10476 5722 10532 5778
rect 10334 5580 10390 5636
rect 10476 5580 10532 5636
rect 10334 5438 10390 5494
rect 10476 5438 10532 5494
rect 10334 5296 10390 5352
rect 10476 5296 10532 5352
rect 10334 5154 10390 5210
rect 10476 5154 10532 5210
rect 10334 5012 10390 5068
rect 10476 5012 10532 5068
rect 10334 4870 10390 4926
rect 10476 4870 10532 4926
rect 10334 4728 10390 4784
rect 10476 4728 10532 4784
rect 10334 4586 10390 4642
rect 10476 4586 10532 4642
rect 10334 4444 10390 4500
rect 10476 4444 10532 4500
rect 10334 4302 10390 4358
rect 10476 4302 10532 4358
rect 10334 4160 10390 4216
rect 10476 4160 10532 4216
rect 10334 4018 10390 4074
rect 10476 4018 10532 4074
rect 10334 3876 10390 3932
rect 10476 3876 10532 3932
rect 10334 3734 10390 3790
rect 10476 3734 10532 3790
rect 10334 3592 10390 3648
rect 10476 3592 10532 3648
rect 10334 3450 10390 3506
rect 10476 3450 10532 3506
rect 10334 3308 10390 3364
rect 10476 3308 10532 3364
rect 10334 3166 10390 3222
rect 10476 3166 10532 3222
rect 10334 3024 10390 3080
rect 10476 3024 10532 3080
rect 10334 2882 10390 2938
rect 10476 2882 10532 2938
rect 10334 2740 10390 2796
rect 10476 2740 10532 2796
rect 10334 2598 10390 2654
rect 10476 2598 10532 2654
rect 10334 2456 10390 2512
rect 10476 2456 10532 2512
rect 10334 2314 10390 2370
rect 10476 2314 10532 2370
rect 10334 2172 10390 2228
rect 10476 2172 10532 2228
rect 10334 2030 10390 2086
rect 10476 2030 10532 2086
rect 10334 1888 10390 1944
rect 10476 1888 10532 1944
rect 10334 1746 10390 1802
rect 10476 1746 10532 1802
rect 10334 1604 10390 1660
rect 10476 1604 10532 1660
rect 10334 1462 10390 1518
rect 10476 1462 10532 1518
rect 10334 1320 10390 1376
rect 10476 1320 10532 1376
rect 10334 1178 10390 1234
rect 10476 1178 10532 1234
rect 10334 1036 10390 1092
rect 10476 1036 10532 1092
rect 10334 894 10390 950
rect 10476 894 10532 950
rect 10334 752 10390 808
rect 10476 752 10532 808
rect 10334 610 10390 666
rect 10476 610 10532 666
rect 10334 468 10390 524
rect 10476 468 10532 524
rect 10731 12254 10787 12310
rect 10873 12254 10929 12310
rect 10731 12112 10787 12168
rect 10873 12112 10929 12168
rect 10731 11970 10787 12026
rect 10873 11970 10929 12026
rect 10731 11828 10787 11884
rect 10873 11828 10929 11884
rect 10731 11686 10787 11742
rect 10873 11686 10929 11742
rect 10731 11544 10787 11600
rect 10873 11544 10929 11600
rect 10731 11402 10787 11458
rect 10873 11402 10929 11458
rect 10731 11260 10787 11316
rect 10873 11260 10929 11316
rect 10731 11118 10787 11174
rect 10873 11118 10929 11174
rect 10731 10976 10787 11032
rect 10873 10976 10929 11032
rect 10731 10834 10787 10890
rect 10873 10834 10929 10890
rect 10731 10692 10787 10748
rect 10873 10692 10929 10748
rect 10731 10550 10787 10606
rect 10873 10550 10929 10606
rect 10731 10408 10787 10464
rect 10873 10408 10929 10464
rect 10731 10266 10787 10322
rect 10873 10266 10929 10322
rect 10731 10124 10787 10180
rect 10873 10124 10929 10180
rect 10731 9982 10787 10038
rect 10873 9982 10929 10038
rect 10731 9840 10787 9896
rect 10873 9840 10929 9896
rect 10731 9698 10787 9754
rect 10873 9698 10929 9754
rect 10731 9556 10787 9612
rect 10873 9556 10929 9612
rect 10731 9414 10787 9470
rect 10873 9414 10929 9470
rect 10731 9272 10787 9328
rect 10873 9272 10929 9328
rect 10731 9130 10787 9186
rect 10873 9130 10929 9186
rect 10731 8988 10787 9044
rect 10873 8988 10929 9044
rect 10731 8846 10787 8902
rect 10873 8846 10929 8902
rect 10731 8704 10787 8760
rect 10873 8704 10929 8760
rect 10731 8562 10787 8618
rect 10873 8562 10929 8618
rect 10731 8420 10787 8476
rect 10873 8420 10929 8476
rect 10731 8278 10787 8334
rect 10873 8278 10929 8334
rect 10731 8136 10787 8192
rect 10873 8136 10929 8192
rect 10731 7994 10787 8050
rect 10873 7994 10929 8050
rect 10731 7852 10787 7908
rect 10873 7852 10929 7908
rect 10731 7710 10787 7766
rect 10873 7710 10929 7766
rect 10731 7568 10787 7624
rect 10873 7568 10929 7624
rect 10731 7426 10787 7482
rect 10873 7426 10929 7482
rect 10731 7284 10787 7340
rect 10873 7284 10929 7340
rect 10731 7142 10787 7198
rect 10873 7142 10929 7198
rect 10731 7000 10787 7056
rect 10873 7000 10929 7056
rect 10731 6858 10787 6914
rect 10873 6858 10929 6914
rect 10731 6716 10787 6772
rect 10873 6716 10929 6772
rect 10731 6574 10787 6630
rect 10873 6574 10929 6630
rect 10731 6432 10787 6488
rect 10873 6432 10929 6488
rect 10731 6290 10787 6346
rect 10873 6290 10929 6346
rect 10731 6148 10787 6204
rect 10873 6148 10929 6204
rect 10731 6006 10787 6062
rect 10873 6006 10929 6062
rect 10731 5864 10787 5920
rect 10873 5864 10929 5920
rect 10731 5722 10787 5778
rect 10873 5722 10929 5778
rect 10731 5580 10787 5636
rect 10873 5580 10929 5636
rect 10731 5438 10787 5494
rect 10873 5438 10929 5494
rect 10731 5296 10787 5352
rect 10873 5296 10929 5352
rect 10731 5154 10787 5210
rect 10873 5154 10929 5210
rect 10731 5012 10787 5068
rect 10873 5012 10929 5068
rect 10731 4870 10787 4926
rect 10873 4870 10929 4926
rect 10731 4728 10787 4784
rect 10873 4728 10929 4784
rect 10731 4586 10787 4642
rect 10873 4586 10929 4642
rect 10731 4444 10787 4500
rect 10873 4444 10929 4500
rect 10731 4302 10787 4358
rect 10873 4302 10929 4358
rect 10731 4160 10787 4216
rect 10873 4160 10929 4216
rect 10731 4018 10787 4074
rect 10873 4018 10929 4074
rect 10731 3876 10787 3932
rect 10873 3876 10929 3932
rect 10731 3734 10787 3790
rect 10873 3734 10929 3790
rect 10731 3592 10787 3648
rect 10873 3592 10929 3648
rect 10731 3450 10787 3506
rect 10873 3450 10929 3506
rect 10731 3308 10787 3364
rect 10873 3308 10929 3364
rect 10731 3166 10787 3222
rect 10873 3166 10929 3222
rect 10731 3024 10787 3080
rect 10873 3024 10929 3080
rect 10731 2882 10787 2938
rect 10873 2882 10929 2938
rect 10731 2740 10787 2796
rect 10873 2740 10929 2796
rect 10731 2598 10787 2654
rect 10873 2598 10929 2654
rect 10731 2456 10787 2512
rect 10873 2456 10929 2512
rect 10731 2314 10787 2370
rect 10873 2314 10929 2370
rect 10731 2172 10787 2228
rect 10873 2172 10929 2228
rect 10731 2030 10787 2086
rect 10873 2030 10929 2086
rect 10731 1888 10787 1944
rect 10873 1888 10929 1944
rect 10731 1746 10787 1802
rect 10873 1746 10929 1802
rect 10731 1604 10787 1660
rect 10873 1604 10929 1660
rect 10731 1462 10787 1518
rect 10873 1462 10929 1518
rect 10731 1320 10787 1376
rect 10873 1320 10929 1376
rect 10731 1178 10787 1234
rect 10873 1178 10929 1234
rect 10731 1036 10787 1092
rect 10873 1036 10929 1092
rect 10731 894 10787 950
rect 10873 894 10929 950
rect 10731 752 10787 808
rect 10873 752 10929 808
rect 10731 610 10787 666
rect 10873 610 10929 666
rect 10731 468 10787 524
rect 10873 468 10929 524
rect 11136 12254 11192 12310
rect 11278 12254 11334 12310
rect 11136 12112 11192 12168
rect 11278 12112 11334 12168
rect 11136 11970 11192 12026
rect 11278 11970 11334 12026
rect 11136 11828 11192 11884
rect 11278 11828 11334 11884
rect 11136 11686 11192 11742
rect 11278 11686 11334 11742
rect 11136 11544 11192 11600
rect 11278 11544 11334 11600
rect 11136 11402 11192 11458
rect 11278 11402 11334 11458
rect 11136 11260 11192 11316
rect 11278 11260 11334 11316
rect 11136 11118 11192 11174
rect 11278 11118 11334 11174
rect 11136 10976 11192 11032
rect 11278 10976 11334 11032
rect 11136 10834 11192 10890
rect 11278 10834 11334 10890
rect 11136 10692 11192 10748
rect 11278 10692 11334 10748
rect 11136 10550 11192 10606
rect 11278 10550 11334 10606
rect 11136 10408 11192 10464
rect 11278 10408 11334 10464
rect 11136 10266 11192 10322
rect 11278 10266 11334 10322
rect 11136 10124 11192 10180
rect 11278 10124 11334 10180
rect 11136 9982 11192 10038
rect 11278 9982 11334 10038
rect 11136 9840 11192 9896
rect 11278 9840 11334 9896
rect 11136 9698 11192 9754
rect 11278 9698 11334 9754
rect 11136 9556 11192 9612
rect 11278 9556 11334 9612
rect 11136 9414 11192 9470
rect 11278 9414 11334 9470
rect 11136 9272 11192 9328
rect 11278 9272 11334 9328
rect 11136 9130 11192 9186
rect 11278 9130 11334 9186
rect 11136 8988 11192 9044
rect 11278 8988 11334 9044
rect 11136 8846 11192 8902
rect 11278 8846 11334 8902
rect 11136 8704 11192 8760
rect 11278 8704 11334 8760
rect 11136 8562 11192 8618
rect 11278 8562 11334 8618
rect 11136 8420 11192 8476
rect 11278 8420 11334 8476
rect 11136 8278 11192 8334
rect 11278 8278 11334 8334
rect 11136 8136 11192 8192
rect 11278 8136 11334 8192
rect 11136 7994 11192 8050
rect 11278 7994 11334 8050
rect 11136 7852 11192 7908
rect 11278 7852 11334 7908
rect 11136 7710 11192 7766
rect 11278 7710 11334 7766
rect 11136 7568 11192 7624
rect 11278 7568 11334 7624
rect 11136 7426 11192 7482
rect 11278 7426 11334 7482
rect 11136 7284 11192 7340
rect 11278 7284 11334 7340
rect 11136 7142 11192 7198
rect 11278 7142 11334 7198
rect 11136 7000 11192 7056
rect 11278 7000 11334 7056
rect 11136 6858 11192 6914
rect 11278 6858 11334 6914
rect 11136 6716 11192 6772
rect 11278 6716 11334 6772
rect 11136 6574 11192 6630
rect 11278 6574 11334 6630
rect 11136 6432 11192 6488
rect 11278 6432 11334 6488
rect 11136 6290 11192 6346
rect 11278 6290 11334 6346
rect 11136 6148 11192 6204
rect 11278 6148 11334 6204
rect 11136 6006 11192 6062
rect 11278 6006 11334 6062
rect 11136 5864 11192 5920
rect 11278 5864 11334 5920
rect 11136 5722 11192 5778
rect 11278 5722 11334 5778
rect 11136 5580 11192 5636
rect 11278 5580 11334 5636
rect 11136 5438 11192 5494
rect 11278 5438 11334 5494
rect 11136 5296 11192 5352
rect 11278 5296 11334 5352
rect 11136 5154 11192 5210
rect 11278 5154 11334 5210
rect 11136 5012 11192 5068
rect 11278 5012 11334 5068
rect 11136 4870 11192 4926
rect 11278 4870 11334 4926
rect 11136 4728 11192 4784
rect 11278 4728 11334 4784
rect 11136 4586 11192 4642
rect 11278 4586 11334 4642
rect 11136 4444 11192 4500
rect 11278 4444 11334 4500
rect 11136 4302 11192 4358
rect 11278 4302 11334 4358
rect 11136 4160 11192 4216
rect 11278 4160 11334 4216
rect 11136 4018 11192 4074
rect 11278 4018 11334 4074
rect 11136 3876 11192 3932
rect 11278 3876 11334 3932
rect 11136 3734 11192 3790
rect 11278 3734 11334 3790
rect 11136 3592 11192 3648
rect 11278 3592 11334 3648
rect 11136 3450 11192 3506
rect 11278 3450 11334 3506
rect 11136 3308 11192 3364
rect 11278 3308 11334 3364
rect 11136 3166 11192 3222
rect 11278 3166 11334 3222
rect 11136 3024 11192 3080
rect 11278 3024 11334 3080
rect 11136 2882 11192 2938
rect 11278 2882 11334 2938
rect 11136 2740 11192 2796
rect 11278 2740 11334 2796
rect 11136 2598 11192 2654
rect 11278 2598 11334 2654
rect 11136 2456 11192 2512
rect 11278 2456 11334 2512
rect 11136 2314 11192 2370
rect 11278 2314 11334 2370
rect 11136 2172 11192 2228
rect 11278 2172 11334 2228
rect 11136 2030 11192 2086
rect 11278 2030 11334 2086
rect 11136 1888 11192 1944
rect 11278 1888 11334 1944
rect 11136 1746 11192 1802
rect 11278 1746 11334 1802
rect 11136 1604 11192 1660
rect 11278 1604 11334 1660
rect 11136 1462 11192 1518
rect 11278 1462 11334 1518
rect 11136 1320 11192 1376
rect 11278 1320 11334 1376
rect 11136 1178 11192 1234
rect 11278 1178 11334 1234
rect 11136 1036 11192 1092
rect 11278 1036 11334 1092
rect 11136 894 11192 950
rect 11278 894 11334 950
rect 11136 752 11192 808
rect 11278 752 11334 808
rect 11136 610 11192 666
rect 11278 610 11334 666
rect 11136 468 11192 524
rect 11278 468 11334 524
rect 11536 12254 11592 12310
rect 11678 12254 11734 12310
rect 11536 12112 11592 12168
rect 11678 12112 11734 12168
rect 11536 11970 11592 12026
rect 11678 11970 11734 12026
rect 11536 11828 11592 11884
rect 11678 11828 11734 11884
rect 11536 11686 11592 11742
rect 11678 11686 11734 11742
rect 11536 11544 11592 11600
rect 11678 11544 11734 11600
rect 11536 11402 11592 11458
rect 11678 11402 11734 11458
rect 11536 11260 11592 11316
rect 11678 11260 11734 11316
rect 11536 11118 11592 11174
rect 11678 11118 11734 11174
rect 11536 10976 11592 11032
rect 11678 10976 11734 11032
rect 11536 10834 11592 10890
rect 11678 10834 11734 10890
rect 11536 10692 11592 10748
rect 11678 10692 11734 10748
rect 11536 10550 11592 10606
rect 11678 10550 11734 10606
rect 11536 10408 11592 10464
rect 11678 10408 11734 10464
rect 11536 10266 11592 10322
rect 11678 10266 11734 10322
rect 11536 10124 11592 10180
rect 11678 10124 11734 10180
rect 11536 9982 11592 10038
rect 11678 9982 11734 10038
rect 11536 9840 11592 9896
rect 11678 9840 11734 9896
rect 11536 9698 11592 9754
rect 11678 9698 11734 9754
rect 11536 9556 11592 9612
rect 11678 9556 11734 9612
rect 11536 9414 11592 9470
rect 11678 9414 11734 9470
rect 11536 9272 11592 9328
rect 11678 9272 11734 9328
rect 11536 9130 11592 9186
rect 11678 9130 11734 9186
rect 11536 8988 11592 9044
rect 11678 8988 11734 9044
rect 11536 8846 11592 8902
rect 11678 8846 11734 8902
rect 11536 8704 11592 8760
rect 11678 8704 11734 8760
rect 11536 8562 11592 8618
rect 11678 8562 11734 8618
rect 11536 8420 11592 8476
rect 11678 8420 11734 8476
rect 11536 8278 11592 8334
rect 11678 8278 11734 8334
rect 11536 8136 11592 8192
rect 11678 8136 11734 8192
rect 11536 7994 11592 8050
rect 11678 7994 11734 8050
rect 11536 7852 11592 7908
rect 11678 7852 11734 7908
rect 11536 7710 11592 7766
rect 11678 7710 11734 7766
rect 11536 7568 11592 7624
rect 11678 7568 11734 7624
rect 11536 7426 11592 7482
rect 11678 7426 11734 7482
rect 11536 7284 11592 7340
rect 11678 7284 11734 7340
rect 11536 7142 11592 7198
rect 11678 7142 11734 7198
rect 11536 7000 11592 7056
rect 11678 7000 11734 7056
rect 11536 6858 11592 6914
rect 11678 6858 11734 6914
rect 11536 6716 11592 6772
rect 11678 6716 11734 6772
rect 11536 6574 11592 6630
rect 11678 6574 11734 6630
rect 11536 6432 11592 6488
rect 11678 6432 11734 6488
rect 11536 6290 11592 6346
rect 11678 6290 11734 6346
rect 11536 6148 11592 6204
rect 11678 6148 11734 6204
rect 11536 6006 11592 6062
rect 11678 6006 11734 6062
rect 11536 5864 11592 5920
rect 11678 5864 11734 5920
rect 11536 5722 11592 5778
rect 11678 5722 11734 5778
rect 11536 5580 11592 5636
rect 11678 5580 11734 5636
rect 11536 5438 11592 5494
rect 11678 5438 11734 5494
rect 11536 5296 11592 5352
rect 11678 5296 11734 5352
rect 11536 5154 11592 5210
rect 11678 5154 11734 5210
rect 11536 5012 11592 5068
rect 11678 5012 11734 5068
rect 11536 4870 11592 4926
rect 11678 4870 11734 4926
rect 11536 4728 11592 4784
rect 11678 4728 11734 4784
rect 11536 4586 11592 4642
rect 11678 4586 11734 4642
rect 11536 4444 11592 4500
rect 11678 4444 11734 4500
rect 11536 4302 11592 4358
rect 11678 4302 11734 4358
rect 11536 4160 11592 4216
rect 11678 4160 11734 4216
rect 11536 4018 11592 4074
rect 11678 4018 11734 4074
rect 11536 3876 11592 3932
rect 11678 3876 11734 3932
rect 11536 3734 11592 3790
rect 11678 3734 11734 3790
rect 11536 3592 11592 3648
rect 11678 3592 11734 3648
rect 11536 3450 11592 3506
rect 11678 3450 11734 3506
rect 11536 3308 11592 3364
rect 11678 3308 11734 3364
rect 11536 3166 11592 3222
rect 11678 3166 11734 3222
rect 11536 3024 11592 3080
rect 11678 3024 11734 3080
rect 11536 2882 11592 2938
rect 11678 2882 11734 2938
rect 11536 2740 11592 2796
rect 11678 2740 11734 2796
rect 11536 2598 11592 2654
rect 11678 2598 11734 2654
rect 11536 2456 11592 2512
rect 11678 2456 11734 2512
rect 11536 2314 11592 2370
rect 11678 2314 11734 2370
rect 11536 2172 11592 2228
rect 11678 2172 11734 2228
rect 11536 2030 11592 2086
rect 11678 2030 11734 2086
rect 11536 1888 11592 1944
rect 11678 1888 11734 1944
rect 11536 1746 11592 1802
rect 11678 1746 11734 1802
rect 11536 1604 11592 1660
rect 11678 1604 11734 1660
rect 11536 1462 11592 1518
rect 11678 1462 11734 1518
rect 11536 1320 11592 1376
rect 11678 1320 11734 1376
rect 11536 1178 11592 1234
rect 11678 1178 11734 1234
rect 11536 1036 11592 1092
rect 11678 1036 11734 1092
rect 11536 894 11592 950
rect 11678 894 11734 950
rect 11536 752 11592 808
rect 11678 752 11734 808
rect 11536 610 11592 666
rect 11678 610 11734 666
rect 11536 468 11592 524
rect 11678 468 11734 524
rect 11941 12254 11997 12310
rect 12083 12254 12139 12310
rect 11941 12112 11997 12168
rect 12083 12112 12139 12168
rect 11941 11970 11997 12026
rect 12083 11970 12139 12026
rect 11941 11828 11997 11884
rect 12083 11828 12139 11884
rect 11941 11686 11997 11742
rect 12083 11686 12139 11742
rect 11941 11544 11997 11600
rect 12083 11544 12139 11600
rect 11941 11402 11997 11458
rect 12083 11402 12139 11458
rect 11941 11260 11997 11316
rect 12083 11260 12139 11316
rect 11941 11118 11997 11174
rect 12083 11118 12139 11174
rect 11941 10976 11997 11032
rect 12083 10976 12139 11032
rect 11941 10834 11997 10890
rect 12083 10834 12139 10890
rect 11941 10692 11997 10748
rect 12083 10692 12139 10748
rect 11941 10550 11997 10606
rect 12083 10550 12139 10606
rect 11941 10408 11997 10464
rect 12083 10408 12139 10464
rect 11941 10266 11997 10322
rect 12083 10266 12139 10322
rect 11941 10124 11997 10180
rect 12083 10124 12139 10180
rect 11941 9982 11997 10038
rect 12083 9982 12139 10038
rect 11941 9840 11997 9896
rect 12083 9840 12139 9896
rect 11941 9698 11997 9754
rect 12083 9698 12139 9754
rect 11941 9556 11997 9612
rect 12083 9556 12139 9612
rect 11941 9414 11997 9470
rect 12083 9414 12139 9470
rect 11941 9272 11997 9328
rect 12083 9272 12139 9328
rect 11941 9130 11997 9186
rect 12083 9130 12139 9186
rect 11941 8988 11997 9044
rect 12083 8988 12139 9044
rect 11941 8846 11997 8902
rect 12083 8846 12139 8902
rect 11941 8704 11997 8760
rect 12083 8704 12139 8760
rect 11941 8562 11997 8618
rect 12083 8562 12139 8618
rect 11941 8420 11997 8476
rect 12083 8420 12139 8476
rect 11941 8278 11997 8334
rect 12083 8278 12139 8334
rect 11941 8136 11997 8192
rect 12083 8136 12139 8192
rect 11941 7994 11997 8050
rect 12083 7994 12139 8050
rect 11941 7852 11997 7908
rect 12083 7852 12139 7908
rect 11941 7710 11997 7766
rect 12083 7710 12139 7766
rect 11941 7568 11997 7624
rect 12083 7568 12139 7624
rect 11941 7426 11997 7482
rect 12083 7426 12139 7482
rect 11941 7284 11997 7340
rect 12083 7284 12139 7340
rect 11941 7142 11997 7198
rect 12083 7142 12139 7198
rect 11941 7000 11997 7056
rect 12083 7000 12139 7056
rect 11941 6858 11997 6914
rect 12083 6858 12139 6914
rect 11941 6716 11997 6772
rect 12083 6716 12139 6772
rect 11941 6574 11997 6630
rect 12083 6574 12139 6630
rect 11941 6432 11997 6488
rect 12083 6432 12139 6488
rect 11941 6290 11997 6346
rect 12083 6290 12139 6346
rect 11941 6148 11997 6204
rect 12083 6148 12139 6204
rect 11941 6006 11997 6062
rect 12083 6006 12139 6062
rect 11941 5864 11997 5920
rect 12083 5864 12139 5920
rect 11941 5722 11997 5778
rect 12083 5722 12139 5778
rect 11941 5580 11997 5636
rect 12083 5580 12139 5636
rect 11941 5438 11997 5494
rect 12083 5438 12139 5494
rect 11941 5296 11997 5352
rect 12083 5296 12139 5352
rect 11941 5154 11997 5210
rect 12083 5154 12139 5210
rect 11941 5012 11997 5068
rect 12083 5012 12139 5068
rect 11941 4870 11997 4926
rect 12083 4870 12139 4926
rect 11941 4728 11997 4784
rect 12083 4728 12139 4784
rect 11941 4586 11997 4642
rect 12083 4586 12139 4642
rect 11941 4444 11997 4500
rect 12083 4444 12139 4500
rect 11941 4302 11997 4358
rect 12083 4302 12139 4358
rect 11941 4160 11997 4216
rect 12083 4160 12139 4216
rect 11941 4018 11997 4074
rect 12083 4018 12139 4074
rect 11941 3876 11997 3932
rect 12083 3876 12139 3932
rect 11941 3734 11997 3790
rect 12083 3734 12139 3790
rect 11941 3592 11997 3648
rect 12083 3592 12139 3648
rect 11941 3450 11997 3506
rect 12083 3450 12139 3506
rect 11941 3308 11997 3364
rect 12083 3308 12139 3364
rect 11941 3166 11997 3222
rect 12083 3166 12139 3222
rect 11941 3024 11997 3080
rect 12083 3024 12139 3080
rect 11941 2882 11997 2938
rect 12083 2882 12139 2938
rect 11941 2740 11997 2796
rect 12083 2740 12139 2796
rect 11941 2598 11997 2654
rect 12083 2598 12139 2654
rect 11941 2456 11997 2512
rect 12083 2456 12139 2512
rect 11941 2314 11997 2370
rect 12083 2314 12139 2370
rect 11941 2172 11997 2228
rect 12083 2172 12139 2228
rect 11941 2030 11997 2086
rect 12083 2030 12139 2086
rect 11941 1888 11997 1944
rect 12083 1888 12139 1944
rect 11941 1746 11997 1802
rect 12083 1746 12139 1802
rect 11941 1604 11997 1660
rect 12083 1604 12139 1660
rect 11941 1462 11997 1518
rect 12083 1462 12139 1518
rect 11941 1320 11997 1376
rect 12083 1320 12139 1376
rect 11941 1178 11997 1234
rect 12083 1178 12139 1234
rect 11941 1036 11997 1092
rect 12083 1036 12139 1092
rect 11941 894 11997 950
rect 12083 894 12139 950
rect 11941 752 11997 808
rect 12083 752 12139 808
rect 11941 610 11997 666
rect 12083 610 12139 666
rect 11941 468 11997 524
rect 12083 468 12139 524
rect 12526 12302 12582 12358
rect 12650 12302 12706 12358
rect 12774 12302 12830 12358
rect 12898 12302 12954 12358
rect 13022 12302 13078 12358
rect 12526 12178 12582 12234
rect 12650 12178 12706 12234
rect 12774 12178 12830 12234
rect 12898 12178 12954 12234
rect 13022 12178 13078 12234
rect 12526 12054 12582 12110
rect 12650 12054 12706 12110
rect 12774 12054 12830 12110
rect 12898 12054 12954 12110
rect 13022 12054 13078 12110
rect 12526 11930 12582 11986
rect 12650 11930 12706 11986
rect 12774 11930 12830 11986
rect 12898 11930 12954 11986
rect 13022 11930 13078 11986
rect 12526 11806 12582 11862
rect 12650 11806 12706 11862
rect 12774 11806 12830 11862
rect 12898 11806 12954 11862
rect 13022 11806 13078 11862
rect 12526 11682 12582 11738
rect 12650 11682 12706 11738
rect 12774 11682 12830 11738
rect 12898 11682 12954 11738
rect 13022 11682 13078 11738
rect 12526 11558 12582 11614
rect 12650 11558 12706 11614
rect 12774 11558 12830 11614
rect 12898 11558 12954 11614
rect 13022 11558 13078 11614
rect 12526 11434 12582 11490
rect 12650 11434 12706 11490
rect 12774 11434 12830 11490
rect 12898 11434 12954 11490
rect 13022 11434 13078 11490
rect 12526 11310 12582 11366
rect 12650 11310 12706 11366
rect 12774 11310 12830 11366
rect 12898 11310 12954 11366
rect 13022 11310 13078 11366
rect 12526 11186 12582 11242
rect 12650 11186 12706 11242
rect 12774 11186 12830 11242
rect 12898 11186 12954 11242
rect 13022 11186 13078 11242
rect 12526 11062 12582 11118
rect 12650 11062 12706 11118
rect 12774 11062 12830 11118
rect 12898 11062 12954 11118
rect 13022 11062 13078 11118
rect 12526 10938 12582 10994
rect 12650 10938 12706 10994
rect 12774 10938 12830 10994
rect 12898 10938 12954 10994
rect 13022 10938 13078 10994
rect 12526 10814 12582 10870
rect 12650 10814 12706 10870
rect 12774 10814 12830 10870
rect 12898 10814 12954 10870
rect 13022 10814 13078 10870
rect 12526 10690 12582 10746
rect 12650 10690 12706 10746
rect 12774 10690 12830 10746
rect 12898 10690 12954 10746
rect 13022 10690 13078 10746
rect 12526 10566 12582 10622
rect 12650 10566 12706 10622
rect 12774 10566 12830 10622
rect 12898 10566 12954 10622
rect 13022 10566 13078 10622
rect 12526 10442 12582 10498
rect 12650 10442 12706 10498
rect 12774 10442 12830 10498
rect 12898 10442 12954 10498
rect 13022 10442 13078 10498
rect 12526 10318 12582 10374
rect 12650 10318 12706 10374
rect 12774 10318 12830 10374
rect 12898 10318 12954 10374
rect 13022 10318 13078 10374
rect 12526 10194 12582 10250
rect 12650 10194 12706 10250
rect 12774 10194 12830 10250
rect 12898 10194 12954 10250
rect 13022 10194 13078 10250
rect 12526 10070 12582 10126
rect 12650 10070 12706 10126
rect 12774 10070 12830 10126
rect 12898 10070 12954 10126
rect 13022 10070 13078 10126
rect 12526 9946 12582 10002
rect 12650 9946 12706 10002
rect 12774 9946 12830 10002
rect 12898 9946 12954 10002
rect 13022 9946 13078 10002
rect 12526 9822 12582 9878
rect 12650 9822 12706 9878
rect 12774 9822 12830 9878
rect 12898 9822 12954 9878
rect 13022 9822 13078 9878
rect 12526 9698 12582 9754
rect 12650 9698 12706 9754
rect 12774 9698 12830 9754
rect 12898 9698 12954 9754
rect 13022 9698 13078 9754
rect 12526 9574 12582 9630
rect 12650 9574 12706 9630
rect 12774 9574 12830 9630
rect 12898 9574 12954 9630
rect 13022 9574 13078 9630
rect 12526 9450 12582 9506
rect 12650 9450 12706 9506
rect 12774 9450 12830 9506
rect 12898 9450 12954 9506
rect 13022 9450 13078 9506
rect 12526 9326 12582 9382
rect 12650 9326 12706 9382
rect 12774 9326 12830 9382
rect 12898 9326 12954 9382
rect 13022 9326 13078 9382
rect 12526 9202 12582 9258
rect 12650 9202 12706 9258
rect 12774 9202 12830 9258
rect 12898 9202 12954 9258
rect 13022 9202 13078 9258
rect 12526 9078 12582 9134
rect 12650 9078 12706 9134
rect 12774 9078 12830 9134
rect 12898 9078 12954 9134
rect 13022 9078 13078 9134
rect 12526 8954 12582 9010
rect 12650 8954 12706 9010
rect 12774 8954 12830 9010
rect 12898 8954 12954 9010
rect 13022 8954 13078 9010
rect 12526 8830 12582 8886
rect 12650 8830 12706 8886
rect 12774 8830 12830 8886
rect 12898 8830 12954 8886
rect 13022 8830 13078 8886
rect 12526 8706 12582 8762
rect 12650 8706 12706 8762
rect 12774 8706 12830 8762
rect 12898 8706 12954 8762
rect 13022 8706 13078 8762
rect 12526 8582 12582 8638
rect 12650 8582 12706 8638
rect 12774 8582 12830 8638
rect 12898 8582 12954 8638
rect 13022 8582 13078 8638
rect 12526 8458 12582 8514
rect 12650 8458 12706 8514
rect 12774 8458 12830 8514
rect 12898 8458 12954 8514
rect 13022 8458 13078 8514
rect 12526 8334 12582 8390
rect 12650 8334 12706 8390
rect 12774 8334 12830 8390
rect 12898 8334 12954 8390
rect 13022 8334 13078 8390
rect 12526 8210 12582 8266
rect 12650 8210 12706 8266
rect 12774 8210 12830 8266
rect 12898 8210 12954 8266
rect 13022 8210 13078 8266
rect 12526 8086 12582 8142
rect 12650 8086 12706 8142
rect 12774 8086 12830 8142
rect 12898 8086 12954 8142
rect 13022 8086 13078 8142
rect 12526 7962 12582 8018
rect 12650 7962 12706 8018
rect 12774 7962 12830 8018
rect 12898 7962 12954 8018
rect 13022 7962 13078 8018
rect 12526 7838 12582 7894
rect 12650 7838 12706 7894
rect 12774 7838 12830 7894
rect 12898 7838 12954 7894
rect 13022 7838 13078 7894
rect 12526 7714 12582 7770
rect 12650 7714 12706 7770
rect 12774 7714 12830 7770
rect 12898 7714 12954 7770
rect 13022 7714 13078 7770
rect 12526 7590 12582 7646
rect 12650 7590 12706 7646
rect 12774 7590 12830 7646
rect 12898 7590 12954 7646
rect 13022 7590 13078 7646
rect 12526 7466 12582 7522
rect 12650 7466 12706 7522
rect 12774 7466 12830 7522
rect 12898 7466 12954 7522
rect 13022 7466 13078 7522
rect 12526 7342 12582 7398
rect 12650 7342 12706 7398
rect 12774 7342 12830 7398
rect 12898 7342 12954 7398
rect 13022 7342 13078 7398
rect 12526 7218 12582 7274
rect 12650 7218 12706 7274
rect 12774 7218 12830 7274
rect 12898 7218 12954 7274
rect 13022 7218 13078 7274
rect 12526 7094 12582 7150
rect 12650 7094 12706 7150
rect 12774 7094 12830 7150
rect 12898 7094 12954 7150
rect 13022 7094 13078 7150
rect 12526 6970 12582 7026
rect 12650 6970 12706 7026
rect 12774 6970 12830 7026
rect 12898 6970 12954 7026
rect 13022 6970 13078 7026
rect 12526 6846 12582 6902
rect 12650 6846 12706 6902
rect 12774 6846 12830 6902
rect 12898 6846 12954 6902
rect 13022 6846 13078 6902
rect 12526 6722 12582 6778
rect 12650 6722 12706 6778
rect 12774 6722 12830 6778
rect 12898 6722 12954 6778
rect 13022 6722 13078 6778
rect 12526 6598 12582 6654
rect 12650 6598 12706 6654
rect 12774 6598 12830 6654
rect 12898 6598 12954 6654
rect 13022 6598 13078 6654
rect 12526 6474 12582 6530
rect 12650 6474 12706 6530
rect 12774 6474 12830 6530
rect 12898 6474 12954 6530
rect 13022 6474 13078 6530
rect 12526 6350 12582 6406
rect 12650 6350 12706 6406
rect 12774 6350 12830 6406
rect 12898 6350 12954 6406
rect 13022 6350 13078 6406
rect 12526 6226 12582 6282
rect 12650 6226 12706 6282
rect 12774 6226 12830 6282
rect 12898 6226 12954 6282
rect 13022 6226 13078 6282
rect 12526 6102 12582 6158
rect 12650 6102 12706 6158
rect 12774 6102 12830 6158
rect 12898 6102 12954 6158
rect 13022 6102 13078 6158
rect 12526 5978 12582 6034
rect 12650 5978 12706 6034
rect 12774 5978 12830 6034
rect 12898 5978 12954 6034
rect 13022 5978 13078 6034
rect 12526 5854 12582 5910
rect 12650 5854 12706 5910
rect 12774 5854 12830 5910
rect 12898 5854 12954 5910
rect 13022 5854 13078 5910
rect 12526 5730 12582 5786
rect 12650 5730 12706 5786
rect 12774 5730 12830 5786
rect 12898 5730 12954 5786
rect 13022 5730 13078 5786
rect 12526 5606 12582 5662
rect 12650 5606 12706 5662
rect 12774 5606 12830 5662
rect 12898 5606 12954 5662
rect 13022 5606 13078 5662
rect 12526 5482 12582 5538
rect 12650 5482 12706 5538
rect 12774 5482 12830 5538
rect 12898 5482 12954 5538
rect 13022 5482 13078 5538
rect 12526 5358 12582 5414
rect 12650 5358 12706 5414
rect 12774 5358 12830 5414
rect 12898 5358 12954 5414
rect 13022 5358 13078 5414
rect 12526 5234 12582 5290
rect 12650 5234 12706 5290
rect 12774 5234 12830 5290
rect 12898 5234 12954 5290
rect 13022 5234 13078 5290
rect 12526 5110 12582 5166
rect 12650 5110 12706 5166
rect 12774 5110 12830 5166
rect 12898 5110 12954 5166
rect 13022 5110 13078 5166
rect 12526 4986 12582 5042
rect 12650 4986 12706 5042
rect 12774 4986 12830 5042
rect 12898 4986 12954 5042
rect 13022 4986 13078 5042
rect 12526 4862 12582 4918
rect 12650 4862 12706 4918
rect 12774 4862 12830 4918
rect 12898 4862 12954 4918
rect 13022 4862 13078 4918
rect 12526 4738 12582 4794
rect 12650 4738 12706 4794
rect 12774 4738 12830 4794
rect 12898 4738 12954 4794
rect 13022 4738 13078 4794
rect 12526 4614 12582 4670
rect 12650 4614 12706 4670
rect 12774 4614 12830 4670
rect 12898 4614 12954 4670
rect 13022 4614 13078 4670
rect 12526 4490 12582 4546
rect 12650 4490 12706 4546
rect 12774 4490 12830 4546
rect 12898 4490 12954 4546
rect 13022 4490 13078 4546
rect 12526 4366 12582 4422
rect 12650 4366 12706 4422
rect 12774 4366 12830 4422
rect 12898 4366 12954 4422
rect 13022 4366 13078 4422
rect 12526 4242 12582 4298
rect 12650 4242 12706 4298
rect 12774 4242 12830 4298
rect 12898 4242 12954 4298
rect 13022 4242 13078 4298
rect 12526 4118 12582 4174
rect 12650 4118 12706 4174
rect 12774 4118 12830 4174
rect 12898 4118 12954 4174
rect 13022 4118 13078 4174
rect 12526 3994 12582 4050
rect 12650 3994 12706 4050
rect 12774 3994 12830 4050
rect 12898 3994 12954 4050
rect 13022 3994 13078 4050
rect 12526 3870 12582 3926
rect 12650 3870 12706 3926
rect 12774 3870 12830 3926
rect 12898 3870 12954 3926
rect 13022 3870 13078 3926
rect 12526 3746 12582 3802
rect 12650 3746 12706 3802
rect 12774 3746 12830 3802
rect 12898 3746 12954 3802
rect 13022 3746 13078 3802
rect 12526 3622 12582 3678
rect 12650 3622 12706 3678
rect 12774 3622 12830 3678
rect 12898 3622 12954 3678
rect 13022 3622 13078 3678
rect 12526 3498 12582 3554
rect 12650 3498 12706 3554
rect 12774 3498 12830 3554
rect 12898 3498 12954 3554
rect 13022 3498 13078 3554
rect 12526 3374 12582 3430
rect 12650 3374 12706 3430
rect 12774 3374 12830 3430
rect 12898 3374 12954 3430
rect 13022 3374 13078 3430
rect 12526 3250 12582 3306
rect 12650 3250 12706 3306
rect 12774 3250 12830 3306
rect 12898 3250 12954 3306
rect 13022 3250 13078 3306
rect 12526 3126 12582 3182
rect 12650 3126 12706 3182
rect 12774 3126 12830 3182
rect 12898 3126 12954 3182
rect 13022 3126 13078 3182
rect 12526 3002 12582 3058
rect 12650 3002 12706 3058
rect 12774 3002 12830 3058
rect 12898 3002 12954 3058
rect 13022 3002 13078 3058
rect 12526 2878 12582 2934
rect 12650 2878 12706 2934
rect 12774 2878 12830 2934
rect 12898 2878 12954 2934
rect 13022 2878 13078 2934
rect 12526 2754 12582 2810
rect 12650 2754 12706 2810
rect 12774 2754 12830 2810
rect 12898 2754 12954 2810
rect 13022 2754 13078 2810
rect 12526 2630 12582 2686
rect 12650 2630 12706 2686
rect 12774 2630 12830 2686
rect 12898 2630 12954 2686
rect 13022 2630 13078 2686
rect 12526 2506 12582 2562
rect 12650 2506 12706 2562
rect 12774 2506 12830 2562
rect 12898 2506 12954 2562
rect 13022 2506 13078 2562
rect 12526 2382 12582 2438
rect 12650 2382 12706 2438
rect 12774 2382 12830 2438
rect 12898 2382 12954 2438
rect 13022 2382 13078 2438
rect 12526 2258 12582 2314
rect 12650 2258 12706 2314
rect 12774 2258 12830 2314
rect 12898 2258 12954 2314
rect 13022 2258 13078 2314
rect 12526 2134 12582 2190
rect 12650 2134 12706 2190
rect 12774 2134 12830 2190
rect 12898 2134 12954 2190
rect 13022 2134 13078 2190
rect 12526 2010 12582 2066
rect 12650 2010 12706 2066
rect 12774 2010 12830 2066
rect 12898 2010 12954 2066
rect 13022 2010 13078 2066
rect 12526 1886 12582 1942
rect 12650 1886 12706 1942
rect 12774 1886 12830 1942
rect 12898 1886 12954 1942
rect 13022 1886 13078 1942
rect 12526 1762 12582 1818
rect 12650 1762 12706 1818
rect 12774 1762 12830 1818
rect 12898 1762 12954 1818
rect 13022 1762 13078 1818
rect 12526 1638 12582 1694
rect 12650 1638 12706 1694
rect 12774 1638 12830 1694
rect 12898 1638 12954 1694
rect 13022 1638 13078 1694
rect 12526 1514 12582 1570
rect 12650 1514 12706 1570
rect 12774 1514 12830 1570
rect 12898 1514 12954 1570
rect 13022 1514 13078 1570
rect 12526 1390 12582 1446
rect 12650 1390 12706 1446
rect 12774 1390 12830 1446
rect 12898 1390 12954 1446
rect 13022 1390 13078 1446
rect 12526 1266 12582 1322
rect 12650 1266 12706 1322
rect 12774 1266 12830 1322
rect 12898 1266 12954 1322
rect 13022 1266 13078 1322
rect 12526 1142 12582 1198
rect 12650 1142 12706 1198
rect 12774 1142 12830 1198
rect 12898 1142 12954 1198
rect 13022 1142 13078 1198
rect 12526 1018 12582 1074
rect 12650 1018 12706 1074
rect 12774 1018 12830 1074
rect 12898 1018 12954 1074
rect 13022 1018 13078 1074
rect 12526 894 12582 950
rect 12650 894 12706 950
rect 12774 894 12830 950
rect 12898 894 12954 950
rect 13022 894 13078 950
rect 12526 770 12582 826
rect 12650 770 12706 826
rect 12774 770 12830 826
rect 12898 770 12954 826
rect 13022 770 13078 826
rect 12526 646 12582 702
rect 12650 646 12706 702
rect 12774 646 12830 702
rect 12898 646 12954 702
rect 13022 646 13078 702
rect 12526 522 12582 578
rect 12650 522 12706 578
rect 12774 522 12830 578
rect 12898 522 12954 578
rect 13022 522 13078 578
rect 12526 398 12582 454
rect 12650 398 12706 454
rect 12774 398 12830 454
rect 12898 398 12954 454
rect 13022 398 13078 454
rect -286 274 -230 330
rect -162 274 -106 330
rect -38 274 18 330
rect 86 274 142 330
rect 210 274 266 330
rect 415 246 471 302
rect 557 246 613 302
rect 699 246 755 302
rect 841 246 897 302
rect 983 246 1039 302
rect 1125 246 1181 302
rect 1267 246 1323 302
rect 1409 246 1465 302
rect 1551 246 1607 302
rect 1693 246 1749 302
rect 1835 246 1891 302
rect 1977 246 2033 302
rect 2119 246 2175 302
rect 2261 246 2317 302
rect 2403 246 2459 302
rect 2545 246 2601 302
rect 2687 246 2743 302
rect 2829 246 2885 302
rect 2971 246 3027 302
rect 3113 246 3169 302
rect 3255 246 3311 302
rect 3397 246 3453 302
rect 3539 246 3595 302
rect 3681 246 3737 302
rect 3823 246 3879 302
rect 3965 246 4021 302
rect 4107 246 4163 302
rect 4249 246 4305 302
rect 4391 246 4447 302
rect 4533 246 4589 302
rect 4675 246 4731 302
rect 4817 246 4873 302
rect 4959 246 5015 302
rect 5101 246 5157 302
rect 5243 246 5299 302
rect 5385 246 5441 302
rect 5527 246 5583 302
rect 5669 246 5725 302
rect 5811 246 5867 302
rect 5953 246 6009 302
rect 6095 246 6151 302
rect 6237 246 6293 302
rect 6379 246 6435 302
rect 6521 246 6577 302
rect 6663 246 6719 302
rect 6805 246 6861 302
rect 6947 246 7003 302
rect 7089 246 7145 302
rect 7231 246 7287 302
rect 7373 246 7429 302
rect 7515 246 7571 302
rect 7657 246 7713 302
rect 7799 246 7855 302
rect 7941 246 7997 302
rect 8083 246 8139 302
rect 8225 246 8281 302
rect 8367 246 8423 302
rect 8509 246 8565 302
rect 8651 246 8707 302
rect 8793 246 8849 302
rect 8935 246 8991 302
rect 9077 246 9133 302
rect 9219 246 9275 302
rect 9361 246 9417 302
rect 9503 246 9559 302
rect 9645 246 9701 302
rect 9787 246 9843 302
rect 9929 246 9985 302
rect 10071 246 10127 302
rect 10213 246 10269 302
rect 10355 246 10411 302
rect 10497 246 10553 302
rect 10639 246 10695 302
rect 10781 246 10837 302
rect 10923 246 10979 302
rect 11065 246 11121 302
rect 11207 246 11263 302
rect 11349 246 11405 302
rect 11491 246 11547 302
rect 11633 246 11689 302
rect 11775 246 11831 302
rect 11917 246 11973 302
rect 12059 246 12115 302
rect 12201 246 12257 302
rect 12343 246 12399 302
rect 12526 274 12582 330
rect 12650 274 12706 330
rect 12774 274 12830 330
rect 12898 274 12954 330
rect 13022 274 13078 330
rect -286 150 -230 206
rect -162 150 -106 206
rect -38 150 18 206
rect 86 150 142 206
rect 210 150 266 206
rect 415 104 471 160
rect 557 104 613 160
rect 699 104 755 160
rect 841 104 897 160
rect 983 104 1039 160
rect 1125 104 1181 160
rect 1267 104 1323 160
rect 1409 104 1465 160
rect 1551 104 1607 160
rect 1693 104 1749 160
rect 1835 104 1891 160
rect 1977 104 2033 160
rect 2119 104 2175 160
rect 2261 104 2317 160
rect 2403 104 2459 160
rect 2545 104 2601 160
rect 2687 104 2743 160
rect 2829 104 2885 160
rect 2971 104 3027 160
rect 3113 104 3169 160
rect 3255 104 3311 160
rect 3397 104 3453 160
rect 3539 104 3595 160
rect 3681 104 3737 160
rect 3823 104 3879 160
rect 3965 104 4021 160
rect 4107 104 4163 160
rect 4249 104 4305 160
rect 4391 104 4447 160
rect 4533 104 4589 160
rect 4675 104 4731 160
rect 4817 104 4873 160
rect 4959 104 5015 160
rect 5101 104 5157 160
rect 5243 104 5299 160
rect 5385 104 5441 160
rect 5527 104 5583 160
rect 5669 104 5725 160
rect 5811 104 5867 160
rect 5953 104 6009 160
rect 6095 104 6151 160
rect 6237 104 6293 160
rect 6379 104 6435 160
rect 6521 104 6577 160
rect 6663 104 6719 160
rect 6805 104 6861 160
rect 6947 104 7003 160
rect 7089 104 7145 160
rect 7231 104 7287 160
rect 7373 104 7429 160
rect 7515 104 7571 160
rect 7657 104 7713 160
rect 7799 104 7855 160
rect 7941 104 7997 160
rect 8083 104 8139 160
rect 8225 104 8281 160
rect 8367 104 8423 160
rect 8509 104 8565 160
rect 8651 104 8707 160
rect 8793 104 8849 160
rect 8935 104 8991 160
rect 9077 104 9133 160
rect 9219 104 9275 160
rect 9361 104 9417 160
rect 9503 104 9559 160
rect 9645 104 9701 160
rect 9787 104 9843 160
rect 9929 104 9985 160
rect 10071 104 10127 160
rect 10213 104 10269 160
rect 10355 104 10411 160
rect 10497 104 10553 160
rect 10639 104 10695 160
rect 10781 104 10837 160
rect 10923 104 10979 160
rect 11065 104 11121 160
rect 11207 104 11263 160
rect 11349 104 11405 160
rect 11491 104 11547 160
rect 11633 104 11689 160
rect 11775 104 11831 160
rect 11917 104 11973 160
rect 12059 104 12115 160
rect 12201 104 12257 160
rect 12343 104 12399 160
rect 12526 150 12582 206
rect 12650 150 12706 206
rect 12774 150 12830 206
rect 12898 150 12954 206
rect 13022 150 13078 206
<< metal3 >>
rect -400 12949 13200 13065
rect -400 12893 -254 12949
rect -198 12893 -130 12949
rect -74 12893 -6 12949
rect 50 12893 118 12949
rect 174 12893 242 12949
rect 298 12893 366 12949
rect 422 12893 490 12949
rect 546 12893 614 12949
rect 670 12893 738 12949
rect 794 12893 862 12949
rect 918 12893 986 12949
rect 1042 12893 1110 12949
rect 1166 12893 1234 12949
rect 1290 12893 1358 12949
rect 1414 12893 1482 12949
rect 1538 12893 1606 12949
rect 1662 12893 1730 12949
rect 1786 12893 1854 12949
rect 1910 12893 1978 12949
rect 2034 12893 2102 12949
rect 2158 12893 2226 12949
rect 2282 12893 2350 12949
rect 2406 12893 2474 12949
rect 2530 12893 2598 12949
rect 2654 12893 2722 12949
rect 2778 12893 2846 12949
rect 2902 12893 2970 12949
rect 3026 12893 3094 12949
rect 3150 12893 3218 12949
rect 3274 12893 3342 12949
rect 3398 12893 3466 12949
rect 3522 12893 3590 12949
rect 3646 12893 3714 12949
rect 3770 12893 3838 12949
rect 3894 12893 3962 12949
rect 4018 12893 4086 12949
rect 4142 12893 4210 12949
rect 4266 12893 4334 12949
rect 4390 12893 4458 12949
rect 4514 12893 4582 12949
rect 4638 12893 4706 12949
rect 4762 12893 4830 12949
rect 4886 12893 4954 12949
rect 5010 12893 5078 12949
rect 5134 12893 5202 12949
rect 5258 12893 5326 12949
rect 5382 12893 5450 12949
rect 5506 12893 5574 12949
rect 5630 12893 5698 12949
rect 5754 12893 5822 12949
rect 5878 12893 5946 12949
rect 6002 12893 6070 12949
rect 6126 12893 6194 12949
rect 6250 12893 6318 12949
rect 6374 12893 6442 12949
rect 6498 12893 6566 12949
rect 6622 12893 6690 12949
rect 6746 12893 6814 12949
rect 6870 12893 6938 12949
rect 6994 12893 7062 12949
rect 7118 12893 7186 12949
rect 7242 12893 7310 12949
rect 7366 12893 7434 12949
rect 7490 12893 7558 12949
rect 7614 12893 7682 12949
rect 7738 12893 7806 12949
rect 7862 12893 7930 12949
rect 7986 12893 8054 12949
rect 8110 12893 8178 12949
rect 8234 12893 8302 12949
rect 8358 12893 8426 12949
rect 8482 12893 8550 12949
rect 8606 12893 8674 12949
rect 8730 12893 8798 12949
rect 8854 12893 8922 12949
rect 8978 12893 9046 12949
rect 9102 12893 9170 12949
rect 9226 12893 9294 12949
rect 9350 12893 9418 12949
rect 9474 12893 9542 12949
rect 9598 12893 9666 12949
rect 9722 12893 9790 12949
rect 9846 12893 9914 12949
rect 9970 12893 10038 12949
rect 10094 12893 10162 12949
rect 10218 12893 10286 12949
rect 10342 12893 10410 12949
rect 10466 12893 10534 12949
rect 10590 12893 10658 12949
rect 10714 12893 10782 12949
rect 10838 12893 10906 12949
rect 10962 12893 11030 12949
rect 11086 12893 11154 12949
rect 11210 12893 11278 12949
rect 11334 12893 11402 12949
rect 11458 12893 11526 12949
rect 11582 12893 11650 12949
rect 11706 12893 11774 12949
rect 11830 12893 11898 12949
rect 11954 12893 12022 12949
rect 12078 12893 12146 12949
rect 12202 12893 12270 12949
rect 12326 12893 12394 12949
rect 12450 12893 12518 12949
rect 12574 12893 12642 12949
rect 12698 12893 12766 12949
rect 12822 12893 12890 12949
rect 12946 12893 13014 12949
rect 13070 12893 13200 12949
rect -400 12825 13200 12893
rect -400 12769 -254 12825
rect -198 12769 -130 12825
rect -74 12769 -6 12825
rect 50 12769 118 12825
rect 174 12769 242 12825
rect 298 12769 366 12825
rect 422 12769 490 12825
rect 546 12769 614 12825
rect 670 12769 738 12825
rect 794 12769 862 12825
rect 918 12769 986 12825
rect 1042 12769 1110 12825
rect 1166 12769 1234 12825
rect 1290 12769 1358 12825
rect 1414 12769 1482 12825
rect 1538 12769 1606 12825
rect 1662 12769 1730 12825
rect 1786 12769 1854 12825
rect 1910 12769 1978 12825
rect 2034 12769 2102 12825
rect 2158 12769 2226 12825
rect 2282 12769 2350 12825
rect 2406 12769 2474 12825
rect 2530 12769 2598 12825
rect 2654 12769 2722 12825
rect 2778 12769 2846 12825
rect 2902 12769 2970 12825
rect 3026 12769 3094 12825
rect 3150 12769 3218 12825
rect 3274 12769 3342 12825
rect 3398 12769 3466 12825
rect 3522 12769 3590 12825
rect 3646 12769 3714 12825
rect 3770 12769 3838 12825
rect 3894 12769 3962 12825
rect 4018 12769 4086 12825
rect 4142 12769 4210 12825
rect 4266 12769 4334 12825
rect 4390 12769 4458 12825
rect 4514 12769 4582 12825
rect 4638 12769 4706 12825
rect 4762 12769 4830 12825
rect 4886 12769 4954 12825
rect 5010 12769 5078 12825
rect 5134 12769 5202 12825
rect 5258 12769 5326 12825
rect 5382 12769 5450 12825
rect 5506 12769 5574 12825
rect 5630 12769 5698 12825
rect 5754 12769 5822 12825
rect 5878 12769 5946 12825
rect 6002 12769 6070 12825
rect 6126 12769 6194 12825
rect 6250 12769 6318 12825
rect 6374 12769 6442 12825
rect 6498 12769 6566 12825
rect 6622 12769 6690 12825
rect 6746 12769 6814 12825
rect 6870 12769 6938 12825
rect 6994 12769 7062 12825
rect 7118 12769 7186 12825
rect 7242 12769 7310 12825
rect 7366 12769 7434 12825
rect 7490 12769 7558 12825
rect 7614 12769 7682 12825
rect 7738 12769 7806 12825
rect 7862 12769 7930 12825
rect 7986 12769 8054 12825
rect 8110 12769 8178 12825
rect 8234 12769 8302 12825
rect 8358 12769 8426 12825
rect 8482 12769 8550 12825
rect 8606 12769 8674 12825
rect 8730 12769 8798 12825
rect 8854 12769 8922 12825
rect 8978 12769 9046 12825
rect 9102 12769 9170 12825
rect 9226 12769 9294 12825
rect 9350 12769 9418 12825
rect 9474 12769 9542 12825
rect 9598 12769 9666 12825
rect 9722 12769 9790 12825
rect 9846 12769 9914 12825
rect 9970 12769 10038 12825
rect 10094 12769 10162 12825
rect 10218 12769 10286 12825
rect 10342 12769 10410 12825
rect 10466 12769 10534 12825
rect 10590 12769 10658 12825
rect 10714 12769 10782 12825
rect 10838 12769 10906 12825
rect 10962 12769 11030 12825
rect 11086 12769 11154 12825
rect 11210 12769 11278 12825
rect 11334 12769 11402 12825
rect 11458 12769 11526 12825
rect 11582 12769 11650 12825
rect 11706 12769 11774 12825
rect 11830 12769 11898 12825
rect 11954 12769 12022 12825
rect 12078 12769 12146 12825
rect 12202 12769 12270 12825
rect 12326 12769 12394 12825
rect 12450 12769 12518 12825
rect 12574 12769 12642 12825
rect 12698 12769 12766 12825
rect 12822 12769 12890 12825
rect 12946 12769 13014 12825
rect 13070 12769 13200 12825
rect -400 12701 13200 12769
rect -400 12645 -254 12701
rect -198 12645 -130 12701
rect -74 12645 -6 12701
rect 50 12645 118 12701
rect 174 12645 242 12701
rect 298 12645 366 12701
rect 422 12645 490 12701
rect 546 12645 614 12701
rect 670 12645 738 12701
rect 794 12645 862 12701
rect 918 12645 986 12701
rect 1042 12645 1110 12701
rect 1166 12645 1234 12701
rect 1290 12645 1358 12701
rect 1414 12645 1482 12701
rect 1538 12645 1606 12701
rect 1662 12645 1730 12701
rect 1786 12645 1854 12701
rect 1910 12645 1978 12701
rect 2034 12645 2102 12701
rect 2158 12645 2226 12701
rect 2282 12645 2350 12701
rect 2406 12645 2474 12701
rect 2530 12645 2598 12701
rect 2654 12645 2722 12701
rect 2778 12645 2846 12701
rect 2902 12645 2970 12701
rect 3026 12645 3094 12701
rect 3150 12645 3218 12701
rect 3274 12645 3342 12701
rect 3398 12645 3466 12701
rect 3522 12645 3590 12701
rect 3646 12645 3714 12701
rect 3770 12645 3838 12701
rect 3894 12645 3962 12701
rect 4018 12645 4086 12701
rect 4142 12645 4210 12701
rect 4266 12645 4334 12701
rect 4390 12645 4458 12701
rect 4514 12645 4582 12701
rect 4638 12645 4706 12701
rect 4762 12645 4830 12701
rect 4886 12645 4954 12701
rect 5010 12645 5078 12701
rect 5134 12645 5202 12701
rect 5258 12645 5326 12701
rect 5382 12645 5450 12701
rect 5506 12645 5574 12701
rect 5630 12645 5698 12701
rect 5754 12645 5822 12701
rect 5878 12645 5946 12701
rect 6002 12645 6070 12701
rect 6126 12645 6194 12701
rect 6250 12645 6318 12701
rect 6374 12645 6442 12701
rect 6498 12645 6566 12701
rect 6622 12645 6690 12701
rect 6746 12645 6814 12701
rect 6870 12645 6938 12701
rect 6994 12645 7062 12701
rect 7118 12645 7186 12701
rect 7242 12645 7310 12701
rect 7366 12645 7434 12701
rect 7490 12645 7558 12701
rect 7614 12645 7682 12701
rect 7738 12645 7806 12701
rect 7862 12645 7930 12701
rect 7986 12645 8054 12701
rect 8110 12645 8178 12701
rect 8234 12645 8302 12701
rect 8358 12645 8426 12701
rect 8482 12645 8550 12701
rect 8606 12645 8674 12701
rect 8730 12645 8798 12701
rect 8854 12645 8922 12701
rect 8978 12645 9046 12701
rect 9102 12645 9170 12701
rect 9226 12645 9294 12701
rect 9350 12645 9418 12701
rect 9474 12645 9542 12701
rect 9598 12645 9666 12701
rect 9722 12645 9790 12701
rect 9846 12645 9914 12701
rect 9970 12645 10038 12701
rect 10094 12645 10162 12701
rect 10218 12645 10286 12701
rect 10342 12645 10410 12701
rect 10466 12645 10534 12701
rect 10590 12645 10658 12701
rect 10714 12645 10782 12701
rect 10838 12645 10906 12701
rect 10962 12645 11030 12701
rect 11086 12645 11154 12701
rect 11210 12645 11278 12701
rect 11334 12645 11402 12701
rect 11458 12645 11526 12701
rect 11582 12645 11650 12701
rect 11706 12645 11774 12701
rect 11830 12645 11898 12701
rect 11954 12645 12022 12701
rect 12078 12645 12146 12701
rect 12202 12645 12270 12701
rect 12326 12645 12394 12701
rect 12450 12645 12518 12701
rect 12574 12645 12642 12701
rect 12698 12645 12766 12701
rect 12822 12645 12890 12701
rect 12946 12645 13014 12701
rect 13070 12645 13200 12701
rect -400 12577 13200 12645
rect -400 12521 -254 12577
rect -198 12521 -130 12577
rect -74 12521 -6 12577
rect 50 12521 118 12577
rect 174 12521 242 12577
rect 298 12521 366 12577
rect 422 12521 490 12577
rect 546 12521 614 12577
rect 670 12521 738 12577
rect 794 12521 862 12577
rect 918 12521 986 12577
rect 1042 12521 1110 12577
rect 1166 12521 1234 12577
rect 1290 12521 1358 12577
rect 1414 12521 1482 12577
rect 1538 12521 1606 12577
rect 1662 12521 1730 12577
rect 1786 12521 1854 12577
rect 1910 12521 1978 12577
rect 2034 12521 2102 12577
rect 2158 12521 2226 12577
rect 2282 12521 2350 12577
rect 2406 12521 2474 12577
rect 2530 12521 2598 12577
rect 2654 12521 2722 12577
rect 2778 12521 2846 12577
rect 2902 12521 2970 12577
rect 3026 12521 3094 12577
rect 3150 12521 3218 12577
rect 3274 12521 3342 12577
rect 3398 12521 3466 12577
rect 3522 12521 3590 12577
rect 3646 12521 3714 12577
rect 3770 12521 3838 12577
rect 3894 12521 3962 12577
rect 4018 12521 4086 12577
rect 4142 12521 4210 12577
rect 4266 12521 4334 12577
rect 4390 12521 4458 12577
rect 4514 12521 4582 12577
rect 4638 12521 4706 12577
rect 4762 12521 4830 12577
rect 4886 12521 4954 12577
rect 5010 12521 5078 12577
rect 5134 12521 5202 12577
rect 5258 12521 5326 12577
rect 5382 12521 5450 12577
rect 5506 12521 5574 12577
rect 5630 12521 5698 12577
rect 5754 12521 5822 12577
rect 5878 12521 5946 12577
rect 6002 12521 6070 12577
rect 6126 12521 6194 12577
rect 6250 12521 6318 12577
rect 6374 12521 6442 12577
rect 6498 12521 6566 12577
rect 6622 12521 6690 12577
rect 6746 12521 6814 12577
rect 6870 12521 6938 12577
rect 6994 12521 7062 12577
rect 7118 12521 7186 12577
rect 7242 12521 7310 12577
rect 7366 12521 7434 12577
rect 7490 12521 7558 12577
rect 7614 12521 7682 12577
rect 7738 12521 7806 12577
rect 7862 12521 7930 12577
rect 7986 12521 8054 12577
rect 8110 12521 8178 12577
rect 8234 12521 8302 12577
rect 8358 12521 8426 12577
rect 8482 12521 8550 12577
rect 8606 12521 8674 12577
rect 8730 12521 8798 12577
rect 8854 12521 8922 12577
rect 8978 12521 9046 12577
rect 9102 12521 9170 12577
rect 9226 12521 9294 12577
rect 9350 12521 9418 12577
rect 9474 12521 9542 12577
rect 9598 12521 9666 12577
rect 9722 12521 9790 12577
rect 9846 12521 9914 12577
rect 9970 12521 10038 12577
rect 10094 12521 10162 12577
rect 10218 12521 10286 12577
rect 10342 12521 10410 12577
rect 10466 12521 10534 12577
rect 10590 12521 10658 12577
rect 10714 12521 10782 12577
rect 10838 12521 10906 12577
rect 10962 12521 11030 12577
rect 11086 12521 11154 12577
rect 11210 12521 11278 12577
rect 11334 12521 11402 12577
rect 11458 12521 11526 12577
rect 11582 12521 11650 12577
rect 11706 12521 11774 12577
rect 11830 12521 11898 12577
rect 11954 12521 12022 12577
rect 12078 12521 12146 12577
rect 12202 12521 12270 12577
rect 12326 12521 12394 12577
rect 12450 12521 12518 12577
rect 12574 12521 12642 12577
rect 12698 12521 12766 12577
rect 12822 12521 12890 12577
rect 12946 12521 13014 12577
rect 13070 12521 13200 12577
rect -400 12400 13200 12521
rect -400 12358 400 12400
rect -400 12302 -286 12358
rect -230 12302 -162 12358
rect -106 12302 -38 12358
rect 18 12302 86 12358
rect 142 12302 210 12358
rect 266 12302 400 12358
rect -400 12234 400 12302
rect -400 12178 -286 12234
rect -230 12178 -162 12234
rect -106 12178 -38 12234
rect 18 12178 86 12234
rect 142 12178 210 12234
rect 266 12178 400 12234
rect -400 12110 400 12178
rect -400 12054 -286 12110
rect -230 12054 -162 12110
rect -106 12054 -38 12110
rect 18 12054 86 12110
rect 142 12054 210 12110
rect 266 12054 400 12110
rect -400 11986 400 12054
rect -400 11930 -286 11986
rect -230 11930 -162 11986
rect -106 11930 -38 11986
rect 18 11930 86 11986
rect 142 11930 210 11986
rect 266 11930 400 11986
rect -400 11862 400 11930
rect -400 11806 -286 11862
rect -230 11806 -162 11862
rect -106 11806 -38 11862
rect 18 11806 86 11862
rect 142 11806 210 11862
rect 266 11806 400 11862
rect -400 11738 400 11806
rect -400 11682 -286 11738
rect -230 11682 -162 11738
rect -106 11682 -38 11738
rect 18 11682 86 11738
rect 142 11682 210 11738
rect 266 11682 400 11738
rect -400 11614 400 11682
rect -400 11558 -286 11614
rect -230 11558 -162 11614
rect -106 11558 -38 11614
rect 18 11558 86 11614
rect 142 11558 210 11614
rect 266 11558 400 11614
rect -400 11490 400 11558
rect -400 11434 -286 11490
rect -230 11434 -162 11490
rect -106 11434 -38 11490
rect 18 11434 86 11490
rect 142 11434 210 11490
rect 266 11434 400 11490
rect -400 11366 400 11434
rect -400 11310 -286 11366
rect -230 11310 -162 11366
rect -106 11310 -38 11366
rect 18 11310 86 11366
rect 142 11310 210 11366
rect 266 11310 400 11366
rect -400 11242 400 11310
rect -400 11186 -286 11242
rect -230 11186 -162 11242
rect -106 11186 -38 11242
rect 18 11186 86 11242
rect 142 11186 210 11242
rect 266 11186 400 11242
rect -400 11118 400 11186
rect -400 11062 -286 11118
rect -230 11062 -162 11118
rect -106 11062 -38 11118
rect 18 11062 86 11118
rect 142 11062 210 11118
rect 266 11062 400 11118
rect -400 10994 400 11062
rect -400 10938 -286 10994
rect -230 10938 -162 10994
rect -106 10938 -38 10994
rect 18 10938 86 10994
rect 142 10938 210 10994
rect 266 10938 400 10994
rect -400 10870 400 10938
rect -400 10814 -286 10870
rect -230 10814 -162 10870
rect -106 10814 -38 10870
rect 18 10814 86 10870
rect 142 10814 210 10870
rect 266 10814 400 10870
rect -400 10746 400 10814
rect -400 10690 -286 10746
rect -230 10690 -162 10746
rect -106 10690 -38 10746
rect 18 10690 86 10746
rect 142 10690 210 10746
rect 266 10690 400 10746
rect -400 10622 400 10690
rect -400 10566 -286 10622
rect -230 10566 -162 10622
rect -106 10566 -38 10622
rect 18 10566 86 10622
rect 142 10566 210 10622
rect 266 10566 400 10622
rect -400 10498 400 10566
rect -400 10442 -286 10498
rect -230 10442 -162 10498
rect -106 10442 -38 10498
rect 18 10442 86 10498
rect 142 10442 210 10498
rect 266 10442 400 10498
rect -400 10374 400 10442
rect -400 10318 -286 10374
rect -230 10318 -162 10374
rect -106 10318 -38 10374
rect 18 10318 86 10374
rect 142 10318 210 10374
rect 266 10318 400 10374
rect -400 10250 400 10318
rect -400 10194 -286 10250
rect -230 10194 -162 10250
rect -106 10194 -38 10250
rect 18 10194 86 10250
rect 142 10194 210 10250
rect 266 10194 400 10250
rect -400 10126 400 10194
rect -400 10070 -286 10126
rect -230 10070 -162 10126
rect -106 10070 -38 10126
rect 18 10070 86 10126
rect 142 10070 210 10126
rect 266 10070 400 10126
rect -400 10002 400 10070
rect -400 9946 -286 10002
rect -230 9946 -162 10002
rect -106 9946 -38 10002
rect 18 9946 86 10002
rect 142 9946 210 10002
rect 266 9946 400 10002
rect -400 9878 400 9946
rect -400 9822 -286 9878
rect -230 9822 -162 9878
rect -106 9822 -38 9878
rect 18 9822 86 9878
rect 142 9822 210 9878
rect 266 9822 400 9878
rect -400 9754 400 9822
rect -400 9698 -286 9754
rect -230 9698 -162 9754
rect -106 9698 -38 9754
rect 18 9698 86 9754
rect 142 9698 210 9754
rect 266 9698 400 9754
rect -400 9630 400 9698
rect -400 9574 -286 9630
rect -230 9574 -162 9630
rect -106 9574 -38 9630
rect 18 9574 86 9630
rect 142 9574 210 9630
rect 266 9574 400 9630
rect -400 9506 400 9574
rect -400 9450 -286 9506
rect -230 9450 -162 9506
rect -106 9450 -38 9506
rect 18 9450 86 9506
rect 142 9450 210 9506
rect 266 9450 400 9506
rect -400 9382 400 9450
rect -400 9326 -286 9382
rect -230 9326 -162 9382
rect -106 9326 -38 9382
rect 18 9326 86 9382
rect 142 9326 210 9382
rect 266 9326 400 9382
rect -400 9258 400 9326
rect -400 9202 -286 9258
rect -230 9202 -162 9258
rect -106 9202 -38 9258
rect 18 9202 86 9258
rect 142 9202 210 9258
rect 266 9202 400 9258
rect -400 9134 400 9202
rect -400 9078 -286 9134
rect -230 9078 -162 9134
rect -106 9078 -38 9134
rect 18 9078 86 9134
rect 142 9078 210 9134
rect 266 9078 400 9134
rect -400 9010 400 9078
rect -400 8954 -286 9010
rect -230 8954 -162 9010
rect -106 8954 -38 9010
rect 18 8954 86 9010
rect 142 8954 210 9010
rect 266 8954 400 9010
rect -400 8886 400 8954
rect -400 8830 -286 8886
rect -230 8830 -162 8886
rect -106 8830 -38 8886
rect 18 8830 86 8886
rect 142 8830 210 8886
rect 266 8830 400 8886
rect -400 8762 400 8830
rect -400 8706 -286 8762
rect -230 8706 -162 8762
rect -106 8706 -38 8762
rect 18 8706 86 8762
rect 142 8706 210 8762
rect 266 8706 400 8762
rect -400 8638 400 8706
rect -400 8582 -286 8638
rect -230 8582 -162 8638
rect -106 8582 -38 8638
rect 18 8582 86 8638
rect 142 8582 210 8638
rect 266 8582 400 8638
rect -400 8514 400 8582
rect -400 8458 -286 8514
rect -230 8458 -162 8514
rect -106 8458 -38 8514
rect 18 8458 86 8514
rect 142 8458 210 8514
rect 266 8458 400 8514
rect -400 8390 400 8458
rect -400 8334 -286 8390
rect -230 8334 -162 8390
rect -106 8334 -38 8390
rect 18 8334 86 8390
rect 142 8334 210 8390
rect 266 8334 400 8390
rect -400 8266 400 8334
rect -400 8210 -286 8266
rect -230 8210 -162 8266
rect -106 8210 -38 8266
rect 18 8210 86 8266
rect 142 8210 210 8266
rect 266 8210 400 8266
rect -400 8142 400 8210
rect -400 8086 -286 8142
rect -230 8086 -162 8142
rect -106 8086 -38 8142
rect 18 8086 86 8142
rect 142 8086 210 8142
rect 266 8086 400 8142
rect -400 8018 400 8086
rect -400 7962 -286 8018
rect -230 7962 -162 8018
rect -106 7962 -38 8018
rect 18 7962 86 8018
rect 142 7962 210 8018
rect 266 7962 400 8018
rect -400 7894 400 7962
rect -400 7838 -286 7894
rect -230 7838 -162 7894
rect -106 7838 -38 7894
rect 18 7838 86 7894
rect 142 7838 210 7894
rect 266 7838 400 7894
rect -400 7770 400 7838
rect -400 7714 -286 7770
rect -230 7714 -162 7770
rect -106 7714 -38 7770
rect 18 7714 86 7770
rect 142 7714 210 7770
rect 266 7714 400 7770
rect -400 7646 400 7714
rect -400 7590 -286 7646
rect -230 7590 -162 7646
rect -106 7590 -38 7646
rect 18 7590 86 7646
rect 142 7590 210 7646
rect 266 7590 400 7646
rect -400 7522 400 7590
rect -400 7466 -286 7522
rect -230 7466 -162 7522
rect -106 7466 -38 7522
rect 18 7466 86 7522
rect 142 7466 210 7522
rect 266 7466 400 7522
rect -400 7398 400 7466
rect -400 7342 -286 7398
rect -230 7342 -162 7398
rect -106 7342 -38 7398
rect 18 7342 86 7398
rect 142 7342 210 7398
rect 266 7342 400 7398
rect -400 7274 400 7342
rect -400 7218 -286 7274
rect -230 7218 -162 7274
rect -106 7218 -38 7274
rect 18 7218 86 7274
rect 142 7218 210 7274
rect 266 7218 400 7274
rect -400 7150 400 7218
rect -400 7094 -286 7150
rect -230 7094 -162 7150
rect -106 7094 -38 7150
rect 18 7094 86 7150
rect 142 7094 210 7150
rect 266 7094 400 7150
rect -400 7026 400 7094
rect -400 6970 -286 7026
rect -230 6970 -162 7026
rect -106 6970 -38 7026
rect 18 6970 86 7026
rect 142 6970 210 7026
rect 266 6970 400 7026
rect -400 6902 400 6970
rect -400 6846 -286 6902
rect -230 6846 -162 6902
rect -106 6846 -38 6902
rect 18 6846 86 6902
rect 142 6846 210 6902
rect 266 6846 400 6902
rect -400 6778 400 6846
rect -400 6722 -286 6778
rect -230 6722 -162 6778
rect -106 6722 -38 6778
rect 18 6722 86 6778
rect 142 6722 210 6778
rect 266 6722 400 6778
rect -400 6654 400 6722
rect -400 6598 -286 6654
rect -230 6598 -162 6654
rect -106 6598 -38 6654
rect 18 6598 86 6654
rect 142 6598 210 6654
rect 266 6598 400 6654
rect -400 6530 400 6598
rect -400 6474 -286 6530
rect -230 6474 -162 6530
rect -106 6474 -38 6530
rect 18 6474 86 6530
rect 142 6474 210 6530
rect 266 6474 400 6530
rect -400 6406 400 6474
rect -400 6350 -286 6406
rect -230 6350 -162 6406
rect -106 6350 -38 6406
rect 18 6350 86 6406
rect 142 6350 210 6406
rect 266 6350 400 6406
rect -400 6282 400 6350
rect -400 6226 -286 6282
rect -230 6226 -162 6282
rect -106 6226 -38 6282
rect 18 6226 86 6282
rect 142 6226 210 6282
rect 266 6226 400 6282
rect -400 6158 400 6226
rect -400 6102 -286 6158
rect -230 6102 -162 6158
rect -106 6102 -38 6158
rect 18 6102 86 6158
rect 142 6102 210 6158
rect 266 6102 400 6158
rect -400 6034 400 6102
rect -400 5978 -286 6034
rect -230 5978 -162 6034
rect -106 5978 -38 6034
rect 18 5978 86 6034
rect 142 5978 210 6034
rect 266 5978 400 6034
rect -400 5910 400 5978
rect -400 5854 -286 5910
rect -230 5854 -162 5910
rect -106 5854 -38 5910
rect 18 5854 86 5910
rect 142 5854 210 5910
rect 266 5854 400 5910
rect -400 5786 400 5854
rect -400 5730 -286 5786
rect -230 5730 -162 5786
rect -106 5730 -38 5786
rect 18 5730 86 5786
rect 142 5730 210 5786
rect 266 5730 400 5786
rect -400 5662 400 5730
rect -400 5606 -286 5662
rect -230 5606 -162 5662
rect -106 5606 -38 5662
rect 18 5606 86 5662
rect 142 5606 210 5662
rect 266 5606 400 5662
rect -400 5538 400 5606
rect -400 5482 -286 5538
rect -230 5482 -162 5538
rect -106 5482 -38 5538
rect 18 5482 86 5538
rect 142 5482 210 5538
rect 266 5482 400 5538
rect -400 5414 400 5482
rect -400 5358 -286 5414
rect -230 5358 -162 5414
rect -106 5358 -38 5414
rect 18 5358 86 5414
rect 142 5358 210 5414
rect 266 5358 400 5414
rect -400 5290 400 5358
rect -400 5234 -286 5290
rect -230 5234 -162 5290
rect -106 5234 -38 5290
rect 18 5234 86 5290
rect 142 5234 210 5290
rect 266 5234 400 5290
rect -400 5166 400 5234
rect -400 5110 -286 5166
rect -230 5110 -162 5166
rect -106 5110 -38 5166
rect 18 5110 86 5166
rect 142 5110 210 5166
rect 266 5110 400 5166
rect -400 5042 400 5110
rect -400 4986 -286 5042
rect -230 4986 -162 5042
rect -106 4986 -38 5042
rect 18 4986 86 5042
rect 142 4986 210 5042
rect 266 4986 400 5042
rect -400 4918 400 4986
rect -400 4862 -286 4918
rect -230 4862 -162 4918
rect -106 4862 -38 4918
rect 18 4862 86 4918
rect 142 4862 210 4918
rect 266 4862 400 4918
rect -400 4794 400 4862
rect -400 4738 -286 4794
rect -230 4738 -162 4794
rect -106 4738 -38 4794
rect 18 4738 86 4794
rect 142 4738 210 4794
rect 266 4738 400 4794
rect -400 4670 400 4738
rect -400 4614 -286 4670
rect -230 4614 -162 4670
rect -106 4614 -38 4670
rect 18 4614 86 4670
rect 142 4614 210 4670
rect 266 4614 400 4670
rect -400 4546 400 4614
rect -400 4490 -286 4546
rect -230 4490 -162 4546
rect -106 4490 -38 4546
rect 18 4490 86 4546
rect 142 4490 210 4546
rect 266 4490 400 4546
rect -400 4422 400 4490
rect -400 4366 -286 4422
rect -230 4366 -162 4422
rect -106 4366 -38 4422
rect 18 4366 86 4422
rect 142 4366 210 4422
rect 266 4366 400 4422
rect -400 4298 400 4366
rect -400 4242 -286 4298
rect -230 4242 -162 4298
rect -106 4242 -38 4298
rect 18 4242 86 4298
rect 142 4242 210 4298
rect 266 4242 400 4298
rect -400 4174 400 4242
rect -400 4118 -286 4174
rect -230 4118 -162 4174
rect -106 4118 -38 4174
rect 18 4118 86 4174
rect 142 4118 210 4174
rect 266 4118 400 4174
rect -400 4050 400 4118
rect -400 3994 -286 4050
rect -230 3994 -162 4050
rect -106 3994 -38 4050
rect 18 3994 86 4050
rect 142 3994 210 4050
rect 266 3994 400 4050
rect -400 3926 400 3994
rect -400 3870 -286 3926
rect -230 3870 -162 3926
rect -106 3870 -38 3926
rect 18 3870 86 3926
rect 142 3870 210 3926
rect 266 3870 400 3926
rect -400 3802 400 3870
rect -400 3746 -286 3802
rect -230 3746 -162 3802
rect -106 3746 -38 3802
rect 18 3746 86 3802
rect 142 3746 210 3802
rect 266 3746 400 3802
rect -400 3678 400 3746
rect -400 3622 -286 3678
rect -230 3622 -162 3678
rect -106 3622 -38 3678
rect 18 3622 86 3678
rect 142 3622 210 3678
rect 266 3622 400 3678
rect -400 3554 400 3622
rect -400 3498 -286 3554
rect -230 3498 -162 3554
rect -106 3498 -38 3554
rect 18 3498 86 3554
rect 142 3498 210 3554
rect 266 3498 400 3554
rect -400 3430 400 3498
rect -400 3374 -286 3430
rect -230 3374 -162 3430
rect -106 3374 -38 3430
rect 18 3374 86 3430
rect 142 3374 210 3430
rect 266 3374 400 3430
rect -400 3306 400 3374
rect -400 3250 -286 3306
rect -230 3250 -162 3306
rect -106 3250 -38 3306
rect 18 3250 86 3306
rect 142 3250 210 3306
rect 266 3250 400 3306
rect -400 3182 400 3250
rect -400 3126 -286 3182
rect -230 3126 -162 3182
rect -106 3126 -38 3182
rect 18 3126 86 3182
rect 142 3126 210 3182
rect 266 3126 400 3182
rect -400 3058 400 3126
rect -400 3002 -286 3058
rect -230 3002 -162 3058
rect -106 3002 -38 3058
rect 18 3002 86 3058
rect 142 3002 210 3058
rect 266 3002 400 3058
rect -400 2934 400 3002
rect -400 2878 -286 2934
rect -230 2878 -162 2934
rect -106 2878 -38 2934
rect 18 2878 86 2934
rect 142 2878 210 2934
rect 266 2878 400 2934
rect -400 2810 400 2878
rect -400 2754 -286 2810
rect -230 2754 -162 2810
rect -106 2754 -38 2810
rect 18 2754 86 2810
rect 142 2754 210 2810
rect 266 2754 400 2810
rect -400 2686 400 2754
rect -400 2630 -286 2686
rect -230 2630 -162 2686
rect -106 2630 -38 2686
rect 18 2630 86 2686
rect 142 2630 210 2686
rect 266 2630 400 2686
rect -400 2562 400 2630
rect -400 2506 -286 2562
rect -230 2506 -162 2562
rect -106 2506 -38 2562
rect 18 2506 86 2562
rect 142 2506 210 2562
rect 266 2506 400 2562
rect -400 2438 400 2506
rect -400 2382 -286 2438
rect -230 2382 -162 2438
rect -106 2382 -38 2438
rect 18 2382 86 2438
rect 142 2382 210 2438
rect 266 2382 400 2438
rect -400 2314 400 2382
rect -400 2258 -286 2314
rect -230 2258 -162 2314
rect -106 2258 -38 2314
rect 18 2258 86 2314
rect 142 2258 210 2314
rect 266 2258 400 2314
rect -400 2190 400 2258
rect -400 2134 -286 2190
rect -230 2134 -162 2190
rect -106 2134 -38 2190
rect 18 2134 86 2190
rect 142 2134 210 2190
rect 266 2134 400 2190
rect -400 2066 400 2134
rect -400 2010 -286 2066
rect -230 2010 -162 2066
rect -106 2010 -38 2066
rect 18 2010 86 2066
rect 142 2010 210 2066
rect 266 2010 400 2066
rect -400 1942 400 2010
rect -400 1886 -286 1942
rect -230 1886 -162 1942
rect -106 1886 -38 1942
rect 18 1886 86 1942
rect 142 1886 210 1942
rect 266 1886 400 1942
rect -400 1818 400 1886
rect -400 1762 -286 1818
rect -230 1762 -162 1818
rect -106 1762 -38 1818
rect 18 1762 86 1818
rect 142 1762 210 1818
rect 266 1762 400 1818
rect -400 1694 400 1762
rect -400 1638 -286 1694
rect -230 1638 -162 1694
rect -106 1638 -38 1694
rect 18 1638 86 1694
rect 142 1638 210 1694
rect 266 1638 400 1694
rect -400 1570 400 1638
rect -400 1514 -286 1570
rect -230 1514 -162 1570
rect -106 1514 -38 1570
rect 18 1514 86 1570
rect 142 1514 210 1570
rect 266 1514 400 1570
rect -400 1446 400 1514
rect -400 1390 -286 1446
rect -230 1390 -162 1446
rect -106 1390 -38 1446
rect 18 1390 86 1446
rect 142 1390 210 1446
rect 266 1390 400 1446
rect -400 1322 400 1390
rect -400 1266 -286 1322
rect -230 1266 -162 1322
rect -106 1266 -38 1322
rect 18 1266 86 1322
rect 142 1266 210 1322
rect 266 1266 400 1322
rect -400 1198 400 1266
rect -400 1142 -286 1198
rect -230 1142 -162 1198
rect -106 1142 -38 1198
rect 18 1142 86 1198
rect 142 1142 210 1198
rect 266 1142 400 1198
rect -400 1074 400 1142
rect -400 1018 -286 1074
rect -230 1018 -162 1074
rect -106 1018 -38 1074
rect 18 1018 86 1074
rect 142 1018 210 1074
rect 266 1018 400 1074
rect -400 950 400 1018
rect -400 894 -286 950
rect -230 894 -162 950
rect -106 894 -38 950
rect 18 894 86 950
rect 142 894 210 950
rect 266 894 400 950
rect -400 826 400 894
rect -400 770 -286 826
rect -230 770 -162 826
rect -106 770 -38 826
rect 18 770 86 826
rect 142 770 210 826
rect 266 770 400 826
rect -400 702 400 770
rect -400 646 -286 702
rect -230 646 -162 702
rect -106 646 -38 702
rect 18 646 86 702
rect 142 646 210 702
rect 266 646 400 702
rect -400 578 400 646
rect -400 522 -286 578
rect -230 522 -162 578
rect -106 522 -38 578
rect 18 522 86 578
rect 142 522 210 578
rect 266 522 400 578
rect -400 454 400 522
rect -400 398 -286 454
rect -230 398 -162 454
rect -106 398 -38 454
rect 18 398 86 454
rect 142 398 210 454
rect 266 400 400 454
rect 668 12310 1008 12400
rect 668 12254 741 12310
rect 797 12254 883 12310
rect 939 12254 1008 12310
rect 668 12168 1008 12254
rect 668 12112 741 12168
rect 797 12112 883 12168
rect 939 12112 1008 12168
rect 668 12026 1008 12112
rect 668 11970 741 12026
rect 797 11970 883 12026
rect 939 11970 1008 12026
rect 668 11884 1008 11970
rect 668 11828 741 11884
rect 797 11828 883 11884
rect 939 11828 1008 11884
rect 668 11742 1008 11828
rect 668 11686 741 11742
rect 797 11686 883 11742
rect 939 11686 1008 11742
rect 668 11600 1008 11686
rect 668 11544 741 11600
rect 797 11544 883 11600
rect 939 11544 1008 11600
rect 668 11458 1008 11544
rect 668 11402 741 11458
rect 797 11402 883 11458
rect 939 11402 1008 11458
rect 668 11316 1008 11402
rect 668 11260 741 11316
rect 797 11260 883 11316
rect 939 11260 1008 11316
rect 668 11174 1008 11260
rect 668 11118 741 11174
rect 797 11118 883 11174
rect 939 11118 1008 11174
rect 668 11032 1008 11118
rect 668 10976 741 11032
rect 797 10976 883 11032
rect 939 10976 1008 11032
rect 668 10890 1008 10976
rect 668 10834 741 10890
rect 797 10834 883 10890
rect 939 10834 1008 10890
rect 668 10748 1008 10834
rect 668 10692 741 10748
rect 797 10692 883 10748
rect 939 10692 1008 10748
rect 668 10606 1008 10692
rect 668 10550 741 10606
rect 797 10550 883 10606
rect 939 10550 1008 10606
rect 668 10464 1008 10550
rect 668 10408 741 10464
rect 797 10408 883 10464
rect 939 10408 1008 10464
rect 668 10322 1008 10408
rect 668 10266 741 10322
rect 797 10266 883 10322
rect 939 10266 1008 10322
rect 668 10180 1008 10266
rect 668 10124 741 10180
rect 797 10124 883 10180
rect 939 10124 1008 10180
rect 668 10038 1008 10124
rect 668 9982 741 10038
rect 797 9982 883 10038
rect 939 9982 1008 10038
rect 668 9896 1008 9982
rect 668 9840 741 9896
rect 797 9840 883 9896
rect 939 9840 1008 9896
rect 668 9754 1008 9840
rect 668 9698 741 9754
rect 797 9698 883 9754
rect 939 9698 1008 9754
rect 668 9612 1008 9698
rect 668 9556 741 9612
rect 797 9556 883 9612
rect 939 9556 1008 9612
rect 668 9470 1008 9556
rect 668 9414 741 9470
rect 797 9414 883 9470
rect 939 9414 1008 9470
rect 668 9328 1008 9414
rect 668 9272 741 9328
rect 797 9272 883 9328
rect 939 9272 1008 9328
rect 668 9186 1008 9272
rect 668 9130 741 9186
rect 797 9130 883 9186
rect 939 9130 1008 9186
rect 668 9044 1008 9130
rect 668 8988 741 9044
rect 797 8988 883 9044
rect 939 8988 1008 9044
rect 668 8902 1008 8988
rect 668 8846 741 8902
rect 797 8846 883 8902
rect 939 8846 1008 8902
rect 668 8760 1008 8846
rect 668 8704 741 8760
rect 797 8704 883 8760
rect 939 8704 1008 8760
rect 668 8618 1008 8704
rect 668 8562 741 8618
rect 797 8562 883 8618
rect 939 8562 1008 8618
rect 668 8476 1008 8562
rect 668 8420 741 8476
rect 797 8420 883 8476
rect 939 8420 1008 8476
rect 668 8334 1008 8420
rect 668 8278 741 8334
rect 797 8278 883 8334
rect 939 8278 1008 8334
rect 668 8192 1008 8278
rect 668 8136 741 8192
rect 797 8136 883 8192
rect 939 8136 1008 8192
rect 668 8050 1008 8136
rect 668 7994 741 8050
rect 797 7994 883 8050
rect 939 7994 1008 8050
rect 668 7908 1008 7994
rect 668 7852 741 7908
rect 797 7852 883 7908
rect 939 7852 1008 7908
rect 668 7766 1008 7852
rect 668 7710 741 7766
rect 797 7710 883 7766
rect 939 7710 1008 7766
rect 668 7624 1008 7710
rect 668 7568 741 7624
rect 797 7568 883 7624
rect 939 7568 1008 7624
rect 668 7482 1008 7568
rect 668 7426 741 7482
rect 797 7426 883 7482
rect 939 7426 1008 7482
rect 668 7340 1008 7426
rect 668 7284 741 7340
rect 797 7284 883 7340
rect 939 7284 1008 7340
rect 668 7198 1008 7284
rect 668 7142 741 7198
rect 797 7142 883 7198
rect 939 7142 1008 7198
rect 668 7056 1008 7142
rect 668 7000 741 7056
rect 797 7000 883 7056
rect 939 7000 1008 7056
rect 668 6914 1008 7000
rect 668 6858 741 6914
rect 797 6858 883 6914
rect 939 6858 1008 6914
rect 668 6772 1008 6858
rect 668 6716 741 6772
rect 797 6716 883 6772
rect 939 6716 1008 6772
rect 668 6630 1008 6716
rect 668 6574 741 6630
rect 797 6574 883 6630
rect 939 6574 1008 6630
rect 668 6488 1008 6574
rect 668 6432 741 6488
rect 797 6432 883 6488
rect 939 6432 1008 6488
rect 668 6346 1008 6432
rect 668 6290 741 6346
rect 797 6290 883 6346
rect 939 6290 1008 6346
rect 668 6204 1008 6290
rect 668 6148 741 6204
rect 797 6148 883 6204
rect 939 6148 1008 6204
rect 668 6062 1008 6148
rect 668 6006 741 6062
rect 797 6006 883 6062
rect 939 6006 1008 6062
rect 668 5920 1008 6006
rect 668 5864 741 5920
rect 797 5864 883 5920
rect 939 5864 1008 5920
rect 668 5778 1008 5864
rect 668 5722 741 5778
rect 797 5722 883 5778
rect 939 5722 1008 5778
rect 668 5636 1008 5722
rect 668 5580 741 5636
rect 797 5580 883 5636
rect 939 5580 1008 5636
rect 668 5494 1008 5580
rect 668 5438 741 5494
rect 797 5438 883 5494
rect 939 5438 1008 5494
rect 668 5352 1008 5438
rect 668 5296 741 5352
rect 797 5296 883 5352
rect 939 5296 1008 5352
rect 668 5210 1008 5296
rect 668 5154 741 5210
rect 797 5154 883 5210
rect 939 5154 1008 5210
rect 668 5068 1008 5154
rect 668 5012 741 5068
rect 797 5012 883 5068
rect 939 5012 1008 5068
rect 668 4926 1008 5012
rect 668 4870 741 4926
rect 797 4870 883 4926
rect 939 4870 1008 4926
rect 668 4784 1008 4870
rect 668 4728 741 4784
rect 797 4728 883 4784
rect 939 4728 1008 4784
rect 668 4642 1008 4728
rect 668 4586 741 4642
rect 797 4586 883 4642
rect 939 4586 1008 4642
rect 668 4500 1008 4586
rect 668 4444 741 4500
rect 797 4444 883 4500
rect 939 4444 1008 4500
rect 668 4358 1008 4444
rect 668 4302 741 4358
rect 797 4302 883 4358
rect 939 4302 1008 4358
rect 668 4216 1008 4302
rect 668 4160 741 4216
rect 797 4160 883 4216
rect 939 4160 1008 4216
rect 668 4074 1008 4160
rect 668 4018 741 4074
rect 797 4018 883 4074
rect 939 4018 1008 4074
rect 668 3932 1008 4018
rect 668 3876 741 3932
rect 797 3876 883 3932
rect 939 3876 1008 3932
rect 668 3790 1008 3876
rect 668 3734 741 3790
rect 797 3734 883 3790
rect 939 3734 1008 3790
rect 668 3648 1008 3734
rect 668 3592 741 3648
rect 797 3592 883 3648
rect 939 3592 1008 3648
rect 668 3506 1008 3592
rect 668 3450 741 3506
rect 797 3450 883 3506
rect 939 3450 1008 3506
rect 668 3364 1008 3450
rect 668 3308 741 3364
rect 797 3308 883 3364
rect 939 3308 1008 3364
rect 668 3222 1008 3308
rect 668 3166 741 3222
rect 797 3166 883 3222
rect 939 3166 1008 3222
rect 668 3080 1008 3166
rect 668 3024 741 3080
rect 797 3024 883 3080
rect 939 3024 1008 3080
rect 668 2938 1008 3024
rect 668 2882 741 2938
rect 797 2882 883 2938
rect 939 2882 1008 2938
rect 668 2796 1008 2882
rect 668 2740 741 2796
rect 797 2740 883 2796
rect 939 2740 1008 2796
rect 668 2654 1008 2740
rect 668 2598 741 2654
rect 797 2598 883 2654
rect 939 2598 1008 2654
rect 668 2512 1008 2598
rect 668 2456 741 2512
rect 797 2456 883 2512
rect 939 2456 1008 2512
rect 668 2370 1008 2456
rect 668 2314 741 2370
rect 797 2314 883 2370
rect 939 2314 1008 2370
rect 668 2228 1008 2314
rect 668 2172 741 2228
rect 797 2172 883 2228
rect 939 2172 1008 2228
rect 668 2086 1008 2172
rect 668 2030 741 2086
rect 797 2030 883 2086
rect 939 2030 1008 2086
rect 668 1944 1008 2030
rect 668 1888 741 1944
rect 797 1888 883 1944
rect 939 1888 1008 1944
rect 668 1802 1008 1888
rect 668 1746 741 1802
rect 797 1746 883 1802
rect 939 1746 1008 1802
rect 668 1660 1008 1746
rect 668 1604 741 1660
rect 797 1604 883 1660
rect 939 1604 1008 1660
rect 668 1518 1008 1604
rect 668 1462 741 1518
rect 797 1462 883 1518
rect 939 1462 1008 1518
rect 668 1376 1008 1462
rect 668 1320 741 1376
rect 797 1320 883 1376
rect 939 1320 1008 1376
rect 668 1234 1008 1320
rect 668 1178 741 1234
rect 797 1178 883 1234
rect 939 1178 1008 1234
rect 668 1092 1008 1178
rect 668 1036 741 1092
rect 797 1036 883 1092
rect 939 1036 1008 1092
rect 668 950 1008 1036
rect 668 894 741 950
rect 797 894 883 950
rect 939 894 1008 950
rect 668 808 1008 894
rect 668 752 741 808
rect 797 752 883 808
rect 939 752 1008 808
rect 668 666 1008 752
rect 668 610 741 666
rect 797 610 883 666
rect 939 610 1008 666
rect 668 524 1008 610
rect 668 468 741 524
rect 797 468 883 524
rect 939 468 1008 524
rect 668 400 1008 468
rect 1068 12310 1408 12400
rect 1068 12254 1142 12310
rect 1198 12254 1284 12310
rect 1340 12254 1408 12310
rect 1068 12168 1408 12254
rect 1068 12112 1142 12168
rect 1198 12112 1284 12168
rect 1340 12112 1408 12168
rect 1068 12026 1408 12112
rect 1068 11970 1142 12026
rect 1198 11970 1284 12026
rect 1340 11970 1408 12026
rect 1068 11884 1408 11970
rect 1068 11828 1142 11884
rect 1198 11828 1284 11884
rect 1340 11828 1408 11884
rect 1068 11742 1408 11828
rect 1068 11686 1142 11742
rect 1198 11686 1284 11742
rect 1340 11686 1408 11742
rect 1068 11600 1408 11686
rect 1068 11544 1142 11600
rect 1198 11544 1284 11600
rect 1340 11544 1408 11600
rect 1068 11458 1408 11544
rect 1068 11402 1142 11458
rect 1198 11402 1284 11458
rect 1340 11402 1408 11458
rect 1068 11316 1408 11402
rect 1068 11260 1142 11316
rect 1198 11260 1284 11316
rect 1340 11260 1408 11316
rect 1068 11174 1408 11260
rect 1068 11118 1142 11174
rect 1198 11118 1284 11174
rect 1340 11118 1408 11174
rect 1068 11032 1408 11118
rect 1068 10976 1142 11032
rect 1198 10976 1284 11032
rect 1340 10976 1408 11032
rect 1068 10890 1408 10976
rect 1068 10834 1142 10890
rect 1198 10834 1284 10890
rect 1340 10834 1408 10890
rect 1068 10748 1408 10834
rect 1068 10692 1142 10748
rect 1198 10692 1284 10748
rect 1340 10692 1408 10748
rect 1068 10606 1408 10692
rect 1068 10550 1142 10606
rect 1198 10550 1284 10606
rect 1340 10550 1408 10606
rect 1068 10464 1408 10550
rect 1068 10408 1142 10464
rect 1198 10408 1284 10464
rect 1340 10408 1408 10464
rect 1068 10322 1408 10408
rect 1068 10266 1142 10322
rect 1198 10266 1284 10322
rect 1340 10266 1408 10322
rect 1068 10180 1408 10266
rect 1068 10124 1142 10180
rect 1198 10124 1284 10180
rect 1340 10124 1408 10180
rect 1068 10038 1408 10124
rect 1068 9982 1142 10038
rect 1198 9982 1284 10038
rect 1340 9982 1408 10038
rect 1068 9896 1408 9982
rect 1068 9840 1142 9896
rect 1198 9840 1284 9896
rect 1340 9840 1408 9896
rect 1068 9754 1408 9840
rect 1068 9698 1142 9754
rect 1198 9698 1284 9754
rect 1340 9698 1408 9754
rect 1068 9612 1408 9698
rect 1068 9556 1142 9612
rect 1198 9556 1284 9612
rect 1340 9556 1408 9612
rect 1068 9470 1408 9556
rect 1068 9414 1142 9470
rect 1198 9414 1284 9470
rect 1340 9414 1408 9470
rect 1068 9328 1408 9414
rect 1068 9272 1142 9328
rect 1198 9272 1284 9328
rect 1340 9272 1408 9328
rect 1068 9186 1408 9272
rect 1068 9130 1142 9186
rect 1198 9130 1284 9186
rect 1340 9130 1408 9186
rect 1068 9044 1408 9130
rect 1068 8988 1142 9044
rect 1198 8988 1284 9044
rect 1340 8988 1408 9044
rect 1068 8902 1408 8988
rect 1068 8846 1142 8902
rect 1198 8846 1284 8902
rect 1340 8846 1408 8902
rect 1068 8760 1408 8846
rect 1068 8704 1142 8760
rect 1198 8704 1284 8760
rect 1340 8704 1408 8760
rect 1068 8618 1408 8704
rect 1068 8562 1142 8618
rect 1198 8562 1284 8618
rect 1340 8562 1408 8618
rect 1068 8476 1408 8562
rect 1068 8420 1142 8476
rect 1198 8420 1284 8476
rect 1340 8420 1408 8476
rect 1068 8334 1408 8420
rect 1068 8278 1142 8334
rect 1198 8278 1284 8334
rect 1340 8278 1408 8334
rect 1068 8192 1408 8278
rect 1068 8136 1142 8192
rect 1198 8136 1284 8192
rect 1340 8136 1408 8192
rect 1068 8050 1408 8136
rect 1068 7994 1142 8050
rect 1198 7994 1284 8050
rect 1340 7994 1408 8050
rect 1068 7908 1408 7994
rect 1068 7852 1142 7908
rect 1198 7852 1284 7908
rect 1340 7852 1408 7908
rect 1068 7766 1408 7852
rect 1068 7710 1142 7766
rect 1198 7710 1284 7766
rect 1340 7710 1408 7766
rect 1068 7624 1408 7710
rect 1068 7568 1142 7624
rect 1198 7568 1284 7624
rect 1340 7568 1408 7624
rect 1068 7482 1408 7568
rect 1068 7426 1142 7482
rect 1198 7426 1284 7482
rect 1340 7426 1408 7482
rect 1068 7340 1408 7426
rect 1068 7284 1142 7340
rect 1198 7284 1284 7340
rect 1340 7284 1408 7340
rect 1068 7198 1408 7284
rect 1068 7142 1142 7198
rect 1198 7142 1284 7198
rect 1340 7142 1408 7198
rect 1068 7056 1408 7142
rect 1068 7000 1142 7056
rect 1198 7000 1284 7056
rect 1340 7000 1408 7056
rect 1068 6914 1408 7000
rect 1068 6858 1142 6914
rect 1198 6858 1284 6914
rect 1340 6858 1408 6914
rect 1068 6772 1408 6858
rect 1068 6716 1142 6772
rect 1198 6716 1284 6772
rect 1340 6716 1408 6772
rect 1068 6630 1408 6716
rect 1068 6574 1142 6630
rect 1198 6574 1284 6630
rect 1340 6574 1408 6630
rect 1068 6488 1408 6574
rect 1068 6432 1142 6488
rect 1198 6432 1284 6488
rect 1340 6432 1408 6488
rect 1068 6346 1408 6432
rect 1068 6290 1142 6346
rect 1198 6290 1284 6346
rect 1340 6290 1408 6346
rect 1068 6204 1408 6290
rect 1068 6148 1142 6204
rect 1198 6148 1284 6204
rect 1340 6148 1408 6204
rect 1068 6062 1408 6148
rect 1068 6006 1142 6062
rect 1198 6006 1284 6062
rect 1340 6006 1408 6062
rect 1068 5920 1408 6006
rect 1068 5864 1142 5920
rect 1198 5864 1284 5920
rect 1340 5864 1408 5920
rect 1068 5778 1408 5864
rect 1068 5722 1142 5778
rect 1198 5722 1284 5778
rect 1340 5722 1408 5778
rect 1068 5636 1408 5722
rect 1068 5580 1142 5636
rect 1198 5580 1284 5636
rect 1340 5580 1408 5636
rect 1068 5494 1408 5580
rect 1068 5438 1142 5494
rect 1198 5438 1284 5494
rect 1340 5438 1408 5494
rect 1068 5352 1408 5438
rect 1068 5296 1142 5352
rect 1198 5296 1284 5352
rect 1340 5296 1408 5352
rect 1068 5210 1408 5296
rect 1068 5154 1142 5210
rect 1198 5154 1284 5210
rect 1340 5154 1408 5210
rect 1068 5068 1408 5154
rect 1068 5012 1142 5068
rect 1198 5012 1284 5068
rect 1340 5012 1408 5068
rect 1068 4926 1408 5012
rect 1068 4870 1142 4926
rect 1198 4870 1284 4926
rect 1340 4870 1408 4926
rect 1068 4784 1408 4870
rect 1068 4728 1142 4784
rect 1198 4728 1284 4784
rect 1340 4728 1408 4784
rect 1068 4642 1408 4728
rect 1068 4586 1142 4642
rect 1198 4586 1284 4642
rect 1340 4586 1408 4642
rect 1068 4500 1408 4586
rect 1068 4444 1142 4500
rect 1198 4444 1284 4500
rect 1340 4444 1408 4500
rect 1068 4358 1408 4444
rect 1068 4302 1142 4358
rect 1198 4302 1284 4358
rect 1340 4302 1408 4358
rect 1068 4216 1408 4302
rect 1068 4160 1142 4216
rect 1198 4160 1284 4216
rect 1340 4160 1408 4216
rect 1068 4074 1408 4160
rect 1068 4018 1142 4074
rect 1198 4018 1284 4074
rect 1340 4018 1408 4074
rect 1068 3932 1408 4018
rect 1068 3876 1142 3932
rect 1198 3876 1284 3932
rect 1340 3876 1408 3932
rect 1068 3790 1408 3876
rect 1068 3734 1142 3790
rect 1198 3734 1284 3790
rect 1340 3734 1408 3790
rect 1068 3648 1408 3734
rect 1068 3592 1142 3648
rect 1198 3592 1284 3648
rect 1340 3592 1408 3648
rect 1068 3506 1408 3592
rect 1068 3450 1142 3506
rect 1198 3450 1284 3506
rect 1340 3450 1408 3506
rect 1068 3364 1408 3450
rect 1068 3308 1142 3364
rect 1198 3308 1284 3364
rect 1340 3308 1408 3364
rect 1068 3222 1408 3308
rect 1068 3166 1142 3222
rect 1198 3166 1284 3222
rect 1340 3166 1408 3222
rect 1068 3080 1408 3166
rect 1068 3024 1142 3080
rect 1198 3024 1284 3080
rect 1340 3024 1408 3080
rect 1068 2938 1408 3024
rect 1068 2882 1142 2938
rect 1198 2882 1284 2938
rect 1340 2882 1408 2938
rect 1068 2796 1408 2882
rect 1068 2740 1142 2796
rect 1198 2740 1284 2796
rect 1340 2740 1408 2796
rect 1068 2654 1408 2740
rect 1068 2598 1142 2654
rect 1198 2598 1284 2654
rect 1340 2598 1408 2654
rect 1068 2512 1408 2598
rect 1068 2456 1142 2512
rect 1198 2456 1284 2512
rect 1340 2456 1408 2512
rect 1068 2370 1408 2456
rect 1068 2314 1142 2370
rect 1198 2314 1284 2370
rect 1340 2314 1408 2370
rect 1068 2228 1408 2314
rect 1068 2172 1142 2228
rect 1198 2172 1284 2228
rect 1340 2172 1408 2228
rect 1068 2086 1408 2172
rect 1068 2030 1142 2086
rect 1198 2030 1284 2086
rect 1340 2030 1408 2086
rect 1068 1944 1408 2030
rect 1068 1888 1142 1944
rect 1198 1888 1284 1944
rect 1340 1888 1408 1944
rect 1068 1802 1408 1888
rect 1068 1746 1142 1802
rect 1198 1746 1284 1802
rect 1340 1746 1408 1802
rect 1068 1660 1408 1746
rect 1068 1604 1142 1660
rect 1198 1604 1284 1660
rect 1340 1604 1408 1660
rect 1068 1518 1408 1604
rect 1068 1462 1142 1518
rect 1198 1462 1284 1518
rect 1340 1462 1408 1518
rect 1068 1376 1408 1462
rect 1068 1320 1142 1376
rect 1198 1320 1284 1376
rect 1340 1320 1408 1376
rect 1068 1234 1408 1320
rect 1068 1178 1142 1234
rect 1198 1178 1284 1234
rect 1340 1178 1408 1234
rect 1068 1092 1408 1178
rect 1068 1036 1142 1092
rect 1198 1036 1284 1092
rect 1340 1036 1408 1092
rect 1068 950 1408 1036
rect 1068 894 1142 950
rect 1198 894 1284 950
rect 1340 894 1408 950
rect 1068 808 1408 894
rect 1068 752 1142 808
rect 1198 752 1284 808
rect 1340 752 1408 808
rect 1068 666 1408 752
rect 1068 610 1142 666
rect 1198 610 1284 666
rect 1340 610 1408 666
rect 1068 524 1408 610
rect 1068 468 1142 524
rect 1198 468 1284 524
rect 1340 468 1408 524
rect 1068 400 1408 468
rect 1468 12310 1808 12400
rect 1468 12254 1542 12310
rect 1598 12254 1684 12310
rect 1740 12254 1808 12310
rect 1468 12168 1808 12254
rect 1468 12112 1542 12168
rect 1598 12112 1684 12168
rect 1740 12112 1808 12168
rect 1468 12026 1808 12112
rect 1468 11970 1542 12026
rect 1598 11970 1684 12026
rect 1740 11970 1808 12026
rect 1468 11884 1808 11970
rect 1468 11828 1542 11884
rect 1598 11828 1684 11884
rect 1740 11828 1808 11884
rect 1468 11742 1808 11828
rect 1468 11686 1542 11742
rect 1598 11686 1684 11742
rect 1740 11686 1808 11742
rect 1468 11600 1808 11686
rect 1468 11544 1542 11600
rect 1598 11544 1684 11600
rect 1740 11544 1808 11600
rect 1468 11458 1808 11544
rect 1468 11402 1542 11458
rect 1598 11402 1684 11458
rect 1740 11402 1808 11458
rect 1468 11316 1808 11402
rect 1468 11260 1542 11316
rect 1598 11260 1684 11316
rect 1740 11260 1808 11316
rect 1468 11174 1808 11260
rect 1468 11118 1542 11174
rect 1598 11118 1684 11174
rect 1740 11118 1808 11174
rect 1468 11032 1808 11118
rect 1468 10976 1542 11032
rect 1598 10976 1684 11032
rect 1740 10976 1808 11032
rect 1468 10890 1808 10976
rect 1468 10834 1542 10890
rect 1598 10834 1684 10890
rect 1740 10834 1808 10890
rect 1468 10748 1808 10834
rect 1468 10692 1542 10748
rect 1598 10692 1684 10748
rect 1740 10692 1808 10748
rect 1468 10606 1808 10692
rect 1468 10550 1542 10606
rect 1598 10550 1684 10606
rect 1740 10550 1808 10606
rect 1468 10464 1808 10550
rect 1468 10408 1542 10464
rect 1598 10408 1684 10464
rect 1740 10408 1808 10464
rect 1468 10322 1808 10408
rect 1468 10266 1542 10322
rect 1598 10266 1684 10322
rect 1740 10266 1808 10322
rect 1468 10180 1808 10266
rect 1468 10124 1542 10180
rect 1598 10124 1684 10180
rect 1740 10124 1808 10180
rect 1468 10038 1808 10124
rect 1468 9982 1542 10038
rect 1598 9982 1684 10038
rect 1740 9982 1808 10038
rect 1468 9896 1808 9982
rect 1468 9840 1542 9896
rect 1598 9840 1684 9896
rect 1740 9840 1808 9896
rect 1468 9754 1808 9840
rect 1468 9698 1542 9754
rect 1598 9698 1684 9754
rect 1740 9698 1808 9754
rect 1468 9612 1808 9698
rect 1468 9556 1542 9612
rect 1598 9556 1684 9612
rect 1740 9556 1808 9612
rect 1468 9470 1808 9556
rect 1468 9414 1542 9470
rect 1598 9414 1684 9470
rect 1740 9414 1808 9470
rect 1468 9328 1808 9414
rect 1468 9272 1542 9328
rect 1598 9272 1684 9328
rect 1740 9272 1808 9328
rect 1468 9186 1808 9272
rect 1468 9130 1542 9186
rect 1598 9130 1684 9186
rect 1740 9130 1808 9186
rect 1468 9044 1808 9130
rect 1468 8988 1542 9044
rect 1598 8988 1684 9044
rect 1740 8988 1808 9044
rect 1468 8902 1808 8988
rect 1468 8846 1542 8902
rect 1598 8846 1684 8902
rect 1740 8846 1808 8902
rect 1468 8760 1808 8846
rect 1468 8704 1542 8760
rect 1598 8704 1684 8760
rect 1740 8704 1808 8760
rect 1468 8618 1808 8704
rect 1468 8562 1542 8618
rect 1598 8562 1684 8618
rect 1740 8562 1808 8618
rect 1468 8476 1808 8562
rect 1468 8420 1542 8476
rect 1598 8420 1684 8476
rect 1740 8420 1808 8476
rect 1468 8334 1808 8420
rect 1468 8278 1542 8334
rect 1598 8278 1684 8334
rect 1740 8278 1808 8334
rect 1468 8192 1808 8278
rect 1468 8136 1542 8192
rect 1598 8136 1684 8192
rect 1740 8136 1808 8192
rect 1468 8050 1808 8136
rect 1468 7994 1542 8050
rect 1598 7994 1684 8050
rect 1740 7994 1808 8050
rect 1468 7908 1808 7994
rect 1468 7852 1542 7908
rect 1598 7852 1684 7908
rect 1740 7852 1808 7908
rect 1468 7766 1808 7852
rect 1468 7710 1542 7766
rect 1598 7710 1684 7766
rect 1740 7710 1808 7766
rect 1468 7624 1808 7710
rect 1468 7568 1542 7624
rect 1598 7568 1684 7624
rect 1740 7568 1808 7624
rect 1468 7482 1808 7568
rect 1468 7426 1542 7482
rect 1598 7426 1684 7482
rect 1740 7426 1808 7482
rect 1468 7340 1808 7426
rect 1468 7284 1542 7340
rect 1598 7284 1684 7340
rect 1740 7284 1808 7340
rect 1468 7198 1808 7284
rect 1468 7142 1542 7198
rect 1598 7142 1684 7198
rect 1740 7142 1808 7198
rect 1468 7056 1808 7142
rect 1468 7000 1542 7056
rect 1598 7000 1684 7056
rect 1740 7000 1808 7056
rect 1468 6914 1808 7000
rect 1468 6858 1542 6914
rect 1598 6858 1684 6914
rect 1740 6858 1808 6914
rect 1468 6772 1808 6858
rect 1468 6716 1542 6772
rect 1598 6716 1684 6772
rect 1740 6716 1808 6772
rect 1468 6630 1808 6716
rect 1468 6574 1542 6630
rect 1598 6574 1684 6630
rect 1740 6574 1808 6630
rect 1468 6488 1808 6574
rect 1468 6432 1542 6488
rect 1598 6432 1684 6488
rect 1740 6432 1808 6488
rect 1468 6346 1808 6432
rect 1468 6290 1542 6346
rect 1598 6290 1684 6346
rect 1740 6290 1808 6346
rect 1468 6204 1808 6290
rect 1468 6148 1542 6204
rect 1598 6148 1684 6204
rect 1740 6148 1808 6204
rect 1468 6062 1808 6148
rect 1468 6006 1542 6062
rect 1598 6006 1684 6062
rect 1740 6006 1808 6062
rect 1468 5920 1808 6006
rect 1468 5864 1542 5920
rect 1598 5864 1684 5920
rect 1740 5864 1808 5920
rect 1468 5778 1808 5864
rect 1468 5722 1542 5778
rect 1598 5722 1684 5778
rect 1740 5722 1808 5778
rect 1468 5636 1808 5722
rect 1468 5580 1542 5636
rect 1598 5580 1684 5636
rect 1740 5580 1808 5636
rect 1468 5494 1808 5580
rect 1468 5438 1542 5494
rect 1598 5438 1684 5494
rect 1740 5438 1808 5494
rect 1468 5352 1808 5438
rect 1468 5296 1542 5352
rect 1598 5296 1684 5352
rect 1740 5296 1808 5352
rect 1468 5210 1808 5296
rect 1468 5154 1542 5210
rect 1598 5154 1684 5210
rect 1740 5154 1808 5210
rect 1468 5068 1808 5154
rect 1468 5012 1542 5068
rect 1598 5012 1684 5068
rect 1740 5012 1808 5068
rect 1468 4926 1808 5012
rect 1468 4870 1542 4926
rect 1598 4870 1684 4926
rect 1740 4870 1808 4926
rect 1468 4784 1808 4870
rect 1468 4728 1542 4784
rect 1598 4728 1684 4784
rect 1740 4728 1808 4784
rect 1468 4642 1808 4728
rect 1468 4586 1542 4642
rect 1598 4586 1684 4642
rect 1740 4586 1808 4642
rect 1468 4500 1808 4586
rect 1468 4444 1542 4500
rect 1598 4444 1684 4500
rect 1740 4444 1808 4500
rect 1468 4358 1808 4444
rect 1468 4302 1542 4358
rect 1598 4302 1684 4358
rect 1740 4302 1808 4358
rect 1468 4216 1808 4302
rect 1468 4160 1542 4216
rect 1598 4160 1684 4216
rect 1740 4160 1808 4216
rect 1468 4074 1808 4160
rect 1468 4018 1542 4074
rect 1598 4018 1684 4074
rect 1740 4018 1808 4074
rect 1468 3932 1808 4018
rect 1468 3876 1542 3932
rect 1598 3876 1684 3932
rect 1740 3876 1808 3932
rect 1468 3790 1808 3876
rect 1468 3734 1542 3790
rect 1598 3734 1684 3790
rect 1740 3734 1808 3790
rect 1468 3648 1808 3734
rect 1468 3592 1542 3648
rect 1598 3592 1684 3648
rect 1740 3592 1808 3648
rect 1468 3506 1808 3592
rect 1468 3450 1542 3506
rect 1598 3450 1684 3506
rect 1740 3450 1808 3506
rect 1468 3364 1808 3450
rect 1468 3308 1542 3364
rect 1598 3308 1684 3364
rect 1740 3308 1808 3364
rect 1468 3222 1808 3308
rect 1468 3166 1542 3222
rect 1598 3166 1684 3222
rect 1740 3166 1808 3222
rect 1468 3080 1808 3166
rect 1468 3024 1542 3080
rect 1598 3024 1684 3080
rect 1740 3024 1808 3080
rect 1468 2938 1808 3024
rect 1468 2882 1542 2938
rect 1598 2882 1684 2938
rect 1740 2882 1808 2938
rect 1468 2796 1808 2882
rect 1468 2740 1542 2796
rect 1598 2740 1684 2796
rect 1740 2740 1808 2796
rect 1468 2654 1808 2740
rect 1468 2598 1542 2654
rect 1598 2598 1684 2654
rect 1740 2598 1808 2654
rect 1468 2512 1808 2598
rect 1468 2456 1542 2512
rect 1598 2456 1684 2512
rect 1740 2456 1808 2512
rect 1468 2370 1808 2456
rect 1468 2314 1542 2370
rect 1598 2314 1684 2370
rect 1740 2314 1808 2370
rect 1468 2228 1808 2314
rect 1468 2172 1542 2228
rect 1598 2172 1684 2228
rect 1740 2172 1808 2228
rect 1468 2086 1808 2172
rect 1468 2030 1542 2086
rect 1598 2030 1684 2086
rect 1740 2030 1808 2086
rect 1468 1944 1808 2030
rect 1468 1888 1542 1944
rect 1598 1888 1684 1944
rect 1740 1888 1808 1944
rect 1468 1802 1808 1888
rect 1468 1746 1542 1802
rect 1598 1746 1684 1802
rect 1740 1746 1808 1802
rect 1468 1660 1808 1746
rect 1468 1604 1542 1660
rect 1598 1604 1684 1660
rect 1740 1604 1808 1660
rect 1468 1518 1808 1604
rect 1468 1462 1542 1518
rect 1598 1462 1684 1518
rect 1740 1462 1808 1518
rect 1468 1376 1808 1462
rect 1468 1320 1542 1376
rect 1598 1320 1684 1376
rect 1740 1320 1808 1376
rect 1468 1234 1808 1320
rect 1468 1178 1542 1234
rect 1598 1178 1684 1234
rect 1740 1178 1808 1234
rect 1468 1092 1808 1178
rect 1468 1036 1542 1092
rect 1598 1036 1684 1092
rect 1740 1036 1808 1092
rect 1468 950 1808 1036
rect 1468 894 1542 950
rect 1598 894 1684 950
rect 1740 894 1808 950
rect 1468 808 1808 894
rect 1468 752 1542 808
rect 1598 752 1684 808
rect 1740 752 1808 808
rect 1468 666 1808 752
rect 1468 610 1542 666
rect 1598 610 1684 666
rect 1740 610 1808 666
rect 1468 524 1808 610
rect 1468 468 1542 524
rect 1598 468 1684 524
rect 1740 468 1808 524
rect 1468 400 1808 468
rect 1868 12310 2208 12400
rect 1868 12254 1939 12310
rect 1995 12254 2081 12310
rect 2137 12254 2208 12310
rect 1868 12168 2208 12254
rect 1868 12112 1939 12168
rect 1995 12112 2081 12168
rect 2137 12112 2208 12168
rect 1868 12026 2208 12112
rect 1868 11970 1939 12026
rect 1995 11970 2081 12026
rect 2137 11970 2208 12026
rect 1868 11884 2208 11970
rect 1868 11828 1939 11884
rect 1995 11828 2081 11884
rect 2137 11828 2208 11884
rect 1868 11742 2208 11828
rect 1868 11686 1939 11742
rect 1995 11686 2081 11742
rect 2137 11686 2208 11742
rect 1868 11600 2208 11686
rect 1868 11544 1939 11600
rect 1995 11544 2081 11600
rect 2137 11544 2208 11600
rect 1868 11458 2208 11544
rect 1868 11402 1939 11458
rect 1995 11402 2081 11458
rect 2137 11402 2208 11458
rect 1868 11316 2208 11402
rect 1868 11260 1939 11316
rect 1995 11260 2081 11316
rect 2137 11260 2208 11316
rect 1868 11174 2208 11260
rect 1868 11118 1939 11174
rect 1995 11118 2081 11174
rect 2137 11118 2208 11174
rect 1868 11032 2208 11118
rect 1868 10976 1939 11032
rect 1995 10976 2081 11032
rect 2137 10976 2208 11032
rect 1868 10890 2208 10976
rect 1868 10834 1939 10890
rect 1995 10834 2081 10890
rect 2137 10834 2208 10890
rect 1868 10748 2208 10834
rect 1868 10692 1939 10748
rect 1995 10692 2081 10748
rect 2137 10692 2208 10748
rect 1868 10606 2208 10692
rect 1868 10550 1939 10606
rect 1995 10550 2081 10606
rect 2137 10550 2208 10606
rect 1868 10464 2208 10550
rect 1868 10408 1939 10464
rect 1995 10408 2081 10464
rect 2137 10408 2208 10464
rect 1868 10322 2208 10408
rect 1868 10266 1939 10322
rect 1995 10266 2081 10322
rect 2137 10266 2208 10322
rect 1868 10180 2208 10266
rect 1868 10124 1939 10180
rect 1995 10124 2081 10180
rect 2137 10124 2208 10180
rect 1868 10038 2208 10124
rect 1868 9982 1939 10038
rect 1995 9982 2081 10038
rect 2137 9982 2208 10038
rect 1868 9896 2208 9982
rect 1868 9840 1939 9896
rect 1995 9840 2081 9896
rect 2137 9840 2208 9896
rect 1868 9754 2208 9840
rect 1868 9698 1939 9754
rect 1995 9698 2081 9754
rect 2137 9698 2208 9754
rect 1868 9612 2208 9698
rect 1868 9556 1939 9612
rect 1995 9556 2081 9612
rect 2137 9556 2208 9612
rect 1868 9470 2208 9556
rect 1868 9414 1939 9470
rect 1995 9414 2081 9470
rect 2137 9414 2208 9470
rect 1868 9328 2208 9414
rect 1868 9272 1939 9328
rect 1995 9272 2081 9328
rect 2137 9272 2208 9328
rect 1868 9186 2208 9272
rect 1868 9130 1939 9186
rect 1995 9130 2081 9186
rect 2137 9130 2208 9186
rect 1868 9044 2208 9130
rect 1868 8988 1939 9044
rect 1995 8988 2081 9044
rect 2137 8988 2208 9044
rect 1868 8902 2208 8988
rect 1868 8846 1939 8902
rect 1995 8846 2081 8902
rect 2137 8846 2208 8902
rect 1868 8760 2208 8846
rect 1868 8704 1939 8760
rect 1995 8704 2081 8760
rect 2137 8704 2208 8760
rect 1868 8618 2208 8704
rect 1868 8562 1939 8618
rect 1995 8562 2081 8618
rect 2137 8562 2208 8618
rect 1868 8476 2208 8562
rect 1868 8420 1939 8476
rect 1995 8420 2081 8476
rect 2137 8420 2208 8476
rect 1868 8334 2208 8420
rect 1868 8278 1939 8334
rect 1995 8278 2081 8334
rect 2137 8278 2208 8334
rect 1868 8192 2208 8278
rect 1868 8136 1939 8192
rect 1995 8136 2081 8192
rect 2137 8136 2208 8192
rect 1868 8050 2208 8136
rect 1868 7994 1939 8050
rect 1995 7994 2081 8050
rect 2137 7994 2208 8050
rect 1868 7908 2208 7994
rect 1868 7852 1939 7908
rect 1995 7852 2081 7908
rect 2137 7852 2208 7908
rect 1868 7766 2208 7852
rect 1868 7710 1939 7766
rect 1995 7710 2081 7766
rect 2137 7710 2208 7766
rect 1868 7624 2208 7710
rect 1868 7568 1939 7624
rect 1995 7568 2081 7624
rect 2137 7568 2208 7624
rect 1868 7482 2208 7568
rect 1868 7426 1939 7482
rect 1995 7426 2081 7482
rect 2137 7426 2208 7482
rect 1868 7340 2208 7426
rect 1868 7284 1939 7340
rect 1995 7284 2081 7340
rect 2137 7284 2208 7340
rect 1868 7198 2208 7284
rect 1868 7142 1939 7198
rect 1995 7142 2081 7198
rect 2137 7142 2208 7198
rect 1868 7056 2208 7142
rect 1868 7000 1939 7056
rect 1995 7000 2081 7056
rect 2137 7000 2208 7056
rect 1868 6914 2208 7000
rect 1868 6858 1939 6914
rect 1995 6858 2081 6914
rect 2137 6858 2208 6914
rect 1868 6772 2208 6858
rect 1868 6716 1939 6772
rect 1995 6716 2081 6772
rect 2137 6716 2208 6772
rect 1868 6630 2208 6716
rect 1868 6574 1939 6630
rect 1995 6574 2081 6630
rect 2137 6574 2208 6630
rect 1868 6488 2208 6574
rect 1868 6432 1939 6488
rect 1995 6432 2081 6488
rect 2137 6432 2208 6488
rect 1868 6346 2208 6432
rect 1868 6290 1939 6346
rect 1995 6290 2081 6346
rect 2137 6290 2208 6346
rect 1868 6204 2208 6290
rect 1868 6148 1939 6204
rect 1995 6148 2081 6204
rect 2137 6148 2208 6204
rect 1868 6062 2208 6148
rect 1868 6006 1939 6062
rect 1995 6006 2081 6062
rect 2137 6006 2208 6062
rect 1868 5920 2208 6006
rect 1868 5864 1939 5920
rect 1995 5864 2081 5920
rect 2137 5864 2208 5920
rect 1868 5778 2208 5864
rect 1868 5722 1939 5778
rect 1995 5722 2081 5778
rect 2137 5722 2208 5778
rect 1868 5636 2208 5722
rect 1868 5580 1939 5636
rect 1995 5580 2081 5636
rect 2137 5580 2208 5636
rect 1868 5494 2208 5580
rect 1868 5438 1939 5494
rect 1995 5438 2081 5494
rect 2137 5438 2208 5494
rect 1868 5352 2208 5438
rect 1868 5296 1939 5352
rect 1995 5296 2081 5352
rect 2137 5296 2208 5352
rect 1868 5210 2208 5296
rect 1868 5154 1939 5210
rect 1995 5154 2081 5210
rect 2137 5154 2208 5210
rect 1868 5068 2208 5154
rect 1868 5012 1939 5068
rect 1995 5012 2081 5068
rect 2137 5012 2208 5068
rect 1868 4926 2208 5012
rect 1868 4870 1939 4926
rect 1995 4870 2081 4926
rect 2137 4870 2208 4926
rect 1868 4784 2208 4870
rect 1868 4728 1939 4784
rect 1995 4728 2081 4784
rect 2137 4728 2208 4784
rect 1868 4642 2208 4728
rect 1868 4586 1939 4642
rect 1995 4586 2081 4642
rect 2137 4586 2208 4642
rect 1868 4500 2208 4586
rect 1868 4444 1939 4500
rect 1995 4444 2081 4500
rect 2137 4444 2208 4500
rect 1868 4358 2208 4444
rect 1868 4302 1939 4358
rect 1995 4302 2081 4358
rect 2137 4302 2208 4358
rect 1868 4216 2208 4302
rect 1868 4160 1939 4216
rect 1995 4160 2081 4216
rect 2137 4160 2208 4216
rect 1868 4074 2208 4160
rect 1868 4018 1939 4074
rect 1995 4018 2081 4074
rect 2137 4018 2208 4074
rect 1868 3932 2208 4018
rect 1868 3876 1939 3932
rect 1995 3876 2081 3932
rect 2137 3876 2208 3932
rect 1868 3790 2208 3876
rect 1868 3734 1939 3790
rect 1995 3734 2081 3790
rect 2137 3734 2208 3790
rect 1868 3648 2208 3734
rect 1868 3592 1939 3648
rect 1995 3592 2081 3648
rect 2137 3592 2208 3648
rect 1868 3506 2208 3592
rect 1868 3450 1939 3506
rect 1995 3450 2081 3506
rect 2137 3450 2208 3506
rect 1868 3364 2208 3450
rect 1868 3308 1939 3364
rect 1995 3308 2081 3364
rect 2137 3308 2208 3364
rect 1868 3222 2208 3308
rect 1868 3166 1939 3222
rect 1995 3166 2081 3222
rect 2137 3166 2208 3222
rect 1868 3080 2208 3166
rect 1868 3024 1939 3080
rect 1995 3024 2081 3080
rect 2137 3024 2208 3080
rect 1868 2938 2208 3024
rect 1868 2882 1939 2938
rect 1995 2882 2081 2938
rect 2137 2882 2208 2938
rect 1868 2796 2208 2882
rect 1868 2740 1939 2796
rect 1995 2740 2081 2796
rect 2137 2740 2208 2796
rect 1868 2654 2208 2740
rect 1868 2598 1939 2654
rect 1995 2598 2081 2654
rect 2137 2598 2208 2654
rect 1868 2512 2208 2598
rect 1868 2456 1939 2512
rect 1995 2456 2081 2512
rect 2137 2456 2208 2512
rect 1868 2370 2208 2456
rect 1868 2314 1939 2370
rect 1995 2314 2081 2370
rect 2137 2314 2208 2370
rect 1868 2228 2208 2314
rect 1868 2172 1939 2228
rect 1995 2172 2081 2228
rect 2137 2172 2208 2228
rect 1868 2086 2208 2172
rect 1868 2030 1939 2086
rect 1995 2030 2081 2086
rect 2137 2030 2208 2086
rect 1868 1944 2208 2030
rect 1868 1888 1939 1944
rect 1995 1888 2081 1944
rect 2137 1888 2208 1944
rect 1868 1802 2208 1888
rect 1868 1746 1939 1802
rect 1995 1746 2081 1802
rect 2137 1746 2208 1802
rect 1868 1660 2208 1746
rect 1868 1604 1939 1660
rect 1995 1604 2081 1660
rect 2137 1604 2208 1660
rect 1868 1518 2208 1604
rect 1868 1462 1939 1518
rect 1995 1462 2081 1518
rect 2137 1462 2208 1518
rect 1868 1376 2208 1462
rect 1868 1320 1939 1376
rect 1995 1320 2081 1376
rect 2137 1320 2208 1376
rect 1868 1234 2208 1320
rect 1868 1178 1939 1234
rect 1995 1178 2081 1234
rect 2137 1178 2208 1234
rect 1868 1092 2208 1178
rect 1868 1036 1939 1092
rect 1995 1036 2081 1092
rect 2137 1036 2208 1092
rect 1868 950 2208 1036
rect 1868 894 1939 950
rect 1995 894 2081 950
rect 2137 894 2208 950
rect 1868 808 2208 894
rect 1868 752 1939 808
rect 1995 752 2081 808
rect 2137 752 2208 808
rect 1868 666 2208 752
rect 1868 610 1939 666
rect 1995 610 2081 666
rect 2137 610 2208 666
rect 1868 524 2208 610
rect 1868 468 1939 524
rect 1995 468 2081 524
rect 2137 468 2208 524
rect 1868 400 2208 468
rect 2268 12310 2608 12400
rect 2268 12254 2336 12310
rect 2392 12254 2478 12310
rect 2534 12254 2608 12310
rect 2268 12168 2608 12254
rect 2268 12112 2336 12168
rect 2392 12112 2478 12168
rect 2534 12112 2608 12168
rect 2268 12026 2608 12112
rect 2268 11970 2336 12026
rect 2392 11970 2478 12026
rect 2534 11970 2608 12026
rect 2268 11884 2608 11970
rect 2268 11828 2336 11884
rect 2392 11828 2478 11884
rect 2534 11828 2608 11884
rect 2268 11742 2608 11828
rect 2268 11686 2336 11742
rect 2392 11686 2478 11742
rect 2534 11686 2608 11742
rect 2268 11600 2608 11686
rect 2268 11544 2336 11600
rect 2392 11544 2478 11600
rect 2534 11544 2608 11600
rect 2268 11458 2608 11544
rect 2268 11402 2336 11458
rect 2392 11402 2478 11458
rect 2534 11402 2608 11458
rect 2268 11316 2608 11402
rect 2268 11260 2336 11316
rect 2392 11260 2478 11316
rect 2534 11260 2608 11316
rect 2268 11174 2608 11260
rect 2268 11118 2336 11174
rect 2392 11118 2478 11174
rect 2534 11118 2608 11174
rect 2268 11032 2608 11118
rect 2268 10976 2336 11032
rect 2392 10976 2478 11032
rect 2534 10976 2608 11032
rect 2268 10890 2608 10976
rect 2268 10834 2336 10890
rect 2392 10834 2478 10890
rect 2534 10834 2608 10890
rect 2268 10748 2608 10834
rect 2268 10692 2336 10748
rect 2392 10692 2478 10748
rect 2534 10692 2608 10748
rect 2268 10606 2608 10692
rect 2268 10550 2336 10606
rect 2392 10550 2478 10606
rect 2534 10550 2608 10606
rect 2268 10464 2608 10550
rect 2268 10408 2336 10464
rect 2392 10408 2478 10464
rect 2534 10408 2608 10464
rect 2268 10322 2608 10408
rect 2268 10266 2336 10322
rect 2392 10266 2478 10322
rect 2534 10266 2608 10322
rect 2268 10180 2608 10266
rect 2268 10124 2336 10180
rect 2392 10124 2478 10180
rect 2534 10124 2608 10180
rect 2268 10038 2608 10124
rect 2268 9982 2336 10038
rect 2392 9982 2478 10038
rect 2534 9982 2608 10038
rect 2268 9896 2608 9982
rect 2268 9840 2336 9896
rect 2392 9840 2478 9896
rect 2534 9840 2608 9896
rect 2268 9754 2608 9840
rect 2268 9698 2336 9754
rect 2392 9698 2478 9754
rect 2534 9698 2608 9754
rect 2268 9612 2608 9698
rect 2268 9556 2336 9612
rect 2392 9556 2478 9612
rect 2534 9556 2608 9612
rect 2268 9470 2608 9556
rect 2268 9414 2336 9470
rect 2392 9414 2478 9470
rect 2534 9414 2608 9470
rect 2268 9328 2608 9414
rect 2268 9272 2336 9328
rect 2392 9272 2478 9328
rect 2534 9272 2608 9328
rect 2268 9186 2608 9272
rect 2268 9130 2336 9186
rect 2392 9130 2478 9186
rect 2534 9130 2608 9186
rect 2268 9044 2608 9130
rect 2268 8988 2336 9044
rect 2392 8988 2478 9044
rect 2534 8988 2608 9044
rect 2268 8902 2608 8988
rect 2268 8846 2336 8902
rect 2392 8846 2478 8902
rect 2534 8846 2608 8902
rect 2268 8760 2608 8846
rect 2268 8704 2336 8760
rect 2392 8704 2478 8760
rect 2534 8704 2608 8760
rect 2268 8618 2608 8704
rect 2268 8562 2336 8618
rect 2392 8562 2478 8618
rect 2534 8562 2608 8618
rect 2268 8476 2608 8562
rect 2268 8420 2336 8476
rect 2392 8420 2478 8476
rect 2534 8420 2608 8476
rect 2268 8334 2608 8420
rect 2268 8278 2336 8334
rect 2392 8278 2478 8334
rect 2534 8278 2608 8334
rect 2268 8192 2608 8278
rect 2268 8136 2336 8192
rect 2392 8136 2478 8192
rect 2534 8136 2608 8192
rect 2268 8050 2608 8136
rect 2268 7994 2336 8050
rect 2392 7994 2478 8050
rect 2534 7994 2608 8050
rect 2268 7908 2608 7994
rect 2268 7852 2336 7908
rect 2392 7852 2478 7908
rect 2534 7852 2608 7908
rect 2268 7766 2608 7852
rect 2268 7710 2336 7766
rect 2392 7710 2478 7766
rect 2534 7710 2608 7766
rect 2268 7624 2608 7710
rect 2268 7568 2336 7624
rect 2392 7568 2478 7624
rect 2534 7568 2608 7624
rect 2268 7482 2608 7568
rect 2268 7426 2336 7482
rect 2392 7426 2478 7482
rect 2534 7426 2608 7482
rect 2268 7340 2608 7426
rect 2268 7284 2336 7340
rect 2392 7284 2478 7340
rect 2534 7284 2608 7340
rect 2268 7198 2608 7284
rect 2268 7142 2336 7198
rect 2392 7142 2478 7198
rect 2534 7142 2608 7198
rect 2268 7056 2608 7142
rect 2268 7000 2336 7056
rect 2392 7000 2478 7056
rect 2534 7000 2608 7056
rect 2268 6914 2608 7000
rect 2268 6858 2336 6914
rect 2392 6858 2478 6914
rect 2534 6858 2608 6914
rect 2268 6772 2608 6858
rect 2268 6716 2336 6772
rect 2392 6716 2478 6772
rect 2534 6716 2608 6772
rect 2268 6630 2608 6716
rect 2268 6574 2336 6630
rect 2392 6574 2478 6630
rect 2534 6574 2608 6630
rect 2268 6488 2608 6574
rect 2268 6432 2336 6488
rect 2392 6432 2478 6488
rect 2534 6432 2608 6488
rect 2268 6346 2608 6432
rect 2268 6290 2336 6346
rect 2392 6290 2478 6346
rect 2534 6290 2608 6346
rect 2268 6204 2608 6290
rect 2268 6148 2336 6204
rect 2392 6148 2478 6204
rect 2534 6148 2608 6204
rect 2268 6062 2608 6148
rect 2268 6006 2336 6062
rect 2392 6006 2478 6062
rect 2534 6006 2608 6062
rect 2268 5920 2608 6006
rect 2268 5864 2336 5920
rect 2392 5864 2478 5920
rect 2534 5864 2608 5920
rect 2268 5778 2608 5864
rect 2268 5722 2336 5778
rect 2392 5722 2478 5778
rect 2534 5722 2608 5778
rect 2268 5636 2608 5722
rect 2268 5580 2336 5636
rect 2392 5580 2478 5636
rect 2534 5580 2608 5636
rect 2268 5494 2608 5580
rect 2268 5438 2336 5494
rect 2392 5438 2478 5494
rect 2534 5438 2608 5494
rect 2268 5352 2608 5438
rect 2268 5296 2336 5352
rect 2392 5296 2478 5352
rect 2534 5296 2608 5352
rect 2268 5210 2608 5296
rect 2268 5154 2336 5210
rect 2392 5154 2478 5210
rect 2534 5154 2608 5210
rect 2268 5068 2608 5154
rect 2268 5012 2336 5068
rect 2392 5012 2478 5068
rect 2534 5012 2608 5068
rect 2268 4926 2608 5012
rect 2268 4870 2336 4926
rect 2392 4870 2478 4926
rect 2534 4870 2608 4926
rect 2268 4784 2608 4870
rect 2268 4728 2336 4784
rect 2392 4728 2478 4784
rect 2534 4728 2608 4784
rect 2268 4642 2608 4728
rect 2268 4586 2336 4642
rect 2392 4586 2478 4642
rect 2534 4586 2608 4642
rect 2268 4500 2608 4586
rect 2268 4444 2336 4500
rect 2392 4444 2478 4500
rect 2534 4444 2608 4500
rect 2268 4358 2608 4444
rect 2268 4302 2336 4358
rect 2392 4302 2478 4358
rect 2534 4302 2608 4358
rect 2268 4216 2608 4302
rect 2268 4160 2336 4216
rect 2392 4160 2478 4216
rect 2534 4160 2608 4216
rect 2268 4074 2608 4160
rect 2268 4018 2336 4074
rect 2392 4018 2478 4074
rect 2534 4018 2608 4074
rect 2268 3932 2608 4018
rect 2268 3876 2336 3932
rect 2392 3876 2478 3932
rect 2534 3876 2608 3932
rect 2268 3790 2608 3876
rect 2268 3734 2336 3790
rect 2392 3734 2478 3790
rect 2534 3734 2608 3790
rect 2268 3648 2608 3734
rect 2268 3592 2336 3648
rect 2392 3592 2478 3648
rect 2534 3592 2608 3648
rect 2268 3506 2608 3592
rect 2268 3450 2336 3506
rect 2392 3450 2478 3506
rect 2534 3450 2608 3506
rect 2268 3364 2608 3450
rect 2268 3308 2336 3364
rect 2392 3308 2478 3364
rect 2534 3308 2608 3364
rect 2268 3222 2608 3308
rect 2268 3166 2336 3222
rect 2392 3166 2478 3222
rect 2534 3166 2608 3222
rect 2268 3080 2608 3166
rect 2268 3024 2336 3080
rect 2392 3024 2478 3080
rect 2534 3024 2608 3080
rect 2268 2938 2608 3024
rect 2268 2882 2336 2938
rect 2392 2882 2478 2938
rect 2534 2882 2608 2938
rect 2268 2796 2608 2882
rect 2268 2740 2336 2796
rect 2392 2740 2478 2796
rect 2534 2740 2608 2796
rect 2268 2654 2608 2740
rect 2268 2598 2336 2654
rect 2392 2598 2478 2654
rect 2534 2598 2608 2654
rect 2268 2512 2608 2598
rect 2268 2456 2336 2512
rect 2392 2456 2478 2512
rect 2534 2456 2608 2512
rect 2268 2370 2608 2456
rect 2268 2314 2336 2370
rect 2392 2314 2478 2370
rect 2534 2314 2608 2370
rect 2268 2228 2608 2314
rect 2268 2172 2336 2228
rect 2392 2172 2478 2228
rect 2534 2172 2608 2228
rect 2268 2086 2608 2172
rect 2268 2030 2336 2086
rect 2392 2030 2478 2086
rect 2534 2030 2608 2086
rect 2268 1944 2608 2030
rect 2268 1888 2336 1944
rect 2392 1888 2478 1944
rect 2534 1888 2608 1944
rect 2268 1802 2608 1888
rect 2268 1746 2336 1802
rect 2392 1746 2478 1802
rect 2534 1746 2608 1802
rect 2268 1660 2608 1746
rect 2268 1604 2336 1660
rect 2392 1604 2478 1660
rect 2534 1604 2608 1660
rect 2268 1518 2608 1604
rect 2268 1462 2336 1518
rect 2392 1462 2478 1518
rect 2534 1462 2608 1518
rect 2268 1376 2608 1462
rect 2268 1320 2336 1376
rect 2392 1320 2478 1376
rect 2534 1320 2608 1376
rect 2268 1234 2608 1320
rect 2268 1178 2336 1234
rect 2392 1178 2478 1234
rect 2534 1178 2608 1234
rect 2268 1092 2608 1178
rect 2268 1036 2336 1092
rect 2392 1036 2478 1092
rect 2534 1036 2608 1092
rect 2268 950 2608 1036
rect 2268 894 2336 950
rect 2392 894 2478 950
rect 2534 894 2608 950
rect 2268 808 2608 894
rect 2268 752 2336 808
rect 2392 752 2478 808
rect 2534 752 2608 808
rect 2268 666 2608 752
rect 2268 610 2336 666
rect 2392 610 2478 666
rect 2534 610 2608 666
rect 2268 524 2608 610
rect 2268 468 2336 524
rect 2392 468 2478 524
rect 2534 468 2608 524
rect 2268 400 2608 468
rect 2668 12310 3008 12400
rect 2668 12254 2740 12310
rect 2796 12254 2882 12310
rect 2938 12254 3008 12310
rect 2668 12168 3008 12254
rect 2668 12112 2740 12168
rect 2796 12112 2882 12168
rect 2938 12112 3008 12168
rect 2668 12026 3008 12112
rect 2668 11970 2740 12026
rect 2796 11970 2882 12026
rect 2938 11970 3008 12026
rect 2668 11884 3008 11970
rect 2668 11828 2740 11884
rect 2796 11828 2882 11884
rect 2938 11828 3008 11884
rect 2668 11742 3008 11828
rect 2668 11686 2740 11742
rect 2796 11686 2882 11742
rect 2938 11686 3008 11742
rect 2668 11600 3008 11686
rect 2668 11544 2740 11600
rect 2796 11544 2882 11600
rect 2938 11544 3008 11600
rect 2668 11458 3008 11544
rect 2668 11402 2740 11458
rect 2796 11402 2882 11458
rect 2938 11402 3008 11458
rect 2668 11316 3008 11402
rect 2668 11260 2740 11316
rect 2796 11260 2882 11316
rect 2938 11260 3008 11316
rect 2668 11174 3008 11260
rect 2668 11118 2740 11174
rect 2796 11118 2882 11174
rect 2938 11118 3008 11174
rect 2668 11032 3008 11118
rect 2668 10976 2740 11032
rect 2796 10976 2882 11032
rect 2938 10976 3008 11032
rect 2668 10890 3008 10976
rect 2668 10834 2740 10890
rect 2796 10834 2882 10890
rect 2938 10834 3008 10890
rect 2668 10748 3008 10834
rect 2668 10692 2740 10748
rect 2796 10692 2882 10748
rect 2938 10692 3008 10748
rect 2668 10606 3008 10692
rect 2668 10550 2740 10606
rect 2796 10550 2882 10606
rect 2938 10550 3008 10606
rect 2668 10464 3008 10550
rect 2668 10408 2740 10464
rect 2796 10408 2882 10464
rect 2938 10408 3008 10464
rect 2668 10322 3008 10408
rect 2668 10266 2740 10322
rect 2796 10266 2882 10322
rect 2938 10266 3008 10322
rect 2668 10180 3008 10266
rect 2668 10124 2740 10180
rect 2796 10124 2882 10180
rect 2938 10124 3008 10180
rect 2668 10038 3008 10124
rect 2668 9982 2740 10038
rect 2796 9982 2882 10038
rect 2938 9982 3008 10038
rect 2668 9896 3008 9982
rect 2668 9840 2740 9896
rect 2796 9840 2882 9896
rect 2938 9840 3008 9896
rect 2668 9754 3008 9840
rect 2668 9698 2740 9754
rect 2796 9698 2882 9754
rect 2938 9698 3008 9754
rect 2668 9612 3008 9698
rect 2668 9556 2740 9612
rect 2796 9556 2882 9612
rect 2938 9556 3008 9612
rect 2668 9470 3008 9556
rect 2668 9414 2740 9470
rect 2796 9414 2882 9470
rect 2938 9414 3008 9470
rect 2668 9328 3008 9414
rect 2668 9272 2740 9328
rect 2796 9272 2882 9328
rect 2938 9272 3008 9328
rect 2668 9186 3008 9272
rect 2668 9130 2740 9186
rect 2796 9130 2882 9186
rect 2938 9130 3008 9186
rect 2668 9044 3008 9130
rect 2668 8988 2740 9044
rect 2796 8988 2882 9044
rect 2938 8988 3008 9044
rect 2668 8902 3008 8988
rect 2668 8846 2740 8902
rect 2796 8846 2882 8902
rect 2938 8846 3008 8902
rect 2668 8760 3008 8846
rect 2668 8704 2740 8760
rect 2796 8704 2882 8760
rect 2938 8704 3008 8760
rect 2668 8618 3008 8704
rect 2668 8562 2740 8618
rect 2796 8562 2882 8618
rect 2938 8562 3008 8618
rect 2668 8476 3008 8562
rect 2668 8420 2740 8476
rect 2796 8420 2882 8476
rect 2938 8420 3008 8476
rect 2668 8334 3008 8420
rect 2668 8278 2740 8334
rect 2796 8278 2882 8334
rect 2938 8278 3008 8334
rect 2668 8192 3008 8278
rect 2668 8136 2740 8192
rect 2796 8136 2882 8192
rect 2938 8136 3008 8192
rect 2668 8050 3008 8136
rect 2668 7994 2740 8050
rect 2796 7994 2882 8050
rect 2938 7994 3008 8050
rect 2668 7908 3008 7994
rect 2668 7852 2740 7908
rect 2796 7852 2882 7908
rect 2938 7852 3008 7908
rect 2668 7766 3008 7852
rect 2668 7710 2740 7766
rect 2796 7710 2882 7766
rect 2938 7710 3008 7766
rect 2668 7624 3008 7710
rect 2668 7568 2740 7624
rect 2796 7568 2882 7624
rect 2938 7568 3008 7624
rect 2668 7482 3008 7568
rect 2668 7426 2740 7482
rect 2796 7426 2882 7482
rect 2938 7426 3008 7482
rect 2668 7340 3008 7426
rect 2668 7284 2740 7340
rect 2796 7284 2882 7340
rect 2938 7284 3008 7340
rect 2668 7198 3008 7284
rect 2668 7142 2740 7198
rect 2796 7142 2882 7198
rect 2938 7142 3008 7198
rect 2668 7056 3008 7142
rect 2668 7000 2740 7056
rect 2796 7000 2882 7056
rect 2938 7000 3008 7056
rect 2668 6914 3008 7000
rect 2668 6858 2740 6914
rect 2796 6858 2882 6914
rect 2938 6858 3008 6914
rect 2668 6772 3008 6858
rect 2668 6716 2740 6772
rect 2796 6716 2882 6772
rect 2938 6716 3008 6772
rect 2668 6630 3008 6716
rect 2668 6574 2740 6630
rect 2796 6574 2882 6630
rect 2938 6574 3008 6630
rect 2668 6488 3008 6574
rect 2668 6432 2740 6488
rect 2796 6432 2882 6488
rect 2938 6432 3008 6488
rect 2668 6346 3008 6432
rect 2668 6290 2740 6346
rect 2796 6290 2882 6346
rect 2938 6290 3008 6346
rect 2668 6204 3008 6290
rect 2668 6148 2740 6204
rect 2796 6148 2882 6204
rect 2938 6148 3008 6204
rect 2668 6062 3008 6148
rect 2668 6006 2740 6062
rect 2796 6006 2882 6062
rect 2938 6006 3008 6062
rect 2668 5920 3008 6006
rect 2668 5864 2740 5920
rect 2796 5864 2882 5920
rect 2938 5864 3008 5920
rect 2668 5778 3008 5864
rect 2668 5722 2740 5778
rect 2796 5722 2882 5778
rect 2938 5722 3008 5778
rect 2668 5636 3008 5722
rect 2668 5580 2740 5636
rect 2796 5580 2882 5636
rect 2938 5580 3008 5636
rect 2668 5494 3008 5580
rect 2668 5438 2740 5494
rect 2796 5438 2882 5494
rect 2938 5438 3008 5494
rect 2668 5352 3008 5438
rect 2668 5296 2740 5352
rect 2796 5296 2882 5352
rect 2938 5296 3008 5352
rect 2668 5210 3008 5296
rect 2668 5154 2740 5210
rect 2796 5154 2882 5210
rect 2938 5154 3008 5210
rect 2668 5068 3008 5154
rect 2668 5012 2740 5068
rect 2796 5012 2882 5068
rect 2938 5012 3008 5068
rect 2668 4926 3008 5012
rect 2668 4870 2740 4926
rect 2796 4870 2882 4926
rect 2938 4870 3008 4926
rect 2668 4784 3008 4870
rect 2668 4728 2740 4784
rect 2796 4728 2882 4784
rect 2938 4728 3008 4784
rect 2668 4642 3008 4728
rect 2668 4586 2740 4642
rect 2796 4586 2882 4642
rect 2938 4586 3008 4642
rect 2668 4500 3008 4586
rect 2668 4444 2740 4500
rect 2796 4444 2882 4500
rect 2938 4444 3008 4500
rect 2668 4358 3008 4444
rect 2668 4302 2740 4358
rect 2796 4302 2882 4358
rect 2938 4302 3008 4358
rect 2668 4216 3008 4302
rect 2668 4160 2740 4216
rect 2796 4160 2882 4216
rect 2938 4160 3008 4216
rect 2668 4074 3008 4160
rect 2668 4018 2740 4074
rect 2796 4018 2882 4074
rect 2938 4018 3008 4074
rect 2668 3932 3008 4018
rect 2668 3876 2740 3932
rect 2796 3876 2882 3932
rect 2938 3876 3008 3932
rect 2668 3790 3008 3876
rect 2668 3734 2740 3790
rect 2796 3734 2882 3790
rect 2938 3734 3008 3790
rect 2668 3648 3008 3734
rect 2668 3592 2740 3648
rect 2796 3592 2882 3648
rect 2938 3592 3008 3648
rect 2668 3506 3008 3592
rect 2668 3450 2740 3506
rect 2796 3450 2882 3506
rect 2938 3450 3008 3506
rect 2668 3364 3008 3450
rect 2668 3308 2740 3364
rect 2796 3308 2882 3364
rect 2938 3308 3008 3364
rect 2668 3222 3008 3308
rect 2668 3166 2740 3222
rect 2796 3166 2882 3222
rect 2938 3166 3008 3222
rect 2668 3080 3008 3166
rect 2668 3024 2740 3080
rect 2796 3024 2882 3080
rect 2938 3024 3008 3080
rect 2668 2938 3008 3024
rect 2668 2882 2740 2938
rect 2796 2882 2882 2938
rect 2938 2882 3008 2938
rect 2668 2796 3008 2882
rect 2668 2740 2740 2796
rect 2796 2740 2882 2796
rect 2938 2740 3008 2796
rect 2668 2654 3008 2740
rect 2668 2598 2740 2654
rect 2796 2598 2882 2654
rect 2938 2598 3008 2654
rect 2668 2512 3008 2598
rect 2668 2456 2740 2512
rect 2796 2456 2882 2512
rect 2938 2456 3008 2512
rect 2668 2370 3008 2456
rect 2668 2314 2740 2370
rect 2796 2314 2882 2370
rect 2938 2314 3008 2370
rect 2668 2228 3008 2314
rect 2668 2172 2740 2228
rect 2796 2172 2882 2228
rect 2938 2172 3008 2228
rect 2668 2086 3008 2172
rect 2668 2030 2740 2086
rect 2796 2030 2882 2086
rect 2938 2030 3008 2086
rect 2668 1944 3008 2030
rect 2668 1888 2740 1944
rect 2796 1888 2882 1944
rect 2938 1888 3008 1944
rect 2668 1802 3008 1888
rect 2668 1746 2740 1802
rect 2796 1746 2882 1802
rect 2938 1746 3008 1802
rect 2668 1660 3008 1746
rect 2668 1604 2740 1660
rect 2796 1604 2882 1660
rect 2938 1604 3008 1660
rect 2668 1518 3008 1604
rect 2668 1462 2740 1518
rect 2796 1462 2882 1518
rect 2938 1462 3008 1518
rect 2668 1376 3008 1462
rect 2668 1320 2740 1376
rect 2796 1320 2882 1376
rect 2938 1320 3008 1376
rect 2668 1234 3008 1320
rect 2668 1178 2740 1234
rect 2796 1178 2882 1234
rect 2938 1178 3008 1234
rect 2668 1092 3008 1178
rect 2668 1036 2740 1092
rect 2796 1036 2882 1092
rect 2938 1036 3008 1092
rect 2668 950 3008 1036
rect 2668 894 2740 950
rect 2796 894 2882 950
rect 2938 894 3008 950
rect 2668 808 3008 894
rect 2668 752 2740 808
rect 2796 752 2882 808
rect 2938 752 3008 808
rect 2668 666 3008 752
rect 2668 610 2740 666
rect 2796 610 2882 666
rect 2938 610 3008 666
rect 2668 524 3008 610
rect 2668 468 2740 524
rect 2796 468 2882 524
rect 2938 468 3008 524
rect 2668 400 3008 468
rect 3068 12310 3408 12400
rect 3068 12254 3136 12310
rect 3192 12254 3278 12310
rect 3334 12254 3408 12310
rect 3068 12168 3408 12254
rect 3068 12112 3136 12168
rect 3192 12112 3278 12168
rect 3334 12112 3408 12168
rect 3068 12026 3408 12112
rect 3068 11970 3136 12026
rect 3192 11970 3278 12026
rect 3334 11970 3408 12026
rect 3068 11884 3408 11970
rect 3068 11828 3136 11884
rect 3192 11828 3278 11884
rect 3334 11828 3408 11884
rect 3068 11742 3408 11828
rect 3068 11686 3136 11742
rect 3192 11686 3278 11742
rect 3334 11686 3408 11742
rect 3068 11600 3408 11686
rect 3068 11544 3136 11600
rect 3192 11544 3278 11600
rect 3334 11544 3408 11600
rect 3068 11458 3408 11544
rect 3068 11402 3136 11458
rect 3192 11402 3278 11458
rect 3334 11402 3408 11458
rect 3068 11316 3408 11402
rect 3068 11260 3136 11316
rect 3192 11260 3278 11316
rect 3334 11260 3408 11316
rect 3068 11174 3408 11260
rect 3068 11118 3136 11174
rect 3192 11118 3278 11174
rect 3334 11118 3408 11174
rect 3068 11032 3408 11118
rect 3068 10976 3136 11032
rect 3192 10976 3278 11032
rect 3334 10976 3408 11032
rect 3068 10890 3408 10976
rect 3068 10834 3136 10890
rect 3192 10834 3278 10890
rect 3334 10834 3408 10890
rect 3068 10748 3408 10834
rect 3068 10692 3136 10748
rect 3192 10692 3278 10748
rect 3334 10692 3408 10748
rect 3068 10606 3408 10692
rect 3068 10550 3136 10606
rect 3192 10550 3278 10606
rect 3334 10550 3408 10606
rect 3068 10464 3408 10550
rect 3068 10408 3136 10464
rect 3192 10408 3278 10464
rect 3334 10408 3408 10464
rect 3068 10322 3408 10408
rect 3068 10266 3136 10322
rect 3192 10266 3278 10322
rect 3334 10266 3408 10322
rect 3068 10180 3408 10266
rect 3068 10124 3136 10180
rect 3192 10124 3278 10180
rect 3334 10124 3408 10180
rect 3068 10038 3408 10124
rect 3068 9982 3136 10038
rect 3192 9982 3278 10038
rect 3334 9982 3408 10038
rect 3068 9896 3408 9982
rect 3068 9840 3136 9896
rect 3192 9840 3278 9896
rect 3334 9840 3408 9896
rect 3068 9754 3408 9840
rect 3068 9698 3136 9754
rect 3192 9698 3278 9754
rect 3334 9698 3408 9754
rect 3068 9612 3408 9698
rect 3068 9556 3136 9612
rect 3192 9556 3278 9612
rect 3334 9556 3408 9612
rect 3068 9470 3408 9556
rect 3068 9414 3136 9470
rect 3192 9414 3278 9470
rect 3334 9414 3408 9470
rect 3068 9328 3408 9414
rect 3068 9272 3136 9328
rect 3192 9272 3278 9328
rect 3334 9272 3408 9328
rect 3068 9186 3408 9272
rect 3068 9130 3136 9186
rect 3192 9130 3278 9186
rect 3334 9130 3408 9186
rect 3068 9044 3408 9130
rect 3068 8988 3136 9044
rect 3192 8988 3278 9044
rect 3334 8988 3408 9044
rect 3068 8902 3408 8988
rect 3068 8846 3136 8902
rect 3192 8846 3278 8902
rect 3334 8846 3408 8902
rect 3068 8760 3408 8846
rect 3068 8704 3136 8760
rect 3192 8704 3278 8760
rect 3334 8704 3408 8760
rect 3068 8618 3408 8704
rect 3068 8562 3136 8618
rect 3192 8562 3278 8618
rect 3334 8562 3408 8618
rect 3068 8476 3408 8562
rect 3068 8420 3136 8476
rect 3192 8420 3278 8476
rect 3334 8420 3408 8476
rect 3068 8334 3408 8420
rect 3068 8278 3136 8334
rect 3192 8278 3278 8334
rect 3334 8278 3408 8334
rect 3068 8192 3408 8278
rect 3068 8136 3136 8192
rect 3192 8136 3278 8192
rect 3334 8136 3408 8192
rect 3068 8050 3408 8136
rect 3068 7994 3136 8050
rect 3192 7994 3278 8050
rect 3334 7994 3408 8050
rect 3068 7908 3408 7994
rect 3068 7852 3136 7908
rect 3192 7852 3278 7908
rect 3334 7852 3408 7908
rect 3068 7766 3408 7852
rect 3068 7710 3136 7766
rect 3192 7710 3278 7766
rect 3334 7710 3408 7766
rect 3068 7624 3408 7710
rect 3068 7568 3136 7624
rect 3192 7568 3278 7624
rect 3334 7568 3408 7624
rect 3068 7482 3408 7568
rect 3068 7426 3136 7482
rect 3192 7426 3278 7482
rect 3334 7426 3408 7482
rect 3068 7340 3408 7426
rect 3068 7284 3136 7340
rect 3192 7284 3278 7340
rect 3334 7284 3408 7340
rect 3068 7198 3408 7284
rect 3068 7142 3136 7198
rect 3192 7142 3278 7198
rect 3334 7142 3408 7198
rect 3068 7056 3408 7142
rect 3068 7000 3136 7056
rect 3192 7000 3278 7056
rect 3334 7000 3408 7056
rect 3068 6914 3408 7000
rect 3068 6858 3136 6914
rect 3192 6858 3278 6914
rect 3334 6858 3408 6914
rect 3068 6772 3408 6858
rect 3068 6716 3136 6772
rect 3192 6716 3278 6772
rect 3334 6716 3408 6772
rect 3068 6630 3408 6716
rect 3068 6574 3136 6630
rect 3192 6574 3278 6630
rect 3334 6574 3408 6630
rect 3068 6488 3408 6574
rect 3068 6432 3136 6488
rect 3192 6432 3278 6488
rect 3334 6432 3408 6488
rect 3068 6346 3408 6432
rect 3068 6290 3136 6346
rect 3192 6290 3278 6346
rect 3334 6290 3408 6346
rect 3068 6204 3408 6290
rect 3068 6148 3136 6204
rect 3192 6148 3278 6204
rect 3334 6148 3408 6204
rect 3068 6062 3408 6148
rect 3068 6006 3136 6062
rect 3192 6006 3278 6062
rect 3334 6006 3408 6062
rect 3068 5920 3408 6006
rect 3068 5864 3136 5920
rect 3192 5864 3278 5920
rect 3334 5864 3408 5920
rect 3068 5778 3408 5864
rect 3068 5722 3136 5778
rect 3192 5722 3278 5778
rect 3334 5722 3408 5778
rect 3068 5636 3408 5722
rect 3068 5580 3136 5636
rect 3192 5580 3278 5636
rect 3334 5580 3408 5636
rect 3068 5494 3408 5580
rect 3068 5438 3136 5494
rect 3192 5438 3278 5494
rect 3334 5438 3408 5494
rect 3068 5352 3408 5438
rect 3068 5296 3136 5352
rect 3192 5296 3278 5352
rect 3334 5296 3408 5352
rect 3068 5210 3408 5296
rect 3068 5154 3136 5210
rect 3192 5154 3278 5210
rect 3334 5154 3408 5210
rect 3068 5068 3408 5154
rect 3068 5012 3136 5068
rect 3192 5012 3278 5068
rect 3334 5012 3408 5068
rect 3068 4926 3408 5012
rect 3068 4870 3136 4926
rect 3192 4870 3278 4926
rect 3334 4870 3408 4926
rect 3068 4784 3408 4870
rect 3068 4728 3136 4784
rect 3192 4728 3278 4784
rect 3334 4728 3408 4784
rect 3068 4642 3408 4728
rect 3068 4586 3136 4642
rect 3192 4586 3278 4642
rect 3334 4586 3408 4642
rect 3068 4500 3408 4586
rect 3068 4444 3136 4500
rect 3192 4444 3278 4500
rect 3334 4444 3408 4500
rect 3068 4358 3408 4444
rect 3068 4302 3136 4358
rect 3192 4302 3278 4358
rect 3334 4302 3408 4358
rect 3068 4216 3408 4302
rect 3068 4160 3136 4216
rect 3192 4160 3278 4216
rect 3334 4160 3408 4216
rect 3068 4074 3408 4160
rect 3068 4018 3136 4074
rect 3192 4018 3278 4074
rect 3334 4018 3408 4074
rect 3068 3932 3408 4018
rect 3068 3876 3136 3932
rect 3192 3876 3278 3932
rect 3334 3876 3408 3932
rect 3068 3790 3408 3876
rect 3068 3734 3136 3790
rect 3192 3734 3278 3790
rect 3334 3734 3408 3790
rect 3068 3648 3408 3734
rect 3068 3592 3136 3648
rect 3192 3592 3278 3648
rect 3334 3592 3408 3648
rect 3068 3506 3408 3592
rect 3068 3450 3136 3506
rect 3192 3450 3278 3506
rect 3334 3450 3408 3506
rect 3068 3364 3408 3450
rect 3068 3308 3136 3364
rect 3192 3308 3278 3364
rect 3334 3308 3408 3364
rect 3068 3222 3408 3308
rect 3068 3166 3136 3222
rect 3192 3166 3278 3222
rect 3334 3166 3408 3222
rect 3068 3080 3408 3166
rect 3068 3024 3136 3080
rect 3192 3024 3278 3080
rect 3334 3024 3408 3080
rect 3068 2938 3408 3024
rect 3068 2882 3136 2938
rect 3192 2882 3278 2938
rect 3334 2882 3408 2938
rect 3068 2796 3408 2882
rect 3068 2740 3136 2796
rect 3192 2740 3278 2796
rect 3334 2740 3408 2796
rect 3068 2654 3408 2740
rect 3068 2598 3136 2654
rect 3192 2598 3278 2654
rect 3334 2598 3408 2654
rect 3068 2512 3408 2598
rect 3068 2456 3136 2512
rect 3192 2456 3278 2512
rect 3334 2456 3408 2512
rect 3068 2370 3408 2456
rect 3068 2314 3136 2370
rect 3192 2314 3278 2370
rect 3334 2314 3408 2370
rect 3068 2228 3408 2314
rect 3068 2172 3136 2228
rect 3192 2172 3278 2228
rect 3334 2172 3408 2228
rect 3068 2086 3408 2172
rect 3068 2030 3136 2086
rect 3192 2030 3278 2086
rect 3334 2030 3408 2086
rect 3068 1944 3408 2030
rect 3068 1888 3136 1944
rect 3192 1888 3278 1944
rect 3334 1888 3408 1944
rect 3068 1802 3408 1888
rect 3068 1746 3136 1802
rect 3192 1746 3278 1802
rect 3334 1746 3408 1802
rect 3068 1660 3408 1746
rect 3068 1604 3136 1660
rect 3192 1604 3278 1660
rect 3334 1604 3408 1660
rect 3068 1518 3408 1604
rect 3068 1462 3136 1518
rect 3192 1462 3278 1518
rect 3334 1462 3408 1518
rect 3068 1376 3408 1462
rect 3068 1320 3136 1376
rect 3192 1320 3278 1376
rect 3334 1320 3408 1376
rect 3068 1234 3408 1320
rect 3068 1178 3136 1234
rect 3192 1178 3278 1234
rect 3334 1178 3408 1234
rect 3068 1092 3408 1178
rect 3068 1036 3136 1092
rect 3192 1036 3278 1092
rect 3334 1036 3408 1092
rect 3068 950 3408 1036
rect 3068 894 3136 950
rect 3192 894 3278 950
rect 3334 894 3408 950
rect 3068 808 3408 894
rect 3068 752 3136 808
rect 3192 752 3278 808
rect 3334 752 3408 808
rect 3068 666 3408 752
rect 3068 610 3136 666
rect 3192 610 3278 666
rect 3334 610 3408 666
rect 3068 524 3408 610
rect 3068 468 3136 524
rect 3192 468 3278 524
rect 3334 468 3408 524
rect 3068 400 3408 468
rect 3468 12310 3808 12400
rect 3468 12254 3536 12310
rect 3592 12254 3678 12310
rect 3734 12254 3808 12310
rect 3468 12168 3808 12254
rect 3468 12112 3536 12168
rect 3592 12112 3678 12168
rect 3734 12112 3808 12168
rect 3468 12026 3808 12112
rect 3468 11970 3536 12026
rect 3592 11970 3678 12026
rect 3734 11970 3808 12026
rect 3468 11884 3808 11970
rect 3468 11828 3536 11884
rect 3592 11828 3678 11884
rect 3734 11828 3808 11884
rect 3468 11742 3808 11828
rect 3468 11686 3536 11742
rect 3592 11686 3678 11742
rect 3734 11686 3808 11742
rect 3468 11600 3808 11686
rect 3468 11544 3536 11600
rect 3592 11544 3678 11600
rect 3734 11544 3808 11600
rect 3468 11458 3808 11544
rect 3468 11402 3536 11458
rect 3592 11402 3678 11458
rect 3734 11402 3808 11458
rect 3468 11316 3808 11402
rect 3468 11260 3536 11316
rect 3592 11260 3678 11316
rect 3734 11260 3808 11316
rect 3468 11174 3808 11260
rect 3468 11118 3536 11174
rect 3592 11118 3678 11174
rect 3734 11118 3808 11174
rect 3468 11032 3808 11118
rect 3468 10976 3536 11032
rect 3592 10976 3678 11032
rect 3734 10976 3808 11032
rect 3468 10890 3808 10976
rect 3468 10834 3536 10890
rect 3592 10834 3678 10890
rect 3734 10834 3808 10890
rect 3468 10748 3808 10834
rect 3468 10692 3536 10748
rect 3592 10692 3678 10748
rect 3734 10692 3808 10748
rect 3468 10606 3808 10692
rect 3468 10550 3536 10606
rect 3592 10550 3678 10606
rect 3734 10550 3808 10606
rect 3468 10464 3808 10550
rect 3468 10408 3536 10464
rect 3592 10408 3678 10464
rect 3734 10408 3808 10464
rect 3468 10322 3808 10408
rect 3468 10266 3536 10322
rect 3592 10266 3678 10322
rect 3734 10266 3808 10322
rect 3468 10180 3808 10266
rect 3468 10124 3536 10180
rect 3592 10124 3678 10180
rect 3734 10124 3808 10180
rect 3468 10038 3808 10124
rect 3468 9982 3536 10038
rect 3592 9982 3678 10038
rect 3734 9982 3808 10038
rect 3468 9896 3808 9982
rect 3468 9840 3536 9896
rect 3592 9840 3678 9896
rect 3734 9840 3808 9896
rect 3468 9754 3808 9840
rect 3468 9698 3536 9754
rect 3592 9698 3678 9754
rect 3734 9698 3808 9754
rect 3468 9612 3808 9698
rect 3468 9556 3536 9612
rect 3592 9556 3678 9612
rect 3734 9556 3808 9612
rect 3468 9470 3808 9556
rect 3468 9414 3536 9470
rect 3592 9414 3678 9470
rect 3734 9414 3808 9470
rect 3468 9328 3808 9414
rect 3468 9272 3536 9328
rect 3592 9272 3678 9328
rect 3734 9272 3808 9328
rect 3468 9186 3808 9272
rect 3468 9130 3536 9186
rect 3592 9130 3678 9186
rect 3734 9130 3808 9186
rect 3468 9044 3808 9130
rect 3468 8988 3536 9044
rect 3592 8988 3678 9044
rect 3734 8988 3808 9044
rect 3468 8902 3808 8988
rect 3468 8846 3536 8902
rect 3592 8846 3678 8902
rect 3734 8846 3808 8902
rect 3468 8760 3808 8846
rect 3468 8704 3536 8760
rect 3592 8704 3678 8760
rect 3734 8704 3808 8760
rect 3468 8618 3808 8704
rect 3468 8562 3536 8618
rect 3592 8562 3678 8618
rect 3734 8562 3808 8618
rect 3468 8476 3808 8562
rect 3468 8420 3536 8476
rect 3592 8420 3678 8476
rect 3734 8420 3808 8476
rect 3468 8334 3808 8420
rect 3468 8278 3536 8334
rect 3592 8278 3678 8334
rect 3734 8278 3808 8334
rect 3468 8192 3808 8278
rect 3468 8136 3536 8192
rect 3592 8136 3678 8192
rect 3734 8136 3808 8192
rect 3468 8050 3808 8136
rect 3468 7994 3536 8050
rect 3592 7994 3678 8050
rect 3734 7994 3808 8050
rect 3468 7908 3808 7994
rect 3468 7852 3536 7908
rect 3592 7852 3678 7908
rect 3734 7852 3808 7908
rect 3468 7766 3808 7852
rect 3468 7710 3536 7766
rect 3592 7710 3678 7766
rect 3734 7710 3808 7766
rect 3468 7624 3808 7710
rect 3468 7568 3536 7624
rect 3592 7568 3678 7624
rect 3734 7568 3808 7624
rect 3468 7482 3808 7568
rect 3468 7426 3536 7482
rect 3592 7426 3678 7482
rect 3734 7426 3808 7482
rect 3468 7340 3808 7426
rect 3468 7284 3536 7340
rect 3592 7284 3678 7340
rect 3734 7284 3808 7340
rect 3468 7198 3808 7284
rect 3468 7142 3536 7198
rect 3592 7142 3678 7198
rect 3734 7142 3808 7198
rect 3468 7056 3808 7142
rect 3468 7000 3536 7056
rect 3592 7000 3678 7056
rect 3734 7000 3808 7056
rect 3468 6914 3808 7000
rect 3468 6858 3536 6914
rect 3592 6858 3678 6914
rect 3734 6858 3808 6914
rect 3468 6772 3808 6858
rect 3468 6716 3536 6772
rect 3592 6716 3678 6772
rect 3734 6716 3808 6772
rect 3468 6630 3808 6716
rect 3468 6574 3536 6630
rect 3592 6574 3678 6630
rect 3734 6574 3808 6630
rect 3468 6488 3808 6574
rect 3468 6432 3536 6488
rect 3592 6432 3678 6488
rect 3734 6432 3808 6488
rect 3468 6346 3808 6432
rect 3468 6290 3536 6346
rect 3592 6290 3678 6346
rect 3734 6290 3808 6346
rect 3468 6204 3808 6290
rect 3468 6148 3536 6204
rect 3592 6148 3678 6204
rect 3734 6148 3808 6204
rect 3468 6062 3808 6148
rect 3468 6006 3536 6062
rect 3592 6006 3678 6062
rect 3734 6006 3808 6062
rect 3468 5920 3808 6006
rect 3468 5864 3536 5920
rect 3592 5864 3678 5920
rect 3734 5864 3808 5920
rect 3468 5778 3808 5864
rect 3468 5722 3536 5778
rect 3592 5722 3678 5778
rect 3734 5722 3808 5778
rect 3468 5636 3808 5722
rect 3468 5580 3536 5636
rect 3592 5580 3678 5636
rect 3734 5580 3808 5636
rect 3468 5494 3808 5580
rect 3468 5438 3536 5494
rect 3592 5438 3678 5494
rect 3734 5438 3808 5494
rect 3468 5352 3808 5438
rect 3468 5296 3536 5352
rect 3592 5296 3678 5352
rect 3734 5296 3808 5352
rect 3468 5210 3808 5296
rect 3468 5154 3536 5210
rect 3592 5154 3678 5210
rect 3734 5154 3808 5210
rect 3468 5068 3808 5154
rect 3468 5012 3536 5068
rect 3592 5012 3678 5068
rect 3734 5012 3808 5068
rect 3468 4926 3808 5012
rect 3468 4870 3536 4926
rect 3592 4870 3678 4926
rect 3734 4870 3808 4926
rect 3468 4784 3808 4870
rect 3468 4728 3536 4784
rect 3592 4728 3678 4784
rect 3734 4728 3808 4784
rect 3468 4642 3808 4728
rect 3468 4586 3536 4642
rect 3592 4586 3678 4642
rect 3734 4586 3808 4642
rect 3468 4500 3808 4586
rect 3468 4444 3536 4500
rect 3592 4444 3678 4500
rect 3734 4444 3808 4500
rect 3468 4358 3808 4444
rect 3468 4302 3536 4358
rect 3592 4302 3678 4358
rect 3734 4302 3808 4358
rect 3468 4216 3808 4302
rect 3468 4160 3536 4216
rect 3592 4160 3678 4216
rect 3734 4160 3808 4216
rect 3468 4074 3808 4160
rect 3468 4018 3536 4074
rect 3592 4018 3678 4074
rect 3734 4018 3808 4074
rect 3468 3932 3808 4018
rect 3468 3876 3536 3932
rect 3592 3876 3678 3932
rect 3734 3876 3808 3932
rect 3468 3790 3808 3876
rect 3468 3734 3536 3790
rect 3592 3734 3678 3790
rect 3734 3734 3808 3790
rect 3468 3648 3808 3734
rect 3468 3592 3536 3648
rect 3592 3592 3678 3648
rect 3734 3592 3808 3648
rect 3468 3506 3808 3592
rect 3468 3450 3536 3506
rect 3592 3450 3678 3506
rect 3734 3450 3808 3506
rect 3468 3364 3808 3450
rect 3468 3308 3536 3364
rect 3592 3308 3678 3364
rect 3734 3308 3808 3364
rect 3468 3222 3808 3308
rect 3468 3166 3536 3222
rect 3592 3166 3678 3222
rect 3734 3166 3808 3222
rect 3468 3080 3808 3166
rect 3468 3024 3536 3080
rect 3592 3024 3678 3080
rect 3734 3024 3808 3080
rect 3468 2938 3808 3024
rect 3468 2882 3536 2938
rect 3592 2882 3678 2938
rect 3734 2882 3808 2938
rect 3468 2796 3808 2882
rect 3468 2740 3536 2796
rect 3592 2740 3678 2796
rect 3734 2740 3808 2796
rect 3468 2654 3808 2740
rect 3468 2598 3536 2654
rect 3592 2598 3678 2654
rect 3734 2598 3808 2654
rect 3468 2512 3808 2598
rect 3468 2456 3536 2512
rect 3592 2456 3678 2512
rect 3734 2456 3808 2512
rect 3468 2370 3808 2456
rect 3468 2314 3536 2370
rect 3592 2314 3678 2370
rect 3734 2314 3808 2370
rect 3468 2228 3808 2314
rect 3468 2172 3536 2228
rect 3592 2172 3678 2228
rect 3734 2172 3808 2228
rect 3468 2086 3808 2172
rect 3468 2030 3536 2086
rect 3592 2030 3678 2086
rect 3734 2030 3808 2086
rect 3468 1944 3808 2030
rect 3468 1888 3536 1944
rect 3592 1888 3678 1944
rect 3734 1888 3808 1944
rect 3468 1802 3808 1888
rect 3468 1746 3536 1802
rect 3592 1746 3678 1802
rect 3734 1746 3808 1802
rect 3468 1660 3808 1746
rect 3468 1604 3536 1660
rect 3592 1604 3678 1660
rect 3734 1604 3808 1660
rect 3468 1518 3808 1604
rect 3468 1462 3536 1518
rect 3592 1462 3678 1518
rect 3734 1462 3808 1518
rect 3468 1376 3808 1462
rect 3468 1320 3536 1376
rect 3592 1320 3678 1376
rect 3734 1320 3808 1376
rect 3468 1234 3808 1320
rect 3468 1178 3536 1234
rect 3592 1178 3678 1234
rect 3734 1178 3808 1234
rect 3468 1092 3808 1178
rect 3468 1036 3536 1092
rect 3592 1036 3678 1092
rect 3734 1036 3808 1092
rect 3468 950 3808 1036
rect 3468 894 3536 950
rect 3592 894 3678 950
rect 3734 894 3808 950
rect 3468 808 3808 894
rect 3468 752 3536 808
rect 3592 752 3678 808
rect 3734 752 3808 808
rect 3468 666 3808 752
rect 3468 610 3536 666
rect 3592 610 3678 666
rect 3734 610 3808 666
rect 3468 524 3808 610
rect 3468 468 3536 524
rect 3592 468 3678 524
rect 3734 468 3808 524
rect 3468 400 3808 468
rect 3868 12310 4208 12400
rect 3868 12254 3933 12310
rect 3989 12254 4075 12310
rect 4131 12254 4208 12310
rect 3868 12168 4208 12254
rect 3868 12112 3933 12168
rect 3989 12112 4075 12168
rect 4131 12112 4208 12168
rect 3868 12026 4208 12112
rect 3868 11970 3933 12026
rect 3989 11970 4075 12026
rect 4131 11970 4208 12026
rect 3868 11884 4208 11970
rect 3868 11828 3933 11884
rect 3989 11828 4075 11884
rect 4131 11828 4208 11884
rect 3868 11742 4208 11828
rect 3868 11686 3933 11742
rect 3989 11686 4075 11742
rect 4131 11686 4208 11742
rect 3868 11600 4208 11686
rect 3868 11544 3933 11600
rect 3989 11544 4075 11600
rect 4131 11544 4208 11600
rect 3868 11458 4208 11544
rect 3868 11402 3933 11458
rect 3989 11402 4075 11458
rect 4131 11402 4208 11458
rect 3868 11316 4208 11402
rect 3868 11260 3933 11316
rect 3989 11260 4075 11316
rect 4131 11260 4208 11316
rect 3868 11174 4208 11260
rect 3868 11118 3933 11174
rect 3989 11118 4075 11174
rect 4131 11118 4208 11174
rect 3868 11032 4208 11118
rect 3868 10976 3933 11032
rect 3989 10976 4075 11032
rect 4131 10976 4208 11032
rect 3868 10890 4208 10976
rect 3868 10834 3933 10890
rect 3989 10834 4075 10890
rect 4131 10834 4208 10890
rect 3868 10748 4208 10834
rect 3868 10692 3933 10748
rect 3989 10692 4075 10748
rect 4131 10692 4208 10748
rect 3868 10606 4208 10692
rect 3868 10550 3933 10606
rect 3989 10550 4075 10606
rect 4131 10550 4208 10606
rect 3868 10464 4208 10550
rect 3868 10408 3933 10464
rect 3989 10408 4075 10464
rect 4131 10408 4208 10464
rect 3868 10322 4208 10408
rect 3868 10266 3933 10322
rect 3989 10266 4075 10322
rect 4131 10266 4208 10322
rect 3868 10180 4208 10266
rect 3868 10124 3933 10180
rect 3989 10124 4075 10180
rect 4131 10124 4208 10180
rect 3868 10038 4208 10124
rect 3868 9982 3933 10038
rect 3989 9982 4075 10038
rect 4131 9982 4208 10038
rect 3868 9896 4208 9982
rect 3868 9840 3933 9896
rect 3989 9840 4075 9896
rect 4131 9840 4208 9896
rect 3868 9754 4208 9840
rect 3868 9698 3933 9754
rect 3989 9698 4075 9754
rect 4131 9698 4208 9754
rect 3868 9612 4208 9698
rect 3868 9556 3933 9612
rect 3989 9556 4075 9612
rect 4131 9556 4208 9612
rect 3868 9470 4208 9556
rect 3868 9414 3933 9470
rect 3989 9414 4075 9470
rect 4131 9414 4208 9470
rect 3868 9328 4208 9414
rect 3868 9272 3933 9328
rect 3989 9272 4075 9328
rect 4131 9272 4208 9328
rect 3868 9186 4208 9272
rect 3868 9130 3933 9186
rect 3989 9130 4075 9186
rect 4131 9130 4208 9186
rect 3868 9044 4208 9130
rect 3868 8988 3933 9044
rect 3989 8988 4075 9044
rect 4131 8988 4208 9044
rect 3868 8902 4208 8988
rect 3868 8846 3933 8902
rect 3989 8846 4075 8902
rect 4131 8846 4208 8902
rect 3868 8760 4208 8846
rect 3868 8704 3933 8760
rect 3989 8704 4075 8760
rect 4131 8704 4208 8760
rect 3868 8618 4208 8704
rect 3868 8562 3933 8618
rect 3989 8562 4075 8618
rect 4131 8562 4208 8618
rect 3868 8476 4208 8562
rect 3868 8420 3933 8476
rect 3989 8420 4075 8476
rect 4131 8420 4208 8476
rect 3868 8334 4208 8420
rect 3868 8278 3933 8334
rect 3989 8278 4075 8334
rect 4131 8278 4208 8334
rect 3868 8192 4208 8278
rect 3868 8136 3933 8192
rect 3989 8136 4075 8192
rect 4131 8136 4208 8192
rect 3868 8050 4208 8136
rect 3868 7994 3933 8050
rect 3989 7994 4075 8050
rect 4131 7994 4208 8050
rect 3868 7908 4208 7994
rect 3868 7852 3933 7908
rect 3989 7852 4075 7908
rect 4131 7852 4208 7908
rect 3868 7766 4208 7852
rect 3868 7710 3933 7766
rect 3989 7710 4075 7766
rect 4131 7710 4208 7766
rect 3868 7624 4208 7710
rect 3868 7568 3933 7624
rect 3989 7568 4075 7624
rect 4131 7568 4208 7624
rect 3868 7482 4208 7568
rect 3868 7426 3933 7482
rect 3989 7426 4075 7482
rect 4131 7426 4208 7482
rect 3868 7340 4208 7426
rect 3868 7284 3933 7340
rect 3989 7284 4075 7340
rect 4131 7284 4208 7340
rect 3868 7198 4208 7284
rect 3868 7142 3933 7198
rect 3989 7142 4075 7198
rect 4131 7142 4208 7198
rect 3868 7056 4208 7142
rect 3868 7000 3933 7056
rect 3989 7000 4075 7056
rect 4131 7000 4208 7056
rect 3868 6914 4208 7000
rect 3868 6858 3933 6914
rect 3989 6858 4075 6914
rect 4131 6858 4208 6914
rect 3868 6772 4208 6858
rect 3868 6716 3933 6772
rect 3989 6716 4075 6772
rect 4131 6716 4208 6772
rect 3868 6630 4208 6716
rect 3868 6574 3933 6630
rect 3989 6574 4075 6630
rect 4131 6574 4208 6630
rect 3868 6488 4208 6574
rect 3868 6432 3933 6488
rect 3989 6432 4075 6488
rect 4131 6432 4208 6488
rect 3868 6346 4208 6432
rect 3868 6290 3933 6346
rect 3989 6290 4075 6346
rect 4131 6290 4208 6346
rect 3868 6204 4208 6290
rect 3868 6148 3933 6204
rect 3989 6148 4075 6204
rect 4131 6148 4208 6204
rect 3868 6062 4208 6148
rect 3868 6006 3933 6062
rect 3989 6006 4075 6062
rect 4131 6006 4208 6062
rect 3868 5920 4208 6006
rect 3868 5864 3933 5920
rect 3989 5864 4075 5920
rect 4131 5864 4208 5920
rect 3868 5778 4208 5864
rect 3868 5722 3933 5778
rect 3989 5722 4075 5778
rect 4131 5722 4208 5778
rect 3868 5636 4208 5722
rect 3868 5580 3933 5636
rect 3989 5580 4075 5636
rect 4131 5580 4208 5636
rect 3868 5494 4208 5580
rect 3868 5438 3933 5494
rect 3989 5438 4075 5494
rect 4131 5438 4208 5494
rect 3868 5352 4208 5438
rect 3868 5296 3933 5352
rect 3989 5296 4075 5352
rect 4131 5296 4208 5352
rect 3868 5210 4208 5296
rect 3868 5154 3933 5210
rect 3989 5154 4075 5210
rect 4131 5154 4208 5210
rect 3868 5068 4208 5154
rect 3868 5012 3933 5068
rect 3989 5012 4075 5068
rect 4131 5012 4208 5068
rect 3868 4926 4208 5012
rect 3868 4870 3933 4926
rect 3989 4870 4075 4926
rect 4131 4870 4208 4926
rect 3868 4784 4208 4870
rect 3868 4728 3933 4784
rect 3989 4728 4075 4784
rect 4131 4728 4208 4784
rect 3868 4642 4208 4728
rect 3868 4586 3933 4642
rect 3989 4586 4075 4642
rect 4131 4586 4208 4642
rect 3868 4500 4208 4586
rect 3868 4444 3933 4500
rect 3989 4444 4075 4500
rect 4131 4444 4208 4500
rect 3868 4358 4208 4444
rect 3868 4302 3933 4358
rect 3989 4302 4075 4358
rect 4131 4302 4208 4358
rect 3868 4216 4208 4302
rect 3868 4160 3933 4216
rect 3989 4160 4075 4216
rect 4131 4160 4208 4216
rect 3868 4074 4208 4160
rect 3868 4018 3933 4074
rect 3989 4018 4075 4074
rect 4131 4018 4208 4074
rect 3868 3932 4208 4018
rect 3868 3876 3933 3932
rect 3989 3876 4075 3932
rect 4131 3876 4208 3932
rect 3868 3790 4208 3876
rect 3868 3734 3933 3790
rect 3989 3734 4075 3790
rect 4131 3734 4208 3790
rect 3868 3648 4208 3734
rect 3868 3592 3933 3648
rect 3989 3592 4075 3648
rect 4131 3592 4208 3648
rect 3868 3506 4208 3592
rect 3868 3450 3933 3506
rect 3989 3450 4075 3506
rect 4131 3450 4208 3506
rect 3868 3364 4208 3450
rect 3868 3308 3933 3364
rect 3989 3308 4075 3364
rect 4131 3308 4208 3364
rect 3868 3222 4208 3308
rect 3868 3166 3933 3222
rect 3989 3166 4075 3222
rect 4131 3166 4208 3222
rect 3868 3080 4208 3166
rect 3868 3024 3933 3080
rect 3989 3024 4075 3080
rect 4131 3024 4208 3080
rect 3868 2938 4208 3024
rect 3868 2882 3933 2938
rect 3989 2882 4075 2938
rect 4131 2882 4208 2938
rect 3868 2796 4208 2882
rect 3868 2740 3933 2796
rect 3989 2740 4075 2796
rect 4131 2740 4208 2796
rect 3868 2654 4208 2740
rect 3868 2598 3933 2654
rect 3989 2598 4075 2654
rect 4131 2598 4208 2654
rect 3868 2512 4208 2598
rect 3868 2456 3933 2512
rect 3989 2456 4075 2512
rect 4131 2456 4208 2512
rect 3868 2370 4208 2456
rect 3868 2314 3933 2370
rect 3989 2314 4075 2370
rect 4131 2314 4208 2370
rect 3868 2228 4208 2314
rect 3868 2172 3933 2228
rect 3989 2172 4075 2228
rect 4131 2172 4208 2228
rect 3868 2086 4208 2172
rect 3868 2030 3933 2086
rect 3989 2030 4075 2086
rect 4131 2030 4208 2086
rect 3868 1944 4208 2030
rect 3868 1888 3933 1944
rect 3989 1888 4075 1944
rect 4131 1888 4208 1944
rect 3868 1802 4208 1888
rect 3868 1746 3933 1802
rect 3989 1746 4075 1802
rect 4131 1746 4208 1802
rect 3868 1660 4208 1746
rect 3868 1604 3933 1660
rect 3989 1604 4075 1660
rect 4131 1604 4208 1660
rect 3868 1518 4208 1604
rect 3868 1462 3933 1518
rect 3989 1462 4075 1518
rect 4131 1462 4208 1518
rect 3868 1376 4208 1462
rect 3868 1320 3933 1376
rect 3989 1320 4075 1376
rect 4131 1320 4208 1376
rect 3868 1234 4208 1320
rect 3868 1178 3933 1234
rect 3989 1178 4075 1234
rect 4131 1178 4208 1234
rect 3868 1092 4208 1178
rect 3868 1036 3933 1092
rect 3989 1036 4075 1092
rect 4131 1036 4208 1092
rect 3868 950 4208 1036
rect 3868 894 3933 950
rect 3989 894 4075 950
rect 4131 894 4208 950
rect 3868 808 4208 894
rect 3868 752 3933 808
rect 3989 752 4075 808
rect 4131 752 4208 808
rect 3868 666 4208 752
rect 3868 610 3933 666
rect 3989 610 4075 666
rect 4131 610 4208 666
rect 3868 524 4208 610
rect 3868 468 3933 524
rect 3989 468 4075 524
rect 4131 468 4208 524
rect 3868 400 4208 468
rect 4268 12310 4608 12400
rect 4268 12254 4338 12310
rect 4394 12254 4480 12310
rect 4536 12254 4608 12310
rect 4268 12168 4608 12254
rect 4268 12112 4338 12168
rect 4394 12112 4480 12168
rect 4536 12112 4608 12168
rect 4268 12026 4608 12112
rect 4268 11970 4338 12026
rect 4394 11970 4480 12026
rect 4536 11970 4608 12026
rect 4268 11884 4608 11970
rect 4268 11828 4338 11884
rect 4394 11828 4480 11884
rect 4536 11828 4608 11884
rect 4268 11742 4608 11828
rect 4268 11686 4338 11742
rect 4394 11686 4480 11742
rect 4536 11686 4608 11742
rect 4268 11600 4608 11686
rect 4268 11544 4338 11600
rect 4394 11544 4480 11600
rect 4536 11544 4608 11600
rect 4268 11458 4608 11544
rect 4268 11402 4338 11458
rect 4394 11402 4480 11458
rect 4536 11402 4608 11458
rect 4268 11316 4608 11402
rect 4268 11260 4338 11316
rect 4394 11260 4480 11316
rect 4536 11260 4608 11316
rect 4268 11174 4608 11260
rect 4268 11118 4338 11174
rect 4394 11118 4480 11174
rect 4536 11118 4608 11174
rect 4268 11032 4608 11118
rect 4268 10976 4338 11032
rect 4394 10976 4480 11032
rect 4536 10976 4608 11032
rect 4268 10890 4608 10976
rect 4268 10834 4338 10890
rect 4394 10834 4480 10890
rect 4536 10834 4608 10890
rect 4268 10748 4608 10834
rect 4268 10692 4338 10748
rect 4394 10692 4480 10748
rect 4536 10692 4608 10748
rect 4268 10606 4608 10692
rect 4268 10550 4338 10606
rect 4394 10550 4480 10606
rect 4536 10550 4608 10606
rect 4268 10464 4608 10550
rect 4268 10408 4338 10464
rect 4394 10408 4480 10464
rect 4536 10408 4608 10464
rect 4268 10322 4608 10408
rect 4268 10266 4338 10322
rect 4394 10266 4480 10322
rect 4536 10266 4608 10322
rect 4268 10180 4608 10266
rect 4268 10124 4338 10180
rect 4394 10124 4480 10180
rect 4536 10124 4608 10180
rect 4268 10038 4608 10124
rect 4268 9982 4338 10038
rect 4394 9982 4480 10038
rect 4536 9982 4608 10038
rect 4268 9896 4608 9982
rect 4268 9840 4338 9896
rect 4394 9840 4480 9896
rect 4536 9840 4608 9896
rect 4268 9754 4608 9840
rect 4268 9698 4338 9754
rect 4394 9698 4480 9754
rect 4536 9698 4608 9754
rect 4268 9612 4608 9698
rect 4268 9556 4338 9612
rect 4394 9556 4480 9612
rect 4536 9556 4608 9612
rect 4268 9470 4608 9556
rect 4268 9414 4338 9470
rect 4394 9414 4480 9470
rect 4536 9414 4608 9470
rect 4268 9328 4608 9414
rect 4268 9272 4338 9328
rect 4394 9272 4480 9328
rect 4536 9272 4608 9328
rect 4268 9186 4608 9272
rect 4268 9130 4338 9186
rect 4394 9130 4480 9186
rect 4536 9130 4608 9186
rect 4268 9044 4608 9130
rect 4268 8988 4338 9044
rect 4394 8988 4480 9044
rect 4536 8988 4608 9044
rect 4268 8902 4608 8988
rect 4268 8846 4338 8902
rect 4394 8846 4480 8902
rect 4536 8846 4608 8902
rect 4268 8760 4608 8846
rect 4268 8704 4338 8760
rect 4394 8704 4480 8760
rect 4536 8704 4608 8760
rect 4268 8618 4608 8704
rect 4268 8562 4338 8618
rect 4394 8562 4480 8618
rect 4536 8562 4608 8618
rect 4268 8476 4608 8562
rect 4268 8420 4338 8476
rect 4394 8420 4480 8476
rect 4536 8420 4608 8476
rect 4268 8334 4608 8420
rect 4268 8278 4338 8334
rect 4394 8278 4480 8334
rect 4536 8278 4608 8334
rect 4268 8192 4608 8278
rect 4268 8136 4338 8192
rect 4394 8136 4480 8192
rect 4536 8136 4608 8192
rect 4268 8050 4608 8136
rect 4268 7994 4338 8050
rect 4394 7994 4480 8050
rect 4536 7994 4608 8050
rect 4268 7908 4608 7994
rect 4268 7852 4338 7908
rect 4394 7852 4480 7908
rect 4536 7852 4608 7908
rect 4268 7766 4608 7852
rect 4268 7710 4338 7766
rect 4394 7710 4480 7766
rect 4536 7710 4608 7766
rect 4268 7624 4608 7710
rect 4268 7568 4338 7624
rect 4394 7568 4480 7624
rect 4536 7568 4608 7624
rect 4268 7482 4608 7568
rect 4268 7426 4338 7482
rect 4394 7426 4480 7482
rect 4536 7426 4608 7482
rect 4268 7340 4608 7426
rect 4268 7284 4338 7340
rect 4394 7284 4480 7340
rect 4536 7284 4608 7340
rect 4268 7198 4608 7284
rect 4268 7142 4338 7198
rect 4394 7142 4480 7198
rect 4536 7142 4608 7198
rect 4268 7056 4608 7142
rect 4268 7000 4338 7056
rect 4394 7000 4480 7056
rect 4536 7000 4608 7056
rect 4268 6914 4608 7000
rect 4268 6858 4338 6914
rect 4394 6858 4480 6914
rect 4536 6858 4608 6914
rect 4268 6772 4608 6858
rect 4268 6716 4338 6772
rect 4394 6716 4480 6772
rect 4536 6716 4608 6772
rect 4268 6630 4608 6716
rect 4268 6574 4338 6630
rect 4394 6574 4480 6630
rect 4536 6574 4608 6630
rect 4268 6488 4608 6574
rect 4268 6432 4338 6488
rect 4394 6432 4480 6488
rect 4536 6432 4608 6488
rect 4268 6346 4608 6432
rect 4268 6290 4338 6346
rect 4394 6290 4480 6346
rect 4536 6290 4608 6346
rect 4268 6204 4608 6290
rect 4268 6148 4338 6204
rect 4394 6148 4480 6204
rect 4536 6148 4608 6204
rect 4268 6062 4608 6148
rect 4268 6006 4338 6062
rect 4394 6006 4480 6062
rect 4536 6006 4608 6062
rect 4268 5920 4608 6006
rect 4268 5864 4338 5920
rect 4394 5864 4480 5920
rect 4536 5864 4608 5920
rect 4268 5778 4608 5864
rect 4268 5722 4338 5778
rect 4394 5722 4480 5778
rect 4536 5722 4608 5778
rect 4268 5636 4608 5722
rect 4268 5580 4338 5636
rect 4394 5580 4480 5636
rect 4536 5580 4608 5636
rect 4268 5494 4608 5580
rect 4268 5438 4338 5494
rect 4394 5438 4480 5494
rect 4536 5438 4608 5494
rect 4268 5352 4608 5438
rect 4268 5296 4338 5352
rect 4394 5296 4480 5352
rect 4536 5296 4608 5352
rect 4268 5210 4608 5296
rect 4268 5154 4338 5210
rect 4394 5154 4480 5210
rect 4536 5154 4608 5210
rect 4268 5068 4608 5154
rect 4268 5012 4338 5068
rect 4394 5012 4480 5068
rect 4536 5012 4608 5068
rect 4268 4926 4608 5012
rect 4268 4870 4338 4926
rect 4394 4870 4480 4926
rect 4536 4870 4608 4926
rect 4268 4784 4608 4870
rect 4268 4728 4338 4784
rect 4394 4728 4480 4784
rect 4536 4728 4608 4784
rect 4268 4642 4608 4728
rect 4268 4586 4338 4642
rect 4394 4586 4480 4642
rect 4536 4586 4608 4642
rect 4268 4500 4608 4586
rect 4268 4444 4338 4500
rect 4394 4444 4480 4500
rect 4536 4444 4608 4500
rect 4268 4358 4608 4444
rect 4268 4302 4338 4358
rect 4394 4302 4480 4358
rect 4536 4302 4608 4358
rect 4268 4216 4608 4302
rect 4268 4160 4338 4216
rect 4394 4160 4480 4216
rect 4536 4160 4608 4216
rect 4268 4074 4608 4160
rect 4268 4018 4338 4074
rect 4394 4018 4480 4074
rect 4536 4018 4608 4074
rect 4268 3932 4608 4018
rect 4268 3876 4338 3932
rect 4394 3876 4480 3932
rect 4536 3876 4608 3932
rect 4268 3790 4608 3876
rect 4268 3734 4338 3790
rect 4394 3734 4480 3790
rect 4536 3734 4608 3790
rect 4268 3648 4608 3734
rect 4268 3592 4338 3648
rect 4394 3592 4480 3648
rect 4536 3592 4608 3648
rect 4268 3506 4608 3592
rect 4268 3450 4338 3506
rect 4394 3450 4480 3506
rect 4536 3450 4608 3506
rect 4268 3364 4608 3450
rect 4268 3308 4338 3364
rect 4394 3308 4480 3364
rect 4536 3308 4608 3364
rect 4268 3222 4608 3308
rect 4268 3166 4338 3222
rect 4394 3166 4480 3222
rect 4536 3166 4608 3222
rect 4268 3080 4608 3166
rect 4268 3024 4338 3080
rect 4394 3024 4480 3080
rect 4536 3024 4608 3080
rect 4268 2938 4608 3024
rect 4268 2882 4338 2938
rect 4394 2882 4480 2938
rect 4536 2882 4608 2938
rect 4268 2796 4608 2882
rect 4268 2740 4338 2796
rect 4394 2740 4480 2796
rect 4536 2740 4608 2796
rect 4268 2654 4608 2740
rect 4268 2598 4338 2654
rect 4394 2598 4480 2654
rect 4536 2598 4608 2654
rect 4268 2512 4608 2598
rect 4268 2456 4338 2512
rect 4394 2456 4480 2512
rect 4536 2456 4608 2512
rect 4268 2370 4608 2456
rect 4268 2314 4338 2370
rect 4394 2314 4480 2370
rect 4536 2314 4608 2370
rect 4268 2228 4608 2314
rect 4268 2172 4338 2228
rect 4394 2172 4480 2228
rect 4536 2172 4608 2228
rect 4268 2086 4608 2172
rect 4268 2030 4338 2086
rect 4394 2030 4480 2086
rect 4536 2030 4608 2086
rect 4268 1944 4608 2030
rect 4268 1888 4338 1944
rect 4394 1888 4480 1944
rect 4536 1888 4608 1944
rect 4268 1802 4608 1888
rect 4268 1746 4338 1802
rect 4394 1746 4480 1802
rect 4536 1746 4608 1802
rect 4268 1660 4608 1746
rect 4268 1604 4338 1660
rect 4394 1604 4480 1660
rect 4536 1604 4608 1660
rect 4268 1518 4608 1604
rect 4268 1462 4338 1518
rect 4394 1462 4480 1518
rect 4536 1462 4608 1518
rect 4268 1376 4608 1462
rect 4268 1320 4338 1376
rect 4394 1320 4480 1376
rect 4536 1320 4608 1376
rect 4268 1234 4608 1320
rect 4268 1178 4338 1234
rect 4394 1178 4480 1234
rect 4536 1178 4608 1234
rect 4268 1092 4608 1178
rect 4268 1036 4338 1092
rect 4394 1036 4480 1092
rect 4536 1036 4608 1092
rect 4268 950 4608 1036
rect 4268 894 4338 950
rect 4394 894 4480 950
rect 4536 894 4608 950
rect 4268 808 4608 894
rect 4268 752 4338 808
rect 4394 752 4480 808
rect 4536 752 4608 808
rect 4268 666 4608 752
rect 4268 610 4338 666
rect 4394 610 4480 666
rect 4536 610 4608 666
rect 4268 524 4608 610
rect 4268 468 4338 524
rect 4394 468 4480 524
rect 4536 468 4608 524
rect 4268 400 4608 468
rect 4668 12310 5008 12400
rect 4668 12254 4738 12310
rect 4794 12254 4880 12310
rect 4936 12254 5008 12310
rect 4668 12168 5008 12254
rect 4668 12112 4738 12168
rect 4794 12112 4880 12168
rect 4936 12112 5008 12168
rect 4668 12026 5008 12112
rect 4668 11970 4738 12026
rect 4794 11970 4880 12026
rect 4936 11970 5008 12026
rect 4668 11884 5008 11970
rect 4668 11828 4738 11884
rect 4794 11828 4880 11884
rect 4936 11828 5008 11884
rect 4668 11742 5008 11828
rect 4668 11686 4738 11742
rect 4794 11686 4880 11742
rect 4936 11686 5008 11742
rect 4668 11600 5008 11686
rect 4668 11544 4738 11600
rect 4794 11544 4880 11600
rect 4936 11544 5008 11600
rect 4668 11458 5008 11544
rect 4668 11402 4738 11458
rect 4794 11402 4880 11458
rect 4936 11402 5008 11458
rect 4668 11316 5008 11402
rect 4668 11260 4738 11316
rect 4794 11260 4880 11316
rect 4936 11260 5008 11316
rect 4668 11174 5008 11260
rect 4668 11118 4738 11174
rect 4794 11118 4880 11174
rect 4936 11118 5008 11174
rect 4668 11032 5008 11118
rect 4668 10976 4738 11032
rect 4794 10976 4880 11032
rect 4936 10976 5008 11032
rect 4668 10890 5008 10976
rect 4668 10834 4738 10890
rect 4794 10834 4880 10890
rect 4936 10834 5008 10890
rect 4668 10748 5008 10834
rect 4668 10692 4738 10748
rect 4794 10692 4880 10748
rect 4936 10692 5008 10748
rect 4668 10606 5008 10692
rect 4668 10550 4738 10606
rect 4794 10550 4880 10606
rect 4936 10550 5008 10606
rect 4668 10464 5008 10550
rect 4668 10408 4738 10464
rect 4794 10408 4880 10464
rect 4936 10408 5008 10464
rect 4668 10322 5008 10408
rect 4668 10266 4738 10322
rect 4794 10266 4880 10322
rect 4936 10266 5008 10322
rect 4668 10180 5008 10266
rect 4668 10124 4738 10180
rect 4794 10124 4880 10180
rect 4936 10124 5008 10180
rect 4668 10038 5008 10124
rect 4668 9982 4738 10038
rect 4794 9982 4880 10038
rect 4936 9982 5008 10038
rect 4668 9896 5008 9982
rect 4668 9840 4738 9896
rect 4794 9840 4880 9896
rect 4936 9840 5008 9896
rect 4668 9754 5008 9840
rect 4668 9698 4738 9754
rect 4794 9698 4880 9754
rect 4936 9698 5008 9754
rect 4668 9612 5008 9698
rect 4668 9556 4738 9612
rect 4794 9556 4880 9612
rect 4936 9556 5008 9612
rect 4668 9470 5008 9556
rect 4668 9414 4738 9470
rect 4794 9414 4880 9470
rect 4936 9414 5008 9470
rect 4668 9328 5008 9414
rect 4668 9272 4738 9328
rect 4794 9272 4880 9328
rect 4936 9272 5008 9328
rect 4668 9186 5008 9272
rect 4668 9130 4738 9186
rect 4794 9130 4880 9186
rect 4936 9130 5008 9186
rect 4668 9044 5008 9130
rect 4668 8988 4738 9044
rect 4794 8988 4880 9044
rect 4936 8988 5008 9044
rect 4668 8902 5008 8988
rect 4668 8846 4738 8902
rect 4794 8846 4880 8902
rect 4936 8846 5008 8902
rect 4668 8760 5008 8846
rect 4668 8704 4738 8760
rect 4794 8704 4880 8760
rect 4936 8704 5008 8760
rect 4668 8618 5008 8704
rect 4668 8562 4738 8618
rect 4794 8562 4880 8618
rect 4936 8562 5008 8618
rect 4668 8476 5008 8562
rect 4668 8420 4738 8476
rect 4794 8420 4880 8476
rect 4936 8420 5008 8476
rect 4668 8334 5008 8420
rect 4668 8278 4738 8334
rect 4794 8278 4880 8334
rect 4936 8278 5008 8334
rect 4668 8192 5008 8278
rect 4668 8136 4738 8192
rect 4794 8136 4880 8192
rect 4936 8136 5008 8192
rect 4668 8050 5008 8136
rect 4668 7994 4738 8050
rect 4794 7994 4880 8050
rect 4936 7994 5008 8050
rect 4668 7908 5008 7994
rect 4668 7852 4738 7908
rect 4794 7852 4880 7908
rect 4936 7852 5008 7908
rect 4668 7766 5008 7852
rect 4668 7710 4738 7766
rect 4794 7710 4880 7766
rect 4936 7710 5008 7766
rect 4668 7624 5008 7710
rect 4668 7568 4738 7624
rect 4794 7568 4880 7624
rect 4936 7568 5008 7624
rect 4668 7482 5008 7568
rect 4668 7426 4738 7482
rect 4794 7426 4880 7482
rect 4936 7426 5008 7482
rect 4668 7340 5008 7426
rect 4668 7284 4738 7340
rect 4794 7284 4880 7340
rect 4936 7284 5008 7340
rect 4668 7198 5008 7284
rect 4668 7142 4738 7198
rect 4794 7142 4880 7198
rect 4936 7142 5008 7198
rect 4668 7056 5008 7142
rect 4668 7000 4738 7056
rect 4794 7000 4880 7056
rect 4936 7000 5008 7056
rect 4668 6914 5008 7000
rect 4668 6858 4738 6914
rect 4794 6858 4880 6914
rect 4936 6858 5008 6914
rect 4668 6772 5008 6858
rect 4668 6716 4738 6772
rect 4794 6716 4880 6772
rect 4936 6716 5008 6772
rect 4668 6630 5008 6716
rect 4668 6574 4738 6630
rect 4794 6574 4880 6630
rect 4936 6574 5008 6630
rect 4668 6488 5008 6574
rect 4668 6432 4738 6488
rect 4794 6432 4880 6488
rect 4936 6432 5008 6488
rect 4668 6346 5008 6432
rect 4668 6290 4738 6346
rect 4794 6290 4880 6346
rect 4936 6290 5008 6346
rect 4668 6204 5008 6290
rect 4668 6148 4738 6204
rect 4794 6148 4880 6204
rect 4936 6148 5008 6204
rect 4668 6062 5008 6148
rect 4668 6006 4738 6062
rect 4794 6006 4880 6062
rect 4936 6006 5008 6062
rect 4668 5920 5008 6006
rect 4668 5864 4738 5920
rect 4794 5864 4880 5920
rect 4936 5864 5008 5920
rect 4668 5778 5008 5864
rect 4668 5722 4738 5778
rect 4794 5722 4880 5778
rect 4936 5722 5008 5778
rect 4668 5636 5008 5722
rect 4668 5580 4738 5636
rect 4794 5580 4880 5636
rect 4936 5580 5008 5636
rect 4668 5494 5008 5580
rect 4668 5438 4738 5494
rect 4794 5438 4880 5494
rect 4936 5438 5008 5494
rect 4668 5352 5008 5438
rect 4668 5296 4738 5352
rect 4794 5296 4880 5352
rect 4936 5296 5008 5352
rect 4668 5210 5008 5296
rect 4668 5154 4738 5210
rect 4794 5154 4880 5210
rect 4936 5154 5008 5210
rect 4668 5068 5008 5154
rect 4668 5012 4738 5068
rect 4794 5012 4880 5068
rect 4936 5012 5008 5068
rect 4668 4926 5008 5012
rect 4668 4870 4738 4926
rect 4794 4870 4880 4926
rect 4936 4870 5008 4926
rect 4668 4784 5008 4870
rect 4668 4728 4738 4784
rect 4794 4728 4880 4784
rect 4936 4728 5008 4784
rect 4668 4642 5008 4728
rect 4668 4586 4738 4642
rect 4794 4586 4880 4642
rect 4936 4586 5008 4642
rect 4668 4500 5008 4586
rect 4668 4444 4738 4500
rect 4794 4444 4880 4500
rect 4936 4444 5008 4500
rect 4668 4358 5008 4444
rect 4668 4302 4738 4358
rect 4794 4302 4880 4358
rect 4936 4302 5008 4358
rect 4668 4216 5008 4302
rect 4668 4160 4738 4216
rect 4794 4160 4880 4216
rect 4936 4160 5008 4216
rect 4668 4074 5008 4160
rect 4668 4018 4738 4074
rect 4794 4018 4880 4074
rect 4936 4018 5008 4074
rect 4668 3932 5008 4018
rect 4668 3876 4738 3932
rect 4794 3876 4880 3932
rect 4936 3876 5008 3932
rect 4668 3790 5008 3876
rect 4668 3734 4738 3790
rect 4794 3734 4880 3790
rect 4936 3734 5008 3790
rect 4668 3648 5008 3734
rect 4668 3592 4738 3648
rect 4794 3592 4880 3648
rect 4936 3592 5008 3648
rect 4668 3506 5008 3592
rect 4668 3450 4738 3506
rect 4794 3450 4880 3506
rect 4936 3450 5008 3506
rect 4668 3364 5008 3450
rect 4668 3308 4738 3364
rect 4794 3308 4880 3364
rect 4936 3308 5008 3364
rect 4668 3222 5008 3308
rect 4668 3166 4738 3222
rect 4794 3166 4880 3222
rect 4936 3166 5008 3222
rect 4668 3080 5008 3166
rect 4668 3024 4738 3080
rect 4794 3024 4880 3080
rect 4936 3024 5008 3080
rect 4668 2938 5008 3024
rect 4668 2882 4738 2938
rect 4794 2882 4880 2938
rect 4936 2882 5008 2938
rect 4668 2796 5008 2882
rect 4668 2740 4738 2796
rect 4794 2740 4880 2796
rect 4936 2740 5008 2796
rect 4668 2654 5008 2740
rect 4668 2598 4738 2654
rect 4794 2598 4880 2654
rect 4936 2598 5008 2654
rect 4668 2512 5008 2598
rect 4668 2456 4738 2512
rect 4794 2456 4880 2512
rect 4936 2456 5008 2512
rect 4668 2370 5008 2456
rect 4668 2314 4738 2370
rect 4794 2314 4880 2370
rect 4936 2314 5008 2370
rect 4668 2228 5008 2314
rect 4668 2172 4738 2228
rect 4794 2172 4880 2228
rect 4936 2172 5008 2228
rect 4668 2086 5008 2172
rect 4668 2030 4738 2086
rect 4794 2030 4880 2086
rect 4936 2030 5008 2086
rect 4668 1944 5008 2030
rect 4668 1888 4738 1944
rect 4794 1888 4880 1944
rect 4936 1888 5008 1944
rect 4668 1802 5008 1888
rect 4668 1746 4738 1802
rect 4794 1746 4880 1802
rect 4936 1746 5008 1802
rect 4668 1660 5008 1746
rect 4668 1604 4738 1660
rect 4794 1604 4880 1660
rect 4936 1604 5008 1660
rect 4668 1518 5008 1604
rect 4668 1462 4738 1518
rect 4794 1462 4880 1518
rect 4936 1462 5008 1518
rect 4668 1376 5008 1462
rect 4668 1320 4738 1376
rect 4794 1320 4880 1376
rect 4936 1320 5008 1376
rect 4668 1234 5008 1320
rect 4668 1178 4738 1234
rect 4794 1178 4880 1234
rect 4936 1178 5008 1234
rect 4668 1092 5008 1178
rect 4668 1036 4738 1092
rect 4794 1036 4880 1092
rect 4936 1036 5008 1092
rect 4668 950 5008 1036
rect 4668 894 4738 950
rect 4794 894 4880 950
rect 4936 894 5008 950
rect 4668 808 5008 894
rect 4668 752 4738 808
rect 4794 752 4880 808
rect 4936 752 5008 808
rect 4668 666 5008 752
rect 4668 610 4738 666
rect 4794 610 4880 666
rect 4936 610 5008 666
rect 4668 524 5008 610
rect 4668 468 4738 524
rect 4794 468 4880 524
rect 4936 468 5008 524
rect 4668 400 5008 468
rect 5068 12310 5408 12400
rect 5068 12254 5143 12310
rect 5199 12254 5285 12310
rect 5341 12254 5408 12310
rect 5068 12168 5408 12254
rect 5068 12112 5143 12168
rect 5199 12112 5285 12168
rect 5341 12112 5408 12168
rect 5068 12026 5408 12112
rect 5068 11970 5143 12026
rect 5199 11970 5285 12026
rect 5341 11970 5408 12026
rect 5068 11884 5408 11970
rect 5068 11828 5143 11884
rect 5199 11828 5285 11884
rect 5341 11828 5408 11884
rect 5068 11742 5408 11828
rect 5068 11686 5143 11742
rect 5199 11686 5285 11742
rect 5341 11686 5408 11742
rect 5068 11600 5408 11686
rect 5068 11544 5143 11600
rect 5199 11544 5285 11600
rect 5341 11544 5408 11600
rect 5068 11458 5408 11544
rect 5068 11402 5143 11458
rect 5199 11402 5285 11458
rect 5341 11402 5408 11458
rect 5068 11316 5408 11402
rect 5068 11260 5143 11316
rect 5199 11260 5285 11316
rect 5341 11260 5408 11316
rect 5068 11174 5408 11260
rect 5068 11118 5143 11174
rect 5199 11118 5285 11174
rect 5341 11118 5408 11174
rect 5068 11032 5408 11118
rect 5068 10976 5143 11032
rect 5199 10976 5285 11032
rect 5341 10976 5408 11032
rect 5068 10890 5408 10976
rect 5068 10834 5143 10890
rect 5199 10834 5285 10890
rect 5341 10834 5408 10890
rect 5068 10748 5408 10834
rect 5068 10692 5143 10748
rect 5199 10692 5285 10748
rect 5341 10692 5408 10748
rect 5068 10606 5408 10692
rect 5068 10550 5143 10606
rect 5199 10550 5285 10606
rect 5341 10550 5408 10606
rect 5068 10464 5408 10550
rect 5068 10408 5143 10464
rect 5199 10408 5285 10464
rect 5341 10408 5408 10464
rect 5068 10322 5408 10408
rect 5068 10266 5143 10322
rect 5199 10266 5285 10322
rect 5341 10266 5408 10322
rect 5068 10180 5408 10266
rect 5068 10124 5143 10180
rect 5199 10124 5285 10180
rect 5341 10124 5408 10180
rect 5068 10038 5408 10124
rect 5068 9982 5143 10038
rect 5199 9982 5285 10038
rect 5341 9982 5408 10038
rect 5068 9896 5408 9982
rect 5068 9840 5143 9896
rect 5199 9840 5285 9896
rect 5341 9840 5408 9896
rect 5068 9754 5408 9840
rect 5068 9698 5143 9754
rect 5199 9698 5285 9754
rect 5341 9698 5408 9754
rect 5068 9612 5408 9698
rect 5068 9556 5143 9612
rect 5199 9556 5285 9612
rect 5341 9556 5408 9612
rect 5068 9470 5408 9556
rect 5068 9414 5143 9470
rect 5199 9414 5285 9470
rect 5341 9414 5408 9470
rect 5068 9328 5408 9414
rect 5068 9272 5143 9328
rect 5199 9272 5285 9328
rect 5341 9272 5408 9328
rect 5068 9186 5408 9272
rect 5068 9130 5143 9186
rect 5199 9130 5285 9186
rect 5341 9130 5408 9186
rect 5068 9044 5408 9130
rect 5068 8988 5143 9044
rect 5199 8988 5285 9044
rect 5341 8988 5408 9044
rect 5068 8902 5408 8988
rect 5068 8846 5143 8902
rect 5199 8846 5285 8902
rect 5341 8846 5408 8902
rect 5068 8760 5408 8846
rect 5068 8704 5143 8760
rect 5199 8704 5285 8760
rect 5341 8704 5408 8760
rect 5068 8618 5408 8704
rect 5068 8562 5143 8618
rect 5199 8562 5285 8618
rect 5341 8562 5408 8618
rect 5068 8476 5408 8562
rect 5068 8420 5143 8476
rect 5199 8420 5285 8476
rect 5341 8420 5408 8476
rect 5068 8334 5408 8420
rect 5068 8278 5143 8334
rect 5199 8278 5285 8334
rect 5341 8278 5408 8334
rect 5068 8192 5408 8278
rect 5068 8136 5143 8192
rect 5199 8136 5285 8192
rect 5341 8136 5408 8192
rect 5068 8050 5408 8136
rect 5068 7994 5143 8050
rect 5199 7994 5285 8050
rect 5341 7994 5408 8050
rect 5068 7908 5408 7994
rect 5068 7852 5143 7908
rect 5199 7852 5285 7908
rect 5341 7852 5408 7908
rect 5068 7766 5408 7852
rect 5068 7710 5143 7766
rect 5199 7710 5285 7766
rect 5341 7710 5408 7766
rect 5068 7624 5408 7710
rect 5068 7568 5143 7624
rect 5199 7568 5285 7624
rect 5341 7568 5408 7624
rect 5068 7482 5408 7568
rect 5068 7426 5143 7482
rect 5199 7426 5285 7482
rect 5341 7426 5408 7482
rect 5068 7340 5408 7426
rect 5068 7284 5143 7340
rect 5199 7284 5285 7340
rect 5341 7284 5408 7340
rect 5068 7198 5408 7284
rect 5068 7142 5143 7198
rect 5199 7142 5285 7198
rect 5341 7142 5408 7198
rect 5068 7056 5408 7142
rect 5068 7000 5143 7056
rect 5199 7000 5285 7056
rect 5341 7000 5408 7056
rect 5068 6914 5408 7000
rect 5068 6858 5143 6914
rect 5199 6858 5285 6914
rect 5341 6858 5408 6914
rect 5068 6772 5408 6858
rect 5068 6716 5143 6772
rect 5199 6716 5285 6772
rect 5341 6716 5408 6772
rect 5068 6630 5408 6716
rect 5068 6574 5143 6630
rect 5199 6574 5285 6630
rect 5341 6574 5408 6630
rect 5068 6488 5408 6574
rect 5068 6432 5143 6488
rect 5199 6432 5285 6488
rect 5341 6432 5408 6488
rect 5068 6346 5408 6432
rect 5068 6290 5143 6346
rect 5199 6290 5285 6346
rect 5341 6290 5408 6346
rect 5068 6204 5408 6290
rect 5068 6148 5143 6204
rect 5199 6148 5285 6204
rect 5341 6148 5408 6204
rect 5068 6062 5408 6148
rect 5068 6006 5143 6062
rect 5199 6006 5285 6062
rect 5341 6006 5408 6062
rect 5068 5920 5408 6006
rect 5068 5864 5143 5920
rect 5199 5864 5285 5920
rect 5341 5864 5408 5920
rect 5068 5778 5408 5864
rect 5068 5722 5143 5778
rect 5199 5722 5285 5778
rect 5341 5722 5408 5778
rect 5068 5636 5408 5722
rect 5068 5580 5143 5636
rect 5199 5580 5285 5636
rect 5341 5580 5408 5636
rect 5068 5494 5408 5580
rect 5068 5438 5143 5494
rect 5199 5438 5285 5494
rect 5341 5438 5408 5494
rect 5068 5352 5408 5438
rect 5068 5296 5143 5352
rect 5199 5296 5285 5352
rect 5341 5296 5408 5352
rect 5068 5210 5408 5296
rect 5068 5154 5143 5210
rect 5199 5154 5285 5210
rect 5341 5154 5408 5210
rect 5068 5068 5408 5154
rect 5068 5012 5143 5068
rect 5199 5012 5285 5068
rect 5341 5012 5408 5068
rect 5068 4926 5408 5012
rect 5068 4870 5143 4926
rect 5199 4870 5285 4926
rect 5341 4870 5408 4926
rect 5068 4784 5408 4870
rect 5068 4728 5143 4784
rect 5199 4728 5285 4784
rect 5341 4728 5408 4784
rect 5068 4642 5408 4728
rect 5068 4586 5143 4642
rect 5199 4586 5285 4642
rect 5341 4586 5408 4642
rect 5068 4500 5408 4586
rect 5068 4444 5143 4500
rect 5199 4444 5285 4500
rect 5341 4444 5408 4500
rect 5068 4358 5408 4444
rect 5068 4302 5143 4358
rect 5199 4302 5285 4358
rect 5341 4302 5408 4358
rect 5068 4216 5408 4302
rect 5068 4160 5143 4216
rect 5199 4160 5285 4216
rect 5341 4160 5408 4216
rect 5068 4074 5408 4160
rect 5068 4018 5143 4074
rect 5199 4018 5285 4074
rect 5341 4018 5408 4074
rect 5068 3932 5408 4018
rect 5068 3876 5143 3932
rect 5199 3876 5285 3932
rect 5341 3876 5408 3932
rect 5068 3790 5408 3876
rect 5068 3734 5143 3790
rect 5199 3734 5285 3790
rect 5341 3734 5408 3790
rect 5068 3648 5408 3734
rect 5068 3592 5143 3648
rect 5199 3592 5285 3648
rect 5341 3592 5408 3648
rect 5068 3506 5408 3592
rect 5068 3450 5143 3506
rect 5199 3450 5285 3506
rect 5341 3450 5408 3506
rect 5068 3364 5408 3450
rect 5068 3308 5143 3364
rect 5199 3308 5285 3364
rect 5341 3308 5408 3364
rect 5068 3222 5408 3308
rect 5068 3166 5143 3222
rect 5199 3166 5285 3222
rect 5341 3166 5408 3222
rect 5068 3080 5408 3166
rect 5068 3024 5143 3080
rect 5199 3024 5285 3080
rect 5341 3024 5408 3080
rect 5068 2938 5408 3024
rect 5068 2882 5143 2938
rect 5199 2882 5285 2938
rect 5341 2882 5408 2938
rect 5068 2796 5408 2882
rect 5068 2740 5143 2796
rect 5199 2740 5285 2796
rect 5341 2740 5408 2796
rect 5068 2654 5408 2740
rect 5068 2598 5143 2654
rect 5199 2598 5285 2654
rect 5341 2598 5408 2654
rect 5068 2512 5408 2598
rect 5068 2456 5143 2512
rect 5199 2456 5285 2512
rect 5341 2456 5408 2512
rect 5068 2370 5408 2456
rect 5068 2314 5143 2370
rect 5199 2314 5285 2370
rect 5341 2314 5408 2370
rect 5068 2228 5408 2314
rect 5068 2172 5143 2228
rect 5199 2172 5285 2228
rect 5341 2172 5408 2228
rect 5068 2086 5408 2172
rect 5068 2030 5143 2086
rect 5199 2030 5285 2086
rect 5341 2030 5408 2086
rect 5068 1944 5408 2030
rect 5068 1888 5143 1944
rect 5199 1888 5285 1944
rect 5341 1888 5408 1944
rect 5068 1802 5408 1888
rect 5068 1746 5143 1802
rect 5199 1746 5285 1802
rect 5341 1746 5408 1802
rect 5068 1660 5408 1746
rect 5068 1604 5143 1660
rect 5199 1604 5285 1660
rect 5341 1604 5408 1660
rect 5068 1518 5408 1604
rect 5068 1462 5143 1518
rect 5199 1462 5285 1518
rect 5341 1462 5408 1518
rect 5068 1376 5408 1462
rect 5068 1320 5143 1376
rect 5199 1320 5285 1376
rect 5341 1320 5408 1376
rect 5068 1234 5408 1320
rect 5068 1178 5143 1234
rect 5199 1178 5285 1234
rect 5341 1178 5408 1234
rect 5068 1092 5408 1178
rect 5068 1036 5143 1092
rect 5199 1036 5285 1092
rect 5341 1036 5408 1092
rect 5068 950 5408 1036
rect 5068 894 5143 950
rect 5199 894 5285 950
rect 5341 894 5408 950
rect 5068 808 5408 894
rect 5068 752 5143 808
rect 5199 752 5285 808
rect 5341 752 5408 808
rect 5068 666 5408 752
rect 5068 610 5143 666
rect 5199 610 5285 666
rect 5341 610 5408 666
rect 5068 524 5408 610
rect 5068 468 5143 524
rect 5199 468 5285 524
rect 5341 468 5408 524
rect 5068 400 5408 468
rect 5468 12310 5808 12400
rect 5468 12254 5540 12310
rect 5596 12254 5682 12310
rect 5738 12254 5808 12310
rect 5468 12168 5808 12254
rect 5468 12112 5540 12168
rect 5596 12112 5682 12168
rect 5738 12112 5808 12168
rect 5468 12026 5808 12112
rect 5468 11970 5540 12026
rect 5596 11970 5682 12026
rect 5738 11970 5808 12026
rect 5468 11884 5808 11970
rect 5468 11828 5540 11884
rect 5596 11828 5682 11884
rect 5738 11828 5808 11884
rect 5468 11742 5808 11828
rect 5468 11686 5540 11742
rect 5596 11686 5682 11742
rect 5738 11686 5808 11742
rect 5468 11600 5808 11686
rect 5468 11544 5540 11600
rect 5596 11544 5682 11600
rect 5738 11544 5808 11600
rect 5468 11458 5808 11544
rect 5468 11402 5540 11458
rect 5596 11402 5682 11458
rect 5738 11402 5808 11458
rect 5468 11316 5808 11402
rect 5468 11260 5540 11316
rect 5596 11260 5682 11316
rect 5738 11260 5808 11316
rect 5468 11174 5808 11260
rect 5468 11118 5540 11174
rect 5596 11118 5682 11174
rect 5738 11118 5808 11174
rect 5468 11032 5808 11118
rect 5468 10976 5540 11032
rect 5596 10976 5682 11032
rect 5738 10976 5808 11032
rect 5468 10890 5808 10976
rect 5468 10834 5540 10890
rect 5596 10834 5682 10890
rect 5738 10834 5808 10890
rect 5468 10748 5808 10834
rect 5468 10692 5540 10748
rect 5596 10692 5682 10748
rect 5738 10692 5808 10748
rect 5468 10606 5808 10692
rect 5468 10550 5540 10606
rect 5596 10550 5682 10606
rect 5738 10550 5808 10606
rect 5468 10464 5808 10550
rect 5468 10408 5540 10464
rect 5596 10408 5682 10464
rect 5738 10408 5808 10464
rect 5468 10322 5808 10408
rect 5468 10266 5540 10322
rect 5596 10266 5682 10322
rect 5738 10266 5808 10322
rect 5468 10180 5808 10266
rect 5468 10124 5540 10180
rect 5596 10124 5682 10180
rect 5738 10124 5808 10180
rect 5468 10038 5808 10124
rect 5468 9982 5540 10038
rect 5596 9982 5682 10038
rect 5738 9982 5808 10038
rect 5468 9896 5808 9982
rect 5468 9840 5540 9896
rect 5596 9840 5682 9896
rect 5738 9840 5808 9896
rect 5468 9754 5808 9840
rect 5468 9698 5540 9754
rect 5596 9698 5682 9754
rect 5738 9698 5808 9754
rect 5468 9612 5808 9698
rect 5468 9556 5540 9612
rect 5596 9556 5682 9612
rect 5738 9556 5808 9612
rect 5468 9470 5808 9556
rect 5468 9414 5540 9470
rect 5596 9414 5682 9470
rect 5738 9414 5808 9470
rect 5468 9328 5808 9414
rect 5468 9272 5540 9328
rect 5596 9272 5682 9328
rect 5738 9272 5808 9328
rect 5468 9186 5808 9272
rect 5468 9130 5540 9186
rect 5596 9130 5682 9186
rect 5738 9130 5808 9186
rect 5468 9044 5808 9130
rect 5468 8988 5540 9044
rect 5596 8988 5682 9044
rect 5738 8988 5808 9044
rect 5468 8902 5808 8988
rect 5468 8846 5540 8902
rect 5596 8846 5682 8902
rect 5738 8846 5808 8902
rect 5468 8760 5808 8846
rect 5468 8704 5540 8760
rect 5596 8704 5682 8760
rect 5738 8704 5808 8760
rect 5468 8618 5808 8704
rect 5468 8562 5540 8618
rect 5596 8562 5682 8618
rect 5738 8562 5808 8618
rect 5468 8476 5808 8562
rect 5468 8420 5540 8476
rect 5596 8420 5682 8476
rect 5738 8420 5808 8476
rect 5468 8334 5808 8420
rect 5468 8278 5540 8334
rect 5596 8278 5682 8334
rect 5738 8278 5808 8334
rect 5468 8192 5808 8278
rect 5468 8136 5540 8192
rect 5596 8136 5682 8192
rect 5738 8136 5808 8192
rect 5468 8050 5808 8136
rect 5468 7994 5540 8050
rect 5596 7994 5682 8050
rect 5738 7994 5808 8050
rect 5468 7908 5808 7994
rect 5468 7852 5540 7908
rect 5596 7852 5682 7908
rect 5738 7852 5808 7908
rect 5468 7766 5808 7852
rect 5468 7710 5540 7766
rect 5596 7710 5682 7766
rect 5738 7710 5808 7766
rect 5468 7624 5808 7710
rect 5468 7568 5540 7624
rect 5596 7568 5682 7624
rect 5738 7568 5808 7624
rect 5468 7482 5808 7568
rect 5468 7426 5540 7482
rect 5596 7426 5682 7482
rect 5738 7426 5808 7482
rect 5468 7340 5808 7426
rect 5468 7284 5540 7340
rect 5596 7284 5682 7340
rect 5738 7284 5808 7340
rect 5468 7198 5808 7284
rect 5468 7142 5540 7198
rect 5596 7142 5682 7198
rect 5738 7142 5808 7198
rect 5468 7056 5808 7142
rect 5468 7000 5540 7056
rect 5596 7000 5682 7056
rect 5738 7000 5808 7056
rect 5468 6914 5808 7000
rect 5468 6858 5540 6914
rect 5596 6858 5682 6914
rect 5738 6858 5808 6914
rect 5468 6772 5808 6858
rect 5468 6716 5540 6772
rect 5596 6716 5682 6772
rect 5738 6716 5808 6772
rect 5468 6630 5808 6716
rect 5468 6574 5540 6630
rect 5596 6574 5682 6630
rect 5738 6574 5808 6630
rect 5468 6488 5808 6574
rect 5468 6432 5540 6488
rect 5596 6432 5682 6488
rect 5738 6432 5808 6488
rect 5468 6346 5808 6432
rect 5468 6290 5540 6346
rect 5596 6290 5682 6346
rect 5738 6290 5808 6346
rect 5468 6204 5808 6290
rect 5468 6148 5540 6204
rect 5596 6148 5682 6204
rect 5738 6148 5808 6204
rect 5468 6062 5808 6148
rect 5468 6006 5540 6062
rect 5596 6006 5682 6062
rect 5738 6006 5808 6062
rect 5468 5920 5808 6006
rect 5468 5864 5540 5920
rect 5596 5864 5682 5920
rect 5738 5864 5808 5920
rect 5468 5778 5808 5864
rect 5468 5722 5540 5778
rect 5596 5722 5682 5778
rect 5738 5722 5808 5778
rect 5468 5636 5808 5722
rect 5468 5580 5540 5636
rect 5596 5580 5682 5636
rect 5738 5580 5808 5636
rect 5468 5494 5808 5580
rect 5468 5438 5540 5494
rect 5596 5438 5682 5494
rect 5738 5438 5808 5494
rect 5468 5352 5808 5438
rect 5468 5296 5540 5352
rect 5596 5296 5682 5352
rect 5738 5296 5808 5352
rect 5468 5210 5808 5296
rect 5468 5154 5540 5210
rect 5596 5154 5682 5210
rect 5738 5154 5808 5210
rect 5468 5068 5808 5154
rect 5468 5012 5540 5068
rect 5596 5012 5682 5068
rect 5738 5012 5808 5068
rect 5468 4926 5808 5012
rect 5468 4870 5540 4926
rect 5596 4870 5682 4926
rect 5738 4870 5808 4926
rect 5468 4784 5808 4870
rect 5468 4728 5540 4784
rect 5596 4728 5682 4784
rect 5738 4728 5808 4784
rect 5468 4642 5808 4728
rect 5468 4586 5540 4642
rect 5596 4586 5682 4642
rect 5738 4586 5808 4642
rect 5468 4500 5808 4586
rect 5468 4444 5540 4500
rect 5596 4444 5682 4500
rect 5738 4444 5808 4500
rect 5468 4358 5808 4444
rect 5468 4302 5540 4358
rect 5596 4302 5682 4358
rect 5738 4302 5808 4358
rect 5468 4216 5808 4302
rect 5468 4160 5540 4216
rect 5596 4160 5682 4216
rect 5738 4160 5808 4216
rect 5468 4074 5808 4160
rect 5468 4018 5540 4074
rect 5596 4018 5682 4074
rect 5738 4018 5808 4074
rect 5468 3932 5808 4018
rect 5468 3876 5540 3932
rect 5596 3876 5682 3932
rect 5738 3876 5808 3932
rect 5468 3790 5808 3876
rect 5468 3734 5540 3790
rect 5596 3734 5682 3790
rect 5738 3734 5808 3790
rect 5468 3648 5808 3734
rect 5468 3592 5540 3648
rect 5596 3592 5682 3648
rect 5738 3592 5808 3648
rect 5468 3506 5808 3592
rect 5468 3450 5540 3506
rect 5596 3450 5682 3506
rect 5738 3450 5808 3506
rect 5468 3364 5808 3450
rect 5468 3308 5540 3364
rect 5596 3308 5682 3364
rect 5738 3308 5808 3364
rect 5468 3222 5808 3308
rect 5468 3166 5540 3222
rect 5596 3166 5682 3222
rect 5738 3166 5808 3222
rect 5468 3080 5808 3166
rect 5468 3024 5540 3080
rect 5596 3024 5682 3080
rect 5738 3024 5808 3080
rect 5468 2938 5808 3024
rect 5468 2882 5540 2938
rect 5596 2882 5682 2938
rect 5738 2882 5808 2938
rect 5468 2796 5808 2882
rect 5468 2740 5540 2796
rect 5596 2740 5682 2796
rect 5738 2740 5808 2796
rect 5468 2654 5808 2740
rect 5468 2598 5540 2654
rect 5596 2598 5682 2654
rect 5738 2598 5808 2654
rect 5468 2512 5808 2598
rect 5468 2456 5540 2512
rect 5596 2456 5682 2512
rect 5738 2456 5808 2512
rect 5468 2370 5808 2456
rect 5468 2314 5540 2370
rect 5596 2314 5682 2370
rect 5738 2314 5808 2370
rect 5468 2228 5808 2314
rect 5468 2172 5540 2228
rect 5596 2172 5682 2228
rect 5738 2172 5808 2228
rect 5468 2086 5808 2172
rect 5468 2030 5540 2086
rect 5596 2030 5682 2086
rect 5738 2030 5808 2086
rect 5468 1944 5808 2030
rect 5468 1888 5540 1944
rect 5596 1888 5682 1944
rect 5738 1888 5808 1944
rect 5468 1802 5808 1888
rect 5468 1746 5540 1802
rect 5596 1746 5682 1802
rect 5738 1746 5808 1802
rect 5468 1660 5808 1746
rect 5468 1604 5540 1660
rect 5596 1604 5682 1660
rect 5738 1604 5808 1660
rect 5468 1518 5808 1604
rect 5468 1462 5540 1518
rect 5596 1462 5682 1518
rect 5738 1462 5808 1518
rect 5468 1376 5808 1462
rect 5468 1320 5540 1376
rect 5596 1320 5682 1376
rect 5738 1320 5808 1376
rect 5468 1234 5808 1320
rect 5468 1178 5540 1234
rect 5596 1178 5682 1234
rect 5738 1178 5808 1234
rect 5468 1092 5808 1178
rect 5468 1036 5540 1092
rect 5596 1036 5682 1092
rect 5738 1036 5808 1092
rect 5468 950 5808 1036
rect 5468 894 5540 950
rect 5596 894 5682 950
rect 5738 894 5808 950
rect 5468 808 5808 894
rect 5468 752 5540 808
rect 5596 752 5682 808
rect 5738 752 5808 808
rect 5468 666 5808 752
rect 5468 610 5540 666
rect 5596 610 5682 666
rect 5738 610 5808 666
rect 5468 524 5808 610
rect 5468 468 5540 524
rect 5596 468 5682 524
rect 5738 468 5808 524
rect 5468 400 5808 468
rect 5868 12310 6208 12400
rect 5868 12254 5937 12310
rect 5993 12254 6079 12310
rect 6135 12254 6208 12310
rect 5868 12168 6208 12254
rect 5868 12112 5937 12168
rect 5993 12112 6079 12168
rect 6135 12112 6208 12168
rect 5868 12026 6208 12112
rect 5868 11970 5937 12026
rect 5993 11970 6079 12026
rect 6135 11970 6208 12026
rect 5868 11884 6208 11970
rect 5868 11828 5937 11884
rect 5993 11828 6079 11884
rect 6135 11828 6208 11884
rect 5868 11742 6208 11828
rect 5868 11686 5937 11742
rect 5993 11686 6079 11742
rect 6135 11686 6208 11742
rect 5868 11600 6208 11686
rect 5868 11544 5937 11600
rect 5993 11544 6079 11600
rect 6135 11544 6208 11600
rect 5868 11458 6208 11544
rect 5868 11402 5937 11458
rect 5993 11402 6079 11458
rect 6135 11402 6208 11458
rect 5868 11316 6208 11402
rect 5868 11260 5937 11316
rect 5993 11260 6079 11316
rect 6135 11260 6208 11316
rect 5868 11174 6208 11260
rect 5868 11118 5937 11174
rect 5993 11118 6079 11174
rect 6135 11118 6208 11174
rect 5868 11032 6208 11118
rect 5868 10976 5937 11032
rect 5993 10976 6079 11032
rect 6135 10976 6208 11032
rect 5868 10890 6208 10976
rect 5868 10834 5937 10890
rect 5993 10834 6079 10890
rect 6135 10834 6208 10890
rect 5868 10748 6208 10834
rect 5868 10692 5937 10748
rect 5993 10692 6079 10748
rect 6135 10692 6208 10748
rect 5868 10606 6208 10692
rect 5868 10550 5937 10606
rect 5993 10550 6079 10606
rect 6135 10550 6208 10606
rect 5868 10464 6208 10550
rect 5868 10408 5937 10464
rect 5993 10408 6079 10464
rect 6135 10408 6208 10464
rect 5868 10322 6208 10408
rect 5868 10266 5937 10322
rect 5993 10266 6079 10322
rect 6135 10266 6208 10322
rect 5868 10180 6208 10266
rect 5868 10124 5937 10180
rect 5993 10124 6079 10180
rect 6135 10124 6208 10180
rect 5868 10038 6208 10124
rect 5868 9982 5937 10038
rect 5993 9982 6079 10038
rect 6135 9982 6208 10038
rect 5868 9896 6208 9982
rect 5868 9840 5937 9896
rect 5993 9840 6079 9896
rect 6135 9840 6208 9896
rect 5868 9754 6208 9840
rect 5868 9698 5937 9754
rect 5993 9698 6079 9754
rect 6135 9698 6208 9754
rect 5868 9612 6208 9698
rect 5868 9556 5937 9612
rect 5993 9556 6079 9612
rect 6135 9556 6208 9612
rect 5868 9470 6208 9556
rect 5868 9414 5937 9470
rect 5993 9414 6079 9470
rect 6135 9414 6208 9470
rect 5868 9328 6208 9414
rect 5868 9272 5937 9328
rect 5993 9272 6079 9328
rect 6135 9272 6208 9328
rect 5868 9186 6208 9272
rect 5868 9130 5937 9186
rect 5993 9130 6079 9186
rect 6135 9130 6208 9186
rect 5868 9044 6208 9130
rect 5868 8988 5937 9044
rect 5993 8988 6079 9044
rect 6135 8988 6208 9044
rect 5868 8902 6208 8988
rect 5868 8846 5937 8902
rect 5993 8846 6079 8902
rect 6135 8846 6208 8902
rect 5868 8760 6208 8846
rect 5868 8704 5937 8760
rect 5993 8704 6079 8760
rect 6135 8704 6208 8760
rect 5868 8618 6208 8704
rect 5868 8562 5937 8618
rect 5993 8562 6079 8618
rect 6135 8562 6208 8618
rect 5868 8476 6208 8562
rect 5868 8420 5937 8476
rect 5993 8420 6079 8476
rect 6135 8420 6208 8476
rect 5868 8334 6208 8420
rect 5868 8278 5937 8334
rect 5993 8278 6079 8334
rect 6135 8278 6208 8334
rect 5868 8192 6208 8278
rect 5868 8136 5937 8192
rect 5993 8136 6079 8192
rect 6135 8136 6208 8192
rect 5868 8050 6208 8136
rect 5868 7994 5937 8050
rect 5993 7994 6079 8050
rect 6135 7994 6208 8050
rect 5868 7908 6208 7994
rect 5868 7852 5937 7908
rect 5993 7852 6079 7908
rect 6135 7852 6208 7908
rect 5868 7766 6208 7852
rect 5868 7710 5937 7766
rect 5993 7710 6079 7766
rect 6135 7710 6208 7766
rect 5868 7624 6208 7710
rect 5868 7568 5937 7624
rect 5993 7568 6079 7624
rect 6135 7568 6208 7624
rect 5868 7482 6208 7568
rect 5868 7426 5937 7482
rect 5993 7426 6079 7482
rect 6135 7426 6208 7482
rect 5868 7340 6208 7426
rect 5868 7284 5937 7340
rect 5993 7284 6079 7340
rect 6135 7284 6208 7340
rect 5868 7198 6208 7284
rect 5868 7142 5937 7198
rect 5993 7142 6079 7198
rect 6135 7142 6208 7198
rect 5868 7056 6208 7142
rect 5868 7000 5937 7056
rect 5993 7000 6079 7056
rect 6135 7000 6208 7056
rect 5868 6914 6208 7000
rect 5868 6858 5937 6914
rect 5993 6858 6079 6914
rect 6135 6858 6208 6914
rect 5868 6772 6208 6858
rect 5868 6716 5937 6772
rect 5993 6716 6079 6772
rect 6135 6716 6208 6772
rect 5868 6630 6208 6716
rect 5868 6574 5937 6630
rect 5993 6574 6079 6630
rect 6135 6574 6208 6630
rect 5868 6488 6208 6574
rect 5868 6432 5937 6488
rect 5993 6432 6079 6488
rect 6135 6432 6208 6488
rect 5868 6346 6208 6432
rect 5868 6290 5937 6346
rect 5993 6290 6079 6346
rect 6135 6290 6208 6346
rect 5868 6204 6208 6290
rect 5868 6148 5937 6204
rect 5993 6148 6079 6204
rect 6135 6148 6208 6204
rect 5868 6062 6208 6148
rect 5868 6006 5937 6062
rect 5993 6006 6079 6062
rect 6135 6006 6208 6062
rect 5868 5920 6208 6006
rect 5868 5864 5937 5920
rect 5993 5864 6079 5920
rect 6135 5864 6208 5920
rect 5868 5778 6208 5864
rect 5868 5722 5937 5778
rect 5993 5722 6079 5778
rect 6135 5722 6208 5778
rect 5868 5636 6208 5722
rect 5868 5580 5937 5636
rect 5993 5580 6079 5636
rect 6135 5580 6208 5636
rect 5868 5494 6208 5580
rect 5868 5438 5937 5494
rect 5993 5438 6079 5494
rect 6135 5438 6208 5494
rect 5868 5352 6208 5438
rect 5868 5296 5937 5352
rect 5993 5296 6079 5352
rect 6135 5296 6208 5352
rect 5868 5210 6208 5296
rect 5868 5154 5937 5210
rect 5993 5154 6079 5210
rect 6135 5154 6208 5210
rect 5868 5068 6208 5154
rect 5868 5012 5937 5068
rect 5993 5012 6079 5068
rect 6135 5012 6208 5068
rect 5868 4926 6208 5012
rect 5868 4870 5937 4926
rect 5993 4870 6079 4926
rect 6135 4870 6208 4926
rect 5868 4784 6208 4870
rect 5868 4728 5937 4784
rect 5993 4728 6079 4784
rect 6135 4728 6208 4784
rect 5868 4642 6208 4728
rect 5868 4586 5937 4642
rect 5993 4586 6079 4642
rect 6135 4586 6208 4642
rect 5868 4500 6208 4586
rect 5868 4444 5937 4500
rect 5993 4444 6079 4500
rect 6135 4444 6208 4500
rect 5868 4358 6208 4444
rect 5868 4302 5937 4358
rect 5993 4302 6079 4358
rect 6135 4302 6208 4358
rect 5868 4216 6208 4302
rect 5868 4160 5937 4216
rect 5993 4160 6079 4216
rect 6135 4160 6208 4216
rect 5868 4074 6208 4160
rect 5868 4018 5937 4074
rect 5993 4018 6079 4074
rect 6135 4018 6208 4074
rect 5868 3932 6208 4018
rect 5868 3876 5937 3932
rect 5993 3876 6079 3932
rect 6135 3876 6208 3932
rect 5868 3790 6208 3876
rect 5868 3734 5937 3790
rect 5993 3734 6079 3790
rect 6135 3734 6208 3790
rect 5868 3648 6208 3734
rect 5868 3592 5937 3648
rect 5993 3592 6079 3648
rect 6135 3592 6208 3648
rect 5868 3506 6208 3592
rect 5868 3450 5937 3506
rect 5993 3450 6079 3506
rect 6135 3450 6208 3506
rect 5868 3364 6208 3450
rect 5868 3308 5937 3364
rect 5993 3308 6079 3364
rect 6135 3308 6208 3364
rect 5868 3222 6208 3308
rect 5868 3166 5937 3222
rect 5993 3166 6079 3222
rect 6135 3166 6208 3222
rect 5868 3080 6208 3166
rect 5868 3024 5937 3080
rect 5993 3024 6079 3080
rect 6135 3024 6208 3080
rect 5868 2938 6208 3024
rect 5868 2882 5937 2938
rect 5993 2882 6079 2938
rect 6135 2882 6208 2938
rect 5868 2796 6208 2882
rect 5868 2740 5937 2796
rect 5993 2740 6079 2796
rect 6135 2740 6208 2796
rect 5868 2654 6208 2740
rect 5868 2598 5937 2654
rect 5993 2598 6079 2654
rect 6135 2598 6208 2654
rect 5868 2512 6208 2598
rect 5868 2456 5937 2512
rect 5993 2456 6079 2512
rect 6135 2456 6208 2512
rect 5868 2370 6208 2456
rect 5868 2314 5937 2370
rect 5993 2314 6079 2370
rect 6135 2314 6208 2370
rect 5868 2228 6208 2314
rect 5868 2172 5937 2228
rect 5993 2172 6079 2228
rect 6135 2172 6208 2228
rect 5868 2086 6208 2172
rect 5868 2030 5937 2086
rect 5993 2030 6079 2086
rect 6135 2030 6208 2086
rect 5868 1944 6208 2030
rect 5868 1888 5937 1944
rect 5993 1888 6079 1944
rect 6135 1888 6208 1944
rect 5868 1802 6208 1888
rect 5868 1746 5937 1802
rect 5993 1746 6079 1802
rect 6135 1746 6208 1802
rect 5868 1660 6208 1746
rect 5868 1604 5937 1660
rect 5993 1604 6079 1660
rect 6135 1604 6208 1660
rect 5868 1518 6208 1604
rect 5868 1462 5937 1518
rect 5993 1462 6079 1518
rect 6135 1462 6208 1518
rect 5868 1376 6208 1462
rect 5868 1320 5937 1376
rect 5993 1320 6079 1376
rect 6135 1320 6208 1376
rect 5868 1234 6208 1320
rect 5868 1178 5937 1234
rect 5993 1178 6079 1234
rect 6135 1178 6208 1234
rect 5868 1092 6208 1178
rect 5868 1036 5937 1092
rect 5993 1036 6079 1092
rect 6135 1036 6208 1092
rect 5868 950 6208 1036
rect 5868 894 5937 950
rect 5993 894 6079 950
rect 6135 894 6208 950
rect 5868 808 6208 894
rect 5868 752 5937 808
rect 5993 752 6079 808
rect 6135 752 6208 808
rect 5868 666 6208 752
rect 5868 610 5937 666
rect 5993 610 6079 666
rect 6135 610 6208 666
rect 5868 524 6208 610
rect 5868 468 5937 524
rect 5993 468 6079 524
rect 6135 468 6208 524
rect 5868 400 6208 468
rect 6268 12310 6608 12400
rect 6268 12254 6340 12310
rect 6396 12254 6482 12310
rect 6538 12254 6608 12310
rect 6268 12168 6608 12254
rect 6268 12112 6340 12168
rect 6396 12112 6482 12168
rect 6538 12112 6608 12168
rect 6268 12026 6608 12112
rect 6268 11970 6340 12026
rect 6396 11970 6482 12026
rect 6538 11970 6608 12026
rect 6268 11884 6608 11970
rect 6268 11828 6340 11884
rect 6396 11828 6482 11884
rect 6538 11828 6608 11884
rect 6268 11742 6608 11828
rect 6268 11686 6340 11742
rect 6396 11686 6482 11742
rect 6538 11686 6608 11742
rect 6268 11600 6608 11686
rect 6268 11544 6340 11600
rect 6396 11544 6482 11600
rect 6538 11544 6608 11600
rect 6268 11458 6608 11544
rect 6268 11402 6340 11458
rect 6396 11402 6482 11458
rect 6538 11402 6608 11458
rect 6268 11316 6608 11402
rect 6268 11260 6340 11316
rect 6396 11260 6482 11316
rect 6538 11260 6608 11316
rect 6268 11174 6608 11260
rect 6268 11118 6340 11174
rect 6396 11118 6482 11174
rect 6538 11118 6608 11174
rect 6268 11032 6608 11118
rect 6268 10976 6340 11032
rect 6396 10976 6482 11032
rect 6538 10976 6608 11032
rect 6268 10890 6608 10976
rect 6268 10834 6340 10890
rect 6396 10834 6482 10890
rect 6538 10834 6608 10890
rect 6268 10748 6608 10834
rect 6268 10692 6340 10748
rect 6396 10692 6482 10748
rect 6538 10692 6608 10748
rect 6268 10606 6608 10692
rect 6268 10550 6340 10606
rect 6396 10550 6482 10606
rect 6538 10550 6608 10606
rect 6268 10464 6608 10550
rect 6268 10408 6340 10464
rect 6396 10408 6482 10464
rect 6538 10408 6608 10464
rect 6268 10322 6608 10408
rect 6268 10266 6340 10322
rect 6396 10266 6482 10322
rect 6538 10266 6608 10322
rect 6268 10180 6608 10266
rect 6268 10124 6340 10180
rect 6396 10124 6482 10180
rect 6538 10124 6608 10180
rect 6268 10038 6608 10124
rect 6268 9982 6340 10038
rect 6396 9982 6482 10038
rect 6538 9982 6608 10038
rect 6268 9896 6608 9982
rect 6268 9840 6340 9896
rect 6396 9840 6482 9896
rect 6538 9840 6608 9896
rect 6268 9754 6608 9840
rect 6268 9698 6340 9754
rect 6396 9698 6482 9754
rect 6538 9698 6608 9754
rect 6268 9612 6608 9698
rect 6268 9556 6340 9612
rect 6396 9556 6482 9612
rect 6538 9556 6608 9612
rect 6268 9470 6608 9556
rect 6268 9414 6340 9470
rect 6396 9414 6482 9470
rect 6538 9414 6608 9470
rect 6268 9328 6608 9414
rect 6268 9272 6340 9328
rect 6396 9272 6482 9328
rect 6538 9272 6608 9328
rect 6268 9186 6608 9272
rect 6268 9130 6340 9186
rect 6396 9130 6482 9186
rect 6538 9130 6608 9186
rect 6268 9044 6608 9130
rect 6268 8988 6340 9044
rect 6396 8988 6482 9044
rect 6538 8988 6608 9044
rect 6268 8902 6608 8988
rect 6268 8846 6340 8902
rect 6396 8846 6482 8902
rect 6538 8846 6608 8902
rect 6268 8760 6608 8846
rect 6268 8704 6340 8760
rect 6396 8704 6482 8760
rect 6538 8704 6608 8760
rect 6268 8618 6608 8704
rect 6268 8562 6340 8618
rect 6396 8562 6482 8618
rect 6538 8562 6608 8618
rect 6268 8476 6608 8562
rect 6268 8420 6340 8476
rect 6396 8420 6482 8476
rect 6538 8420 6608 8476
rect 6268 8334 6608 8420
rect 6268 8278 6340 8334
rect 6396 8278 6482 8334
rect 6538 8278 6608 8334
rect 6268 8192 6608 8278
rect 6268 8136 6340 8192
rect 6396 8136 6482 8192
rect 6538 8136 6608 8192
rect 6268 8050 6608 8136
rect 6268 7994 6340 8050
rect 6396 7994 6482 8050
rect 6538 7994 6608 8050
rect 6268 7908 6608 7994
rect 6268 7852 6340 7908
rect 6396 7852 6482 7908
rect 6538 7852 6608 7908
rect 6268 7766 6608 7852
rect 6268 7710 6340 7766
rect 6396 7710 6482 7766
rect 6538 7710 6608 7766
rect 6268 7624 6608 7710
rect 6268 7568 6340 7624
rect 6396 7568 6482 7624
rect 6538 7568 6608 7624
rect 6268 7482 6608 7568
rect 6268 7426 6340 7482
rect 6396 7426 6482 7482
rect 6538 7426 6608 7482
rect 6268 7340 6608 7426
rect 6268 7284 6340 7340
rect 6396 7284 6482 7340
rect 6538 7284 6608 7340
rect 6268 7198 6608 7284
rect 6268 7142 6340 7198
rect 6396 7142 6482 7198
rect 6538 7142 6608 7198
rect 6268 7056 6608 7142
rect 6268 7000 6340 7056
rect 6396 7000 6482 7056
rect 6538 7000 6608 7056
rect 6268 6914 6608 7000
rect 6268 6858 6340 6914
rect 6396 6858 6482 6914
rect 6538 6858 6608 6914
rect 6268 6772 6608 6858
rect 6268 6716 6340 6772
rect 6396 6716 6482 6772
rect 6538 6716 6608 6772
rect 6268 6630 6608 6716
rect 6268 6574 6340 6630
rect 6396 6574 6482 6630
rect 6538 6574 6608 6630
rect 6268 6488 6608 6574
rect 6268 6432 6340 6488
rect 6396 6432 6482 6488
rect 6538 6432 6608 6488
rect 6268 6346 6608 6432
rect 6268 6290 6340 6346
rect 6396 6290 6482 6346
rect 6538 6290 6608 6346
rect 6268 6204 6608 6290
rect 6268 6148 6340 6204
rect 6396 6148 6482 6204
rect 6538 6148 6608 6204
rect 6268 6062 6608 6148
rect 6268 6006 6340 6062
rect 6396 6006 6482 6062
rect 6538 6006 6608 6062
rect 6268 5920 6608 6006
rect 6268 5864 6340 5920
rect 6396 5864 6482 5920
rect 6538 5864 6608 5920
rect 6268 5778 6608 5864
rect 6268 5722 6340 5778
rect 6396 5722 6482 5778
rect 6538 5722 6608 5778
rect 6268 5636 6608 5722
rect 6268 5580 6340 5636
rect 6396 5580 6482 5636
rect 6538 5580 6608 5636
rect 6268 5494 6608 5580
rect 6268 5438 6340 5494
rect 6396 5438 6482 5494
rect 6538 5438 6608 5494
rect 6268 5352 6608 5438
rect 6268 5296 6340 5352
rect 6396 5296 6482 5352
rect 6538 5296 6608 5352
rect 6268 5210 6608 5296
rect 6268 5154 6340 5210
rect 6396 5154 6482 5210
rect 6538 5154 6608 5210
rect 6268 5068 6608 5154
rect 6268 5012 6340 5068
rect 6396 5012 6482 5068
rect 6538 5012 6608 5068
rect 6268 4926 6608 5012
rect 6268 4870 6340 4926
rect 6396 4870 6482 4926
rect 6538 4870 6608 4926
rect 6268 4784 6608 4870
rect 6268 4728 6340 4784
rect 6396 4728 6482 4784
rect 6538 4728 6608 4784
rect 6268 4642 6608 4728
rect 6268 4586 6340 4642
rect 6396 4586 6482 4642
rect 6538 4586 6608 4642
rect 6268 4500 6608 4586
rect 6268 4444 6340 4500
rect 6396 4444 6482 4500
rect 6538 4444 6608 4500
rect 6268 4358 6608 4444
rect 6268 4302 6340 4358
rect 6396 4302 6482 4358
rect 6538 4302 6608 4358
rect 6268 4216 6608 4302
rect 6268 4160 6340 4216
rect 6396 4160 6482 4216
rect 6538 4160 6608 4216
rect 6268 4074 6608 4160
rect 6268 4018 6340 4074
rect 6396 4018 6482 4074
rect 6538 4018 6608 4074
rect 6268 3932 6608 4018
rect 6268 3876 6340 3932
rect 6396 3876 6482 3932
rect 6538 3876 6608 3932
rect 6268 3790 6608 3876
rect 6268 3734 6340 3790
rect 6396 3734 6482 3790
rect 6538 3734 6608 3790
rect 6268 3648 6608 3734
rect 6268 3592 6340 3648
rect 6396 3592 6482 3648
rect 6538 3592 6608 3648
rect 6268 3506 6608 3592
rect 6268 3450 6340 3506
rect 6396 3450 6482 3506
rect 6538 3450 6608 3506
rect 6268 3364 6608 3450
rect 6268 3308 6340 3364
rect 6396 3308 6482 3364
rect 6538 3308 6608 3364
rect 6268 3222 6608 3308
rect 6268 3166 6340 3222
rect 6396 3166 6482 3222
rect 6538 3166 6608 3222
rect 6268 3080 6608 3166
rect 6268 3024 6340 3080
rect 6396 3024 6482 3080
rect 6538 3024 6608 3080
rect 6268 2938 6608 3024
rect 6268 2882 6340 2938
rect 6396 2882 6482 2938
rect 6538 2882 6608 2938
rect 6268 2796 6608 2882
rect 6268 2740 6340 2796
rect 6396 2740 6482 2796
rect 6538 2740 6608 2796
rect 6268 2654 6608 2740
rect 6268 2598 6340 2654
rect 6396 2598 6482 2654
rect 6538 2598 6608 2654
rect 6268 2512 6608 2598
rect 6268 2456 6340 2512
rect 6396 2456 6482 2512
rect 6538 2456 6608 2512
rect 6268 2370 6608 2456
rect 6268 2314 6340 2370
rect 6396 2314 6482 2370
rect 6538 2314 6608 2370
rect 6268 2228 6608 2314
rect 6268 2172 6340 2228
rect 6396 2172 6482 2228
rect 6538 2172 6608 2228
rect 6268 2086 6608 2172
rect 6268 2030 6340 2086
rect 6396 2030 6482 2086
rect 6538 2030 6608 2086
rect 6268 1944 6608 2030
rect 6268 1888 6340 1944
rect 6396 1888 6482 1944
rect 6538 1888 6608 1944
rect 6268 1802 6608 1888
rect 6268 1746 6340 1802
rect 6396 1746 6482 1802
rect 6538 1746 6608 1802
rect 6268 1660 6608 1746
rect 6268 1604 6340 1660
rect 6396 1604 6482 1660
rect 6538 1604 6608 1660
rect 6268 1518 6608 1604
rect 6268 1462 6340 1518
rect 6396 1462 6482 1518
rect 6538 1462 6608 1518
rect 6268 1376 6608 1462
rect 6268 1320 6340 1376
rect 6396 1320 6482 1376
rect 6538 1320 6608 1376
rect 6268 1234 6608 1320
rect 6268 1178 6340 1234
rect 6396 1178 6482 1234
rect 6538 1178 6608 1234
rect 6268 1092 6608 1178
rect 6268 1036 6340 1092
rect 6396 1036 6482 1092
rect 6538 1036 6608 1092
rect 6268 950 6608 1036
rect 6268 894 6340 950
rect 6396 894 6482 950
rect 6538 894 6608 950
rect 6268 808 6608 894
rect 6268 752 6340 808
rect 6396 752 6482 808
rect 6538 752 6608 808
rect 6268 666 6608 752
rect 6268 610 6340 666
rect 6396 610 6482 666
rect 6538 610 6608 666
rect 6268 524 6608 610
rect 6268 468 6340 524
rect 6396 468 6482 524
rect 6538 468 6608 524
rect 6268 400 6608 468
rect 6668 12310 7008 12400
rect 6668 12254 6742 12310
rect 6798 12254 6884 12310
rect 6940 12254 7008 12310
rect 6668 12168 7008 12254
rect 6668 12112 6742 12168
rect 6798 12112 6884 12168
rect 6940 12112 7008 12168
rect 6668 12026 7008 12112
rect 6668 11970 6742 12026
rect 6798 11970 6884 12026
rect 6940 11970 7008 12026
rect 6668 11884 7008 11970
rect 6668 11828 6742 11884
rect 6798 11828 6884 11884
rect 6940 11828 7008 11884
rect 6668 11742 7008 11828
rect 6668 11686 6742 11742
rect 6798 11686 6884 11742
rect 6940 11686 7008 11742
rect 6668 11600 7008 11686
rect 6668 11544 6742 11600
rect 6798 11544 6884 11600
rect 6940 11544 7008 11600
rect 6668 11458 7008 11544
rect 6668 11402 6742 11458
rect 6798 11402 6884 11458
rect 6940 11402 7008 11458
rect 6668 11316 7008 11402
rect 6668 11260 6742 11316
rect 6798 11260 6884 11316
rect 6940 11260 7008 11316
rect 6668 11174 7008 11260
rect 6668 11118 6742 11174
rect 6798 11118 6884 11174
rect 6940 11118 7008 11174
rect 6668 11032 7008 11118
rect 6668 10976 6742 11032
rect 6798 10976 6884 11032
rect 6940 10976 7008 11032
rect 6668 10890 7008 10976
rect 6668 10834 6742 10890
rect 6798 10834 6884 10890
rect 6940 10834 7008 10890
rect 6668 10748 7008 10834
rect 6668 10692 6742 10748
rect 6798 10692 6884 10748
rect 6940 10692 7008 10748
rect 6668 10606 7008 10692
rect 6668 10550 6742 10606
rect 6798 10550 6884 10606
rect 6940 10550 7008 10606
rect 6668 10464 7008 10550
rect 6668 10408 6742 10464
rect 6798 10408 6884 10464
rect 6940 10408 7008 10464
rect 6668 10322 7008 10408
rect 6668 10266 6742 10322
rect 6798 10266 6884 10322
rect 6940 10266 7008 10322
rect 6668 10180 7008 10266
rect 6668 10124 6742 10180
rect 6798 10124 6884 10180
rect 6940 10124 7008 10180
rect 6668 10038 7008 10124
rect 6668 9982 6742 10038
rect 6798 9982 6884 10038
rect 6940 9982 7008 10038
rect 6668 9896 7008 9982
rect 6668 9840 6742 9896
rect 6798 9840 6884 9896
rect 6940 9840 7008 9896
rect 6668 9754 7008 9840
rect 6668 9698 6742 9754
rect 6798 9698 6884 9754
rect 6940 9698 7008 9754
rect 6668 9612 7008 9698
rect 6668 9556 6742 9612
rect 6798 9556 6884 9612
rect 6940 9556 7008 9612
rect 6668 9470 7008 9556
rect 6668 9414 6742 9470
rect 6798 9414 6884 9470
rect 6940 9414 7008 9470
rect 6668 9328 7008 9414
rect 6668 9272 6742 9328
rect 6798 9272 6884 9328
rect 6940 9272 7008 9328
rect 6668 9186 7008 9272
rect 6668 9130 6742 9186
rect 6798 9130 6884 9186
rect 6940 9130 7008 9186
rect 6668 9044 7008 9130
rect 6668 8988 6742 9044
rect 6798 8988 6884 9044
rect 6940 8988 7008 9044
rect 6668 8902 7008 8988
rect 6668 8846 6742 8902
rect 6798 8846 6884 8902
rect 6940 8846 7008 8902
rect 6668 8760 7008 8846
rect 6668 8704 6742 8760
rect 6798 8704 6884 8760
rect 6940 8704 7008 8760
rect 6668 8618 7008 8704
rect 6668 8562 6742 8618
rect 6798 8562 6884 8618
rect 6940 8562 7008 8618
rect 6668 8476 7008 8562
rect 6668 8420 6742 8476
rect 6798 8420 6884 8476
rect 6940 8420 7008 8476
rect 6668 8334 7008 8420
rect 6668 8278 6742 8334
rect 6798 8278 6884 8334
rect 6940 8278 7008 8334
rect 6668 8192 7008 8278
rect 6668 8136 6742 8192
rect 6798 8136 6884 8192
rect 6940 8136 7008 8192
rect 6668 8050 7008 8136
rect 6668 7994 6742 8050
rect 6798 7994 6884 8050
rect 6940 7994 7008 8050
rect 6668 7908 7008 7994
rect 6668 7852 6742 7908
rect 6798 7852 6884 7908
rect 6940 7852 7008 7908
rect 6668 7766 7008 7852
rect 6668 7710 6742 7766
rect 6798 7710 6884 7766
rect 6940 7710 7008 7766
rect 6668 7624 7008 7710
rect 6668 7568 6742 7624
rect 6798 7568 6884 7624
rect 6940 7568 7008 7624
rect 6668 7482 7008 7568
rect 6668 7426 6742 7482
rect 6798 7426 6884 7482
rect 6940 7426 7008 7482
rect 6668 7340 7008 7426
rect 6668 7284 6742 7340
rect 6798 7284 6884 7340
rect 6940 7284 7008 7340
rect 6668 7198 7008 7284
rect 6668 7142 6742 7198
rect 6798 7142 6884 7198
rect 6940 7142 7008 7198
rect 6668 7056 7008 7142
rect 6668 7000 6742 7056
rect 6798 7000 6884 7056
rect 6940 7000 7008 7056
rect 6668 6914 7008 7000
rect 6668 6858 6742 6914
rect 6798 6858 6884 6914
rect 6940 6858 7008 6914
rect 6668 6772 7008 6858
rect 6668 6716 6742 6772
rect 6798 6716 6884 6772
rect 6940 6716 7008 6772
rect 6668 6630 7008 6716
rect 6668 6574 6742 6630
rect 6798 6574 6884 6630
rect 6940 6574 7008 6630
rect 6668 6488 7008 6574
rect 6668 6432 6742 6488
rect 6798 6432 6884 6488
rect 6940 6432 7008 6488
rect 6668 6346 7008 6432
rect 6668 6290 6742 6346
rect 6798 6290 6884 6346
rect 6940 6290 7008 6346
rect 6668 6204 7008 6290
rect 6668 6148 6742 6204
rect 6798 6148 6884 6204
rect 6940 6148 7008 6204
rect 6668 6062 7008 6148
rect 6668 6006 6742 6062
rect 6798 6006 6884 6062
rect 6940 6006 7008 6062
rect 6668 5920 7008 6006
rect 6668 5864 6742 5920
rect 6798 5864 6884 5920
rect 6940 5864 7008 5920
rect 6668 5778 7008 5864
rect 6668 5722 6742 5778
rect 6798 5722 6884 5778
rect 6940 5722 7008 5778
rect 6668 5636 7008 5722
rect 6668 5580 6742 5636
rect 6798 5580 6884 5636
rect 6940 5580 7008 5636
rect 6668 5494 7008 5580
rect 6668 5438 6742 5494
rect 6798 5438 6884 5494
rect 6940 5438 7008 5494
rect 6668 5352 7008 5438
rect 6668 5296 6742 5352
rect 6798 5296 6884 5352
rect 6940 5296 7008 5352
rect 6668 5210 7008 5296
rect 6668 5154 6742 5210
rect 6798 5154 6884 5210
rect 6940 5154 7008 5210
rect 6668 5068 7008 5154
rect 6668 5012 6742 5068
rect 6798 5012 6884 5068
rect 6940 5012 7008 5068
rect 6668 4926 7008 5012
rect 6668 4870 6742 4926
rect 6798 4870 6884 4926
rect 6940 4870 7008 4926
rect 6668 4784 7008 4870
rect 6668 4728 6742 4784
rect 6798 4728 6884 4784
rect 6940 4728 7008 4784
rect 6668 4642 7008 4728
rect 6668 4586 6742 4642
rect 6798 4586 6884 4642
rect 6940 4586 7008 4642
rect 6668 4500 7008 4586
rect 6668 4444 6742 4500
rect 6798 4444 6884 4500
rect 6940 4444 7008 4500
rect 6668 4358 7008 4444
rect 6668 4302 6742 4358
rect 6798 4302 6884 4358
rect 6940 4302 7008 4358
rect 6668 4216 7008 4302
rect 6668 4160 6742 4216
rect 6798 4160 6884 4216
rect 6940 4160 7008 4216
rect 6668 4074 7008 4160
rect 6668 4018 6742 4074
rect 6798 4018 6884 4074
rect 6940 4018 7008 4074
rect 6668 3932 7008 4018
rect 6668 3876 6742 3932
rect 6798 3876 6884 3932
rect 6940 3876 7008 3932
rect 6668 3790 7008 3876
rect 6668 3734 6742 3790
rect 6798 3734 6884 3790
rect 6940 3734 7008 3790
rect 6668 3648 7008 3734
rect 6668 3592 6742 3648
rect 6798 3592 6884 3648
rect 6940 3592 7008 3648
rect 6668 3506 7008 3592
rect 6668 3450 6742 3506
rect 6798 3450 6884 3506
rect 6940 3450 7008 3506
rect 6668 3364 7008 3450
rect 6668 3308 6742 3364
rect 6798 3308 6884 3364
rect 6940 3308 7008 3364
rect 6668 3222 7008 3308
rect 6668 3166 6742 3222
rect 6798 3166 6884 3222
rect 6940 3166 7008 3222
rect 6668 3080 7008 3166
rect 6668 3024 6742 3080
rect 6798 3024 6884 3080
rect 6940 3024 7008 3080
rect 6668 2938 7008 3024
rect 6668 2882 6742 2938
rect 6798 2882 6884 2938
rect 6940 2882 7008 2938
rect 6668 2796 7008 2882
rect 6668 2740 6742 2796
rect 6798 2740 6884 2796
rect 6940 2740 7008 2796
rect 6668 2654 7008 2740
rect 6668 2598 6742 2654
rect 6798 2598 6884 2654
rect 6940 2598 7008 2654
rect 6668 2512 7008 2598
rect 6668 2456 6742 2512
rect 6798 2456 6884 2512
rect 6940 2456 7008 2512
rect 6668 2370 7008 2456
rect 6668 2314 6742 2370
rect 6798 2314 6884 2370
rect 6940 2314 7008 2370
rect 6668 2228 7008 2314
rect 6668 2172 6742 2228
rect 6798 2172 6884 2228
rect 6940 2172 7008 2228
rect 6668 2086 7008 2172
rect 6668 2030 6742 2086
rect 6798 2030 6884 2086
rect 6940 2030 7008 2086
rect 6668 1944 7008 2030
rect 6668 1888 6742 1944
rect 6798 1888 6884 1944
rect 6940 1888 7008 1944
rect 6668 1802 7008 1888
rect 6668 1746 6742 1802
rect 6798 1746 6884 1802
rect 6940 1746 7008 1802
rect 6668 1660 7008 1746
rect 6668 1604 6742 1660
rect 6798 1604 6884 1660
rect 6940 1604 7008 1660
rect 6668 1518 7008 1604
rect 6668 1462 6742 1518
rect 6798 1462 6884 1518
rect 6940 1462 7008 1518
rect 6668 1376 7008 1462
rect 6668 1320 6742 1376
rect 6798 1320 6884 1376
rect 6940 1320 7008 1376
rect 6668 1234 7008 1320
rect 6668 1178 6742 1234
rect 6798 1178 6884 1234
rect 6940 1178 7008 1234
rect 6668 1092 7008 1178
rect 6668 1036 6742 1092
rect 6798 1036 6884 1092
rect 6940 1036 7008 1092
rect 6668 950 7008 1036
rect 6668 894 6742 950
rect 6798 894 6884 950
rect 6940 894 7008 950
rect 6668 808 7008 894
rect 6668 752 6742 808
rect 6798 752 6884 808
rect 6940 752 7008 808
rect 6668 666 7008 752
rect 6668 610 6742 666
rect 6798 610 6884 666
rect 6940 610 7008 666
rect 6668 524 7008 610
rect 6668 468 6742 524
rect 6798 468 6884 524
rect 6940 468 7008 524
rect 6668 400 7008 468
rect 7068 12310 7408 12400
rect 7068 12254 7145 12310
rect 7201 12254 7287 12310
rect 7343 12254 7408 12310
rect 7068 12168 7408 12254
rect 7068 12112 7145 12168
rect 7201 12112 7287 12168
rect 7343 12112 7408 12168
rect 7068 12026 7408 12112
rect 7068 11970 7145 12026
rect 7201 11970 7287 12026
rect 7343 11970 7408 12026
rect 7068 11884 7408 11970
rect 7068 11828 7145 11884
rect 7201 11828 7287 11884
rect 7343 11828 7408 11884
rect 7068 11742 7408 11828
rect 7068 11686 7145 11742
rect 7201 11686 7287 11742
rect 7343 11686 7408 11742
rect 7068 11600 7408 11686
rect 7068 11544 7145 11600
rect 7201 11544 7287 11600
rect 7343 11544 7408 11600
rect 7068 11458 7408 11544
rect 7068 11402 7145 11458
rect 7201 11402 7287 11458
rect 7343 11402 7408 11458
rect 7068 11316 7408 11402
rect 7068 11260 7145 11316
rect 7201 11260 7287 11316
rect 7343 11260 7408 11316
rect 7068 11174 7408 11260
rect 7068 11118 7145 11174
rect 7201 11118 7287 11174
rect 7343 11118 7408 11174
rect 7068 11032 7408 11118
rect 7068 10976 7145 11032
rect 7201 10976 7287 11032
rect 7343 10976 7408 11032
rect 7068 10890 7408 10976
rect 7068 10834 7145 10890
rect 7201 10834 7287 10890
rect 7343 10834 7408 10890
rect 7068 10748 7408 10834
rect 7068 10692 7145 10748
rect 7201 10692 7287 10748
rect 7343 10692 7408 10748
rect 7068 10606 7408 10692
rect 7068 10550 7145 10606
rect 7201 10550 7287 10606
rect 7343 10550 7408 10606
rect 7068 10464 7408 10550
rect 7068 10408 7145 10464
rect 7201 10408 7287 10464
rect 7343 10408 7408 10464
rect 7068 10322 7408 10408
rect 7068 10266 7145 10322
rect 7201 10266 7287 10322
rect 7343 10266 7408 10322
rect 7068 10180 7408 10266
rect 7068 10124 7145 10180
rect 7201 10124 7287 10180
rect 7343 10124 7408 10180
rect 7068 10038 7408 10124
rect 7068 9982 7145 10038
rect 7201 9982 7287 10038
rect 7343 9982 7408 10038
rect 7068 9896 7408 9982
rect 7068 9840 7145 9896
rect 7201 9840 7287 9896
rect 7343 9840 7408 9896
rect 7068 9754 7408 9840
rect 7068 9698 7145 9754
rect 7201 9698 7287 9754
rect 7343 9698 7408 9754
rect 7068 9612 7408 9698
rect 7068 9556 7145 9612
rect 7201 9556 7287 9612
rect 7343 9556 7408 9612
rect 7068 9470 7408 9556
rect 7068 9414 7145 9470
rect 7201 9414 7287 9470
rect 7343 9414 7408 9470
rect 7068 9328 7408 9414
rect 7068 9272 7145 9328
rect 7201 9272 7287 9328
rect 7343 9272 7408 9328
rect 7068 9186 7408 9272
rect 7068 9130 7145 9186
rect 7201 9130 7287 9186
rect 7343 9130 7408 9186
rect 7068 9044 7408 9130
rect 7068 8988 7145 9044
rect 7201 8988 7287 9044
rect 7343 8988 7408 9044
rect 7068 8902 7408 8988
rect 7068 8846 7145 8902
rect 7201 8846 7287 8902
rect 7343 8846 7408 8902
rect 7068 8760 7408 8846
rect 7068 8704 7145 8760
rect 7201 8704 7287 8760
rect 7343 8704 7408 8760
rect 7068 8618 7408 8704
rect 7068 8562 7145 8618
rect 7201 8562 7287 8618
rect 7343 8562 7408 8618
rect 7068 8476 7408 8562
rect 7068 8420 7145 8476
rect 7201 8420 7287 8476
rect 7343 8420 7408 8476
rect 7068 8334 7408 8420
rect 7068 8278 7145 8334
rect 7201 8278 7287 8334
rect 7343 8278 7408 8334
rect 7068 8192 7408 8278
rect 7068 8136 7145 8192
rect 7201 8136 7287 8192
rect 7343 8136 7408 8192
rect 7068 8050 7408 8136
rect 7068 7994 7145 8050
rect 7201 7994 7287 8050
rect 7343 7994 7408 8050
rect 7068 7908 7408 7994
rect 7068 7852 7145 7908
rect 7201 7852 7287 7908
rect 7343 7852 7408 7908
rect 7068 7766 7408 7852
rect 7068 7710 7145 7766
rect 7201 7710 7287 7766
rect 7343 7710 7408 7766
rect 7068 7624 7408 7710
rect 7068 7568 7145 7624
rect 7201 7568 7287 7624
rect 7343 7568 7408 7624
rect 7068 7482 7408 7568
rect 7068 7426 7145 7482
rect 7201 7426 7287 7482
rect 7343 7426 7408 7482
rect 7068 7340 7408 7426
rect 7068 7284 7145 7340
rect 7201 7284 7287 7340
rect 7343 7284 7408 7340
rect 7068 7198 7408 7284
rect 7068 7142 7145 7198
rect 7201 7142 7287 7198
rect 7343 7142 7408 7198
rect 7068 7056 7408 7142
rect 7068 7000 7145 7056
rect 7201 7000 7287 7056
rect 7343 7000 7408 7056
rect 7068 6914 7408 7000
rect 7068 6858 7145 6914
rect 7201 6858 7287 6914
rect 7343 6858 7408 6914
rect 7068 6772 7408 6858
rect 7068 6716 7145 6772
rect 7201 6716 7287 6772
rect 7343 6716 7408 6772
rect 7068 6630 7408 6716
rect 7068 6574 7145 6630
rect 7201 6574 7287 6630
rect 7343 6574 7408 6630
rect 7068 6488 7408 6574
rect 7068 6432 7145 6488
rect 7201 6432 7287 6488
rect 7343 6432 7408 6488
rect 7068 6346 7408 6432
rect 7068 6290 7145 6346
rect 7201 6290 7287 6346
rect 7343 6290 7408 6346
rect 7068 6204 7408 6290
rect 7068 6148 7145 6204
rect 7201 6148 7287 6204
rect 7343 6148 7408 6204
rect 7068 6062 7408 6148
rect 7068 6006 7145 6062
rect 7201 6006 7287 6062
rect 7343 6006 7408 6062
rect 7068 5920 7408 6006
rect 7068 5864 7145 5920
rect 7201 5864 7287 5920
rect 7343 5864 7408 5920
rect 7068 5778 7408 5864
rect 7068 5722 7145 5778
rect 7201 5722 7287 5778
rect 7343 5722 7408 5778
rect 7068 5636 7408 5722
rect 7068 5580 7145 5636
rect 7201 5580 7287 5636
rect 7343 5580 7408 5636
rect 7068 5494 7408 5580
rect 7068 5438 7145 5494
rect 7201 5438 7287 5494
rect 7343 5438 7408 5494
rect 7068 5352 7408 5438
rect 7068 5296 7145 5352
rect 7201 5296 7287 5352
rect 7343 5296 7408 5352
rect 7068 5210 7408 5296
rect 7068 5154 7145 5210
rect 7201 5154 7287 5210
rect 7343 5154 7408 5210
rect 7068 5068 7408 5154
rect 7068 5012 7145 5068
rect 7201 5012 7287 5068
rect 7343 5012 7408 5068
rect 7068 4926 7408 5012
rect 7068 4870 7145 4926
rect 7201 4870 7287 4926
rect 7343 4870 7408 4926
rect 7068 4784 7408 4870
rect 7068 4728 7145 4784
rect 7201 4728 7287 4784
rect 7343 4728 7408 4784
rect 7068 4642 7408 4728
rect 7068 4586 7145 4642
rect 7201 4586 7287 4642
rect 7343 4586 7408 4642
rect 7068 4500 7408 4586
rect 7068 4444 7145 4500
rect 7201 4444 7287 4500
rect 7343 4444 7408 4500
rect 7068 4358 7408 4444
rect 7068 4302 7145 4358
rect 7201 4302 7287 4358
rect 7343 4302 7408 4358
rect 7068 4216 7408 4302
rect 7068 4160 7145 4216
rect 7201 4160 7287 4216
rect 7343 4160 7408 4216
rect 7068 4074 7408 4160
rect 7068 4018 7145 4074
rect 7201 4018 7287 4074
rect 7343 4018 7408 4074
rect 7068 3932 7408 4018
rect 7068 3876 7145 3932
rect 7201 3876 7287 3932
rect 7343 3876 7408 3932
rect 7068 3790 7408 3876
rect 7068 3734 7145 3790
rect 7201 3734 7287 3790
rect 7343 3734 7408 3790
rect 7068 3648 7408 3734
rect 7068 3592 7145 3648
rect 7201 3592 7287 3648
rect 7343 3592 7408 3648
rect 7068 3506 7408 3592
rect 7068 3450 7145 3506
rect 7201 3450 7287 3506
rect 7343 3450 7408 3506
rect 7068 3364 7408 3450
rect 7068 3308 7145 3364
rect 7201 3308 7287 3364
rect 7343 3308 7408 3364
rect 7068 3222 7408 3308
rect 7068 3166 7145 3222
rect 7201 3166 7287 3222
rect 7343 3166 7408 3222
rect 7068 3080 7408 3166
rect 7068 3024 7145 3080
rect 7201 3024 7287 3080
rect 7343 3024 7408 3080
rect 7068 2938 7408 3024
rect 7068 2882 7145 2938
rect 7201 2882 7287 2938
rect 7343 2882 7408 2938
rect 7068 2796 7408 2882
rect 7068 2740 7145 2796
rect 7201 2740 7287 2796
rect 7343 2740 7408 2796
rect 7068 2654 7408 2740
rect 7068 2598 7145 2654
rect 7201 2598 7287 2654
rect 7343 2598 7408 2654
rect 7068 2512 7408 2598
rect 7068 2456 7145 2512
rect 7201 2456 7287 2512
rect 7343 2456 7408 2512
rect 7068 2370 7408 2456
rect 7068 2314 7145 2370
rect 7201 2314 7287 2370
rect 7343 2314 7408 2370
rect 7068 2228 7408 2314
rect 7068 2172 7145 2228
rect 7201 2172 7287 2228
rect 7343 2172 7408 2228
rect 7068 2086 7408 2172
rect 7068 2030 7145 2086
rect 7201 2030 7287 2086
rect 7343 2030 7408 2086
rect 7068 1944 7408 2030
rect 7068 1888 7145 1944
rect 7201 1888 7287 1944
rect 7343 1888 7408 1944
rect 7068 1802 7408 1888
rect 7068 1746 7145 1802
rect 7201 1746 7287 1802
rect 7343 1746 7408 1802
rect 7068 1660 7408 1746
rect 7068 1604 7145 1660
rect 7201 1604 7287 1660
rect 7343 1604 7408 1660
rect 7068 1518 7408 1604
rect 7068 1462 7145 1518
rect 7201 1462 7287 1518
rect 7343 1462 7408 1518
rect 7068 1376 7408 1462
rect 7068 1320 7145 1376
rect 7201 1320 7287 1376
rect 7343 1320 7408 1376
rect 7068 1234 7408 1320
rect 7068 1178 7145 1234
rect 7201 1178 7287 1234
rect 7343 1178 7408 1234
rect 7068 1092 7408 1178
rect 7068 1036 7145 1092
rect 7201 1036 7287 1092
rect 7343 1036 7408 1092
rect 7068 950 7408 1036
rect 7068 894 7145 950
rect 7201 894 7287 950
rect 7343 894 7408 950
rect 7068 808 7408 894
rect 7068 752 7145 808
rect 7201 752 7287 808
rect 7343 752 7408 808
rect 7068 666 7408 752
rect 7068 610 7145 666
rect 7201 610 7287 666
rect 7343 610 7408 666
rect 7068 524 7408 610
rect 7068 468 7145 524
rect 7201 468 7287 524
rect 7343 468 7408 524
rect 7068 400 7408 468
rect 7468 12310 7808 12400
rect 7468 12254 7539 12310
rect 7595 12254 7681 12310
rect 7737 12254 7808 12310
rect 7468 12168 7808 12254
rect 7468 12112 7539 12168
rect 7595 12112 7681 12168
rect 7737 12112 7808 12168
rect 7468 12026 7808 12112
rect 7468 11970 7539 12026
rect 7595 11970 7681 12026
rect 7737 11970 7808 12026
rect 7468 11884 7808 11970
rect 7468 11828 7539 11884
rect 7595 11828 7681 11884
rect 7737 11828 7808 11884
rect 7468 11742 7808 11828
rect 7468 11686 7539 11742
rect 7595 11686 7681 11742
rect 7737 11686 7808 11742
rect 7468 11600 7808 11686
rect 7468 11544 7539 11600
rect 7595 11544 7681 11600
rect 7737 11544 7808 11600
rect 7468 11458 7808 11544
rect 7468 11402 7539 11458
rect 7595 11402 7681 11458
rect 7737 11402 7808 11458
rect 7468 11316 7808 11402
rect 7468 11260 7539 11316
rect 7595 11260 7681 11316
rect 7737 11260 7808 11316
rect 7468 11174 7808 11260
rect 7468 11118 7539 11174
rect 7595 11118 7681 11174
rect 7737 11118 7808 11174
rect 7468 11032 7808 11118
rect 7468 10976 7539 11032
rect 7595 10976 7681 11032
rect 7737 10976 7808 11032
rect 7468 10890 7808 10976
rect 7468 10834 7539 10890
rect 7595 10834 7681 10890
rect 7737 10834 7808 10890
rect 7468 10748 7808 10834
rect 7468 10692 7539 10748
rect 7595 10692 7681 10748
rect 7737 10692 7808 10748
rect 7468 10606 7808 10692
rect 7468 10550 7539 10606
rect 7595 10550 7681 10606
rect 7737 10550 7808 10606
rect 7468 10464 7808 10550
rect 7468 10408 7539 10464
rect 7595 10408 7681 10464
rect 7737 10408 7808 10464
rect 7468 10322 7808 10408
rect 7468 10266 7539 10322
rect 7595 10266 7681 10322
rect 7737 10266 7808 10322
rect 7468 10180 7808 10266
rect 7468 10124 7539 10180
rect 7595 10124 7681 10180
rect 7737 10124 7808 10180
rect 7468 10038 7808 10124
rect 7468 9982 7539 10038
rect 7595 9982 7681 10038
rect 7737 9982 7808 10038
rect 7468 9896 7808 9982
rect 7468 9840 7539 9896
rect 7595 9840 7681 9896
rect 7737 9840 7808 9896
rect 7468 9754 7808 9840
rect 7468 9698 7539 9754
rect 7595 9698 7681 9754
rect 7737 9698 7808 9754
rect 7468 9612 7808 9698
rect 7468 9556 7539 9612
rect 7595 9556 7681 9612
rect 7737 9556 7808 9612
rect 7468 9470 7808 9556
rect 7468 9414 7539 9470
rect 7595 9414 7681 9470
rect 7737 9414 7808 9470
rect 7468 9328 7808 9414
rect 7468 9272 7539 9328
rect 7595 9272 7681 9328
rect 7737 9272 7808 9328
rect 7468 9186 7808 9272
rect 7468 9130 7539 9186
rect 7595 9130 7681 9186
rect 7737 9130 7808 9186
rect 7468 9044 7808 9130
rect 7468 8988 7539 9044
rect 7595 8988 7681 9044
rect 7737 8988 7808 9044
rect 7468 8902 7808 8988
rect 7468 8846 7539 8902
rect 7595 8846 7681 8902
rect 7737 8846 7808 8902
rect 7468 8760 7808 8846
rect 7468 8704 7539 8760
rect 7595 8704 7681 8760
rect 7737 8704 7808 8760
rect 7468 8618 7808 8704
rect 7468 8562 7539 8618
rect 7595 8562 7681 8618
rect 7737 8562 7808 8618
rect 7468 8476 7808 8562
rect 7468 8420 7539 8476
rect 7595 8420 7681 8476
rect 7737 8420 7808 8476
rect 7468 8334 7808 8420
rect 7468 8278 7539 8334
rect 7595 8278 7681 8334
rect 7737 8278 7808 8334
rect 7468 8192 7808 8278
rect 7468 8136 7539 8192
rect 7595 8136 7681 8192
rect 7737 8136 7808 8192
rect 7468 8050 7808 8136
rect 7468 7994 7539 8050
rect 7595 7994 7681 8050
rect 7737 7994 7808 8050
rect 7468 7908 7808 7994
rect 7468 7852 7539 7908
rect 7595 7852 7681 7908
rect 7737 7852 7808 7908
rect 7468 7766 7808 7852
rect 7468 7710 7539 7766
rect 7595 7710 7681 7766
rect 7737 7710 7808 7766
rect 7468 7624 7808 7710
rect 7468 7568 7539 7624
rect 7595 7568 7681 7624
rect 7737 7568 7808 7624
rect 7468 7482 7808 7568
rect 7468 7426 7539 7482
rect 7595 7426 7681 7482
rect 7737 7426 7808 7482
rect 7468 7340 7808 7426
rect 7468 7284 7539 7340
rect 7595 7284 7681 7340
rect 7737 7284 7808 7340
rect 7468 7198 7808 7284
rect 7468 7142 7539 7198
rect 7595 7142 7681 7198
rect 7737 7142 7808 7198
rect 7468 7056 7808 7142
rect 7468 7000 7539 7056
rect 7595 7000 7681 7056
rect 7737 7000 7808 7056
rect 7468 6914 7808 7000
rect 7468 6858 7539 6914
rect 7595 6858 7681 6914
rect 7737 6858 7808 6914
rect 7468 6772 7808 6858
rect 7468 6716 7539 6772
rect 7595 6716 7681 6772
rect 7737 6716 7808 6772
rect 7468 6630 7808 6716
rect 7468 6574 7539 6630
rect 7595 6574 7681 6630
rect 7737 6574 7808 6630
rect 7468 6488 7808 6574
rect 7468 6432 7539 6488
rect 7595 6432 7681 6488
rect 7737 6432 7808 6488
rect 7468 6346 7808 6432
rect 7468 6290 7539 6346
rect 7595 6290 7681 6346
rect 7737 6290 7808 6346
rect 7468 6204 7808 6290
rect 7468 6148 7539 6204
rect 7595 6148 7681 6204
rect 7737 6148 7808 6204
rect 7468 6062 7808 6148
rect 7468 6006 7539 6062
rect 7595 6006 7681 6062
rect 7737 6006 7808 6062
rect 7468 5920 7808 6006
rect 7468 5864 7539 5920
rect 7595 5864 7681 5920
rect 7737 5864 7808 5920
rect 7468 5778 7808 5864
rect 7468 5722 7539 5778
rect 7595 5722 7681 5778
rect 7737 5722 7808 5778
rect 7468 5636 7808 5722
rect 7468 5580 7539 5636
rect 7595 5580 7681 5636
rect 7737 5580 7808 5636
rect 7468 5494 7808 5580
rect 7468 5438 7539 5494
rect 7595 5438 7681 5494
rect 7737 5438 7808 5494
rect 7468 5352 7808 5438
rect 7468 5296 7539 5352
rect 7595 5296 7681 5352
rect 7737 5296 7808 5352
rect 7468 5210 7808 5296
rect 7468 5154 7539 5210
rect 7595 5154 7681 5210
rect 7737 5154 7808 5210
rect 7468 5068 7808 5154
rect 7468 5012 7539 5068
rect 7595 5012 7681 5068
rect 7737 5012 7808 5068
rect 7468 4926 7808 5012
rect 7468 4870 7539 4926
rect 7595 4870 7681 4926
rect 7737 4870 7808 4926
rect 7468 4784 7808 4870
rect 7468 4728 7539 4784
rect 7595 4728 7681 4784
rect 7737 4728 7808 4784
rect 7468 4642 7808 4728
rect 7468 4586 7539 4642
rect 7595 4586 7681 4642
rect 7737 4586 7808 4642
rect 7468 4500 7808 4586
rect 7468 4444 7539 4500
rect 7595 4444 7681 4500
rect 7737 4444 7808 4500
rect 7468 4358 7808 4444
rect 7468 4302 7539 4358
rect 7595 4302 7681 4358
rect 7737 4302 7808 4358
rect 7468 4216 7808 4302
rect 7468 4160 7539 4216
rect 7595 4160 7681 4216
rect 7737 4160 7808 4216
rect 7468 4074 7808 4160
rect 7468 4018 7539 4074
rect 7595 4018 7681 4074
rect 7737 4018 7808 4074
rect 7468 3932 7808 4018
rect 7468 3876 7539 3932
rect 7595 3876 7681 3932
rect 7737 3876 7808 3932
rect 7468 3790 7808 3876
rect 7468 3734 7539 3790
rect 7595 3734 7681 3790
rect 7737 3734 7808 3790
rect 7468 3648 7808 3734
rect 7468 3592 7539 3648
rect 7595 3592 7681 3648
rect 7737 3592 7808 3648
rect 7468 3506 7808 3592
rect 7468 3450 7539 3506
rect 7595 3450 7681 3506
rect 7737 3450 7808 3506
rect 7468 3364 7808 3450
rect 7468 3308 7539 3364
rect 7595 3308 7681 3364
rect 7737 3308 7808 3364
rect 7468 3222 7808 3308
rect 7468 3166 7539 3222
rect 7595 3166 7681 3222
rect 7737 3166 7808 3222
rect 7468 3080 7808 3166
rect 7468 3024 7539 3080
rect 7595 3024 7681 3080
rect 7737 3024 7808 3080
rect 7468 2938 7808 3024
rect 7468 2882 7539 2938
rect 7595 2882 7681 2938
rect 7737 2882 7808 2938
rect 7468 2796 7808 2882
rect 7468 2740 7539 2796
rect 7595 2740 7681 2796
rect 7737 2740 7808 2796
rect 7468 2654 7808 2740
rect 7468 2598 7539 2654
rect 7595 2598 7681 2654
rect 7737 2598 7808 2654
rect 7468 2512 7808 2598
rect 7468 2456 7539 2512
rect 7595 2456 7681 2512
rect 7737 2456 7808 2512
rect 7468 2370 7808 2456
rect 7468 2314 7539 2370
rect 7595 2314 7681 2370
rect 7737 2314 7808 2370
rect 7468 2228 7808 2314
rect 7468 2172 7539 2228
rect 7595 2172 7681 2228
rect 7737 2172 7808 2228
rect 7468 2086 7808 2172
rect 7468 2030 7539 2086
rect 7595 2030 7681 2086
rect 7737 2030 7808 2086
rect 7468 1944 7808 2030
rect 7468 1888 7539 1944
rect 7595 1888 7681 1944
rect 7737 1888 7808 1944
rect 7468 1802 7808 1888
rect 7468 1746 7539 1802
rect 7595 1746 7681 1802
rect 7737 1746 7808 1802
rect 7468 1660 7808 1746
rect 7468 1604 7539 1660
rect 7595 1604 7681 1660
rect 7737 1604 7808 1660
rect 7468 1518 7808 1604
rect 7468 1462 7539 1518
rect 7595 1462 7681 1518
rect 7737 1462 7808 1518
rect 7468 1376 7808 1462
rect 7468 1320 7539 1376
rect 7595 1320 7681 1376
rect 7737 1320 7808 1376
rect 7468 1234 7808 1320
rect 7468 1178 7539 1234
rect 7595 1178 7681 1234
rect 7737 1178 7808 1234
rect 7468 1092 7808 1178
rect 7468 1036 7539 1092
rect 7595 1036 7681 1092
rect 7737 1036 7808 1092
rect 7468 950 7808 1036
rect 7468 894 7539 950
rect 7595 894 7681 950
rect 7737 894 7808 950
rect 7468 808 7808 894
rect 7468 752 7539 808
rect 7595 752 7681 808
rect 7737 752 7808 808
rect 7468 666 7808 752
rect 7468 610 7539 666
rect 7595 610 7681 666
rect 7737 610 7808 666
rect 7468 524 7808 610
rect 7468 468 7539 524
rect 7595 468 7681 524
rect 7737 468 7808 524
rect 7468 400 7808 468
rect 7868 12310 8208 12400
rect 7868 12254 7940 12310
rect 7996 12254 8082 12310
rect 8138 12254 8208 12310
rect 7868 12168 8208 12254
rect 7868 12112 7940 12168
rect 7996 12112 8082 12168
rect 8138 12112 8208 12168
rect 7868 12026 8208 12112
rect 7868 11970 7940 12026
rect 7996 11970 8082 12026
rect 8138 11970 8208 12026
rect 7868 11884 8208 11970
rect 7868 11828 7940 11884
rect 7996 11828 8082 11884
rect 8138 11828 8208 11884
rect 7868 11742 8208 11828
rect 7868 11686 7940 11742
rect 7996 11686 8082 11742
rect 8138 11686 8208 11742
rect 7868 11600 8208 11686
rect 7868 11544 7940 11600
rect 7996 11544 8082 11600
rect 8138 11544 8208 11600
rect 7868 11458 8208 11544
rect 7868 11402 7940 11458
rect 7996 11402 8082 11458
rect 8138 11402 8208 11458
rect 7868 11316 8208 11402
rect 7868 11260 7940 11316
rect 7996 11260 8082 11316
rect 8138 11260 8208 11316
rect 7868 11174 8208 11260
rect 7868 11118 7940 11174
rect 7996 11118 8082 11174
rect 8138 11118 8208 11174
rect 7868 11032 8208 11118
rect 7868 10976 7940 11032
rect 7996 10976 8082 11032
rect 8138 10976 8208 11032
rect 7868 10890 8208 10976
rect 7868 10834 7940 10890
rect 7996 10834 8082 10890
rect 8138 10834 8208 10890
rect 7868 10748 8208 10834
rect 7868 10692 7940 10748
rect 7996 10692 8082 10748
rect 8138 10692 8208 10748
rect 7868 10606 8208 10692
rect 7868 10550 7940 10606
rect 7996 10550 8082 10606
rect 8138 10550 8208 10606
rect 7868 10464 8208 10550
rect 7868 10408 7940 10464
rect 7996 10408 8082 10464
rect 8138 10408 8208 10464
rect 7868 10322 8208 10408
rect 7868 10266 7940 10322
rect 7996 10266 8082 10322
rect 8138 10266 8208 10322
rect 7868 10180 8208 10266
rect 7868 10124 7940 10180
rect 7996 10124 8082 10180
rect 8138 10124 8208 10180
rect 7868 10038 8208 10124
rect 7868 9982 7940 10038
rect 7996 9982 8082 10038
rect 8138 9982 8208 10038
rect 7868 9896 8208 9982
rect 7868 9840 7940 9896
rect 7996 9840 8082 9896
rect 8138 9840 8208 9896
rect 7868 9754 8208 9840
rect 7868 9698 7940 9754
rect 7996 9698 8082 9754
rect 8138 9698 8208 9754
rect 7868 9612 8208 9698
rect 7868 9556 7940 9612
rect 7996 9556 8082 9612
rect 8138 9556 8208 9612
rect 7868 9470 8208 9556
rect 7868 9414 7940 9470
rect 7996 9414 8082 9470
rect 8138 9414 8208 9470
rect 7868 9328 8208 9414
rect 7868 9272 7940 9328
rect 7996 9272 8082 9328
rect 8138 9272 8208 9328
rect 7868 9186 8208 9272
rect 7868 9130 7940 9186
rect 7996 9130 8082 9186
rect 8138 9130 8208 9186
rect 7868 9044 8208 9130
rect 7868 8988 7940 9044
rect 7996 8988 8082 9044
rect 8138 8988 8208 9044
rect 7868 8902 8208 8988
rect 7868 8846 7940 8902
rect 7996 8846 8082 8902
rect 8138 8846 8208 8902
rect 7868 8760 8208 8846
rect 7868 8704 7940 8760
rect 7996 8704 8082 8760
rect 8138 8704 8208 8760
rect 7868 8618 8208 8704
rect 7868 8562 7940 8618
rect 7996 8562 8082 8618
rect 8138 8562 8208 8618
rect 7868 8476 8208 8562
rect 7868 8420 7940 8476
rect 7996 8420 8082 8476
rect 8138 8420 8208 8476
rect 7868 8334 8208 8420
rect 7868 8278 7940 8334
rect 7996 8278 8082 8334
rect 8138 8278 8208 8334
rect 7868 8192 8208 8278
rect 7868 8136 7940 8192
rect 7996 8136 8082 8192
rect 8138 8136 8208 8192
rect 7868 8050 8208 8136
rect 7868 7994 7940 8050
rect 7996 7994 8082 8050
rect 8138 7994 8208 8050
rect 7868 7908 8208 7994
rect 7868 7852 7940 7908
rect 7996 7852 8082 7908
rect 8138 7852 8208 7908
rect 7868 7766 8208 7852
rect 7868 7710 7940 7766
rect 7996 7710 8082 7766
rect 8138 7710 8208 7766
rect 7868 7624 8208 7710
rect 7868 7568 7940 7624
rect 7996 7568 8082 7624
rect 8138 7568 8208 7624
rect 7868 7482 8208 7568
rect 7868 7426 7940 7482
rect 7996 7426 8082 7482
rect 8138 7426 8208 7482
rect 7868 7340 8208 7426
rect 7868 7284 7940 7340
rect 7996 7284 8082 7340
rect 8138 7284 8208 7340
rect 7868 7198 8208 7284
rect 7868 7142 7940 7198
rect 7996 7142 8082 7198
rect 8138 7142 8208 7198
rect 7868 7056 8208 7142
rect 7868 7000 7940 7056
rect 7996 7000 8082 7056
rect 8138 7000 8208 7056
rect 7868 6914 8208 7000
rect 7868 6858 7940 6914
rect 7996 6858 8082 6914
rect 8138 6858 8208 6914
rect 7868 6772 8208 6858
rect 7868 6716 7940 6772
rect 7996 6716 8082 6772
rect 8138 6716 8208 6772
rect 7868 6630 8208 6716
rect 7868 6574 7940 6630
rect 7996 6574 8082 6630
rect 8138 6574 8208 6630
rect 7868 6488 8208 6574
rect 7868 6432 7940 6488
rect 7996 6432 8082 6488
rect 8138 6432 8208 6488
rect 7868 6346 8208 6432
rect 7868 6290 7940 6346
rect 7996 6290 8082 6346
rect 8138 6290 8208 6346
rect 7868 6204 8208 6290
rect 7868 6148 7940 6204
rect 7996 6148 8082 6204
rect 8138 6148 8208 6204
rect 7868 6062 8208 6148
rect 7868 6006 7940 6062
rect 7996 6006 8082 6062
rect 8138 6006 8208 6062
rect 7868 5920 8208 6006
rect 7868 5864 7940 5920
rect 7996 5864 8082 5920
rect 8138 5864 8208 5920
rect 7868 5778 8208 5864
rect 7868 5722 7940 5778
rect 7996 5722 8082 5778
rect 8138 5722 8208 5778
rect 7868 5636 8208 5722
rect 7868 5580 7940 5636
rect 7996 5580 8082 5636
rect 8138 5580 8208 5636
rect 7868 5494 8208 5580
rect 7868 5438 7940 5494
rect 7996 5438 8082 5494
rect 8138 5438 8208 5494
rect 7868 5352 8208 5438
rect 7868 5296 7940 5352
rect 7996 5296 8082 5352
rect 8138 5296 8208 5352
rect 7868 5210 8208 5296
rect 7868 5154 7940 5210
rect 7996 5154 8082 5210
rect 8138 5154 8208 5210
rect 7868 5068 8208 5154
rect 7868 5012 7940 5068
rect 7996 5012 8082 5068
rect 8138 5012 8208 5068
rect 7868 4926 8208 5012
rect 7868 4870 7940 4926
rect 7996 4870 8082 4926
rect 8138 4870 8208 4926
rect 7868 4784 8208 4870
rect 7868 4728 7940 4784
rect 7996 4728 8082 4784
rect 8138 4728 8208 4784
rect 7868 4642 8208 4728
rect 7868 4586 7940 4642
rect 7996 4586 8082 4642
rect 8138 4586 8208 4642
rect 7868 4500 8208 4586
rect 7868 4444 7940 4500
rect 7996 4444 8082 4500
rect 8138 4444 8208 4500
rect 7868 4358 8208 4444
rect 7868 4302 7940 4358
rect 7996 4302 8082 4358
rect 8138 4302 8208 4358
rect 7868 4216 8208 4302
rect 7868 4160 7940 4216
rect 7996 4160 8082 4216
rect 8138 4160 8208 4216
rect 7868 4074 8208 4160
rect 7868 4018 7940 4074
rect 7996 4018 8082 4074
rect 8138 4018 8208 4074
rect 7868 3932 8208 4018
rect 7868 3876 7940 3932
rect 7996 3876 8082 3932
rect 8138 3876 8208 3932
rect 7868 3790 8208 3876
rect 7868 3734 7940 3790
rect 7996 3734 8082 3790
rect 8138 3734 8208 3790
rect 7868 3648 8208 3734
rect 7868 3592 7940 3648
rect 7996 3592 8082 3648
rect 8138 3592 8208 3648
rect 7868 3506 8208 3592
rect 7868 3450 7940 3506
rect 7996 3450 8082 3506
rect 8138 3450 8208 3506
rect 7868 3364 8208 3450
rect 7868 3308 7940 3364
rect 7996 3308 8082 3364
rect 8138 3308 8208 3364
rect 7868 3222 8208 3308
rect 7868 3166 7940 3222
rect 7996 3166 8082 3222
rect 8138 3166 8208 3222
rect 7868 3080 8208 3166
rect 7868 3024 7940 3080
rect 7996 3024 8082 3080
rect 8138 3024 8208 3080
rect 7868 2938 8208 3024
rect 7868 2882 7940 2938
rect 7996 2882 8082 2938
rect 8138 2882 8208 2938
rect 7868 2796 8208 2882
rect 7868 2740 7940 2796
rect 7996 2740 8082 2796
rect 8138 2740 8208 2796
rect 7868 2654 8208 2740
rect 7868 2598 7940 2654
rect 7996 2598 8082 2654
rect 8138 2598 8208 2654
rect 7868 2512 8208 2598
rect 7868 2456 7940 2512
rect 7996 2456 8082 2512
rect 8138 2456 8208 2512
rect 7868 2370 8208 2456
rect 7868 2314 7940 2370
rect 7996 2314 8082 2370
rect 8138 2314 8208 2370
rect 7868 2228 8208 2314
rect 7868 2172 7940 2228
rect 7996 2172 8082 2228
rect 8138 2172 8208 2228
rect 7868 2086 8208 2172
rect 7868 2030 7940 2086
rect 7996 2030 8082 2086
rect 8138 2030 8208 2086
rect 7868 1944 8208 2030
rect 7868 1888 7940 1944
rect 7996 1888 8082 1944
rect 8138 1888 8208 1944
rect 7868 1802 8208 1888
rect 7868 1746 7940 1802
rect 7996 1746 8082 1802
rect 8138 1746 8208 1802
rect 7868 1660 8208 1746
rect 7868 1604 7940 1660
rect 7996 1604 8082 1660
rect 8138 1604 8208 1660
rect 7868 1518 8208 1604
rect 7868 1462 7940 1518
rect 7996 1462 8082 1518
rect 8138 1462 8208 1518
rect 7868 1376 8208 1462
rect 7868 1320 7940 1376
rect 7996 1320 8082 1376
rect 8138 1320 8208 1376
rect 7868 1234 8208 1320
rect 7868 1178 7940 1234
rect 7996 1178 8082 1234
rect 8138 1178 8208 1234
rect 7868 1092 8208 1178
rect 7868 1036 7940 1092
rect 7996 1036 8082 1092
rect 8138 1036 8208 1092
rect 7868 950 8208 1036
rect 7868 894 7940 950
rect 7996 894 8082 950
rect 8138 894 8208 950
rect 7868 808 8208 894
rect 7868 752 7940 808
rect 7996 752 8082 808
rect 8138 752 8208 808
rect 7868 666 8208 752
rect 7868 610 7940 666
rect 7996 610 8082 666
rect 8138 610 8208 666
rect 7868 524 8208 610
rect 7868 468 7940 524
rect 7996 468 8082 524
rect 8138 468 8208 524
rect 7868 400 8208 468
rect 8268 12310 8608 12400
rect 8268 12254 8340 12310
rect 8396 12254 8482 12310
rect 8538 12254 8608 12310
rect 8268 12168 8608 12254
rect 8268 12112 8340 12168
rect 8396 12112 8482 12168
rect 8538 12112 8608 12168
rect 8268 12026 8608 12112
rect 8268 11970 8340 12026
rect 8396 11970 8482 12026
rect 8538 11970 8608 12026
rect 8268 11884 8608 11970
rect 8268 11828 8340 11884
rect 8396 11828 8482 11884
rect 8538 11828 8608 11884
rect 8268 11742 8608 11828
rect 8268 11686 8340 11742
rect 8396 11686 8482 11742
rect 8538 11686 8608 11742
rect 8268 11600 8608 11686
rect 8268 11544 8340 11600
rect 8396 11544 8482 11600
rect 8538 11544 8608 11600
rect 8268 11458 8608 11544
rect 8268 11402 8340 11458
rect 8396 11402 8482 11458
rect 8538 11402 8608 11458
rect 8268 11316 8608 11402
rect 8268 11260 8340 11316
rect 8396 11260 8482 11316
rect 8538 11260 8608 11316
rect 8268 11174 8608 11260
rect 8268 11118 8340 11174
rect 8396 11118 8482 11174
rect 8538 11118 8608 11174
rect 8268 11032 8608 11118
rect 8268 10976 8340 11032
rect 8396 10976 8482 11032
rect 8538 10976 8608 11032
rect 8268 10890 8608 10976
rect 8268 10834 8340 10890
rect 8396 10834 8482 10890
rect 8538 10834 8608 10890
rect 8268 10748 8608 10834
rect 8268 10692 8340 10748
rect 8396 10692 8482 10748
rect 8538 10692 8608 10748
rect 8268 10606 8608 10692
rect 8268 10550 8340 10606
rect 8396 10550 8482 10606
rect 8538 10550 8608 10606
rect 8268 10464 8608 10550
rect 8268 10408 8340 10464
rect 8396 10408 8482 10464
rect 8538 10408 8608 10464
rect 8268 10322 8608 10408
rect 8268 10266 8340 10322
rect 8396 10266 8482 10322
rect 8538 10266 8608 10322
rect 8268 10180 8608 10266
rect 8268 10124 8340 10180
rect 8396 10124 8482 10180
rect 8538 10124 8608 10180
rect 8268 10038 8608 10124
rect 8268 9982 8340 10038
rect 8396 9982 8482 10038
rect 8538 9982 8608 10038
rect 8268 9896 8608 9982
rect 8268 9840 8340 9896
rect 8396 9840 8482 9896
rect 8538 9840 8608 9896
rect 8268 9754 8608 9840
rect 8268 9698 8340 9754
rect 8396 9698 8482 9754
rect 8538 9698 8608 9754
rect 8268 9612 8608 9698
rect 8268 9556 8340 9612
rect 8396 9556 8482 9612
rect 8538 9556 8608 9612
rect 8268 9470 8608 9556
rect 8268 9414 8340 9470
rect 8396 9414 8482 9470
rect 8538 9414 8608 9470
rect 8268 9328 8608 9414
rect 8268 9272 8340 9328
rect 8396 9272 8482 9328
rect 8538 9272 8608 9328
rect 8268 9186 8608 9272
rect 8268 9130 8340 9186
rect 8396 9130 8482 9186
rect 8538 9130 8608 9186
rect 8268 9044 8608 9130
rect 8268 8988 8340 9044
rect 8396 8988 8482 9044
rect 8538 8988 8608 9044
rect 8268 8902 8608 8988
rect 8268 8846 8340 8902
rect 8396 8846 8482 8902
rect 8538 8846 8608 8902
rect 8268 8760 8608 8846
rect 8268 8704 8340 8760
rect 8396 8704 8482 8760
rect 8538 8704 8608 8760
rect 8268 8618 8608 8704
rect 8268 8562 8340 8618
rect 8396 8562 8482 8618
rect 8538 8562 8608 8618
rect 8268 8476 8608 8562
rect 8268 8420 8340 8476
rect 8396 8420 8482 8476
rect 8538 8420 8608 8476
rect 8268 8334 8608 8420
rect 8268 8278 8340 8334
rect 8396 8278 8482 8334
rect 8538 8278 8608 8334
rect 8268 8192 8608 8278
rect 8268 8136 8340 8192
rect 8396 8136 8482 8192
rect 8538 8136 8608 8192
rect 8268 8050 8608 8136
rect 8268 7994 8340 8050
rect 8396 7994 8482 8050
rect 8538 7994 8608 8050
rect 8268 7908 8608 7994
rect 8268 7852 8340 7908
rect 8396 7852 8482 7908
rect 8538 7852 8608 7908
rect 8268 7766 8608 7852
rect 8268 7710 8340 7766
rect 8396 7710 8482 7766
rect 8538 7710 8608 7766
rect 8268 7624 8608 7710
rect 8268 7568 8340 7624
rect 8396 7568 8482 7624
rect 8538 7568 8608 7624
rect 8268 7482 8608 7568
rect 8268 7426 8340 7482
rect 8396 7426 8482 7482
rect 8538 7426 8608 7482
rect 8268 7340 8608 7426
rect 8268 7284 8340 7340
rect 8396 7284 8482 7340
rect 8538 7284 8608 7340
rect 8268 7198 8608 7284
rect 8268 7142 8340 7198
rect 8396 7142 8482 7198
rect 8538 7142 8608 7198
rect 8268 7056 8608 7142
rect 8268 7000 8340 7056
rect 8396 7000 8482 7056
rect 8538 7000 8608 7056
rect 8268 6914 8608 7000
rect 8268 6858 8340 6914
rect 8396 6858 8482 6914
rect 8538 6858 8608 6914
rect 8268 6772 8608 6858
rect 8268 6716 8340 6772
rect 8396 6716 8482 6772
rect 8538 6716 8608 6772
rect 8268 6630 8608 6716
rect 8268 6574 8340 6630
rect 8396 6574 8482 6630
rect 8538 6574 8608 6630
rect 8268 6488 8608 6574
rect 8268 6432 8340 6488
rect 8396 6432 8482 6488
rect 8538 6432 8608 6488
rect 8268 6346 8608 6432
rect 8268 6290 8340 6346
rect 8396 6290 8482 6346
rect 8538 6290 8608 6346
rect 8268 6204 8608 6290
rect 8268 6148 8340 6204
rect 8396 6148 8482 6204
rect 8538 6148 8608 6204
rect 8268 6062 8608 6148
rect 8268 6006 8340 6062
rect 8396 6006 8482 6062
rect 8538 6006 8608 6062
rect 8268 5920 8608 6006
rect 8268 5864 8340 5920
rect 8396 5864 8482 5920
rect 8538 5864 8608 5920
rect 8268 5778 8608 5864
rect 8268 5722 8340 5778
rect 8396 5722 8482 5778
rect 8538 5722 8608 5778
rect 8268 5636 8608 5722
rect 8268 5580 8340 5636
rect 8396 5580 8482 5636
rect 8538 5580 8608 5636
rect 8268 5494 8608 5580
rect 8268 5438 8340 5494
rect 8396 5438 8482 5494
rect 8538 5438 8608 5494
rect 8268 5352 8608 5438
rect 8268 5296 8340 5352
rect 8396 5296 8482 5352
rect 8538 5296 8608 5352
rect 8268 5210 8608 5296
rect 8268 5154 8340 5210
rect 8396 5154 8482 5210
rect 8538 5154 8608 5210
rect 8268 5068 8608 5154
rect 8268 5012 8340 5068
rect 8396 5012 8482 5068
rect 8538 5012 8608 5068
rect 8268 4926 8608 5012
rect 8268 4870 8340 4926
rect 8396 4870 8482 4926
rect 8538 4870 8608 4926
rect 8268 4784 8608 4870
rect 8268 4728 8340 4784
rect 8396 4728 8482 4784
rect 8538 4728 8608 4784
rect 8268 4642 8608 4728
rect 8268 4586 8340 4642
rect 8396 4586 8482 4642
rect 8538 4586 8608 4642
rect 8268 4500 8608 4586
rect 8268 4444 8340 4500
rect 8396 4444 8482 4500
rect 8538 4444 8608 4500
rect 8268 4358 8608 4444
rect 8268 4302 8340 4358
rect 8396 4302 8482 4358
rect 8538 4302 8608 4358
rect 8268 4216 8608 4302
rect 8268 4160 8340 4216
rect 8396 4160 8482 4216
rect 8538 4160 8608 4216
rect 8268 4074 8608 4160
rect 8268 4018 8340 4074
rect 8396 4018 8482 4074
rect 8538 4018 8608 4074
rect 8268 3932 8608 4018
rect 8268 3876 8340 3932
rect 8396 3876 8482 3932
rect 8538 3876 8608 3932
rect 8268 3790 8608 3876
rect 8268 3734 8340 3790
rect 8396 3734 8482 3790
rect 8538 3734 8608 3790
rect 8268 3648 8608 3734
rect 8268 3592 8340 3648
rect 8396 3592 8482 3648
rect 8538 3592 8608 3648
rect 8268 3506 8608 3592
rect 8268 3450 8340 3506
rect 8396 3450 8482 3506
rect 8538 3450 8608 3506
rect 8268 3364 8608 3450
rect 8268 3308 8340 3364
rect 8396 3308 8482 3364
rect 8538 3308 8608 3364
rect 8268 3222 8608 3308
rect 8268 3166 8340 3222
rect 8396 3166 8482 3222
rect 8538 3166 8608 3222
rect 8268 3080 8608 3166
rect 8268 3024 8340 3080
rect 8396 3024 8482 3080
rect 8538 3024 8608 3080
rect 8268 2938 8608 3024
rect 8268 2882 8340 2938
rect 8396 2882 8482 2938
rect 8538 2882 8608 2938
rect 8268 2796 8608 2882
rect 8268 2740 8340 2796
rect 8396 2740 8482 2796
rect 8538 2740 8608 2796
rect 8268 2654 8608 2740
rect 8268 2598 8340 2654
rect 8396 2598 8482 2654
rect 8538 2598 8608 2654
rect 8268 2512 8608 2598
rect 8268 2456 8340 2512
rect 8396 2456 8482 2512
rect 8538 2456 8608 2512
rect 8268 2370 8608 2456
rect 8268 2314 8340 2370
rect 8396 2314 8482 2370
rect 8538 2314 8608 2370
rect 8268 2228 8608 2314
rect 8268 2172 8340 2228
rect 8396 2172 8482 2228
rect 8538 2172 8608 2228
rect 8268 2086 8608 2172
rect 8268 2030 8340 2086
rect 8396 2030 8482 2086
rect 8538 2030 8608 2086
rect 8268 1944 8608 2030
rect 8268 1888 8340 1944
rect 8396 1888 8482 1944
rect 8538 1888 8608 1944
rect 8268 1802 8608 1888
rect 8268 1746 8340 1802
rect 8396 1746 8482 1802
rect 8538 1746 8608 1802
rect 8268 1660 8608 1746
rect 8268 1604 8340 1660
rect 8396 1604 8482 1660
rect 8538 1604 8608 1660
rect 8268 1518 8608 1604
rect 8268 1462 8340 1518
rect 8396 1462 8482 1518
rect 8538 1462 8608 1518
rect 8268 1376 8608 1462
rect 8268 1320 8340 1376
rect 8396 1320 8482 1376
rect 8538 1320 8608 1376
rect 8268 1234 8608 1320
rect 8268 1178 8340 1234
rect 8396 1178 8482 1234
rect 8538 1178 8608 1234
rect 8268 1092 8608 1178
rect 8268 1036 8340 1092
rect 8396 1036 8482 1092
rect 8538 1036 8608 1092
rect 8268 950 8608 1036
rect 8268 894 8340 950
rect 8396 894 8482 950
rect 8538 894 8608 950
rect 8268 808 8608 894
rect 8268 752 8340 808
rect 8396 752 8482 808
rect 8538 752 8608 808
rect 8268 666 8608 752
rect 8268 610 8340 666
rect 8396 610 8482 666
rect 8538 610 8608 666
rect 8268 524 8608 610
rect 8268 468 8340 524
rect 8396 468 8482 524
rect 8538 468 8608 524
rect 8268 400 8608 468
rect 8668 12310 9008 12400
rect 8668 12254 8737 12310
rect 8793 12254 8879 12310
rect 8935 12254 9008 12310
rect 8668 12168 9008 12254
rect 8668 12112 8737 12168
rect 8793 12112 8879 12168
rect 8935 12112 9008 12168
rect 8668 12026 9008 12112
rect 8668 11970 8737 12026
rect 8793 11970 8879 12026
rect 8935 11970 9008 12026
rect 8668 11884 9008 11970
rect 8668 11828 8737 11884
rect 8793 11828 8879 11884
rect 8935 11828 9008 11884
rect 8668 11742 9008 11828
rect 8668 11686 8737 11742
rect 8793 11686 8879 11742
rect 8935 11686 9008 11742
rect 8668 11600 9008 11686
rect 8668 11544 8737 11600
rect 8793 11544 8879 11600
rect 8935 11544 9008 11600
rect 8668 11458 9008 11544
rect 8668 11402 8737 11458
rect 8793 11402 8879 11458
rect 8935 11402 9008 11458
rect 8668 11316 9008 11402
rect 8668 11260 8737 11316
rect 8793 11260 8879 11316
rect 8935 11260 9008 11316
rect 8668 11174 9008 11260
rect 8668 11118 8737 11174
rect 8793 11118 8879 11174
rect 8935 11118 9008 11174
rect 8668 11032 9008 11118
rect 8668 10976 8737 11032
rect 8793 10976 8879 11032
rect 8935 10976 9008 11032
rect 8668 10890 9008 10976
rect 8668 10834 8737 10890
rect 8793 10834 8879 10890
rect 8935 10834 9008 10890
rect 8668 10748 9008 10834
rect 8668 10692 8737 10748
rect 8793 10692 8879 10748
rect 8935 10692 9008 10748
rect 8668 10606 9008 10692
rect 8668 10550 8737 10606
rect 8793 10550 8879 10606
rect 8935 10550 9008 10606
rect 8668 10464 9008 10550
rect 8668 10408 8737 10464
rect 8793 10408 8879 10464
rect 8935 10408 9008 10464
rect 8668 10322 9008 10408
rect 8668 10266 8737 10322
rect 8793 10266 8879 10322
rect 8935 10266 9008 10322
rect 8668 10180 9008 10266
rect 8668 10124 8737 10180
rect 8793 10124 8879 10180
rect 8935 10124 9008 10180
rect 8668 10038 9008 10124
rect 8668 9982 8737 10038
rect 8793 9982 8879 10038
rect 8935 9982 9008 10038
rect 8668 9896 9008 9982
rect 8668 9840 8737 9896
rect 8793 9840 8879 9896
rect 8935 9840 9008 9896
rect 8668 9754 9008 9840
rect 8668 9698 8737 9754
rect 8793 9698 8879 9754
rect 8935 9698 9008 9754
rect 8668 9612 9008 9698
rect 8668 9556 8737 9612
rect 8793 9556 8879 9612
rect 8935 9556 9008 9612
rect 8668 9470 9008 9556
rect 8668 9414 8737 9470
rect 8793 9414 8879 9470
rect 8935 9414 9008 9470
rect 8668 9328 9008 9414
rect 8668 9272 8737 9328
rect 8793 9272 8879 9328
rect 8935 9272 9008 9328
rect 8668 9186 9008 9272
rect 8668 9130 8737 9186
rect 8793 9130 8879 9186
rect 8935 9130 9008 9186
rect 8668 9044 9008 9130
rect 8668 8988 8737 9044
rect 8793 8988 8879 9044
rect 8935 8988 9008 9044
rect 8668 8902 9008 8988
rect 8668 8846 8737 8902
rect 8793 8846 8879 8902
rect 8935 8846 9008 8902
rect 8668 8760 9008 8846
rect 8668 8704 8737 8760
rect 8793 8704 8879 8760
rect 8935 8704 9008 8760
rect 8668 8618 9008 8704
rect 8668 8562 8737 8618
rect 8793 8562 8879 8618
rect 8935 8562 9008 8618
rect 8668 8476 9008 8562
rect 8668 8420 8737 8476
rect 8793 8420 8879 8476
rect 8935 8420 9008 8476
rect 8668 8334 9008 8420
rect 8668 8278 8737 8334
rect 8793 8278 8879 8334
rect 8935 8278 9008 8334
rect 8668 8192 9008 8278
rect 8668 8136 8737 8192
rect 8793 8136 8879 8192
rect 8935 8136 9008 8192
rect 8668 8050 9008 8136
rect 8668 7994 8737 8050
rect 8793 7994 8879 8050
rect 8935 7994 9008 8050
rect 8668 7908 9008 7994
rect 8668 7852 8737 7908
rect 8793 7852 8879 7908
rect 8935 7852 9008 7908
rect 8668 7766 9008 7852
rect 8668 7710 8737 7766
rect 8793 7710 8879 7766
rect 8935 7710 9008 7766
rect 8668 7624 9008 7710
rect 8668 7568 8737 7624
rect 8793 7568 8879 7624
rect 8935 7568 9008 7624
rect 8668 7482 9008 7568
rect 8668 7426 8737 7482
rect 8793 7426 8879 7482
rect 8935 7426 9008 7482
rect 8668 7340 9008 7426
rect 8668 7284 8737 7340
rect 8793 7284 8879 7340
rect 8935 7284 9008 7340
rect 8668 7198 9008 7284
rect 8668 7142 8737 7198
rect 8793 7142 8879 7198
rect 8935 7142 9008 7198
rect 8668 7056 9008 7142
rect 8668 7000 8737 7056
rect 8793 7000 8879 7056
rect 8935 7000 9008 7056
rect 8668 6914 9008 7000
rect 8668 6858 8737 6914
rect 8793 6858 8879 6914
rect 8935 6858 9008 6914
rect 8668 6772 9008 6858
rect 8668 6716 8737 6772
rect 8793 6716 8879 6772
rect 8935 6716 9008 6772
rect 8668 6630 9008 6716
rect 8668 6574 8737 6630
rect 8793 6574 8879 6630
rect 8935 6574 9008 6630
rect 8668 6488 9008 6574
rect 8668 6432 8737 6488
rect 8793 6432 8879 6488
rect 8935 6432 9008 6488
rect 8668 6346 9008 6432
rect 8668 6290 8737 6346
rect 8793 6290 8879 6346
rect 8935 6290 9008 6346
rect 8668 6204 9008 6290
rect 8668 6148 8737 6204
rect 8793 6148 8879 6204
rect 8935 6148 9008 6204
rect 8668 6062 9008 6148
rect 8668 6006 8737 6062
rect 8793 6006 8879 6062
rect 8935 6006 9008 6062
rect 8668 5920 9008 6006
rect 8668 5864 8737 5920
rect 8793 5864 8879 5920
rect 8935 5864 9008 5920
rect 8668 5778 9008 5864
rect 8668 5722 8737 5778
rect 8793 5722 8879 5778
rect 8935 5722 9008 5778
rect 8668 5636 9008 5722
rect 8668 5580 8737 5636
rect 8793 5580 8879 5636
rect 8935 5580 9008 5636
rect 8668 5494 9008 5580
rect 8668 5438 8737 5494
rect 8793 5438 8879 5494
rect 8935 5438 9008 5494
rect 8668 5352 9008 5438
rect 8668 5296 8737 5352
rect 8793 5296 8879 5352
rect 8935 5296 9008 5352
rect 8668 5210 9008 5296
rect 8668 5154 8737 5210
rect 8793 5154 8879 5210
rect 8935 5154 9008 5210
rect 8668 5068 9008 5154
rect 8668 5012 8737 5068
rect 8793 5012 8879 5068
rect 8935 5012 9008 5068
rect 8668 4926 9008 5012
rect 8668 4870 8737 4926
rect 8793 4870 8879 4926
rect 8935 4870 9008 4926
rect 8668 4784 9008 4870
rect 8668 4728 8737 4784
rect 8793 4728 8879 4784
rect 8935 4728 9008 4784
rect 8668 4642 9008 4728
rect 8668 4586 8737 4642
rect 8793 4586 8879 4642
rect 8935 4586 9008 4642
rect 8668 4500 9008 4586
rect 8668 4444 8737 4500
rect 8793 4444 8879 4500
rect 8935 4444 9008 4500
rect 8668 4358 9008 4444
rect 8668 4302 8737 4358
rect 8793 4302 8879 4358
rect 8935 4302 9008 4358
rect 8668 4216 9008 4302
rect 8668 4160 8737 4216
rect 8793 4160 8879 4216
rect 8935 4160 9008 4216
rect 8668 4074 9008 4160
rect 8668 4018 8737 4074
rect 8793 4018 8879 4074
rect 8935 4018 9008 4074
rect 8668 3932 9008 4018
rect 8668 3876 8737 3932
rect 8793 3876 8879 3932
rect 8935 3876 9008 3932
rect 8668 3790 9008 3876
rect 8668 3734 8737 3790
rect 8793 3734 8879 3790
rect 8935 3734 9008 3790
rect 8668 3648 9008 3734
rect 8668 3592 8737 3648
rect 8793 3592 8879 3648
rect 8935 3592 9008 3648
rect 8668 3506 9008 3592
rect 8668 3450 8737 3506
rect 8793 3450 8879 3506
rect 8935 3450 9008 3506
rect 8668 3364 9008 3450
rect 8668 3308 8737 3364
rect 8793 3308 8879 3364
rect 8935 3308 9008 3364
rect 8668 3222 9008 3308
rect 8668 3166 8737 3222
rect 8793 3166 8879 3222
rect 8935 3166 9008 3222
rect 8668 3080 9008 3166
rect 8668 3024 8737 3080
rect 8793 3024 8879 3080
rect 8935 3024 9008 3080
rect 8668 2938 9008 3024
rect 8668 2882 8737 2938
rect 8793 2882 8879 2938
rect 8935 2882 9008 2938
rect 8668 2796 9008 2882
rect 8668 2740 8737 2796
rect 8793 2740 8879 2796
rect 8935 2740 9008 2796
rect 8668 2654 9008 2740
rect 8668 2598 8737 2654
rect 8793 2598 8879 2654
rect 8935 2598 9008 2654
rect 8668 2512 9008 2598
rect 8668 2456 8737 2512
rect 8793 2456 8879 2512
rect 8935 2456 9008 2512
rect 8668 2370 9008 2456
rect 8668 2314 8737 2370
rect 8793 2314 8879 2370
rect 8935 2314 9008 2370
rect 8668 2228 9008 2314
rect 8668 2172 8737 2228
rect 8793 2172 8879 2228
rect 8935 2172 9008 2228
rect 8668 2086 9008 2172
rect 8668 2030 8737 2086
rect 8793 2030 8879 2086
rect 8935 2030 9008 2086
rect 8668 1944 9008 2030
rect 8668 1888 8737 1944
rect 8793 1888 8879 1944
rect 8935 1888 9008 1944
rect 8668 1802 9008 1888
rect 8668 1746 8737 1802
rect 8793 1746 8879 1802
rect 8935 1746 9008 1802
rect 8668 1660 9008 1746
rect 8668 1604 8737 1660
rect 8793 1604 8879 1660
rect 8935 1604 9008 1660
rect 8668 1518 9008 1604
rect 8668 1462 8737 1518
rect 8793 1462 8879 1518
rect 8935 1462 9008 1518
rect 8668 1376 9008 1462
rect 8668 1320 8737 1376
rect 8793 1320 8879 1376
rect 8935 1320 9008 1376
rect 8668 1234 9008 1320
rect 8668 1178 8737 1234
rect 8793 1178 8879 1234
rect 8935 1178 9008 1234
rect 8668 1092 9008 1178
rect 8668 1036 8737 1092
rect 8793 1036 8879 1092
rect 8935 1036 9008 1092
rect 8668 950 9008 1036
rect 8668 894 8737 950
rect 8793 894 8879 950
rect 8935 894 9008 950
rect 8668 808 9008 894
rect 8668 752 8737 808
rect 8793 752 8879 808
rect 8935 752 9008 808
rect 8668 666 9008 752
rect 8668 610 8737 666
rect 8793 610 8879 666
rect 8935 610 9008 666
rect 8668 524 9008 610
rect 8668 468 8737 524
rect 8793 468 8879 524
rect 8935 468 9008 524
rect 8668 400 9008 468
rect 9068 12310 9408 12400
rect 9068 12254 9134 12310
rect 9190 12254 9276 12310
rect 9332 12254 9408 12310
rect 9068 12168 9408 12254
rect 9068 12112 9134 12168
rect 9190 12112 9276 12168
rect 9332 12112 9408 12168
rect 9068 12026 9408 12112
rect 9068 11970 9134 12026
rect 9190 11970 9276 12026
rect 9332 11970 9408 12026
rect 9068 11884 9408 11970
rect 9068 11828 9134 11884
rect 9190 11828 9276 11884
rect 9332 11828 9408 11884
rect 9068 11742 9408 11828
rect 9068 11686 9134 11742
rect 9190 11686 9276 11742
rect 9332 11686 9408 11742
rect 9068 11600 9408 11686
rect 9068 11544 9134 11600
rect 9190 11544 9276 11600
rect 9332 11544 9408 11600
rect 9068 11458 9408 11544
rect 9068 11402 9134 11458
rect 9190 11402 9276 11458
rect 9332 11402 9408 11458
rect 9068 11316 9408 11402
rect 9068 11260 9134 11316
rect 9190 11260 9276 11316
rect 9332 11260 9408 11316
rect 9068 11174 9408 11260
rect 9068 11118 9134 11174
rect 9190 11118 9276 11174
rect 9332 11118 9408 11174
rect 9068 11032 9408 11118
rect 9068 10976 9134 11032
rect 9190 10976 9276 11032
rect 9332 10976 9408 11032
rect 9068 10890 9408 10976
rect 9068 10834 9134 10890
rect 9190 10834 9276 10890
rect 9332 10834 9408 10890
rect 9068 10748 9408 10834
rect 9068 10692 9134 10748
rect 9190 10692 9276 10748
rect 9332 10692 9408 10748
rect 9068 10606 9408 10692
rect 9068 10550 9134 10606
rect 9190 10550 9276 10606
rect 9332 10550 9408 10606
rect 9068 10464 9408 10550
rect 9068 10408 9134 10464
rect 9190 10408 9276 10464
rect 9332 10408 9408 10464
rect 9068 10322 9408 10408
rect 9068 10266 9134 10322
rect 9190 10266 9276 10322
rect 9332 10266 9408 10322
rect 9068 10180 9408 10266
rect 9068 10124 9134 10180
rect 9190 10124 9276 10180
rect 9332 10124 9408 10180
rect 9068 10038 9408 10124
rect 9068 9982 9134 10038
rect 9190 9982 9276 10038
rect 9332 9982 9408 10038
rect 9068 9896 9408 9982
rect 9068 9840 9134 9896
rect 9190 9840 9276 9896
rect 9332 9840 9408 9896
rect 9068 9754 9408 9840
rect 9068 9698 9134 9754
rect 9190 9698 9276 9754
rect 9332 9698 9408 9754
rect 9068 9612 9408 9698
rect 9068 9556 9134 9612
rect 9190 9556 9276 9612
rect 9332 9556 9408 9612
rect 9068 9470 9408 9556
rect 9068 9414 9134 9470
rect 9190 9414 9276 9470
rect 9332 9414 9408 9470
rect 9068 9328 9408 9414
rect 9068 9272 9134 9328
rect 9190 9272 9276 9328
rect 9332 9272 9408 9328
rect 9068 9186 9408 9272
rect 9068 9130 9134 9186
rect 9190 9130 9276 9186
rect 9332 9130 9408 9186
rect 9068 9044 9408 9130
rect 9068 8988 9134 9044
rect 9190 8988 9276 9044
rect 9332 8988 9408 9044
rect 9068 8902 9408 8988
rect 9068 8846 9134 8902
rect 9190 8846 9276 8902
rect 9332 8846 9408 8902
rect 9068 8760 9408 8846
rect 9068 8704 9134 8760
rect 9190 8704 9276 8760
rect 9332 8704 9408 8760
rect 9068 8618 9408 8704
rect 9068 8562 9134 8618
rect 9190 8562 9276 8618
rect 9332 8562 9408 8618
rect 9068 8476 9408 8562
rect 9068 8420 9134 8476
rect 9190 8420 9276 8476
rect 9332 8420 9408 8476
rect 9068 8334 9408 8420
rect 9068 8278 9134 8334
rect 9190 8278 9276 8334
rect 9332 8278 9408 8334
rect 9068 8192 9408 8278
rect 9068 8136 9134 8192
rect 9190 8136 9276 8192
rect 9332 8136 9408 8192
rect 9068 8050 9408 8136
rect 9068 7994 9134 8050
rect 9190 7994 9276 8050
rect 9332 7994 9408 8050
rect 9068 7908 9408 7994
rect 9068 7852 9134 7908
rect 9190 7852 9276 7908
rect 9332 7852 9408 7908
rect 9068 7766 9408 7852
rect 9068 7710 9134 7766
rect 9190 7710 9276 7766
rect 9332 7710 9408 7766
rect 9068 7624 9408 7710
rect 9068 7568 9134 7624
rect 9190 7568 9276 7624
rect 9332 7568 9408 7624
rect 9068 7482 9408 7568
rect 9068 7426 9134 7482
rect 9190 7426 9276 7482
rect 9332 7426 9408 7482
rect 9068 7340 9408 7426
rect 9068 7284 9134 7340
rect 9190 7284 9276 7340
rect 9332 7284 9408 7340
rect 9068 7198 9408 7284
rect 9068 7142 9134 7198
rect 9190 7142 9276 7198
rect 9332 7142 9408 7198
rect 9068 7056 9408 7142
rect 9068 7000 9134 7056
rect 9190 7000 9276 7056
rect 9332 7000 9408 7056
rect 9068 6914 9408 7000
rect 9068 6858 9134 6914
rect 9190 6858 9276 6914
rect 9332 6858 9408 6914
rect 9068 6772 9408 6858
rect 9068 6716 9134 6772
rect 9190 6716 9276 6772
rect 9332 6716 9408 6772
rect 9068 6630 9408 6716
rect 9068 6574 9134 6630
rect 9190 6574 9276 6630
rect 9332 6574 9408 6630
rect 9068 6488 9408 6574
rect 9068 6432 9134 6488
rect 9190 6432 9276 6488
rect 9332 6432 9408 6488
rect 9068 6346 9408 6432
rect 9068 6290 9134 6346
rect 9190 6290 9276 6346
rect 9332 6290 9408 6346
rect 9068 6204 9408 6290
rect 9068 6148 9134 6204
rect 9190 6148 9276 6204
rect 9332 6148 9408 6204
rect 9068 6062 9408 6148
rect 9068 6006 9134 6062
rect 9190 6006 9276 6062
rect 9332 6006 9408 6062
rect 9068 5920 9408 6006
rect 9068 5864 9134 5920
rect 9190 5864 9276 5920
rect 9332 5864 9408 5920
rect 9068 5778 9408 5864
rect 9068 5722 9134 5778
rect 9190 5722 9276 5778
rect 9332 5722 9408 5778
rect 9068 5636 9408 5722
rect 9068 5580 9134 5636
rect 9190 5580 9276 5636
rect 9332 5580 9408 5636
rect 9068 5494 9408 5580
rect 9068 5438 9134 5494
rect 9190 5438 9276 5494
rect 9332 5438 9408 5494
rect 9068 5352 9408 5438
rect 9068 5296 9134 5352
rect 9190 5296 9276 5352
rect 9332 5296 9408 5352
rect 9068 5210 9408 5296
rect 9068 5154 9134 5210
rect 9190 5154 9276 5210
rect 9332 5154 9408 5210
rect 9068 5068 9408 5154
rect 9068 5012 9134 5068
rect 9190 5012 9276 5068
rect 9332 5012 9408 5068
rect 9068 4926 9408 5012
rect 9068 4870 9134 4926
rect 9190 4870 9276 4926
rect 9332 4870 9408 4926
rect 9068 4784 9408 4870
rect 9068 4728 9134 4784
rect 9190 4728 9276 4784
rect 9332 4728 9408 4784
rect 9068 4642 9408 4728
rect 9068 4586 9134 4642
rect 9190 4586 9276 4642
rect 9332 4586 9408 4642
rect 9068 4500 9408 4586
rect 9068 4444 9134 4500
rect 9190 4444 9276 4500
rect 9332 4444 9408 4500
rect 9068 4358 9408 4444
rect 9068 4302 9134 4358
rect 9190 4302 9276 4358
rect 9332 4302 9408 4358
rect 9068 4216 9408 4302
rect 9068 4160 9134 4216
rect 9190 4160 9276 4216
rect 9332 4160 9408 4216
rect 9068 4074 9408 4160
rect 9068 4018 9134 4074
rect 9190 4018 9276 4074
rect 9332 4018 9408 4074
rect 9068 3932 9408 4018
rect 9068 3876 9134 3932
rect 9190 3876 9276 3932
rect 9332 3876 9408 3932
rect 9068 3790 9408 3876
rect 9068 3734 9134 3790
rect 9190 3734 9276 3790
rect 9332 3734 9408 3790
rect 9068 3648 9408 3734
rect 9068 3592 9134 3648
rect 9190 3592 9276 3648
rect 9332 3592 9408 3648
rect 9068 3506 9408 3592
rect 9068 3450 9134 3506
rect 9190 3450 9276 3506
rect 9332 3450 9408 3506
rect 9068 3364 9408 3450
rect 9068 3308 9134 3364
rect 9190 3308 9276 3364
rect 9332 3308 9408 3364
rect 9068 3222 9408 3308
rect 9068 3166 9134 3222
rect 9190 3166 9276 3222
rect 9332 3166 9408 3222
rect 9068 3080 9408 3166
rect 9068 3024 9134 3080
rect 9190 3024 9276 3080
rect 9332 3024 9408 3080
rect 9068 2938 9408 3024
rect 9068 2882 9134 2938
rect 9190 2882 9276 2938
rect 9332 2882 9408 2938
rect 9068 2796 9408 2882
rect 9068 2740 9134 2796
rect 9190 2740 9276 2796
rect 9332 2740 9408 2796
rect 9068 2654 9408 2740
rect 9068 2598 9134 2654
rect 9190 2598 9276 2654
rect 9332 2598 9408 2654
rect 9068 2512 9408 2598
rect 9068 2456 9134 2512
rect 9190 2456 9276 2512
rect 9332 2456 9408 2512
rect 9068 2370 9408 2456
rect 9068 2314 9134 2370
rect 9190 2314 9276 2370
rect 9332 2314 9408 2370
rect 9068 2228 9408 2314
rect 9068 2172 9134 2228
rect 9190 2172 9276 2228
rect 9332 2172 9408 2228
rect 9068 2086 9408 2172
rect 9068 2030 9134 2086
rect 9190 2030 9276 2086
rect 9332 2030 9408 2086
rect 9068 1944 9408 2030
rect 9068 1888 9134 1944
rect 9190 1888 9276 1944
rect 9332 1888 9408 1944
rect 9068 1802 9408 1888
rect 9068 1746 9134 1802
rect 9190 1746 9276 1802
rect 9332 1746 9408 1802
rect 9068 1660 9408 1746
rect 9068 1604 9134 1660
rect 9190 1604 9276 1660
rect 9332 1604 9408 1660
rect 9068 1518 9408 1604
rect 9068 1462 9134 1518
rect 9190 1462 9276 1518
rect 9332 1462 9408 1518
rect 9068 1376 9408 1462
rect 9068 1320 9134 1376
rect 9190 1320 9276 1376
rect 9332 1320 9408 1376
rect 9068 1234 9408 1320
rect 9068 1178 9134 1234
rect 9190 1178 9276 1234
rect 9332 1178 9408 1234
rect 9068 1092 9408 1178
rect 9068 1036 9134 1092
rect 9190 1036 9276 1092
rect 9332 1036 9408 1092
rect 9068 950 9408 1036
rect 9068 894 9134 950
rect 9190 894 9276 950
rect 9332 894 9408 950
rect 9068 808 9408 894
rect 9068 752 9134 808
rect 9190 752 9276 808
rect 9332 752 9408 808
rect 9068 666 9408 752
rect 9068 610 9134 666
rect 9190 610 9276 666
rect 9332 610 9408 666
rect 9068 524 9408 610
rect 9068 468 9134 524
rect 9190 468 9276 524
rect 9332 468 9408 524
rect 9068 400 9408 468
rect 9468 12310 9808 12400
rect 9468 12254 9538 12310
rect 9594 12254 9680 12310
rect 9736 12254 9808 12310
rect 9468 12168 9808 12254
rect 9468 12112 9538 12168
rect 9594 12112 9680 12168
rect 9736 12112 9808 12168
rect 9468 12026 9808 12112
rect 9468 11970 9538 12026
rect 9594 11970 9680 12026
rect 9736 11970 9808 12026
rect 9468 11884 9808 11970
rect 9468 11828 9538 11884
rect 9594 11828 9680 11884
rect 9736 11828 9808 11884
rect 9468 11742 9808 11828
rect 9468 11686 9538 11742
rect 9594 11686 9680 11742
rect 9736 11686 9808 11742
rect 9468 11600 9808 11686
rect 9468 11544 9538 11600
rect 9594 11544 9680 11600
rect 9736 11544 9808 11600
rect 9468 11458 9808 11544
rect 9468 11402 9538 11458
rect 9594 11402 9680 11458
rect 9736 11402 9808 11458
rect 9468 11316 9808 11402
rect 9468 11260 9538 11316
rect 9594 11260 9680 11316
rect 9736 11260 9808 11316
rect 9468 11174 9808 11260
rect 9468 11118 9538 11174
rect 9594 11118 9680 11174
rect 9736 11118 9808 11174
rect 9468 11032 9808 11118
rect 9468 10976 9538 11032
rect 9594 10976 9680 11032
rect 9736 10976 9808 11032
rect 9468 10890 9808 10976
rect 9468 10834 9538 10890
rect 9594 10834 9680 10890
rect 9736 10834 9808 10890
rect 9468 10748 9808 10834
rect 9468 10692 9538 10748
rect 9594 10692 9680 10748
rect 9736 10692 9808 10748
rect 9468 10606 9808 10692
rect 9468 10550 9538 10606
rect 9594 10550 9680 10606
rect 9736 10550 9808 10606
rect 9468 10464 9808 10550
rect 9468 10408 9538 10464
rect 9594 10408 9680 10464
rect 9736 10408 9808 10464
rect 9468 10322 9808 10408
rect 9468 10266 9538 10322
rect 9594 10266 9680 10322
rect 9736 10266 9808 10322
rect 9468 10180 9808 10266
rect 9468 10124 9538 10180
rect 9594 10124 9680 10180
rect 9736 10124 9808 10180
rect 9468 10038 9808 10124
rect 9468 9982 9538 10038
rect 9594 9982 9680 10038
rect 9736 9982 9808 10038
rect 9468 9896 9808 9982
rect 9468 9840 9538 9896
rect 9594 9840 9680 9896
rect 9736 9840 9808 9896
rect 9468 9754 9808 9840
rect 9468 9698 9538 9754
rect 9594 9698 9680 9754
rect 9736 9698 9808 9754
rect 9468 9612 9808 9698
rect 9468 9556 9538 9612
rect 9594 9556 9680 9612
rect 9736 9556 9808 9612
rect 9468 9470 9808 9556
rect 9468 9414 9538 9470
rect 9594 9414 9680 9470
rect 9736 9414 9808 9470
rect 9468 9328 9808 9414
rect 9468 9272 9538 9328
rect 9594 9272 9680 9328
rect 9736 9272 9808 9328
rect 9468 9186 9808 9272
rect 9468 9130 9538 9186
rect 9594 9130 9680 9186
rect 9736 9130 9808 9186
rect 9468 9044 9808 9130
rect 9468 8988 9538 9044
rect 9594 8988 9680 9044
rect 9736 8988 9808 9044
rect 9468 8902 9808 8988
rect 9468 8846 9538 8902
rect 9594 8846 9680 8902
rect 9736 8846 9808 8902
rect 9468 8760 9808 8846
rect 9468 8704 9538 8760
rect 9594 8704 9680 8760
rect 9736 8704 9808 8760
rect 9468 8618 9808 8704
rect 9468 8562 9538 8618
rect 9594 8562 9680 8618
rect 9736 8562 9808 8618
rect 9468 8476 9808 8562
rect 9468 8420 9538 8476
rect 9594 8420 9680 8476
rect 9736 8420 9808 8476
rect 9468 8334 9808 8420
rect 9468 8278 9538 8334
rect 9594 8278 9680 8334
rect 9736 8278 9808 8334
rect 9468 8192 9808 8278
rect 9468 8136 9538 8192
rect 9594 8136 9680 8192
rect 9736 8136 9808 8192
rect 9468 8050 9808 8136
rect 9468 7994 9538 8050
rect 9594 7994 9680 8050
rect 9736 7994 9808 8050
rect 9468 7908 9808 7994
rect 9468 7852 9538 7908
rect 9594 7852 9680 7908
rect 9736 7852 9808 7908
rect 9468 7766 9808 7852
rect 9468 7710 9538 7766
rect 9594 7710 9680 7766
rect 9736 7710 9808 7766
rect 9468 7624 9808 7710
rect 9468 7568 9538 7624
rect 9594 7568 9680 7624
rect 9736 7568 9808 7624
rect 9468 7482 9808 7568
rect 9468 7426 9538 7482
rect 9594 7426 9680 7482
rect 9736 7426 9808 7482
rect 9468 7340 9808 7426
rect 9468 7284 9538 7340
rect 9594 7284 9680 7340
rect 9736 7284 9808 7340
rect 9468 7198 9808 7284
rect 9468 7142 9538 7198
rect 9594 7142 9680 7198
rect 9736 7142 9808 7198
rect 9468 7056 9808 7142
rect 9468 7000 9538 7056
rect 9594 7000 9680 7056
rect 9736 7000 9808 7056
rect 9468 6914 9808 7000
rect 9468 6858 9538 6914
rect 9594 6858 9680 6914
rect 9736 6858 9808 6914
rect 9468 6772 9808 6858
rect 9468 6716 9538 6772
rect 9594 6716 9680 6772
rect 9736 6716 9808 6772
rect 9468 6630 9808 6716
rect 9468 6574 9538 6630
rect 9594 6574 9680 6630
rect 9736 6574 9808 6630
rect 9468 6488 9808 6574
rect 9468 6432 9538 6488
rect 9594 6432 9680 6488
rect 9736 6432 9808 6488
rect 9468 6346 9808 6432
rect 9468 6290 9538 6346
rect 9594 6290 9680 6346
rect 9736 6290 9808 6346
rect 9468 6204 9808 6290
rect 9468 6148 9538 6204
rect 9594 6148 9680 6204
rect 9736 6148 9808 6204
rect 9468 6062 9808 6148
rect 9468 6006 9538 6062
rect 9594 6006 9680 6062
rect 9736 6006 9808 6062
rect 9468 5920 9808 6006
rect 9468 5864 9538 5920
rect 9594 5864 9680 5920
rect 9736 5864 9808 5920
rect 9468 5778 9808 5864
rect 9468 5722 9538 5778
rect 9594 5722 9680 5778
rect 9736 5722 9808 5778
rect 9468 5636 9808 5722
rect 9468 5580 9538 5636
rect 9594 5580 9680 5636
rect 9736 5580 9808 5636
rect 9468 5494 9808 5580
rect 9468 5438 9538 5494
rect 9594 5438 9680 5494
rect 9736 5438 9808 5494
rect 9468 5352 9808 5438
rect 9468 5296 9538 5352
rect 9594 5296 9680 5352
rect 9736 5296 9808 5352
rect 9468 5210 9808 5296
rect 9468 5154 9538 5210
rect 9594 5154 9680 5210
rect 9736 5154 9808 5210
rect 9468 5068 9808 5154
rect 9468 5012 9538 5068
rect 9594 5012 9680 5068
rect 9736 5012 9808 5068
rect 9468 4926 9808 5012
rect 9468 4870 9538 4926
rect 9594 4870 9680 4926
rect 9736 4870 9808 4926
rect 9468 4784 9808 4870
rect 9468 4728 9538 4784
rect 9594 4728 9680 4784
rect 9736 4728 9808 4784
rect 9468 4642 9808 4728
rect 9468 4586 9538 4642
rect 9594 4586 9680 4642
rect 9736 4586 9808 4642
rect 9468 4500 9808 4586
rect 9468 4444 9538 4500
rect 9594 4444 9680 4500
rect 9736 4444 9808 4500
rect 9468 4358 9808 4444
rect 9468 4302 9538 4358
rect 9594 4302 9680 4358
rect 9736 4302 9808 4358
rect 9468 4216 9808 4302
rect 9468 4160 9538 4216
rect 9594 4160 9680 4216
rect 9736 4160 9808 4216
rect 9468 4074 9808 4160
rect 9468 4018 9538 4074
rect 9594 4018 9680 4074
rect 9736 4018 9808 4074
rect 9468 3932 9808 4018
rect 9468 3876 9538 3932
rect 9594 3876 9680 3932
rect 9736 3876 9808 3932
rect 9468 3790 9808 3876
rect 9468 3734 9538 3790
rect 9594 3734 9680 3790
rect 9736 3734 9808 3790
rect 9468 3648 9808 3734
rect 9468 3592 9538 3648
rect 9594 3592 9680 3648
rect 9736 3592 9808 3648
rect 9468 3506 9808 3592
rect 9468 3450 9538 3506
rect 9594 3450 9680 3506
rect 9736 3450 9808 3506
rect 9468 3364 9808 3450
rect 9468 3308 9538 3364
rect 9594 3308 9680 3364
rect 9736 3308 9808 3364
rect 9468 3222 9808 3308
rect 9468 3166 9538 3222
rect 9594 3166 9680 3222
rect 9736 3166 9808 3222
rect 9468 3080 9808 3166
rect 9468 3024 9538 3080
rect 9594 3024 9680 3080
rect 9736 3024 9808 3080
rect 9468 2938 9808 3024
rect 9468 2882 9538 2938
rect 9594 2882 9680 2938
rect 9736 2882 9808 2938
rect 9468 2796 9808 2882
rect 9468 2740 9538 2796
rect 9594 2740 9680 2796
rect 9736 2740 9808 2796
rect 9468 2654 9808 2740
rect 9468 2598 9538 2654
rect 9594 2598 9680 2654
rect 9736 2598 9808 2654
rect 9468 2512 9808 2598
rect 9468 2456 9538 2512
rect 9594 2456 9680 2512
rect 9736 2456 9808 2512
rect 9468 2370 9808 2456
rect 9468 2314 9538 2370
rect 9594 2314 9680 2370
rect 9736 2314 9808 2370
rect 9468 2228 9808 2314
rect 9468 2172 9538 2228
rect 9594 2172 9680 2228
rect 9736 2172 9808 2228
rect 9468 2086 9808 2172
rect 9468 2030 9538 2086
rect 9594 2030 9680 2086
rect 9736 2030 9808 2086
rect 9468 1944 9808 2030
rect 9468 1888 9538 1944
rect 9594 1888 9680 1944
rect 9736 1888 9808 1944
rect 9468 1802 9808 1888
rect 9468 1746 9538 1802
rect 9594 1746 9680 1802
rect 9736 1746 9808 1802
rect 9468 1660 9808 1746
rect 9468 1604 9538 1660
rect 9594 1604 9680 1660
rect 9736 1604 9808 1660
rect 9468 1518 9808 1604
rect 9468 1462 9538 1518
rect 9594 1462 9680 1518
rect 9736 1462 9808 1518
rect 9468 1376 9808 1462
rect 9468 1320 9538 1376
rect 9594 1320 9680 1376
rect 9736 1320 9808 1376
rect 9468 1234 9808 1320
rect 9468 1178 9538 1234
rect 9594 1178 9680 1234
rect 9736 1178 9808 1234
rect 9468 1092 9808 1178
rect 9468 1036 9538 1092
rect 9594 1036 9680 1092
rect 9736 1036 9808 1092
rect 9468 950 9808 1036
rect 9468 894 9538 950
rect 9594 894 9680 950
rect 9736 894 9808 950
rect 9468 808 9808 894
rect 9468 752 9538 808
rect 9594 752 9680 808
rect 9736 752 9808 808
rect 9468 666 9808 752
rect 9468 610 9538 666
rect 9594 610 9680 666
rect 9736 610 9808 666
rect 9468 524 9808 610
rect 9468 468 9538 524
rect 9594 468 9680 524
rect 9736 468 9808 524
rect 9468 400 9808 468
rect 9868 12310 10208 12400
rect 9868 12254 9934 12310
rect 9990 12254 10076 12310
rect 10132 12254 10208 12310
rect 9868 12168 10208 12254
rect 9868 12112 9934 12168
rect 9990 12112 10076 12168
rect 10132 12112 10208 12168
rect 9868 12026 10208 12112
rect 9868 11970 9934 12026
rect 9990 11970 10076 12026
rect 10132 11970 10208 12026
rect 9868 11884 10208 11970
rect 9868 11828 9934 11884
rect 9990 11828 10076 11884
rect 10132 11828 10208 11884
rect 9868 11742 10208 11828
rect 9868 11686 9934 11742
rect 9990 11686 10076 11742
rect 10132 11686 10208 11742
rect 9868 11600 10208 11686
rect 9868 11544 9934 11600
rect 9990 11544 10076 11600
rect 10132 11544 10208 11600
rect 9868 11458 10208 11544
rect 9868 11402 9934 11458
rect 9990 11402 10076 11458
rect 10132 11402 10208 11458
rect 9868 11316 10208 11402
rect 9868 11260 9934 11316
rect 9990 11260 10076 11316
rect 10132 11260 10208 11316
rect 9868 11174 10208 11260
rect 9868 11118 9934 11174
rect 9990 11118 10076 11174
rect 10132 11118 10208 11174
rect 9868 11032 10208 11118
rect 9868 10976 9934 11032
rect 9990 10976 10076 11032
rect 10132 10976 10208 11032
rect 9868 10890 10208 10976
rect 9868 10834 9934 10890
rect 9990 10834 10076 10890
rect 10132 10834 10208 10890
rect 9868 10748 10208 10834
rect 9868 10692 9934 10748
rect 9990 10692 10076 10748
rect 10132 10692 10208 10748
rect 9868 10606 10208 10692
rect 9868 10550 9934 10606
rect 9990 10550 10076 10606
rect 10132 10550 10208 10606
rect 9868 10464 10208 10550
rect 9868 10408 9934 10464
rect 9990 10408 10076 10464
rect 10132 10408 10208 10464
rect 9868 10322 10208 10408
rect 9868 10266 9934 10322
rect 9990 10266 10076 10322
rect 10132 10266 10208 10322
rect 9868 10180 10208 10266
rect 9868 10124 9934 10180
rect 9990 10124 10076 10180
rect 10132 10124 10208 10180
rect 9868 10038 10208 10124
rect 9868 9982 9934 10038
rect 9990 9982 10076 10038
rect 10132 9982 10208 10038
rect 9868 9896 10208 9982
rect 9868 9840 9934 9896
rect 9990 9840 10076 9896
rect 10132 9840 10208 9896
rect 9868 9754 10208 9840
rect 9868 9698 9934 9754
rect 9990 9698 10076 9754
rect 10132 9698 10208 9754
rect 9868 9612 10208 9698
rect 9868 9556 9934 9612
rect 9990 9556 10076 9612
rect 10132 9556 10208 9612
rect 9868 9470 10208 9556
rect 9868 9414 9934 9470
rect 9990 9414 10076 9470
rect 10132 9414 10208 9470
rect 9868 9328 10208 9414
rect 9868 9272 9934 9328
rect 9990 9272 10076 9328
rect 10132 9272 10208 9328
rect 9868 9186 10208 9272
rect 9868 9130 9934 9186
rect 9990 9130 10076 9186
rect 10132 9130 10208 9186
rect 9868 9044 10208 9130
rect 9868 8988 9934 9044
rect 9990 8988 10076 9044
rect 10132 8988 10208 9044
rect 9868 8902 10208 8988
rect 9868 8846 9934 8902
rect 9990 8846 10076 8902
rect 10132 8846 10208 8902
rect 9868 8760 10208 8846
rect 9868 8704 9934 8760
rect 9990 8704 10076 8760
rect 10132 8704 10208 8760
rect 9868 8618 10208 8704
rect 9868 8562 9934 8618
rect 9990 8562 10076 8618
rect 10132 8562 10208 8618
rect 9868 8476 10208 8562
rect 9868 8420 9934 8476
rect 9990 8420 10076 8476
rect 10132 8420 10208 8476
rect 9868 8334 10208 8420
rect 9868 8278 9934 8334
rect 9990 8278 10076 8334
rect 10132 8278 10208 8334
rect 9868 8192 10208 8278
rect 9868 8136 9934 8192
rect 9990 8136 10076 8192
rect 10132 8136 10208 8192
rect 9868 8050 10208 8136
rect 9868 7994 9934 8050
rect 9990 7994 10076 8050
rect 10132 7994 10208 8050
rect 9868 7908 10208 7994
rect 9868 7852 9934 7908
rect 9990 7852 10076 7908
rect 10132 7852 10208 7908
rect 9868 7766 10208 7852
rect 9868 7710 9934 7766
rect 9990 7710 10076 7766
rect 10132 7710 10208 7766
rect 9868 7624 10208 7710
rect 9868 7568 9934 7624
rect 9990 7568 10076 7624
rect 10132 7568 10208 7624
rect 9868 7482 10208 7568
rect 9868 7426 9934 7482
rect 9990 7426 10076 7482
rect 10132 7426 10208 7482
rect 9868 7340 10208 7426
rect 9868 7284 9934 7340
rect 9990 7284 10076 7340
rect 10132 7284 10208 7340
rect 9868 7198 10208 7284
rect 9868 7142 9934 7198
rect 9990 7142 10076 7198
rect 10132 7142 10208 7198
rect 9868 7056 10208 7142
rect 9868 7000 9934 7056
rect 9990 7000 10076 7056
rect 10132 7000 10208 7056
rect 9868 6914 10208 7000
rect 9868 6858 9934 6914
rect 9990 6858 10076 6914
rect 10132 6858 10208 6914
rect 9868 6772 10208 6858
rect 9868 6716 9934 6772
rect 9990 6716 10076 6772
rect 10132 6716 10208 6772
rect 9868 6630 10208 6716
rect 9868 6574 9934 6630
rect 9990 6574 10076 6630
rect 10132 6574 10208 6630
rect 9868 6488 10208 6574
rect 9868 6432 9934 6488
rect 9990 6432 10076 6488
rect 10132 6432 10208 6488
rect 9868 6346 10208 6432
rect 9868 6290 9934 6346
rect 9990 6290 10076 6346
rect 10132 6290 10208 6346
rect 9868 6204 10208 6290
rect 9868 6148 9934 6204
rect 9990 6148 10076 6204
rect 10132 6148 10208 6204
rect 9868 6062 10208 6148
rect 9868 6006 9934 6062
rect 9990 6006 10076 6062
rect 10132 6006 10208 6062
rect 9868 5920 10208 6006
rect 9868 5864 9934 5920
rect 9990 5864 10076 5920
rect 10132 5864 10208 5920
rect 9868 5778 10208 5864
rect 9868 5722 9934 5778
rect 9990 5722 10076 5778
rect 10132 5722 10208 5778
rect 9868 5636 10208 5722
rect 9868 5580 9934 5636
rect 9990 5580 10076 5636
rect 10132 5580 10208 5636
rect 9868 5494 10208 5580
rect 9868 5438 9934 5494
rect 9990 5438 10076 5494
rect 10132 5438 10208 5494
rect 9868 5352 10208 5438
rect 9868 5296 9934 5352
rect 9990 5296 10076 5352
rect 10132 5296 10208 5352
rect 9868 5210 10208 5296
rect 9868 5154 9934 5210
rect 9990 5154 10076 5210
rect 10132 5154 10208 5210
rect 9868 5068 10208 5154
rect 9868 5012 9934 5068
rect 9990 5012 10076 5068
rect 10132 5012 10208 5068
rect 9868 4926 10208 5012
rect 9868 4870 9934 4926
rect 9990 4870 10076 4926
rect 10132 4870 10208 4926
rect 9868 4784 10208 4870
rect 9868 4728 9934 4784
rect 9990 4728 10076 4784
rect 10132 4728 10208 4784
rect 9868 4642 10208 4728
rect 9868 4586 9934 4642
rect 9990 4586 10076 4642
rect 10132 4586 10208 4642
rect 9868 4500 10208 4586
rect 9868 4444 9934 4500
rect 9990 4444 10076 4500
rect 10132 4444 10208 4500
rect 9868 4358 10208 4444
rect 9868 4302 9934 4358
rect 9990 4302 10076 4358
rect 10132 4302 10208 4358
rect 9868 4216 10208 4302
rect 9868 4160 9934 4216
rect 9990 4160 10076 4216
rect 10132 4160 10208 4216
rect 9868 4074 10208 4160
rect 9868 4018 9934 4074
rect 9990 4018 10076 4074
rect 10132 4018 10208 4074
rect 9868 3932 10208 4018
rect 9868 3876 9934 3932
rect 9990 3876 10076 3932
rect 10132 3876 10208 3932
rect 9868 3790 10208 3876
rect 9868 3734 9934 3790
rect 9990 3734 10076 3790
rect 10132 3734 10208 3790
rect 9868 3648 10208 3734
rect 9868 3592 9934 3648
rect 9990 3592 10076 3648
rect 10132 3592 10208 3648
rect 9868 3506 10208 3592
rect 9868 3450 9934 3506
rect 9990 3450 10076 3506
rect 10132 3450 10208 3506
rect 9868 3364 10208 3450
rect 9868 3308 9934 3364
rect 9990 3308 10076 3364
rect 10132 3308 10208 3364
rect 9868 3222 10208 3308
rect 9868 3166 9934 3222
rect 9990 3166 10076 3222
rect 10132 3166 10208 3222
rect 9868 3080 10208 3166
rect 9868 3024 9934 3080
rect 9990 3024 10076 3080
rect 10132 3024 10208 3080
rect 9868 2938 10208 3024
rect 9868 2882 9934 2938
rect 9990 2882 10076 2938
rect 10132 2882 10208 2938
rect 9868 2796 10208 2882
rect 9868 2740 9934 2796
rect 9990 2740 10076 2796
rect 10132 2740 10208 2796
rect 9868 2654 10208 2740
rect 9868 2598 9934 2654
rect 9990 2598 10076 2654
rect 10132 2598 10208 2654
rect 9868 2512 10208 2598
rect 9868 2456 9934 2512
rect 9990 2456 10076 2512
rect 10132 2456 10208 2512
rect 9868 2370 10208 2456
rect 9868 2314 9934 2370
rect 9990 2314 10076 2370
rect 10132 2314 10208 2370
rect 9868 2228 10208 2314
rect 9868 2172 9934 2228
rect 9990 2172 10076 2228
rect 10132 2172 10208 2228
rect 9868 2086 10208 2172
rect 9868 2030 9934 2086
rect 9990 2030 10076 2086
rect 10132 2030 10208 2086
rect 9868 1944 10208 2030
rect 9868 1888 9934 1944
rect 9990 1888 10076 1944
rect 10132 1888 10208 1944
rect 9868 1802 10208 1888
rect 9868 1746 9934 1802
rect 9990 1746 10076 1802
rect 10132 1746 10208 1802
rect 9868 1660 10208 1746
rect 9868 1604 9934 1660
rect 9990 1604 10076 1660
rect 10132 1604 10208 1660
rect 9868 1518 10208 1604
rect 9868 1462 9934 1518
rect 9990 1462 10076 1518
rect 10132 1462 10208 1518
rect 9868 1376 10208 1462
rect 9868 1320 9934 1376
rect 9990 1320 10076 1376
rect 10132 1320 10208 1376
rect 9868 1234 10208 1320
rect 9868 1178 9934 1234
rect 9990 1178 10076 1234
rect 10132 1178 10208 1234
rect 9868 1092 10208 1178
rect 9868 1036 9934 1092
rect 9990 1036 10076 1092
rect 10132 1036 10208 1092
rect 9868 950 10208 1036
rect 9868 894 9934 950
rect 9990 894 10076 950
rect 10132 894 10208 950
rect 9868 808 10208 894
rect 9868 752 9934 808
rect 9990 752 10076 808
rect 10132 752 10208 808
rect 9868 666 10208 752
rect 9868 610 9934 666
rect 9990 610 10076 666
rect 10132 610 10208 666
rect 9868 524 10208 610
rect 9868 468 9934 524
rect 9990 468 10076 524
rect 10132 468 10208 524
rect 9868 400 10208 468
rect 10268 12310 10608 12400
rect 10268 12254 10334 12310
rect 10390 12254 10476 12310
rect 10532 12254 10608 12310
rect 10268 12168 10608 12254
rect 10268 12112 10334 12168
rect 10390 12112 10476 12168
rect 10532 12112 10608 12168
rect 10268 12026 10608 12112
rect 10268 11970 10334 12026
rect 10390 11970 10476 12026
rect 10532 11970 10608 12026
rect 10268 11884 10608 11970
rect 10268 11828 10334 11884
rect 10390 11828 10476 11884
rect 10532 11828 10608 11884
rect 10268 11742 10608 11828
rect 10268 11686 10334 11742
rect 10390 11686 10476 11742
rect 10532 11686 10608 11742
rect 10268 11600 10608 11686
rect 10268 11544 10334 11600
rect 10390 11544 10476 11600
rect 10532 11544 10608 11600
rect 10268 11458 10608 11544
rect 10268 11402 10334 11458
rect 10390 11402 10476 11458
rect 10532 11402 10608 11458
rect 10268 11316 10608 11402
rect 10268 11260 10334 11316
rect 10390 11260 10476 11316
rect 10532 11260 10608 11316
rect 10268 11174 10608 11260
rect 10268 11118 10334 11174
rect 10390 11118 10476 11174
rect 10532 11118 10608 11174
rect 10268 11032 10608 11118
rect 10268 10976 10334 11032
rect 10390 10976 10476 11032
rect 10532 10976 10608 11032
rect 10268 10890 10608 10976
rect 10268 10834 10334 10890
rect 10390 10834 10476 10890
rect 10532 10834 10608 10890
rect 10268 10748 10608 10834
rect 10268 10692 10334 10748
rect 10390 10692 10476 10748
rect 10532 10692 10608 10748
rect 10268 10606 10608 10692
rect 10268 10550 10334 10606
rect 10390 10550 10476 10606
rect 10532 10550 10608 10606
rect 10268 10464 10608 10550
rect 10268 10408 10334 10464
rect 10390 10408 10476 10464
rect 10532 10408 10608 10464
rect 10268 10322 10608 10408
rect 10268 10266 10334 10322
rect 10390 10266 10476 10322
rect 10532 10266 10608 10322
rect 10268 10180 10608 10266
rect 10268 10124 10334 10180
rect 10390 10124 10476 10180
rect 10532 10124 10608 10180
rect 10268 10038 10608 10124
rect 10268 9982 10334 10038
rect 10390 9982 10476 10038
rect 10532 9982 10608 10038
rect 10268 9896 10608 9982
rect 10268 9840 10334 9896
rect 10390 9840 10476 9896
rect 10532 9840 10608 9896
rect 10268 9754 10608 9840
rect 10268 9698 10334 9754
rect 10390 9698 10476 9754
rect 10532 9698 10608 9754
rect 10268 9612 10608 9698
rect 10268 9556 10334 9612
rect 10390 9556 10476 9612
rect 10532 9556 10608 9612
rect 10268 9470 10608 9556
rect 10268 9414 10334 9470
rect 10390 9414 10476 9470
rect 10532 9414 10608 9470
rect 10268 9328 10608 9414
rect 10268 9272 10334 9328
rect 10390 9272 10476 9328
rect 10532 9272 10608 9328
rect 10268 9186 10608 9272
rect 10268 9130 10334 9186
rect 10390 9130 10476 9186
rect 10532 9130 10608 9186
rect 10268 9044 10608 9130
rect 10268 8988 10334 9044
rect 10390 8988 10476 9044
rect 10532 8988 10608 9044
rect 10268 8902 10608 8988
rect 10268 8846 10334 8902
rect 10390 8846 10476 8902
rect 10532 8846 10608 8902
rect 10268 8760 10608 8846
rect 10268 8704 10334 8760
rect 10390 8704 10476 8760
rect 10532 8704 10608 8760
rect 10268 8618 10608 8704
rect 10268 8562 10334 8618
rect 10390 8562 10476 8618
rect 10532 8562 10608 8618
rect 10268 8476 10608 8562
rect 10268 8420 10334 8476
rect 10390 8420 10476 8476
rect 10532 8420 10608 8476
rect 10268 8334 10608 8420
rect 10268 8278 10334 8334
rect 10390 8278 10476 8334
rect 10532 8278 10608 8334
rect 10268 8192 10608 8278
rect 10268 8136 10334 8192
rect 10390 8136 10476 8192
rect 10532 8136 10608 8192
rect 10268 8050 10608 8136
rect 10268 7994 10334 8050
rect 10390 7994 10476 8050
rect 10532 7994 10608 8050
rect 10268 7908 10608 7994
rect 10268 7852 10334 7908
rect 10390 7852 10476 7908
rect 10532 7852 10608 7908
rect 10268 7766 10608 7852
rect 10268 7710 10334 7766
rect 10390 7710 10476 7766
rect 10532 7710 10608 7766
rect 10268 7624 10608 7710
rect 10268 7568 10334 7624
rect 10390 7568 10476 7624
rect 10532 7568 10608 7624
rect 10268 7482 10608 7568
rect 10268 7426 10334 7482
rect 10390 7426 10476 7482
rect 10532 7426 10608 7482
rect 10268 7340 10608 7426
rect 10268 7284 10334 7340
rect 10390 7284 10476 7340
rect 10532 7284 10608 7340
rect 10268 7198 10608 7284
rect 10268 7142 10334 7198
rect 10390 7142 10476 7198
rect 10532 7142 10608 7198
rect 10268 7056 10608 7142
rect 10268 7000 10334 7056
rect 10390 7000 10476 7056
rect 10532 7000 10608 7056
rect 10268 6914 10608 7000
rect 10268 6858 10334 6914
rect 10390 6858 10476 6914
rect 10532 6858 10608 6914
rect 10268 6772 10608 6858
rect 10268 6716 10334 6772
rect 10390 6716 10476 6772
rect 10532 6716 10608 6772
rect 10268 6630 10608 6716
rect 10268 6574 10334 6630
rect 10390 6574 10476 6630
rect 10532 6574 10608 6630
rect 10268 6488 10608 6574
rect 10268 6432 10334 6488
rect 10390 6432 10476 6488
rect 10532 6432 10608 6488
rect 10268 6346 10608 6432
rect 10268 6290 10334 6346
rect 10390 6290 10476 6346
rect 10532 6290 10608 6346
rect 10268 6204 10608 6290
rect 10268 6148 10334 6204
rect 10390 6148 10476 6204
rect 10532 6148 10608 6204
rect 10268 6062 10608 6148
rect 10268 6006 10334 6062
rect 10390 6006 10476 6062
rect 10532 6006 10608 6062
rect 10268 5920 10608 6006
rect 10268 5864 10334 5920
rect 10390 5864 10476 5920
rect 10532 5864 10608 5920
rect 10268 5778 10608 5864
rect 10268 5722 10334 5778
rect 10390 5722 10476 5778
rect 10532 5722 10608 5778
rect 10268 5636 10608 5722
rect 10268 5580 10334 5636
rect 10390 5580 10476 5636
rect 10532 5580 10608 5636
rect 10268 5494 10608 5580
rect 10268 5438 10334 5494
rect 10390 5438 10476 5494
rect 10532 5438 10608 5494
rect 10268 5352 10608 5438
rect 10268 5296 10334 5352
rect 10390 5296 10476 5352
rect 10532 5296 10608 5352
rect 10268 5210 10608 5296
rect 10268 5154 10334 5210
rect 10390 5154 10476 5210
rect 10532 5154 10608 5210
rect 10268 5068 10608 5154
rect 10268 5012 10334 5068
rect 10390 5012 10476 5068
rect 10532 5012 10608 5068
rect 10268 4926 10608 5012
rect 10268 4870 10334 4926
rect 10390 4870 10476 4926
rect 10532 4870 10608 4926
rect 10268 4784 10608 4870
rect 10268 4728 10334 4784
rect 10390 4728 10476 4784
rect 10532 4728 10608 4784
rect 10268 4642 10608 4728
rect 10268 4586 10334 4642
rect 10390 4586 10476 4642
rect 10532 4586 10608 4642
rect 10268 4500 10608 4586
rect 10268 4444 10334 4500
rect 10390 4444 10476 4500
rect 10532 4444 10608 4500
rect 10268 4358 10608 4444
rect 10268 4302 10334 4358
rect 10390 4302 10476 4358
rect 10532 4302 10608 4358
rect 10268 4216 10608 4302
rect 10268 4160 10334 4216
rect 10390 4160 10476 4216
rect 10532 4160 10608 4216
rect 10268 4074 10608 4160
rect 10268 4018 10334 4074
rect 10390 4018 10476 4074
rect 10532 4018 10608 4074
rect 10268 3932 10608 4018
rect 10268 3876 10334 3932
rect 10390 3876 10476 3932
rect 10532 3876 10608 3932
rect 10268 3790 10608 3876
rect 10268 3734 10334 3790
rect 10390 3734 10476 3790
rect 10532 3734 10608 3790
rect 10268 3648 10608 3734
rect 10268 3592 10334 3648
rect 10390 3592 10476 3648
rect 10532 3592 10608 3648
rect 10268 3506 10608 3592
rect 10268 3450 10334 3506
rect 10390 3450 10476 3506
rect 10532 3450 10608 3506
rect 10268 3364 10608 3450
rect 10268 3308 10334 3364
rect 10390 3308 10476 3364
rect 10532 3308 10608 3364
rect 10268 3222 10608 3308
rect 10268 3166 10334 3222
rect 10390 3166 10476 3222
rect 10532 3166 10608 3222
rect 10268 3080 10608 3166
rect 10268 3024 10334 3080
rect 10390 3024 10476 3080
rect 10532 3024 10608 3080
rect 10268 2938 10608 3024
rect 10268 2882 10334 2938
rect 10390 2882 10476 2938
rect 10532 2882 10608 2938
rect 10268 2796 10608 2882
rect 10268 2740 10334 2796
rect 10390 2740 10476 2796
rect 10532 2740 10608 2796
rect 10268 2654 10608 2740
rect 10268 2598 10334 2654
rect 10390 2598 10476 2654
rect 10532 2598 10608 2654
rect 10268 2512 10608 2598
rect 10268 2456 10334 2512
rect 10390 2456 10476 2512
rect 10532 2456 10608 2512
rect 10268 2370 10608 2456
rect 10268 2314 10334 2370
rect 10390 2314 10476 2370
rect 10532 2314 10608 2370
rect 10268 2228 10608 2314
rect 10268 2172 10334 2228
rect 10390 2172 10476 2228
rect 10532 2172 10608 2228
rect 10268 2086 10608 2172
rect 10268 2030 10334 2086
rect 10390 2030 10476 2086
rect 10532 2030 10608 2086
rect 10268 1944 10608 2030
rect 10268 1888 10334 1944
rect 10390 1888 10476 1944
rect 10532 1888 10608 1944
rect 10268 1802 10608 1888
rect 10268 1746 10334 1802
rect 10390 1746 10476 1802
rect 10532 1746 10608 1802
rect 10268 1660 10608 1746
rect 10268 1604 10334 1660
rect 10390 1604 10476 1660
rect 10532 1604 10608 1660
rect 10268 1518 10608 1604
rect 10268 1462 10334 1518
rect 10390 1462 10476 1518
rect 10532 1462 10608 1518
rect 10268 1376 10608 1462
rect 10268 1320 10334 1376
rect 10390 1320 10476 1376
rect 10532 1320 10608 1376
rect 10268 1234 10608 1320
rect 10268 1178 10334 1234
rect 10390 1178 10476 1234
rect 10532 1178 10608 1234
rect 10268 1092 10608 1178
rect 10268 1036 10334 1092
rect 10390 1036 10476 1092
rect 10532 1036 10608 1092
rect 10268 950 10608 1036
rect 10268 894 10334 950
rect 10390 894 10476 950
rect 10532 894 10608 950
rect 10268 808 10608 894
rect 10268 752 10334 808
rect 10390 752 10476 808
rect 10532 752 10608 808
rect 10268 666 10608 752
rect 10268 610 10334 666
rect 10390 610 10476 666
rect 10532 610 10608 666
rect 10268 524 10608 610
rect 10268 468 10334 524
rect 10390 468 10476 524
rect 10532 468 10608 524
rect 10268 400 10608 468
rect 10668 12310 11008 12400
rect 10668 12254 10731 12310
rect 10787 12254 10873 12310
rect 10929 12254 11008 12310
rect 10668 12168 11008 12254
rect 10668 12112 10731 12168
rect 10787 12112 10873 12168
rect 10929 12112 11008 12168
rect 10668 12026 11008 12112
rect 10668 11970 10731 12026
rect 10787 11970 10873 12026
rect 10929 11970 11008 12026
rect 10668 11884 11008 11970
rect 10668 11828 10731 11884
rect 10787 11828 10873 11884
rect 10929 11828 11008 11884
rect 10668 11742 11008 11828
rect 10668 11686 10731 11742
rect 10787 11686 10873 11742
rect 10929 11686 11008 11742
rect 10668 11600 11008 11686
rect 10668 11544 10731 11600
rect 10787 11544 10873 11600
rect 10929 11544 11008 11600
rect 10668 11458 11008 11544
rect 10668 11402 10731 11458
rect 10787 11402 10873 11458
rect 10929 11402 11008 11458
rect 10668 11316 11008 11402
rect 10668 11260 10731 11316
rect 10787 11260 10873 11316
rect 10929 11260 11008 11316
rect 10668 11174 11008 11260
rect 10668 11118 10731 11174
rect 10787 11118 10873 11174
rect 10929 11118 11008 11174
rect 10668 11032 11008 11118
rect 10668 10976 10731 11032
rect 10787 10976 10873 11032
rect 10929 10976 11008 11032
rect 10668 10890 11008 10976
rect 10668 10834 10731 10890
rect 10787 10834 10873 10890
rect 10929 10834 11008 10890
rect 10668 10748 11008 10834
rect 10668 10692 10731 10748
rect 10787 10692 10873 10748
rect 10929 10692 11008 10748
rect 10668 10606 11008 10692
rect 10668 10550 10731 10606
rect 10787 10550 10873 10606
rect 10929 10550 11008 10606
rect 10668 10464 11008 10550
rect 10668 10408 10731 10464
rect 10787 10408 10873 10464
rect 10929 10408 11008 10464
rect 10668 10322 11008 10408
rect 10668 10266 10731 10322
rect 10787 10266 10873 10322
rect 10929 10266 11008 10322
rect 10668 10180 11008 10266
rect 10668 10124 10731 10180
rect 10787 10124 10873 10180
rect 10929 10124 11008 10180
rect 10668 10038 11008 10124
rect 10668 9982 10731 10038
rect 10787 9982 10873 10038
rect 10929 9982 11008 10038
rect 10668 9896 11008 9982
rect 10668 9840 10731 9896
rect 10787 9840 10873 9896
rect 10929 9840 11008 9896
rect 10668 9754 11008 9840
rect 10668 9698 10731 9754
rect 10787 9698 10873 9754
rect 10929 9698 11008 9754
rect 10668 9612 11008 9698
rect 10668 9556 10731 9612
rect 10787 9556 10873 9612
rect 10929 9556 11008 9612
rect 10668 9470 11008 9556
rect 10668 9414 10731 9470
rect 10787 9414 10873 9470
rect 10929 9414 11008 9470
rect 10668 9328 11008 9414
rect 10668 9272 10731 9328
rect 10787 9272 10873 9328
rect 10929 9272 11008 9328
rect 10668 9186 11008 9272
rect 10668 9130 10731 9186
rect 10787 9130 10873 9186
rect 10929 9130 11008 9186
rect 10668 9044 11008 9130
rect 10668 8988 10731 9044
rect 10787 8988 10873 9044
rect 10929 8988 11008 9044
rect 10668 8902 11008 8988
rect 10668 8846 10731 8902
rect 10787 8846 10873 8902
rect 10929 8846 11008 8902
rect 10668 8760 11008 8846
rect 10668 8704 10731 8760
rect 10787 8704 10873 8760
rect 10929 8704 11008 8760
rect 10668 8618 11008 8704
rect 10668 8562 10731 8618
rect 10787 8562 10873 8618
rect 10929 8562 11008 8618
rect 10668 8476 11008 8562
rect 10668 8420 10731 8476
rect 10787 8420 10873 8476
rect 10929 8420 11008 8476
rect 10668 8334 11008 8420
rect 10668 8278 10731 8334
rect 10787 8278 10873 8334
rect 10929 8278 11008 8334
rect 10668 8192 11008 8278
rect 10668 8136 10731 8192
rect 10787 8136 10873 8192
rect 10929 8136 11008 8192
rect 10668 8050 11008 8136
rect 10668 7994 10731 8050
rect 10787 7994 10873 8050
rect 10929 7994 11008 8050
rect 10668 7908 11008 7994
rect 10668 7852 10731 7908
rect 10787 7852 10873 7908
rect 10929 7852 11008 7908
rect 10668 7766 11008 7852
rect 10668 7710 10731 7766
rect 10787 7710 10873 7766
rect 10929 7710 11008 7766
rect 10668 7624 11008 7710
rect 10668 7568 10731 7624
rect 10787 7568 10873 7624
rect 10929 7568 11008 7624
rect 10668 7482 11008 7568
rect 10668 7426 10731 7482
rect 10787 7426 10873 7482
rect 10929 7426 11008 7482
rect 10668 7340 11008 7426
rect 10668 7284 10731 7340
rect 10787 7284 10873 7340
rect 10929 7284 11008 7340
rect 10668 7198 11008 7284
rect 10668 7142 10731 7198
rect 10787 7142 10873 7198
rect 10929 7142 11008 7198
rect 10668 7056 11008 7142
rect 10668 7000 10731 7056
rect 10787 7000 10873 7056
rect 10929 7000 11008 7056
rect 10668 6914 11008 7000
rect 10668 6858 10731 6914
rect 10787 6858 10873 6914
rect 10929 6858 11008 6914
rect 10668 6772 11008 6858
rect 10668 6716 10731 6772
rect 10787 6716 10873 6772
rect 10929 6716 11008 6772
rect 10668 6630 11008 6716
rect 10668 6574 10731 6630
rect 10787 6574 10873 6630
rect 10929 6574 11008 6630
rect 10668 6488 11008 6574
rect 10668 6432 10731 6488
rect 10787 6432 10873 6488
rect 10929 6432 11008 6488
rect 10668 6346 11008 6432
rect 10668 6290 10731 6346
rect 10787 6290 10873 6346
rect 10929 6290 11008 6346
rect 10668 6204 11008 6290
rect 10668 6148 10731 6204
rect 10787 6148 10873 6204
rect 10929 6148 11008 6204
rect 10668 6062 11008 6148
rect 10668 6006 10731 6062
rect 10787 6006 10873 6062
rect 10929 6006 11008 6062
rect 10668 5920 11008 6006
rect 10668 5864 10731 5920
rect 10787 5864 10873 5920
rect 10929 5864 11008 5920
rect 10668 5778 11008 5864
rect 10668 5722 10731 5778
rect 10787 5722 10873 5778
rect 10929 5722 11008 5778
rect 10668 5636 11008 5722
rect 10668 5580 10731 5636
rect 10787 5580 10873 5636
rect 10929 5580 11008 5636
rect 10668 5494 11008 5580
rect 10668 5438 10731 5494
rect 10787 5438 10873 5494
rect 10929 5438 11008 5494
rect 10668 5352 11008 5438
rect 10668 5296 10731 5352
rect 10787 5296 10873 5352
rect 10929 5296 11008 5352
rect 10668 5210 11008 5296
rect 10668 5154 10731 5210
rect 10787 5154 10873 5210
rect 10929 5154 11008 5210
rect 10668 5068 11008 5154
rect 10668 5012 10731 5068
rect 10787 5012 10873 5068
rect 10929 5012 11008 5068
rect 10668 4926 11008 5012
rect 10668 4870 10731 4926
rect 10787 4870 10873 4926
rect 10929 4870 11008 4926
rect 10668 4784 11008 4870
rect 10668 4728 10731 4784
rect 10787 4728 10873 4784
rect 10929 4728 11008 4784
rect 10668 4642 11008 4728
rect 10668 4586 10731 4642
rect 10787 4586 10873 4642
rect 10929 4586 11008 4642
rect 10668 4500 11008 4586
rect 10668 4444 10731 4500
rect 10787 4444 10873 4500
rect 10929 4444 11008 4500
rect 10668 4358 11008 4444
rect 10668 4302 10731 4358
rect 10787 4302 10873 4358
rect 10929 4302 11008 4358
rect 10668 4216 11008 4302
rect 10668 4160 10731 4216
rect 10787 4160 10873 4216
rect 10929 4160 11008 4216
rect 10668 4074 11008 4160
rect 10668 4018 10731 4074
rect 10787 4018 10873 4074
rect 10929 4018 11008 4074
rect 10668 3932 11008 4018
rect 10668 3876 10731 3932
rect 10787 3876 10873 3932
rect 10929 3876 11008 3932
rect 10668 3790 11008 3876
rect 10668 3734 10731 3790
rect 10787 3734 10873 3790
rect 10929 3734 11008 3790
rect 10668 3648 11008 3734
rect 10668 3592 10731 3648
rect 10787 3592 10873 3648
rect 10929 3592 11008 3648
rect 10668 3506 11008 3592
rect 10668 3450 10731 3506
rect 10787 3450 10873 3506
rect 10929 3450 11008 3506
rect 10668 3364 11008 3450
rect 10668 3308 10731 3364
rect 10787 3308 10873 3364
rect 10929 3308 11008 3364
rect 10668 3222 11008 3308
rect 10668 3166 10731 3222
rect 10787 3166 10873 3222
rect 10929 3166 11008 3222
rect 10668 3080 11008 3166
rect 10668 3024 10731 3080
rect 10787 3024 10873 3080
rect 10929 3024 11008 3080
rect 10668 2938 11008 3024
rect 10668 2882 10731 2938
rect 10787 2882 10873 2938
rect 10929 2882 11008 2938
rect 10668 2796 11008 2882
rect 10668 2740 10731 2796
rect 10787 2740 10873 2796
rect 10929 2740 11008 2796
rect 10668 2654 11008 2740
rect 10668 2598 10731 2654
rect 10787 2598 10873 2654
rect 10929 2598 11008 2654
rect 10668 2512 11008 2598
rect 10668 2456 10731 2512
rect 10787 2456 10873 2512
rect 10929 2456 11008 2512
rect 10668 2370 11008 2456
rect 10668 2314 10731 2370
rect 10787 2314 10873 2370
rect 10929 2314 11008 2370
rect 10668 2228 11008 2314
rect 10668 2172 10731 2228
rect 10787 2172 10873 2228
rect 10929 2172 11008 2228
rect 10668 2086 11008 2172
rect 10668 2030 10731 2086
rect 10787 2030 10873 2086
rect 10929 2030 11008 2086
rect 10668 1944 11008 2030
rect 10668 1888 10731 1944
rect 10787 1888 10873 1944
rect 10929 1888 11008 1944
rect 10668 1802 11008 1888
rect 10668 1746 10731 1802
rect 10787 1746 10873 1802
rect 10929 1746 11008 1802
rect 10668 1660 11008 1746
rect 10668 1604 10731 1660
rect 10787 1604 10873 1660
rect 10929 1604 11008 1660
rect 10668 1518 11008 1604
rect 10668 1462 10731 1518
rect 10787 1462 10873 1518
rect 10929 1462 11008 1518
rect 10668 1376 11008 1462
rect 10668 1320 10731 1376
rect 10787 1320 10873 1376
rect 10929 1320 11008 1376
rect 10668 1234 11008 1320
rect 10668 1178 10731 1234
rect 10787 1178 10873 1234
rect 10929 1178 11008 1234
rect 10668 1092 11008 1178
rect 10668 1036 10731 1092
rect 10787 1036 10873 1092
rect 10929 1036 11008 1092
rect 10668 950 11008 1036
rect 10668 894 10731 950
rect 10787 894 10873 950
rect 10929 894 11008 950
rect 10668 808 11008 894
rect 10668 752 10731 808
rect 10787 752 10873 808
rect 10929 752 11008 808
rect 10668 666 11008 752
rect 10668 610 10731 666
rect 10787 610 10873 666
rect 10929 610 11008 666
rect 10668 524 11008 610
rect 10668 468 10731 524
rect 10787 468 10873 524
rect 10929 468 11008 524
rect 10668 400 11008 468
rect 11068 12310 11408 12400
rect 11068 12254 11136 12310
rect 11192 12254 11278 12310
rect 11334 12254 11408 12310
rect 11068 12168 11408 12254
rect 11068 12112 11136 12168
rect 11192 12112 11278 12168
rect 11334 12112 11408 12168
rect 11068 12026 11408 12112
rect 11068 11970 11136 12026
rect 11192 11970 11278 12026
rect 11334 11970 11408 12026
rect 11068 11884 11408 11970
rect 11068 11828 11136 11884
rect 11192 11828 11278 11884
rect 11334 11828 11408 11884
rect 11068 11742 11408 11828
rect 11068 11686 11136 11742
rect 11192 11686 11278 11742
rect 11334 11686 11408 11742
rect 11068 11600 11408 11686
rect 11068 11544 11136 11600
rect 11192 11544 11278 11600
rect 11334 11544 11408 11600
rect 11068 11458 11408 11544
rect 11068 11402 11136 11458
rect 11192 11402 11278 11458
rect 11334 11402 11408 11458
rect 11068 11316 11408 11402
rect 11068 11260 11136 11316
rect 11192 11260 11278 11316
rect 11334 11260 11408 11316
rect 11068 11174 11408 11260
rect 11068 11118 11136 11174
rect 11192 11118 11278 11174
rect 11334 11118 11408 11174
rect 11068 11032 11408 11118
rect 11068 10976 11136 11032
rect 11192 10976 11278 11032
rect 11334 10976 11408 11032
rect 11068 10890 11408 10976
rect 11068 10834 11136 10890
rect 11192 10834 11278 10890
rect 11334 10834 11408 10890
rect 11068 10748 11408 10834
rect 11068 10692 11136 10748
rect 11192 10692 11278 10748
rect 11334 10692 11408 10748
rect 11068 10606 11408 10692
rect 11068 10550 11136 10606
rect 11192 10550 11278 10606
rect 11334 10550 11408 10606
rect 11068 10464 11408 10550
rect 11068 10408 11136 10464
rect 11192 10408 11278 10464
rect 11334 10408 11408 10464
rect 11068 10322 11408 10408
rect 11068 10266 11136 10322
rect 11192 10266 11278 10322
rect 11334 10266 11408 10322
rect 11068 10180 11408 10266
rect 11068 10124 11136 10180
rect 11192 10124 11278 10180
rect 11334 10124 11408 10180
rect 11068 10038 11408 10124
rect 11068 9982 11136 10038
rect 11192 9982 11278 10038
rect 11334 9982 11408 10038
rect 11068 9896 11408 9982
rect 11068 9840 11136 9896
rect 11192 9840 11278 9896
rect 11334 9840 11408 9896
rect 11068 9754 11408 9840
rect 11068 9698 11136 9754
rect 11192 9698 11278 9754
rect 11334 9698 11408 9754
rect 11068 9612 11408 9698
rect 11068 9556 11136 9612
rect 11192 9556 11278 9612
rect 11334 9556 11408 9612
rect 11068 9470 11408 9556
rect 11068 9414 11136 9470
rect 11192 9414 11278 9470
rect 11334 9414 11408 9470
rect 11068 9328 11408 9414
rect 11068 9272 11136 9328
rect 11192 9272 11278 9328
rect 11334 9272 11408 9328
rect 11068 9186 11408 9272
rect 11068 9130 11136 9186
rect 11192 9130 11278 9186
rect 11334 9130 11408 9186
rect 11068 9044 11408 9130
rect 11068 8988 11136 9044
rect 11192 8988 11278 9044
rect 11334 8988 11408 9044
rect 11068 8902 11408 8988
rect 11068 8846 11136 8902
rect 11192 8846 11278 8902
rect 11334 8846 11408 8902
rect 11068 8760 11408 8846
rect 11068 8704 11136 8760
rect 11192 8704 11278 8760
rect 11334 8704 11408 8760
rect 11068 8618 11408 8704
rect 11068 8562 11136 8618
rect 11192 8562 11278 8618
rect 11334 8562 11408 8618
rect 11068 8476 11408 8562
rect 11068 8420 11136 8476
rect 11192 8420 11278 8476
rect 11334 8420 11408 8476
rect 11068 8334 11408 8420
rect 11068 8278 11136 8334
rect 11192 8278 11278 8334
rect 11334 8278 11408 8334
rect 11068 8192 11408 8278
rect 11068 8136 11136 8192
rect 11192 8136 11278 8192
rect 11334 8136 11408 8192
rect 11068 8050 11408 8136
rect 11068 7994 11136 8050
rect 11192 7994 11278 8050
rect 11334 7994 11408 8050
rect 11068 7908 11408 7994
rect 11068 7852 11136 7908
rect 11192 7852 11278 7908
rect 11334 7852 11408 7908
rect 11068 7766 11408 7852
rect 11068 7710 11136 7766
rect 11192 7710 11278 7766
rect 11334 7710 11408 7766
rect 11068 7624 11408 7710
rect 11068 7568 11136 7624
rect 11192 7568 11278 7624
rect 11334 7568 11408 7624
rect 11068 7482 11408 7568
rect 11068 7426 11136 7482
rect 11192 7426 11278 7482
rect 11334 7426 11408 7482
rect 11068 7340 11408 7426
rect 11068 7284 11136 7340
rect 11192 7284 11278 7340
rect 11334 7284 11408 7340
rect 11068 7198 11408 7284
rect 11068 7142 11136 7198
rect 11192 7142 11278 7198
rect 11334 7142 11408 7198
rect 11068 7056 11408 7142
rect 11068 7000 11136 7056
rect 11192 7000 11278 7056
rect 11334 7000 11408 7056
rect 11068 6914 11408 7000
rect 11068 6858 11136 6914
rect 11192 6858 11278 6914
rect 11334 6858 11408 6914
rect 11068 6772 11408 6858
rect 11068 6716 11136 6772
rect 11192 6716 11278 6772
rect 11334 6716 11408 6772
rect 11068 6630 11408 6716
rect 11068 6574 11136 6630
rect 11192 6574 11278 6630
rect 11334 6574 11408 6630
rect 11068 6488 11408 6574
rect 11068 6432 11136 6488
rect 11192 6432 11278 6488
rect 11334 6432 11408 6488
rect 11068 6346 11408 6432
rect 11068 6290 11136 6346
rect 11192 6290 11278 6346
rect 11334 6290 11408 6346
rect 11068 6204 11408 6290
rect 11068 6148 11136 6204
rect 11192 6148 11278 6204
rect 11334 6148 11408 6204
rect 11068 6062 11408 6148
rect 11068 6006 11136 6062
rect 11192 6006 11278 6062
rect 11334 6006 11408 6062
rect 11068 5920 11408 6006
rect 11068 5864 11136 5920
rect 11192 5864 11278 5920
rect 11334 5864 11408 5920
rect 11068 5778 11408 5864
rect 11068 5722 11136 5778
rect 11192 5722 11278 5778
rect 11334 5722 11408 5778
rect 11068 5636 11408 5722
rect 11068 5580 11136 5636
rect 11192 5580 11278 5636
rect 11334 5580 11408 5636
rect 11068 5494 11408 5580
rect 11068 5438 11136 5494
rect 11192 5438 11278 5494
rect 11334 5438 11408 5494
rect 11068 5352 11408 5438
rect 11068 5296 11136 5352
rect 11192 5296 11278 5352
rect 11334 5296 11408 5352
rect 11068 5210 11408 5296
rect 11068 5154 11136 5210
rect 11192 5154 11278 5210
rect 11334 5154 11408 5210
rect 11068 5068 11408 5154
rect 11068 5012 11136 5068
rect 11192 5012 11278 5068
rect 11334 5012 11408 5068
rect 11068 4926 11408 5012
rect 11068 4870 11136 4926
rect 11192 4870 11278 4926
rect 11334 4870 11408 4926
rect 11068 4784 11408 4870
rect 11068 4728 11136 4784
rect 11192 4728 11278 4784
rect 11334 4728 11408 4784
rect 11068 4642 11408 4728
rect 11068 4586 11136 4642
rect 11192 4586 11278 4642
rect 11334 4586 11408 4642
rect 11068 4500 11408 4586
rect 11068 4444 11136 4500
rect 11192 4444 11278 4500
rect 11334 4444 11408 4500
rect 11068 4358 11408 4444
rect 11068 4302 11136 4358
rect 11192 4302 11278 4358
rect 11334 4302 11408 4358
rect 11068 4216 11408 4302
rect 11068 4160 11136 4216
rect 11192 4160 11278 4216
rect 11334 4160 11408 4216
rect 11068 4074 11408 4160
rect 11068 4018 11136 4074
rect 11192 4018 11278 4074
rect 11334 4018 11408 4074
rect 11068 3932 11408 4018
rect 11068 3876 11136 3932
rect 11192 3876 11278 3932
rect 11334 3876 11408 3932
rect 11068 3790 11408 3876
rect 11068 3734 11136 3790
rect 11192 3734 11278 3790
rect 11334 3734 11408 3790
rect 11068 3648 11408 3734
rect 11068 3592 11136 3648
rect 11192 3592 11278 3648
rect 11334 3592 11408 3648
rect 11068 3506 11408 3592
rect 11068 3450 11136 3506
rect 11192 3450 11278 3506
rect 11334 3450 11408 3506
rect 11068 3364 11408 3450
rect 11068 3308 11136 3364
rect 11192 3308 11278 3364
rect 11334 3308 11408 3364
rect 11068 3222 11408 3308
rect 11068 3166 11136 3222
rect 11192 3166 11278 3222
rect 11334 3166 11408 3222
rect 11068 3080 11408 3166
rect 11068 3024 11136 3080
rect 11192 3024 11278 3080
rect 11334 3024 11408 3080
rect 11068 2938 11408 3024
rect 11068 2882 11136 2938
rect 11192 2882 11278 2938
rect 11334 2882 11408 2938
rect 11068 2796 11408 2882
rect 11068 2740 11136 2796
rect 11192 2740 11278 2796
rect 11334 2740 11408 2796
rect 11068 2654 11408 2740
rect 11068 2598 11136 2654
rect 11192 2598 11278 2654
rect 11334 2598 11408 2654
rect 11068 2512 11408 2598
rect 11068 2456 11136 2512
rect 11192 2456 11278 2512
rect 11334 2456 11408 2512
rect 11068 2370 11408 2456
rect 11068 2314 11136 2370
rect 11192 2314 11278 2370
rect 11334 2314 11408 2370
rect 11068 2228 11408 2314
rect 11068 2172 11136 2228
rect 11192 2172 11278 2228
rect 11334 2172 11408 2228
rect 11068 2086 11408 2172
rect 11068 2030 11136 2086
rect 11192 2030 11278 2086
rect 11334 2030 11408 2086
rect 11068 1944 11408 2030
rect 11068 1888 11136 1944
rect 11192 1888 11278 1944
rect 11334 1888 11408 1944
rect 11068 1802 11408 1888
rect 11068 1746 11136 1802
rect 11192 1746 11278 1802
rect 11334 1746 11408 1802
rect 11068 1660 11408 1746
rect 11068 1604 11136 1660
rect 11192 1604 11278 1660
rect 11334 1604 11408 1660
rect 11068 1518 11408 1604
rect 11068 1462 11136 1518
rect 11192 1462 11278 1518
rect 11334 1462 11408 1518
rect 11068 1376 11408 1462
rect 11068 1320 11136 1376
rect 11192 1320 11278 1376
rect 11334 1320 11408 1376
rect 11068 1234 11408 1320
rect 11068 1178 11136 1234
rect 11192 1178 11278 1234
rect 11334 1178 11408 1234
rect 11068 1092 11408 1178
rect 11068 1036 11136 1092
rect 11192 1036 11278 1092
rect 11334 1036 11408 1092
rect 11068 950 11408 1036
rect 11068 894 11136 950
rect 11192 894 11278 950
rect 11334 894 11408 950
rect 11068 808 11408 894
rect 11068 752 11136 808
rect 11192 752 11278 808
rect 11334 752 11408 808
rect 11068 666 11408 752
rect 11068 610 11136 666
rect 11192 610 11278 666
rect 11334 610 11408 666
rect 11068 524 11408 610
rect 11068 468 11136 524
rect 11192 468 11278 524
rect 11334 468 11408 524
rect 11068 400 11408 468
rect 11468 12310 11808 12400
rect 11468 12254 11536 12310
rect 11592 12254 11678 12310
rect 11734 12254 11808 12310
rect 11468 12168 11808 12254
rect 11468 12112 11536 12168
rect 11592 12112 11678 12168
rect 11734 12112 11808 12168
rect 11468 12026 11808 12112
rect 11468 11970 11536 12026
rect 11592 11970 11678 12026
rect 11734 11970 11808 12026
rect 11468 11884 11808 11970
rect 11468 11828 11536 11884
rect 11592 11828 11678 11884
rect 11734 11828 11808 11884
rect 11468 11742 11808 11828
rect 11468 11686 11536 11742
rect 11592 11686 11678 11742
rect 11734 11686 11808 11742
rect 11468 11600 11808 11686
rect 11468 11544 11536 11600
rect 11592 11544 11678 11600
rect 11734 11544 11808 11600
rect 11468 11458 11808 11544
rect 11468 11402 11536 11458
rect 11592 11402 11678 11458
rect 11734 11402 11808 11458
rect 11468 11316 11808 11402
rect 11468 11260 11536 11316
rect 11592 11260 11678 11316
rect 11734 11260 11808 11316
rect 11468 11174 11808 11260
rect 11468 11118 11536 11174
rect 11592 11118 11678 11174
rect 11734 11118 11808 11174
rect 11468 11032 11808 11118
rect 11468 10976 11536 11032
rect 11592 10976 11678 11032
rect 11734 10976 11808 11032
rect 11468 10890 11808 10976
rect 11468 10834 11536 10890
rect 11592 10834 11678 10890
rect 11734 10834 11808 10890
rect 11468 10748 11808 10834
rect 11468 10692 11536 10748
rect 11592 10692 11678 10748
rect 11734 10692 11808 10748
rect 11468 10606 11808 10692
rect 11468 10550 11536 10606
rect 11592 10550 11678 10606
rect 11734 10550 11808 10606
rect 11468 10464 11808 10550
rect 11468 10408 11536 10464
rect 11592 10408 11678 10464
rect 11734 10408 11808 10464
rect 11468 10322 11808 10408
rect 11468 10266 11536 10322
rect 11592 10266 11678 10322
rect 11734 10266 11808 10322
rect 11468 10180 11808 10266
rect 11468 10124 11536 10180
rect 11592 10124 11678 10180
rect 11734 10124 11808 10180
rect 11468 10038 11808 10124
rect 11468 9982 11536 10038
rect 11592 9982 11678 10038
rect 11734 9982 11808 10038
rect 11468 9896 11808 9982
rect 11468 9840 11536 9896
rect 11592 9840 11678 9896
rect 11734 9840 11808 9896
rect 11468 9754 11808 9840
rect 11468 9698 11536 9754
rect 11592 9698 11678 9754
rect 11734 9698 11808 9754
rect 11468 9612 11808 9698
rect 11468 9556 11536 9612
rect 11592 9556 11678 9612
rect 11734 9556 11808 9612
rect 11468 9470 11808 9556
rect 11468 9414 11536 9470
rect 11592 9414 11678 9470
rect 11734 9414 11808 9470
rect 11468 9328 11808 9414
rect 11468 9272 11536 9328
rect 11592 9272 11678 9328
rect 11734 9272 11808 9328
rect 11468 9186 11808 9272
rect 11468 9130 11536 9186
rect 11592 9130 11678 9186
rect 11734 9130 11808 9186
rect 11468 9044 11808 9130
rect 11468 8988 11536 9044
rect 11592 8988 11678 9044
rect 11734 8988 11808 9044
rect 11468 8902 11808 8988
rect 11468 8846 11536 8902
rect 11592 8846 11678 8902
rect 11734 8846 11808 8902
rect 11468 8760 11808 8846
rect 11468 8704 11536 8760
rect 11592 8704 11678 8760
rect 11734 8704 11808 8760
rect 11468 8618 11808 8704
rect 11468 8562 11536 8618
rect 11592 8562 11678 8618
rect 11734 8562 11808 8618
rect 11468 8476 11808 8562
rect 11468 8420 11536 8476
rect 11592 8420 11678 8476
rect 11734 8420 11808 8476
rect 11468 8334 11808 8420
rect 11468 8278 11536 8334
rect 11592 8278 11678 8334
rect 11734 8278 11808 8334
rect 11468 8192 11808 8278
rect 11468 8136 11536 8192
rect 11592 8136 11678 8192
rect 11734 8136 11808 8192
rect 11468 8050 11808 8136
rect 11468 7994 11536 8050
rect 11592 7994 11678 8050
rect 11734 7994 11808 8050
rect 11468 7908 11808 7994
rect 11468 7852 11536 7908
rect 11592 7852 11678 7908
rect 11734 7852 11808 7908
rect 11468 7766 11808 7852
rect 11468 7710 11536 7766
rect 11592 7710 11678 7766
rect 11734 7710 11808 7766
rect 11468 7624 11808 7710
rect 11468 7568 11536 7624
rect 11592 7568 11678 7624
rect 11734 7568 11808 7624
rect 11468 7482 11808 7568
rect 11468 7426 11536 7482
rect 11592 7426 11678 7482
rect 11734 7426 11808 7482
rect 11468 7340 11808 7426
rect 11468 7284 11536 7340
rect 11592 7284 11678 7340
rect 11734 7284 11808 7340
rect 11468 7198 11808 7284
rect 11468 7142 11536 7198
rect 11592 7142 11678 7198
rect 11734 7142 11808 7198
rect 11468 7056 11808 7142
rect 11468 7000 11536 7056
rect 11592 7000 11678 7056
rect 11734 7000 11808 7056
rect 11468 6914 11808 7000
rect 11468 6858 11536 6914
rect 11592 6858 11678 6914
rect 11734 6858 11808 6914
rect 11468 6772 11808 6858
rect 11468 6716 11536 6772
rect 11592 6716 11678 6772
rect 11734 6716 11808 6772
rect 11468 6630 11808 6716
rect 11468 6574 11536 6630
rect 11592 6574 11678 6630
rect 11734 6574 11808 6630
rect 11468 6488 11808 6574
rect 11468 6432 11536 6488
rect 11592 6432 11678 6488
rect 11734 6432 11808 6488
rect 11468 6346 11808 6432
rect 11468 6290 11536 6346
rect 11592 6290 11678 6346
rect 11734 6290 11808 6346
rect 11468 6204 11808 6290
rect 11468 6148 11536 6204
rect 11592 6148 11678 6204
rect 11734 6148 11808 6204
rect 11468 6062 11808 6148
rect 11468 6006 11536 6062
rect 11592 6006 11678 6062
rect 11734 6006 11808 6062
rect 11468 5920 11808 6006
rect 11468 5864 11536 5920
rect 11592 5864 11678 5920
rect 11734 5864 11808 5920
rect 11468 5778 11808 5864
rect 11468 5722 11536 5778
rect 11592 5722 11678 5778
rect 11734 5722 11808 5778
rect 11468 5636 11808 5722
rect 11468 5580 11536 5636
rect 11592 5580 11678 5636
rect 11734 5580 11808 5636
rect 11468 5494 11808 5580
rect 11468 5438 11536 5494
rect 11592 5438 11678 5494
rect 11734 5438 11808 5494
rect 11468 5352 11808 5438
rect 11468 5296 11536 5352
rect 11592 5296 11678 5352
rect 11734 5296 11808 5352
rect 11468 5210 11808 5296
rect 11468 5154 11536 5210
rect 11592 5154 11678 5210
rect 11734 5154 11808 5210
rect 11468 5068 11808 5154
rect 11468 5012 11536 5068
rect 11592 5012 11678 5068
rect 11734 5012 11808 5068
rect 11468 4926 11808 5012
rect 11468 4870 11536 4926
rect 11592 4870 11678 4926
rect 11734 4870 11808 4926
rect 11468 4784 11808 4870
rect 11468 4728 11536 4784
rect 11592 4728 11678 4784
rect 11734 4728 11808 4784
rect 11468 4642 11808 4728
rect 11468 4586 11536 4642
rect 11592 4586 11678 4642
rect 11734 4586 11808 4642
rect 11468 4500 11808 4586
rect 11468 4444 11536 4500
rect 11592 4444 11678 4500
rect 11734 4444 11808 4500
rect 11468 4358 11808 4444
rect 11468 4302 11536 4358
rect 11592 4302 11678 4358
rect 11734 4302 11808 4358
rect 11468 4216 11808 4302
rect 11468 4160 11536 4216
rect 11592 4160 11678 4216
rect 11734 4160 11808 4216
rect 11468 4074 11808 4160
rect 11468 4018 11536 4074
rect 11592 4018 11678 4074
rect 11734 4018 11808 4074
rect 11468 3932 11808 4018
rect 11468 3876 11536 3932
rect 11592 3876 11678 3932
rect 11734 3876 11808 3932
rect 11468 3790 11808 3876
rect 11468 3734 11536 3790
rect 11592 3734 11678 3790
rect 11734 3734 11808 3790
rect 11468 3648 11808 3734
rect 11468 3592 11536 3648
rect 11592 3592 11678 3648
rect 11734 3592 11808 3648
rect 11468 3506 11808 3592
rect 11468 3450 11536 3506
rect 11592 3450 11678 3506
rect 11734 3450 11808 3506
rect 11468 3364 11808 3450
rect 11468 3308 11536 3364
rect 11592 3308 11678 3364
rect 11734 3308 11808 3364
rect 11468 3222 11808 3308
rect 11468 3166 11536 3222
rect 11592 3166 11678 3222
rect 11734 3166 11808 3222
rect 11468 3080 11808 3166
rect 11468 3024 11536 3080
rect 11592 3024 11678 3080
rect 11734 3024 11808 3080
rect 11468 2938 11808 3024
rect 11468 2882 11536 2938
rect 11592 2882 11678 2938
rect 11734 2882 11808 2938
rect 11468 2796 11808 2882
rect 11468 2740 11536 2796
rect 11592 2740 11678 2796
rect 11734 2740 11808 2796
rect 11468 2654 11808 2740
rect 11468 2598 11536 2654
rect 11592 2598 11678 2654
rect 11734 2598 11808 2654
rect 11468 2512 11808 2598
rect 11468 2456 11536 2512
rect 11592 2456 11678 2512
rect 11734 2456 11808 2512
rect 11468 2370 11808 2456
rect 11468 2314 11536 2370
rect 11592 2314 11678 2370
rect 11734 2314 11808 2370
rect 11468 2228 11808 2314
rect 11468 2172 11536 2228
rect 11592 2172 11678 2228
rect 11734 2172 11808 2228
rect 11468 2086 11808 2172
rect 11468 2030 11536 2086
rect 11592 2030 11678 2086
rect 11734 2030 11808 2086
rect 11468 1944 11808 2030
rect 11468 1888 11536 1944
rect 11592 1888 11678 1944
rect 11734 1888 11808 1944
rect 11468 1802 11808 1888
rect 11468 1746 11536 1802
rect 11592 1746 11678 1802
rect 11734 1746 11808 1802
rect 11468 1660 11808 1746
rect 11468 1604 11536 1660
rect 11592 1604 11678 1660
rect 11734 1604 11808 1660
rect 11468 1518 11808 1604
rect 11468 1462 11536 1518
rect 11592 1462 11678 1518
rect 11734 1462 11808 1518
rect 11468 1376 11808 1462
rect 11468 1320 11536 1376
rect 11592 1320 11678 1376
rect 11734 1320 11808 1376
rect 11468 1234 11808 1320
rect 11468 1178 11536 1234
rect 11592 1178 11678 1234
rect 11734 1178 11808 1234
rect 11468 1092 11808 1178
rect 11468 1036 11536 1092
rect 11592 1036 11678 1092
rect 11734 1036 11808 1092
rect 11468 950 11808 1036
rect 11468 894 11536 950
rect 11592 894 11678 950
rect 11734 894 11808 950
rect 11468 808 11808 894
rect 11468 752 11536 808
rect 11592 752 11678 808
rect 11734 752 11808 808
rect 11468 666 11808 752
rect 11468 610 11536 666
rect 11592 610 11678 666
rect 11734 610 11808 666
rect 11468 524 11808 610
rect 11468 468 11536 524
rect 11592 468 11678 524
rect 11734 468 11808 524
rect 11468 400 11808 468
rect 11868 12310 12208 12400
rect 11868 12254 11941 12310
rect 11997 12254 12083 12310
rect 12139 12254 12208 12310
rect 11868 12168 12208 12254
rect 11868 12112 11941 12168
rect 11997 12112 12083 12168
rect 12139 12112 12208 12168
rect 11868 12026 12208 12112
rect 11868 11970 11941 12026
rect 11997 11970 12083 12026
rect 12139 11970 12208 12026
rect 11868 11884 12208 11970
rect 11868 11828 11941 11884
rect 11997 11828 12083 11884
rect 12139 11828 12208 11884
rect 11868 11742 12208 11828
rect 11868 11686 11941 11742
rect 11997 11686 12083 11742
rect 12139 11686 12208 11742
rect 11868 11600 12208 11686
rect 11868 11544 11941 11600
rect 11997 11544 12083 11600
rect 12139 11544 12208 11600
rect 11868 11458 12208 11544
rect 11868 11402 11941 11458
rect 11997 11402 12083 11458
rect 12139 11402 12208 11458
rect 11868 11316 12208 11402
rect 11868 11260 11941 11316
rect 11997 11260 12083 11316
rect 12139 11260 12208 11316
rect 11868 11174 12208 11260
rect 11868 11118 11941 11174
rect 11997 11118 12083 11174
rect 12139 11118 12208 11174
rect 11868 11032 12208 11118
rect 11868 10976 11941 11032
rect 11997 10976 12083 11032
rect 12139 10976 12208 11032
rect 11868 10890 12208 10976
rect 11868 10834 11941 10890
rect 11997 10834 12083 10890
rect 12139 10834 12208 10890
rect 11868 10748 12208 10834
rect 11868 10692 11941 10748
rect 11997 10692 12083 10748
rect 12139 10692 12208 10748
rect 11868 10606 12208 10692
rect 11868 10550 11941 10606
rect 11997 10550 12083 10606
rect 12139 10550 12208 10606
rect 11868 10464 12208 10550
rect 11868 10408 11941 10464
rect 11997 10408 12083 10464
rect 12139 10408 12208 10464
rect 11868 10322 12208 10408
rect 11868 10266 11941 10322
rect 11997 10266 12083 10322
rect 12139 10266 12208 10322
rect 11868 10180 12208 10266
rect 11868 10124 11941 10180
rect 11997 10124 12083 10180
rect 12139 10124 12208 10180
rect 11868 10038 12208 10124
rect 11868 9982 11941 10038
rect 11997 9982 12083 10038
rect 12139 9982 12208 10038
rect 11868 9896 12208 9982
rect 11868 9840 11941 9896
rect 11997 9840 12083 9896
rect 12139 9840 12208 9896
rect 11868 9754 12208 9840
rect 11868 9698 11941 9754
rect 11997 9698 12083 9754
rect 12139 9698 12208 9754
rect 11868 9612 12208 9698
rect 11868 9556 11941 9612
rect 11997 9556 12083 9612
rect 12139 9556 12208 9612
rect 11868 9470 12208 9556
rect 11868 9414 11941 9470
rect 11997 9414 12083 9470
rect 12139 9414 12208 9470
rect 11868 9328 12208 9414
rect 11868 9272 11941 9328
rect 11997 9272 12083 9328
rect 12139 9272 12208 9328
rect 11868 9186 12208 9272
rect 11868 9130 11941 9186
rect 11997 9130 12083 9186
rect 12139 9130 12208 9186
rect 11868 9044 12208 9130
rect 11868 8988 11941 9044
rect 11997 8988 12083 9044
rect 12139 8988 12208 9044
rect 11868 8902 12208 8988
rect 11868 8846 11941 8902
rect 11997 8846 12083 8902
rect 12139 8846 12208 8902
rect 11868 8760 12208 8846
rect 11868 8704 11941 8760
rect 11997 8704 12083 8760
rect 12139 8704 12208 8760
rect 11868 8618 12208 8704
rect 11868 8562 11941 8618
rect 11997 8562 12083 8618
rect 12139 8562 12208 8618
rect 11868 8476 12208 8562
rect 11868 8420 11941 8476
rect 11997 8420 12083 8476
rect 12139 8420 12208 8476
rect 11868 8334 12208 8420
rect 11868 8278 11941 8334
rect 11997 8278 12083 8334
rect 12139 8278 12208 8334
rect 11868 8192 12208 8278
rect 11868 8136 11941 8192
rect 11997 8136 12083 8192
rect 12139 8136 12208 8192
rect 11868 8050 12208 8136
rect 11868 7994 11941 8050
rect 11997 7994 12083 8050
rect 12139 7994 12208 8050
rect 11868 7908 12208 7994
rect 11868 7852 11941 7908
rect 11997 7852 12083 7908
rect 12139 7852 12208 7908
rect 11868 7766 12208 7852
rect 11868 7710 11941 7766
rect 11997 7710 12083 7766
rect 12139 7710 12208 7766
rect 11868 7624 12208 7710
rect 11868 7568 11941 7624
rect 11997 7568 12083 7624
rect 12139 7568 12208 7624
rect 11868 7482 12208 7568
rect 11868 7426 11941 7482
rect 11997 7426 12083 7482
rect 12139 7426 12208 7482
rect 11868 7340 12208 7426
rect 11868 7284 11941 7340
rect 11997 7284 12083 7340
rect 12139 7284 12208 7340
rect 11868 7198 12208 7284
rect 11868 7142 11941 7198
rect 11997 7142 12083 7198
rect 12139 7142 12208 7198
rect 11868 7056 12208 7142
rect 11868 7000 11941 7056
rect 11997 7000 12083 7056
rect 12139 7000 12208 7056
rect 11868 6914 12208 7000
rect 11868 6858 11941 6914
rect 11997 6858 12083 6914
rect 12139 6858 12208 6914
rect 11868 6772 12208 6858
rect 11868 6716 11941 6772
rect 11997 6716 12083 6772
rect 12139 6716 12208 6772
rect 11868 6630 12208 6716
rect 11868 6574 11941 6630
rect 11997 6574 12083 6630
rect 12139 6574 12208 6630
rect 11868 6488 12208 6574
rect 11868 6432 11941 6488
rect 11997 6432 12083 6488
rect 12139 6432 12208 6488
rect 11868 6346 12208 6432
rect 11868 6290 11941 6346
rect 11997 6290 12083 6346
rect 12139 6290 12208 6346
rect 11868 6204 12208 6290
rect 11868 6148 11941 6204
rect 11997 6148 12083 6204
rect 12139 6148 12208 6204
rect 11868 6062 12208 6148
rect 11868 6006 11941 6062
rect 11997 6006 12083 6062
rect 12139 6006 12208 6062
rect 11868 5920 12208 6006
rect 11868 5864 11941 5920
rect 11997 5864 12083 5920
rect 12139 5864 12208 5920
rect 11868 5778 12208 5864
rect 11868 5722 11941 5778
rect 11997 5722 12083 5778
rect 12139 5722 12208 5778
rect 11868 5636 12208 5722
rect 11868 5580 11941 5636
rect 11997 5580 12083 5636
rect 12139 5580 12208 5636
rect 11868 5494 12208 5580
rect 11868 5438 11941 5494
rect 11997 5438 12083 5494
rect 12139 5438 12208 5494
rect 11868 5352 12208 5438
rect 11868 5296 11941 5352
rect 11997 5296 12083 5352
rect 12139 5296 12208 5352
rect 11868 5210 12208 5296
rect 11868 5154 11941 5210
rect 11997 5154 12083 5210
rect 12139 5154 12208 5210
rect 11868 5068 12208 5154
rect 11868 5012 11941 5068
rect 11997 5012 12083 5068
rect 12139 5012 12208 5068
rect 11868 4926 12208 5012
rect 11868 4870 11941 4926
rect 11997 4870 12083 4926
rect 12139 4870 12208 4926
rect 11868 4784 12208 4870
rect 11868 4728 11941 4784
rect 11997 4728 12083 4784
rect 12139 4728 12208 4784
rect 11868 4642 12208 4728
rect 11868 4586 11941 4642
rect 11997 4586 12083 4642
rect 12139 4586 12208 4642
rect 11868 4500 12208 4586
rect 11868 4444 11941 4500
rect 11997 4444 12083 4500
rect 12139 4444 12208 4500
rect 11868 4358 12208 4444
rect 11868 4302 11941 4358
rect 11997 4302 12083 4358
rect 12139 4302 12208 4358
rect 11868 4216 12208 4302
rect 11868 4160 11941 4216
rect 11997 4160 12083 4216
rect 12139 4160 12208 4216
rect 11868 4074 12208 4160
rect 11868 4018 11941 4074
rect 11997 4018 12083 4074
rect 12139 4018 12208 4074
rect 11868 3932 12208 4018
rect 11868 3876 11941 3932
rect 11997 3876 12083 3932
rect 12139 3876 12208 3932
rect 11868 3790 12208 3876
rect 11868 3734 11941 3790
rect 11997 3734 12083 3790
rect 12139 3734 12208 3790
rect 11868 3648 12208 3734
rect 11868 3592 11941 3648
rect 11997 3592 12083 3648
rect 12139 3592 12208 3648
rect 11868 3506 12208 3592
rect 11868 3450 11941 3506
rect 11997 3450 12083 3506
rect 12139 3450 12208 3506
rect 11868 3364 12208 3450
rect 11868 3308 11941 3364
rect 11997 3308 12083 3364
rect 12139 3308 12208 3364
rect 11868 3222 12208 3308
rect 11868 3166 11941 3222
rect 11997 3166 12083 3222
rect 12139 3166 12208 3222
rect 11868 3080 12208 3166
rect 11868 3024 11941 3080
rect 11997 3024 12083 3080
rect 12139 3024 12208 3080
rect 11868 2938 12208 3024
rect 11868 2882 11941 2938
rect 11997 2882 12083 2938
rect 12139 2882 12208 2938
rect 11868 2796 12208 2882
rect 11868 2740 11941 2796
rect 11997 2740 12083 2796
rect 12139 2740 12208 2796
rect 11868 2654 12208 2740
rect 11868 2598 11941 2654
rect 11997 2598 12083 2654
rect 12139 2598 12208 2654
rect 11868 2512 12208 2598
rect 11868 2456 11941 2512
rect 11997 2456 12083 2512
rect 12139 2456 12208 2512
rect 11868 2370 12208 2456
rect 11868 2314 11941 2370
rect 11997 2314 12083 2370
rect 12139 2314 12208 2370
rect 11868 2228 12208 2314
rect 11868 2172 11941 2228
rect 11997 2172 12083 2228
rect 12139 2172 12208 2228
rect 11868 2086 12208 2172
rect 11868 2030 11941 2086
rect 11997 2030 12083 2086
rect 12139 2030 12208 2086
rect 11868 1944 12208 2030
rect 11868 1888 11941 1944
rect 11997 1888 12083 1944
rect 12139 1888 12208 1944
rect 11868 1802 12208 1888
rect 11868 1746 11941 1802
rect 11997 1746 12083 1802
rect 12139 1746 12208 1802
rect 11868 1660 12208 1746
rect 11868 1604 11941 1660
rect 11997 1604 12083 1660
rect 12139 1604 12208 1660
rect 11868 1518 12208 1604
rect 11868 1462 11941 1518
rect 11997 1462 12083 1518
rect 12139 1462 12208 1518
rect 11868 1376 12208 1462
rect 11868 1320 11941 1376
rect 11997 1320 12083 1376
rect 12139 1320 12208 1376
rect 11868 1234 12208 1320
rect 11868 1178 11941 1234
rect 11997 1178 12083 1234
rect 12139 1178 12208 1234
rect 11868 1092 12208 1178
rect 11868 1036 11941 1092
rect 11997 1036 12083 1092
rect 12139 1036 12208 1092
rect 11868 950 12208 1036
rect 11868 894 11941 950
rect 11997 894 12083 950
rect 12139 894 12208 950
rect 11868 808 12208 894
rect 11868 752 11941 808
rect 11997 752 12083 808
rect 12139 752 12208 808
rect 11868 666 12208 752
rect 11868 610 11941 666
rect 11997 610 12083 666
rect 12139 610 12208 666
rect 11868 524 12208 610
rect 11868 468 11941 524
rect 11997 468 12083 524
rect 12139 468 12208 524
rect 11868 400 12208 468
rect 12400 12358 13200 12400
rect 12400 12302 12526 12358
rect 12582 12302 12650 12358
rect 12706 12302 12774 12358
rect 12830 12302 12898 12358
rect 12954 12302 13022 12358
rect 13078 12302 13200 12358
rect 12400 12234 13200 12302
rect 12400 12178 12526 12234
rect 12582 12178 12650 12234
rect 12706 12178 12774 12234
rect 12830 12178 12898 12234
rect 12954 12178 13022 12234
rect 13078 12178 13200 12234
rect 12400 12110 13200 12178
rect 12400 12054 12526 12110
rect 12582 12054 12650 12110
rect 12706 12054 12774 12110
rect 12830 12054 12898 12110
rect 12954 12054 13022 12110
rect 13078 12054 13200 12110
rect 12400 11986 13200 12054
rect 12400 11930 12526 11986
rect 12582 11930 12650 11986
rect 12706 11930 12774 11986
rect 12830 11930 12898 11986
rect 12954 11930 13022 11986
rect 13078 11930 13200 11986
rect 12400 11862 13200 11930
rect 12400 11806 12526 11862
rect 12582 11806 12650 11862
rect 12706 11806 12774 11862
rect 12830 11806 12898 11862
rect 12954 11806 13022 11862
rect 13078 11806 13200 11862
rect 12400 11738 13200 11806
rect 12400 11682 12526 11738
rect 12582 11682 12650 11738
rect 12706 11682 12774 11738
rect 12830 11682 12898 11738
rect 12954 11682 13022 11738
rect 13078 11682 13200 11738
rect 12400 11614 13200 11682
rect 12400 11558 12526 11614
rect 12582 11558 12650 11614
rect 12706 11558 12774 11614
rect 12830 11558 12898 11614
rect 12954 11558 13022 11614
rect 13078 11558 13200 11614
rect 12400 11490 13200 11558
rect 12400 11434 12526 11490
rect 12582 11434 12650 11490
rect 12706 11434 12774 11490
rect 12830 11434 12898 11490
rect 12954 11434 13022 11490
rect 13078 11434 13200 11490
rect 12400 11366 13200 11434
rect 12400 11310 12526 11366
rect 12582 11310 12650 11366
rect 12706 11310 12774 11366
rect 12830 11310 12898 11366
rect 12954 11310 13022 11366
rect 13078 11310 13200 11366
rect 12400 11242 13200 11310
rect 12400 11186 12526 11242
rect 12582 11186 12650 11242
rect 12706 11186 12774 11242
rect 12830 11186 12898 11242
rect 12954 11186 13022 11242
rect 13078 11186 13200 11242
rect 12400 11118 13200 11186
rect 12400 11062 12526 11118
rect 12582 11062 12650 11118
rect 12706 11062 12774 11118
rect 12830 11062 12898 11118
rect 12954 11062 13022 11118
rect 13078 11062 13200 11118
rect 12400 10994 13200 11062
rect 12400 10938 12526 10994
rect 12582 10938 12650 10994
rect 12706 10938 12774 10994
rect 12830 10938 12898 10994
rect 12954 10938 13022 10994
rect 13078 10938 13200 10994
rect 12400 10870 13200 10938
rect 12400 10814 12526 10870
rect 12582 10814 12650 10870
rect 12706 10814 12774 10870
rect 12830 10814 12898 10870
rect 12954 10814 13022 10870
rect 13078 10814 13200 10870
rect 12400 10746 13200 10814
rect 12400 10690 12526 10746
rect 12582 10690 12650 10746
rect 12706 10690 12774 10746
rect 12830 10690 12898 10746
rect 12954 10690 13022 10746
rect 13078 10690 13200 10746
rect 12400 10622 13200 10690
rect 12400 10566 12526 10622
rect 12582 10566 12650 10622
rect 12706 10566 12774 10622
rect 12830 10566 12898 10622
rect 12954 10566 13022 10622
rect 13078 10566 13200 10622
rect 12400 10498 13200 10566
rect 12400 10442 12526 10498
rect 12582 10442 12650 10498
rect 12706 10442 12774 10498
rect 12830 10442 12898 10498
rect 12954 10442 13022 10498
rect 13078 10442 13200 10498
rect 12400 10374 13200 10442
rect 12400 10318 12526 10374
rect 12582 10318 12650 10374
rect 12706 10318 12774 10374
rect 12830 10318 12898 10374
rect 12954 10318 13022 10374
rect 13078 10318 13200 10374
rect 12400 10250 13200 10318
rect 12400 10194 12526 10250
rect 12582 10194 12650 10250
rect 12706 10194 12774 10250
rect 12830 10194 12898 10250
rect 12954 10194 13022 10250
rect 13078 10194 13200 10250
rect 12400 10126 13200 10194
rect 12400 10070 12526 10126
rect 12582 10070 12650 10126
rect 12706 10070 12774 10126
rect 12830 10070 12898 10126
rect 12954 10070 13022 10126
rect 13078 10070 13200 10126
rect 12400 10002 13200 10070
rect 12400 9946 12526 10002
rect 12582 9946 12650 10002
rect 12706 9946 12774 10002
rect 12830 9946 12898 10002
rect 12954 9946 13022 10002
rect 13078 9946 13200 10002
rect 12400 9878 13200 9946
rect 12400 9822 12526 9878
rect 12582 9822 12650 9878
rect 12706 9822 12774 9878
rect 12830 9822 12898 9878
rect 12954 9822 13022 9878
rect 13078 9822 13200 9878
rect 12400 9754 13200 9822
rect 12400 9698 12526 9754
rect 12582 9698 12650 9754
rect 12706 9698 12774 9754
rect 12830 9698 12898 9754
rect 12954 9698 13022 9754
rect 13078 9698 13200 9754
rect 12400 9630 13200 9698
rect 12400 9574 12526 9630
rect 12582 9574 12650 9630
rect 12706 9574 12774 9630
rect 12830 9574 12898 9630
rect 12954 9574 13022 9630
rect 13078 9574 13200 9630
rect 12400 9506 13200 9574
rect 12400 9450 12526 9506
rect 12582 9450 12650 9506
rect 12706 9450 12774 9506
rect 12830 9450 12898 9506
rect 12954 9450 13022 9506
rect 13078 9450 13200 9506
rect 12400 9382 13200 9450
rect 12400 9326 12526 9382
rect 12582 9326 12650 9382
rect 12706 9326 12774 9382
rect 12830 9326 12898 9382
rect 12954 9326 13022 9382
rect 13078 9326 13200 9382
rect 12400 9258 13200 9326
rect 12400 9202 12526 9258
rect 12582 9202 12650 9258
rect 12706 9202 12774 9258
rect 12830 9202 12898 9258
rect 12954 9202 13022 9258
rect 13078 9202 13200 9258
rect 12400 9134 13200 9202
rect 12400 9078 12526 9134
rect 12582 9078 12650 9134
rect 12706 9078 12774 9134
rect 12830 9078 12898 9134
rect 12954 9078 13022 9134
rect 13078 9078 13200 9134
rect 12400 9010 13200 9078
rect 12400 8954 12526 9010
rect 12582 8954 12650 9010
rect 12706 8954 12774 9010
rect 12830 8954 12898 9010
rect 12954 8954 13022 9010
rect 13078 8954 13200 9010
rect 12400 8886 13200 8954
rect 12400 8830 12526 8886
rect 12582 8830 12650 8886
rect 12706 8830 12774 8886
rect 12830 8830 12898 8886
rect 12954 8830 13022 8886
rect 13078 8830 13200 8886
rect 12400 8762 13200 8830
rect 12400 8706 12526 8762
rect 12582 8706 12650 8762
rect 12706 8706 12774 8762
rect 12830 8706 12898 8762
rect 12954 8706 13022 8762
rect 13078 8706 13200 8762
rect 12400 8638 13200 8706
rect 12400 8582 12526 8638
rect 12582 8582 12650 8638
rect 12706 8582 12774 8638
rect 12830 8582 12898 8638
rect 12954 8582 13022 8638
rect 13078 8582 13200 8638
rect 12400 8514 13200 8582
rect 12400 8458 12526 8514
rect 12582 8458 12650 8514
rect 12706 8458 12774 8514
rect 12830 8458 12898 8514
rect 12954 8458 13022 8514
rect 13078 8458 13200 8514
rect 12400 8390 13200 8458
rect 12400 8334 12526 8390
rect 12582 8334 12650 8390
rect 12706 8334 12774 8390
rect 12830 8334 12898 8390
rect 12954 8334 13022 8390
rect 13078 8334 13200 8390
rect 12400 8266 13200 8334
rect 12400 8210 12526 8266
rect 12582 8210 12650 8266
rect 12706 8210 12774 8266
rect 12830 8210 12898 8266
rect 12954 8210 13022 8266
rect 13078 8210 13200 8266
rect 12400 8142 13200 8210
rect 12400 8086 12526 8142
rect 12582 8086 12650 8142
rect 12706 8086 12774 8142
rect 12830 8086 12898 8142
rect 12954 8086 13022 8142
rect 13078 8086 13200 8142
rect 12400 8018 13200 8086
rect 12400 7962 12526 8018
rect 12582 7962 12650 8018
rect 12706 7962 12774 8018
rect 12830 7962 12898 8018
rect 12954 7962 13022 8018
rect 13078 7962 13200 8018
rect 12400 7894 13200 7962
rect 12400 7838 12526 7894
rect 12582 7838 12650 7894
rect 12706 7838 12774 7894
rect 12830 7838 12898 7894
rect 12954 7838 13022 7894
rect 13078 7838 13200 7894
rect 12400 7770 13200 7838
rect 12400 7714 12526 7770
rect 12582 7714 12650 7770
rect 12706 7714 12774 7770
rect 12830 7714 12898 7770
rect 12954 7714 13022 7770
rect 13078 7714 13200 7770
rect 12400 7646 13200 7714
rect 12400 7590 12526 7646
rect 12582 7590 12650 7646
rect 12706 7590 12774 7646
rect 12830 7590 12898 7646
rect 12954 7590 13022 7646
rect 13078 7590 13200 7646
rect 12400 7522 13200 7590
rect 12400 7466 12526 7522
rect 12582 7466 12650 7522
rect 12706 7466 12774 7522
rect 12830 7466 12898 7522
rect 12954 7466 13022 7522
rect 13078 7466 13200 7522
rect 12400 7398 13200 7466
rect 12400 7342 12526 7398
rect 12582 7342 12650 7398
rect 12706 7342 12774 7398
rect 12830 7342 12898 7398
rect 12954 7342 13022 7398
rect 13078 7342 13200 7398
rect 12400 7274 13200 7342
rect 12400 7218 12526 7274
rect 12582 7218 12650 7274
rect 12706 7218 12774 7274
rect 12830 7218 12898 7274
rect 12954 7218 13022 7274
rect 13078 7218 13200 7274
rect 12400 7150 13200 7218
rect 12400 7094 12526 7150
rect 12582 7094 12650 7150
rect 12706 7094 12774 7150
rect 12830 7094 12898 7150
rect 12954 7094 13022 7150
rect 13078 7094 13200 7150
rect 12400 7026 13200 7094
rect 12400 6970 12526 7026
rect 12582 6970 12650 7026
rect 12706 6970 12774 7026
rect 12830 6970 12898 7026
rect 12954 6970 13022 7026
rect 13078 6970 13200 7026
rect 12400 6902 13200 6970
rect 12400 6846 12526 6902
rect 12582 6846 12650 6902
rect 12706 6846 12774 6902
rect 12830 6846 12898 6902
rect 12954 6846 13022 6902
rect 13078 6846 13200 6902
rect 12400 6778 13200 6846
rect 12400 6722 12526 6778
rect 12582 6722 12650 6778
rect 12706 6722 12774 6778
rect 12830 6722 12898 6778
rect 12954 6722 13022 6778
rect 13078 6722 13200 6778
rect 12400 6654 13200 6722
rect 12400 6598 12526 6654
rect 12582 6598 12650 6654
rect 12706 6598 12774 6654
rect 12830 6598 12898 6654
rect 12954 6598 13022 6654
rect 13078 6598 13200 6654
rect 12400 6530 13200 6598
rect 12400 6474 12526 6530
rect 12582 6474 12650 6530
rect 12706 6474 12774 6530
rect 12830 6474 12898 6530
rect 12954 6474 13022 6530
rect 13078 6474 13200 6530
rect 12400 6406 13200 6474
rect 12400 6350 12526 6406
rect 12582 6350 12650 6406
rect 12706 6350 12774 6406
rect 12830 6350 12898 6406
rect 12954 6350 13022 6406
rect 13078 6350 13200 6406
rect 12400 6282 13200 6350
rect 12400 6226 12526 6282
rect 12582 6226 12650 6282
rect 12706 6226 12774 6282
rect 12830 6226 12898 6282
rect 12954 6226 13022 6282
rect 13078 6226 13200 6282
rect 12400 6158 13200 6226
rect 12400 6102 12526 6158
rect 12582 6102 12650 6158
rect 12706 6102 12774 6158
rect 12830 6102 12898 6158
rect 12954 6102 13022 6158
rect 13078 6102 13200 6158
rect 12400 6034 13200 6102
rect 12400 5978 12526 6034
rect 12582 5978 12650 6034
rect 12706 5978 12774 6034
rect 12830 5978 12898 6034
rect 12954 5978 13022 6034
rect 13078 5978 13200 6034
rect 12400 5910 13200 5978
rect 12400 5854 12526 5910
rect 12582 5854 12650 5910
rect 12706 5854 12774 5910
rect 12830 5854 12898 5910
rect 12954 5854 13022 5910
rect 13078 5854 13200 5910
rect 12400 5786 13200 5854
rect 12400 5730 12526 5786
rect 12582 5730 12650 5786
rect 12706 5730 12774 5786
rect 12830 5730 12898 5786
rect 12954 5730 13022 5786
rect 13078 5730 13200 5786
rect 12400 5662 13200 5730
rect 12400 5606 12526 5662
rect 12582 5606 12650 5662
rect 12706 5606 12774 5662
rect 12830 5606 12898 5662
rect 12954 5606 13022 5662
rect 13078 5606 13200 5662
rect 12400 5538 13200 5606
rect 12400 5482 12526 5538
rect 12582 5482 12650 5538
rect 12706 5482 12774 5538
rect 12830 5482 12898 5538
rect 12954 5482 13022 5538
rect 13078 5482 13200 5538
rect 12400 5414 13200 5482
rect 12400 5358 12526 5414
rect 12582 5358 12650 5414
rect 12706 5358 12774 5414
rect 12830 5358 12898 5414
rect 12954 5358 13022 5414
rect 13078 5358 13200 5414
rect 12400 5290 13200 5358
rect 12400 5234 12526 5290
rect 12582 5234 12650 5290
rect 12706 5234 12774 5290
rect 12830 5234 12898 5290
rect 12954 5234 13022 5290
rect 13078 5234 13200 5290
rect 12400 5166 13200 5234
rect 12400 5110 12526 5166
rect 12582 5110 12650 5166
rect 12706 5110 12774 5166
rect 12830 5110 12898 5166
rect 12954 5110 13022 5166
rect 13078 5110 13200 5166
rect 12400 5042 13200 5110
rect 12400 4986 12526 5042
rect 12582 4986 12650 5042
rect 12706 4986 12774 5042
rect 12830 4986 12898 5042
rect 12954 4986 13022 5042
rect 13078 4986 13200 5042
rect 12400 4918 13200 4986
rect 12400 4862 12526 4918
rect 12582 4862 12650 4918
rect 12706 4862 12774 4918
rect 12830 4862 12898 4918
rect 12954 4862 13022 4918
rect 13078 4862 13200 4918
rect 12400 4794 13200 4862
rect 12400 4738 12526 4794
rect 12582 4738 12650 4794
rect 12706 4738 12774 4794
rect 12830 4738 12898 4794
rect 12954 4738 13022 4794
rect 13078 4738 13200 4794
rect 12400 4670 13200 4738
rect 12400 4614 12526 4670
rect 12582 4614 12650 4670
rect 12706 4614 12774 4670
rect 12830 4614 12898 4670
rect 12954 4614 13022 4670
rect 13078 4614 13200 4670
rect 12400 4546 13200 4614
rect 12400 4490 12526 4546
rect 12582 4490 12650 4546
rect 12706 4490 12774 4546
rect 12830 4490 12898 4546
rect 12954 4490 13022 4546
rect 13078 4490 13200 4546
rect 12400 4422 13200 4490
rect 12400 4366 12526 4422
rect 12582 4366 12650 4422
rect 12706 4366 12774 4422
rect 12830 4366 12898 4422
rect 12954 4366 13022 4422
rect 13078 4366 13200 4422
rect 12400 4298 13200 4366
rect 12400 4242 12526 4298
rect 12582 4242 12650 4298
rect 12706 4242 12774 4298
rect 12830 4242 12898 4298
rect 12954 4242 13022 4298
rect 13078 4242 13200 4298
rect 12400 4174 13200 4242
rect 12400 4118 12526 4174
rect 12582 4118 12650 4174
rect 12706 4118 12774 4174
rect 12830 4118 12898 4174
rect 12954 4118 13022 4174
rect 13078 4118 13200 4174
rect 12400 4050 13200 4118
rect 12400 3994 12526 4050
rect 12582 3994 12650 4050
rect 12706 3994 12774 4050
rect 12830 3994 12898 4050
rect 12954 3994 13022 4050
rect 13078 3994 13200 4050
rect 12400 3926 13200 3994
rect 12400 3870 12526 3926
rect 12582 3870 12650 3926
rect 12706 3870 12774 3926
rect 12830 3870 12898 3926
rect 12954 3870 13022 3926
rect 13078 3870 13200 3926
rect 12400 3802 13200 3870
rect 12400 3746 12526 3802
rect 12582 3746 12650 3802
rect 12706 3746 12774 3802
rect 12830 3746 12898 3802
rect 12954 3746 13022 3802
rect 13078 3746 13200 3802
rect 12400 3678 13200 3746
rect 12400 3622 12526 3678
rect 12582 3622 12650 3678
rect 12706 3622 12774 3678
rect 12830 3622 12898 3678
rect 12954 3622 13022 3678
rect 13078 3622 13200 3678
rect 12400 3554 13200 3622
rect 12400 3498 12526 3554
rect 12582 3498 12650 3554
rect 12706 3498 12774 3554
rect 12830 3498 12898 3554
rect 12954 3498 13022 3554
rect 13078 3498 13200 3554
rect 12400 3430 13200 3498
rect 12400 3374 12526 3430
rect 12582 3374 12650 3430
rect 12706 3374 12774 3430
rect 12830 3374 12898 3430
rect 12954 3374 13022 3430
rect 13078 3374 13200 3430
rect 12400 3306 13200 3374
rect 12400 3250 12526 3306
rect 12582 3250 12650 3306
rect 12706 3250 12774 3306
rect 12830 3250 12898 3306
rect 12954 3250 13022 3306
rect 13078 3250 13200 3306
rect 12400 3182 13200 3250
rect 12400 3126 12526 3182
rect 12582 3126 12650 3182
rect 12706 3126 12774 3182
rect 12830 3126 12898 3182
rect 12954 3126 13022 3182
rect 13078 3126 13200 3182
rect 12400 3058 13200 3126
rect 12400 3002 12526 3058
rect 12582 3002 12650 3058
rect 12706 3002 12774 3058
rect 12830 3002 12898 3058
rect 12954 3002 13022 3058
rect 13078 3002 13200 3058
rect 12400 2934 13200 3002
rect 12400 2878 12526 2934
rect 12582 2878 12650 2934
rect 12706 2878 12774 2934
rect 12830 2878 12898 2934
rect 12954 2878 13022 2934
rect 13078 2878 13200 2934
rect 12400 2810 13200 2878
rect 12400 2754 12526 2810
rect 12582 2754 12650 2810
rect 12706 2754 12774 2810
rect 12830 2754 12898 2810
rect 12954 2754 13022 2810
rect 13078 2754 13200 2810
rect 12400 2686 13200 2754
rect 12400 2630 12526 2686
rect 12582 2630 12650 2686
rect 12706 2630 12774 2686
rect 12830 2630 12898 2686
rect 12954 2630 13022 2686
rect 13078 2630 13200 2686
rect 12400 2562 13200 2630
rect 12400 2506 12526 2562
rect 12582 2506 12650 2562
rect 12706 2506 12774 2562
rect 12830 2506 12898 2562
rect 12954 2506 13022 2562
rect 13078 2506 13200 2562
rect 12400 2438 13200 2506
rect 12400 2382 12526 2438
rect 12582 2382 12650 2438
rect 12706 2382 12774 2438
rect 12830 2382 12898 2438
rect 12954 2382 13022 2438
rect 13078 2382 13200 2438
rect 12400 2314 13200 2382
rect 12400 2258 12526 2314
rect 12582 2258 12650 2314
rect 12706 2258 12774 2314
rect 12830 2258 12898 2314
rect 12954 2258 13022 2314
rect 13078 2258 13200 2314
rect 12400 2190 13200 2258
rect 12400 2134 12526 2190
rect 12582 2134 12650 2190
rect 12706 2134 12774 2190
rect 12830 2134 12898 2190
rect 12954 2134 13022 2190
rect 13078 2134 13200 2190
rect 12400 2066 13200 2134
rect 12400 2010 12526 2066
rect 12582 2010 12650 2066
rect 12706 2010 12774 2066
rect 12830 2010 12898 2066
rect 12954 2010 13022 2066
rect 13078 2010 13200 2066
rect 12400 1942 13200 2010
rect 12400 1886 12526 1942
rect 12582 1886 12650 1942
rect 12706 1886 12774 1942
rect 12830 1886 12898 1942
rect 12954 1886 13022 1942
rect 13078 1886 13200 1942
rect 12400 1818 13200 1886
rect 12400 1762 12526 1818
rect 12582 1762 12650 1818
rect 12706 1762 12774 1818
rect 12830 1762 12898 1818
rect 12954 1762 13022 1818
rect 13078 1762 13200 1818
rect 12400 1694 13200 1762
rect 12400 1638 12526 1694
rect 12582 1638 12650 1694
rect 12706 1638 12774 1694
rect 12830 1638 12898 1694
rect 12954 1638 13022 1694
rect 13078 1638 13200 1694
rect 12400 1570 13200 1638
rect 12400 1514 12526 1570
rect 12582 1514 12650 1570
rect 12706 1514 12774 1570
rect 12830 1514 12898 1570
rect 12954 1514 13022 1570
rect 13078 1514 13200 1570
rect 12400 1446 13200 1514
rect 12400 1390 12526 1446
rect 12582 1390 12650 1446
rect 12706 1390 12774 1446
rect 12830 1390 12898 1446
rect 12954 1390 13022 1446
rect 13078 1390 13200 1446
rect 12400 1322 13200 1390
rect 12400 1266 12526 1322
rect 12582 1266 12650 1322
rect 12706 1266 12774 1322
rect 12830 1266 12898 1322
rect 12954 1266 13022 1322
rect 13078 1266 13200 1322
rect 12400 1198 13200 1266
rect 12400 1142 12526 1198
rect 12582 1142 12650 1198
rect 12706 1142 12774 1198
rect 12830 1142 12898 1198
rect 12954 1142 13022 1198
rect 13078 1142 13200 1198
rect 12400 1074 13200 1142
rect 12400 1018 12526 1074
rect 12582 1018 12650 1074
rect 12706 1018 12774 1074
rect 12830 1018 12898 1074
rect 12954 1018 13022 1074
rect 13078 1018 13200 1074
rect 12400 950 13200 1018
rect 12400 894 12526 950
rect 12582 894 12650 950
rect 12706 894 12774 950
rect 12830 894 12898 950
rect 12954 894 13022 950
rect 13078 894 13200 950
rect 12400 826 13200 894
rect 12400 770 12526 826
rect 12582 770 12650 826
rect 12706 770 12774 826
rect 12830 770 12898 826
rect 12954 770 13022 826
rect 13078 770 13200 826
rect 12400 702 13200 770
rect 12400 646 12526 702
rect 12582 646 12650 702
rect 12706 646 12774 702
rect 12830 646 12898 702
rect 12954 646 13022 702
rect 13078 646 13200 702
rect 12400 578 13200 646
rect 12400 522 12526 578
rect 12582 522 12650 578
rect 12706 522 12774 578
rect 12830 522 12898 578
rect 12954 522 13022 578
rect 13078 522 13200 578
rect 12400 454 13200 522
rect 12400 400 12526 454
rect 266 398 12526 400
rect 12582 398 12650 454
rect 12706 398 12774 454
rect 12830 398 12898 454
rect 12954 398 13022 454
rect 13078 398 13200 454
rect -400 330 13200 398
rect -400 274 -286 330
rect -230 274 -162 330
rect -106 274 -38 330
rect 18 274 86 330
rect 142 274 210 330
rect 266 302 12526 330
rect 266 274 415 302
rect -400 246 415 274
rect 471 246 557 302
rect 613 246 699 302
rect 755 246 841 302
rect 897 246 983 302
rect 1039 246 1125 302
rect 1181 246 1267 302
rect 1323 246 1409 302
rect 1465 246 1551 302
rect 1607 246 1693 302
rect 1749 246 1835 302
rect 1891 246 1977 302
rect 2033 246 2119 302
rect 2175 246 2261 302
rect 2317 246 2403 302
rect 2459 246 2545 302
rect 2601 246 2687 302
rect 2743 246 2829 302
rect 2885 246 2971 302
rect 3027 246 3113 302
rect 3169 246 3255 302
rect 3311 246 3397 302
rect 3453 246 3539 302
rect 3595 246 3681 302
rect 3737 246 3823 302
rect 3879 246 3965 302
rect 4021 246 4107 302
rect 4163 246 4249 302
rect 4305 246 4391 302
rect 4447 246 4533 302
rect 4589 246 4675 302
rect 4731 246 4817 302
rect 4873 246 4959 302
rect 5015 246 5101 302
rect 5157 246 5243 302
rect 5299 246 5385 302
rect 5441 246 5527 302
rect 5583 246 5669 302
rect 5725 246 5811 302
rect 5867 246 5953 302
rect 6009 246 6095 302
rect 6151 246 6237 302
rect 6293 246 6379 302
rect 6435 246 6521 302
rect 6577 246 6663 302
rect 6719 246 6805 302
rect 6861 246 6947 302
rect 7003 246 7089 302
rect 7145 246 7231 302
rect 7287 246 7373 302
rect 7429 246 7515 302
rect 7571 246 7657 302
rect 7713 246 7799 302
rect 7855 246 7941 302
rect 7997 246 8083 302
rect 8139 246 8225 302
rect 8281 246 8367 302
rect 8423 246 8509 302
rect 8565 246 8651 302
rect 8707 246 8793 302
rect 8849 246 8935 302
rect 8991 246 9077 302
rect 9133 246 9219 302
rect 9275 246 9361 302
rect 9417 246 9503 302
rect 9559 246 9645 302
rect 9701 246 9787 302
rect 9843 246 9929 302
rect 9985 246 10071 302
rect 10127 246 10213 302
rect 10269 246 10355 302
rect 10411 246 10497 302
rect 10553 246 10639 302
rect 10695 246 10781 302
rect 10837 246 10923 302
rect 10979 246 11065 302
rect 11121 246 11207 302
rect 11263 246 11349 302
rect 11405 246 11491 302
rect 11547 246 11633 302
rect 11689 246 11775 302
rect 11831 246 11917 302
rect 11973 246 12059 302
rect 12115 246 12201 302
rect 12257 246 12343 302
rect 12399 274 12526 302
rect 12582 274 12650 330
rect 12706 274 12774 330
rect 12830 274 12898 330
rect 12954 274 13022 330
rect 13078 274 13200 330
rect 12399 246 13200 274
rect -400 206 13200 246
rect -400 150 -286 206
rect -230 150 -162 206
rect -106 150 -38 206
rect 18 150 86 206
rect 142 150 210 206
rect 266 160 12526 206
rect 266 150 415 160
rect -400 104 415 150
rect 471 104 557 160
rect 613 104 699 160
rect 755 104 841 160
rect 897 104 983 160
rect 1039 104 1125 160
rect 1181 104 1267 160
rect 1323 104 1409 160
rect 1465 104 1551 160
rect 1607 104 1693 160
rect 1749 104 1835 160
rect 1891 104 1977 160
rect 2033 104 2119 160
rect 2175 104 2261 160
rect 2317 104 2403 160
rect 2459 104 2545 160
rect 2601 104 2687 160
rect 2743 104 2829 160
rect 2885 104 2971 160
rect 3027 104 3113 160
rect 3169 104 3255 160
rect 3311 104 3397 160
rect 3453 104 3539 160
rect 3595 104 3681 160
rect 3737 104 3823 160
rect 3879 104 3965 160
rect 4021 104 4107 160
rect 4163 104 4249 160
rect 4305 104 4391 160
rect 4447 104 4533 160
rect 4589 104 4675 160
rect 4731 104 4817 160
rect 4873 104 4959 160
rect 5015 104 5101 160
rect 5157 104 5243 160
rect 5299 104 5385 160
rect 5441 104 5527 160
rect 5583 104 5669 160
rect 5725 104 5811 160
rect 5867 104 5953 160
rect 6009 104 6095 160
rect 6151 104 6237 160
rect 6293 104 6379 160
rect 6435 104 6521 160
rect 6577 104 6663 160
rect 6719 104 6805 160
rect 6861 104 6947 160
rect 7003 104 7089 160
rect 7145 104 7231 160
rect 7287 104 7373 160
rect 7429 104 7515 160
rect 7571 104 7657 160
rect 7713 104 7799 160
rect 7855 104 7941 160
rect 7997 104 8083 160
rect 8139 104 8225 160
rect 8281 104 8367 160
rect 8423 104 8509 160
rect 8565 104 8651 160
rect 8707 104 8793 160
rect 8849 104 8935 160
rect 8991 104 9077 160
rect 9133 104 9219 160
rect 9275 104 9361 160
rect 9417 104 9503 160
rect 9559 104 9645 160
rect 9701 104 9787 160
rect 9843 104 9929 160
rect 9985 104 10071 160
rect 10127 104 10213 160
rect 10269 104 10355 160
rect 10411 104 10497 160
rect 10553 104 10639 160
rect 10695 104 10781 160
rect 10837 104 10923 160
rect 10979 104 11065 160
rect 11121 104 11207 160
rect 11263 104 11349 160
rect 11405 104 11491 160
rect 11547 104 11633 160
rect 11689 104 11775 160
rect 11831 104 11917 160
rect 11973 104 12059 160
rect 12115 104 12201 160
rect 12257 104 12343 160
rect 12399 150 12526 160
rect 12582 150 12650 206
rect 12706 150 12774 206
rect 12830 150 12898 206
rect 12954 150 13022 206
rect 13078 150 13200 206
rect 12399 104 13200 150
rect -400 0 13200 104
<< via3 >>
rect -254 12893 -198 12949
rect -130 12893 -74 12949
rect -6 12893 50 12949
rect 118 12893 174 12949
rect 242 12893 298 12949
rect 366 12893 422 12949
rect 490 12893 546 12949
rect 614 12893 670 12949
rect 738 12893 794 12949
rect 862 12893 918 12949
rect 986 12893 1042 12949
rect 1110 12893 1166 12949
rect 1234 12893 1290 12949
rect 1358 12893 1414 12949
rect 1482 12893 1538 12949
rect 1606 12893 1662 12949
rect 1730 12893 1786 12949
rect 1854 12893 1910 12949
rect 1978 12893 2034 12949
rect 2102 12893 2158 12949
rect 2226 12893 2282 12949
rect 2350 12893 2406 12949
rect 2474 12893 2530 12949
rect 2598 12893 2654 12949
rect 2722 12893 2778 12949
rect 2846 12893 2902 12949
rect 2970 12893 3026 12949
rect 3094 12893 3150 12949
rect 3218 12893 3274 12949
rect 3342 12893 3398 12949
rect 3466 12893 3522 12949
rect 3590 12893 3646 12949
rect 3714 12893 3770 12949
rect 3838 12893 3894 12949
rect 3962 12893 4018 12949
rect 4086 12893 4142 12949
rect 4210 12893 4266 12949
rect 4334 12893 4390 12949
rect 4458 12893 4514 12949
rect 4582 12893 4638 12949
rect 4706 12893 4762 12949
rect 4830 12893 4886 12949
rect 4954 12893 5010 12949
rect 5078 12893 5134 12949
rect 5202 12893 5258 12949
rect 5326 12893 5382 12949
rect 5450 12893 5506 12949
rect 5574 12893 5630 12949
rect 5698 12893 5754 12949
rect 5822 12893 5878 12949
rect 5946 12893 6002 12949
rect 6070 12893 6126 12949
rect 6194 12893 6250 12949
rect 6318 12893 6374 12949
rect 6442 12893 6498 12949
rect 6566 12893 6622 12949
rect 6690 12893 6746 12949
rect 6814 12893 6870 12949
rect 6938 12893 6994 12949
rect 7062 12893 7118 12949
rect 7186 12893 7242 12949
rect 7310 12893 7366 12949
rect 7434 12893 7490 12949
rect 7558 12893 7614 12949
rect 7682 12893 7738 12949
rect 7806 12893 7862 12949
rect 7930 12893 7986 12949
rect 8054 12893 8110 12949
rect 8178 12893 8234 12949
rect 8302 12893 8358 12949
rect 8426 12893 8482 12949
rect 8550 12893 8606 12949
rect 8674 12893 8730 12949
rect 8798 12893 8854 12949
rect 8922 12893 8978 12949
rect 9046 12893 9102 12949
rect 9170 12893 9226 12949
rect 9294 12893 9350 12949
rect 9418 12893 9474 12949
rect 9542 12893 9598 12949
rect 9666 12893 9722 12949
rect 9790 12893 9846 12949
rect 9914 12893 9970 12949
rect 10038 12893 10094 12949
rect 10162 12893 10218 12949
rect 10286 12893 10342 12949
rect 10410 12893 10466 12949
rect 10534 12893 10590 12949
rect 10658 12893 10714 12949
rect 10782 12893 10838 12949
rect 10906 12893 10962 12949
rect 11030 12893 11086 12949
rect 11154 12893 11210 12949
rect 11278 12893 11334 12949
rect 11402 12893 11458 12949
rect 11526 12893 11582 12949
rect 11650 12893 11706 12949
rect 11774 12893 11830 12949
rect 11898 12893 11954 12949
rect 12022 12893 12078 12949
rect 12146 12893 12202 12949
rect 12270 12893 12326 12949
rect 12394 12893 12450 12949
rect 12518 12893 12574 12949
rect 12642 12893 12698 12949
rect 12766 12893 12822 12949
rect 12890 12893 12946 12949
rect 13014 12893 13070 12949
rect -254 12769 -198 12825
rect -130 12769 -74 12825
rect -6 12769 50 12825
rect 118 12769 174 12825
rect 242 12769 298 12825
rect 366 12769 422 12825
rect 490 12769 546 12825
rect 614 12769 670 12825
rect 738 12769 794 12825
rect 862 12769 918 12825
rect 986 12769 1042 12825
rect 1110 12769 1166 12825
rect 1234 12769 1290 12825
rect 1358 12769 1414 12825
rect 1482 12769 1538 12825
rect 1606 12769 1662 12825
rect 1730 12769 1786 12825
rect 1854 12769 1910 12825
rect 1978 12769 2034 12825
rect 2102 12769 2158 12825
rect 2226 12769 2282 12825
rect 2350 12769 2406 12825
rect 2474 12769 2530 12825
rect 2598 12769 2654 12825
rect 2722 12769 2778 12825
rect 2846 12769 2902 12825
rect 2970 12769 3026 12825
rect 3094 12769 3150 12825
rect 3218 12769 3274 12825
rect 3342 12769 3398 12825
rect 3466 12769 3522 12825
rect 3590 12769 3646 12825
rect 3714 12769 3770 12825
rect 3838 12769 3894 12825
rect 3962 12769 4018 12825
rect 4086 12769 4142 12825
rect 4210 12769 4266 12825
rect 4334 12769 4390 12825
rect 4458 12769 4514 12825
rect 4582 12769 4638 12825
rect 4706 12769 4762 12825
rect 4830 12769 4886 12825
rect 4954 12769 5010 12825
rect 5078 12769 5134 12825
rect 5202 12769 5258 12825
rect 5326 12769 5382 12825
rect 5450 12769 5506 12825
rect 5574 12769 5630 12825
rect 5698 12769 5754 12825
rect 5822 12769 5878 12825
rect 5946 12769 6002 12825
rect 6070 12769 6126 12825
rect 6194 12769 6250 12825
rect 6318 12769 6374 12825
rect 6442 12769 6498 12825
rect 6566 12769 6622 12825
rect 6690 12769 6746 12825
rect 6814 12769 6870 12825
rect 6938 12769 6994 12825
rect 7062 12769 7118 12825
rect 7186 12769 7242 12825
rect 7310 12769 7366 12825
rect 7434 12769 7490 12825
rect 7558 12769 7614 12825
rect 7682 12769 7738 12825
rect 7806 12769 7862 12825
rect 7930 12769 7986 12825
rect 8054 12769 8110 12825
rect 8178 12769 8234 12825
rect 8302 12769 8358 12825
rect 8426 12769 8482 12825
rect 8550 12769 8606 12825
rect 8674 12769 8730 12825
rect 8798 12769 8854 12825
rect 8922 12769 8978 12825
rect 9046 12769 9102 12825
rect 9170 12769 9226 12825
rect 9294 12769 9350 12825
rect 9418 12769 9474 12825
rect 9542 12769 9598 12825
rect 9666 12769 9722 12825
rect 9790 12769 9846 12825
rect 9914 12769 9970 12825
rect 10038 12769 10094 12825
rect 10162 12769 10218 12825
rect 10286 12769 10342 12825
rect 10410 12769 10466 12825
rect 10534 12769 10590 12825
rect 10658 12769 10714 12825
rect 10782 12769 10838 12825
rect 10906 12769 10962 12825
rect 11030 12769 11086 12825
rect 11154 12769 11210 12825
rect 11278 12769 11334 12825
rect 11402 12769 11458 12825
rect 11526 12769 11582 12825
rect 11650 12769 11706 12825
rect 11774 12769 11830 12825
rect 11898 12769 11954 12825
rect 12022 12769 12078 12825
rect 12146 12769 12202 12825
rect 12270 12769 12326 12825
rect 12394 12769 12450 12825
rect 12518 12769 12574 12825
rect 12642 12769 12698 12825
rect 12766 12769 12822 12825
rect 12890 12769 12946 12825
rect 13014 12769 13070 12825
rect -254 12645 -198 12701
rect -130 12645 -74 12701
rect -6 12645 50 12701
rect 118 12645 174 12701
rect 242 12645 298 12701
rect 366 12645 422 12701
rect 490 12645 546 12701
rect 614 12645 670 12701
rect 738 12645 794 12701
rect 862 12645 918 12701
rect 986 12645 1042 12701
rect 1110 12645 1166 12701
rect 1234 12645 1290 12701
rect 1358 12645 1414 12701
rect 1482 12645 1538 12701
rect 1606 12645 1662 12701
rect 1730 12645 1786 12701
rect 1854 12645 1910 12701
rect 1978 12645 2034 12701
rect 2102 12645 2158 12701
rect 2226 12645 2282 12701
rect 2350 12645 2406 12701
rect 2474 12645 2530 12701
rect 2598 12645 2654 12701
rect 2722 12645 2778 12701
rect 2846 12645 2902 12701
rect 2970 12645 3026 12701
rect 3094 12645 3150 12701
rect 3218 12645 3274 12701
rect 3342 12645 3398 12701
rect 3466 12645 3522 12701
rect 3590 12645 3646 12701
rect 3714 12645 3770 12701
rect 3838 12645 3894 12701
rect 3962 12645 4018 12701
rect 4086 12645 4142 12701
rect 4210 12645 4266 12701
rect 4334 12645 4390 12701
rect 4458 12645 4514 12701
rect 4582 12645 4638 12701
rect 4706 12645 4762 12701
rect 4830 12645 4886 12701
rect 4954 12645 5010 12701
rect 5078 12645 5134 12701
rect 5202 12645 5258 12701
rect 5326 12645 5382 12701
rect 5450 12645 5506 12701
rect 5574 12645 5630 12701
rect 5698 12645 5754 12701
rect 5822 12645 5878 12701
rect 5946 12645 6002 12701
rect 6070 12645 6126 12701
rect 6194 12645 6250 12701
rect 6318 12645 6374 12701
rect 6442 12645 6498 12701
rect 6566 12645 6622 12701
rect 6690 12645 6746 12701
rect 6814 12645 6870 12701
rect 6938 12645 6994 12701
rect 7062 12645 7118 12701
rect 7186 12645 7242 12701
rect 7310 12645 7366 12701
rect 7434 12645 7490 12701
rect 7558 12645 7614 12701
rect 7682 12645 7738 12701
rect 7806 12645 7862 12701
rect 7930 12645 7986 12701
rect 8054 12645 8110 12701
rect 8178 12645 8234 12701
rect 8302 12645 8358 12701
rect 8426 12645 8482 12701
rect 8550 12645 8606 12701
rect 8674 12645 8730 12701
rect 8798 12645 8854 12701
rect 8922 12645 8978 12701
rect 9046 12645 9102 12701
rect 9170 12645 9226 12701
rect 9294 12645 9350 12701
rect 9418 12645 9474 12701
rect 9542 12645 9598 12701
rect 9666 12645 9722 12701
rect 9790 12645 9846 12701
rect 9914 12645 9970 12701
rect 10038 12645 10094 12701
rect 10162 12645 10218 12701
rect 10286 12645 10342 12701
rect 10410 12645 10466 12701
rect 10534 12645 10590 12701
rect 10658 12645 10714 12701
rect 10782 12645 10838 12701
rect 10906 12645 10962 12701
rect 11030 12645 11086 12701
rect 11154 12645 11210 12701
rect 11278 12645 11334 12701
rect 11402 12645 11458 12701
rect 11526 12645 11582 12701
rect 11650 12645 11706 12701
rect 11774 12645 11830 12701
rect 11898 12645 11954 12701
rect 12022 12645 12078 12701
rect 12146 12645 12202 12701
rect 12270 12645 12326 12701
rect 12394 12645 12450 12701
rect 12518 12645 12574 12701
rect 12642 12645 12698 12701
rect 12766 12645 12822 12701
rect 12890 12645 12946 12701
rect 13014 12645 13070 12701
rect -254 12521 -198 12577
rect -130 12521 -74 12577
rect -6 12521 50 12577
rect 118 12521 174 12577
rect 242 12521 298 12577
rect 366 12521 422 12577
rect 490 12521 546 12577
rect 614 12521 670 12577
rect 738 12521 794 12577
rect 862 12521 918 12577
rect 986 12521 1042 12577
rect 1110 12521 1166 12577
rect 1234 12521 1290 12577
rect 1358 12521 1414 12577
rect 1482 12521 1538 12577
rect 1606 12521 1662 12577
rect 1730 12521 1786 12577
rect 1854 12521 1910 12577
rect 1978 12521 2034 12577
rect 2102 12521 2158 12577
rect 2226 12521 2282 12577
rect 2350 12521 2406 12577
rect 2474 12521 2530 12577
rect 2598 12521 2654 12577
rect 2722 12521 2778 12577
rect 2846 12521 2902 12577
rect 2970 12521 3026 12577
rect 3094 12521 3150 12577
rect 3218 12521 3274 12577
rect 3342 12521 3398 12577
rect 3466 12521 3522 12577
rect 3590 12521 3646 12577
rect 3714 12521 3770 12577
rect 3838 12521 3894 12577
rect 3962 12521 4018 12577
rect 4086 12521 4142 12577
rect 4210 12521 4266 12577
rect 4334 12521 4390 12577
rect 4458 12521 4514 12577
rect 4582 12521 4638 12577
rect 4706 12521 4762 12577
rect 4830 12521 4886 12577
rect 4954 12521 5010 12577
rect 5078 12521 5134 12577
rect 5202 12521 5258 12577
rect 5326 12521 5382 12577
rect 5450 12521 5506 12577
rect 5574 12521 5630 12577
rect 5698 12521 5754 12577
rect 5822 12521 5878 12577
rect 5946 12521 6002 12577
rect 6070 12521 6126 12577
rect 6194 12521 6250 12577
rect 6318 12521 6374 12577
rect 6442 12521 6498 12577
rect 6566 12521 6622 12577
rect 6690 12521 6746 12577
rect 6814 12521 6870 12577
rect 6938 12521 6994 12577
rect 7062 12521 7118 12577
rect 7186 12521 7242 12577
rect 7310 12521 7366 12577
rect 7434 12521 7490 12577
rect 7558 12521 7614 12577
rect 7682 12521 7738 12577
rect 7806 12521 7862 12577
rect 7930 12521 7986 12577
rect 8054 12521 8110 12577
rect 8178 12521 8234 12577
rect 8302 12521 8358 12577
rect 8426 12521 8482 12577
rect 8550 12521 8606 12577
rect 8674 12521 8730 12577
rect 8798 12521 8854 12577
rect 8922 12521 8978 12577
rect 9046 12521 9102 12577
rect 9170 12521 9226 12577
rect 9294 12521 9350 12577
rect 9418 12521 9474 12577
rect 9542 12521 9598 12577
rect 9666 12521 9722 12577
rect 9790 12521 9846 12577
rect 9914 12521 9970 12577
rect 10038 12521 10094 12577
rect 10162 12521 10218 12577
rect 10286 12521 10342 12577
rect 10410 12521 10466 12577
rect 10534 12521 10590 12577
rect 10658 12521 10714 12577
rect 10782 12521 10838 12577
rect 10906 12521 10962 12577
rect 11030 12521 11086 12577
rect 11154 12521 11210 12577
rect 11278 12521 11334 12577
rect 11402 12521 11458 12577
rect 11526 12521 11582 12577
rect 11650 12521 11706 12577
rect 11774 12521 11830 12577
rect 11898 12521 11954 12577
rect 12022 12521 12078 12577
rect 12146 12521 12202 12577
rect 12270 12521 12326 12577
rect 12394 12521 12450 12577
rect 12518 12521 12574 12577
rect 12642 12521 12698 12577
rect 12766 12521 12822 12577
rect 12890 12521 12946 12577
rect 13014 12521 13070 12577
rect -286 12302 -230 12358
rect -162 12302 -106 12358
rect -38 12302 18 12358
rect 86 12302 142 12358
rect 210 12302 266 12358
rect -286 12178 -230 12234
rect -162 12178 -106 12234
rect -38 12178 18 12234
rect 86 12178 142 12234
rect 210 12178 266 12234
rect -286 12054 -230 12110
rect -162 12054 -106 12110
rect -38 12054 18 12110
rect 86 12054 142 12110
rect 210 12054 266 12110
rect -286 11930 -230 11986
rect -162 11930 -106 11986
rect -38 11930 18 11986
rect 86 11930 142 11986
rect 210 11930 266 11986
rect -286 11806 -230 11862
rect -162 11806 -106 11862
rect -38 11806 18 11862
rect 86 11806 142 11862
rect 210 11806 266 11862
rect -286 11682 -230 11738
rect -162 11682 -106 11738
rect -38 11682 18 11738
rect 86 11682 142 11738
rect 210 11682 266 11738
rect -286 11558 -230 11614
rect -162 11558 -106 11614
rect -38 11558 18 11614
rect 86 11558 142 11614
rect 210 11558 266 11614
rect -286 11434 -230 11490
rect -162 11434 -106 11490
rect -38 11434 18 11490
rect 86 11434 142 11490
rect 210 11434 266 11490
rect -286 11310 -230 11366
rect -162 11310 -106 11366
rect -38 11310 18 11366
rect 86 11310 142 11366
rect 210 11310 266 11366
rect -286 11186 -230 11242
rect -162 11186 -106 11242
rect -38 11186 18 11242
rect 86 11186 142 11242
rect 210 11186 266 11242
rect -286 11062 -230 11118
rect -162 11062 -106 11118
rect -38 11062 18 11118
rect 86 11062 142 11118
rect 210 11062 266 11118
rect -286 10938 -230 10994
rect -162 10938 -106 10994
rect -38 10938 18 10994
rect 86 10938 142 10994
rect 210 10938 266 10994
rect -286 10814 -230 10870
rect -162 10814 -106 10870
rect -38 10814 18 10870
rect 86 10814 142 10870
rect 210 10814 266 10870
rect -286 10690 -230 10746
rect -162 10690 -106 10746
rect -38 10690 18 10746
rect 86 10690 142 10746
rect 210 10690 266 10746
rect -286 10566 -230 10622
rect -162 10566 -106 10622
rect -38 10566 18 10622
rect 86 10566 142 10622
rect 210 10566 266 10622
rect -286 10442 -230 10498
rect -162 10442 -106 10498
rect -38 10442 18 10498
rect 86 10442 142 10498
rect 210 10442 266 10498
rect -286 10318 -230 10374
rect -162 10318 -106 10374
rect -38 10318 18 10374
rect 86 10318 142 10374
rect 210 10318 266 10374
rect -286 10194 -230 10250
rect -162 10194 -106 10250
rect -38 10194 18 10250
rect 86 10194 142 10250
rect 210 10194 266 10250
rect -286 10070 -230 10126
rect -162 10070 -106 10126
rect -38 10070 18 10126
rect 86 10070 142 10126
rect 210 10070 266 10126
rect -286 9946 -230 10002
rect -162 9946 -106 10002
rect -38 9946 18 10002
rect 86 9946 142 10002
rect 210 9946 266 10002
rect -286 9822 -230 9878
rect -162 9822 -106 9878
rect -38 9822 18 9878
rect 86 9822 142 9878
rect 210 9822 266 9878
rect -286 9698 -230 9754
rect -162 9698 -106 9754
rect -38 9698 18 9754
rect 86 9698 142 9754
rect 210 9698 266 9754
rect -286 9574 -230 9630
rect -162 9574 -106 9630
rect -38 9574 18 9630
rect 86 9574 142 9630
rect 210 9574 266 9630
rect -286 9450 -230 9506
rect -162 9450 -106 9506
rect -38 9450 18 9506
rect 86 9450 142 9506
rect 210 9450 266 9506
rect -286 9326 -230 9382
rect -162 9326 -106 9382
rect -38 9326 18 9382
rect 86 9326 142 9382
rect 210 9326 266 9382
rect -286 9202 -230 9258
rect -162 9202 -106 9258
rect -38 9202 18 9258
rect 86 9202 142 9258
rect 210 9202 266 9258
rect -286 9078 -230 9134
rect -162 9078 -106 9134
rect -38 9078 18 9134
rect 86 9078 142 9134
rect 210 9078 266 9134
rect -286 8954 -230 9010
rect -162 8954 -106 9010
rect -38 8954 18 9010
rect 86 8954 142 9010
rect 210 8954 266 9010
rect -286 8830 -230 8886
rect -162 8830 -106 8886
rect -38 8830 18 8886
rect 86 8830 142 8886
rect 210 8830 266 8886
rect -286 8706 -230 8762
rect -162 8706 -106 8762
rect -38 8706 18 8762
rect 86 8706 142 8762
rect 210 8706 266 8762
rect -286 8582 -230 8638
rect -162 8582 -106 8638
rect -38 8582 18 8638
rect 86 8582 142 8638
rect 210 8582 266 8638
rect -286 8458 -230 8514
rect -162 8458 -106 8514
rect -38 8458 18 8514
rect 86 8458 142 8514
rect 210 8458 266 8514
rect -286 8334 -230 8390
rect -162 8334 -106 8390
rect -38 8334 18 8390
rect 86 8334 142 8390
rect 210 8334 266 8390
rect -286 8210 -230 8266
rect -162 8210 -106 8266
rect -38 8210 18 8266
rect 86 8210 142 8266
rect 210 8210 266 8266
rect -286 8086 -230 8142
rect -162 8086 -106 8142
rect -38 8086 18 8142
rect 86 8086 142 8142
rect 210 8086 266 8142
rect -286 7962 -230 8018
rect -162 7962 -106 8018
rect -38 7962 18 8018
rect 86 7962 142 8018
rect 210 7962 266 8018
rect -286 7838 -230 7894
rect -162 7838 -106 7894
rect -38 7838 18 7894
rect 86 7838 142 7894
rect 210 7838 266 7894
rect -286 7714 -230 7770
rect -162 7714 -106 7770
rect -38 7714 18 7770
rect 86 7714 142 7770
rect 210 7714 266 7770
rect -286 7590 -230 7646
rect -162 7590 -106 7646
rect -38 7590 18 7646
rect 86 7590 142 7646
rect 210 7590 266 7646
rect -286 7466 -230 7522
rect -162 7466 -106 7522
rect -38 7466 18 7522
rect 86 7466 142 7522
rect 210 7466 266 7522
rect -286 7342 -230 7398
rect -162 7342 -106 7398
rect -38 7342 18 7398
rect 86 7342 142 7398
rect 210 7342 266 7398
rect -286 7218 -230 7274
rect -162 7218 -106 7274
rect -38 7218 18 7274
rect 86 7218 142 7274
rect 210 7218 266 7274
rect -286 7094 -230 7150
rect -162 7094 -106 7150
rect -38 7094 18 7150
rect 86 7094 142 7150
rect 210 7094 266 7150
rect -286 6970 -230 7026
rect -162 6970 -106 7026
rect -38 6970 18 7026
rect 86 6970 142 7026
rect 210 6970 266 7026
rect -286 6846 -230 6902
rect -162 6846 -106 6902
rect -38 6846 18 6902
rect 86 6846 142 6902
rect 210 6846 266 6902
rect -286 6722 -230 6778
rect -162 6722 -106 6778
rect -38 6722 18 6778
rect 86 6722 142 6778
rect 210 6722 266 6778
rect -286 6598 -230 6654
rect -162 6598 -106 6654
rect -38 6598 18 6654
rect 86 6598 142 6654
rect 210 6598 266 6654
rect -286 6474 -230 6530
rect -162 6474 -106 6530
rect -38 6474 18 6530
rect 86 6474 142 6530
rect 210 6474 266 6530
rect -286 6350 -230 6406
rect -162 6350 -106 6406
rect -38 6350 18 6406
rect 86 6350 142 6406
rect 210 6350 266 6406
rect -286 6226 -230 6282
rect -162 6226 -106 6282
rect -38 6226 18 6282
rect 86 6226 142 6282
rect 210 6226 266 6282
rect -286 6102 -230 6158
rect -162 6102 -106 6158
rect -38 6102 18 6158
rect 86 6102 142 6158
rect 210 6102 266 6158
rect -286 5978 -230 6034
rect -162 5978 -106 6034
rect -38 5978 18 6034
rect 86 5978 142 6034
rect 210 5978 266 6034
rect -286 5854 -230 5910
rect -162 5854 -106 5910
rect -38 5854 18 5910
rect 86 5854 142 5910
rect 210 5854 266 5910
rect -286 5730 -230 5786
rect -162 5730 -106 5786
rect -38 5730 18 5786
rect 86 5730 142 5786
rect 210 5730 266 5786
rect -286 5606 -230 5662
rect -162 5606 -106 5662
rect -38 5606 18 5662
rect 86 5606 142 5662
rect 210 5606 266 5662
rect -286 5482 -230 5538
rect -162 5482 -106 5538
rect -38 5482 18 5538
rect 86 5482 142 5538
rect 210 5482 266 5538
rect -286 5358 -230 5414
rect -162 5358 -106 5414
rect -38 5358 18 5414
rect 86 5358 142 5414
rect 210 5358 266 5414
rect -286 5234 -230 5290
rect -162 5234 -106 5290
rect -38 5234 18 5290
rect 86 5234 142 5290
rect 210 5234 266 5290
rect -286 5110 -230 5166
rect -162 5110 -106 5166
rect -38 5110 18 5166
rect 86 5110 142 5166
rect 210 5110 266 5166
rect -286 4986 -230 5042
rect -162 4986 -106 5042
rect -38 4986 18 5042
rect 86 4986 142 5042
rect 210 4986 266 5042
rect -286 4862 -230 4918
rect -162 4862 -106 4918
rect -38 4862 18 4918
rect 86 4862 142 4918
rect 210 4862 266 4918
rect -286 4738 -230 4794
rect -162 4738 -106 4794
rect -38 4738 18 4794
rect 86 4738 142 4794
rect 210 4738 266 4794
rect -286 4614 -230 4670
rect -162 4614 -106 4670
rect -38 4614 18 4670
rect 86 4614 142 4670
rect 210 4614 266 4670
rect -286 4490 -230 4546
rect -162 4490 -106 4546
rect -38 4490 18 4546
rect 86 4490 142 4546
rect 210 4490 266 4546
rect -286 4366 -230 4422
rect -162 4366 -106 4422
rect -38 4366 18 4422
rect 86 4366 142 4422
rect 210 4366 266 4422
rect -286 4242 -230 4298
rect -162 4242 -106 4298
rect -38 4242 18 4298
rect 86 4242 142 4298
rect 210 4242 266 4298
rect -286 4118 -230 4174
rect -162 4118 -106 4174
rect -38 4118 18 4174
rect 86 4118 142 4174
rect 210 4118 266 4174
rect -286 3994 -230 4050
rect -162 3994 -106 4050
rect -38 3994 18 4050
rect 86 3994 142 4050
rect 210 3994 266 4050
rect -286 3870 -230 3926
rect -162 3870 -106 3926
rect -38 3870 18 3926
rect 86 3870 142 3926
rect 210 3870 266 3926
rect -286 3746 -230 3802
rect -162 3746 -106 3802
rect -38 3746 18 3802
rect 86 3746 142 3802
rect 210 3746 266 3802
rect -286 3622 -230 3678
rect -162 3622 -106 3678
rect -38 3622 18 3678
rect 86 3622 142 3678
rect 210 3622 266 3678
rect -286 3498 -230 3554
rect -162 3498 -106 3554
rect -38 3498 18 3554
rect 86 3498 142 3554
rect 210 3498 266 3554
rect -286 3374 -230 3430
rect -162 3374 -106 3430
rect -38 3374 18 3430
rect 86 3374 142 3430
rect 210 3374 266 3430
rect -286 3250 -230 3306
rect -162 3250 -106 3306
rect -38 3250 18 3306
rect 86 3250 142 3306
rect 210 3250 266 3306
rect -286 3126 -230 3182
rect -162 3126 -106 3182
rect -38 3126 18 3182
rect 86 3126 142 3182
rect 210 3126 266 3182
rect -286 3002 -230 3058
rect -162 3002 -106 3058
rect -38 3002 18 3058
rect 86 3002 142 3058
rect 210 3002 266 3058
rect -286 2878 -230 2934
rect -162 2878 -106 2934
rect -38 2878 18 2934
rect 86 2878 142 2934
rect 210 2878 266 2934
rect -286 2754 -230 2810
rect -162 2754 -106 2810
rect -38 2754 18 2810
rect 86 2754 142 2810
rect 210 2754 266 2810
rect -286 2630 -230 2686
rect -162 2630 -106 2686
rect -38 2630 18 2686
rect 86 2630 142 2686
rect 210 2630 266 2686
rect -286 2506 -230 2562
rect -162 2506 -106 2562
rect -38 2506 18 2562
rect 86 2506 142 2562
rect 210 2506 266 2562
rect -286 2382 -230 2438
rect -162 2382 -106 2438
rect -38 2382 18 2438
rect 86 2382 142 2438
rect 210 2382 266 2438
rect -286 2258 -230 2314
rect -162 2258 -106 2314
rect -38 2258 18 2314
rect 86 2258 142 2314
rect 210 2258 266 2314
rect -286 2134 -230 2190
rect -162 2134 -106 2190
rect -38 2134 18 2190
rect 86 2134 142 2190
rect 210 2134 266 2190
rect -286 2010 -230 2066
rect -162 2010 -106 2066
rect -38 2010 18 2066
rect 86 2010 142 2066
rect 210 2010 266 2066
rect -286 1886 -230 1942
rect -162 1886 -106 1942
rect -38 1886 18 1942
rect 86 1886 142 1942
rect 210 1886 266 1942
rect -286 1762 -230 1818
rect -162 1762 -106 1818
rect -38 1762 18 1818
rect 86 1762 142 1818
rect 210 1762 266 1818
rect -286 1638 -230 1694
rect -162 1638 -106 1694
rect -38 1638 18 1694
rect 86 1638 142 1694
rect 210 1638 266 1694
rect -286 1514 -230 1570
rect -162 1514 -106 1570
rect -38 1514 18 1570
rect 86 1514 142 1570
rect 210 1514 266 1570
rect -286 1390 -230 1446
rect -162 1390 -106 1446
rect -38 1390 18 1446
rect 86 1390 142 1446
rect 210 1390 266 1446
rect -286 1266 -230 1322
rect -162 1266 -106 1322
rect -38 1266 18 1322
rect 86 1266 142 1322
rect 210 1266 266 1322
rect -286 1142 -230 1198
rect -162 1142 -106 1198
rect -38 1142 18 1198
rect 86 1142 142 1198
rect 210 1142 266 1198
rect -286 1018 -230 1074
rect -162 1018 -106 1074
rect -38 1018 18 1074
rect 86 1018 142 1074
rect 210 1018 266 1074
rect -286 894 -230 950
rect -162 894 -106 950
rect -38 894 18 950
rect 86 894 142 950
rect 210 894 266 950
rect -286 770 -230 826
rect -162 770 -106 826
rect -38 770 18 826
rect 86 770 142 826
rect 210 770 266 826
rect -286 646 -230 702
rect -162 646 -106 702
rect -38 646 18 702
rect 86 646 142 702
rect 210 646 266 702
rect -286 522 -230 578
rect -162 522 -106 578
rect -38 522 18 578
rect 86 522 142 578
rect 210 522 266 578
rect -286 398 -230 454
rect -162 398 -106 454
rect -38 398 18 454
rect 86 398 142 454
rect 210 398 266 454
rect 741 12254 797 12310
rect 883 12254 939 12310
rect 741 12112 797 12168
rect 883 12112 939 12168
rect 741 11970 797 12026
rect 883 11970 939 12026
rect 741 11828 797 11884
rect 883 11828 939 11884
rect 741 11686 797 11742
rect 883 11686 939 11742
rect 741 11544 797 11600
rect 883 11544 939 11600
rect 741 11402 797 11458
rect 883 11402 939 11458
rect 741 11260 797 11316
rect 883 11260 939 11316
rect 741 11118 797 11174
rect 883 11118 939 11174
rect 741 10976 797 11032
rect 883 10976 939 11032
rect 741 10834 797 10890
rect 883 10834 939 10890
rect 741 10692 797 10748
rect 883 10692 939 10748
rect 741 10550 797 10606
rect 883 10550 939 10606
rect 741 10408 797 10464
rect 883 10408 939 10464
rect 741 10266 797 10322
rect 883 10266 939 10322
rect 741 10124 797 10180
rect 883 10124 939 10180
rect 741 9982 797 10038
rect 883 9982 939 10038
rect 741 9840 797 9896
rect 883 9840 939 9896
rect 741 9698 797 9754
rect 883 9698 939 9754
rect 741 9556 797 9612
rect 883 9556 939 9612
rect 741 9414 797 9470
rect 883 9414 939 9470
rect 741 9272 797 9328
rect 883 9272 939 9328
rect 741 9130 797 9186
rect 883 9130 939 9186
rect 741 8988 797 9044
rect 883 8988 939 9044
rect 741 8846 797 8902
rect 883 8846 939 8902
rect 741 8704 797 8760
rect 883 8704 939 8760
rect 741 8562 797 8618
rect 883 8562 939 8618
rect 741 8420 797 8476
rect 883 8420 939 8476
rect 741 8278 797 8334
rect 883 8278 939 8334
rect 741 8136 797 8192
rect 883 8136 939 8192
rect 741 7994 797 8050
rect 883 7994 939 8050
rect 741 7852 797 7908
rect 883 7852 939 7908
rect 741 7710 797 7766
rect 883 7710 939 7766
rect 741 7568 797 7624
rect 883 7568 939 7624
rect 741 7426 797 7482
rect 883 7426 939 7482
rect 741 7284 797 7340
rect 883 7284 939 7340
rect 741 7142 797 7198
rect 883 7142 939 7198
rect 741 7000 797 7056
rect 883 7000 939 7056
rect 741 6858 797 6914
rect 883 6858 939 6914
rect 741 6716 797 6772
rect 883 6716 939 6772
rect 741 6574 797 6630
rect 883 6574 939 6630
rect 741 6432 797 6488
rect 883 6432 939 6488
rect 741 6290 797 6346
rect 883 6290 939 6346
rect 741 6148 797 6204
rect 883 6148 939 6204
rect 741 6006 797 6062
rect 883 6006 939 6062
rect 741 5864 797 5920
rect 883 5864 939 5920
rect 741 5722 797 5778
rect 883 5722 939 5778
rect 741 5580 797 5636
rect 883 5580 939 5636
rect 741 5438 797 5494
rect 883 5438 939 5494
rect 741 5296 797 5352
rect 883 5296 939 5352
rect 741 5154 797 5210
rect 883 5154 939 5210
rect 741 5012 797 5068
rect 883 5012 939 5068
rect 741 4870 797 4926
rect 883 4870 939 4926
rect 741 4728 797 4784
rect 883 4728 939 4784
rect 741 4586 797 4642
rect 883 4586 939 4642
rect 741 4444 797 4500
rect 883 4444 939 4500
rect 741 4302 797 4358
rect 883 4302 939 4358
rect 741 4160 797 4216
rect 883 4160 939 4216
rect 741 4018 797 4074
rect 883 4018 939 4074
rect 741 3876 797 3932
rect 883 3876 939 3932
rect 741 3734 797 3790
rect 883 3734 939 3790
rect 741 3592 797 3648
rect 883 3592 939 3648
rect 741 3450 797 3506
rect 883 3450 939 3506
rect 741 3308 797 3364
rect 883 3308 939 3364
rect 741 3166 797 3222
rect 883 3166 939 3222
rect 741 3024 797 3080
rect 883 3024 939 3080
rect 741 2882 797 2938
rect 883 2882 939 2938
rect 741 2740 797 2796
rect 883 2740 939 2796
rect 741 2598 797 2654
rect 883 2598 939 2654
rect 741 2456 797 2512
rect 883 2456 939 2512
rect 741 2314 797 2370
rect 883 2314 939 2370
rect 741 2172 797 2228
rect 883 2172 939 2228
rect 741 2030 797 2086
rect 883 2030 939 2086
rect 741 1888 797 1944
rect 883 1888 939 1944
rect 741 1746 797 1802
rect 883 1746 939 1802
rect 741 1604 797 1660
rect 883 1604 939 1660
rect 741 1462 797 1518
rect 883 1462 939 1518
rect 741 1320 797 1376
rect 883 1320 939 1376
rect 741 1178 797 1234
rect 883 1178 939 1234
rect 741 1036 797 1092
rect 883 1036 939 1092
rect 741 894 797 950
rect 883 894 939 950
rect 741 752 797 808
rect 883 752 939 808
rect 741 610 797 666
rect 883 610 939 666
rect 741 468 797 524
rect 883 468 939 524
rect 1142 12254 1198 12310
rect 1284 12254 1340 12310
rect 1142 12112 1198 12168
rect 1284 12112 1340 12168
rect 1142 11970 1198 12026
rect 1284 11970 1340 12026
rect 1142 11828 1198 11884
rect 1284 11828 1340 11884
rect 1142 11686 1198 11742
rect 1284 11686 1340 11742
rect 1142 11544 1198 11600
rect 1284 11544 1340 11600
rect 1142 11402 1198 11458
rect 1284 11402 1340 11458
rect 1142 11260 1198 11316
rect 1284 11260 1340 11316
rect 1142 11118 1198 11174
rect 1284 11118 1340 11174
rect 1142 10976 1198 11032
rect 1284 10976 1340 11032
rect 1142 10834 1198 10890
rect 1284 10834 1340 10890
rect 1142 10692 1198 10748
rect 1284 10692 1340 10748
rect 1142 10550 1198 10606
rect 1284 10550 1340 10606
rect 1142 10408 1198 10464
rect 1284 10408 1340 10464
rect 1142 10266 1198 10322
rect 1284 10266 1340 10322
rect 1142 10124 1198 10180
rect 1284 10124 1340 10180
rect 1142 9982 1198 10038
rect 1284 9982 1340 10038
rect 1142 9840 1198 9896
rect 1284 9840 1340 9896
rect 1142 9698 1198 9754
rect 1284 9698 1340 9754
rect 1142 9556 1198 9612
rect 1284 9556 1340 9612
rect 1142 9414 1198 9470
rect 1284 9414 1340 9470
rect 1142 9272 1198 9328
rect 1284 9272 1340 9328
rect 1142 9130 1198 9186
rect 1284 9130 1340 9186
rect 1142 8988 1198 9044
rect 1284 8988 1340 9044
rect 1142 8846 1198 8902
rect 1284 8846 1340 8902
rect 1142 8704 1198 8760
rect 1284 8704 1340 8760
rect 1142 8562 1198 8618
rect 1284 8562 1340 8618
rect 1142 8420 1198 8476
rect 1284 8420 1340 8476
rect 1142 8278 1198 8334
rect 1284 8278 1340 8334
rect 1142 8136 1198 8192
rect 1284 8136 1340 8192
rect 1142 7994 1198 8050
rect 1284 7994 1340 8050
rect 1142 7852 1198 7908
rect 1284 7852 1340 7908
rect 1142 7710 1198 7766
rect 1284 7710 1340 7766
rect 1142 7568 1198 7624
rect 1284 7568 1340 7624
rect 1142 7426 1198 7482
rect 1284 7426 1340 7482
rect 1142 7284 1198 7340
rect 1284 7284 1340 7340
rect 1142 7142 1198 7198
rect 1284 7142 1340 7198
rect 1142 7000 1198 7056
rect 1284 7000 1340 7056
rect 1142 6858 1198 6914
rect 1284 6858 1340 6914
rect 1142 6716 1198 6772
rect 1284 6716 1340 6772
rect 1142 6574 1198 6630
rect 1284 6574 1340 6630
rect 1142 6432 1198 6488
rect 1284 6432 1340 6488
rect 1142 6290 1198 6346
rect 1284 6290 1340 6346
rect 1142 6148 1198 6204
rect 1284 6148 1340 6204
rect 1142 6006 1198 6062
rect 1284 6006 1340 6062
rect 1142 5864 1198 5920
rect 1284 5864 1340 5920
rect 1142 5722 1198 5778
rect 1284 5722 1340 5778
rect 1142 5580 1198 5636
rect 1284 5580 1340 5636
rect 1142 5438 1198 5494
rect 1284 5438 1340 5494
rect 1142 5296 1198 5352
rect 1284 5296 1340 5352
rect 1142 5154 1198 5210
rect 1284 5154 1340 5210
rect 1142 5012 1198 5068
rect 1284 5012 1340 5068
rect 1142 4870 1198 4926
rect 1284 4870 1340 4926
rect 1142 4728 1198 4784
rect 1284 4728 1340 4784
rect 1142 4586 1198 4642
rect 1284 4586 1340 4642
rect 1142 4444 1198 4500
rect 1284 4444 1340 4500
rect 1142 4302 1198 4358
rect 1284 4302 1340 4358
rect 1142 4160 1198 4216
rect 1284 4160 1340 4216
rect 1142 4018 1198 4074
rect 1284 4018 1340 4074
rect 1142 3876 1198 3932
rect 1284 3876 1340 3932
rect 1142 3734 1198 3790
rect 1284 3734 1340 3790
rect 1142 3592 1198 3648
rect 1284 3592 1340 3648
rect 1142 3450 1198 3506
rect 1284 3450 1340 3506
rect 1142 3308 1198 3364
rect 1284 3308 1340 3364
rect 1142 3166 1198 3222
rect 1284 3166 1340 3222
rect 1142 3024 1198 3080
rect 1284 3024 1340 3080
rect 1142 2882 1198 2938
rect 1284 2882 1340 2938
rect 1142 2740 1198 2796
rect 1284 2740 1340 2796
rect 1142 2598 1198 2654
rect 1284 2598 1340 2654
rect 1142 2456 1198 2512
rect 1284 2456 1340 2512
rect 1142 2314 1198 2370
rect 1284 2314 1340 2370
rect 1142 2172 1198 2228
rect 1284 2172 1340 2228
rect 1142 2030 1198 2086
rect 1284 2030 1340 2086
rect 1142 1888 1198 1944
rect 1284 1888 1340 1944
rect 1142 1746 1198 1802
rect 1284 1746 1340 1802
rect 1142 1604 1198 1660
rect 1284 1604 1340 1660
rect 1142 1462 1198 1518
rect 1284 1462 1340 1518
rect 1142 1320 1198 1376
rect 1284 1320 1340 1376
rect 1142 1178 1198 1234
rect 1284 1178 1340 1234
rect 1142 1036 1198 1092
rect 1284 1036 1340 1092
rect 1142 894 1198 950
rect 1284 894 1340 950
rect 1142 752 1198 808
rect 1284 752 1340 808
rect 1142 610 1198 666
rect 1284 610 1340 666
rect 1142 468 1198 524
rect 1284 468 1340 524
rect 1542 12254 1598 12310
rect 1684 12254 1740 12310
rect 1542 12112 1598 12168
rect 1684 12112 1740 12168
rect 1542 11970 1598 12026
rect 1684 11970 1740 12026
rect 1542 11828 1598 11884
rect 1684 11828 1740 11884
rect 1542 11686 1598 11742
rect 1684 11686 1740 11742
rect 1542 11544 1598 11600
rect 1684 11544 1740 11600
rect 1542 11402 1598 11458
rect 1684 11402 1740 11458
rect 1542 11260 1598 11316
rect 1684 11260 1740 11316
rect 1542 11118 1598 11174
rect 1684 11118 1740 11174
rect 1542 10976 1598 11032
rect 1684 10976 1740 11032
rect 1542 10834 1598 10890
rect 1684 10834 1740 10890
rect 1542 10692 1598 10748
rect 1684 10692 1740 10748
rect 1542 10550 1598 10606
rect 1684 10550 1740 10606
rect 1542 10408 1598 10464
rect 1684 10408 1740 10464
rect 1542 10266 1598 10322
rect 1684 10266 1740 10322
rect 1542 10124 1598 10180
rect 1684 10124 1740 10180
rect 1542 9982 1598 10038
rect 1684 9982 1740 10038
rect 1542 9840 1598 9896
rect 1684 9840 1740 9896
rect 1542 9698 1598 9754
rect 1684 9698 1740 9754
rect 1542 9556 1598 9612
rect 1684 9556 1740 9612
rect 1542 9414 1598 9470
rect 1684 9414 1740 9470
rect 1542 9272 1598 9328
rect 1684 9272 1740 9328
rect 1542 9130 1598 9186
rect 1684 9130 1740 9186
rect 1542 8988 1598 9044
rect 1684 8988 1740 9044
rect 1542 8846 1598 8902
rect 1684 8846 1740 8902
rect 1542 8704 1598 8760
rect 1684 8704 1740 8760
rect 1542 8562 1598 8618
rect 1684 8562 1740 8618
rect 1542 8420 1598 8476
rect 1684 8420 1740 8476
rect 1542 8278 1598 8334
rect 1684 8278 1740 8334
rect 1542 8136 1598 8192
rect 1684 8136 1740 8192
rect 1542 7994 1598 8050
rect 1684 7994 1740 8050
rect 1542 7852 1598 7908
rect 1684 7852 1740 7908
rect 1542 7710 1598 7766
rect 1684 7710 1740 7766
rect 1542 7568 1598 7624
rect 1684 7568 1740 7624
rect 1542 7426 1598 7482
rect 1684 7426 1740 7482
rect 1542 7284 1598 7340
rect 1684 7284 1740 7340
rect 1542 7142 1598 7198
rect 1684 7142 1740 7198
rect 1542 7000 1598 7056
rect 1684 7000 1740 7056
rect 1542 6858 1598 6914
rect 1684 6858 1740 6914
rect 1542 6716 1598 6772
rect 1684 6716 1740 6772
rect 1542 6574 1598 6630
rect 1684 6574 1740 6630
rect 1542 6432 1598 6488
rect 1684 6432 1740 6488
rect 1542 6290 1598 6346
rect 1684 6290 1740 6346
rect 1542 6148 1598 6204
rect 1684 6148 1740 6204
rect 1542 6006 1598 6062
rect 1684 6006 1740 6062
rect 1542 5864 1598 5920
rect 1684 5864 1740 5920
rect 1542 5722 1598 5778
rect 1684 5722 1740 5778
rect 1542 5580 1598 5636
rect 1684 5580 1740 5636
rect 1542 5438 1598 5494
rect 1684 5438 1740 5494
rect 1542 5296 1598 5352
rect 1684 5296 1740 5352
rect 1542 5154 1598 5210
rect 1684 5154 1740 5210
rect 1542 5012 1598 5068
rect 1684 5012 1740 5068
rect 1542 4870 1598 4926
rect 1684 4870 1740 4926
rect 1542 4728 1598 4784
rect 1684 4728 1740 4784
rect 1542 4586 1598 4642
rect 1684 4586 1740 4642
rect 1542 4444 1598 4500
rect 1684 4444 1740 4500
rect 1542 4302 1598 4358
rect 1684 4302 1740 4358
rect 1542 4160 1598 4216
rect 1684 4160 1740 4216
rect 1542 4018 1598 4074
rect 1684 4018 1740 4074
rect 1542 3876 1598 3932
rect 1684 3876 1740 3932
rect 1542 3734 1598 3790
rect 1684 3734 1740 3790
rect 1542 3592 1598 3648
rect 1684 3592 1740 3648
rect 1542 3450 1598 3506
rect 1684 3450 1740 3506
rect 1542 3308 1598 3364
rect 1684 3308 1740 3364
rect 1542 3166 1598 3222
rect 1684 3166 1740 3222
rect 1542 3024 1598 3080
rect 1684 3024 1740 3080
rect 1542 2882 1598 2938
rect 1684 2882 1740 2938
rect 1542 2740 1598 2796
rect 1684 2740 1740 2796
rect 1542 2598 1598 2654
rect 1684 2598 1740 2654
rect 1542 2456 1598 2512
rect 1684 2456 1740 2512
rect 1542 2314 1598 2370
rect 1684 2314 1740 2370
rect 1542 2172 1598 2228
rect 1684 2172 1740 2228
rect 1542 2030 1598 2086
rect 1684 2030 1740 2086
rect 1542 1888 1598 1944
rect 1684 1888 1740 1944
rect 1542 1746 1598 1802
rect 1684 1746 1740 1802
rect 1542 1604 1598 1660
rect 1684 1604 1740 1660
rect 1542 1462 1598 1518
rect 1684 1462 1740 1518
rect 1542 1320 1598 1376
rect 1684 1320 1740 1376
rect 1542 1178 1598 1234
rect 1684 1178 1740 1234
rect 1542 1036 1598 1092
rect 1684 1036 1740 1092
rect 1542 894 1598 950
rect 1684 894 1740 950
rect 1542 752 1598 808
rect 1684 752 1740 808
rect 1542 610 1598 666
rect 1684 610 1740 666
rect 1542 468 1598 524
rect 1684 468 1740 524
rect 1939 12254 1995 12310
rect 2081 12254 2137 12310
rect 1939 12112 1995 12168
rect 2081 12112 2137 12168
rect 1939 11970 1995 12026
rect 2081 11970 2137 12026
rect 1939 11828 1995 11884
rect 2081 11828 2137 11884
rect 1939 11686 1995 11742
rect 2081 11686 2137 11742
rect 1939 11544 1995 11600
rect 2081 11544 2137 11600
rect 1939 11402 1995 11458
rect 2081 11402 2137 11458
rect 1939 11260 1995 11316
rect 2081 11260 2137 11316
rect 1939 11118 1995 11174
rect 2081 11118 2137 11174
rect 1939 10976 1995 11032
rect 2081 10976 2137 11032
rect 1939 10834 1995 10890
rect 2081 10834 2137 10890
rect 1939 10692 1995 10748
rect 2081 10692 2137 10748
rect 1939 10550 1995 10606
rect 2081 10550 2137 10606
rect 1939 10408 1995 10464
rect 2081 10408 2137 10464
rect 1939 10266 1995 10322
rect 2081 10266 2137 10322
rect 1939 10124 1995 10180
rect 2081 10124 2137 10180
rect 1939 9982 1995 10038
rect 2081 9982 2137 10038
rect 1939 9840 1995 9896
rect 2081 9840 2137 9896
rect 1939 9698 1995 9754
rect 2081 9698 2137 9754
rect 1939 9556 1995 9612
rect 2081 9556 2137 9612
rect 1939 9414 1995 9470
rect 2081 9414 2137 9470
rect 1939 9272 1995 9328
rect 2081 9272 2137 9328
rect 1939 9130 1995 9186
rect 2081 9130 2137 9186
rect 1939 8988 1995 9044
rect 2081 8988 2137 9044
rect 1939 8846 1995 8902
rect 2081 8846 2137 8902
rect 1939 8704 1995 8760
rect 2081 8704 2137 8760
rect 1939 8562 1995 8618
rect 2081 8562 2137 8618
rect 1939 8420 1995 8476
rect 2081 8420 2137 8476
rect 1939 8278 1995 8334
rect 2081 8278 2137 8334
rect 1939 8136 1995 8192
rect 2081 8136 2137 8192
rect 1939 7994 1995 8050
rect 2081 7994 2137 8050
rect 1939 7852 1995 7908
rect 2081 7852 2137 7908
rect 1939 7710 1995 7766
rect 2081 7710 2137 7766
rect 1939 7568 1995 7624
rect 2081 7568 2137 7624
rect 1939 7426 1995 7482
rect 2081 7426 2137 7482
rect 1939 7284 1995 7340
rect 2081 7284 2137 7340
rect 1939 7142 1995 7198
rect 2081 7142 2137 7198
rect 1939 7000 1995 7056
rect 2081 7000 2137 7056
rect 1939 6858 1995 6914
rect 2081 6858 2137 6914
rect 1939 6716 1995 6772
rect 2081 6716 2137 6772
rect 1939 6574 1995 6630
rect 2081 6574 2137 6630
rect 1939 6432 1995 6488
rect 2081 6432 2137 6488
rect 1939 6290 1995 6346
rect 2081 6290 2137 6346
rect 1939 6148 1995 6204
rect 2081 6148 2137 6204
rect 1939 6006 1995 6062
rect 2081 6006 2137 6062
rect 1939 5864 1995 5920
rect 2081 5864 2137 5920
rect 1939 5722 1995 5778
rect 2081 5722 2137 5778
rect 1939 5580 1995 5636
rect 2081 5580 2137 5636
rect 1939 5438 1995 5494
rect 2081 5438 2137 5494
rect 1939 5296 1995 5352
rect 2081 5296 2137 5352
rect 1939 5154 1995 5210
rect 2081 5154 2137 5210
rect 1939 5012 1995 5068
rect 2081 5012 2137 5068
rect 1939 4870 1995 4926
rect 2081 4870 2137 4926
rect 1939 4728 1995 4784
rect 2081 4728 2137 4784
rect 1939 4586 1995 4642
rect 2081 4586 2137 4642
rect 1939 4444 1995 4500
rect 2081 4444 2137 4500
rect 1939 4302 1995 4358
rect 2081 4302 2137 4358
rect 1939 4160 1995 4216
rect 2081 4160 2137 4216
rect 1939 4018 1995 4074
rect 2081 4018 2137 4074
rect 1939 3876 1995 3932
rect 2081 3876 2137 3932
rect 1939 3734 1995 3790
rect 2081 3734 2137 3790
rect 1939 3592 1995 3648
rect 2081 3592 2137 3648
rect 1939 3450 1995 3506
rect 2081 3450 2137 3506
rect 1939 3308 1995 3364
rect 2081 3308 2137 3364
rect 1939 3166 1995 3222
rect 2081 3166 2137 3222
rect 1939 3024 1995 3080
rect 2081 3024 2137 3080
rect 1939 2882 1995 2938
rect 2081 2882 2137 2938
rect 1939 2740 1995 2796
rect 2081 2740 2137 2796
rect 1939 2598 1995 2654
rect 2081 2598 2137 2654
rect 1939 2456 1995 2512
rect 2081 2456 2137 2512
rect 1939 2314 1995 2370
rect 2081 2314 2137 2370
rect 1939 2172 1995 2228
rect 2081 2172 2137 2228
rect 1939 2030 1995 2086
rect 2081 2030 2137 2086
rect 1939 1888 1995 1944
rect 2081 1888 2137 1944
rect 1939 1746 1995 1802
rect 2081 1746 2137 1802
rect 1939 1604 1995 1660
rect 2081 1604 2137 1660
rect 1939 1462 1995 1518
rect 2081 1462 2137 1518
rect 1939 1320 1995 1376
rect 2081 1320 2137 1376
rect 1939 1178 1995 1234
rect 2081 1178 2137 1234
rect 1939 1036 1995 1092
rect 2081 1036 2137 1092
rect 1939 894 1995 950
rect 2081 894 2137 950
rect 1939 752 1995 808
rect 2081 752 2137 808
rect 1939 610 1995 666
rect 2081 610 2137 666
rect 1939 468 1995 524
rect 2081 468 2137 524
rect 2336 12254 2392 12310
rect 2478 12254 2534 12310
rect 2336 12112 2392 12168
rect 2478 12112 2534 12168
rect 2336 11970 2392 12026
rect 2478 11970 2534 12026
rect 2336 11828 2392 11884
rect 2478 11828 2534 11884
rect 2336 11686 2392 11742
rect 2478 11686 2534 11742
rect 2336 11544 2392 11600
rect 2478 11544 2534 11600
rect 2336 11402 2392 11458
rect 2478 11402 2534 11458
rect 2336 11260 2392 11316
rect 2478 11260 2534 11316
rect 2336 11118 2392 11174
rect 2478 11118 2534 11174
rect 2336 10976 2392 11032
rect 2478 10976 2534 11032
rect 2336 10834 2392 10890
rect 2478 10834 2534 10890
rect 2336 10692 2392 10748
rect 2478 10692 2534 10748
rect 2336 10550 2392 10606
rect 2478 10550 2534 10606
rect 2336 10408 2392 10464
rect 2478 10408 2534 10464
rect 2336 10266 2392 10322
rect 2478 10266 2534 10322
rect 2336 10124 2392 10180
rect 2478 10124 2534 10180
rect 2336 9982 2392 10038
rect 2478 9982 2534 10038
rect 2336 9840 2392 9896
rect 2478 9840 2534 9896
rect 2336 9698 2392 9754
rect 2478 9698 2534 9754
rect 2336 9556 2392 9612
rect 2478 9556 2534 9612
rect 2336 9414 2392 9470
rect 2478 9414 2534 9470
rect 2336 9272 2392 9328
rect 2478 9272 2534 9328
rect 2336 9130 2392 9186
rect 2478 9130 2534 9186
rect 2336 8988 2392 9044
rect 2478 8988 2534 9044
rect 2336 8846 2392 8902
rect 2478 8846 2534 8902
rect 2336 8704 2392 8760
rect 2478 8704 2534 8760
rect 2336 8562 2392 8618
rect 2478 8562 2534 8618
rect 2336 8420 2392 8476
rect 2478 8420 2534 8476
rect 2336 8278 2392 8334
rect 2478 8278 2534 8334
rect 2336 8136 2392 8192
rect 2478 8136 2534 8192
rect 2336 7994 2392 8050
rect 2478 7994 2534 8050
rect 2336 7852 2392 7908
rect 2478 7852 2534 7908
rect 2336 7710 2392 7766
rect 2478 7710 2534 7766
rect 2336 7568 2392 7624
rect 2478 7568 2534 7624
rect 2336 7426 2392 7482
rect 2478 7426 2534 7482
rect 2336 7284 2392 7340
rect 2478 7284 2534 7340
rect 2336 7142 2392 7198
rect 2478 7142 2534 7198
rect 2336 7000 2392 7056
rect 2478 7000 2534 7056
rect 2336 6858 2392 6914
rect 2478 6858 2534 6914
rect 2336 6716 2392 6772
rect 2478 6716 2534 6772
rect 2336 6574 2392 6630
rect 2478 6574 2534 6630
rect 2336 6432 2392 6488
rect 2478 6432 2534 6488
rect 2336 6290 2392 6346
rect 2478 6290 2534 6346
rect 2336 6148 2392 6204
rect 2478 6148 2534 6204
rect 2336 6006 2392 6062
rect 2478 6006 2534 6062
rect 2336 5864 2392 5920
rect 2478 5864 2534 5920
rect 2336 5722 2392 5778
rect 2478 5722 2534 5778
rect 2336 5580 2392 5636
rect 2478 5580 2534 5636
rect 2336 5438 2392 5494
rect 2478 5438 2534 5494
rect 2336 5296 2392 5352
rect 2478 5296 2534 5352
rect 2336 5154 2392 5210
rect 2478 5154 2534 5210
rect 2336 5012 2392 5068
rect 2478 5012 2534 5068
rect 2336 4870 2392 4926
rect 2478 4870 2534 4926
rect 2336 4728 2392 4784
rect 2478 4728 2534 4784
rect 2336 4586 2392 4642
rect 2478 4586 2534 4642
rect 2336 4444 2392 4500
rect 2478 4444 2534 4500
rect 2336 4302 2392 4358
rect 2478 4302 2534 4358
rect 2336 4160 2392 4216
rect 2478 4160 2534 4216
rect 2336 4018 2392 4074
rect 2478 4018 2534 4074
rect 2336 3876 2392 3932
rect 2478 3876 2534 3932
rect 2336 3734 2392 3790
rect 2478 3734 2534 3790
rect 2336 3592 2392 3648
rect 2478 3592 2534 3648
rect 2336 3450 2392 3506
rect 2478 3450 2534 3506
rect 2336 3308 2392 3364
rect 2478 3308 2534 3364
rect 2336 3166 2392 3222
rect 2478 3166 2534 3222
rect 2336 3024 2392 3080
rect 2478 3024 2534 3080
rect 2336 2882 2392 2938
rect 2478 2882 2534 2938
rect 2336 2740 2392 2796
rect 2478 2740 2534 2796
rect 2336 2598 2392 2654
rect 2478 2598 2534 2654
rect 2336 2456 2392 2512
rect 2478 2456 2534 2512
rect 2336 2314 2392 2370
rect 2478 2314 2534 2370
rect 2336 2172 2392 2228
rect 2478 2172 2534 2228
rect 2336 2030 2392 2086
rect 2478 2030 2534 2086
rect 2336 1888 2392 1944
rect 2478 1888 2534 1944
rect 2336 1746 2392 1802
rect 2478 1746 2534 1802
rect 2336 1604 2392 1660
rect 2478 1604 2534 1660
rect 2336 1462 2392 1518
rect 2478 1462 2534 1518
rect 2336 1320 2392 1376
rect 2478 1320 2534 1376
rect 2336 1178 2392 1234
rect 2478 1178 2534 1234
rect 2336 1036 2392 1092
rect 2478 1036 2534 1092
rect 2336 894 2392 950
rect 2478 894 2534 950
rect 2336 752 2392 808
rect 2478 752 2534 808
rect 2336 610 2392 666
rect 2478 610 2534 666
rect 2336 468 2392 524
rect 2478 468 2534 524
rect 2740 12254 2796 12310
rect 2882 12254 2938 12310
rect 2740 12112 2796 12168
rect 2882 12112 2938 12168
rect 2740 11970 2796 12026
rect 2882 11970 2938 12026
rect 2740 11828 2796 11884
rect 2882 11828 2938 11884
rect 2740 11686 2796 11742
rect 2882 11686 2938 11742
rect 2740 11544 2796 11600
rect 2882 11544 2938 11600
rect 2740 11402 2796 11458
rect 2882 11402 2938 11458
rect 2740 11260 2796 11316
rect 2882 11260 2938 11316
rect 2740 11118 2796 11174
rect 2882 11118 2938 11174
rect 2740 10976 2796 11032
rect 2882 10976 2938 11032
rect 2740 10834 2796 10890
rect 2882 10834 2938 10890
rect 2740 10692 2796 10748
rect 2882 10692 2938 10748
rect 2740 10550 2796 10606
rect 2882 10550 2938 10606
rect 2740 10408 2796 10464
rect 2882 10408 2938 10464
rect 2740 10266 2796 10322
rect 2882 10266 2938 10322
rect 2740 10124 2796 10180
rect 2882 10124 2938 10180
rect 2740 9982 2796 10038
rect 2882 9982 2938 10038
rect 2740 9840 2796 9896
rect 2882 9840 2938 9896
rect 2740 9698 2796 9754
rect 2882 9698 2938 9754
rect 2740 9556 2796 9612
rect 2882 9556 2938 9612
rect 2740 9414 2796 9470
rect 2882 9414 2938 9470
rect 2740 9272 2796 9328
rect 2882 9272 2938 9328
rect 2740 9130 2796 9186
rect 2882 9130 2938 9186
rect 2740 8988 2796 9044
rect 2882 8988 2938 9044
rect 2740 8846 2796 8902
rect 2882 8846 2938 8902
rect 2740 8704 2796 8760
rect 2882 8704 2938 8760
rect 2740 8562 2796 8618
rect 2882 8562 2938 8618
rect 2740 8420 2796 8476
rect 2882 8420 2938 8476
rect 2740 8278 2796 8334
rect 2882 8278 2938 8334
rect 2740 8136 2796 8192
rect 2882 8136 2938 8192
rect 2740 7994 2796 8050
rect 2882 7994 2938 8050
rect 2740 7852 2796 7908
rect 2882 7852 2938 7908
rect 2740 7710 2796 7766
rect 2882 7710 2938 7766
rect 2740 7568 2796 7624
rect 2882 7568 2938 7624
rect 2740 7426 2796 7482
rect 2882 7426 2938 7482
rect 2740 7284 2796 7340
rect 2882 7284 2938 7340
rect 2740 7142 2796 7198
rect 2882 7142 2938 7198
rect 2740 7000 2796 7056
rect 2882 7000 2938 7056
rect 2740 6858 2796 6914
rect 2882 6858 2938 6914
rect 2740 6716 2796 6772
rect 2882 6716 2938 6772
rect 2740 6574 2796 6630
rect 2882 6574 2938 6630
rect 2740 6432 2796 6488
rect 2882 6432 2938 6488
rect 2740 6290 2796 6346
rect 2882 6290 2938 6346
rect 2740 6148 2796 6204
rect 2882 6148 2938 6204
rect 2740 6006 2796 6062
rect 2882 6006 2938 6062
rect 2740 5864 2796 5920
rect 2882 5864 2938 5920
rect 2740 5722 2796 5778
rect 2882 5722 2938 5778
rect 2740 5580 2796 5636
rect 2882 5580 2938 5636
rect 2740 5438 2796 5494
rect 2882 5438 2938 5494
rect 2740 5296 2796 5352
rect 2882 5296 2938 5352
rect 2740 5154 2796 5210
rect 2882 5154 2938 5210
rect 2740 5012 2796 5068
rect 2882 5012 2938 5068
rect 2740 4870 2796 4926
rect 2882 4870 2938 4926
rect 2740 4728 2796 4784
rect 2882 4728 2938 4784
rect 2740 4586 2796 4642
rect 2882 4586 2938 4642
rect 2740 4444 2796 4500
rect 2882 4444 2938 4500
rect 2740 4302 2796 4358
rect 2882 4302 2938 4358
rect 2740 4160 2796 4216
rect 2882 4160 2938 4216
rect 2740 4018 2796 4074
rect 2882 4018 2938 4074
rect 2740 3876 2796 3932
rect 2882 3876 2938 3932
rect 2740 3734 2796 3790
rect 2882 3734 2938 3790
rect 2740 3592 2796 3648
rect 2882 3592 2938 3648
rect 2740 3450 2796 3506
rect 2882 3450 2938 3506
rect 2740 3308 2796 3364
rect 2882 3308 2938 3364
rect 2740 3166 2796 3222
rect 2882 3166 2938 3222
rect 2740 3024 2796 3080
rect 2882 3024 2938 3080
rect 2740 2882 2796 2938
rect 2882 2882 2938 2938
rect 2740 2740 2796 2796
rect 2882 2740 2938 2796
rect 2740 2598 2796 2654
rect 2882 2598 2938 2654
rect 2740 2456 2796 2512
rect 2882 2456 2938 2512
rect 2740 2314 2796 2370
rect 2882 2314 2938 2370
rect 2740 2172 2796 2228
rect 2882 2172 2938 2228
rect 2740 2030 2796 2086
rect 2882 2030 2938 2086
rect 2740 1888 2796 1944
rect 2882 1888 2938 1944
rect 2740 1746 2796 1802
rect 2882 1746 2938 1802
rect 2740 1604 2796 1660
rect 2882 1604 2938 1660
rect 2740 1462 2796 1518
rect 2882 1462 2938 1518
rect 2740 1320 2796 1376
rect 2882 1320 2938 1376
rect 2740 1178 2796 1234
rect 2882 1178 2938 1234
rect 2740 1036 2796 1092
rect 2882 1036 2938 1092
rect 2740 894 2796 950
rect 2882 894 2938 950
rect 2740 752 2796 808
rect 2882 752 2938 808
rect 2740 610 2796 666
rect 2882 610 2938 666
rect 2740 468 2796 524
rect 2882 468 2938 524
rect 3136 12254 3192 12310
rect 3278 12254 3334 12310
rect 3136 12112 3192 12168
rect 3278 12112 3334 12168
rect 3136 11970 3192 12026
rect 3278 11970 3334 12026
rect 3136 11828 3192 11884
rect 3278 11828 3334 11884
rect 3136 11686 3192 11742
rect 3278 11686 3334 11742
rect 3136 11544 3192 11600
rect 3278 11544 3334 11600
rect 3136 11402 3192 11458
rect 3278 11402 3334 11458
rect 3136 11260 3192 11316
rect 3278 11260 3334 11316
rect 3136 11118 3192 11174
rect 3278 11118 3334 11174
rect 3136 10976 3192 11032
rect 3278 10976 3334 11032
rect 3136 10834 3192 10890
rect 3278 10834 3334 10890
rect 3136 10692 3192 10748
rect 3278 10692 3334 10748
rect 3136 10550 3192 10606
rect 3278 10550 3334 10606
rect 3136 10408 3192 10464
rect 3278 10408 3334 10464
rect 3136 10266 3192 10322
rect 3278 10266 3334 10322
rect 3136 10124 3192 10180
rect 3278 10124 3334 10180
rect 3136 9982 3192 10038
rect 3278 9982 3334 10038
rect 3136 9840 3192 9896
rect 3278 9840 3334 9896
rect 3136 9698 3192 9754
rect 3278 9698 3334 9754
rect 3136 9556 3192 9612
rect 3278 9556 3334 9612
rect 3136 9414 3192 9470
rect 3278 9414 3334 9470
rect 3136 9272 3192 9328
rect 3278 9272 3334 9328
rect 3136 9130 3192 9186
rect 3278 9130 3334 9186
rect 3136 8988 3192 9044
rect 3278 8988 3334 9044
rect 3136 8846 3192 8902
rect 3278 8846 3334 8902
rect 3136 8704 3192 8760
rect 3278 8704 3334 8760
rect 3136 8562 3192 8618
rect 3278 8562 3334 8618
rect 3136 8420 3192 8476
rect 3278 8420 3334 8476
rect 3136 8278 3192 8334
rect 3278 8278 3334 8334
rect 3136 8136 3192 8192
rect 3278 8136 3334 8192
rect 3136 7994 3192 8050
rect 3278 7994 3334 8050
rect 3136 7852 3192 7908
rect 3278 7852 3334 7908
rect 3136 7710 3192 7766
rect 3278 7710 3334 7766
rect 3136 7568 3192 7624
rect 3278 7568 3334 7624
rect 3136 7426 3192 7482
rect 3278 7426 3334 7482
rect 3136 7284 3192 7340
rect 3278 7284 3334 7340
rect 3136 7142 3192 7198
rect 3278 7142 3334 7198
rect 3136 7000 3192 7056
rect 3278 7000 3334 7056
rect 3136 6858 3192 6914
rect 3278 6858 3334 6914
rect 3136 6716 3192 6772
rect 3278 6716 3334 6772
rect 3136 6574 3192 6630
rect 3278 6574 3334 6630
rect 3136 6432 3192 6488
rect 3278 6432 3334 6488
rect 3136 6290 3192 6346
rect 3278 6290 3334 6346
rect 3136 6148 3192 6204
rect 3278 6148 3334 6204
rect 3136 6006 3192 6062
rect 3278 6006 3334 6062
rect 3136 5864 3192 5920
rect 3278 5864 3334 5920
rect 3136 5722 3192 5778
rect 3278 5722 3334 5778
rect 3136 5580 3192 5636
rect 3278 5580 3334 5636
rect 3136 5438 3192 5494
rect 3278 5438 3334 5494
rect 3136 5296 3192 5352
rect 3278 5296 3334 5352
rect 3136 5154 3192 5210
rect 3278 5154 3334 5210
rect 3136 5012 3192 5068
rect 3278 5012 3334 5068
rect 3136 4870 3192 4926
rect 3278 4870 3334 4926
rect 3136 4728 3192 4784
rect 3278 4728 3334 4784
rect 3136 4586 3192 4642
rect 3278 4586 3334 4642
rect 3136 4444 3192 4500
rect 3278 4444 3334 4500
rect 3136 4302 3192 4358
rect 3278 4302 3334 4358
rect 3136 4160 3192 4216
rect 3278 4160 3334 4216
rect 3136 4018 3192 4074
rect 3278 4018 3334 4074
rect 3136 3876 3192 3932
rect 3278 3876 3334 3932
rect 3136 3734 3192 3790
rect 3278 3734 3334 3790
rect 3136 3592 3192 3648
rect 3278 3592 3334 3648
rect 3136 3450 3192 3506
rect 3278 3450 3334 3506
rect 3136 3308 3192 3364
rect 3278 3308 3334 3364
rect 3136 3166 3192 3222
rect 3278 3166 3334 3222
rect 3136 3024 3192 3080
rect 3278 3024 3334 3080
rect 3136 2882 3192 2938
rect 3278 2882 3334 2938
rect 3136 2740 3192 2796
rect 3278 2740 3334 2796
rect 3136 2598 3192 2654
rect 3278 2598 3334 2654
rect 3136 2456 3192 2512
rect 3278 2456 3334 2512
rect 3136 2314 3192 2370
rect 3278 2314 3334 2370
rect 3136 2172 3192 2228
rect 3278 2172 3334 2228
rect 3136 2030 3192 2086
rect 3278 2030 3334 2086
rect 3136 1888 3192 1944
rect 3278 1888 3334 1944
rect 3136 1746 3192 1802
rect 3278 1746 3334 1802
rect 3136 1604 3192 1660
rect 3278 1604 3334 1660
rect 3136 1462 3192 1518
rect 3278 1462 3334 1518
rect 3136 1320 3192 1376
rect 3278 1320 3334 1376
rect 3136 1178 3192 1234
rect 3278 1178 3334 1234
rect 3136 1036 3192 1092
rect 3278 1036 3334 1092
rect 3136 894 3192 950
rect 3278 894 3334 950
rect 3136 752 3192 808
rect 3278 752 3334 808
rect 3136 610 3192 666
rect 3278 610 3334 666
rect 3136 468 3192 524
rect 3278 468 3334 524
rect 3536 12254 3592 12310
rect 3678 12254 3734 12310
rect 3536 12112 3592 12168
rect 3678 12112 3734 12168
rect 3536 11970 3592 12026
rect 3678 11970 3734 12026
rect 3536 11828 3592 11884
rect 3678 11828 3734 11884
rect 3536 11686 3592 11742
rect 3678 11686 3734 11742
rect 3536 11544 3592 11600
rect 3678 11544 3734 11600
rect 3536 11402 3592 11458
rect 3678 11402 3734 11458
rect 3536 11260 3592 11316
rect 3678 11260 3734 11316
rect 3536 11118 3592 11174
rect 3678 11118 3734 11174
rect 3536 10976 3592 11032
rect 3678 10976 3734 11032
rect 3536 10834 3592 10890
rect 3678 10834 3734 10890
rect 3536 10692 3592 10748
rect 3678 10692 3734 10748
rect 3536 10550 3592 10606
rect 3678 10550 3734 10606
rect 3536 10408 3592 10464
rect 3678 10408 3734 10464
rect 3536 10266 3592 10322
rect 3678 10266 3734 10322
rect 3536 10124 3592 10180
rect 3678 10124 3734 10180
rect 3536 9982 3592 10038
rect 3678 9982 3734 10038
rect 3536 9840 3592 9896
rect 3678 9840 3734 9896
rect 3536 9698 3592 9754
rect 3678 9698 3734 9754
rect 3536 9556 3592 9612
rect 3678 9556 3734 9612
rect 3536 9414 3592 9470
rect 3678 9414 3734 9470
rect 3536 9272 3592 9328
rect 3678 9272 3734 9328
rect 3536 9130 3592 9186
rect 3678 9130 3734 9186
rect 3536 8988 3592 9044
rect 3678 8988 3734 9044
rect 3536 8846 3592 8902
rect 3678 8846 3734 8902
rect 3536 8704 3592 8760
rect 3678 8704 3734 8760
rect 3536 8562 3592 8618
rect 3678 8562 3734 8618
rect 3536 8420 3592 8476
rect 3678 8420 3734 8476
rect 3536 8278 3592 8334
rect 3678 8278 3734 8334
rect 3536 8136 3592 8192
rect 3678 8136 3734 8192
rect 3536 7994 3592 8050
rect 3678 7994 3734 8050
rect 3536 7852 3592 7908
rect 3678 7852 3734 7908
rect 3536 7710 3592 7766
rect 3678 7710 3734 7766
rect 3536 7568 3592 7624
rect 3678 7568 3734 7624
rect 3536 7426 3592 7482
rect 3678 7426 3734 7482
rect 3536 7284 3592 7340
rect 3678 7284 3734 7340
rect 3536 7142 3592 7198
rect 3678 7142 3734 7198
rect 3536 7000 3592 7056
rect 3678 7000 3734 7056
rect 3536 6858 3592 6914
rect 3678 6858 3734 6914
rect 3536 6716 3592 6772
rect 3678 6716 3734 6772
rect 3536 6574 3592 6630
rect 3678 6574 3734 6630
rect 3536 6432 3592 6488
rect 3678 6432 3734 6488
rect 3536 6290 3592 6346
rect 3678 6290 3734 6346
rect 3536 6148 3592 6204
rect 3678 6148 3734 6204
rect 3536 6006 3592 6062
rect 3678 6006 3734 6062
rect 3536 5864 3592 5920
rect 3678 5864 3734 5920
rect 3536 5722 3592 5778
rect 3678 5722 3734 5778
rect 3536 5580 3592 5636
rect 3678 5580 3734 5636
rect 3536 5438 3592 5494
rect 3678 5438 3734 5494
rect 3536 5296 3592 5352
rect 3678 5296 3734 5352
rect 3536 5154 3592 5210
rect 3678 5154 3734 5210
rect 3536 5012 3592 5068
rect 3678 5012 3734 5068
rect 3536 4870 3592 4926
rect 3678 4870 3734 4926
rect 3536 4728 3592 4784
rect 3678 4728 3734 4784
rect 3536 4586 3592 4642
rect 3678 4586 3734 4642
rect 3536 4444 3592 4500
rect 3678 4444 3734 4500
rect 3536 4302 3592 4358
rect 3678 4302 3734 4358
rect 3536 4160 3592 4216
rect 3678 4160 3734 4216
rect 3536 4018 3592 4074
rect 3678 4018 3734 4074
rect 3536 3876 3592 3932
rect 3678 3876 3734 3932
rect 3536 3734 3592 3790
rect 3678 3734 3734 3790
rect 3536 3592 3592 3648
rect 3678 3592 3734 3648
rect 3536 3450 3592 3506
rect 3678 3450 3734 3506
rect 3536 3308 3592 3364
rect 3678 3308 3734 3364
rect 3536 3166 3592 3222
rect 3678 3166 3734 3222
rect 3536 3024 3592 3080
rect 3678 3024 3734 3080
rect 3536 2882 3592 2938
rect 3678 2882 3734 2938
rect 3536 2740 3592 2796
rect 3678 2740 3734 2796
rect 3536 2598 3592 2654
rect 3678 2598 3734 2654
rect 3536 2456 3592 2512
rect 3678 2456 3734 2512
rect 3536 2314 3592 2370
rect 3678 2314 3734 2370
rect 3536 2172 3592 2228
rect 3678 2172 3734 2228
rect 3536 2030 3592 2086
rect 3678 2030 3734 2086
rect 3536 1888 3592 1944
rect 3678 1888 3734 1944
rect 3536 1746 3592 1802
rect 3678 1746 3734 1802
rect 3536 1604 3592 1660
rect 3678 1604 3734 1660
rect 3536 1462 3592 1518
rect 3678 1462 3734 1518
rect 3536 1320 3592 1376
rect 3678 1320 3734 1376
rect 3536 1178 3592 1234
rect 3678 1178 3734 1234
rect 3536 1036 3592 1092
rect 3678 1036 3734 1092
rect 3536 894 3592 950
rect 3678 894 3734 950
rect 3536 752 3592 808
rect 3678 752 3734 808
rect 3536 610 3592 666
rect 3678 610 3734 666
rect 3536 468 3592 524
rect 3678 468 3734 524
rect 3933 12254 3989 12310
rect 4075 12254 4131 12310
rect 3933 12112 3989 12168
rect 4075 12112 4131 12168
rect 3933 11970 3989 12026
rect 4075 11970 4131 12026
rect 3933 11828 3989 11884
rect 4075 11828 4131 11884
rect 3933 11686 3989 11742
rect 4075 11686 4131 11742
rect 3933 11544 3989 11600
rect 4075 11544 4131 11600
rect 3933 11402 3989 11458
rect 4075 11402 4131 11458
rect 3933 11260 3989 11316
rect 4075 11260 4131 11316
rect 3933 11118 3989 11174
rect 4075 11118 4131 11174
rect 3933 10976 3989 11032
rect 4075 10976 4131 11032
rect 3933 10834 3989 10890
rect 4075 10834 4131 10890
rect 3933 10692 3989 10748
rect 4075 10692 4131 10748
rect 3933 10550 3989 10606
rect 4075 10550 4131 10606
rect 3933 10408 3989 10464
rect 4075 10408 4131 10464
rect 3933 10266 3989 10322
rect 4075 10266 4131 10322
rect 3933 10124 3989 10180
rect 4075 10124 4131 10180
rect 3933 9982 3989 10038
rect 4075 9982 4131 10038
rect 3933 9840 3989 9896
rect 4075 9840 4131 9896
rect 3933 9698 3989 9754
rect 4075 9698 4131 9754
rect 3933 9556 3989 9612
rect 4075 9556 4131 9612
rect 3933 9414 3989 9470
rect 4075 9414 4131 9470
rect 3933 9272 3989 9328
rect 4075 9272 4131 9328
rect 3933 9130 3989 9186
rect 4075 9130 4131 9186
rect 3933 8988 3989 9044
rect 4075 8988 4131 9044
rect 3933 8846 3989 8902
rect 4075 8846 4131 8902
rect 3933 8704 3989 8760
rect 4075 8704 4131 8760
rect 3933 8562 3989 8618
rect 4075 8562 4131 8618
rect 3933 8420 3989 8476
rect 4075 8420 4131 8476
rect 3933 8278 3989 8334
rect 4075 8278 4131 8334
rect 3933 8136 3989 8192
rect 4075 8136 4131 8192
rect 3933 7994 3989 8050
rect 4075 7994 4131 8050
rect 3933 7852 3989 7908
rect 4075 7852 4131 7908
rect 3933 7710 3989 7766
rect 4075 7710 4131 7766
rect 3933 7568 3989 7624
rect 4075 7568 4131 7624
rect 3933 7426 3989 7482
rect 4075 7426 4131 7482
rect 3933 7284 3989 7340
rect 4075 7284 4131 7340
rect 3933 7142 3989 7198
rect 4075 7142 4131 7198
rect 3933 7000 3989 7056
rect 4075 7000 4131 7056
rect 3933 6858 3989 6914
rect 4075 6858 4131 6914
rect 3933 6716 3989 6772
rect 4075 6716 4131 6772
rect 3933 6574 3989 6630
rect 4075 6574 4131 6630
rect 3933 6432 3989 6488
rect 4075 6432 4131 6488
rect 3933 6290 3989 6346
rect 4075 6290 4131 6346
rect 3933 6148 3989 6204
rect 4075 6148 4131 6204
rect 3933 6006 3989 6062
rect 4075 6006 4131 6062
rect 3933 5864 3989 5920
rect 4075 5864 4131 5920
rect 3933 5722 3989 5778
rect 4075 5722 4131 5778
rect 3933 5580 3989 5636
rect 4075 5580 4131 5636
rect 3933 5438 3989 5494
rect 4075 5438 4131 5494
rect 3933 5296 3989 5352
rect 4075 5296 4131 5352
rect 3933 5154 3989 5210
rect 4075 5154 4131 5210
rect 3933 5012 3989 5068
rect 4075 5012 4131 5068
rect 3933 4870 3989 4926
rect 4075 4870 4131 4926
rect 3933 4728 3989 4784
rect 4075 4728 4131 4784
rect 3933 4586 3989 4642
rect 4075 4586 4131 4642
rect 3933 4444 3989 4500
rect 4075 4444 4131 4500
rect 3933 4302 3989 4358
rect 4075 4302 4131 4358
rect 3933 4160 3989 4216
rect 4075 4160 4131 4216
rect 3933 4018 3989 4074
rect 4075 4018 4131 4074
rect 3933 3876 3989 3932
rect 4075 3876 4131 3932
rect 3933 3734 3989 3790
rect 4075 3734 4131 3790
rect 3933 3592 3989 3648
rect 4075 3592 4131 3648
rect 3933 3450 3989 3506
rect 4075 3450 4131 3506
rect 3933 3308 3989 3364
rect 4075 3308 4131 3364
rect 3933 3166 3989 3222
rect 4075 3166 4131 3222
rect 3933 3024 3989 3080
rect 4075 3024 4131 3080
rect 3933 2882 3989 2938
rect 4075 2882 4131 2938
rect 3933 2740 3989 2796
rect 4075 2740 4131 2796
rect 3933 2598 3989 2654
rect 4075 2598 4131 2654
rect 3933 2456 3989 2512
rect 4075 2456 4131 2512
rect 3933 2314 3989 2370
rect 4075 2314 4131 2370
rect 3933 2172 3989 2228
rect 4075 2172 4131 2228
rect 3933 2030 3989 2086
rect 4075 2030 4131 2086
rect 3933 1888 3989 1944
rect 4075 1888 4131 1944
rect 3933 1746 3989 1802
rect 4075 1746 4131 1802
rect 3933 1604 3989 1660
rect 4075 1604 4131 1660
rect 3933 1462 3989 1518
rect 4075 1462 4131 1518
rect 3933 1320 3989 1376
rect 4075 1320 4131 1376
rect 3933 1178 3989 1234
rect 4075 1178 4131 1234
rect 3933 1036 3989 1092
rect 4075 1036 4131 1092
rect 3933 894 3989 950
rect 4075 894 4131 950
rect 3933 752 3989 808
rect 4075 752 4131 808
rect 3933 610 3989 666
rect 4075 610 4131 666
rect 3933 468 3989 524
rect 4075 468 4131 524
rect 4338 12254 4394 12310
rect 4480 12254 4536 12310
rect 4338 12112 4394 12168
rect 4480 12112 4536 12168
rect 4338 11970 4394 12026
rect 4480 11970 4536 12026
rect 4338 11828 4394 11884
rect 4480 11828 4536 11884
rect 4338 11686 4394 11742
rect 4480 11686 4536 11742
rect 4338 11544 4394 11600
rect 4480 11544 4536 11600
rect 4338 11402 4394 11458
rect 4480 11402 4536 11458
rect 4338 11260 4394 11316
rect 4480 11260 4536 11316
rect 4338 11118 4394 11174
rect 4480 11118 4536 11174
rect 4338 10976 4394 11032
rect 4480 10976 4536 11032
rect 4338 10834 4394 10890
rect 4480 10834 4536 10890
rect 4338 10692 4394 10748
rect 4480 10692 4536 10748
rect 4338 10550 4394 10606
rect 4480 10550 4536 10606
rect 4338 10408 4394 10464
rect 4480 10408 4536 10464
rect 4338 10266 4394 10322
rect 4480 10266 4536 10322
rect 4338 10124 4394 10180
rect 4480 10124 4536 10180
rect 4338 9982 4394 10038
rect 4480 9982 4536 10038
rect 4338 9840 4394 9896
rect 4480 9840 4536 9896
rect 4338 9698 4394 9754
rect 4480 9698 4536 9754
rect 4338 9556 4394 9612
rect 4480 9556 4536 9612
rect 4338 9414 4394 9470
rect 4480 9414 4536 9470
rect 4338 9272 4394 9328
rect 4480 9272 4536 9328
rect 4338 9130 4394 9186
rect 4480 9130 4536 9186
rect 4338 8988 4394 9044
rect 4480 8988 4536 9044
rect 4338 8846 4394 8902
rect 4480 8846 4536 8902
rect 4338 8704 4394 8760
rect 4480 8704 4536 8760
rect 4338 8562 4394 8618
rect 4480 8562 4536 8618
rect 4338 8420 4394 8476
rect 4480 8420 4536 8476
rect 4338 8278 4394 8334
rect 4480 8278 4536 8334
rect 4338 8136 4394 8192
rect 4480 8136 4536 8192
rect 4338 7994 4394 8050
rect 4480 7994 4536 8050
rect 4338 7852 4394 7908
rect 4480 7852 4536 7908
rect 4338 7710 4394 7766
rect 4480 7710 4536 7766
rect 4338 7568 4394 7624
rect 4480 7568 4536 7624
rect 4338 7426 4394 7482
rect 4480 7426 4536 7482
rect 4338 7284 4394 7340
rect 4480 7284 4536 7340
rect 4338 7142 4394 7198
rect 4480 7142 4536 7198
rect 4338 7000 4394 7056
rect 4480 7000 4536 7056
rect 4338 6858 4394 6914
rect 4480 6858 4536 6914
rect 4338 6716 4394 6772
rect 4480 6716 4536 6772
rect 4338 6574 4394 6630
rect 4480 6574 4536 6630
rect 4338 6432 4394 6488
rect 4480 6432 4536 6488
rect 4338 6290 4394 6346
rect 4480 6290 4536 6346
rect 4338 6148 4394 6204
rect 4480 6148 4536 6204
rect 4338 6006 4394 6062
rect 4480 6006 4536 6062
rect 4338 5864 4394 5920
rect 4480 5864 4536 5920
rect 4338 5722 4394 5778
rect 4480 5722 4536 5778
rect 4338 5580 4394 5636
rect 4480 5580 4536 5636
rect 4338 5438 4394 5494
rect 4480 5438 4536 5494
rect 4338 5296 4394 5352
rect 4480 5296 4536 5352
rect 4338 5154 4394 5210
rect 4480 5154 4536 5210
rect 4338 5012 4394 5068
rect 4480 5012 4536 5068
rect 4338 4870 4394 4926
rect 4480 4870 4536 4926
rect 4338 4728 4394 4784
rect 4480 4728 4536 4784
rect 4338 4586 4394 4642
rect 4480 4586 4536 4642
rect 4338 4444 4394 4500
rect 4480 4444 4536 4500
rect 4338 4302 4394 4358
rect 4480 4302 4536 4358
rect 4338 4160 4394 4216
rect 4480 4160 4536 4216
rect 4338 4018 4394 4074
rect 4480 4018 4536 4074
rect 4338 3876 4394 3932
rect 4480 3876 4536 3932
rect 4338 3734 4394 3790
rect 4480 3734 4536 3790
rect 4338 3592 4394 3648
rect 4480 3592 4536 3648
rect 4338 3450 4394 3506
rect 4480 3450 4536 3506
rect 4338 3308 4394 3364
rect 4480 3308 4536 3364
rect 4338 3166 4394 3222
rect 4480 3166 4536 3222
rect 4338 3024 4394 3080
rect 4480 3024 4536 3080
rect 4338 2882 4394 2938
rect 4480 2882 4536 2938
rect 4338 2740 4394 2796
rect 4480 2740 4536 2796
rect 4338 2598 4394 2654
rect 4480 2598 4536 2654
rect 4338 2456 4394 2512
rect 4480 2456 4536 2512
rect 4338 2314 4394 2370
rect 4480 2314 4536 2370
rect 4338 2172 4394 2228
rect 4480 2172 4536 2228
rect 4338 2030 4394 2086
rect 4480 2030 4536 2086
rect 4338 1888 4394 1944
rect 4480 1888 4536 1944
rect 4338 1746 4394 1802
rect 4480 1746 4536 1802
rect 4338 1604 4394 1660
rect 4480 1604 4536 1660
rect 4338 1462 4394 1518
rect 4480 1462 4536 1518
rect 4338 1320 4394 1376
rect 4480 1320 4536 1376
rect 4338 1178 4394 1234
rect 4480 1178 4536 1234
rect 4338 1036 4394 1092
rect 4480 1036 4536 1092
rect 4338 894 4394 950
rect 4480 894 4536 950
rect 4338 752 4394 808
rect 4480 752 4536 808
rect 4338 610 4394 666
rect 4480 610 4536 666
rect 4338 468 4394 524
rect 4480 468 4536 524
rect 4738 12254 4794 12310
rect 4880 12254 4936 12310
rect 4738 12112 4794 12168
rect 4880 12112 4936 12168
rect 4738 11970 4794 12026
rect 4880 11970 4936 12026
rect 4738 11828 4794 11884
rect 4880 11828 4936 11884
rect 4738 11686 4794 11742
rect 4880 11686 4936 11742
rect 4738 11544 4794 11600
rect 4880 11544 4936 11600
rect 4738 11402 4794 11458
rect 4880 11402 4936 11458
rect 4738 11260 4794 11316
rect 4880 11260 4936 11316
rect 4738 11118 4794 11174
rect 4880 11118 4936 11174
rect 4738 10976 4794 11032
rect 4880 10976 4936 11032
rect 4738 10834 4794 10890
rect 4880 10834 4936 10890
rect 4738 10692 4794 10748
rect 4880 10692 4936 10748
rect 4738 10550 4794 10606
rect 4880 10550 4936 10606
rect 4738 10408 4794 10464
rect 4880 10408 4936 10464
rect 4738 10266 4794 10322
rect 4880 10266 4936 10322
rect 4738 10124 4794 10180
rect 4880 10124 4936 10180
rect 4738 9982 4794 10038
rect 4880 9982 4936 10038
rect 4738 9840 4794 9896
rect 4880 9840 4936 9896
rect 4738 9698 4794 9754
rect 4880 9698 4936 9754
rect 4738 9556 4794 9612
rect 4880 9556 4936 9612
rect 4738 9414 4794 9470
rect 4880 9414 4936 9470
rect 4738 9272 4794 9328
rect 4880 9272 4936 9328
rect 4738 9130 4794 9186
rect 4880 9130 4936 9186
rect 4738 8988 4794 9044
rect 4880 8988 4936 9044
rect 4738 8846 4794 8902
rect 4880 8846 4936 8902
rect 4738 8704 4794 8760
rect 4880 8704 4936 8760
rect 4738 8562 4794 8618
rect 4880 8562 4936 8618
rect 4738 8420 4794 8476
rect 4880 8420 4936 8476
rect 4738 8278 4794 8334
rect 4880 8278 4936 8334
rect 4738 8136 4794 8192
rect 4880 8136 4936 8192
rect 4738 7994 4794 8050
rect 4880 7994 4936 8050
rect 4738 7852 4794 7908
rect 4880 7852 4936 7908
rect 4738 7710 4794 7766
rect 4880 7710 4936 7766
rect 4738 7568 4794 7624
rect 4880 7568 4936 7624
rect 4738 7426 4794 7482
rect 4880 7426 4936 7482
rect 4738 7284 4794 7340
rect 4880 7284 4936 7340
rect 4738 7142 4794 7198
rect 4880 7142 4936 7198
rect 4738 7000 4794 7056
rect 4880 7000 4936 7056
rect 4738 6858 4794 6914
rect 4880 6858 4936 6914
rect 4738 6716 4794 6772
rect 4880 6716 4936 6772
rect 4738 6574 4794 6630
rect 4880 6574 4936 6630
rect 4738 6432 4794 6488
rect 4880 6432 4936 6488
rect 4738 6290 4794 6346
rect 4880 6290 4936 6346
rect 4738 6148 4794 6204
rect 4880 6148 4936 6204
rect 4738 6006 4794 6062
rect 4880 6006 4936 6062
rect 4738 5864 4794 5920
rect 4880 5864 4936 5920
rect 4738 5722 4794 5778
rect 4880 5722 4936 5778
rect 4738 5580 4794 5636
rect 4880 5580 4936 5636
rect 4738 5438 4794 5494
rect 4880 5438 4936 5494
rect 4738 5296 4794 5352
rect 4880 5296 4936 5352
rect 4738 5154 4794 5210
rect 4880 5154 4936 5210
rect 4738 5012 4794 5068
rect 4880 5012 4936 5068
rect 4738 4870 4794 4926
rect 4880 4870 4936 4926
rect 4738 4728 4794 4784
rect 4880 4728 4936 4784
rect 4738 4586 4794 4642
rect 4880 4586 4936 4642
rect 4738 4444 4794 4500
rect 4880 4444 4936 4500
rect 4738 4302 4794 4358
rect 4880 4302 4936 4358
rect 4738 4160 4794 4216
rect 4880 4160 4936 4216
rect 4738 4018 4794 4074
rect 4880 4018 4936 4074
rect 4738 3876 4794 3932
rect 4880 3876 4936 3932
rect 4738 3734 4794 3790
rect 4880 3734 4936 3790
rect 4738 3592 4794 3648
rect 4880 3592 4936 3648
rect 4738 3450 4794 3506
rect 4880 3450 4936 3506
rect 4738 3308 4794 3364
rect 4880 3308 4936 3364
rect 4738 3166 4794 3222
rect 4880 3166 4936 3222
rect 4738 3024 4794 3080
rect 4880 3024 4936 3080
rect 4738 2882 4794 2938
rect 4880 2882 4936 2938
rect 4738 2740 4794 2796
rect 4880 2740 4936 2796
rect 4738 2598 4794 2654
rect 4880 2598 4936 2654
rect 4738 2456 4794 2512
rect 4880 2456 4936 2512
rect 4738 2314 4794 2370
rect 4880 2314 4936 2370
rect 4738 2172 4794 2228
rect 4880 2172 4936 2228
rect 4738 2030 4794 2086
rect 4880 2030 4936 2086
rect 4738 1888 4794 1944
rect 4880 1888 4936 1944
rect 4738 1746 4794 1802
rect 4880 1746 4936 1802
rect 4738 1604 4794 1660
rect 4880 1604 4936 1660
rect 4738 1462 4794 1518
rect 4880 1462 4936 1518
rect 4738 1320 4794 1376
rect 4880 1320 4936 1376
rect 4738 1178 4794 1234
rect 4880 1178 4936 1234
rect 4738 1036 4794 1092
rect 4880 1036 4936 1092
rect 4738 894 4794 950
rect 4880 894 4936 950
rect 4738 752 4794 808
rect 4880 752 4936 808
rect 4738 610 4794 666
rect 4880 610 4936 666
rect 4738 468 4794 524
rect 4880 468 4936 524
rect 5143 12254 5199 12310
rect 5285 12254 5341 12310
rect 5143 12112 5199 12168
rect 5285 12112 5341 12168
rect 5143 11970 5199 12026
rect 5285 11970 5341 12026
rect 5143 11828 5199 11884
rect 5285 11828 5341 11884
rect 5143 11686 5199 11742
rect 5285 11686 5341 11742
rect 5143 11544 5199 11600
rect 5285 11544 5341 11600
rect 5143 11402 5199 11458
rect 5285 11402 5341 11458
rect 5143 11260 5199 11316
rect 5285 11260 5341 11316
rect 5143 11118 5199 11174
rect 5285 11118 5341 11174
rect 5143 10976 5199 11032
rect 5285 10976 5341 11032
rect 5143 10834 5199 10890
rect 5285 10834 5341 10890
rect 5143 10692 5199 10748
rect 5285 10692 5341 10748
rect 5143 10550 5199 10606
rect 5285 10550 5341 10606
rect 5143 10408 5199 10464
rect 5285 10408 5341 10464
rect 5143 10266 5199 10322
rect 5285 10266 5341 10322
rect 5143 10124 5199 10180
rect 5285 10124 5341 10180
rect 5143 9982 5199 10038
rect 5285 9982 5341 10038
rect 5143 9840 5199 9896
rect 5285 9840 5341 9896
rect 5143 9698 5199 9754
rect 5285 9698 5341 9754
rect 5143 9556 5199 9612
rect 5285 9556 5341 9612
rect 5143 9414 5199 9470
rect 5285 9414 5341 9470
rect 5143 9272 5199 9328
rect 5285 9272 5341 9328
rect 5143 9130 5199 9186
rect 5285 9130 5341 9186
rect 5143 8988 5199 9044
rect 5285 8988 5341 9044
rect 5143 8846 5199 8902
rect 5285 8846 5341 8902
rect 5143 8704 5199 8760
rect 5285 8704 5341 8760
rect 5143 8562 5199 8618
rect 5285 8562 5341 8618
rect 5143 8420 5199 8476
rect 5285 8420 5341 8476
rect 5143 8278 5199 8334
rect 5285 8278 5341 8334
rect 5143 8136 5199 8192
rect 5285 8136 5341 8192
rect 5143 7994 5199 8050
rect 5285 7994 5341 8050
rect 5143 7852 5199 7908
rect 5285 7852 5341 7908
rect 5143 7710 5199 7766
rect 5285 7710 5341 7766
rect 5143 7568 5199 7624
rect 5285 7568 5341 7624
rect 5143 7426 5199 7482
rect 5285 7426 5341 7482
rect 5143 7284 5199 7340
rect 5285 7284 5341 7340
rect 5143 7142 5199 7198
rect 5285 7142 5341 7198
rect 5143 7000 5199 7056
rect 5285 7000 5341 7056
rect 5143 6858 5199 6914
rect 5285 6858 5341 6914
rect 5143 6716 5199 6772
rect 5285 6716 5341 6772
rect 5143 6574 5199 6630
rect 5285 6574 5341 6630
rect 5143 6432 5199 6488
rect 5285 6432 5341 6488
rect 5143 6290 5199 6346
rect 5285 6290 5341 6346
rect 5143 6148 5199 6204
rect 5285 6148 5341 6204
rect 5143 6006 5199 6062
rect 5285 6006 5341 6062
rect 5143 5864 5199 5920
rect 5285 5864 5341 5920
rect 5143 5722 5199 5778
rect 5285 5722 5341 5778
rect 5143 5580 5199 5636
rect 5285 5580 5341 5636
rect 5143 5438 5199 5494
rect 5285 5438 5341 5494
rect 5143 5296 5199 5352
rect 5285 5296 5341 5352
rect 5143 5154 5199 5210
rect 5285 5154 5341 5210
rect 5143 5012 5199 5068
rect 5285 5012 5341 5068
rect 5143 4870 5199 4926
rect 5285 4870 5341 4926
rect 5143 4728 5199 4784
rect 5285 4728 5341 4784
rect 5143 4586 5199 4642
rect 5285 4586 5341 4642
rect 5143 4444 5199 4500
rect 5285 4444 5341 4500
rect 5143 4302 5199 4358
rect 5285 4302 5341 4358
rect 5143 4160 5199 4216
rect 5285 4160 5341 4216
rect 5143 4018 5199 4074
rect 5285 4018 5341 4074
rect 5143 3876 5199 3932
rect 5285 3876 5341 3932
rect 5143 3734 5199 3790
rect 5285 3734 5341 3790
rect 5143 3592 5199 3648
rect 5285 3592 5341 3648
rect 5143 3450 5199 3506
rect 5285 3450 5341 3506
rect 5143 3308 5199 3364
rect 5285 3308 5341 3364
rect 5143 3166 5199 3222
rect 5285 3166 5341 3222
rect 5143 3024 5199 3080
rect 5285 3024 5341 3080
rect 5143 2882 5199 2938
rect 5285 2882 5341 2938
rect 5143 2740 5199 2796
rect 5285 2740 5341 2796
rect 5143 2598 5199 2654
rect 5285 2598 5341 2654
rect 5143 2456 5199 2512
rect 5285 2456 5341 2512
rect 5143 2314 5199 2370
rect 5285 2314 5341 2370
rect 5143 2172 5199 2228
rect 5285 2172 5341 2228
rect 5143 2030 5199 2086
rect 5285 2030 5341 2086
rect 5143 1888 5199 1944
rect 5285 1888 5341 1944
rect 5143 1746 5199 1802
rect 5285 1746 5341 1802
rect 5143 1604 5199 1660
rect 5285 1604 5341 1660
rect 5143 1462 5199 1518
rect 5285 1462 5341 1518
rect 5143 1320 5199 1376
rect 5285 1320 5341 1376
rect 5143 1178 5199 1234
rect 5285 1178 5341 1234
rect 5143 1036 5199 1092
rect 5285 1036 5341 1092
rect 5143 894 5199 950
rect 5285 894 5341 950
rect 5143 752 5199 808
rect 5285 752 5341 808
rect 5143 610 5199 666
rect 5285 610 5341 666
rect 5143 468 5199 524
rect 5285 468 5341 524
rect 5540 12254 5596 12310
rect 5682 12254 5738 12310
rect 5540 12112 5596 12168
rect 5682 12112 5738 12168
rect 5540 11970 5596 12026
rect 5682 11970 5738 12026
rect 5540 11828 5596 11884
rect 5682 11828 5738 11884
rect 5540 11686 5596 11742
rect 5682 11686 5738 11742
rect 5540 11544 5596 11600
rect 5682 11544 5738 11600
rect 5540 11402 5596 11458
rect 5682 11402 5738 11458
rect 5540 11260 5596 11316
rect 5682 11260 5738 11316
rect 5540 11118 5596 11174
rect 5682 11118 5738 11174
rect 5540 10976 5596 11032
rect 5682 10976 5738 11032
rect 5540 10834 5596 10890
rect 5682 10834 5738 10890
rect 5540 10692 5596 10748
rect 5682 10692 5738 10748
rect 5540 10550 5596 10606
rect 5682 10550 5738 10606
rect 5540 10408 5596 10464
rect 5682 10408 5738 10464
rect 5540 10266 5596 10322
rect 5682 10266 5738 10322
rect 5540 10124 5596 10180
rect 5682 10124 5738 10180
rect 5540 9982 5596 10038
rect 5682 9982 5738 10038
rect 5540 9840 5596 9896
rect 5682 9840 5738 9896
rect 5540 9698 5596 9754
rect 5682 9698 5738 9754
rect 5540 9556 5596 9612
rect 5682 9556 5738 9612
rect 5540 9414 5596 9470
rect 5682 9414 5738 9470
rect 5540 9272 5596 9328
rect 5682 9272 5738 9328
rect 5540 9130 5596 9186
rect 5682 9130 5738 9186
rect 5540 8988 5596 9044
rect 5682 8988 5738 9044
rect 5540 8846 5596 8902
rect 5682 8846 5738 8902
rect 5540 8704 5596 8760
rect 5682 8704 5738 8760
rect 5540 8562 5596 8618
rect 5682 8562 5738 8618
rect 5540 8420 5596 8476
rect 5682 8420 5738 8476
rect 5540 8278 5596 8334
rect 5682 8278 5738 8334
rect 5540 8136 5596 8192
rect 5682 8136 5738 8192
rect 5540 7994 5596 8050
rect 5682 7994 5738 8050
rect 5540 7852 5596 7908
rect 5682 7852 5738 7908
rect 5540 7710 5596 7766
rect 5682 7710 5738 7766
rect 5540 7568 5596 7624
rect 5682 7568 5738 7624
rect 5540 7426 5596 7482
rect 5682 7426 5738 7482
rect 5540 7284 5596 7340
rect 5682 7284 5738 7340
rect 5540 7142 5596 7198
rect 5682 7142 5738 7198
rect 5540 7000 5596 7056
rect 5682 7000 5738 7056
rect 5540 6858 5596 6914
rect 5682 6858 5738 6914
rect 5540 6716 5596 6772
rect 5682 6716 5738 6772
rect 5540 6574 5596 6630
rect 5682 6574 5738 6630
rect 5540 6432 5596 6488
rect 5682 6432 5738 6488
rect 5540 6290 5596 6346
rect 5682 6290 5738 6346
rect 5540 6148 5596 6204
rect 5682 6148 5738 6204
rect 5540 6006 5596 6062
rect 5682 6006 5738 6062
rect 5540 5864 5596 5920
rect 5682 5864 5738 5920
rect 5540 5722 5596 5778
rect 5682 5722 5738 5778
rect 5540 5580 5596 5636
rect 5682 5580 5738 5636
rect 5540 5438 5596 5494
rect 5682 5438 5738 5494
rect 5540 5296 5596 5352
rect 5682 5296 5738 5352
rect 5540 5154 5596 5210
rect 5682 5154 5738 5210
rect 5540 5012 5596 5068
rect 5682 5012 5738 5068
rect 5540 4870 5596 4926
rect 5682 4870 5738 4926
rect 5540 4728 5596 4784
rect 5682 4728 5738 4784
rect 5540 4586 5596 4642
rect 5682 4586 5738 4642
rect 5540 4444 5596 4500
rect 5682 4444 5738 4500
rect 5540 4302 5596 4358
rect 5682 4302 5738 4358
rect 5540 4160 5596 4216
rect 5682 4160 5738 4216
rect 5540 4018 5596 4074
rect 5682 4018 5738 4074
rect 5540 3876 5596 3932
rect 5682 3876 5738 3932
rect 5540 3734 5596 3790
rect 5682 3734 5738 3790
rect 5540 3592 5596 3648
rect 5682 3592 5738 3648
rect 5540 3450 5596 3506
rect 5682 3450 5738 3506
rect 5540 3308 5596 3364
rect 5682 3308 5738 3364
rect 5540 3166 5596 3222
rect 5682 3166 5738 3222
rect 5540 3024 5596 3080
rect 5682 3024 5738 3080
rect 5540 2882 5596 2938
rect 5682 2882 5738 2938
rect 5540 2740 5596 2796
rect 5682 2740 5738 2796
rect 5540 2598 5596 2654
rect 5682 2598 5738 2654
rect 5540 2456 5596 2512
rect 5682 2456 5738 2512
rect 5540 2314 5596 2370
rect 5682 2314 5738 2370
rect 5540 2172 5596 2228
rect 5682 2172 5738 2228
rect 5540 2030 5596 2086
rect 5682 2030 5738 2086
rect 5540 1888 5596 1944
rect 5682 1888 5738 1944
rect 5540 1746 5596 1802
rect 5682 1746 5738 1802
rect 5540 1604 5596 1660
rect 5682 1604 5738 1660
rect 5540 1462 5596 1518
rect 5682 1462 5738 1518
rect 5540 1320 5596 1376
rect 5682 1320 5738 1376
rect 5540 1178 5596 1234
rect 5682 1178 5738 1234
rect 5540 1036 5596 1092
rect 5682 1036 5738 1092
rect 5540 894 5596 950
rect 5682 894 5738 950
rect 5540 752 5596 808
rect 5682 752 5738 808
rect 5540 610 5596 666
rect 5682 610 5738 666
rect 5540 468 5596 524
rect 5682 468 5738 524
rect 5937 12254 5993 12310
rect 6079 12254 6135 12310
rect 5937 12112 5993 12168
rect 6079 12112 6135 12168
rect 5937 11970 5993 12026
rect 6079 11970 6135 12026
rect 5937 11828 5993 11884
rect 6079 11828 6135 11884
rect 5937 11686 5993 11742
rect 6079 11686 6135 11742
rect 5937 11544 5993 11600
rect 6079 11544 6135 11600
rect 5937 11402 5993 11458
rect 6079 11402 6135 11458
rect 5937 11260 5993 11316
rect 6079 11260 6135 11316
rect 5937 11118 5993 11174
rect 6079 11118 6135 11174
rect 5937 10976 5993 11032
rect 6079 10976 6135 11032
rect 5937 10834 5993 10890
rect 6079 10834 6135 10890
rect 5937 10692 5993 10748
rect 6079 10692 6135 10748
rect 5937 10550 5993 10606
rect 6079 10550 6135 10606
rect 5937 10408 5993 10464
rect 6079 10408 6135 10464
rect 5937 10266 5993 10322
rect 6079 10266 6135 10322
rect 5937 10124 5993 10180
rect 6079 10124 6135 10180
rect 5937 9982 5993 10038
rect 6079 9982 6135 10038
rect 5937 9840 5993 9896
rect 6079 9840 6135 9896
rect 5937 9698 5993 9754
rect 6079 9698 6135 9754
rect 5937 9556 5993 9612
rect 6079 9556 6135 9612
rect 5937 9414 5993 9470
rect 6079 9414 6135 9470
rect 5937 9272 5993 9328
rect 6079 9272 6135 9328
rect 5937 9130 5993 9186
rect 6079 9130 6135 9186
rect 5937 8988 5993 9044
rect 6079 8988 6135 9044
rect 5937 8846 5993 8902
rect 6079 8846 6135 8902
rect 5937 8704 5993 8760
rect 6079 8704 6135 8760
rect 5937 8562 5993 8618
rect 6079 8562 6135 8618
rect 5937 8420 5993 8476
rect 6079 8420 6135 8476
rect 5937 8278 5993 8334
rect 6079 8278 6135 8334
rect 5937 8136 5993 8192
rect 6079 8136 6135 8192
rect 5937 7994 5993 8050
rect 6079 7994 6135 8050
rect 5937 7852 5993 7908
rect 6079 7852 6135 7908
rect 5937 7710 5993 7766
rect 6079 7710 6135 7766
rect 5937 7568 5993 7624
rect 6079 7568 6135 7624
rect 5937 7426 5993 7482
rect 6079 7426 6135 7482
rect 5937 7284 5993 7340
rect 6079 7284 6135 7340
rect 5937 7142 5993 7198
rect 6079 7142 6135 7198
rect 5937 7000 5993 7056
rect 6079 7000 6135 7056
rect 5937 6858 5993 6914
rect 6079 6858 6135 6914
rect 5937 6716 5993 6772
rect 6079 6716 6135 6772
rect 5937 6574 5993 6630
rect 6079 6574 6135 6630
rect 5937 6432 5993 6488
rect 6079 6432 6135 6488
rect 5937 6290 5993 6346
rect 6079 6290 6135 6346
rect 5937 6148 5993 6204
rect 6079 6148 6135 6204
rect 5937 6006 5993 6062
rect 6079 6006 6135 6062
rect 5937 5864 5993 5920
rect 6079 5864 6135 5920
rect 5937 5722 5993 5778
rect 6079 5722 6135 5778
rect 5937 5580 5993 5636
rect 6079 5580 6135 5636
rect 5937 5438 5993 5494
rect 6079 5438 6135 5494
rect 5937 5296 5993 5352
rect 6079 5296 6135 5352
rect 5937 5154 5993 5210
rect 6079 5154 6135 5210
rect 5937 5012 5993 5068
rect 6079 5012 6135 5068
rect 5937 4870 5993 4926
rect 6079 4870 6135 4926
rect 5937 4728 5993 4784
rect 6079 4728 6135 4784
rect 5937 4586 5993 4642
rect 6079 4586 6135 4642
rect 5937 4444 5993 4500
rect 6079 4444 6135 4500
rect 5937 4302 5993 4358
rect 6079 4302 6135 4358
rect 5937 4160 5993 4216
rect 6079 4160 6135 4216
rect 5937 4018 5993 4074
rect 6079 4018 6135 4074
rect 5937 3876 5993 3932
rect 6079 3876 6135 3932
rect 5937 3734 5993 3790
rect 6079 3734 6135 3790
rect 5937 3592 5993 3648
rect 6079 3592 6135 3648
rect 5937 3450 5993 3506
rect 6079 3450 6135 3506
rect 5937 3308 5993 3364
rect 6079 3308 6135 3364
rect 5937 3166 5993 3222
rect 6079 3166 6135 3222
rect 5937 3024 5993 3080
rect 6079 3024 6135 3080
rect 5937 2882 5993 2938
rect 6079 2882 6135 2938
rect 5937 2740 5993 2796
rect 6079 2740 6135 2796
rect 5937 2598 5993 2654
rect 6079 2598 6135 2654
rect 5937 2456 5993 2512
rect 6079 2456 6135 2512
rect 5937 2314 5993 2370
rect 6079 2314 6135 2370
rect 5937 2172 5993 2228
rect 6079 2172 6135 2228
rect 5937 2030 5993 2086
rect 6079 2030 6135 2086
rect 5937 1888 5993 1944
rect 6079 1888 6135 1944
rect 5937 1746 5993 1802
rect 6079 1746 6135 1802
rect 5937 1604 5993 1660
rect 6079 1604 6135 1660
rect 5937 1462 5993 1518
rect 6079 1462 6135 1518
rect 5937 1320 5993 1376
rect 6079 1320 6135 1376
rect 5937 1178 5993 1234
rect 6079 1178 6135 1234
rect 5937 1036 5993 1092
rect 6079 1036 6135 1092
rect 5937 894 5993 950
rect 6079 894 6135 950
rect 5937 752 5993 808
rect 6079 752 6135 808
rect 5937 610 5993 666
rect 6079 610 6135 666
rect 5937 468 5993 524
rect 6079 468 6135 524
rect 6340 12254 6396 12310
rect 6482 12254 6538 12310
rect 6340 12112 6396 12168
rect 6482 12112 6538 12168
rect 6340 11970 6396 12026
rect 6482 11970 6538 12026
rect 6340 11828 6396 11884
rect 6482 11828 6538 11884
rect 6340 11686 6396 11742
rect 6482 11686 6538 11742
rect 6340 11544 6396 11600
rect 6482 11544 6538 11600
rect 6340 11402 6396 11458
rect 6482 11402 6538 11458
rect 6340 11260 6396 11316
rect 6482 11260 6538 11316
rect 6340 11118 6396 11174
rect 6482 11118 6538 11174
rect 6340 10976 6396 11032
rect 6482 10976 6538 11032
rect 6340 10834 6396 10890
rect 6482 10834 6538 10890
rect 6340 10692 6396 10748
rect 6482 10692 6538 10748
rect 6340 10550 6396 10606
rect 6482 10550 6538 10606
rect 6340 10408 6396 10464
rect 6482 10408 6538 10464
rect 6340 10266 6396 10322
rect 6482 10266 6538 10322
rect 6340 10124 6396 10180
rect 6482 10124 6538 10180
rect 6340 9982 6396 10038
rect 6482 9982 6538 10038
rect 6340 9840 6396 9896
rect 6482 9840 6538 9896
rect 6340 9698 6396 9754
rect 6482 9698 6538 9754
rect 6340 9556 6396 9612
rect 6482 9556 6538 9612
rect 6340 9414 6396 9470
rect 6482 9414 6538 9470
rect 6340 9272 6396 9328
rect 6482 9272 6538 9328
rect 6340 9130 6396 9186
rect 6482 9130 6538 9186
rect 6340 8988 6396 9044
rect 6482 8988 6538 9044
rect 6340 8846 6396 8902
rect 6482 8846 6538 8902
rect 6340 8704 6396 8760
rect 6482 8704 6538 8760
rect 6340 8562 6396 8618
rect 6482 8562 6538 8618
rect 6340 8420 6396 8476
rect 6482 8420 6538 8476
rect 6340 8278 6396 8334
rect 6482 8278 6538 8334
rect 6340 8136 6396 8192
rect 6482 8136 6538 8192
rect 6340 7994 6396 8050
rect 6482 7994 6538 8050
rect 6340 7852 6396 7908
rect 6482 7852 6538 7908
rect 6340 7710 6396 7766
rect 6482 7710 6538 7766
rect 6340 7568 6396 7624
rect 6482 7568 6538 7624
rect 6340 7426 6396 7482
rect 6482 7426 6538 7482
rect 6340 7284 6396 7340
rect 6482 7284 6538 7340
rect 6340 7142 6396 7198
rect 6482 7142 6538 7198
rect 6340 7000 6396 7056
rect 6482 7000 6538 7056
rect 6340 6858 6396 6914
rect 6482 6858 6538 6914
rect 6340 6716 6396 6772
rect 6482 6716 6538 6772
rect 6340 6574 6396 6630
rect 6482 6574 6538 6630
rect 6340 6432 6396 6488
rect 6482 6432 6538 6488
rect 6340 6290 6396 6346
rect 6482 6290 6538 6346
rect 6340 6148 6396 6204
rect 6482 6148 6538 6204
rect 6340 6006 6396 6062
rect 6482 6006 6538 6062
rect 6340 5864 6396 5920
rect 6482 5864 6538 5920
rect 6340 5722 6396 5778
rect 6482 5722 6538 5778
rect 6340 5580 6396 5636
rect 6482 5580 6538 5636
rect 6340 5438 6396 5494
rect 6482 5438 6538 5494
rect 6340 5296 6396 5352
rect 6482 5296 6538 5352
rect 6340 5154 6396 5210
rect 6482 5154 6538 5210
rect 6340 5012 6396 5068
rect 6482 5012 6538 5068
rect 6340 4870 6396 4926
rect 6482 4870 6538 4926
rect 6340 4728 6396 4784
rect 6482 4728 6538 4784
rect 6340 4586 6396 4642
rect 6482 4586 6538 4642
rect 6340 4444 6396 4500
rect 6482 4444 6538 4500
rect 6340 4302 6396 4358
rect 6482 4302 6538 4358
rect 6340 4160 6396 4216
rect 6482 4160 6538 4216
rect 6340 4018 6396 4074
rect 6482 4018 6538 4074
rect 6340 3876 6396 3932
rect 6482 3876 6538 3932
rect 6340 3734 6396 3790
rect 6482 3734 6538 3790
rect 6340 3592 6396 3648
rect 6482 3592 6538 3648
rect 6340 3450 6396 3506
rect 6482 3450 6538 3506
rect 6340 3308 6396 3364
rect 6482 3308 6538 3364
rect 6340 3166 6396 3222
rect 6482 3166 6538 3222
rect 6340 3024 6396 3080
rect 6482 3024 6538 3080
rect 6340 2882 6396 2938
rect 6482 2882 6538 2938
rect 6340 2740 6396 2796
rect 6482 2740 6538 2796
rect 6340 2598 6396 2654
rect 6482 2598 6538 2654
rect 6340 2456 6396 2512
rect 6482 2456 6538 2512
rect 6340 2314 6396 2370
rect 6482 2314 6538 2370
rect 6340 2172 6396 2228
rect 6482 2172 6538 2228
rect 6340 2030 6396 2086
rect 6482 2030 6538 2086
rect 6340 1888 6396 1944
rect 6482 1888 6538 1944
rect 6340 1746 6396 1802
rect 6482 1746 6538 1802
rect 6340 1604 6396 1660
rect 6482 1604 6538 1660
rect 6340 1462 6396 1518
rect 6482 1462 6538 1518
rect 6340 1320 6396 1376
rect 6482 1320 6538 1376
rect 6340 1178 6396 1234
rect 6482 1178 6538 1234
rect 6340 1036 6396 1092
rect 6482 1036 6538 1092
rect 6340 894 6396 950
rect 6482 894 6538 950
rect 6340 752 6396 808
rect 6482 752 6538 808
rect 6340 610 6396 666
rect 6482 610 6538 666
rect 6340 468 6396 524
rect 6482 468 6538 524
rect 6742 12254 6798 12310
rect 6884 12254 6940 12310
rect 6742 12112 6798 12168
rect 6884 12112 6940 12168
rect 6742 11970 6798 12026
rect 6884 11970 6940 12026
rect 6742 11828 6798 11884
rect 6884 11828 6940 11884
rect 6742 11686 6798 11742
rect 6884 11686 6940 11742
rect 6742 11544 6798 11600
rect 6884 11544 6940 11600
rect 6742 11402 6798 11458
rect 6884 11402 6940 11458
rect 6742 11260 6798 11316
rect 6884 11260 6940 11316
rect 6742 11118 6798 11174
rect 6884 11118 6940 11174
rect 6742 10976 6798 11032
rect 6884 10976 6940 11032
rect 6742 10834 6798 10890
rect 6884 10834 6940 10890
rect 6742 10692 6798 10748
rect 6884 10692 6940 10748
rect 6742 10550 6798 10606
rect 6884 10550 6940 10606
rect 6742 10408 6798 10464
rect 6884 10408 6940 10464
rect 6742 10266 6798 10322
rect 6884 10266 6940 10322
rect 6742 10124 6798 10180
rect 6884 10124 6940 10180
rect 6742 9982 6798 10038
rect 6884 9982 6940 10038
rect 6742 9840 6798 9896
rect 6884 9840 6940 9896
rect 6742 9698 6798 9754
rect 6884 9698 6940 9754
rect 6742 9556 6798 9612
rect 6884 9556 6940 9612
rect 6742 9414 6798 9470
rect 6884 9414 6940 9470
rect 6742 9272 6798 9328
rect 6884 9272 6940 9328
rect 6742 9130 6798 9186
rect 6884 9130 6940 9186
rect 6742 8988 6798 9044
rect 6884 8988 6940 9044
rect 6742 8846 6798 8902
rect 6884 8846 6940 8902
rect 6742 8704 6798 8760
rect 6884 8704 6940 8760
rect 6742 8562 6798 8618
rect 6884 8562 6940 8618
rect 6742 8420 6798 8476
rect 6884 8420 6940 8476
rect 6742 8278 6798 8334
rect 6884 8278 6940 8334
rect 6742 8136 6798 8192
rect 6884 8136 6940 8192
rect 6742 7994 6798 8050
rect 6884 7994 6940 8050
rect 6742 7852 6798 7908
rect 6884 7852 6940 7908
rect 6742 7710 6798 7766
rect 6884 7710 6940 7766
rect 6742 7568 6798 7624
rect 6884 7568 6940 7624
rect 6742 7426 6798 7482
rect 6884 7426 6940 7482
rect 6742 7284 6798 7340
rect 6884 7284 6940 7340
rect 6742 7142 6798 7198
rect 6884 7142 6940 7198
rect 6742 7000 6798 7056
rect 6884 7000 6940 7056
rect 6742 6858 6798 6914
rect 6884 6858 6940 6914
rect 6742 6716 6798 6772
rect 6884 6716 6940 6772
rect 6742 6574 6798 6630
rect 6884 6574 6940 6630
rect 6742 6432 6798 6488
rect 6884 6432 6940 6488
rect 6742 6290 6798 6346
rect 6884 6290 6940 6346
rect 6742 6148 6798 6204
rect 6884 6148 6940 6204
rect 6742 6006 6798 6062
rect 6884 6006 6940 6062
rect 6742 5864 6798 5920
rect 6884 5864 6940 5920
rect 6742 5722 6798 5778
rect 6884 5722 6940 5778
rect 6742 5580 6798 5636
rect 6884 5580 6940 5636
rect 6742 5438 6798 5494
rect 6884 5438 6940 5494
rect 6742 5296 6798 5352
rect 6884 5296 6940 5352
rect 6742 5154 6798 5210
rect 6884 5154 6940 5210
rect 6742 5012 6798 5068
rect 6884 5012 6940 5068
rect 6742 4870 6798 4926
rect 6884 4870 6940 4926
rect 6742 4728 6798 4784
rect 6884 4728 6940 4784
rect 6742 4586 6798 4642
rect 6884 4586 6940 4642
rect 6742 4444 6798 4500
rect 6884 4444 6940 4500
rect 6742 4302 6798 4358
rect 6884 4302 6940 4358
rect 6742 4160 6798 4216
rect 6884 4160 6940 4216
rect 6742 4018 6798 4074
rect 6884 4018 6940 4074
rect 6742 3876 6798 3932
rect 6884 3876 6940 3932
rect 6742 3734 6798 3790
rect 6884 3734 6940 3790
rect 6742 3592 6798 3648
rect 6884 3592 6940 3648
rect 6742 3450 6798 3506
rect 6884 3450 6940 3506
rect 6742 3308 6798 3364
rect 6884 3308 6940 3364
rect 6742 3166 6798 3222
rect 6884 3166 6940 3222
rect 6742 3024 6798 3080
rect 6884 3024 6940 3080
rect 6742 2882 6798 2938
rect 6884 2882 6940 2938
rect 6742 2740 6798 2796
rect 6884 2740 6940 2796
rect 6742 2598 6798 2654
rect 6884 2598 6940 2654
rect 6742 2456 6798 2512
rect 6884 2456 6940 2512
rect 6742 2314 6798 2370
rect 6884 2314 6940 2370
rect 6742 2172 6798 2228
rect 6884 2172 6940 2228
rect 6742 2030 6798 2086
rect 6884 2030 6940 2086
rect 6742 1888 6798 1944
rect 6884 1888 6940 1944
rect 6742 1746 6798 1802
rect 6884 1746 6940 1802
rect 6742 1604 6798 1660
rect 6884 1604 6940 1660
rect 6742 1462 6798 1518
rect 6884 1462 6940 1518
rect 6742 1320 6798 1376
rect 6884 1320 6940 1376
rect 6742 1178 6798 1234
rect 6884 1178 6940 1234
rect 6742 1036 6798 1092
rect 6884 1036 6940 1092
rect 6742 894 6798 950
rect 6884 894 6940 950
rect 6742 752 6798 808
rect 6884 752 6940 808
rect 6742 610 6798 666
rect 6884 610 6940 666
rect 6742 468 6798 524
rect 6884 468 6940 524
rect 7145 12254 7201 12310
rect 7287 12254 7343 12310
rect 7145 12112 7201 12168
rect 7287 12112 7343 12168
rect 7145 11970 7201 12026
rect 7287 11970 7343 12026
rect 7145 11828 7201 11884
rect 7287 11828 7343 11884
rect 7145 11686 7201 11742
rect 7287 11686 7343 11742
rect 7145 11544 7201 11600
rect 7287 11544 7343 11600
rect 7145 11402 7201 11458
rect 7287 11402 7343 11458
rect 7145 11260 7201 11316
rect 7287 11260 7343 11316
rect 7145 11118 7201 11174
rect 7287 11118 7343 11174
rect 7145 10976 7201 11032
rect 7287 10976 7343 11032
rect 7145 10834 7201 10890
rect 7287 10834 7343 10890
rect 7145 10692 7201 10748
rect 7287 10692 7343 10748
rect 7145 10550 7201 10606
rect 7287 10550 7343 10606
rect 7145 10408 7201 10464
rect 7287 10408 7343 10464
rect 7145 10266 7201 10322
rect 7287 10266 7343 10322
rect 7145 10124 7201 10180
rect 7287 10124 7343 10180
rect 7145 9982 7201 10038
rect 7287 9982 7343 10038
rect 7145 9840 7201 9896
rect 7287 9840 7343 9896
rect 7145 9698 7201 9754
rect 7287 9698 7343 9754
rect 7145 9556 7201 9612
rect 7287 9556 7343 9612
rect 7145 9414 7201 9470
rect 7287 9414 7343 9470
rect 7145 9272 7201 9328
rect 7287 9272 7343 9328
rect 7145 9130 7201 9186
rect 7287 9130 7343 9186
rect 7145 8988 7201 9044
rect 7287 8988 7343 9044
rect 7145 8846 7201 8902
rect 7287 8846 7343 8902
rect 7145 8704 7201 8760
rect 7287 8704 7343 8760
rect 7145 8562 7201 8618
rect 7287 8562 7343 8618
rect 7145 8420 7201 8476
rect 7287 8420 7343 8476
rect 7145 8278 7201 8334
rect 7287 8278 7343 8334
rect 7145 8136 7201 8192
rect 7287 8136 7343 8192
rect 7145 7994 7201 8050
rect 7287 7994 7343 8050
rect 7145 7852 7201 7908
rect 7287 7852 7343 7908
rect 7145 7710 7201 7766
rect 7287 7710 7343 7766
rect 7145 7568 7201 7624
rect 7287 7568 7343 7624
rect 7145 7426 7201 7482
rect 7287 7426 7343 7482
rect 7145 7284 7201 7340
rect 7287 7284 7343 7340
rect 7145 7142 7201 7198
rect 7287 7142 7343 7198
rect 7145 7000 7201 7056
rect 7287 7000 7343 7056
rect 7145 6858 7201 6914
rect 7287 6858 7343 6914
rect 7145 6716 7201 6772
rect 7287 6716 7343 6772
rect 7145 6574 7201 6630
rect 7287 6574 7343 6630
rect 7145 6432 7201 6488
rect 7287 6432 7343 6488
rect 7145 6290 7201 6346
rect 7287 6290 7343 6346
rect 7145 6148 7201 6204
rect 7287 6148 7343 6204
rect 7145 6006 7201 6062
rect 7287 6006 7343 6062
rect 7145 5864 7201 5920
rect 7287 5864 7343 5920
rect 7145 5722 7201 5778
rect 7287 5722 7343 5778
rect 7145 5580 7201 5636
rect 7287 5580 7343 5636
rect 7145 5438 7201 5494
rect 7287 5438 7343 5494
rect 7145 5296 7201 5352
rect 7287 5296 7343 5352
rect 7145 5154 7201 5210
rect 7287 5154 7343 5210
rect 7145 5012 7201 5068
rect 7287 5012 7343 5068
rect 7145 4870 7201 4926
rect 7287 4870 7343 4926
rect 7145 4728 7201 4784
rect 7287 4728 7343 4784
rect 7145 4586 7201 4642
rect 7287 4586 7343 4642
rect 7145 4444 7201 4500
rect 7287 4444 7343 4500
rect 7145 4302 7201 4358
rect 7287 4302 7343 4358
rect 7145 4160 7201 4216
rect 7287 4160 7343 4216
rect 7145 4018 7201 4074
rect 7287 4018 7343 4074
rect 7145 3876 7201 3932
rect 7287 3876 7343 3932
rect 7145 3734 7201 3790
rect 7287 3734 7343 3790
rect 7145 3592 7201 3648
rect 7287 3592 7343 3648
rect 7145 3450 7201 3506
rect 7287 3450 7343 3506
rect 7145 3308 7201 3364
rect 7287 3308 7343 3364
rect 7145 3166 7201 3222
rect 7287 3166 7343 3222
rect 7145 3024 7201 3080
rect 7287 3024 7343 3080
rect 7145 2882 7201 2938
rect 7287 2882 7343 2938
rect 7145 2740 7201 2796
rect 7287 2740 7343 2796
rect 7145 2598 7201 2654
rect 7287 2598 7343 2654
rect 7145 2456 7201 2512
rect 7287 2456 7343 2512
rect 7145 2314 7201 2370
rect 7287 2314 7343 2370
rect 7145 2172 7201 2228
rect 7287 2172 7343 2228
rect 7145 2030 7201 2086
rect 7287 2030 7343 2086
rect 7145 1888 7201 1944
rect 7287 1888 7343 1944
rect 7145 1746 7201 1802
rect 7287 1746 7343 1802
rect 7145 1604 7201 1660
rect 7287 1604 7343 1660
rect 7145 1462 7201 1518
rect 7287 1462 7343 1518
rect 7145 1320 7201 1376
rect 7287 1320 7343 1376
rect 7145 1178 7201 1234
rect 7287 1178 7343 1234
rect 7145 1036 7201 1092
rect 7287 1036 7343 1092
rect 7145 894 7201 950
rect 7287 894 7343 950
rect 7145 752 7201 808
rect 7287 752 7343 808
rect 7145 610 7201 666
rect 7287 610 7343 666
rect 7145 468 7201 524
rect 7287 468 7343 524
rect 7539 12254 7595 12310
rect 7681 12254 7737 12310
rect 7539 12112 7595 12168
rect 7681 12112 7737 12168
rect 7539 11970 7595 12026
rect 7681 11970 7737 12026
rect 7539 11828 7595 11884
rect 7681 11828 7737 11884
rect 7539 11686 7595 11742
rect 7681 11686 7737 11742
rect 7539 11544 7595 11600
rect 7681 11544 7737 11600
rect 7539 11402 7595 11458
rect 7681 11402 7737 11458
rect 7539 11260 7595 11316
rect 7681 11260 7737 11316
rect 7539 11118 7595 11174
rect 7681 11118 7737 11174
rect 7539 10976 7595 11032
rect 7681 10976 7737 11032
rect 7539 10834 7595 10890
rect 7681 10834 7737 10890
rect 7539 10692 7595 10748
rect 7681 10692 7737 10748
rect 7539 10550 7595 10606
rect 7681 10550 7737 10606
rect 7539 10408 7595 10464
rect 7681 10408 7737 10464
rect 7539 10266 7595 10322
rect 7681 10266 7737 10322
rect 7539 10124 7595 10180
rect 7681 10124 7737 10180
rect 7539 9982 7595 10038
rect 7681 9982 7737 10038
rect 7539 9840 7595 9896
rect 7681 9840 7737 9896
rect 7539 9698 7595 9754
rect 7681 9698 7737 9754
rect 7539 9556 7595 9612
rect 7681 9556 7737 9612
rect 7539 9414 7595 9470
rect 7681 9414 7737 9470
rect 7539 9272 7595 9328
rect 7681 9272 7737 9328
rect 7539 9130 7595 9186
rect 7681 9130 7737 9186
rect 7539 8988 7595 9044
rect 7681 8988 7737 9044
rect 7539 8846 7595 8902
rect 7681 8846 7737 8902
rect 7539 8704 7595 8760
rect 7681 8704 7737 8760
rect 7539 8562 7595 8618
rect 7681 8562 7737 8618
rect 7539 8420 7595 8476
rect 7681 8420 7737 8476
rect 7539 8278 7595 8334
rect 7681 8278 7737 8334
rect 7539 8136 7595 8192
rect 7681 8136 7737 8192
rect 7539 7994 7595 8050
rect 7681 7994 7737 8050
rect 7539 7852 7595 7908
rect 7681 7852 7737 7908
rect 7539 7710 7595 7766
rect 7681 7710 7737 7766
rect 7539 7568 7595 7624
rect 7681 7568 7737 7624
rect 7539 7426 7595 7482
rect 7681 7426 7737 7482
rect 7539 7284 7595 7340
rect 7681 7284 7737 7340
rect 7539 7142 7595 7198
rect 7681 7142 7737 7198
rect 7539 7000 7595 7056
rect 7681 7000 7737 7056
rect 7539 6858 7595 6914
rect 7681 6858 7737 6914
rect 7539 6716 7595 6772
rect 7681 6716 7737 6772
rect 7539 6574 7595 6630
rect 7681 6574 7737 6630
rect 7539 6432 7595 6488
rect 7681 6432 7737 6488
rect 7539 6290 7595 6346
rect 7681 6290 7737 6346
rect 7539 6148 7595 6204
rect 7681 6148 7737 6204
rect 7539 6006 7595 6062
rect 7681 6006 7737 6062
rect 7539 5864 7595 5920
rect 7681 5864 7737 5920
rect 7539 5722 7595 5778
rect 7681 5722 7737 5778
rect 7539 5580 7595 5636
rect 7681 5580 7737 5636
rect 7539 5438 7595 5494
rect 7681 5438 7737 5494
rect 7539 5296 7595 5352
rect 7681 5296 7737 5352
rect 7539 5154 7595 5210
rect 7681 5154 7737 5210
rect 7539 5012 7595 5068
rect 7681 5012 7737 5068
rect 7539 4870 7595 4926
rect 7681 4870 7737 4926
rect 7539 4728 7595 4784
rect 7681 4728 7737 4784
rect 7539 4586 7595 4642
rect 7681 4586 7737 4642
rect 7539 4444 7595 4500
rect 7681 4444 7737 4500
rect 7539 4302 7595 4358
rect 7681 4302 7737 4358
rect 7539 4160 7595 4216
rect 7681 4160 7737 4216
rect 7539 4018 7595 4074
rect 7681 4018 7737 4074
rect 7539 3876 7595 3932
rect 7681 3876 7737 3932
rect 7539 3734 7595 3790
rect 7681 3734 7737 3790
rect 7539 3592 7595 3648
rect 7681 3592 7737 3648
rect 7539 3450 7595 3506
rect 7681 3450 7737 3506
rect 7539 3308 7595 3364
rect 7681 3308 7737 3364
rect 7539 3166 7595 3222
rect 7681 3166 7737 3222
rect 7539 3024 7595 3080
rect 7681 3024 7737 3080
rect 7539 2882 7595 2938
rect 7681 2882 7737 2938
rect 7539 2740 7595 2796
rect 7681 2740 7737 2796
rect 7539 2598 7595 2654
rect 7681 2598 7737 2654
rect 7539 2456 7595 2512
rect 7681 2456 7737 2512
rect 7539 2314 7595 2370
rect 7681 2314 7737 2370
rect 7539 2172 7595 2228
rect 7681 2172 7737 2228
rect 7539 2030 7595 2086
rect 7681 2030 7737 2086
rect 7539 1888 7595 1944
rect 7681 1888 7737 1944
rect 7539 1746 7595 1802
rect 7681 1746 7737 1802
rect 7539 1604 7595 1660
rect 7681 1604 7737 1660
rect 7539 1462 7595 1518
rect 7681 1462 7737 1518
rect 7539 1320 7595 1376
rect 7681 1320 7737 1376
rect 7539 1178 7595 1234
rect 7681 1178 7737 1234
rect 7539 1036 7595 1092
rect 7681 1036 7737 1092
rect 7539 894 7595 950
rect 7681 894 7737 950
rect 7539 752 7595 808
rect 7681 752 7737 808
rect 7539 610 7595 666
rect 7681 610 7737 666
rect 7539 468 7595 524
rect 7681 468 7737 524
rect 7940 12254 7996 12310
rect 8082 12254 8138 12310
rect 7940 12112 7996 12168
rect 8082 12112 8138 12168
rect 7940 11970 7996 12026
rect 8082 11970 8138 12026
rect 7940 11828 7996 11884
rect 8082 11828 8138 11884
rect 7940 11686 7996 11742
rect 8082 11686 8138 11742
rect 7940 11544 7996 11600
rect 8082 11544 8138 11600
rect 7940 11402 7996 11458
rect 8082 11402 8138 11458
rect 7940 11260 7996 11316
rect 8082 11260 8138 11316
rect 7940 11118 7996 11174
rect 8082 11118 8138 11174
rect 7940 10976 7996 11032
rect 8082 10976 8138 11032
rect 7940 10834 7996 10890
rect 8082 10834 8138 10890
rect 7940 10692 7996 10748
rect 8082 10692 8138 10748
rect 7940 10550 7996 10606
rect 8082 10550 8138 10606
rect 7940 10408 7996 10464
rect 8082 10408 8138 10464
rect 7940 10266 7996 10322
rect 8082 10266 8138 10322
rect 7940 10124 7996 10180
rect 8082 10124 8138 10180
rect 7940 9982 7996 10038
rect 8082 9982 8138 10038
rect 7940 9840 7996 9896
rect 8082 9840 8138 9896
rect 7940 9698 7996 9754
rect 8082 9698 8138 9754
rect 7940 9556 7996 9612
rect 8082 9556 8138 9612
rect 7940 9414 7996 9470
rect 8082 9414 8138 9470
rect 7940 9272 7996 9328
rect 8082 9272 8138 9328
rect 7940 9130 7996 9186
rect 8082 9130 8138 9186
rect 7940 8988 7996 9044
rect 8082 8988 8138 9044
rect 7940 8846 7996 8902
rect 8082 8846 8138 8902
rect 7940 8704 7996 8760
rect 8082 8704 8138 8760
rect 7940 8562 7996 8618
rect 8082 8562 8138 8618
rect 7940 8420 7996 8476
rect 8082 8420 8138 8476
rect 7940 8278 7996 8334
rect 8082 8278 8138 8334
rect 7940 8136 7996 8192
rect 8082 8136 8138 8192
rect 7940 7994 7996 8050
rect 8082 7994 8138 8050
rect 7940 7852 7996 7908
rect 8082 7852 8138 7908
rect 7940 7710 7996 7766
rect 8082 7710 8138 7766
rect 7940 7568 7996 7624
rect 8082 7568 8138 7624
rect 7940 7426 7996 7482
rect 8082 7426 8138 7482
rect 7940 7284 7996 7340
rect 8082 7284 8138 7340
rect 7940 7142 7996 7198
rect 8082 7142 8138 7198
rect 7940 7000 7996 7056
rect 8082 7000 8138 7056
rect 7940 6858 7996 6914
rect 8082 6858 8138 6914
rect 7940 6716 7996 6772
rect 8082 6716 8138 6772
rect 7940 6574 7996 6630
rect 8082 6574 8138 6630
rect 7940 6432 7996 6488
rect 8082 6432 8138 6488
rect 7940 6290 7996 6346
rect 8082 6290 8138 6346
rect 7940 6148 7996 6204
rect 8082 6148 8138 6204
rect 7940 6006 7996 6062
rect 8082 6006 8138 6062
rect 7940 5864 7996 5920
rect 8082 5864 8138 5920
rect 7940 5722 7996 5778
rect 8082 5722 8138 5778
rect 7940 5580 7996 5636
rect 8082 5580 8138 5636
rect 7940 5438 7996 5494
rect 8082 5438 8138 5494
rect 7940 5296 7996 5352
rect 8082 5296 8138 5352
rect 7940 5154 7996 5210
rect 8082 5154 8138 5210
rect 7940 5012 7996 5068
rect 8082 5012 8138 5068
rect 7940 4870 7996 4926
rect 8082 4870 8138 4926
rect 7940 4728 7996 4784
rect 8082 4728 8138 4784
rect 7940 4586 7996 4642
rect 8082 4586 8138 4642
rect 7940 4444 7996 4500
rect 8082 4444 8138 4500
rect 7940 4302 7996 4358
rect 8082 4302 8138 4358
rect 7940 4160 7996 4216
rect 8082 4160 8138 4216
rect 7940 4018 7996 4074
rect 8082 4018 8138 4074
rect 7940 3876 7996 3932
rect 8082 3876 8138 3932
rect 7940 3734 7996 3790
rect 8082 3734 8138 3790
rect 7940 3592 7996 3648
rect 8082 3592 8138 3648
rect 7940 3450 7996 3506
rect 8082 3450 8138 3506
rect 7940 3308 7996 3364
rect 8082 3308 8138 3364
rect 7940 3166 7996 3222
rect 8082 3166 8138 3222
rect 7940 3024 7996 3080
rect 8082 3024 8138 3080
rect 7940 2882 7996 2938
rect 8082 2882 8138 2938
rect 7940 2740 7996 2796
rect 8082 2740 8138 2796
rect 7940 2598 7996 2654
rect 8082 2598 8138 2654
rect 7940 2456 7996 2512
rect 8082 2456 8138 2512
rect 7940 2314 7996 2370
rect 8082 2314 8138 2370
rect 7940 2172 7996 2228
rect 8082 2172 8138 2228
rect 7940 2030 7996 2086
rect 8082 2030 8138 2086
rect 7940 1888 7996 1944
rect 8082 1888 8138 1944
rect 7940 1746 7996 1802
rect 8082 1746 8138 1802
rect 7940 1604 7996 1660
rect 8082 1604 8138 1660
rect 7940 1462 7996 1518
rect 8082 1462 8138 1518
rect 7940 1320 7996 1376
rect 8082 1320 8138 1376
rect 7940 1178 7996 1234
rect 8082 1178 8138 1234
rect 7940 1036 7996 1092
rect 8082 1036 8138 1092
rect 7940 894 7996 950
rect 8082 894 8138 950
rect 7940 752 7996 808
rect 8082 752 8138 808
rect 7940 610 7996 666
rect 8082 610 8138 666
rect 7940 468 7996 524
rect 8082 468 8138 524
rect 8340 12254 8396 12310
rect 8482 12254 8538 12310
rect 8340 12112 8396 12168
rect 8482 12112 8538 12168
rect 8340 11970 8396 12026
rect 8482 11970 8538 12026
rect 8340 11828 8396 11884
rect 8482 11828 8538 11884
rect 8340 11686 8396 11742
rect 8482 11686 8538 11742
rect 8340 11544 8396 11600
rect 8482 11544 8538 11600
rect 8340 11402 8396 11458
rect 8482 11402 8538 11458
rect 8340 11260 8396 11316
rect 8482 11260 8538 11316
rect 8340 11118 8396 11174
rect 8482 11118 8538 11174
rect 8340 10976 8396 11032
rect 8482 10976 8538 11032
rect 8340 10834 8396 10890
rect 8482 10834 8538 10890
rect 8340 10692 8396 10748
rect 8482 10692 8538 10748
rect 8340 10550 8396 10606
rect 8482 10550 8538 10606
rect 8340 10408 8396 10464
rect 8482 10408 8538 10464
rect 8340 10266 8396 10322
rect 8482 10266 8538 10322
rect 8340 10124 8396 10180
rect 8482 10124 8538 10180
rect 8340 9982 8396 10038
rect 8482 9982 8538 10038
rect 8340 9840 8396 9896
rect 8482 9840 8538 9896
rect 8340 9698 8396 9754
rect 8482 9698 8538 9754
rect 8340 9556 8396 9612
rect 8482 9556 8538 9612
rect 8340 9414 8396 9470
rect 8482 9414 8538 9470
rect 8340 9272 8396 9328
rect 8482 9272 8538 9328
rect 8340 9130 8396 9186
rect 8482 9130 8538 9186
rect 8340 8988 8396 9044
rect 8482 8988 8538 9044
rect 8340 8846 8396 8902
rect 8482 8846 8538 8902
rect 8340 8704 8396 8760
rect 8482 8704 8538 8760
rect 8340 8562 8396 8618
rect 8482 8562 8538 8618
rect 8340 8420 8396 8476
rect 8482 8420 8538 8476
rect 8340 8278 8396 8334
rect 8482 8278 8538 8334
rect 8340 8136 8396 8192
rect 8482 8136 8538 8192
rect 8340 7994 8396 8050
rect 8482 7994 8538 8050
rect 8340 7852 8396 7908
rect 8482 7852 8538 7908
rect 8340 7710 8396 7766
rect 8482 7710 8538 7766
rect 8340 7568 8396 7624
rect 8482 7568 8538 7624
rect 8340 7426 8396 7482
rect 8482 7426 8538 7482
rect 8340 7284 8396 7340
rect 8482 7284 8538 7340
rect 8340 7142 8396 7198
rect 8482 7142 8538 7198
rect 8340 7000 8396 7056
rect 8482 7000 8538 7056
rect 8340 6858 8396 6914
rect 8482 6858 8538 6914
rect 8340 6716 8396 6772
rect 8482 6716 8538 6772
rect 8340 6574 8396 6630
rect 8482 6574 8538 6630
rect 8340 6432 8396 6488
rect 8482 6432 8538 6488
rect 8340 6290 8396 6346
rect 8482 6290 8538 6346
rect 8340 6148 8396 6204
rect 8482 6148 8538 6204
rect 8340 6006 8396 6062
rect 8482 6006 8538 6062
rect 8340 5864 8396 5920
rect 8482 5864 8538 5920
rect 8340 5722 8396 5778
rect 8482 5722 8538 5778
rect 8340 5580 8396 5636
rect 8482 5580 8538 5636
rect 8340 5438 8396 5494
rect 8482 5438 8538 5494
rect 8340 5296 8396 5352
rect 8482 5296 8538 5352
rect 8340 5154 8396 5210
rect 8482 5154 8538 5210
rect 8340 5012 8396 5068
rect 8482 5012 8538 5068
rect 8340 4870 8396 4926
rect 8482 4870 8538 4926
rect 8340 4728 8396 4784
rect 8482 4728 8538 4784
rect 8340 4586 8396 4642
rect 8482 4586 8538 4642
rect 8340 4444 8396 4500
rect 8482 4444 8538 4500
rect 8340 4302 8396 4358
rect 8482 4302 8538 4358
rect 8340 4160 8396 4216
rect 8482 4160 8538 4216
rect 8340 4018 8396 4074
rect 8482 4018 8538 4074
rect 8340 3876 8396 3932
rect 8482 3876 8538 3932
rect 8340 3734 8396 3790
rect 8482 3734 8538 3790
rect 8340 3592 8396 3648
rect 8482 3592 8538 3648
rect 8340 3450 8396 3506
rect 8482 3450 8538 3506
rect 8340 3308 8396 3364
rect 8482 3308 8538 3364
rect 8340 3166 8396 3222
rect 8482 3166 8538 3222
rect 8340 3024 8396 3080
rect 8482 3024 8538 3080
rect 8340 2882 8396 2938
rect 8482 2882 8538 2938
rect 8340 2740 8396 2796
rect 8482 2740 8538 2796
rect 8340 2598 8396 2654
rect 8482 2598 8538 2654
rect 8340 2456 8396 2512
rect 8482 2456 8538 2512
rect 8340 2314 8396 2370
rect 8482 2314 8538 2370
rect 8340 2172 8396 2228
rect 8482 2172 8538 2228
rect 8340 2030 8396 2086
rect 8482 2030 8538 2086
rect 8340 1888 8396 1944
rect 8482 1888 8538 1944
rect 8340 1746 8396 1802
rect 8482 1746 8538 1802
rect 8340 1604 8396 1660
rect 8482 1604 8538 1660
rect 8340 1462 8396 1518
rect 8482 1462 8538 1518
rect 8340 1320 8396 1376
rect 8482 1320 8538 1376
rect 8340 1178 8396 1234
rect 8482 1178 8538 1234
rect 8340 1036 8396 1092
rect 8482 1036 8538 1092
rect 8340 894 8396 950
rect 8482 894 8538 950
rect 8340 752 8396 808
rect 8482 752 8538 808
rect 8340 610 8396 666
rect 8482 610 8538 666
rect 8340 468 8396 524
rect 8482 468 8538 524
rect 8737 12254 8793 12310
rect 8879 12254 8935 12310
rect 8737 12112 8793 12168
rect 8879 12112 8935 12168
rect 8737 11970 8793 12026
rect 8879 11970 8935 12026
rect 8737 11828 8793 11884
rect 8879 11828 8935 11884
rect 8737 11686 8793 11742
rect 8879 11686 8935 11742
rect 8737 11544 8793 11600
rect 8879 11544 8935 11600
rect 8737 11402 8793 11458
rect 8879 11402 8935 11458
rect 8737 11260 8793 11316
rect 8879 11260 8935 11316
rect 8737 11118 8793 11174
rect 8879 11118 8935 11174
rect 8737 10976 8793 11032
rect 8879 10976 8935 11032
rect 8737 10834 8793 10890
rect 8879 10834 8935 10890
rect 8737 10692 8793 10748
rect 8879 10692 8935 10748
rect 8737 10550 8793 10606
rect 8879 10550 8935 10606
rect 8737 10408 8793 10464
rect 8879 10408 8935 10464
rect 8737 10266 8793 10322
rect 8879 10266 8935 10322
rect 8737 10124 8793 10180
rect 8879 10124 8935 10180
rect 8737 9982 8793 10038
rect 8879 9982 8935 10038
rect 8737 9840 8793 9896
rect 8879 9840 8935 9896
rect 8737 9698 8793 9754
rect 8879 9698 8935 9754
rect 8737 9556 8793 9612
rect 8879 9556 8935 9612
rect 8737 9414 8793 9470
rect 8879 9414 8935 9470
rect 8737 9272 8793 9328
rect 8879 9272 8935 9328
rect 8737 9130 8793 9186
rect 8879 9130 8935 9186
rect 8737 8988 8793 9044
rect 8879 8988 8935 9044
rect 8737 8846 8793 8902
rect 8879 8846 8935 8902
rect 8737 8704 8793 8760
rect 8879 8704 8935 8760
rect 8737 8562 8793 8618
rect 8879 8562 8935 8618
rect 8737 8420 8793 8476
rect 8879 8420 8935 8476
rect 8737 8278 8793 8334
rect 8879 8278 8935 8334
rect 8737 8136 8793 8192
rect 8879 8136 8935 8192
rect 8737 7994 8793 8050
rect 8879 7994 8935 8050
rect 8737 7852 8793 7908
rect 8879 7852 8935 7908
rect 8737 7710 8793 7766
rect 8879 7710 8935 7766
rect 8737 7568 8793 7624
rect 8879 7568 8935 7624
rect 8737 7426 8793 7482
rect 8879 7426 8935 7482
rect 8737 7284 8793 7340
rect 8879 7284 8935 7340
rect 8737 7142 8793 7198
rect 8879 7142 8935 7198
rect 8737 7000 8793 7056
rect 8879 7000 8935 7056
rect 8737 6858 8793 6914
rect 8879 6858 8935 6914
rect 8737 6716 8793 6772
rect 8879 6716 8935 6772
rect 8737 6574 8793 6630
rect 8879 6574 8935 6630
rect 8737 6432 8793 6488
rect 8879 6432 8935 6488
rect 8737 6290 8793 6346
rect 8879 6290 8935 6346
rect 8737 6148 8793 6204
rect 8879 6148 8935 6204
rect 8737 6006 8793 6062
rect 8879 6006 8935 6062
rect 8737 5864 8793 5920
rect 8879 5864 8935 5920
rect 8737 5722 8793 5778
rect 8879 5722 8935 5778
rect 8737 5580 8793 5636
rect 8879 5580 8935 5636
rect 8737 5438 8793 5494
rect 8879 5438 8935 5494
rect 8737 5296 8793 5352
rect 8879 5296 8935 5352
rect 8737 5154 8793 5210
rect 8879 5154 8935 5210
rect 8737 5012 8793 5068
rect 8879 5012 8935 5068
rect 8737 4870 8793 4926
rect 8879 4870 8935 4926
rect 8737 4728 8793 4784
rect 8879 4728 8935 4784
rect 8737 4586 8793 4642
rect 8879 4586 8935 4642
rect 8737 4444 8793 4500
rect 8879 4444 8935 4500
rect 8737 4302 8793 4358
rect 8879 4302 8935 4358
rect 8737 4160 8793 4216
rect 8879 4160 8935 4216
rect 8737 4018 8793 4074
rect 8879 4018 8935 4074
rect 8737 3876 8793 3932
rect 8879 3876 8935 3932
rect 8737 3734 8793 3790
rect 8879 3734 8935 3790
rect 8737 3592 8793 3648
rect 8879 3592 8935 3648
rect 8737 3450 8793 3506
rect 8879 3450 8935 3506
rect 8737 3308 8793 3364
rect 8879 3308 8935 3364
rect 8737 3166 8793 3222
rect 8879 3166 8935 3222
rect 8737 3024 8793 3080
rect 8879 3024 8935 3080
rect 8737 2882 8793 2938
rect 8879 2882 8935 2938
rect 8737 2740 8793 2796
rect 8879 2740 8935 2796
rect 8737 2598 8793 2654
rect 8879 2598 8935 2654
rect 8737 2456 8793 2512
rect 8879 2456 8935 2512
rect 8737 2314 8793 2370
rect 8879 2314 8935 2370
rect 8737 2172 8793 2228
rect 8879 2172 8935 2228
rect 8737 2030 8793 2086
rect 8879 2030 8935 2086
rect 8737 1888 8793 1944
rect 8879 1888 8935 1944
rect 8737 1746 8793 1802
rect 8879 1746 8935 1802
rect 8737 1604 8793 1660
rect 8879 1604 8935 1660
rect 8737 1462 8793 1518
rect 8879 1462 8935 1518
rect 8737 1320 8793 1376
rect 8879 1320 8935 1376
rect 8737 1178 8793 1234
rect 8879 1178 8935 1234
rect 8737 1036 8793 1092
rect 8879 1036 8935 1092
rect 8737 894 8793 950
rect 8879 894 8935 950
rect 8737 752 8793 808
rect 8879 752 8935 808
rect 8737 610 8793 666
rect 8879 610 8935 666
rect 8737 468 8793 524
rect 8879 468 8935 524
rect 9134 12254 9190 12310
rect 9276 12254 9332 12310
rect 9134 12112 9190 12168
rect 9276 12112 9332 12168
rect 9134 11970 9190 12026
rect 9276 11970 9332 12026
rect 9134 11828 9190 11884
rect 9276 11828 9332 11884
rect 9134 11686 9190 11742
rect 9276 11686 9332 11742
rect 9134 11544 9190 11600
rect 9276 11544 9332 11600
rect 9134 11402 9190 11458
rect 9276 11402 9332 11458
rect 9134 11260 9190 11316
rect 9276 11260 9332 11316
rect 9134 11118 9190 11174
rect 9276 11118 9332 11174
rect 9134 10976 9190 11032
rect 9276 10976 9332 11032
rect 9134 10834 9190 10890
rect 9276 10834 9332 10890
rect 9134 10692 9190 10748
rect 9276 10692 9332 10748
rect 9134 10550 9190 10606
rect 9276 10550 9332 10606
rect 9134 10408 9190 10464
rect 9276 10408 9332 10464
rect 9134 10266 9190 10322
rect 9276 10266 9332 10322
rect 9134 10124 9190 10180
rect 9276 10124 9332 10180
rect 9134 9982 9190 10038
rect 9276 9982 9332 10038
rect 9134 9840 9190 9896
rect 9276 9840 9332 9896
rect 9134 9698 9190 9754
rect 9276 9698 9332 9754
rect 9134 9556 9190 9612
rect 9276 9556 9332 9612
rect 9134 9414 9190 9470
rect 9276 9414 9332 9470
rect 9134 9272 9190 9328
rect 9276 9272 9332 9328
rect 9134 9130 9190 9186
rect 9276 9130 9332 9186
rect 9134 8988 9190 9044
rect 9276 8988 9332 9044
rect 9134 8846 9190 8902
rect 9276 8846 9332 8902
rect 9134 8704 9190 8760
rect 9276 8704 9332 8760
rect 9134 8562 9190 8618
rect 9276 8562 9332 8618
rect 9134 8420 9190 8476
rect 9276 8420 9332 8476
rect 9134 8278 9190 8334
rect 9276 8278 9332 8334
rect 9134 8136 9190 8192
rect 9276 8136 9332 8192
rect 9134 7994 9190 8050
rect 9276 7994 9332 8050
rect 9134 7852 9190 7908
rect 9276 7852 9332 7908
rect 9134 7710 9190 7766
rect 9276 7710 9332 7766
rect 9134 7568 9190 7624
rect 9276 7568 9332 7624
rect 9134 7426 9190 7482
rect 9276 7426 9332 7482
rect 9134 7284 9190 7340
rect 9276 7284 9332 7340
rect 9134 7142 9190 7198
rect 9276 7142 9332 7198
rect 9134 7000 9190 7056
rect 9276 7000 9332 7056
rect 9134 6858 9190 6914
rect 9276 6858 9332 6914
rect 9134 6716 9190 6772
rect 9276 6716 9332 6772
rect 9134 6574 9190 6630
rect 9276 6574 9332 6630
rect 9134 6432 9190 6488
rect 9276 6432 9332 6488
rect 9134 6290 9190 6346
rect 9276 6290 9332 6346
rect 9134 6148 9190 6204
rect 9276 6148 9332 6204
rect 9134 6006 9190 6062
rect 9276 6006 9332 6062
rect 9134 5864 9190 5920
rect 9276 5864 9332 5920
rect 9134 5722 9190 5778
rect 9276 5722 9332 5778
rect 9134 5580 9190 5636
rect 9276 5580 9332 5636
rect 9134 5438 9190 5494
rect 9276 5438 9332 5494
rect 9134 5296 9190 5352
rect 9276 5296 9332 5352
rect 9134 5154 9190 5210
rect 9276 5154 9332 5210
rect 9134 5012 9190 5068
rect 9276 5012 9332 5068
rect 9134 4870 9190 4926
rect 9276 4870 9332 4926
rect 9134 4728 9190 4784
rect 9276 4728 9332 4784
rect 9134 4586 9190 4642
rect 9276 4586 9332 4642
rect 9134 4444 9190 4500
rect 9276 4444 9332 4500
rect 9134 4302 9190 4358
rect 9276 4302 9332 4358
rect 9134 4160 9190 4216
rect 9276 4160 9332 4216
rect 9134 4018 9190 4074
rect 9276 4018 9332 4074
rect 9134 3876 9190 3932
rect 9276 3876 9332 3932
rect 9134 3734 9190 3790
rect 9276 3734 9332 3790
rect 9134 3592 9190 3648
rect 9276 3592 9332 3648
rect 9134 3450 9190 3506
rect 9276 3450 9332 3506
rect 9134 3308 9190 3364
rect 9276 3308 9332 3364
rect 9134 3166 9190 3222
rect 9276 3166 9332 3222
rect 9134 3024 9190 3080
rect 9276 3024 9332 3080
rect 9134 2882 9190 2938
rect 9276 2882 9332 2938
rect 9134 2740 9190 2796
rect 9276 2740 9332 2796
rect 9134 2598 9190 2654
rect 9276 2598 9332 2654
rect 9134 2456 9190 2512
rect 9276 2456 9332 2512
rect 9134 2314 9190 2370
rect 9276 2314 9332 2370
rect 9134 2172 9190 2228
rect 9276 2172 9332 2228
rect 9134 2030 9190 2086
rect 9276 2030 9332 2086
rect 9134 1888 9190 1944
rect 9276 1888 9332 1944
rect 9134 1746 9190 1802
rect 9276 1746 9332 1802
rect 9134 1604 9190 1660
rect 9276 1604 9332 1660
rect 9134 1462 9190 1518
rect 9276 1462 9332 1518
rect 9134 1320 9190 1376
rect 9276 1320 9332 1376
rect 9134 1178 9190 1234
rect 9276 1178 9332 1234
rect 9134 1036 9190 1092
rect 9276 1036 9332 1092
rect 9134 894 9190 950
rect 9276 894 9332 950
rect 9134 752 9190 808
rect 9276 752 9332 808
rect 9134 610 9190 666
rect 9276 610 9332 666
rect 9134 468 9190 524
rect 9276 468 9332 524
rect 9538 12254 9594 12310
rect 9680 12254 9736 12310
rect 9538 12112 9594 12168
rect 9680 12112 9736 12168
rect 9538 11970 9594 12026
rect 9680 11970 9736 12026
rect 9538 11828 9594 11884
rect 9680 11828 9736 11884
rect 9538 11686 9594 11742
rect 9680 11686 9736 11742
rect 9538 11544 9594 11600
rect 9680 11544 9736 11600
rect 9538 11402 9594 11458
rect 9680 11402 9736 11458
rect 9538 11260 9594 11316
rect 9680 11260 9736 11316
rect 9538 11118 9594 11174
rect 9680 11118 9736 11174
rect 9538 10976 9594 11032
rect 9680 10976 9736 11032
rect 9538 10834 9594 10890
rect 9680 10834 9736 10890
rect 9538 10692 9594 10748
rect 9680 10692 9736 10748
rect 9538 10550 9594 10606
rect 9680 10550 9736 10606
rect 9538 10408 9594 10464
rect 9680 10408 9736 10464
rect 9538 10266 9594 10322
rect 9680 10266 9736 10322
rect 9538 10124 9594 10180
rect 9680 10124 9736 10180
rect 9538 9982 9594 10038
rect 9680 9982 9736 10038
rect 9538 9840 9594 9896
rect 9680 9840 9736 9896
rect 9538 9698 9594 9754
rect 9680 9698 9736 9754
rect 9538 9556 9594 9612
rect 9680 9556 9736 9612
rect 9538 9414 9594 9470
rect 9680 9414 9736 9470
rect 9538 9272 9594 9328
rect 9680 9272 9736 9328
rect 9538 9130 9594 9186
rect 9680 9130 9736 9186
rect 9538 8988 9594 9044
rect 9680 8988 9736 9044
rect 9538 8846 9594 8902
rect 9680 8846 9736 8902
rect 9538 8704 9594 8760
rect 9680 8704 9736 8760
rect 9538 8562 9594 8618
rect 9680 8562 9736 8618
rect 9538 8420 9594 8476
rect 9680 8420 9736 8476
rect 9538 8278 9594 8334
rect 9680 8278 9736 8334
rect 9538 8136 9594 8192
rect 9680 8136 9736 8192
rect 9538 7994 9594 8050
rect 9680 7994 9736 8050
rect 9538 7852 9594 7908
rect 9680 7852 9736 7908
rect 9538 7710 9594 7766
rect 9680 7710 9736 7766
rect 9538 7568 9594 7624
rect 9680 7568 9736 7624
rect 9538 7426 9594 7482
rect 9680 7426 9736 7482
rect 9538 7284 9594 7340
rect 9680 7284 9736 7340
rect 9538 7142 9594 7198
rect 9680 7142 9736 7198
rect 9538 7000 9594 7056
rect 9680 7000 9736 7056
rect 9538 6858 9594 6914
rect 9680 6858 9736 6914
rect 9538 6716 9594 6772
rect 9680 6716 9736 6772
rect 9538 6574 9594 6630
rect 9680 6574 9736 6630
rect 9538 6432 9594 6488
rect 9680 6432 9736 6488
rect 9538 6290 9594 6346
rect 9680 6290 9736 6346
rect 9538 6148 9594 6204
rect 9680 6148 9736 6204
rect 9538 6006 9594 6062
rect 9680 6006 9736 6062
rect 9538 5864 9594 5920
rect 9680 5864 9736 5920
rect 9538 5722 9594 5778
rect 9680 5722 9736 5778
rect 9538 5580 9594 5636
rect 9680 5580 9736 5636
rect 9538 5438 9594 5494
rect 9680 5438 9736 5494
rect 9538 5296 9594 5352
rect 9680 5296 9736 5352
rect 9538 5154 9594 5210
rect 9680 5154 9736 5210
rect 9538 5012 9594 5068
rect 9680 5012 9736 5068
rect 9538 4870 9594 4926
rect 9680 4870 9736 4926
rect 9538 4728 9594 4784
rect 9680 4728 9736 4784
rect 9538 4586 9594 4642
rect 9680 4586 9736 4642
rect 9538 4444 9594 4500
rect 9680 4444 9736 4500
rect 9538 4302 9594 4358
rect 9680 4302 9736 4358
rect 9538 4160 9594 4216
rect 9680 4160 9736 4216
rect 9538 4018 9594 4074
rect 9680 4018 9736 4074
rect 9538 3876 9594 3932
rect 9680 3876 9736 3932
rect 9538 3734 9594 3790
rect 9680 3734 9736 3790
rect 9538 3592 9594 3648
rect 9680 3592 9736 3648
rect 9538 3450 9594 3506
rect 9680 3450 9736 3506
rect 9538 3308 9594 3364
rect 9680 3308 9736 3364
rect 9538 3166 9594 3222
rect 9680 3166 9736 3222
rect 9538 3024 9594 3080
rect 9680 3024 9736 3080
rect 9538 2882 9594 2938
rect 9680 2882 9736 2938
rect 9538 2740 9594 2796
rect 9680 2740 9736 2796
rect 9538 2598 9594 2654
rect 9680 2598 9736 2654
rect 9538 2456 9594 2512
rect 9680 2456 9736 2512
rect 9538 2314 9594 2370
rect 9680 2314 9736 2370
rect 9538 2172 9594 2228
rect 9680 2172 9736 2228
rect 9538 2030 9594 2086
rect 9680 2030 9736 2086
rect 9538 1888 9594 1944
rect 9680 1888 9736 1944
rect 9538 1746 9594 1802
rect 9680 1746 9736 1802
rect 9538 1604 9594 1660
rect 9680 1604 9736 1660
rect 9538 1462 9594 1518
rect 9680 1462 9736 1518
rect 9538 1320 9594 1376
rect 9680 1320 9736 1376
rect 9538 1178 9594 1234
rect 9680 1178 9736 1234
rect 9538 1036 9594 1092
rect 9680 1036 9736 1092
rect 9538 894 9594 950
rect 9680 894 9736 950
rect 9538 752 9594 808
rect 9680 752 9736 808
rect 9538 610 9594 666
rect 9680 610 9736 666
rect 9538 468 9594 524
rect 9680 468 9736 524
rect 9934 12254 9990 12310
rect 10076 12254 10132 12310
rect 9934 12112 9990 12168
rect 10076 12112 10132 12168
rect 9934 11970 9990 12026
rect 10076 11970 10132 12026
rect 9934 11828 9990 11884
rect 10076 11828 10132 11884
rect 9934 11686 9990 11742
rect 10076 11686 10132 11742
rect 9934 11544 9990 11600
rect 10076 11544 10132 11600
rect 9934 11402 9990 11458
rect 10076 11402 10132 11458
rect 9934 11260 9990 11316
rect 10076 11260 10132 11316
rect 9934 11118 9990 11174
rect 10076 11118 10132 11174
rect 9934 10976 9990 11032
rect 10076 10976 10132 11032
rect 9934 10834 9990 10890
rect 10076 10834 10132 10890
rect 9934 10692 9990 10748
rect 10076 10692 10132 10748
rect 9934 10550 9990 10606
rect 10076 10550 10132 10606
rect 9934 10408 9990 10464
rect 10076 10408 10132 10464
rect 9934 10266 9990 10322
rect 10076 10266 10132 10322
rect 9934 10124 9990 10180
rect 10076 10124 10132 10180
rect 9934 9982 9990 10038
rect 10076 9982 10132 10038
rect 9934 9840 9990 9896
rect 10076 9840 10132 9896
rect 9934 9698 9990 9754
rect 10076 9698 10132 9754
rect 9934 9556 9990 9612
rect 10076 9556 10132 9612
rect 9934 9414 9990 9470
rect 10076 9414 10132 9470
rect 9934 9272 9990 9328
rect 10076 9272 10132 9328
rect 9934 9130 9990 9186
rect 10076 9130 10132 9186
rect 9934 8988 9990 9044
rect 10076 8988 10132 9044
rect 9934 8846 9990 8902
rect 10076 8846 10132 8902
rect 9934 8704 9990 8760
rect 10076 8704 10132 8760
rect 9934 8562 9990 8618
rect 10076 8562 10132 8618
rect 9934 8420 9990 8476
rect 10076 8420 10132 8476
rect 9934 8278 9990 8334
rect 10076 8278 10132 8334
rect 9934 8136 9990 8192
rect 10076 8136 10132 8192
rect 9934 7994 9990 8050
rect 10076 7994 10132 8050
rect 9934 7852 9990 7908
rect 10076 7852 10132 7908
rect 9934 7710 9990 7766
rect 10076 7710 10132 7766
rect 9934 7568 9990 7624
rect 10076 7568 10132 7624
rect 9934 7426 9990 7482
rect 10076 7426 10132 7482
rect 9934 7284 9990 7340
rect 10076 7284 10132 7340
rect 9934 7142 9990 7198
rect 10076 7142 10132 7198
rect 9934 7000 9990 7056
rect 10076 7000 10132 7056
rect 9934 6858 9990 6914
rect 10076 6858 10132 6914
rect 9934 6716 9990 6772
rect 10076 6716 10132 6772
rect 9934 6574 9990 6630
rect 10076 6574 10132 6630
rect 9934 6432 9990 6488
rect 10076 6432 10132 6488
rect 9934 6290 9990 6346
rect 10076 6290 10132 6346
rect 9934 6148 9990 6204
rect 10076 6148 10132 6204
rect 9934 6006 9990 6062
rect 10076 6006 10132 6062
rect 9934 5864 9990 5920
rect 10076 5864 10132 5920
rect 9934 5722 9990 5778
rect 10076 5722 10132 5778
rect 9934 5580 9990 5636
rect 10076 5580 10132 5636
rect 9934 5438 9990 5494
rect 10076 5438 10132 5494
rect 9934 5296 9990 5352
rect 10076 5296 10132 5352
rect 9934 5154 9990 5210
rect 10076 5154 10132 5210
rect 9934 5012 9990 5068
rect 10076 5012 10132 5068
rect 9934 4870 9990 4926
rect 10076 4870 10132 4926
rect 9934 4728 9990 4784
rect 10076 4728 10132 4784
rect 9934 4586 9990 4642
rect 10076 4586 10132 4642
rect 9934 4444 9990 4500
rect 10076 4444 10132 4500
rect 9934 4302 9990 4358
rect 10076 4302 10132 4358
rect 9934 4160 9990 4216
rect 10076 4160 10132 4216
rect 9934 4018 9990 4074
rect 10076 4018 10132 4074
rect 9934 3876 9990 3932
rect 10076 3876 10132 3932
rect 9934 3734 9990 3790
rect 10076 3734 10132 3790
rect 9934 3592 9990 3648
rect 10076 3592 10132 3648
rect 9934 3450 9990 3506
rect 10076 3450 10132 3506
rect 9934 3308 9990 3364
rect 10076 3308 10132 3364
rect 9934 3166 9990 3222
rect 10076 3166 10132 3222
rect 9934 3024 9990 3080
rect 10076 3024 10132 3080
rect 9934 2882 9990 2938
rect 10076 2882 10132 2938
rect 9934 2740 9990 2796
rect 10076 2740 10132 2796
rect 9934 2598 9990 2654
rect 10076 2598 10132 2654
rect 9934 2456 9990 2512
rect 10076 2456 10132 2512
rect 9934 2314 9990 2370
rect 10076 2314 10132 2370
rect 9934 2172 9990 2228
rect 10076 2172 10132 2228
rect 9934 2030 9990 2086
rect 10076 2030 10132 2086
rect 9934 1888 9990 1944
rect 10076 1888 10132 1944
rect 9934 1746 9990 1802
rect 10076 1746 10132 1802
rect 9934 1604 9990 1660
rect 10076 1604 10132 1660
rect 9934 1462 9990 1518
rect 10076 1462 10132 1518
rect 9934 1320 9990 1376
rect 10076 1320 10132 1376
rect 9934 1178 9990 1234
rect 10076 1178 10132 1234
rect 9934 1036 9990 1092
rect 10076 1036 10132 1092
rect 9934 894 9990 950
rect 10076 894 10132 950
rect 9934 752 9990 808
rect 10076 752 10132 808
rect 9934 610 9990 666
rect 10076 610 10132 666
rect 9934 468 9990 524
rect 10076 468 10132 524
rect 10334 12254 10390 12310
rect 10476 12254 10532 12310
rect 10334 12112 10390 12168
rect 10476 12112 10532 12168
rect 10334 11970 10390 12026
rect 10476 11970 10532 12026
rect 10334 11828 10390 11884
rect 10476 11828 10532 11884
rect 10334 11686 10390 11742
rect 10476 11686 10532 11742
rect 10334 11544 10390 11600
rect 10476 11544 10532 11600
rect 10334 11402 10390 11458
rect 10476 11402 10532 11458
rect 10334 11260 10390 11316
rect 10476 11260 10532 11316
rect 10334 11118 10390 11174
rect 10476 11118 10532 11174
rect 10334 10976 10390 11032
rect 10476 10976 10532 11032
rect 10334 10834 10390 10890
rect 10476 10834 10532 10890
rect 10334 10692 10390 10748
rect 10476 10692 10532 10748
rect 10334 10550 10390 10606
rect 10476 10550 10532 10606
rect 10334 10408 10390 10464
rect 10476 10408 10532 10464
rect 10334 10266 10390 10322
rect 10476 10266 10532 10322
rect 10334 10124 10390 10180
rect 10476 10124 10532 10180
rect 10334 9982 10390 10038
rect 10476 9982 10532 10038
rect 10334 9840 10390 9896
rect 10476 9840 10532 9896
rect 10334 9698 10390 9754
rect 10476 9698 10532 9754
rect 10334 9556 10390 9612
rect 10476 9556 10532 9612
rect 10334 9414 10390 9470
rect 10476 9414 10532 9470
rect 10334 9272 10390 9328
rect 10476 9272 10532 9328
rect 10334 9130 10390 9186
rect 10476 9130 10532 9186
rect 10334 8988 10390 9044
rect 10476 8988 10532 9044
rect 10334 8846 10390 8902
rect 10476 8846 10532 8902
rect 10334 8704 10390 8760
rect 10476 8704 10532 8760
rect 10334 8562 10390 8618
rect 10476 8562 10532 8618
rect 10334 8420 10390 8476
rect 10476 8420 10532 8476
rect 10334 8278 10390 8334
rect 10476 8278 10532 8334
rect 10334 8136 10390 8192
rect 10476 8136 10532 8192
rect 10334 7994 10390 8050
rect 10476 7994 10532 8050
rect 10334 7852 10390 7908
rect 10476 7852 10532 7908
rect 10334 7710 10390 7766
rect 10476 7710 10532 7766
rect 10334 7568 10390 7624
rect 10476 7568 10532 7624
rect 10334 7426 10390 7482
rect 10476 7426 10532 7482
rect 10334 7284 10390 7340
rect 10476 7284 10532 7340
rect 10334 7142 10390 7198
rect 10476 7142 10532 7198
rect 10334 7000 10390 7056
rect 10476 7000 10532 7056
rect 10334 6858 10390 6914
rect 10476 6858 10532 6914
rect 10334 6716 10390 6772
rect 10476 6716 10532 6772
rect 10334 6574 10390 6630
rect 10476 6574 10532 6630
rect 10334 6432 10390 6488
rect 10476 6432 10532 6488
rect 10334 6290 10390 6346
rect 10476 6290 10532 6346
rect 10334 6148 10390 6204
rect 10476 6148 10532 6204
rect 10334 6006 10390 6062
rect 10476 6006 10532 6062
rect 10334 5864 10390 5920
rect 10476 5864 10532 5920
rect 10334 5722 10390 5778
rect 10476 5722 10532 5778
rect 10334 5580 10390 5636
rect 10476 5580 10532 5636
rect 10334 5438 10390 5494
rect 10476 5438 10532 5494
rect 10334 5296 10390 5352
rect 10476 5296 10532 5352
rect 10334 5154 10390 5210
rect 10476 5154 10532 5210
rect 10334 5012 10390 5068
rect 10476 5012 10532 5068
rect 10334 4870 10390 4926
rect 10476 4870 10532 4926
rect 10334 4728 10390 4784
rect 10476 4728 10532 4784
rect 10334 4586 10390 4642
rect 10476 4586 10532 4642
rect 10334 4444 10390 4500
rect 10476 4444 10532 4500
rect 10334 4302 10390 4358
rect 10476 4302 10532 4358
rect 10334 4160 10390 4216
rect 10476 4160 10532 4216
rect 10334 4018 10390 4074
rect 10476 4018 10532 4074
rect 10334 3876 10390 3932
rect 10476 3876 10532 3932
rect 10334 3734 10390 3790
rect 10476 3734 10532 3790
rect 10334 3592 10390 3648
rect 10476 3592 10532 3648
rect 10334 3450 10390 3506
rect 10476 3450 10532 3506
rect 10334 3308 10390 3364
rect 10476 3308 10532 3364
rect 10334 3166 10390 3222
rect 10476 3166 10532 3222
rect 10334 3024 10390 3080
rect 10476 3024 10532 3080
rect 10334 2882 10390 2938
rect 10476 2882 10532 2938
rect 10334 2740 10390 2796
rect 10476 2740 10532 2796
rect 10334 2598 10390 2654
rect 10476 2598 10532 2654
rect 10334 2456 10390 2512
rect 10476 2456 10532 2512
rect 10334 2314 10390 2370
rect 10476 2314 10532 2370
rect 10334 2172 10390 2228
rect 10476 2172 10532 2228
rect 10334 2030 10390 2086
rect 10476 2030 10532 2086
rect 10334 1888 10390 1944
rect 10476 1888 10532 1944
rect 10334 1746 10390 1802
rect 10476 1746 10532 1802
rect 10334 1604 10390 1660
rect 10476 1604 10532 1660
rect 10334 1462 10390 1518
rect 10476 1462 10532 1518
rect 10334 1320 10390 1376
rect 10476 1320 10532 1376
rect 10334 1178 10390 1234
rect 10476 1178 10532 1234
rect 10334 1036 10390 1092
rect 10476 1036 10532 1092
rect 10334 894 10390 950
rect 10476 894 10532 950
rect 10334 752 10390 808
rect 10476 752 10532 808
rect 10334 610 10390 666
rect 10476 610 10532 666
rect 10334 468 10390 524
rect 10476 468 10532 524
rect 10731 12254 10787 12310
rect 10873 12254 10929 12310
rect 10731 12112 10787 12168
rect 10873 12112 10929 12168
rect 10731 11970 10787 12026
rect 10873 11970 10929 12026
rect 10731 11828 10787 11884
rect 10873 11828 10929 11884
rect 10731 11686 10787 11742
rect 10873 11686 10929 11742
rect 10731 11544 10787 11600
rect 10873 11544 10929 11600
rect 10731 11402 10787 11458
rect 10873 11402 10929 11458
rect 10731 11260 10787 11316
rect 10873 11260 10929 11316
rect 10731 11118 10787 11174
rect 10873 11118 10929 11174
rect 10731 10976 10787 11032
rect 10873 10976 10929 11032
rect 10731 10834 10787 10890
rect 10873 10834 10929 10890
rect 10731 10692 10787 10748
rect 10873 10692 10929 10748
rect 10731 10550 10787 10606
rect 10873 10550 10929 10606
rect 10731 10408 10787 10464
rect 10873 10408 10929 10464
rect 10731 10266 10787 10322
rect 10873 10266 10929 10322
rect 10731 10124 10787 10180
rect 10873 10124 10929 10180
rect 10731 9982 10787 10038
rect 10873 9982 10929 10038
rect 10731 9840 10787 9896
rect 10873 9840 10929 9896
rect 10731 9698 10787 9754
rect 10873 9698 10929 9754
rect 10731 9556 10787 9612
rect 10873 9556 10929 9612
rect 10731 9414 10787 9470
rect 10873 9414 10929 9470
rect 10731 9272 10787 9328
rect 10873 9272 10929 9328
rect 10731 9130 10787 9186
rect 10873 9130 10929 9186
rect 10731 8988 10787 9044
rect 10873 8988 10929 9044
rect 10731 8846 10787 8902
rect 10873 8846 10929 8902
rect 10731 8704 10787 8760
rect 10873 8704 10929 8760
rect 10731 8562 10787 8618
rect 10873 8562 10929 8618
rect 10731 8420 10787 8476
rect 10873 8420 10929 8476
rect 10731 8278 10787 8334
rect 10873 8278 10929 8334
rect 10731 8136 10787 8192
rect 10873 8136 10929 8192
rect 10731 7994 10787 8050
rect 10873 7994 10929 8050
rect 10731 7852 10787 7908
rect 10873 7852 10929 7908
rect 10731 7710 10787 7766
rect 10873 7710 10929 7766
rect 10731 7568 10787 7624
rect 10873 7568 10929 7624
rect 10731 7426 10787 7482
rect 10873 7426 10929 7482
rect 10731 7284 10787 7340
rect 10873 7284 10929 7340
rect 10731 7142 10787 7198
rect 10873 7142 10929 7198
rect 10731 7000 10787 7056
rect 10873 7000 10929 7056
rect 10731 6858 10787 6914
rect 10873 6858 10929 6914
rect 10731 6716 10787 6772
rect 10873 6716 10929 6772
rect 10731 6574 10787 6630
rect 10873 6574 10929 6630
rect 10731 6432 10787 6488
rect 10873 6432 10929 6488
rect 10731 6290 10787 6346
rect 10873 6290 10929 6346
rect 10731 6148 10787 6204
rect 10873 6148 10929 6204
rect 10731 6006 10787 6062
rect 10873 6006 10929 6062
rect 10731 5864 10787 5920
rect 10873 5864 10929 5920
rect 10731 5722 10787 5778
rect 10873 5722 10929 5778
rect 10731 5580 10787 5636
rect 10873 5580 10929 5636
rect 10731 5438 10787 5494
rect 10873 5438 10929 5494
rect 10731 5296 10787 5352
rect 10873 5296 10929 5352
rect 10731 5154 10787 5210
rect 10873 5154 10929 5210
rect 10731 5012 10787 5068
rect 10873 5012 10929 5068
rect 10731 4870 10787 4926
rect 10873 4870 10929 4926
rect 10731 4728 10787 4784
rect 10873 4728 10929 4784
rect 10731 4586 10787 4642
rect 10873 4586 10929 4642
rect 10731 4444 10787 4500
rect 10873 4444 10929 4500
rect 10731 4302 10787 4358
rect 10873 4302 10929 4358
rect 10731 4160 10787 4216
rect 10873 4160 10929 4216
rect 10731 4018 10787 4074
rect 10873 4018 10929 4074
rect 10731 3876 10787 3932
rect 10873 3876 10929 3932
rect 10731 3734 10787 3790
rect 10873 3734 10929 3790
rect 10731 3592 10787 3648
rect 10873 3592 10929 3648
rect 10731 3450 10787 3506
rect 10873 3450 10929 3506
rect 10731 3308 10787 3364
rect 10873 3308 10929 3364
rect 10731 3166 10787 3222
rect 10873 3166 10929 3222
rect 10731 3024 10787 3080
rect 10873 3024 10929 3080
rect 10731 2882 10787 2938
rect 10873 2882 10929 2938
rect 10731 2740 10787 2796
rect 10873 2740 10929 2796
rect 10731 2598 10787 2654
rect 10873 2598 10929 2654
rect 10731 2456 10787 2512
rect 10873 2456 10929 2512
rect 10731 2314 10787 2370
rect 10873 2314 10929 2370
rect 10731 2172 10787 2228
rect 10873 2172 10929 2228
rect 10731 2030 10787 2086
rect 10873 2030 10929 2086
rect 10731 1888 10787 1944
rect 10873 1888 10929 1944
rect 10731 1746 10787 1802
rect 10873 1746 10929 1802
rect 10731 1604 10787 1660
rect 10873 1604 10929 1660
rect 10731 1462 10787 1518
rect 10873 1462 10929 1518
rect 10731 1320 10787 1376
rect 10873 1320 10929 1376
rect 10731 1178 10787 1234
rect 10873 1178 10929 1234
rect 10731 1036 10787 1092
rect 10873 1036 10929 1092
rect 10731 894 10787 950
rect 10873 894 10929 950
rect 10731 752 10787 808
rect 10873 752 10929 808
rect 10731 610 10787 666
rect 10873 610 10929 666
rect 10731 468 10787 524
rect 10873 468 10929 524
rect 11136 12254 11192 12310
rect 11278 12254 11334 12310
rect 11136 12112 11192 12168
rect 11278 12112 11334 12168
rect 11136 11970 11192 12026
rect 11278 11970 11334 12026
rect 11136 11828 11192 11884
rect 11278 11828 11334 11884
rect 11136 11686 11192 11742
rect 11278 11686 11334 11742
rect 11136 11544 11192 11600
rect 11278 11544 11334 11600
rect 11136 11402 11192 11458
rect 11278 11402 11334 11458
rect 11136 11260 11192 11316
rect 11278 11260 11334 11316
rect 11136 11118 11192 11174
rect 11278 11118 11334 11174
rect 11136 10976 11192 11032
rect 11278 10976 11334 11032
rect 11136 10834 11192 10890
rect 11278 10834 11334 10890
rect 11136 10692 11192 10748
rect 11278 10692 11334 10748
rect 11136 10550 11192 10606
rect 11278 10550 11334 10606
rect 11136 10408 11192 10464
rect 11278 10408 11334 10464
rect 11136 10266 11192 10322
rect 11278 10266 11334 10322
rect 11136 10124 11192 10180
rect 11278 10124 11334 10180
rect 11136 9982 11192 10038
rect 11278 9982 11334 10038
rect 11136 9840 11192 9896
rect 11278 9840 11334 9896
rect 11136 9698 11192 9754
rect 11278 9698 11334 9754
rect 11136 9556 11192 9612
rect 11278 9556 11334 9612
rect 11136 9414 11192 9470
rect 11278 9414 11334 9470
rect 11136 9272 11192 9328
rect 11278 9272 11334 9328
rect 11136 9130 11192 9186
rect 11278 9130 11334 9186
rect 11136 8988 11192 9044
rect 11278 8988 11334 9044
rect 11136 8846 11192 8902
rect 11278 8846 11334 8902
rect 11136 8704 11192 8760
rect 11278 8704 11334 8760
rect 11136 8562 11192 8618
rect 11278 8562 11334 8618
rect 11136 8420 11192 8476
rect 11278 8420 11334 8476
rect 11136 8278 11192 8334
rect 11278 8278 11334 8334
rect 11136 8136 11192 8192
rect 11278 8136 11334 8192
rect 11136 7994 11192 8050
rect 11278 7994 11334 8050
rect 11136 7852 11192 7908
rect 11278 7852 11334 7908
rect 11136 7710 11192 7766
rect 11278 7710 11334 7766
rect 11136 7568 11192 7624
rect 11278 7568 11334 7624
rect 11136 7426 11192 7482
rect 11278 7426 11334 7482
rect 11136 7284 11192 7340
rect 11278 7284 11334 7340
rect 11136 7142 11192 7198
rect 11278 7142 11334 7198
rect 11136 7000 11192 7056
rect 11278 7000 11334 7056
rect 11136 6858 11192 6914
rect 11278 6858 11334 6914
rect 11136 6716 11192 6772
rect 11278 6716 11334 6772
rect 11136 6574 11192 6630
rect 11278 6574 11334 6630
rect 11136 6432 11192 6488
rect 11278 6432 11334 6488
rect 11136 6290 11192 6346
rect 11278 6290 11334 6346
rect 11136 6148 11192 6204
rect 11278 6148 11334 6204
rect 11136 6006 11192 6062
rect 11278 6006 11334 6062
rect 11136 5864 11192 5920
rect 11278 5864 11334 5920
rect 11136 5722 11192 5778
rect 11278 5722 11334 5778
rect 11136 5580 11192 5636
rect 11278 5580 11334 5636
rect 11136 5438 11192 5494
rect 11278 5438 11334 5494
rect 11136 5296 11192 5352
rect 11278 5296 11334 5352
rect 11136 5154 11192 5210
rect 11278 5154 11334 5210
rect 11136 5012 11192 5068
rect 11278 5012 11334 5068
rect 11136 4870 11192 4926
rect 11278 4870 11334 4926
rect 11136 4728 11192 4784
rect 11278 4728 11334 4784
rect 11136 4586 11192 4642
rect 11278 4586 11334 4642
rect 11136 4444 11192 4500
rect 11278 4444 11334 4500
rect 11136 4302 11192 4358
rect 11278 4302 11334 4358
rect 11136 4160 11192 4216
rect 11278 4160 11334 4216
rect 11136 4018 11192 4074
rect 11278 4018 11334 4074
rect 11136 3876 11192 3932
rect 11278 3876 11334 3932
rect 11136 3734 11192 3790
rect 11278 3734 11334 3790
rect 11136 3592 11192 3648
rect 11278 3592 11334 3648
rect 11136 3450 11192 3506
rect 11278 3450 11334 3506
rect 11136 3308 11192 3364
rect 11278 3308 11334 3364
rect 11136 3166 11192 3222
rect 11278 3166 11334 3222
rect 11136 3024 11192 3080
rect 11278 3024 11334 3080
rect 11136 2882 11192 2938
rect 11278 2882 11334 2938
rect 11136 2740 11192 2796
rect 11278 2740 11334 2796
rect 11136 2598 11192 2654
rect 11278 2598 11334 2654
rect 11136 2456 11192 2512
rect 11278 2456 11334 2512
rect 11136 2314 11192 2370
rect 11278 2314 11334 2370
rect 11136 2172 11192 2228
rect 11278 2172 11334 2228
rect 11136 2030 11192 2086
rect 11278 2030 11334 2086
rect 11136 1888 11192 1944
rect 11278 1888 11334 1944
rect 11136 1746 11192 1802
rect 11278 1746 11334 1802
rect 11136 1604 11192 1660
rect 11278 1604 11334 1660
rect 11136 1462 11192 1518
rect 11278 1462 11334 1518
rect 11136 1320 11192 1376
rect 11278 1320 11334 1376
rect 11136 1178 11192 1234
rect 11278 1178 11334 1234
rect 11136 1036 11192 1092
rect 11278 1036 11334 1092
rect 11136 894 11192 950
rect 11278 894 11334 950
rect 11136 752 11192 808
rect 11278 752 11334 808
rect 11136 610 11192 666
rect 11278 610 11334 666
rect 11136 468 11192 524
rect 11278 468 11334 524
rect 11536 12254 11592 12310
rect 11678 12254 11734 12310
rect 11536 12112 11592 12168
rect 11678 12112 11734 12168
rect 11536 11970 11592 12026
rect 11678 11970 11734 12026
rect 11536 11828 11592 11884
rect 11678 11828 11734 11884
rect 11536 11686 11592 11742
rect 11678 11686 11734 11742
rect 11536 11544 11592 11600
rect 11678 11544 11734 11600
rect 11536 11402 11592 11458
rect 11678 11402 11734 11458
rect 11536 11260 11592 11316
rect 11678 11260 11734 11316
rect 11536 11118 11592 11174
rect 11678 11118 11734 11174
rect 11536 10976 11592 11032
rect 11678 10976 11734 11032
rect 11536 10834 11592 10890
rect 11678 10834 11734 10890
rect 11536 10692 11592 10748
rect 11678 10692 11734 10748
rect 11536 10550 11592 10606
rect 11678 10550 11734 10606
rect 11536 10408 11592 10464
rect 11678 10408 11734 10464
rect 11536 10266 11592 10322
rect 11678 10266 11734 10322
rect 11536 10124 11592 10180
rect 11678 10124 11734 10180
rect 11536 9982 11592 10038
rect 11678 9982 11734 10038
rect 11536 9840 11592 9896
rect 11678 9840 11734 9896
rect 11536 9698 11592 9754
rect 11678 9698 11734 9754
rect 11536 9556 11592 9612
rect 11678 9556 11734 9612
rect 11536 9414 11592 9470
rect 11678 9414 11734 9470
rect 11536 9272 11592 9328
rect 11678 9272 11734 9328
rect 11536 9130 11592 9186
rect 11678 9130 11734 9186
rect 11536 8988 11592 9044
rect 11678 8988 11734 9044
rect 11536 8846 11592 8902
rect 11678 8846 11734 8902
rect 11536 8704 11592 8760
rect 11678 8704 11734 8760
rect 11536 8562 11592 8618
rect 11678 8562 11734 8618
rect 11536 8420 11592 8476
rect 11678 8420 11734 8476
rect 11536 8278 11592 8334
rect 11678 8278 11734 8334
rect 11536 8136 11592 8192
rect 11678 8136 11734 8192
rect 11536 7994 11592 8050
rect 11678 7994 11734 8050
rect 11536 7852 11592 7908
rect 11678 7852 11734 7908
rect 11536 7710 11592 7766
rect 11678 7710 11734 7766
rect 11536 7568 11592 7624
rect 11678 7568 11734 7624
rect 11536 7426 11592 7482
rect 11678 7426 11734 7482
rect 11536 7284 11592 7340
rect 11678 7284 11734 7340
rect 11536 7142 11592 7198
rect 11678 7142 11734 7198
rect 11536 7000 11592 7056
rect 11678 7000 11734 7056
rect 11536 6858 11592 6914
rect 11678 6858 11734 6914
rect 11536 6716 11592 6772
rect 11678 6716 11734 6772
rect 11536 6574 11592 6630
rect 11678 6574 11734 6630
rect 11536 6432 11592 6488
rect 11678 6432 11734 6488
rect 11536 6290 11592 6346
rect 11678 6290 11734 6346
rect 11536 6148 11592 6204
rect 11678 6148 11734 6204
rect 11536 6006 11592 6062
rect 11678 6006 11734 6062
rect 11536 5864 11592 5920
rect 11678 5864 11734 5920
rect 11536 5722 11592 5778
rect 11678 5722 11734 5778
rect 11536 5580 11592 5636
rect 11678 5580 11734 5636
rect 11536 5438 11592 5494
rect 11678 5438 11734 5494
rect 11536 5296 11592 5352
rect 11678 5296 11734 5352
rect 11536 5154 11592 5210
rect 11678 5154 11734 5210
rect 11536 5012 11592 5068
rect 11678 5012 11734 5068
rect 11536 4870 11592 4926
rect 11678 4870 11734 4926
rect 11536 4728 11592 4784
rect 11678 4728 11734 4784
rect 11536 4586 11592 4642
rect 11678 4586 11734 4642
rect 11536 4444 11592 4500
rect 11678 4444 11734 4500
rect 11536 4302 11592 4358
rect 11678 4302 11734 4358
rect 11536 4160 11592 4216
rect 11678 4160 11734 4216
rect 11536 4018 11592 4074
rect 11678 4018 11734 4074
rect 11536 3876 11592 3932
rect 11678 3876 11734 3932
rect 11536 3734 11592 3790
rect 11678 3734 11734 3790
rect 11536 3592 11592 3648
rect 11678 3592 11734 3648
rect 11536 3450 11592 3506
rect 11678 3450 11734 3506
rect 11536 3308 11592 3364
rect 11678 3308 11734 3364
rect 11536 3166 11592 3222
rect 11678 3166 11734 3222
rect 11536 3024 11592 3080
rect 11678 3024 11734 3080
rect 11536 2882 11592 2938
rect 11678 2882 11734 2938
rect 11536 2740 11592 2796
rect 11678 2740 11734 2796
rect 11536 2598 11592 2654
rect 11678 2598 11734 2654
rect 11536 2456 11592 2512
rect 11678 2456 11734 2512
rect 11536 2314 11592 2370
rect 11678 2314 11734 2370
rect 11536 2172 11592 2228
rect 11678 2172 11734 2228
rect 11536 2030 11592 2086
rect 11678 2030 11734 2086
rect 11536 1888 11592 1944
rect 11678 1888 11734 1944
rect 11536 1746 11592 1802
rect 11678 1746 11734 1802
rect 11536 1604 11592 1660
rect 11678 1604 11734 1660
rect 11536 1462 11592 1518
rect 11678 1462 11734 1518
rect 11536 1320 11592 1376
rect 11678 1320 11734 1376
rect 11536 1178 11592 1234
rect 11678 1178 11734 1234
rect 11536 1036 11592 1092
rect 11678 1036 11734 1092
rect 11536 894 11592 950
rect 11678 894 11734 950
rect 11536 752 11592 808
rect 11678 752 11734 808
rect 11536 610 11592 666
rect 11678 610 11734 666
rect 11536 468 11592 524
rect 11678 468 11734 524
rect 11941 12254 11997 12310
rect 12083 12254 12139 12310
rect 11941 12112 11997 12168
rect 12083 12112 12139 12168
rect 11941 11970 11997 12026
rect 12083 11970 12139 12026
rect 11941 11828 11997 11884
rect 12083 11828 12139 11884
rect 11941 11686 11997 11742
rect 12083 11686 12139 11742
rect 11941 11544 11997 11600
rect 12083 11544 12139 11600
rect 11941 11402 11997 11458
rect 12083 11402 12139 11458
rect 11941 11260 11997 11316
rect 12083 11260 12139 11316
rect 11941 11118 11997 11174
rect 12083 11118 12139 11174
rect 11941 10976 11997 11032
rect 12083 10976 12139 11032
rect 11941 10834 11997 10890
rect 12083 10834 12139 10890
rect 11941 10692 11997 10748
rect 12083 10692 12139 10748
rect 11941 10550 11997 10606
rect 12083 10550 12139 10606
rect 11941 10408 11997 10464
rect 12083 10408 12139 10464
rect 11941 10266 11997 10322
rect 12083 10266 12139 10322
rect 11941 10124 11997 10180
rect 12083 10124 12139 10180
rect 11941 9982 11997 10038
rect 12083 9982 12139 10038
rect 11941 9840 11997 9896
rect 12083 9840 12139 9896
rect 11941 9698 11997 9754
rect 12083 9698 12139 9754
rect 11941 9556 11997 9612
rect 12083 9556 12139 9612
rect 11941 9414 11997 9470
rect 12083 9414 12139 9470
rect 11941 9272 11997 9328
rect 12083 9272 12139 9328
rect 11941 9130 11997 9186
rect 12083 9130 12139 9186
rect 11941 8988 11997 9044
rect 12083 8988 12139 9044
rect 11941 8846 11997 8902
rect 12083 8846 12139 8902
rect 11941 8704 11997 8760
rect 12083 8704 12139 8760
rect 11941 8562 11997 8618
rect 12083 8562 12139 8618
rect 11941 8420 11997 8476
rect 12083 8420 12139 8476
rect 11941 8278 11997 8334
rect 12083 8278 12139 8334
rect 11941 8136 11997 8192
rect 12083 8136 12139 8192
rect 11941 7994 11997 8050
rect 12083 7994 12139 8050
rect 11941 7852 11997 7908
rect 12083 7852 12139 7908
rect 11941 7710 11997 7766
rect 12083 7710 12139 7766
rect 11941 7568 11997 7624
rect 12083 7568 12139 7624
rect 11941 7426 11997 7482
rect 12083 7426 12139 7482
rect 11941 7284 11997 7340
rect 12083 7284 12139 7340
rect 11941 7142 11997 7198
rect 12083 7142 12139 7198
rect 11941 7000 11997 7056
rect 12083 7000 12139 7056
rect 11941 6858 11997 6914
rect 12083 6858 12139 6914
rect 11941 6716 11997 6772
rect 12083 6716 12139 6772
rect 11941 6574 11997 6630
rect 12083 6574 12139 6630
rect 11941 6432 11997 6488
rect 12083 6432 12139 6488
rect 11941 6290 11997 6346
rect 12083 6290 12139 6346
rect 11941 6148 11997 6204
rect 12083 6148 12139 6204
rect 11941 6006 11997 6062
rect 12083 6006 12139 6062
rect 11941 5864 11997 5920
rect 12083 5864 12139 5920
rect 11941 5722 11997 5778
rect 12083 5722 12139 5778
rect 11941 5580 11997 5636
rect 12083 5580 12139 5636
rect 11941 5438 11997 5494
rect 12083 5438 12139 5494
rect 11941 5296 11997 5352
rect 12083 5296 12139 5352
rect 11941 5154 11997 5210
rect 12083 5154 12139 5210
rect 11941 5012 11997 5068
rect 12083 5012 12139 5068
rect 11941 4870 11997 4926
rect 12083 4870 12139 4926
rect 11941 4728 11997 4784
rect 12083 4728 12139 4784
rect 11941 4586 11997 4642
rect 12083 4586 12139 4642
rect 11941 4444 11997 4500
rect 12083 4444 12139 4500
rect 11941 4302 11997 4358
rect 12083 4302 12139 4358
rect 11941 4160 11997 4216
rect 12083 4160 12139 4216
rect 11941 4018 11997 4074
rect 12083 4018 12139 4074
rect 11941 3876 11997 3932
rect 12083 3876 12139 3932
rect 11941 3734 11997 3790
rect 12083 3734 12139 3790
rect 11941 3592 11997 3648
rect 12083 3592 12139 3648
rect 11941 3450 11997 3506
rect 12083 3450 12139 3506
rect 11941 3308 11997 3364
rect 12083 3308 12139 3364
rect 11941 3166 11997 3222
rect 12083 3166 12139 3222
rect 11941 3024 11997 3080
rect 12083 3024 12139 3080
rect 11941 2882 11997 2938
rect 12083 2882 12139 2938
rect 11941 2740 11997 2796
rect 12083 2740 12139 2796
rect 11941 2598 11997 2654
rect 12083 2598 12139 2654
rect 11941 2456 11997 2512
rect 12083 2456 12139 2512
rect 11941 2314 11997 2370
rect 12083 2314 12139 2370
rect 11941 2172 11997 2228
rect 12083 2172 12139 2228
rect 11941 2030 11997 2086
rect 12083 2030 12139 2086
rect 11941 1888 11997 1944
rect 12083 1888 12139 1944
rect 11941 1746 11997 1802
rect 12083 1746 12139 1802
rect 11941 1604 11997 1660
rect 12083 1604 12139 1660
rect 11941 1462 11997 1518
rect 12083 1462 12139 1518
rect 11941 1320 11997 1376
rect 12083 1320 12139 1376
rect 11941 1178 11997 1234
rect 12083 1178 12139 1234
rect 11941 1036 11997 1092
rect 12083 1036 12139 1092
rect 11941 894 11997 950
rect 12083 894 12139 950
rect 11941 752 11997 808
rect 12083 752 12139 808
rect 11941 610 11997 666
rect 12083 610 12139 666
rect 11941 468 11997 524
rect 12083 468 12139 524
rect 12526 12302 12582 12358
rect 12650 12302 12706 12358
rect 12774 12302 12830 12358
rect 12898 12302 12954 12358
rect 13022 12302 13078 12358
rect 12526 12178 12582 12234
rect 12650 12178 12706 12234
rect 12774 12178 12830 12234
rect 12898 12178 12954 12234
rect 13022 12178 13078 12234
rect 12526 12054 12582 12110
rect 12650 12054 12706 12110
rect 12774 12054 12830 12110
rect 12898 12054 12954 12110
rect 13022 12054 13078 12110
rect 12526 11930 12582 11986
rect 12650 11930 12706 11986
rect 12774 11930 12830 11986
rect 12898 11930 12954 11986
rect 13022 11930 13078 11986
rect 12526 11806 12582 11862
rect 12650 11806 12706 11862
rect 12774 11806 12830 11862
rect 12898 11806 12954 11862
rect 13022 11806 13078 11862
rect 12526 11682 12582 11738
rect 12650 11682 12706 11738
rect 12774 11682 12830 11738
rect 12898 11682 12954 11738
rect 13022 11682 13078 11738
rect 12526 11558 12582 11614
rect 12650 11558 12706 11614
rect 12774 11558 12830 11614
rect 12898 11558 12954 11614
rect 13022 11558 13078 11614
rect 12526 11434 12582 11490
rect 12650 11434 12706 11490
rect 12774 11434 12830 11490
rect 12898 11434 12954 11490
rect 13022 11434 13078 11490
rect 12526 11310 12582 11366
rect 12650 11310 12706 11366
rect 12774 11310 12830 11366
rect 12898 11310 12954 11366
rect 13022 11310 13078 11366
rect 12526 11186 12582 11242
rect 12650 11186 12706 11242
rect 12774 11186 12830 11242
rect 12898 11186 12954 11242
rect 13022 11186 13078 11242
rect 12526 11062 12582 11118
rect 12650 11062 12706 11118
rect 12774 11062 12830 11118
rect 12898 11062 12954 11118
rect 13022 11062 13078 11118
rect 12526 10938 12582 10994
rect 12650 10938 12706 10994
rect 12774 10938 12830 10994
rect 12898 10938 12954 10994
rect 13022 10938 13078 10994
rect 12526 10814 12582 10870
rect 12650 10814 12706 10870
rect 12774 10814 12830 10870
rect 12898 10814 12954 10870
rect 13022 10814 13078 10870
rect 12526 10690 12582 10746
rect 12650 10690 12706 10746
rect 12774 10690 12830 10746
rect 12898 10690 12954 10746
rect 13022 10690 13078 10746
rect 12526 10566 12582 10622
rect 12650 10566 12706 10622
rect 12774 10566 12830 10622
rect 12898 10566 12954 10622
rect 13022 10566 13078 10622
rect 12526 10442 12582 10498
rect 12650 10442 12706 10498
rect 12774 10442 12830 10498
rect 12898 10442 12954 10498
rect 13022 10442 13078 10498
rect 12526 10318 12582 10374
rect 12650 10318 12706 10374
rect 12774 10318 12830 10374
rect 12898 10318 12954 10374
rect 13022 10318 13078 10374
rect 12526 10194 12582 10250
rect 12650 10194 12706 10250
rect 12774 10194 12830 10250
rect 12898 10194 12954 10250
rect 13022 10194 13078 10250
rect 12526 10070 12582 10126
rect 12650 10070 12706 10126
rect 12774 10070 12830 10126
rect 12898 10070 12954 10126
rect 13022 10070 13078 10126
rect 12526 9946 12582 10002
rect 12650 9946 12706 10002
rect 12774 9946 12830 10002
rect 12898 9946 12954 10002
rect 13022 9946 13078 10002
rect 12526 9822 12582 9878
rect 12650 9822 12706 9878
rect 12774 9822 12830 9878
rect 12898 9822 12954 9878
rect 13022 9822 13078 9878
rect 12526 9698 12582 9754
rect 12650 9698 12706 9754
rect 12774 9698 12830 9754
rect 12898 9698 12954 9754
rect 13022 9698 13078 9754
rect 12526 9574 12582 9630
rect 12650 9574 12706 9630
rect 12774 9574 12830 9630
rect 12898 9574 12954 9630
rect 13022 9574 13078 9630
rect 12526 9450 12582 9506
rect 12650 9450 12706 9506
rect 12774 9450 12830 9506
rect 12898 9450 12954 9506
rect 13022 9450 13078 9506
rect 12526 9326 12582 9382
rect 12650 9326 12706 9382
rect 12774 9326 12830 9382
rect 12898 9326 12954 9382
rect 13022 9326 13078 9382
rect 12526 9202 12582 9258
rect 12650 9202 12706 9258
rect 12774 9202 12830 9258
rect 12898 9202 12954 9258
rect 13022 9202 13078 9258
rect 12526 9078 12582 9134
rect 12650 9078 12706 9134
rect 12774 9078 12830 9134
rect 12898 9078 12954 9134
rect 13022 9078 13078 9134
rect 12526 8954 12582 9010
rect 12650 8954 12706 9010
rect 12774 8954 12830 9010
rect 12898 8954 12954 9010
rect 13022 8954 13078 9010
rect 12526 8830 12582 8886
rect 12650 8830 12706 8886
rect 12774 8830 12830 8886
rect 12898 8830 12954 8886
rect 13022 8830 13078 8886
rect 12526 8706 12582 8762
rect 12650 8706 12706 8762
rect 12774 8706 12830 8762
rect 12898 8706 12954 8762
rect 13022 8706 13078 8762
rect 12526 8582 12582 8638
rect 12650 8582 12706 8638
rect 12774 8582 12830 8638
rect 12898 8582 12954 8638
rect 13022 8582 13078 8638
rect 12526 8458 12582 8514
rect 12650 8458 12706 8514
rect 12774 8458 12830 8514
rect 12898 8458 12954 8514
rect 13022 8458 13078 8514
rect 12526 8334 12582 8390
rect 12650 8334 12706 8390
rect 12774 8334 12830 8390
rect 12898 8334 12954 8390
rect 13022 8334 13078 8390
rect 12526 8210 12582 8266
rect 12650 8210 12706 8266
rect 12774 8210 12830 8266
rect 12898 8210 12954 8266
rect 13022 8210 13078 8266
rect 12526 8086 12582 8142
rect 12650 8086 12706 8142
rect 12774 8086 12830 8142
rect 12898 8086 12954 8142
rect 13022 8086 13078 8142
rect 12526 7962 12582 8018
rect 12650 7962 12706 8018
rect 12774 7962 12830 8018
rect 12898 7962 12954 8018
rect 13022 7962 13078 8018
rect 12526 7838 12582 7894
rect 12650 7838 12706 7894
rect 12774 7838 12830 7894
rect 12898 7838 12954 7894
rect 13022 7838 13078 7894
rect 12526 7714 12582 7770
rect 12650 7714 12706 7770
rect 12774 7714 12830 7770
rect 12898 7714 12954 7770
rect 13022 7714 13078 7770
rect 12526 7590 12582 7646
rect 12650 7590 12706 7646
rect 12774 7590 12830 7646
rect 12898 7590 12954 7646
rect 13022 7590 13078 7646
rect 12526 7466 12582 7522
rect 12650 7466 12706 7522
rect 12774 7466 12830 7522
rect 12898 7466 12954 7522
rect 13022 7466 13078 7522
rect 12526 7342 12582 7398
rect 12650 7342 12706 7398
rect 12774 7342 12830 7398
rect 12898 7342 12954 7398
rect 13022 7342 13078 7398
rect 12526 7218 12582 7274
rect 12650 7218 12706 7274
rect 12774 7218 12830 7274
rect 12898 7218 12954 7274
rect 13022 7218 13078 7274
rect 12526 7094 12582 7150
rect 12650 7094 12706 7150
rect 12774 7094 12830 7150
rect 12898 7094 12954 7150
rect 13022 7094 13078 7150
rect 12526 6970 12582 7026
rect 12650 6970 12706 7026
rect 12774 6970 12830 7026
rect 12898 6970 12954 7026
rect 13022 6970 13078 7026
rect 12526 6846 12582 6902
rect 12650 6846 12706 6902
rect 12774 6846 12830 6902
rect 12898 6846 12954 6902
rect 13022 6846 13078 6902
rect 12526 6722 12582 6778
rect 12650 6722 12706 6778
rect 12774 6722 12830 6778
rect 12898 6722 12954 6778
rect 13022 6722 13078 6778
rect 12526 6598 12582 6654
rect 12650 6598 12706 6654
rect 12774 6598 12830 6654
rect 12898 6598 12954 6654
rect 13022 6598 13078 6654
rect 12526 6474 12582 6530
rect 12650 6474 12706 6530
rect 12774 6474 12830 6530
rect 12898 6474 12954 6530
rect 13022 6474 13078 6530
rect 12526 6350 12582 6406
rect 12650 6350 12706 6406
rect 12774 6350 12830 6406
rect 12898 6350 12954 6406
rect 13022 6350 13078 6406
rect 12526 6226 12582 6282
rect 12650 6226 12706 6282
rect 12774 6226 12830 6282
rect 12898 6226 12954 6282
rect 13022 6226 13078 6282
rect 12526 6102 12582 6158
rect 12650 6102 12706 6158
rect 12774 6102 12830 6158
rect 12898 6102 12954 6158
rect 13022 6102 13078 6158
rect 12526 5978 12582 6034
rect 12650 5978 12706 6034
rect 12774 5978 12830 6034
rect 12898 5978 12954 6034
rect 13022 5978 13078 6034
rect 12526 5854 12582 5910
rect 12650 5854 12706 5910
rect 12774 5854 12830 5910
rect 12898 5854 12954 5910
rect 13022 5854 13078 5910
rect 12526 5730 12582 5786
rect 12650 5730 12706 5786
rect 12774 5730 12830 5786
rect 12898 5730 12954 5786
rect 13022 5730 13078 5786
rect 12526 5606 12582 5662
rect 12650 5606 12706 5662
rect 12774 5606 12830 5662
rect 12898 5606 12954 5662
rect 13022 5606 13078 5662
rect 12526 5482 12582 5538
rect 12650 5482 12706 5538
rect 12774 5482 12830 5538
rect 12898 5482 12954 5538
rect 13022 5482 13078 5538
rect 12526 5358 12582 5414
rect 12650 5358 12706 5414
rect 12774 5358 12830 5414
rect 12898 5358 12954 5414
rect 13022 5358 13078 5414
rect 12526 5234 12582 5290
rect 12650 5234 12706 5290
rect 12774 5234 12830 5290
rect 12898 5234 12954 5290
rect 13022 5234 13078 5290
rect 12526 5110 12582 5166
rect 12650 5110 12706 5166
rect 12774 5110 12830 5166
rect 12898 5110 12954 5166
rect 13022 5110 13078 5166
rect 12526 4986 12582 5042
rect 12650 4986 12706 5042
rect 12774 4986 12830 5042
rect 12898 4986 12954 5042
rect 13022 4986 13078 5042
rect 12526 4862 12582 4918
rect 12650 4862 12706 4918
rect 12774 4862 12830 4918
rect 12898 4862 12954 4918
rect 13022 4862 13078 4918
rect 12526 4738 12582 4794
rect 12650 4738 12706 4794
rect 12774 4738 12830 4794
rect 12898 4738 12954 4794
rect 13022 4738 13078 4794
rect 12526 4614 12582 4670
rect 12650 4614 12706 4670
rect 12774 4614 12830 4670
rect 12898 4614 12954 4670
rect 13022 4614 13078 4670
rect 12526 4490 12582 4546
rect 12650 4490 12706 4546
rect 12774 4490 12830 4546
rect 12898 4490 12954 4546
rect 13022 4490 13078 4546
rect 12526 4366 12582 4422
rect 12650 4366 12706 4422
rect 12774 4366 12830 4422
rect 12898 4366 12954 4422
rect 13022 4366 13078 4422
rect 12526 4242 12582 4298
rect 12650 4242 12706 4298
rect 12774 4242 12830 4298
rect 12898 4242 12954 4298
rect 13022 4242 13078 4298
rect 12526 4118 12582 4174
rect 12650 4118 12706 4174
rect 12774 4118 12830 4174
rect 12898 4118 12954 4174
rect 13022 4118 13078 4174
rect 12526 3994 12582 4050
rect 12650 3994 12706 4050
rect 12774 3994 12830 4050
rect 12898 3994 12954 4050
rect 13022 3994 13078 4050
rect 12526 3870 12582 3926
rect 12650 3870 12706 3926
rect 12774 3870 12830 3926
rect 12898 3870 12954 3926
rect 13022 3870 13078 3926
rect 12526 3746 12582 3802
rect 12650 3746 12706 3802
rect 12774 3746 12830 3802
rect 12898 3746 12954 3802
rect 13022 3746 13078 3802
rect 12526 3622 12582 3678
rect 12650 3622 12706 3678
rect 12774 3622 12830 3678
rect 12898 3622 12954 3678
rect 13022 3622 13078 3678
rect 12526 3498 12582 3554
rect 12650 3498 12706 3554
rect 12774 3498 12830 3554
rect 12898 3498 12954 3554
rect 13022 3498 13078 3554
rect 12526 3374 12582 3430
rect 12650 3374 12706 3430
rect 12774 3374 12830 3430
rect 12898 3374 12954 3430
rect 13022 3374 13078 3430
rect 12526 3250 12582 3306
rect 12650 3250 12706 3306
rect 12774 3250 12830 3306
rect 12898 3250 12954 3306
rect 13022 3250 13078 3306
rect 12526 3126 12582 3182
rect 12650 3126 12706 3182
rect 12774 3126 12830 3182
rect 12898 3126 12954 3182
rect 13022 3126 13078 3182
rect 12526 3002 12582 3058
rect 12650 3002 12706 3058
rect 12774 3002 12830 3058
rect 12898 3002 12954 3058
rect 13022 3002 13078 3058
rect 12526 2878 12582 2934
rect 12650 2878 12706 2934
rect 12774 2878 12830 2934
rect 12898 2878 12954 2934
rect 13022 2878 13078 2934
rect 12526 2754 12582 2810
rect 12650 2754 12706 2810
rect 12774 2754 12830 2810
rect 12898 2754 12954 2810
rect 13022 2754 13078 2810
rect 12526 2630 12582 2686
rect 12650 2630 12706 2686
rect 12774 2630 12830 2686
rect 12898 2630 12954 2686
rect 13022 2630 13078 2686
rect 12526 2506 12582 2562
rect 12650 2506 12706 2562
rect 12774 2506 12830 2562
rect 12898 2506 12954 2562
rect 13022 2506 13078 2562
rect 12526 2382 12582 2438
rect 12650 2382 12706 2438
rect 12774 2382 12830 2438
rect 12898 2382 12954 2438
rect 13022 2382 13078 2438
rect 12526 2258 12582 2314
rect 12650 2258 12706 2314
rect 12774 2258 12830 2314
rect 12898 2258 12954 2314
rect 13022 2258 13078 2314
rect 12526 2134 12582 2190
rect 12650 2134 12706 2190
rect 12774 2134 12830 2190
rect 12898 2134 12954 2190
rect 13022 2134 13078 2190
rect 12526 2010 12582 2066
rect 12650 2010 12706 2066
rect 12774 2010 12830 2066
rect 12898 2010 12954 2066
rect 13022 2010 13078 2066
rect 12526 1886 12582 1942
rect 12650 1886 12706 1942
rect 12774 1886 12830 1942
rect 12898 1886 12954 1942
rect 13022 1886 13078 1942
rect 12526 1762 12582 1818
rect 12650 1762 12706 1818
rect 12774 1762 12830 1818
rect 12898 1762 12954 1818
rect 13022 1762 13078 1818
rect 12526 1638 12582 1694
rect 12650 1638 12706 1694
rect 12774 1638 12830 1694
rect 12898 1638 12954 1694
rect 13022 1638 13078 1694
rect 12526 1514 12582 1570
rect 12650 1514 12706 1570
rect 12774 1514 12830 1570
rect 12898 1514 12954 1570
rect 13022 1514 13078 1570
rect 12526 1390 12582 1446
rect 12650 1390 12706 1446
rect 12774 1390 12830 1446
rect 12898 1390 12954 1446
rect 13022 1390 13078 1446
rect 12526 1266 12582 1322
rect 12650 1266 12706 1322
rect 12774 1266 12830 1322
rect 12898 1266 12954 1322
rect 13022 1266 13078 1322
rect 12526 1142 12582 1198
rect 12650 1142 12706 1198
rect 12774 1142 12830 1198
rect 12898 1142 12954 1198
rect 13022 1142 13078 1198
rect 12526 1018 12582 1074
rect 12650 1018 12706 1074
rect 12774 1018 12830 1074
rect 12898 1018 12954 1074
rect 13022 1018 13078 1074
rect 12526 894 12582 950
rect 12650 894 12706 950
rect 12774 894 12830 950
rect 12898 894 12954 950
rect 13022 894 13078 950
rect 12526 770 12582 826
rect 12650 770 12706 826
rect 12774 770 12830 826
rect 12898 770 12954 826
rect 13022 770 13078 826
rect 12526 646 12582 702
rect 12650 646 12706 702
rect 12774 646 12830 702
rect 12898 646 12954 702
rect 13022 646 13078 702
rect 12526 522 12582 578
rect 12650 522 12706 578
rect 12774 522 12830 578
rect 12898 522 12954 578
rect 13022 522 13078 578
rect 12526 398 12582 454
rect 12650 398 12706 454
rect 12774 398 12830 454
rect 12898 398 12954 454
rect 13022 398 13078 454
rect -286 274 -230 330
rect -162 274 -106 330
rect -38 274 18 330
rect 86 274 142 330
rect 210 274 266 330
rect 415 246 471 302
rect 557 246 613 302
rect 699 246 755 302
rect 841 246 897 302
rect 983 246 1039 302
rect 1125 246 1181 302
rect 1267 246 1323 302
rect 1409 246 1465 302
rect 1551 246 1607 302
rect 1693 246 1749 302
rect 1835 246 1891 302
rect 1977 246 2033 302
rect 2119 246 2175 302
rect 2261 246 2317 302
rect 2403 246 2459 302
rect 2545 246 2601 302
rect 2687 246 2743 302
rect 2829 246 2885 302
rect 2971 246 3027 302
rect 3113 246 3169 302
rect 3255 246 3311 302
rect 3397 246 3453 302
rect 3539 246 3595 302
rect 3681 246 3737 302
rect 3823 246 3879 302
rect 3965 246 4021 302
rect 4107 246 4163 302
rect 4249 246 4305 302
rect 4391 246 4447 302
rect 4533 246 4589 302
rect 4675 246 4731 302
rect 4817 246 4873 302
rect 4959 246 5015 302
rect 5101 246 5157 302
rect 5243 246 5299 302
rect 5385 246 5441 302
rect 5527 246 5583 302
rect 5669 246 5725 302
rect 5811 246 5867 302
rect 5953 246 6009 302
rect 6095 246 6151 302
rect 6237 246 6293 302
rect 6379 246 6435 302
rect 6521 246 6577 302
rect 6663 246 6719 302
rect 6805 246 6861 302
rect 6947 246 7003 302
rect 7089 246 7145 302
rect 7231 246 7287 302
rect 7373 246 7429 302
rect 7515 246 7571 302
rect 7657 246 7713 302
rect 7799 246 7855 302
rect 7941 246 7997 302
rect 8083 246 8139 302
rect 8225 246 8281 302
rect 8367 246 8423 302
rect 8509 246 8565 302
rect 8651 246 8707 302
rect 8793 246 8849 302
rect 8935 246 8991 302
rect 9077 246 9133 302
rect 9219 246 9275 302
rect 9361 246 9417 302
rect 9503 246 9559 302
rect 9645 246 9701 302
rect 9787 246 9843 302
rect 9929 246 9985 302
rect 10071 246 10127 302
rect 10213 246 10269 302
rect 10355 246 10411 302
rect 10497 246 10553 302
rect 10639 246 10695 302
rect 10781 246 10837 302
rect 10923 246 10979 302
rect 11065 246 11121 302
rect 11207 246 11263 302
rect 11349 246 11405 302
rect 11491 246 11547 302
rect 11633 246 11689 302
rect 11775 246 11831 302
rect 11917 246 11973 302
rect 12059 246 12115 302
rect 12201 246 12257 302
rect 12343 246 12399 302
rect 12526 274 12582 330
rect 12650 274 12706 330
rect 12774 274 12830 330
rect 12898 274 12954 330
rect 13022 274 13078 330
rect -286 150 -230 206
rect -162 150 -106 206
rect -38 150 18 206
rect 86 150 142 206
rect 210 150 266 206
rect 415 104 471 160
rect 557 104 613 160
rect 699 104 755 160
rect 841 104 897 160
rect 983 104 1039 160
rect 1125 104 1181 160
rect 1267 104 1323 160
rect 1409 104 1465 160
rect 1551 104 1607 160
rect 1693 104 1749 160
rect 1835 104 1891 160
rect 1977 104 2033 160
rect 2119 104 2175 160
rect 2261 104 2317 160
rect 2403 104 2459 160
rect 2545 104 2601 160
rect 2687 104 2743 160
rect 2829 104 2885 160
rect 2971 104 3027 160
rect 3113 104 3169 160
rect 3255 104 3311 160
rect 3397 104 3453 160
rect 3539 104 3595 160
rect 3681 104 3737 160
rect 3823 104 3879 160
rect 3965 104 4021 160
rect 4107 104 4163 160
rect 4249 104 4305 160
rect 4391 104 4447 160
rect 4533 104 4589 160
rect 4675 104 4731 160
rect 4817 104 4873 160
rect 4959 104 5015 160
rect 5101 104 5157 160
rect 5243 104 5299 160
rect 5385 104 5441 160
rect 5527 104 5583 160
rect 5669 104 5725 160
rect 5811 104 5867 160
rect 5953 104 6009 160
rect 6095 104 6151 160
rect 6237 104 6293 160
rect 6379 104 6435 160
rect 6521 104 6577 160
rect 6663 104 6719 160
rect 6805 104 6861 160
rect 6947 104 7003 160
rect 7089 104 7145 160
rect 7231 104 7287 160
rect 7373 104 7429 160
rect 7515 104 7571 160
rect 7657 104 7713 160
rect 7799 104 7855 160
rect 7941 104 7997 160
rect 8083 104 8139 160
rect 8225 104 8281 160
rect 8367 104 8423 160
rect 8509 104 8565 160
rect 8651 104 8707 160
rect 8793 104 8849 160
rect 8935 104 8991 160
rect 9077 104 9133 160
rect 9219 104 9275 160
rect 9361 104 9417 160
rect 9503 104 9559 160
rect 9645 104 9701 160
rect 9787 104 9843 160
rect 9929 104 9985 160
rect 10071 104 10127 160
rect 10213 104 10269 160
rect 10355 104 10411 160
rect 10497 104 10553 160
rect 10639 104 10695 160
rect 10781 104 10837 160
rect 10923 104 10979 160
rect 11065 104 11121 160
rect 11207 104 11263 160
rect 11349 104 11405 160
rect 11491 104 11547 160
rect 11633 104 11689 160
rect 11775 104 11831 160
rect 11917 104 11973 160
rect 12059 104 12115 160
rect 12201 104 12257 160
rect 12343 104 12399 160
rect 12526 150 12582 206
rect 12650 150 12706 206
rect 12774 150 12830 206
rect 12898 150 12954 206
rect 13022 150 13078 206
<< metal4 >>
rect -400 12949 13200 13065
rect -400 12893 -254 12949
rect -198 12893 -130 12949
rect -74 12893 -6 12949
rect 50 12893 118 12949
rect 174 12893 242 12949
rect 298 12893 366 12949
rect 422 12893 490 12949
rect 546 12893 614 12949
rect 670 12893 738 12949
rect 794 12893 862 12949
rect 918 12893 986 12949
rect 1042 12893 1110 12949
rect 1166 12893 1234 12949
rect 1290 12893 1358 12949
rect 1414 12893 1482 12949
rect 1538 12893 1606 12949
rect 1662 12893 1730 12949
rect 1786 12893 1854 12949
rect 1910 12893 1978 12949
rect 2034 12893 2102 12949
rect 2158 12893 2226 12949
rect 2282 12893 2350 12949
rect 2406 12893 2474 12949
rect 2530 12893 2598 12949
rect 2654 12893 2722 12949
rect 2778 12893 2846 12949
rect 2902 12893 2970 12949
rect 3026 12893 3094 12949
rect 3150 12893 3218 12949
rect 3274 12893 3342 12949
rect 3398 12893 3466 12949
rect 3522 12893 3590 12949
rect 3646 12893 3714 12949
rect 3770 12893 3838 12949
rect 3894 12893 3962 12949
rect 4018 12893 4086 12949
rect 4142 12893 4210 12949
rect 4266 12893 4334 12949
rect 4390 12893 4458 12949
rect 4514 12893 4582 12949
rect 4638 12893 4706 12949
rect 4762 12893 4830 12949
rect 4886 12893 4954 12949
rect 5010 12893 5078 12949
rect 5134 12893 5202 12949
rect 5258 12893 5326 12949
rect 5382 12893 5450 12949
rect 5506 12893 5574 12949
rect 5630 12893 5698 12949
rect 5754 12893 5822 12949
rect 5878 12893 5946 12949
rect 6002 12893 6070 12949
rect 6126 12893 6194 12949
rect 6250 12893 6318 12949
rect 6374 12893 6442 12949
rect 6498 12893 6566 12949
rect 6622 12893 6690 12949
rect 6746 12893 6814 12949
rect 6870 12893 6938 12949
rect 6994 12893 7062 12949
rect 7118 12893 7186 12949
rect 7242 12893 7310 12949
rect 7366 12893 7434 12949
rect 7490 12893 7558 12949
rect 7614 12893 7682 12949
rect 7738 12893 7806 12949
rect 7862 12893 7930 12949
rect 7986 12893 8054 12949
rect 8110 12893 8178 12949
rect 8234 12893 8302 12949
rect 8358 12893 8426 12949
rect 8482 12893 8550 12949
rect 8606 12893 8674 12949
rect 8730 12893 8798 12949
rect 8854 12893 8922 12949
rect 8978 12893 9046 12949
rect 9102 12893 9170 12949
rect 9226 12893 9294 12949
rect 9350 12893 9418 12949
rect 9474 12893 9542 12949
rect 9598 12893 9666 12949
rect 9722 12893 9790 12949
rect 9846 12893 9914 12949
rect 9970 12893 10038 12949
rect 10094 12893 10162 12949
rect 10218 12893 10286 12949
rect 10342 12893 10410 12949
rect 10466 12893 10534 12949
rect 10590 12893 10658 12949
rect 10714 12893 10782 12949
rect 10838 12893 10906 12949
rect 10962 12893 11030 12949
rect 11086 12893 11154 12949
rect 11210 12893 11278 12949
rect 11334 12893 11402 12949
rect 11458 12893 11526 12949
rect 11582 12893 11650 12949
rect 11706 12893 11774 12949
rect 11830 12893 11898 12949
rect 11954 12893 12022 12949
rect 12078 12893 12146 12949
rect 12202 12893 12270 12949
rect 12326 12893 12394 12949
rect 12450 12893 12518 12949
rect 12574 12893 12642 12949
rect 12698 12893 12766 12949
rect 12822 12893 12890 12949
rect 12946 12893 13014 12949
rect 13070 12893 13200 12949
rect -400 12825 13200 12893
rect -400 12769 -254 12825
rect -198 12769 -130 12825
rect -74 12769 -6 12825
rect 50 12769 118 12825
rect 174 12769 242 12825
rect 298 12769 366 12825
rect 422 12769 490 12825
rect 546 12769 614 12825
rect 670 12769 738 12825
rect 794 12769 862 12825
rect 918 12769 986 12825
rect 1042 12769 1110 12825
rect 1166 12769 1234 12825
rect 1290 12769 1358 12825
rect 1414 12769 1482 12825
rect 1538 12769 1606 12825
rect 1662 12769 1730 12825
rect 1786 12769 1854 12825
rect 1910 12769 1978 12825
rect 2034 12769 2102 12825
rect 2158 12769 2226 12825
rect 2282 12769 2350 12825
rect 2406 12769 2474 12825
rect 2530 12769 2598 12825
rect 2654 12769 2722 12825
rect 2778 12769 2846 12825
rect 2902 12769 2970 12825
rect 3026 12769 3094 12825
rect 3150 12769 3218 12825
rect 3274 12769 3342 12825
rect 3398 12769 3466 12825
rect 3522 12769 3590 12825
rect 3646 12769 3714 12825
rect 3770 12769 3838 12825
rect 3894 12769 3962 12825
rect 4018 12769 4086 12825
rect 4142 12769 4210 12825
rect 4266 12769 4334 12825
rect 4390 12769 4458 12825
rect 4514 12769 4582 12825
rect 4638 12769 4706 12825
rect 4762 12769 4830 12825
rect 4886 12769 4954 12825
rect 5010 12769 5078 12825
rect 5134 12769 5202 12825
rect 5258 12769 5326 12825
rect 5382 12769 5450 12825
rect 5506 12769 5574 12825
rect 5630 12769 5698 12825
rect 5754 12769 5822 12825
rect 5878 12769 5946 12825
rect 6002 12769 6070 12825
rect 6126 12769 6194 12825
rect 6250 12769 6318 12825
rect 6374 12769 6442 12825
rect 6498 12769 6566 12825
rect 6622 12769 6690 12825
rect 6746 12769 6814 12825
rect 6870 12769 6938 12825
rect 6994 12769 7062 12825
rect 7118 12769 7186 12825
rect 7242 12769 7310 12825
rect 7366 12769 7434 12825
rect 7490 12769 7558 12825
rect 7614 12769 7682 12825
rect 7738 12769 7806 12825
rect 7862 12769 7930 12825
rect 7986 12769 8054 12825
rect 8110 12769 8178 12825
rect 8234 12769 8302 12825
rect 8358 12769 8426 12825
rect 8482 12769 8550 12825
rect 8606 12769 8674 12825
rect 8730 12769 8798 12825
rect 8854 12769 8922 12825
rect 8978 12769 9046 12825
rect 9102 12769 9170 12825
rect 9226 12769 9294 12825
rect 9350 12769 9418 12825
rect 9474 12769 9542 12825
rect 9598 12769 9666 12825
rect 9722 12769 9790 12825
rect 9846 12769 9914 12825
rect 9970 12769 10038 12825
rect 10094 12769 10162 12825
rect 10218 12769 10286 12825
rect 10342 12769 10410 12825
rect 10466 12769 10534 12825
rect 10590 12769 10658 12825
rect 10714 12769 10782 12825
rect 10838 12769 10906 12825
rect 10962 12769 11030 12825
rect 11086 12769 11154 12825
rect 11210 12769 11278 12825
rect 11334 12769 11402 12825
rect 11458 12769 11526 12825
rect 11582 12769 11650 12825
rect 11706 12769 11774 12825
rect 11830 12769 11898 12825
rect 11954 12769 12022 12825
rect 12078 12769 12146 12825
rect 12202 12769 12270 12825
rect 12326 12769 12394 12825
rect 12450 12769 12518 12825
rect 12574 12769 12642 12825
rect 12698 12769 12766 12825
rect 12822 12769 12890 12825
rect 12946 12769 13014 12825
rect 13070 12769 13200 12825
rect -400 12701 13200 12769
rect -400 12645 -254 12701
rect -198 12645 -130 12701
rect -74 12645 -6 12701
rect 50 12645 118 12701
rect 174 12645 242 12701
rect 298 12645 366 12701
rect 422 12645 490 12701
rect 546 12645 614 12701
rect 670 12645 738 12701
rect 794 12645 862 12701
rect 918 12645 986 12701
rect 1042 12645 1110 12701
rect 1166 12645 1234 12701
rect 1290 12645 1358 12701
rect 1414 12645 1482 12701
rect 1538 12645 1606 12701
rect 1662 12645 1730 12701
rect 1786 12645 1854 12701
rect 1910 12645 1978 12701
rect 2034 12645 2102 12701
rect 2158 12645 2226 12701
rect 2282 12645 2350 12701
rect 2406 12645 2474 12701
rect 2530 12645 2598 12701
rect 2654 12645 2722 12701
rect 2778 12645 2846 12701
rect 2902 12645 2970 12701
rect 3026 12645 3094 12701
rect 3150 12645 3218 12701
rect 3274 12645 3342 12701
rect 3398 12645 3466 12701
rect 3522 12645 3590 12701
rect 3646 12645 3714 12701
rect 3770 12645 3838 12701
rect 3894 12645 3962 12701
rect 4018 12645 4086 12701
rect 4142 12645 4210 12701
rect 4266 12645 4334 12701
rect 4390 12645 4458 12701
rect 4514 12645 4582 12701
rect 4638 12645 4706 12701
rect 4762 12645 4830 12701
rect 4886 12645 4954 12701
rect 5010 12645 5078 12701
rect 5134 12645 5202 12701
rect 5258 12645 5326 12701
rect 5382 12645 5450 12701
rect 5506 12645 5574 12701
rect 5630 12645 5698 12701
rect 5754 12645 5822 12701
rect 5878 12645 5946 12701
rect 6002 12645 6070 12701
rect 6126 12645 6194 12701
rect 6250 12645 6318 12701
rect 6374 12645 6442 12701
rect 6498 12645 6566 12701
rect 6622 12645 6690 12701
rect 6746 12645 6814 12701
rect 6870 12645 6938 12701
rect 6994 12645 7062 12701
rect 7118 12645 7186 12701
rect 7242 12645 7310 12701
rect 7366 12645 7434 12701
rect 7490 12645 7558 12701
rect 7614 12645 7682 12701
rect 7738 12645 7806 12701
rect 7862 12645 7930 12701
rect 7986 12645 8054 12701
rect 8110 12645 8178 12701
rect 8234 12645 8302 12701
rect 8358 12645 8426 12701
rect 8482 12645 8550 12701
rect 8606 12645 8674 12701
rect 8730 12645 8798 12701
rect 8854 12645 8922 12701
rect 8978 12645 9046 12701
rect 9102 12645 9170 12701
rect 9226 12645 9294 12701
rect 9350 12645 9418 12701
rect 9474 12645 9542 12701
rect 9598 12645 9666 12701
rect 9722 12645 9790 12701
rect 9846 12645 9914 12701
rect 9970 12645 10038 12701
rect 10094 12645 10162 12701
rect 10218 12645 10286 12701
rect 10342 12645 10410 12701
rect 10466 12645 10534 12701
rect 10590 12645 10658 12701
rect 10714 12645 10782 12701
rect 10838 12645 10906 12701
rect 10962 12645 11030 12701
rect 11086 12645 11154 12701
rect 11210 12645 11278 12701
rect 11334 12645 11402 12701
rect 11458 12645 11526 12701
rect 11582 12645 11650 12701
rect 11706 12645 11774 12701
rect 11830 12645 11898 12701
rect 11954 12645 12022 12701
rect 12078 12645 12146 12701
rect 12202 12645 12270 12701
rect 12326 12645 12394 12701
rect 12450 12645 12518 12701
rect 12574 12645 12642 12701
rect 12698 12645 12766 12701
rect 12822 12645 12890 12701
rect 12946 12645 13014 12701
rect 13070 12645 13200 12701
rect -400 12577 13200 12645
rect -400 12521 -254 12577
rect -198 12521 -130 12577
rect -74 12521 -6 12577
rect 50 12521 118 12577
rect 174 12521 242 12577
rect 298 12521 366 12577
rect 422 12521 490 12577
rect 546 12521 614 12577
rect 670 12521 738 12577
rect 794 12521 862 12577
rect 918 12521 986 12577
rect 1042 12521 1110 12577
rect 1166 12521 1234 12577
rect 1290 12521 1358 12577
rect 1414 12521 1482 12577
rect 1538 12521 1606 12577
rect 1662 12521 1730 12577
rect 1786 12521 1854 12577
rect 1910 12521 1978 12577
rect 2034 12521 2102 12577
rect 2158 12521 2226 12577
rect 2282 12521 2350 12577
rect 2406 12521 2474 12577
rect 2530 12521 2598 12577
rect 2654 12521 2722 12577
rect 2778 12521 2846 12577
rect 2902 12521 2970 12577
rect 3026 12521 3094 12577
rect 3150 12521 3218 12577
rect 3274 12521 3342 12577
rect 3398 12521 3466 12577
rect 3522 12521 3590 12577
rect 3646 12521 3714 12577
rect 3770 12521 3838 12577
rect 3894 12521 3962 12577
rect 4018 12521 4086 12577
rect 4142 12521 4210 12577
rect 4266 12521 4334 12577
rect 4390 12521 4458 12577
rect 4514 12521 4582 12577
rect 4638 12521 4706 12577
rect 4762 12521 4830 12577
rect 4886 12521 4954 12577
rect 5010 12521 5078 12577
rect 5134 12521 5202 12577
rect 5258 12521 5326 12577
rect 5382 12521 5450 12577
rect 5506 12521 5574 12577
rect 5630 12521 5698 12577
rect 5754 12521 5822 12577
rect 5878 12521 5946 12577
rect 6002 12521 6070 12577
rect 6126 12521 6194 12577
rect 6250 12521 6318 12577
rect 6374 12521 6442 12577
rect 6498 12521 6566 12577
rect 6622 12521 6690 12577
rect 6746 12521 6814 12577
rect 6870 12521 6938 12577
rect 6994 12521 7062 12577
rect 7118 12521 7186 12577
rect 7242 12521 7310 12577
rect 7366 12521 7434 12577
rect 7490 12521 7558 12577
rect 7614 12521 7682 12577
rect 7738 12521 7806 12577
rect 7862 12521 7930 12577
rect 7986 12521 8054 12577
rect 8110 12521 8178 12577
rect 8234 12521 8302 12577
rect 8358 12521 8426 12577
rect 8482 12521 8550 12577
rect 8606 12521 8674 12577
rect 8730 12521 8798 12577
rect 8854 12521 8922 12577
rect 8978 12521 9046 12577
rect 9102 12521 9170 12577
rect 9226 12521 9294 12577
rect 9350 12521 9418 12577
rect 9474 12521 9542 12577
rect 9598 12521 9666 12577
rect 9722 12521 9790 12577
rect 9846 12521 9914 12577
rect 9970 12521 10038 12577
rect 10094 12521 10162 12577
rect 10218 12521 10286 12577
rect 10342 12521 10410 12577
rect 10466 12521 10534 12577
rect 10590 12521 10658 12577
rect 10714 12521 10782 12577
rect 10838 12521 10906 12577
rect 10962 12521 11030 12577
rect 11086 12521 11154 12577
rect 11210 12521 11278 12577
rect 11334 12521 11402 12577
rect 11458 12521 11526 12577
rect 11582 12521 11650 12577
rect 11706 12521 11774 12577
rect 11830 12521 11898 12577
rect 11954 12521 12022 12577
rect 12078 12521 12146 12577
rect 12202 12521 12270 12577
rect 12326 12521 12394 12577
rect 12450 12521 12518 12577
rect 12574 12521 12642 12577
rect 12698 12521 12766 12577
rect 12822 12521 12890 12577
rect 12946 12521 13014 12577
rect 13070 12521 13200 12577
rect -400 12358 13200 12521
rect -400 12302 -286 12358
rect -230 12302 -162 12358
rect -106 12302 -38 12358
rect 18 12302 86 12358
rect 142 12302 210 12358
rect 266 12310 12526 12358
rect 266 12302 741 12310
rect -400 12254 741 12302
rect 797 12254 883 12310
rect 939 12254 1142 12310
rect 1198 12254 1284 12310
rect 1340 12254 1542 12310
rect 1598 12254 1684 12310
rect 1740 12254 1939 12310
rect 1995 12254 2081 12310
rect 2137 12254 2336 12310
rect 2392 12254 2478 12310
rect 2534 12254 2740 12310
rect 2796 12254 2882 12310
rect 2938 12254 3136 12310
rect 3192 12254 3278 12310
rect 3334 12254 3536 12310
rect 3592 12254 3678 12310
rect 3734 12254 3933 12310
rect 3989 12254 4075 12310
rect 4131 12254 4338 12310
rect 4394 12254 4480 12310
rect 4536 12254 4738 12310
rect 4794 12254 4880 12310
rect 4936 12254 5143 12310
rect 5199 12254 5285 12310
rect 5341 12254 5540 12310
rect 5596 12254 5682 12310
rect 5738 12254 5937 12310
rect 5993 12254 6079 12310
rect 6135 12254 6340 12310
rect 6396 12254 6482 12310
rect 6538 12254 6742 12310
rect 6798 12254 6884 12310
rect 6940 12254 7145 12310
rect 7201 12254 7287 12310
rect 7343 12254 7539 12310
rect 7595 12254 7681 12310
rect 7737 12254 7940 12310
rect 7996 12254 8082 12310
rect 8138 12254 8340 12310
rect 8396 12254 8482 12310
rect 8538 12254 8737 12310
rect 8793 12254 8879 12310
rect 8935 12254 9134 12310
rect 9190 12254 9276 12310
rect 9332 12254 9538 12310
rect 9594 12254 9680 12310
rect 9736 12254 9934 12310
rect 9990 12254 10076 12310
rect 10132 12254 10334 12310
rect 10390 12254 10476 12310
rect 10532 12254 10731 12310
rect 10787 12254 10873 12310
rect 10929 12254 11136 12310
rect 11192 12254 11278 12310
rect 11334 12254 11536 12310
rect 11592 12254 11678 12310
rect 11734 12254 11941 12310
rect 11997 12254 12083 12310
rect 12139 12302 12526 12310
rect 12582 12302 12650 12358
rect 12706 12302 12774 12358
rect 12830 12302 12898 12358
rect 12954 12302 13022 12358
rect 13078 12302 13200 12358
rect 12139 12254 13200 12302
rect -400 12234 13200 12254
rect -400 12178 -286 12234
rect -230 12178 -162 12234
rect -106 12178 -38 12234
rect 18 12178 86 12234
rect 142 12178 210 12234
rect 266 12178 12526 12234
rect 12582 12178 12650 12234
rect 12706 12178 12774 12234
rect 12830 12178 12898 12234
rect 12954 12178 13022 12234
rect 13078 12178 13200 12234
rect -400 12168 13200 12178
rect -400 12112 741 12168
rect 797 12112 883 12168
rect 939 12112 1142 12168
rect 1198 12112 1284 12168
rect 1340 12112 1542 12168
rect 1598 12112 1684 12168
rect 1740 12112 1939 12168
rect 1995 12112 2081 12168
rect 2137 12112 2336 12168
rect 2392 12112 2478 12168
rect 2534 12112 2740 12168
rect 2796 12112 2882 12168
rect 2938 12112 3136 12168
rect 3192 12112 3278 12168
rect 3334 12112 3536 12168
rect 3592 12112 3678 12168
rect 3734 12112 3933 12168
rect 3989 12112 4075 12168
rect 4131 12112 4338 12168
rect 4394 12112 4480 12168
rect 4536 12112 4738 12168
rect 4794 12112 4880 12168
rect 4936 12112 5143 12168
rect 5199 12112 5285 12168
rect 5341 12112 5540 12168
rect 5596 12112 5682 12168
rect 5738 12112 5937 12168
rect 5993 12112 6079 12168
rect 6135 12112 6340 12168
rect 6396 12112 6482 12168
rect 6538 12112 6742 12168
rect 6798 12112 6884 12168
rect 6940 12112 7145 12168
rect 7201 12112 7287 12168
rect 7343 12112 7539 12168
rect 7595 12112 7681 12168
rect 7737 12112 7940 12168
rect 7996 12112 8082 12168
rect 8138 12112 8340 12168
rect 8396 12112 8482 12168
rect 8538 12112 8737 12168
rect 8793 12112 8879 12168
rect 8935 12112 9134 12168
rect 9190 12112 9276 12168
rect 9332 12112 9538 12168
rect 9594 12112 9680 12168
rect 9736 12112 9934 12168
rect 9990 12112 10076 12168
rect 10132 12112 10334 12168
rect 10390 12112 10476 12168
rect 10532 12112 10731 12168
rect 10787 12112 10873 12168
rect 10929 12112 11136 12168
rect 11192 12112 11278 12168
rect 11334 12112 11536 12168
rect 11592 12112 11678 12168
rect 11734 12112 11941 12168
rect 11997 12112 12083 12168
rect 12139 12112 13200 12168
rect -400 12110 13200 12112
rect -400 12054 -286 12110
rect -230 12054 -162 12110
rect -106 12054 -38 12110
rect 18 12054 86 12110
rect 142 12054 210 12110
rect 266 12054 12526 12110
rect 12582 12054 12650 12110
rect 12706 12054 12774 12110
rect 12830 12054 12898 12110
rect 12954 12054 13022 12110
rect 13078 12054 13200 12110
rect -400 12026 13200 12054
rect -400 11986 741 12026
rect -400 11930 -286 11986
rect -230 11930 -162 11986
rect -106 11930 -38 11986
rect 18 11930 86 11986
rect 142 11930 210 11986
rect 266 11970 741 11986
rect 797 11970 883 12026
rect 939 11970 1142 12026
rect 1198 11970 1284 12026
rect 1340 11970 1542 12026
rect 1598 11970 1684 12026
rect 1740 11970 1939 12026
rect 1995 11970 2081 12026
rect 2137 11970 2336 12026
rect 2392 11970 2478 12026
rect 2534 11970 2740 12026
rect 2796 11970 2882 12026
rect 2938 11970 3136 12026
rect 3192 11970 3278 12026
rect 3334 11970 3536 12026
rect 3592 11970 3678 12026
rect 3734 11970 3933 12026
rect 3989 11970 4075 12026
rect 4131 11970 4338 12026
rect 4394 11970 4480 12026
rect 4536 11970 4738 12026
rect 4794 11970 4880 12026
rect 4936 11970 5143 12026
rect 5199 11970 5285 12026
rect 5341 11970 5540 12026
rect 5596 11970 5682 12026
rect 5738 11970 5937 12026
rect 5993 11970 6079 12026
rect 6135 11970 6340 12026
rect 6396 11970 6482 12026
rect 6538 11970 6742 12026
rect 6798 11970 6884 12026
rect 6940 11970 7145 12026
rect 7201 11970 7287 12026
rect 7343 11970 7539 12026
rect 7595 11970 7681 12026
rect 7737 11970 7940 12026
rect 7996 11970 8082 12026
rect 8138 11970 8340 12026
rect 8396 11970 8482 12026
rect 8538 11970 8737 12026
rect 8793 11970 8879 12026
rect 8935 11970 9134 12026
rect 9190 11970 9276 12026
rect 9332 11970 9538 12026
rect 9594 11970 9680 12026
rect 9736 11970 9934 12026
rect 9990 11970 10076 12026
rect 10132 11970 10334 12026
rect 10390 11970 10476 12026
rect 10532 11970 10731 12026
rect 10787 11970 10873 12026
rect 10929 11970 11136 12026
rect 11192 11970 11278 12026
rect 11334 11970 11536 12026
rect 11592 11970 11678 12026
rect 11734 11970 11941 12026
rect 11997 11970 12083 12026
rect 12139 11986 13200 12026
rect 12139 11970 12526 11986
rect 266 11930 12526 11970
rect 12582 11930 12650 11986
rect 12706 11930 12774 11986
rect 12830 11930 12898 11986
rect 12954 11930 13022 11986
rect 13078 11930 13200 11986
rect -400 11884 13200 11930
rect -400 11862 741 11884
rect -400 11806 -286 11862
rect -230 11806 -162 11862
rect -106 11806 -38 11862
rect 18 11806 86 11862
rect 142 11806 210 11862
rect 266 11828 741 11862
rect 797 11828 883 11884
rect 939 11828 1142 11884
rect 1198 11828 1284 11884
rect 1340 11828 1542 11884
rect 1598 11828 1684 11884
rect 1740 11828 1939 11884
rect 1995 11828 2081 11884
rect 2137 11828 2336 11884
rect 2392 11828 2478 11884
rect 2534 11828 2740 11884
rect 2796 11828 2882 11884
rect 2938 11828 3136 11884
rect 3192 11828 3278 11884
rect 3334 11828 3536 11884
rect 3592 11828 3678 11884
rect 3734 11828 3933 11884
rect 3989 11828 4075 11884
rect 4131 11828 4338 11884
rect 4394 11828 4480 11884
rect 4536 11828 4738 11884
rect 4794 11828 4880 11884
rect 4936 11828 5143 11884
rect 5199 11828 5285 11884
rect 5341 11828 5540 11884
rect 5596 11828 5682 11884
rect 5738 11828 5937 11884
rect 5993 11828 6079 11884
rect 6135 11828 6340 11884
rect 6396 11828 6482 11884
rect 6538 11828 6742 11884
rect 6798 11828 6884 11884
rect 6940 11828 7145 11884
rect 7201 11828 7287 11884
rect 7343 11828 7539 11884
rect 7595 11828 7681 11884
rect 7737 11828 7940 11884
rect 7996 11828 8082 11884
rect 8138 11828 8340 11884
rect 8396 11828 8482 11884
rect 8538 11828 8737 11884
rect 8793 11828 8879 11884
rect 8935 11828 9134 11884
rect 9190 11828 9276 11884
rect 9332 11828 9538 11884
rect 9594 11828 9680 11884
rect 9736 11828 9934 11884
rect 9990 11828 10076 11884
rect 10132 11828 10334 11884
rect 10390 11828 10476 11884
rect 10532 11828 10731 11884
rect 10787 11828 10873 11884
rect 10929 11828 11136 11884
rect 11192 11828 11278 11884
rect 11334 11828 11536 11884
rect 11592 11828 11678 11884
rect 11734 11828 11941 11884
rect 11997 11828 12083 11884
rect 12139 11862 13200 11884
rect 12139 11828 12526 11862
rect 266 11806 12526 11828
rect 12582 11806 12650 11862
rect 12706 11806 12774 11862
rect 12830 11806 12898 11862
rect 12954 11806 13022 11862
rect 13078 11806 13200 11862
rect -400 11742 13200 11806
rect -400 11738 741 11742
rect -400 11682 -286 11738
rect -230 11682 -162 11738
rect -106 11682 -38 11738
rect 18 11682 86 11738
rect 142 11682 210 11738
rect 266 11686 741 11738
rect 797 11686 883 11742
rect 939 11686 1142 11742
rect 1198 11686 1284 11742
rect 1340 11686 1542 11742
rect 1598 11686 1684 11742
rect 1740 11686 1939 11742
rect 1995 11686 2081 11742
rect 2137 11686 2336 11742
rect 2392 11686 2478 11742
rect 2534 11686 2740 11742
rect 2796 11686 2882 11742
rect 2938 11686 3136 11742
rect 3192 11686 3278 11742
rect 3334 11686 3536 11742
rect 3592 11686 3678 11742
rect 3734 11686 3933 11742
rect 3989 11686 4075 11742
rect 4131 11686 4338 11742
rect 4394 11686 4480 11742
rect 4536 11686 4738 11742
rect 4794 11686 4880 11742
rect 4936 11686 5143 11742
rect 5199 11686 5285 11742
rect 5341 11686 5540 11742
rect 5596 11686 5682 11742
rect 5738 11686 5937 11742
rect 5993 11686 6079 11742
rect 6135 11686 6340 11742
rect 6396 11686 6482 11742
rect 6538 11686 6742 11742
rect 6798 11686 6884 11742
rect 6940 11686 7145 11742
rect 7201 11686 7287 11742
rect 7343 11686 7539 11742
rect 7595 11686 7681 11742
rect 7737 11686 7940 11742
rect 7996 11686 8082 11742
rect 8138 11686 8340 11742
rect 8396 11686 8482 11742
rect 8538 11686 8737 11742
rect 8793 11686 8879 11742
rect 8935 11686 9134 11742
rect 9190 11686 9276 11742
rect 9332 11686 9538 11742
rect 9594 11686 9680 11742
rect 9736 11686 9934 11742
rect 9990 11686 10076 11742
rect 10132 11686 10334 11742
rect 10390 11686 10476 11742
rect 10532 11686 10731 11742
rect 10787 11686 10873 11742
rect 10929 11686 11136 11742
rect 11192 11686 11278 11742
rect 11334 11686 11536 11742
rect 11592 11686 11678 11742
rect 11734 11686 11941 11742
rect 11997 11686 12083 11742
rect 12139 11738 13200 11742
rect 12139 11686 12526 11738
rect 266 11682 12526 11686
rect 12582 11682 12650 11738
rect 12706 11682 12774 11738
rect 12830 11682 12898 11738
rect 12954 11682 13022 11738
rect 13078 11682 13200 11738
rect -400 11614 13200 11682
rect -400 11558 -286 11614
rect -230 11558 -162 11614
rect -106 11558 -38 11614
rect 18 11558 86 11614
rect 142 11558 210 11614
rect 266 11600 12526 11614
rect 266 11558 741 11600
rect -400 11544 741 11558
rect 797 11544 883 11600
rect 939 11544 1142 11600
rect 1198 11544 1284 11600
rect 1340 11544 1542 11600
rect 1598 11544 1684 11600
rect 1740 11544 1939 11600
rect 1995 11544 2081 11600
rect 2137 11544 2336 11600
rect 2392 11544 2478 11600
rect 2534 11544 2740 11600
rect 2796 11544 2882 11600
rect 2938 11544 3136 11600
rect 3192 11544 3278 11600
rect 3334 11544 3536 11600
rect 3592 11544 3678 11600
rect 3734 11544 3933 11600
rect 3989 11544 4075 11600
rect 4131 11544 4338 11600
rect 4394 11544 4480 11600
rect 4536 11544 4738 11600
rect 4794 11544 4880 11600
rect 4936 11544 5143 11600
rect 5199 11544 5285 11600
rect 5341 11544 5540 11600
rect 5596 11544 5682 11600
rect 5738 11544 5937 11600
rect 5993 11544 6079 11600
rect 6135 11544 6340 11600
rect 6396 11544 6482 11600
rect 6538 11544 6742 11600
rect 6798 11544 6884 11600
rect 6940 11544 7145 11600
rect 7201 11544 7287 11600
rect 7343 11544 7539 11600
rect 7595 11544 7681 11600
rect 7737 11544 7940 11600
rect 7996 11544 8082 11600
rect 8138 11544 8340 11600
rect 8396 11544 8482 11600
rect 8538 11544 8737 11600
rect 8793 11544 8879 11600
rect 8935 11544 9134 11600
rect 9190 11544 9276 11600
rect 9332 11544 9538 11600
rect 9594 11544 9680 11600
rect 9736 11544 9934 11600
rect 9990 11544 10076 11600
rect 10132 11544 10334 11600
rect 10390 11544 10476 11600
rect 10532 11544 10731 11600
rect 10787 11544 10873 11600
rect 10929 11544 11136 11600
rect 11192 11544 11278 11600
rect 11334 11544 11536 11600
rect 11592 11544 11678 11600
rect 11734 11544 11941 11600
rect 11997 11544 12083 11600
rect 12139 11558 12526 11600
rect 12582 11558 12650 11614
rect 12706 11558 12774 11614
rect 12830 11558 12898 11614
rect 12954 11558 13022 11614
rect 13078 11558 13200 11614
rect 12139 11544 13200 11558
rect -400 11490 13200 11544
rect -400 11434 -286 11490
rect -230 11434 -162 11490
rect -106 11434 -38 11490
rect 18 11434 86 11490
rect 142 11434 210 11490
rect 266 11458 12526 11490
rect 266 11434 741 11458
rect -400 11402 741 11434
rect 797 11402 883 11458
rect 939 11402 1142 11458
rect 1198 11402 1284 11458
rect 1340 11402 1542 11458
rect 1598 11402 1684 11458
rect 1740 11402 1939 11458
rect 1995 11402 2081 11458
rect 2137 11402 2336 11458
rect 2392 11402 2478 11458
rect 2534 11402 2740 11458
rect 2796 11402 2882 11458
rect 2938 11402 3136 11458
rect 3192 11402 3278 11458
rect 3334 11402 3536 11458
rect 3592 11402 3678 11458
rect 3734 11402 3933 11458
rect 3989 11402 4075 11458
rect 4131 11402 4338 11458
rect 4394 11402 4480 11458
rect 4536 11402 4738 11458
rect 4794 11402 4880 11458
rect 4936 11402 5143 11458
rect 5199 11402 5285 11458
rect 5341 11402 5540 11458
rect 5596 11402 5682 11458
rect 5738 11402 5937 11458
rect 5993 11402 6079 11458
rect 6135 11402 6340 11458
rect 6396 11402 6482 11458
rect 6538 11402 6742 11458
rect 6798 11402 6884 11458
rect 6940 11402 7145 11458
rect 7201 11402 7287 11458
rect 7343 11402 7539 11458
rect 7595 11402 7681 11458
rect 7737 11402 7940 11458
rect 7996 11402 8082 11458
rect 8138 11402 8340 11458
rect 8396 11402 8482 11458
rect 8538 11402 8737 11458
rect 8793 11402 8879 11458
rect 8935 11402 9134 11458
rect 9190 11402 9276 11458
rect 9332 11402 9538 11458
rect 9594 11402 9680 11458
rect 9736 11402 9934 11458
rect 9990 11402 10076 11458
rect 10132 11402 10334 11458
rect 10390 11402 10476 11458
rect 10532 11402 10731 11458
rect 10787 11402 10873 11458
rect 10929 11402 11136 11458
rect 11192 11402 11278 11458
rect 11334 11402 11536 11458
rect 11592 11402 11678 11458
rect 11734 11402 11941 11458
rect 11997 11402 12083 11458
rect 12139 11434 12526 11458
rect 12582 11434 12650 11490
rect 12706 11434 12774 11490
rect 12830 11434 12898 11490
rect 12954 11434 13022 11490
rect 13078 11434 13200 11490
rect 12139 11402 13200 11434
rect -400 11366 13200 11402
rect -400 11310 -286 11366
rect -230 11310 -162 11366
rect -106 11310 -38 11366
rect 18 11310 86 11366
rect 142 11310 210 11366
rect 266 11316 12526 11366
rect 266 11310 741 11316
rect -400 11260 741 11310
rect 797 11260 883 11316
rect 939 11260 1142 11316
rect 1198 11260 1284 11316
rect 1340 11260 1542 11316
rect 1598 11260 1684 11316
rect 1740 11260 1939 11316
rect 1995 11260 2081 11316
rect 2137 11260 2336 11316
rect 2392 11260 2478 11316
rect 2534 11260 2740 11316
rect 2796 11260 2882 11316
rect 2938 11260 3136 11316
rect 3192 11260 3278 11316
rect 3334 11260 3536 11316
rect 3592 11260 3678 11316
rect 3734 11260 3933 11316
rect 3989 11260 4075 11316
rect 4131 11260 4338 11316
rect 4394 11260 4480 11316
rect 4536 11260 4738 11316
rect 4794 11260 4880 11316
rect 4936 11260 5143 11316
rect 5199 11260 5285 11316
rect 5341 11260 5540 11316
rect 5596 11260 5682 11316
rect 5738 11260 5937 11316
rect 5993 11260 6079 11316
rect 6135 11260 6340 11316
rect 6396 11260 6482 11316
rect 6538 11260 6742 11316
rect 6798 11260 6884 11316
rect 6940 11260 7145 11316
rect 7201 11260 7287 11316
rect 7343 11260 7539 11316
rect 7595 11260 7681 11316
rect 7737 11260 7940 11316
rect 7996 11260 8082 11316
rect 8138 11260 8340 11316
rect 8396 11260 8482 11316
rect 8538 11260 8737 11316
rect 8793 11260 8879 11316
rect 8935 11260 9134 11316
rect 9190 11260 9276 11316
rect 9332 11260 9538 11316
rect 9594 11260 9680 11316
rect 9736 11260 9934 11316
rect 9990 11260 10076 11316
rect 10132 11260 10334 11316
rect 10390 11260 10476 11316
rect 10532 11260 10731 11316
rect 10787 11260 10873 11316
rect 10929 11260 11136 11316
rect 11192 11260 11278 11316
rect 11334 11260 11536 11316
rect 11592 11260 11678 11316
rect 11734 11260 11941 11316
rect 11997 11260 12083 11316
rect 12139 11310 12526 11316
rect 12582 11310 12650 11366
rect 12706 11310 12774 11366
rect 12830 11310 12898 11366
rect 12954 11310 13022 11366
rect 13078 11310 13200 11366
rect 12139 11260 13200 11310
rect -400 11242 13200 11260
rect -400 11186 -286 11242
rect -230 11186 -162 11242
rect -106 11186 -38 11242
rect 18 11186 86 11242
rect 142 11186 210 11242
rect 266 11186 12526 11242
rect 12582 11186 12650 11242
rect 12706 11186 12774 11242
rect 12830 11186 12898 11242
rect 12954 11186 13022 11242
rect 13078 11186 13200 11242
rect -400 11174 13200 11186
rect -400 11118 741 11174
rect 797 11118 883 11174
rect 939 11118 1142 11174
rect 1198 11118 1284 11174
rect 1340 11118 1542 11174
rect 1598 11118 1684 11174
rect 1740 11118 1939 11174
rect 1995 11118 2081 11174
rect 2137 11118 2336 11174
rect 2392 11118 2478 11174
rect 2534 11118 2740 11174
rect 2796 11118 2882 11174
rect 2938 11118 3136 11174
rect 3192 11118 3278 11174
rect 3334 11118 3536 11174
rect 3592 11118 3678 11174
rect 3734 11118 3933 11174
rect 3989 11118 4075 11174
rect 4131 11118 4338 11174
rect 4394 11118 4480 11174
rect 4536 11118 4738 11174
rect 4794 11118 4880 11174
rect 4936 11118 5143 11174
rect 5199 11118 5285 11174
rect 5341 11118 5540 11174
rect 5596 11118 5682 11174
rect 5738 11118 5937 11174
rect 5993 11118 6079 11174
rect 6135 11118 6340 11174
rect 6396 11118 6482 11174
rect 6538 11118 6742 11174
rect 6798 11118 6884 11174
rect 6940 11118 7145 11174
rect 7201 11118 7287 11174
rect 7343 11118 7539 11174
rect 7595 11118 7681 11174
rect 7737 11118 7940 11174
rect 7996 11118 8082 11174
rect 8138 11118 8340 11174
rect 8396 11118 8482 11174
rect 8538 11118 8737 11174
rect 8793 11118 8879 11174
rect 8935 11118 9134 11174
rect 9190 11118 9276 11174
rect 9332 11118 9538 11174
rect 9594 11118 9680 11174
rect 9736 11118 9934 11174
rect 9990 11118 10076 11174
rect 10132 11118 10334 11174
rect 10390 11118 10476 11174
rect 10532 11118 10731 11174
rect 10787 11118 10873 11174
rect 10929 11118 11136 11174
rect 11192 11118 11278 11174
rect 11334 11118 11536 11174
rect 11592 11118 11678 11174
rect 11734 11118 11941 11174
rect 11997 11118 12083 11174
rect 12139 11118 13200 11174
rect -400 11062 -286 11118
rect -230 11062 -162 11118
rect -106 11062 -38 11118
rect 18 11062 86 11118
rect 142 11062 210 11118
rect 266 11062 12526 11118
rect 12582 11062 12650 11118
rect 12706 11062 12774 11118
rect 12830 11062 12898 11118
rect 12954 11062 13022 11118
rect 13078 11062 13200 11118
rect -400 11032 13200 11062
rect -400 10994 741 11032
rect -400 10938 -286 10994
rect -230 10938 -162 10994
rect -106 10938 -38 10994
rect 18 10938 86 10994
rect 142 10938 210 10994
rect 266 10976 741 10994
rect 797 10976 883 11032
rect 939 10976 1142 11032
rect 1198 10976 1284 11032
rect 1340 10976 1542 11032
rect 1598 10976 1684 11032
rect 1740 10976 1939 11032
rect 1995 10976 2081 11032
rect 2137 10976 2336 11032
rect 2392 10976 2478 11032
rect 2534 10976 2740 11032
rect 2796 10976 2882 11032
rect 2938 10976 3136 11032
rect 3192 10976 3278 11032
rect 3334 10976 3536 11032
rect 3592 10976 3678 11032
rect 3734 10976 3933 11032
rect 3989 10976 4075 11032
rect 4131 10976 4338 11032
rect 4394 10976 4480 11032
rect 4536 10976 4738 11032
rect 4794 10976 4880 11032
rect 4936 10976 5143 11032
rect 5199 10976 5285 11032
rect 5341 10976 5540 11032
rect 5596 10976 5682 11032
rect 5738 10976 5937 11032
rect 5993 10976 6079 11032
rect 6135 10976 6340 11032
rect 6396 10976 6482 11032
rect 6538 10976 6742 11032
rect 6798 10976 6884 11032
rect 6940 10976 7145 11032
rect 7201 10976 7287 11032
rect 7343 10976 7539 11032
rect 7595 10976 7681 11032
rect 7737 10976 7940 11032
rect 7996 10976 8082 11032
rect 8138 10976 8340 11032
rect 8396 10976 8482 11032
rect 8538 10976 8737 11032
rect 8793 10976 8879 11032
rect 8935 10976 9134 11032
rect 9190 10976 9276 11032
rect 9332 10976 9538 11032
rect 9594 10976 9680 11032
rect 9736 10976 9934 11032
rect 9990 10976 10076 11032
rect 10132 10976 10334 11032
rect 10390 10976 10476 11032
rect 10532 10976 10731 11032
rect 10787 10976 10873 11032
rect 10929 10976 11136 11032
rect 11192 10976 11278 11032
rect 11334 10976 11536 11032
rect 11592 10976 11678 11032
rect 11734 10976 11941 11032
rect 11997 10976 12083 11032
rect 12139 10994 13200 11032
rect 12139 10976 12526 10994
rect 266 10938 12526 10976
rect 12582 10938 12650 10994
rect 12706 10938 12774 10994
rect 12830 10938 12898 10994
rect 12954 10938 13022 10994
rect 13078 10938 13200 10994
rect -400 10890 13200 10938
rect -400 10870 741 10890
rect -400 10814 -286 10870
rect -230 10814 -162 10870
rect -106 10814 -38 10870
rect 18 10814 86 10870
rect 142 10814 210 10870
rect 266 10834 741 10870
rect 797 10834 883 10890
rect 939 10834 1142 10890
rect 1198 10834 1284 10890
rect 1340 10834 1542 10890
rect 1598 10834 1684 10890
rect 1740 10834 1939 10890
rect 1995 10834 2081 10890
rect 2137 10834 2336 10890
rect 2392 10834 2478 10890
rect 2534 10834 2740 10890
rect 2796 10834 2882 10890
rect 2938 10834 3136 10890
rect 3192 10834 3278 10890
rect 3334 10834 3536 10890
rect 3592 10834 3678 10890
rect 3734 10834 3933 10890
rect 3989 10834 4075 10890
rect 4131 10834 4338 10890
rect 4394 10834 4480 10890
rect 4536 10834 4738 10890
rect 4794 10834 4880 10890
rect 4936 10834 5143 10890
rect 5199 10834 5285 10890
rect 5341 10834 5540 10890
rect 5596 10834 5682 10890
rect 5738 10834 5937 10890
rect 5993 10834 6079 10890
rect 6135 10834 6340 10890
rect 6396 10834 6482 10890
rect 6538 10834 6742 10890
rect 6798 10834 6884 10890
rect 6940 10834 7145 10890
rect 7201 10834 7287 10890
rect 7343 10834 7539 10890
rect 7595 10834 7681 10890
rect 7737 10834 7940 10890
rect 7996 10834 8082 10890
rect 8138 10834 8340 10890
rect 8396 10834 8482 10890
rect 8538 10834 8737 10890
rect 8793 10834 8879 10890
rect 8935 10834 9134 10890
rect 9190 10834 9276 10890
rect 9332 10834 9538 10890
rect 9594 10834 9680 10890
rect 9736 10834 9934 10890
rect 9990 10834 10076 10890
rect 10132 10834 10334 10890
rect 10390 10834 10476 10890
rect 10532 10834 10731 10890
rect 10787 10834 10873 10890
rect 10929 10834 11136 10890
rect 11192 10834 11278 10890
rect 11334 10834 11536 10890
rect 11592 10834 11678 10890
rect 11734 10834 11941 10890
rect 11997 10834 12083 10890
rect 12139 10870 13200 10890
rect 12139 10834 12526 10870
rect 266 10814 12526 10834
rect 12582 10814 12650 10870
rect 12706 10814 12774 10870
rect 12830 10814 12898 10870
rect 12954 10814 13022 10870
rect 13078 10814 13200 10870
rect -400 10748 13200 10814
rect -400 10746 741 10748
rect -400 10690 -286 10746
rect -230 10690 -162 10746
rect -106 10690 -38 10746
rect 18 10690 86 10746
rect 142 10690 210 10746
rect 266 10692 741 10746
rect 797 10692 883 10748
rect 939 10692 1142 10748
rect 1198 10692 1284 10748
rect 1340 10692 1542 10748
rect 1598 10692 1684 10748
rect 1740 10692 1939 10748
rect 1995 10692 2081 10748
rect 2137 10692 2336 10748
rect 2392 10692 2478 10748
rect 2534 10692 2740 10748
rect 2796 10692 2882 10748
rect 2938 10692 3136 10748
rect 3192 10692 3278 10748
rect 3334 10692 3536 10748
rect 3592 10692 3678 10748
rect 3734 10692 3933 10748
rect 3989 10692 4075 10748
rect 4131 10692 4338 10748
rect 4394 10692 4480 10748
rect 4536 10692 4738 10748
rect 4794 10692 4880 10748
rect 4936 10692 5143 10748
rect 5199 10692 5285 10748
rect 5341 10692 5540 10748
rect 5596 10692 5682 10748
rect 5738 10692 5937 10748
rect 5993 10692 6079 10748
rect 6135 10692 6340 10748
rect 6396 10692 6482 10748
rect 6538 10692 6742 10748
rect 6798 10692 6884 10748
rect 6940 10692 7145 10748
rect 7201 10692 7287 10748
rect 7343 10692 7539 10748
rect 7595 10692 7681 10748
rect 7737 10692 7940 10748
rect 7996 10692 8082 10748
rect 8138 10692 8340 10748
rect 8396 10692 8482 10748
rect 8538 10692 8737 10748
rect 8793 10692 8879 10748
rect 8935 10692 9134 10748
rect 9190 10692 9276 10748
rect 9332 10692 9538 10748
rect 9594 10692 9680 10748
rect 9736 10692 9934 10748
rect 9990 10692 10076 10748
rect 10132 10692 10334 10748
rect 10390 10692 10476 10748
rect 10532 10692 10731 10748
rect 10787 10692 10873 10748
rect 10929 10692 11136 10748
rect 11192 10692 11278 10748
rect 11334 10692 11536 10748
rect 11592 10692 11678 10748
rect 11734 10692 11941 10748
rect 11997 10692 12083 10748
rect 12139 10746 13200 10748
rect 12139 10692 12526 10746
rect 266 10690 12526 10692
rect 12582 10690 12650 10746
rect 12706 10690 12774 10746
rect 12830 10690 12898 10746
rect 12954 10690 13022 10746
rect 13078 10690 13200 10746
rect -400 10622 13200 10690
rect -400 10566 -286 10622
rect -230 10566 -162 10622
rect -106 10566 -38 10622
rect 18 10566 86 10622
rect 142 10566 210 10622
rect 266 10606 12526 10622
rect 266 10566 741 10606
rect -400 10550 741 10566
rect 797 10550 883 10606
rect 939 10550 1142 10606
rect 1198 10550 1284 10606
rect 1340 10550 1542 10606
rect 1598 10550 1684 10606
rect 1740 10550 1939 10606
rect 1995 10550 2081 10606
rect 2137 10550 2336 10606
rect 2392 10550 2478 10606
rect 2534 10550 2740 10606
rect 2796 10550 2882 10606
rect 2938 10550 3136 10606
rect 3192 10550 3278 10606
rect 3334 10550 3536 10606
rect 3592 10550 3678 10606
rect 3734 10550 3933 10606
rect 3989 10550 4075 10606
rect 4131 10550 4338 10606
rect 4394 10550 4480 10606
rect 4536 10550 4738 10606
rect 4794 10550 4880 10606
rect 4936 10550 5143 10606
rect 5199 10550 5285 10606
rect 5341 10550 5540 10606
rect 5596 10550 5682 10606
rect 5738 10550 5937 10606
rect 5993 10550 6079 10606
rect 6135 10550 6340 10606
rect 6396 10550 6482 10606
rect 6538 10550 6742 10606
rect 6798 10550 6884 10606
rect 6940 10550 7145 10606
rect 7201 10550 7287 10606
rect 7343 10550 7539 10606
rect 7595 10550 7681 10606
rect 7737 10550 7940 10606
rect 7996 10550 8082 10606
rect 8138 10550 8340 10606
rect 8396 10550 8482 10606
rect 8538 10550 8737 10606
rect 8793 10550 8879 10606
rect 8935 10550 9134 10606
rect 9190 10550 9276 10606
rect 9332 10550 9538 10606
rect 9594 10550 9680 10606
rect 9736 10550 9934 10606
rect 9990 10550 10076 10606
rect 10132 10550 10334 10606
rect 10390 10550 10476 10606
rect 10532 10550 10731 10606
rect 10787 10550 10873 10606
rect 10929 10550 11136 10606
rect 11192 10550 11278 10606
rect 11334 10550 11536 10606
rect 11592 10550 11678 10606
rect 11734 10550 11941 10606
rect 11997 10550 12083 10606
rect 12139 10566 12526 10606
rect 12582 10566 12650 10622
rect 12706 10566 12774 10622
rect 12830 10566 12898 10622
rect 12954 10566 13022 10622
rect 13078 10566 13200 10622
rect 12139 10550 13200 10566
rect -400 10498 13200 10550
rect -400 10442 -286 10498
rect -230 10442 -162 10498
rect -106 10442 -38 10498
rect 18 10442 86 10498
rect 142 10442 210 10498
rect 266 10464 12526 10498
rect 266 10442 741 10464
rect -400 10408 741 10442
rect 797 10408 883 10464
rect 939 10408 1142 10464
rect 1198 10408 1284 10464
rect 1340 10408 1542 10464
rect 1598 10408 1684 10464
rect 1740 10408 1939 10464
rect 1995 10408 2081 10464
rect 2137 10408 2336 10464
rect 2392 10408 2478 10464
rect 2534 10408 2740 10464
rect 2796 10408 2882 10464
rect 2938 10408 3136 10464
rect 3192 10408 3278 10464
rect 3334 10408 3536 10464
rect 3592 10408 3678 10464
rect 3734 10408 3933 10464
rect 3989 10408 4075 10464
rect 4131 10408 4338 10464
rect 4394 10408 4480 10464
rect 4536 10408 4738 10464
rect 4794 10408 4880 10464
rect 4936 10408 5143 10464
rect 5199 10408 5285 10464
rect 5341 10408 5540 10464
rect 5596 10408 5682 10464
rect 5738 10408 5937 10464
rect 5993 10408 6079 10464
rect 6135 10408 6340 10464
rect 6396 10408 6482 10464
rect 6538 10408 6742 10464
rect 6798 10408 6884 10464
rect 6940 10408 7145 10464
rect 7201 10408 7287 10464
rect 7343 10408 7539 10464
rect 7595 10408 7681 10464
rect 7737 10408 7940 10464
rect 7996 10408 8082 10464
rect 8138 10408 8340 10464
rect 8396 10408 8482 10464
rect 8538 10408 8737 10464
rect 8793 10408 8879 10464
rect 8935 10408 9134 10464
rect 9190 10408 9276 10464
rect 9332 10408 9538 10464
rect 9594 10408 9680 10464
rect 9736 10408 9934 10464
rect 9990 10408 10076 10464
rect 10132 10408 10334 10464
rect 10390 10408 10476 10464
rect 10532 10408 10731 10464
rect 10787 10408 10873 10464
rect 10929 10408 11136 10464
rect 11192 10408 11278 10464
rect 11334 10408 11536 10464
rect 11592 10408 11678 10464
rect 11734 10408 11941 10464
rect 11997 10408 12083 10464
rect 12139 10442 12526 10464
rect 12582 10442 12650 10498
rect 12706 10442 12774 10498
rect 12830 10442 12898 10498
rect 12954 10442 13022 10498
rect 13078 10442 13200 10498
rect 12139 10408 13200 10442
rect -400 10374 13200 10408
rect -400 10318 -286 10374
rect -230 10318 -162 10374
rect -106 10318 -38 10374
rect 18 10318 86 10374
rect 142 10318 210 10374
rect 266 10322 12526 10374
rect 266 10318 741 10322
rect -400 10266 741 10318
rect 797 10266 883 10322
rect 939 10266 1142 10322
rect 1198 10266 1284 10322
rect 1340 10266 1542 10322
rect 1598 10266 1684 10322
rect 1740 10266 1939 10322
rect 1995 10266 2081 10322
rect 2137 10266 2336 10322
rect 2392 10266 2478 10322
rect 2534 10266 2740 10322
rect 2796 10266 2882 10322
rect 2938 10266 3136 10322
rect 3192 10266 3278 10322
rect 3334 10266 3536 10322
rect 3592 10266 3678 10322
rect 3734 10266 3933 10322
rect 3989 10266 4075 10322
rect 4131 10266 4338 10322
rect 4394 10266 4480 10322
rect 4536 10266 4738 10322
rect 4794 10266 4880 10322
rect 4936 10266 5143 10322
rect 5199 10266 5285 10322
rect 5341 10266 5540 10322
rect 5596 10266 5682 10322
rect 5738 10266 5937 10322
rect 5993 10266 6079 10322
rect 6135 10266 6340 10322
rect 6396 10266 6482 10322
rect 6538 10266 6742 10322
rect 6798 10266 6884 10322
rect 6940 10266 7145 10322
rect 7201 10266 7287 10322
rect 7343 10266 7539 10322
rect 7595 10266 7681 10322
rect 7737 10266 7940 10322
rect 7996 10266 8082 10322
rect 8138 10266 8340 10322
rect 8396 10266 8482 10322
rect 8538 10266 8737 10322
rect 8793 10266 8879 10322
rect 8935 10266 9134 10322
rect 9190 10266 9276 10322
rect 9332 10266 9538 10322
rect 9594 10266 9680 10322
rect 9736 10266 9934 10322
rect 9990 10266 10076 10322
rect 10132 10266 10334 10322
rect 10390 10266 10476 10322
rect 10532 10266 10731 10322
rect 10787 10266 10873 10322
rect 10929 10266 11136 10322
rect 11192 10266 11278 10322
rect 11334 10266 11536 10322
rect 11592 10266 11678 10322
rect 11734 10266 11941 10322
rect 11997 10266 12083 10322
rect 12139 10318 12526 10322
rect 12582 10318 12650 10374
rect 12706 10318 12774 10374
rect 12830 10318 12898 10374
rect 12954 10318 13022 10374
rect 13078 10318 13200 10374
rect 12139 10266 13200 10318
rect -400 10250 13200 10266
rect -400 10194 -286 10250
rect -230 10194 -162 10250
rect -106 10194 -38 10250
rect 18 10194 86 10250
rect 142 10194 210 10250
rect 266 10194 12526 10250
rect 12582 10194 12650 10250
rect 12706 10194 12774 10250
rect 12830 10194 12898 10250
rect 12954 10194 13022 10250
rect 13078 10194 13200 10250
rect -400 10180 13200 10194
rect -400 10126 741 10180
rect -400 10070 -286 10126
rect -230 10070 -162 10126
rect -106 10070 -38 10126
rect 18 10070 86 10126
rect 142 10070 210 10126
rect 266 10124 741 10126
rect 797 10124 883 10180
rect 939 10124 1142 10180
rect 1198 10124 1284 10180
rect 1340 10124 1542 10180
rect 1598 10124 1684 10180
rect 1740 10124 1939 10180
rect 1995 10124 2081 10180
rect 2137 10124 2336 10180
rect 2392 10124 2478 10180
rect 2534 10124 2740 10180
rect 2796 10124 2882 10180
rect 2938 10124 3136 10180
rect 3192 10124 3278 10180
rect 3334 10124 3536 10180
rect 3592 10124 3678 10180
rect 3734 10124 3933 10180
rect 3989 10124 4075 10180
rect 4131 10124 4338 10180
rect 4394 10124 4480 10180
rect 4536 10124 4738 10180
rect 4794 10124 4880 10180
rect 4936 10124 5143 10180
rect 5199 10124 5285 10180
rect 5341 10124 5540 10180
rect 5596 10124 5682 10180
rect 5738 10124 5937 10180
rect 5993 10124 6079 10180
rect 6135 10124 6340 10180
rect 6396 10124 6482 10180
rect 6538 10124 6742 10180
rect 6798 10124 6884 10180
rect 6940 10124 7145 10180
rect 7201 10124 7287 10180
rect 7343 10124 7539 10180
rect 7595 10124 7681 10180
rect 7737 10124 7940 10180
rect 7996 10124 8082 10180
rect 8138 10124 8340 10180
rect 8396 10124 8482 10180
rect 8538 10124 8737 10180
rect 8793 10124 8879 10180
rect 8935 10124 9134 10180
rect 9190 10124 9276 10180
rect 9332 10124 9538 10180
rect 9594 10124 9680 10180
rect 9736 10124 9934 10180
rect 9990 10124 10076 10180
rect 10132 10124 10334 10180
rect 10390 10124 10476 10180
rect 10532 10124 10731 10180
rect 10787 10124 10873 10180
rect 10929 10124 11136 10180
rect 11192 10124 11278 10180
rect 11334 10124 11536 10180
rect 11592 10124 11678 10180
rect 11734 10124 11941 10180
rect 11997 10124 12083 10180
rect 12139 10126 13200 10180
rect 12139 10124 12526 10126
rect 266 10070 12526 10124
rect 12582 10070 12650 10126
rect 12706 10070 12774 10126
rect 12830 10070 12898 10126
rect 12954 10070 13022 10126
rect 13078 10070 13200 10126
rect -400 10038 13200 10070
rect -400 10002 741 10038
rect -400 9946 -286 10002
rect -230 9946 -162 10002
rect -106 9946 -38 10002
rect 18 9946 86 10002
rect 142 9946 210 10002
rect 266 9982 741 10002
rect 797 9982 883 10038
rect 939 9982 1142 10038
rect 1198 9982 1284 10038
rect 1340 9982 1542 10038
rect 1598 9982 1684 10038
rect 1740 9982 1939 10038
rect 1995 9982 2081 10038
rect 2137 9982 2336 10038
rect 2392 9982 2478 10038
rect 2534 9982 2740 10038
rect 2796 9982 2882 10038
rect 2938 9982 3136 10038
rect 3192 9982 3278 10038
rect 3334 9982 3536 10038
rect 3592 9982 3678 10038
rect 3734 9982 3933 10038
rect 3989 9982 4075 10038
rect 4131 9982 4338 10038
rect 4394 9982 4480 10038
rect 4536 9982 4738 10038
rect 4794 9982 4880 10038
rect 4936 9982 5143 10038
rect 5199 9982 5285 10038
rect 5341 9982 5540 10038
rect 5596 9982 5682 10038
rect 5738 9982 5937 10038
rect 5993 9982 6079 10038
rect 6135 9982 6340 10038
rect 6396 9982 6482 10038
rect 6538 9982 6742 10038
rect 6798 9982 6884 10038
rect 6940 9982 7145 10038
rect 7201 9982 7287 10038
rect 7343 9982 7539 10038
rect 7595 9982 7681 10038
rect 7737 9982 7940 10038
rect 7996 9982 8082 10038
rect 8138 9982 8340 10038
rect 8396 9982 8482 10038
rect 8538 9982 8737 10038
rect 8793 9982 8879 10038
rect 8935 9982 9134 10038
rect 9190 9982 9276 10038
rect 9332 9982 9538 10038
rect 9594 9982 9680 10038
rect 9736 9982 9934 10038
rect 9990 9982 10076 10038
rect 10132 9982 10334 10038
rect 10390 9982 10476 10038
rect 10532 9982 10731 10038
rect 10787 9982 10873 10038
rect 10929 9982 11136 10038
rect 11192 9982 11278 10038
rect 11334 9982 11536 10038
rect 11592 9982 11678 10038
rect 11734 9982 11941 10038
rect 11997 9982 12083 10038
rect 12139 10002 13200 10038
rect 12139 9982 12526 10002
rect 266 9946 12526 9982
rect 12582 9946 12650 10002
rect 12706 9946 12774 10002
rect 12830 9946 12898 10002
rect 12954 9946 13022 10002
rect 13078 9946 13200 10002
rect -400 9896 13200 9946
rect -400 9878 741 9896
rect -400 9822 -286 9878
rect -230 9822 -162 9878
rect -106 9822 -38 9878
rect 18 9822 86 9878
rect 142 9822 210 9878
rect 266 9840 741 9878
rect 797 9840 883 9896
rect 939 9840 1142 9896
rect 1198 9840 1284 9896
rect 1340 9840 1542 9896
rect 1598 9840 1684 9896
rect 1740 9840 1939 9896
rect 1995 9840 2081 9896
rect 2137 9840 2336 9896
rect 2392 9840 2478 9896
rect 2534 9840 2740 9896
rect 2796 9840 2882 9896
rect 2938 9840 3136 9896
rect 3192 9840 3278 9896
rect 3334 9840 3536 9896
rect 3592 9840 3678 9896
rect 3734 9840 3933 9896
rect 3989 9840 4075 9896
rect 4131 9840 4338 9896
rect 4394 9840 4480 9896
rect 4536 9840 4738 9896
rect 4794 9840 4880 9896
rect 4936 9840 5143 9896
rect 5199 9840 5285 9896
rect 5341 9840 5540 9896
rect 5596 9840 5682 9896
rect 5738 9840 5937 9896
rect 5993 9840 6079 9896
rect 6135 9840 6340 9896
rect 6396 9840 6482 9896
rect 6538 9840 6742 9896
rect 6798 9840 6884 9896
rect 6940 9840 7145 9896
rect 7201 9840 7287 9896
rect 7343 9840 7539 9896
rect 7595 9840 7681 9896
rect 7737 9840 7940 9896
rect 7996 9840 8082 9896
rect 8138 9840 8340 9896
rect 8396 9840 8482 9896
rect 8538 9840 8737 9896
rect 8793 9840 8879 9896
rect 8935 9840 9134 9896
rect 9190 9840 9276 9896
rect 9332 9840 9538 9896
rect 9594 9840 9680 9896
rect 9736 9840 9934 9896
rect 9990 9840 10076 9896
rect 10132 9840 10334 9896
rect 10390 9840 10476 9896
rect 10532 9840 10731 9896
rect 10787 9840 10873 9896
rect 10929 9840 11136 9896
rect 11192 9840 11278 9896
rect 11334 9840 11536 9896
rect 11592 9840 11678 9896
rect 11734 9840 11941 9896
rect 11997 9840 12083 9896
rect 12139 9878 13200 9896
rect 12139 9840 12526 9878
rect 266 9822 12526 9840
rect 12582 9822 12650 9878
rect 12706 9822 12774 9878
rect 12830 9822 12898 9878
rect 12954 9822 13022 9878
rect 13078 9822 13200 9878
rect -400 9754 13200 9822
rect -400 9698 -286 9754
rect -230 9698 -162 9754
rect -106 9698 -38 9754
rect 18 9698 86 9754
rect 142 9698 210 9754
rect 266 9698 741 9754
rect 797 9698 883 9754
rect 939 9698 1142 9754
rect 1198 9698 1284 9754
rect 1340 9698 1542 9754
rect 1598 9698 1684 9754
rect 1740 9698 1939 9754
rect 1995 9698 2081 9754
rect 2137 9698 2336 9754
rect 2392 9698 2478 9754
rect 2534 9698 2740 9754
rect 2796 9698 2882 9754
rect 2938 9698 3136 9754
rect 3192 9698 3278 9754
rect 3334 9698 3536 9754
rect 3592 9698 3678 9754
rect 3734 9698 3933 9754
rect 3989 9698 4075 9754
rect 4131 9698 4338 9754
rect 4394 9698 4480 9754
rect 4536 9698 4738 9754
rect 4794 9698 4880 9754
rect 4936 9698 5143 9754
rect 5199 9698 5285 9754
rect 5341 9698 5540 9754
rect 5596 9698 5682 9754
rect 5738 9698 5937 9754
rect 5993 9698 6079 9754
rect 6135 9698 6340 9754
rect 6396 9698 6482 9754
rect 6538 9698 6742 9754
rect 6798 9698 6884 9754
rect 6940 9698 7145 9754
rect 7201 9698 7287 9754
rect 7343 9698 7539 9754
rect 7595 9698 7681 9754
rect 7737 9698 7940 9754
rect 7996 9698 8082 9754
rect 8138 9698 8340 9754
rect 8396 9698 8482 9754
rect 8538 9698 8737 9754
rect 8793 9698 8879 9754
rect 8935 9698 9134 9754
rect 9190 9698 9276 9754
rect 9332 9698 9538 9754
rect 9594 9698 9680 9754
rect 9736 9698 9934 9754
rect 9990 9698 10076 9754
rect 10132 9698 10334 9754
rect 10390 9698 10476 9754
rect 10532 9698 10731 9754
rect 10787 9698 10873 9754
rect 10929 9698 11136 9754
rect 11192 9698 11278 9754
rect 11334 9698 11536 9754
rect 11592 9698 11678 9754
rect 11734 9698 11941 9754
rect 11997 9698 12083 9754
rect 12139 9698 12526 9754
rect 12582 9698 12650 9754
rect 12706 9698 12774 9754
rect 12830 9698 12898 9754
rect 12954 9698 13022 9754
rect 13078 9698 13200 9754
rect -400 9630 13200 9698
rect -400 9574 -286 9630
rect -230 9574 -162 9630
rect -106 9574 -38 9630
rect 18 9574 86 9630
rect 142 9574 210 9630
rect 266 9612 12526 9630
rect 266 9574 741 9612
rect -400 9556 741 9574
rect 797 9556 883 9612
rect 939 9556 1142 9612
rect 1198 9556 1284 9612
rect 1340 9556 1542 9612
rect 1598 9556 1684 9612
rect 1740 9556 1939 9612
rect 1995 9556 2081 9612
rect 2137 9556 2336 9612
rect 2392 9556 2478 9612
rect 2534 9556 2740 9612
rect 2796 9556 2882 9612
rect 2938 9556 3136 9612
rect 3192 9556 3278 9612
rect 3334 9556 3536 9612
rect 3592 9556 3678 9612
rect 3734 9556 3933 9612
rect 3989 9556 4075 9612
rect 4131 9556 4338 9612
rect 4394 9556 4480 9612
rect 4536 9556 4738 9612
rect 4794 9556 4880 9612
rect 4936 9556 5143 9612
rect 5199 9556 5285 9612
rect 5341 9556 5540 9612
rect 5596 9556 5682 9612
rect 5738 9556 5937 9612
rect 5993 9556 6079 9612
rect 6135 9556 6340 9612
rect 6396 9556 6482 9612
rect 6538 9556 6742 9612
rect 6798 9556 6884 9612
rect 6940 9556 7145 9612
rect 7201 9556 7287 9612
rect 7343 9556 7539 9612
rect 7595 9556 7681 9612
rect 7737 9556 7940 9612
rect 7996 9556 8082 9612
rect 8138 9556 8340 9612
rect 8396 9556 8482 9612
rect 8538 9556 8737 9612
rect 8793 9556 8879 9612
rect 8935 9556 9134 9612
rect 9190 9556 9276 9612
rect 9332 9556 9538 9612
rect 9594 9556 9680 9612
rect 9736 9556 9934 9612
rect 9990 9556 10076 9612
rect 10132 9556 10334 9612
rect 10390 9556 10476 9612
rect 10532 9556 10731 9612
rect 10787 9556 10873 9612
rect 10929 9556 11136 9612
rect 11192 9556 11278 9612
rect 11334 9556 11536 9612
rect 11592 9556 11678 9612
rect 11734 9556 11941 9612
rect 11997 9556 12083 9612
rect 12139 9574 12526 9612
rect 12582 9574 12650 9630
rect 12706 9574 12774 9630
rect 12830 9574 12898 9630
rect 12954 9574 13022 9630
rect 13078 9574 13200 9630
rect 12139 9556 13200 9574
rect -400 9506 13200 9556
rect -400 9450 -286 9506
rect -230 9450 -162 9506
rect -106 9450 -38 9506
rect 18 9450 86 9506
rect 142 9450 210 9506
rect 266 9470 12526 9506
rect 266 9450 741 9470
rect -400 9414 741 9450
rect 797 9414 883 9470
rect 939 9414 1142 9470
rect 1198 9414 1284 9470
rect 1340 9414 1542 9470
rect 1598 9414 1684 9470
rect 1740 9414 1939 9470
rect 1995 9414 2081 9470
rect 2137 9414 2336 9470
rect 2392 9414 2478 9470
rect 2534 9414 2740 9470
rect 2796 9414 2882 9470
rect 2938 9414 3136 9470
rect 3192 9414 3278 9470
rect 3334 9414 3536 9470
rect 3592 9414 3678 9470
rect 3734 9414 3933 9470
rect 3989 9414 4075 9470
rect 4131 9414 4338 9470
rect 4394 9414 4480 9470
rect 4536 9414 4738 9470
rect 4794 9414 4880 9470
rect 4936 9414 5143 9470
rect 5199 9414 5285 9470
rect 5341 9414 5540 9470
rect 5596 9414 5682 9470
rect 5738 9414 5937 9470
rect 5993 9414 6079 9470
rect 6135 9414 6340 9470
rect 6396 9414 6482 9470
rect 6538 9414 6742 9470
rect 6798 9414 6884 9470
rect 6940 9414 7145 9470
rect 7201 9414 7287 9470
rect 7343 9414 7539 9470
rect 7595 9414 7681 9470
rect 7737 9414 7940 9470
rect 7996 9414 8082 9470
rect 8138 9414 8340 9470
rect 8396 9414 8482 9470
rect 8538 9414 8737 9470
rect 8793 9414 8879 9470
rect 8935 9414 9134 9470
rect 9190 9414 9276 9470
rect 9332 9414 9538 9470
rect 9594 9414 9680 9470
rect 9736 9414 9934 9470
rect 9990 9414 10076 9470
rect 10132 9414 10334 9470
rect 10390 9414 10476 9470
rect 10532 9414 10731 9470
rect 10787 9414 10873 9470
rect 10929 9414 11136 9470
rect 11192 9414 11278 9470
rect 11334 9414 11536 9470
rect 11592 9414 11678 9470
rect 11734 9414 11941 9470
rect 11997 9414 12083 9470
rect 12139 9450 12526 9470
rect 12582 9450 12650 9506
rect 12706 9450 12774 9506
rect 12830 9450 12898 9506
rect 12954 9450 13022 9506
rect 13078 9450 13200 9506
rect 12139 9414 13200 9450
rect -400 9382 13200 9414
rect -400 9326 -286 9382
rect -230 9326 -162 9382
rect -106 9326 -38 9382
rect 18 9326 86 9382
rect 142 9326 210 9382
rect 266 9328 12526 9382
rect 266 9326 741 9328
rect -400 9272 741 9326
rect 797 9272 883 9328
rect 939 9272 1142 9328
rect 1198 9272 1284 9328
rect 1340 9272 1542 9328
rect 1598 9272 1684 9328
rect 1740 9272 1939 9328
rect 1995 9272 2081 9328
rect 2137 9272 2336 9328
rect 2392 9272 2478 9328
rect 2534 9272 2740 9328
rect 2796 9272 2882 9328
rect 2938 9272 3136 9328
rect 3192 9272 3278 9328
rect 3334 9272 3536 9328
rect 3592 9272 3678 9328
rect 3734 9272 3933 9328
rect 3989 9272 4075 9328
rect 4131 9272 4338 9328
rect 4394 9272 4480 9328
rect 4536 9272 4738 9328
rect 4794 9272 4880 9328
rect 4936 9272 5143 9328
rect 5199 9272 5285 9328
rect 5341 9272 5540 9328
rect 5596 9272 5682 9328
rect 5738 9272 5937 9328
rect 5993 9272 6079 9328
rect 6135 9272 6340 9328
rect 6396 9272 6482 9328
rect 6538 9272 6742 9328
rect 6798 9272 6884 9328
rect 6940 9272 7145 9328
rect 7201 9272 7287 9328
rect 7343 9272 7539 9328
rect 7595 9272 7681 9328
rect 7737 9272 7940 9328
rect 7996 9272 8082 9328
rect 8138 9272 8340 9328
rect 8396 9272 8482 9328
rect 8538 9272 8737 9328
rect 8793 9272 8879 9328
rect 8935 9272 9134 9328
rect 9190 9272 9276 9328
rect 9332 9272 9538 9328
rect 9594 9272 9680 9328
rect 9736 9272 9934 9328
rect 9990 9272 10076 9328
rect 10132 9272 10334 9328
rect 10390 9272 10476 9328
rect 10532 9272 10731 9328
rect 10787 9272 10873 9328
rect 10929 9272 11136 9328
rect 11192 9272 11278 9328
rect 11334 9272 11536 9328
rect 11592 9272 11678 9328
rect 11734 9272 11941 9328
rect 11997 9272 12083 9328
rect 12139 9326 12526 9328
rect 12582 9326 12650 9382
rect 12706 9326 12774 9382
rect 12830 9326 12898 9382
rect 12954 9326 13022 9382
rect 13078 9326 13200 9382
rect 12139 9272 13200 9326
rect -400 9258 13200 9272
rect -400 9202 -286 9258
rect -230 9202 -162 9258
rect -106 9202 -38 9258
rect 18 9202 86 9258
rect 142 9202 210 9258
rect 266 9202 12526 9258
rect 12582 9202 12650 9258
rect 12706 9202 12774 9258
rect 12830 9202 12898 9258
rect 12954 9202 13022 9258
rect 13078 9202 13200 9258
rect -400 9186 13200 9202
rect -400 9134 741 9186
rect -400 9078 -286 9134
rect -230 9078 -162 9134
rect -106 9078 -38 9134
rect 18 9078 86 9134
rect 142 9078 210 9134
rect 266 9130 741 9134
rect 797 9130 883 9186
rect 939 9130 1142 9186
rect 1198 9130 1284 9186
rect 1340 9130 1542 9186
rect 1598 9130 1684 9186
rect 1740 9130 1939 9186
rect 1995 9130 2081 9186
rect 2137 9130 2336 9186
rect 2392 9130 2478 9186
rect 2534 9130 2740 9186
rect 2796 9130 2882 9186
rect 2938 9130 3136 9186
rect 3192 9130 3278 9186
rect 3334 9130 3536 9186
rect 3592 9130 3678 9186
rect 3734 9130 3933 9186
rect 3989 9130 4075 9186
rect 4131 9130 4338 9186
rect 4394 9130 4480 9186
rect 4536 9130 4738 9186
rect 4794 9130 4880 9186
rect 4936 9130 5143 9186
rect 5199 9130 5285 9186
rect 5341 9130 5540 9186
rect 5596 9130 5682 9186
rect 5738 9130 5937 9186
rect 5993 9130 6079 9186
rect 6135 9130 6340 9186
rect 6396 9130 6482 9186
rect 6538 9130 6742 9186
rect 6798 9130 6884 9186
rect 6940 9130 7145 9186
rect 7201 9130 7287 9186
rect 7343 9130 7539 9186
rect 7595 9130 7681 9186
rect 7737 9130 7940 9186
rect 7996 9130 8082 9186
rect 8138 9130 8340 9186
rect 8396 9130 8482 9186
rect 8538 9130 8737 9186
rect 8793 9130 8879 9186
rect 8935 9130 9134 9186
rect 9190 9130 9276 9186
rect 9332 9130 9538 9186
rect 9594 9130 9680 9186
rect 9736 9130 9934 9186
rect 9990 9130 10076 9186
rect 10132 9130 10334 9186
rect 10390 9130 10476 9186
rect 10532 9130 10731 9186
rect 10787 9130 10873 9186
rect 10929 9130 11136 9186
rect 11192 9130 11278 9186
rect 11334 9130 11536 9186
rect 11592 9130 11678 9186
rect 11734 9130 11941 9186
rect 11997 9130 12083 9186
rect 12139 9134 13200 9186
rect 12139 9130 12526 9134
rect 266 9078 12526 9130
rect 12582 9078 12650 9134
rect 12706 9078 12774 9134
rect 12830 9078 12898 9134
rect 12954 9078 13022 9134
rect 13078 9078 13200 9134
rect -400 9044 13200 9078
rect -400 9010 741 9044
rect -400 8954 -286 9010
rect -230 8954 -162 9010
rect -106 8954 -38 9010
rect 18 8954 86 9010
rect 142 8954 210 9010
rect 266 8988 741 9010
rect 797 8988 883 9044
rect 939 8988 1142 9044
rect 1198 8988 1284 9044
rect 1340 8988 1542 9044
rect 1598 8988 1684 9044
rect 1740 8988 1939 9044
rect 1995 8988 2081 9044
rect 2137 8988 2336 9044
rect 2392 8988 2478 9044
rect 2534 8988 2740 9044
rect 2796 8988 2882 9044
rect 2938 8988 3136 9044
rect 3192 8988 3278 9044
rect 3334 8988 3536 9044
rect 3592 8988 3678 9044
rect 3734 8988 3933 9044
rect 3989 8988 4075 9044
rect 4131 8988 4338 9044
rect 4394 8988 4480 9044
rect 4536 8988 4738 9044
rect 4794 8988 4880 9044
rect 4936 8988 5143 9044
rect 5199 8988 5285 9044
rect 5341 8988 5540 9044
rect 5596 8988 5682 9044
rect 5738 8988 5937 9044
rect 5993 8988 6079 9044
rect 6135 8988 6340 9044
rect 6396 8988 6482 9044
rect 6538 8988 6742 9044
rect 6798 8988 6884 9044
rect 6940 8988 7145 9044
rect 7201 8988 7287 9044
rect 7343 8988 7539 9044
rect 7595 8988 7681 9044
rect 7737 8988 7940 9044
rect 7996 8988 8082 9044
rect 8138 8988 8340 9044
rect 8396 8988 8482 9044
rect 8538 8988 8737 9044
rect 8793 8988 8879 9044
rect 8935 8988 9134 9044
rect 9190 8988 9276 9044
rect 9332 8988 9538 9044
rect 9594 8988 9680 9044
rect 9736 8988 9934 9044
rect 9990 8988 10076 9044
rect 10132 8988 10334 9044
rect 10390 8988 10476 9044
rect 10532 8988 10731 9044
rect 10787 8988 10873 9044
rect 10929 8988 11136 9044
rect 11192 8988 11278 9044
rect 11334 8988 11536 9044
rect 11592 8988 11678 9044
rect 11734 8988 11941 9044
rect 11997 8988 12083 9044
rect 12139 9010 13200 9044
rect 12139 8988 12526 9010
rect 266 8954 12526 8988
rect 12582 8954 12650 9010
rect 12706 8954 12774 9010
rect 12830 8954 12898 9010
rect 12954 8954 13022 9010
rect 13078 8954 13200 9010
rect -400 8902 13200 8954
rect -400 8886 741 8902
rect -400 8830 -286 8886
rect -230 8830 -162 8886
rect -106 8830 -38 8886
rect 18 8830 86 8886
rect 142 8830 210 8886
rect 266 8846 741 8886
rect 797 8846 883 8902
rect 939 8846 1142 8902
rect 1198 8846 1284 8902
rect 1340 8846 1542 8902
rect 1598 8846 1684 8902
rect 1740 8846 1939 8902
rect 1995 8846 2081 8902
rect 2137 8846 2336 8902
rect 2392 8846 2478 8902
rect 2534 8846 2740 8902
rect 2796 8846 2882 8902
rect 2938 8846 3136 8902
rect 3192 8846 3278 8902
rect 3334 8846 3536 8902
rect 3592 8846 3678 8902
rect 3734 8846 3933 8902
rect 3989 8846 4075 8902
rect 4131 8846 4338 8902
rect 4394 8846 4480 8902
rect 4536 8846 4738 8902
rect 4794 8846 4880 8902
rect 4936 8846 5143 8902
rect 5199 8846 5285 8902
rect 5341 8846 5540 8902
rect 5596 8846 5682 8902
rect 5738 8846 5937 8902
rect 5993 8846 6079 8902
rect 6135 8846 6340 8902
rect 6396 8846 6482 8902
rect 6538 8846 6742 8902
rect 6798 8846 6884 8902
rect 6940 8846 7145 8902
rect 7201 8846 7287 8902
rect 7343 8846 7539 8902
rect 7595 8846 7681 8902
rect 7737 8846 7940 8902
rect 7996 8846 8082 8902
rect 8138 8846 8340 8902
rect 8396 8846 8482 8902
rect 8538 8846 8737 8902
rect 8793 8846 8879 8902
rect 8935 8846 9134 8902
rect 9190 8846 9276 8902
rect 9332 8846 9538 8902
rect 9594 8846 9680 8902
rect 9736 8846 9934 8902
rect 9990 8846 10076 8902
rect 10132 8846 10334 8902
rect 10390 8846 10476 8902
rect 10532 8846 10731 8902
rect 10787 8846 10873 8902
rect 10929 8846 11136 8902
rect 11192 8846 11278 8902
rect 11334 8846 11536 8902
rect 11592 8846 11678 8902
rect 11734 8846 11941 8902
rect 11997 8846 12083 8902
rect 12139 8886 13200 8902
rect 12139 8846 12526 8886
rect 266 8830 12526 8846
rect 12582 8830 12650 8886
rect 12706 8830 12774 8886
rect 12830 8830 12898 8886
rect 12954 8830 13022 8886
rect 13078 8830 13200 8886
rect -400 8762 13200 8830
rect -400 8706 -286 8762
rect -230 8706 -162 8762
rect -106 8706 -38 8762
rect 18 8706 86 8762
rect 142 8706 210 8762
rect 266 8760 12526 8762
rect 266 8706 741 8760
rect -400 8704 741 8706
rect 797 8704 883 8760
rect 939 8704 1142 8760
rect 1198 8704 1284 8760
rect 1340 8704 1542 8760
rect 1598 8704 1684 8760
rect 1740 8704 1939 8760
rect 1995 8704 2081 8760
rect 2137 8704 2336 8760
rect 2392 8704 2478 8760
rect 2534 8704 2740 8760
rect 2796 8704 2882 8760
rect 2938 8704 3136 8760
rect 3192 8704 3278 8760
rect 3334 8704 3536 8760
rect 3592 8704 3678 8760
rect 3734 8704 3933 8760
rect 3989 8704 4075 8760
rect 4131 8704 4338 8760
rect 4394 8704 4480 8760
rect 4536 8704 4738 8760
rect 4794 8704 4880 8760
rect 4936 8704 5143 8760
rect 5199 8704 5285 8760
rect 5341 8704 5540 8760
rect 5596 8704 5682 8760
rect 5738 8704 5937 8760
rect 5993 8704 6079 8760
rect 6135 8704 6340 8760
rect 6396 8704 6482 8760
rect 6538 8704 6742 8760
rect 6798 8704 6884 8760
rect 6940 8704 7145 8760
rect 7201 8704 7287 8760
rect 7343 8704 7539 8760
rect 7595 8704 7681 8760
rect 7737 8704 7940 8760
rect 7996 8704 8082 8760
rect 8138 8704 8340 8760
rect 8396 8704 8482 8760
rect 8538 8704 8737 8760
rect 8793 8704 8879 8760
rect 8935 8704 9134 8760
rect 9190 8704 9276 8760
rect 9332 8704 9538 8760
rect 9594 8704 9680 8760
rect 9736 8704 9934 8760
rect 9990 8704 10076 8760
rect 10132 8704 10334 8760
rect 10390 8704 10476 8760
rect 10532 8704 10731 8760
rect 10787 8704 10873 8760
rect 10929 8704 11136 8760
rect 11192 8704 11278 8760
rect 11334 8704 11536 8760
rect 11592 8704 11678 8760
rect 11734 8704 11941 8760
rect 11997 8704 12083 8760
rect 12139 8706 12526 8760
rect 12582 8706 12650 8762
rect 12706 8706 12774 8762
rect 12830 8706 12898 8762
rect 12954 8706 13022 8762
rect 13078 8706 13200 8762
rect 12139 8704 13200 8706
rect -400 8638 13200 8704
rect -400 8582 -286 8638
rect -230 8582 -162 8638
rect -106 8582 -38 8638
rect 18 8582 86 8638
rect 142 8582 210 8638
rect 266 8618 12526 8638
rect 266 8582 741 8618
rect -400 8562 741 8582
rect 797 8562 883 8618
rect 939 8562 1142 8618
rect 1198 8562 1284 8618
rect 1340 8562 1542 8618
rect 1598 8562 1684 8618
rect 1740 8562 1939 8618
rect 1995 8562 2081 8618
rect 2137 8562 2336 8618
rect 2392 8562 2478 8618
rect 2534 8562 2740 8618
rect 2796 8562 2882 8618
rect 2938 8562 3136 8618
rect 3192 8562 3278 8618
rect 3334 8562 3536 8618
rect 3592 8562 3678 8618
rect 3734 8562 3933 8618
rect 3989 8562 4075 8618
rect 4131 8562 4338 8618
rect 4394 8562 4480 8618
rect 4536 8562 4738 8618
rect 4794 8562 4880 8618
rect 4936 8562 5143 8618
rect 5199 8562 5285 8618
rect 5341 8562 5540 8618
rect 5596 8562 5682 8618
rect 5738 8562 5937 8618
rect 5993 8562 6079 8618
rect 6135 8562 6340 8618
rect 6396 8562 6482 8618
rect 6538 8562 6742 8618
rect 6798 8562 6884 8618
rect 6940 8562 7145 8618
rect 7201 8562 7287 8618
rect 7343 8562 7539 8618
rect 7595 8562 7681 8618
rect 7737 8562 7940 8618
rect 7996 8562 8082 8618
rect 8138 8562 8340 8618
rect 8396 8562 8482 8618
rect 8538 8562 8737 8618
rect 8793 8562 8879 8618
rect 8935 8562 9134 8618
rect 9190 8562 9276 8618
rect 9332 8562 9538 8618
rect 9594 8562 9680 8618
rect 9736 8562 9934 8618
rect 9990 8562 10076 8618
rect 10132 8562 10334 8618
rect 10390 8562 10476 8618
rect 10532 8562 10731 8618
rect 10787 8562 10873 8618
rect 10929 8562 11136 8618
rect 11192 8562 11278 8618
rect 11334 8562 11536 8618
rect 11592 8562 11678 8618
rect 11734 8562 11941 8618
rect 11997 8562 12083 8618
rect 12139 8582 12526 8618
rect 12582 8582 12650 8638
rect 12706 8582 12774 8638
rect 12830 8582 12898 8638
rect 12954 8582 13022 8638
rect 13078 8582 13200 8638
rect 12139 8562 13200 8582
rect -400 8514 13200 8562
rect -400 8458 -286 8514
rect -230 8458 -162 8514
rect -106 8458 -38 8514
rect 18 8458 86 8514
rect 142 8458 210 8514
rect 266 8476 12526 8514
rect 266 8458 741 8476
rect -400 8420 741 8458
rect 797 8420 883 8476
rect 939 8420 1142 8476
rect 1198 8420 1284 8476
rect 1340 8420 1542 8476
rect 1598 8420 1684 8476
rect 1740 8420 1939 8476
rect 1995 8420 2081 8476
rect 2137 8420 2336 8476
rect 2392 8420 2478 8476
rect 2534 8420 2740 8476
rect 2796 8420 2882 8476
rect 2938 8420 3136 8476
rect 3192 8420 3278 8476
rect 3334 8420 3536 8476
rect 3592 8420 3678 8476
rect 3734 8420 3933 8476
rect 3989 8420 4075 8476
rect 4131 8420 4338 8476
rect 4394 8420 4480 8476
rect 4536 8420 4738 8476
rect 4794 8420 4880 8476
rect 4936 8420 5143 8476
rect 5199 8420 5285 8476
rect 5341 8420 5540 8476
rect 5596 8420 5682 8476
rect 5738 8420 5937 8476
rect 5993 8420 6079 8476
rect 6135 8420 6340 8476
rect 6396 8420 6482 8476
rect 6538 8420 6742 8476
rect 6798 8420 6884 8476
rect 6940 8420 7145 8476
rect 7201 8420 7287 8476
rect 7343 8420 7539 8476
rect 7595 8420 7681 8476
rect 7737 8420 7940 8476
rect 7996 8420 8082 8476
rect 8138 8420 8340 8476
rect 8396 8420 8482 8476
rect 8538 8420 8737 8476
rect 8793 8420 8879 8476
rect 8935 8420 9134 8476
rect 9190 8420 9276 8476
rect 9332 8420 9538 8476
rect 9594 8420 9680 8476
rect 9736 8420 9934 8476
rect 9990 8420 10076 8476
rect 10132 8420 10334 8476
rect 10390 8420 10476 8476
rect 10532 8420 10731 8476
rect 10787 8420 10873 8476
rect 10929 8420 11136 8476
rect 11192 8420 11278 8476
rect 11334 8420 11536 8476
rect 11592 8420 11678 8476
rect 11734 8420 11941 8476
rect 11997 8420 12083 8476
rect 12139 8458 12526 8476
rect 12582 8458 12650 8514
rect 12706 8458 12774 8514
rect 12830 8458 12898 8514
rect 12954 8458 13022 8514
rect 13078 8458 13200 8514
rect 12139 8420 13200 8458
rect -400 8390 13200 8420
rect -400 8334 -286 8390
rect -230 8334 -162 8390
rect -106 8334 -38 8390
rect 18 8334 86 8390
rect 142 8334 210 8390
rect 266 8334 12526 8390
rect 12582 8334 12650 8390
rect 12706 8334 12774 8390
rect 12830 8334 12898 8390
rect 12954 8334 13022 8390
rect 13078 8334 13200 8390
rect -400 8278 741 8334
rect 797 8278 883 8334
rect 939 8278 1142 8334
rect 1198 8278 1284 8334
rect 1340 8278 1542 8334
rect 1598 8278 1684 8334
rect 1740 8278 1939 8334
rect 1995 8278 2081 8334
rect 2137 8278 2336 8334
rect 2392 8278 2478 8334
rect 2534 8278 2740 8334
rect 2796 8278 2882 8334
rect 2938 8278 3136 8334
rect 3192 8278 3278 8334
rect 3334 8278 3536 8334
rect 3592 8278 3678 8334
rect 3734 8278 3933 8334
rect 3989 8278 4075 8334
rect 4131 8278 4338 8334
rect 4394 8278 4480 8334
rect 4536 8278 4738 8334
rect 4794 8278 4880 8334
rect 4936 8278 5143 8334
rect 5199 8278 5285 8334
rect 5341 8278 5540 8334
rect 5596 8278 5682 8334
rect 5738 8278 5937 8334
rect 5993 8278 6079 8334
rect 6135 8278 6340 8334
rect 6396 8278 6482 8334
rect 6538 8278 6742 8334
rect 6798 8278 6884 8334
rect 6940 8278 7145 8334
rect 7201 8278 7287 8334
rect 7343 8278 7539 8334
rect 7595 8278 7681 8334
rect 7737 8278 7940 8334
rect 7996 8278 8082 8334
rect 8138 8278 8340 8334
rect 8396 8278 8482 8334
rect 8538 8278 8737 8334
rect 8793 8278 8879 8334
rect 8935 8278 9134 8334
rect 9190 8278 9276 8334
rect 9332 8278 9538 8334
rect 9594 8278 9680 8334
rect 9736 8278 9934 8334
rect 9990 8278 10076 8334
rect 10132 8278 10334 8334
rect 10390 8278 10476 8334
rect 10532 8278 10731 8334
rect 10787 8278 10873 8334
rect 10929 8278 11136 8334
rect 11192 8278 11278 8334
rect 11334 8278 11536 8334
rect 11592 8278 11678 8334
rect 11734 8278 11941 8334
rect 11997 8278 12083 8334
rect 12139 8278 13200 8334
rect -400 8266 13200 8278
rect -400 8210 -286 8266
rect -230 8210 -162 8266
rect -106 8210 -38 8266
rect 18 8210 86 8266
rect 142 8210 210 8266
rect 266 8210 12526 8266
rect 12582 8210 12650 8266
rect 12706 8210 12774 8266
rect 12830 8210 12898 8266
rect 12954 8210 13022 8266
rect 13078 8210 13200 8266
rect -400 8192 13200 8210
rect -400 8142 741 8192
rect -400 8086 -286 8142
rect -230 8086 -162 8142
rect -106 8086 -38 8142
rect 18 8086 86 8142
rect 142 8086 210 8142
rect 266 8136 741 8142
rect 797 8136 883 8192
rect 939 8136 1142 8192
rect 1198 8136 1284 8192
rect 1340 8136 1542 8192
rect 1598 8136 1684 8192
rect 1740 8136 1939 8192
rect 1995 8136 2081 8192
rect 2137 8136 2336 8192
rect 2392 8136 2478 8192
rect 2534 8136 2740 8192
rect 2796 8136 2882 8192
rect 2938 8136 3136 8192
rect 3192 8136 3278 8192
rect 3334 8136 3536 8192
rect 3592 8136 3678 8192
rect 3734 8136 3933 8192
rect 3989 8136 4075 8192
rect 4131 8136 4338 8192
rect 4394 8136 4480 8192
rect 4536 8136 4738 8192
rect 4794 8136 4880 8192
rect 4936 8136 5143 8192
rect 5199 8136 5285 8192
rect 5341 8136 5540 8192
rect 5596 8136 5682 8192
rect 5738 8136 5937 8192
rect 5993 8136 6079 8192
rect 6135 8136 6340 8192
rect 6396 8136 6482 8192
rect 6538 8136 6742 8192
rect 6798 8136 6884 8192
rect 6940 8136 7145 8192
rect 7201 8136 7287 8192
rect 7343 8136 7539 8192
rect 7595 8136 7681 8192
rect 7737 8136 7940 8192
rect 7996 8136 8082 8192
rect 8138 8136 8340 8192
rect 8396 8136 8482 8192
rect 8538 8136 8737 8192
rect 8793 8136 8879 8192
rect 8935 8136 9134 8192
rect 9190 8136 9276 8192
rect 9332 8136 9538 8192
rect 9594 8136 9680 8192
rect 9736 8136 9934 8192
rect 9990 8136 10076 8192
rect 10132 8136 10334 8192
rect 10390 8136 10476 8192
rect 10532 8136 10731 8192
rect 10787 8136 10873 8192
rect 10929 8136 11136 8192
rect 11192 8136 11278 8192
rect 11334 8136 11536 8192
rect 11592 8136 11678 8192
rect 11734 8136 11941 8192
rect 11997 8136 12083 8192
rect 12139 8142 13200 8192
rect 12139 8136 12526 8142
rect 266 8086 12526 8136
rect 12582 8086 12650 8142
rect 12706 8086 12774 8142
rect 12830 8086 12898 8142
rect 12954 8086 13022 8142
rect 13078 8086 13200 8142
rect -400 8050 13200 8086
rect -400 8018 741 8050
rect -400 7962 -286 8018
rect -230 7962 -162 8018
rect -106 7962 -38 8018
rect 18 7962 86 8018
rect 142 7962 210 8018
rect 266 7994 741 8018
rect 797 7994 883 8050
rect 939 7994 1142 8050
rect 1198 7994 1284 8050
rect 1340 7994 1542 8050
rect 1598 7994 1684 8050
rect 1740 7994 1939 8050
rect 1995 7994 2081 8050
rect 2137 7994 2336 8050
rect 2392 7994 2478 8050
rect 2534 7994 2740 8050
rect 2796 7994 2882 8050
rect 2938 7994 3136 8050
rect 3192 7994 3278 8050
rect 3334 7994 3536 8050
rect 3592 7994 3678 8050
rect 3734 7994 3933 8050
rect 3989 7994 4075 8050
rect 4131 7994 4338 8050
rect 4394 7994 4480 8050
rect 4536 7994 4738 8050
rect 4794 7994 4880 8050
rect 4936 7994 5143 8050
rect 5199 7994 5285 8050
rect 5341 7994 5540 8050
rect 5596 7994 5682 8050
rect 5738 7994 5937 8050
rect 5993 7994 6079 8050
rect 6135 7994 6340 8050
rect 6396 7994 6482 8050
rect 6538 7994 6742 8050
rect 6798 7994 6884 8050
rect 6940 7994 7145 8050
rect 7201 7994 7287 8050
rect 7343 7994 7539 8050
rect 7595 7994 7681 8050
rect 7737 7994 7940 8050
rect 7996 7994 8082 8050
rect 8138 7994 8340 8050
rect 8396 7994 8482 8050
rect 8538 7994 8737 8050
rect 8793 7994 8879 8050
rect 8935 7994 9134 8050
rect 9190 7994 9276 8050
rect 9332 7994 9538 8050
rect 9594 7994 9680 8050
rect 9736 7994 9934 8050
rect 9990 7994 10076 8050
rect 10132 7994 10334 8050
rect 10390 7994 10476 8050
rect 10532 7994 10731 8050
rect 10787 7994 10873 8050
rect 10929 7994 11136 8050
rect 11192 7994 11278 8050
rect 11334 7994 11536 8050
rect 11592 7994 11678 8050
rect 11734 7994 11941 8050
rect 11997 7994 12083 8050
rect 12139 8018 13200 8050
rect 12139 7994 12526 8018
rect 266 7962 12526 7994
rect 12582 7962 12650 8018
rect 12706 7962 12774 8018
rect 12830 7962 12898 8018
rect 12954 7962 13022 8018
rect 13078 7962 13200 8018
rect -400 7908 13200 7962
rect -400 7894 741 7908
rect -400 7838 -286 7894
rect -230 7838 -162 7894
rect -106 7838 -38 7894
rect 18 7838 86 7894
rect 142 7838 210 7894
rect 266 7852 741 7894
rect 797 7852 883 7908
rect 939 7852 1142 7908
rect 1198 7852 1284 7908
rect 1340 7852 1542 7908
rect 1598 7852 1684 7908
rect 1740 7852 1939 7908
rect 1995 7852 2081 7908
rect 2137 7852 2336 7908
rect 2392 7852 2478 7908
rect 2534 7852 2740 7908
rect 2796 7852 2882 7908
rect 2938 7852 3136 7908
rect 3192 7852 3278 7908
rect 3334 7852 3536 7908
rect 3592 7852 3678 7908
rect 3734 7852 3933 7908
rect 3989 7852 4075 7908
rect 4131 7852 4338 7908
rect 4394 7852 4480 7908
rect 4536 7852 4738 7908
rect 4794 7852 4880 7908
rect 4936 7852 5143 7908
rect 5199 7852 5285 7908
rect 5341 7852 5540 7908
rect 5596 7852 5682 7908
rect 5738 7852 5937 7908
rect 5993 7852 6079 7908
rect 6135 7852 6340 7908
rect 6396 7852 6482 7908
rect 6538 7852 6742 7908
rect 6798 7852 6884 7908
rect 6940 7852 7145 7908
rect 7201 7852 7287 7908
rect 7343 7852 7539 7908
rect 7595 7852 7681 7908
rect 7737 7852 7940 7908
rect 7996 7852 8082 7908
rect 8138 7852 8340 7908
rect 8396 7852 8482 7908
rect 8538 7852 8737 7908
rect 8793 7852 8879 7908
rect 8935 7852 9134 7908
rect 9190 7852 9276 7908
rect 9332 7852 9538 7908
rect 9594 7852 9680 7908
rect 9736 7852 9934 7908
rect 9990 7852 10076 7908
rect 10132 7852 10334 7908
rect 10390 7852 10476 7908
rect 10532 7852 10731 7908
rect 10787 7852 10873 7908
rect 10929 7852 11136 7908
rect 11192 7852 11278 7908
rect 11334 7852 11536 7908
rect 11592 7852 11678 7908
rect 11734 7852 11941 7908
rect 11997 7852 12083 7908
rect 12139 7894 13200 7908
rect 12139 7852 12526 7894
rect 266 7838 12526 7852
rect 12582 7838 12650 7894
rect 12706 7838 12774 7894
rect 12830 7838 12898 7894
rect 12954 7838 13022 7894
rect 13078 7838 13200 7894
rect -400 7770 13200 7838
rect -400 7714 -286 7770
rect -230 7714 -162 7770
rect -106 7714 -38 7770
rect 18 7714 86 7770
rect 142 7714 210 7770
rect 266 7766 12526 7770
rect 266 7714 741 7766
rect -400 7710 741 7714
rect 797 7710 883 7766
rect 939 7710 1142 7766
rect 1198 7710 1284 7766
rect 1340 7710 1542 7766
rect 1598 7710 1684 7766
rect 1740 7710 1939 7766
rect 1995 7710 2081 7766
rect 2137 7710 2336 7766
rect 2392 7710 2478 7766
rect 2534 7710 2740 7766
rect 2796 7710 2882 7766
rect 2938 7710 3136 7766
rect 3192 7710 3278 7766
rect 3334 7710 3536 7766
rect 3592 7710 3678 7766
rect 3734 7710 3933 7766
rect 3989 7710 4075 7766
rect 4131 7710 4338 7766
rect 4394 7710 4480 7766
rect 4536 7710 4738 7766
rect 4794 7710 4880 7766
rect 4936 7710 5143 7766
rect 5199 7710 5285 7766
rect 5341 7710 5540 7766
rect 5596 7710 5682 7766
rect 5738 7710 5937 7766
rect 5993 7710 6079 7766
rect 6135 7710 6340 7766
rect 6396 7710 6482 7766
rect 6538 7710 6742 7766
rect 6798 7710 6884 7766
rect 6940 7710 7145 7766
rect 7201 7710 7287 7766
rect 7343 7710 7539 7766
rect 7595 7710 7681 7766
rect 7737 7710 7940 7766
rect 7996 7710 8082 7766
rect 8138 7710 8340 7766
rect 8396 7710 8482 7766
rect 8538 7710 8737 7766
rect 8793 7710 8879 7766
rect 8935 7710 9134 7766
rect 9190 7710 9276 7766
rect 9332 7710 9538 7766
rect 9594 7710 9680 7766
rect 9736 7710 9934 7766
rect 9990 7710 10076 7766
rect 10132 7710 10334 7766
rect 10390 7710 10476 7766
rect 10532 7710 10731 7766
rect 10787 7710 10873 7766
rect 10929 7710 11136 7766
rect 11192 7710 11278 7766
rect 11334 7710 11536 7766
rect 11592 7710 11678 7766
rect 11734 7710 11941 7766
rect 11997 7710 12083 7766
rect 12139 7714 12526 7766
rect 12582 7714 12650 7770
rect 12706 7714 12774 7770
rect 12830 7714 12898 7770
rect 12954 7714 13022 7770
rect 13078 7714 13200 7770
rect 12139 7710 13200 7714
rect -400 7646 13200 7710
rect -400 7590 -286 7646
rect -230 7590 -162 7646
rect -106 7590 -38 7646
rect 18 7590 86 7646
rect 142 7590 210 7646
rect 266 7624 12526 7646
rect 266 7590 741 7624
rect -400 7568 741 7590
rect 797 7568 883 7624
rect 939 7568 1142 7624
rect 1198 7568 1284 7624
rect 1340 7568 1542 7624
rect 1598 7568 1684 7624
rect 1740 7568 1939 7624
rect 1995 7568 2081 7624
rect 2137 7568 2336 7624
rect 2392 7568 2478 7624
rect 2534 7568 2740 7624
rect 2796 7568 2882 7624
rect 2938 7568 3136 7624
rect 3192 7568 3278 7624
rect 3334 7568 3536 7624
rect 3592 7568 3678 7624
rect 3734 7568 3933 7624
rect 3989 7568 4075 7624
rect 4131 7568 4338 7624
rect 4394 7568 4480 7624
rect 4536 7568 4738 7624
rect 4794 7568 4880 7624
rect 4936 7568 5143 7624
rect 5199 7568 5285 7624
rect 5341 7568 5540 7624
rect 5596 7568 5682 7624
rect 5738 7568 5937 7624
rect 5993 7568 6079 7624
rect 6135 7568 6340 7624
rect 6396 7568 6482 7624
rect 6538 7568 6742 7624
rect 6798 7568 6884 7624
rect 6940 7568 7145 7624
rect 7201 7568 7287 7624
rect 7343 7568 7539 7624
rect 7595 7568 7681 7624
rect 7737 7568 7940 7624
rect 7996 7568 8082 7624
rect 8138 7568 8340 7624
rect 8396 7568 8482 7624
rect 8538 7568 8737 7624
rect 8793 7568 8879 7624
rect 8935 7568 9134 7624
rect 9190 7568 9276 7624
rect 9332 7568 9538 7624
rect 9594 7568 9680 7624
rect 9736 7568 9934 7624
rect 9990 7568 10076 7624
rect 10132 7568 10334 7624
rect 10390 7568 10476 7624
rect 10532 7568 10731 7624
rect 10787 7568 10873 7624
rect 10929 7568 11136 7624
rect 11192 7568 11278 7624
rect 11334 7568 11536 7624
rect 11592 7568 11678 7624
rect 11734 7568 11941 7624
rect 11997 7568 12083 7624
rect 12139 7590 12526 7624
rect 12582 7590 12650 7646
rect 12706 7590 12774 7646
rect 12830 7590 12898 7646
rect 12954 7590 13022 7646
rect 13078 7590 13200 7646
rect 12139 7568 13200 7590
rect -400 7522 13200 7568
rect -400 7466 -286 7522
rect -230 7466 -162 7522
rect -106 7466 -38 7522
rect 18 7466 86 7522
rect 142 7466 210 7522
rect 266 7482 12526 7522
rect 266 7466 741 7482
rect -400 7426 741 7466
rect 797 7426 883 7482
rect 939 7426 1142 7482
rect 1198 7426 1284 7482
rect 1340 7426 1542 7482
rect 1598 7426 1684 7482
rect 1740 7426 1939 7482
rect 1995 7426 2081 7482
rect 2137 7426 2336 7482
rect 2392 7426 2478 7482
rect 2534 7426 2740 7482
rect 2796 7426 2882 7482
rect 2938 7426 3136 7482
rect 3192 7426 3278 7482
rect 3334 7426 3536 7482
rect 3592 7426 3678 7482
rect 3734 7426 3933 7482
rect 3989 7426 4075 7482
rect 4131 7426 4338 7482
rect 4394 7426 4480 7482
rect 4536 7426 4738 7482
rect 4794 7426 4880 7482
rect 4936 7426 5143 7482
rect 5199 7426 5285 7482
rect 5341 7426 5540 7482
rect 5596 7426 5682 7482
rect 5738 7426 5937 7482
rect 5993 7426 6079 7482
rect 6135 7426 6340 7482
rect 6396 7426 6482 7482
rect 6538 7426 6742 7482
rect 6798 7426 6884 7482
rect 6940 7426 7145 7482
rect 7201 7426 7287 7482
rect 7343 7426 7539 7482
rect 7595 7426 7681 7482
rect 7737 7426 7940 7482
rect 7996 7426 8082 7482
rect 8138 7426 8340 7482
rect 8396 7426 8482 7482
rect 8538 7426 8737 7482
rect 8793 7426 8879 7482
rect 8935 7426 9134 7482
rect 9190 7426 9276 7482
rect 9332 7426 9538 7482
rect 9594 7426 9680 7482
rect 9736 7426 9934 7482
rect 9990 7426 10076 7482
rect 10132 7426 10334 7482
rect 10390 7426 10476 7482
rect 10532 7426 10731 7482
rect 10787 7426 10873 7482
rect 10929 7426 11136 7482
rect 11192 7426 11278 7482
rect 11334 7426 11536 7482
rect 11592 7426 11678 7482
rect 11734 7426 11941 7482
rect 11997 7426 12083 7482
rect 12139 7466 12526 7482
rect 12582 7466 12650 7522
rect 12706 7466 12774 7522
rect 12830 7466 12898 7522
rect 12954 7466 13022 7522
rect 13078 7466 13200 7522
rect 12139 7426 13200 7466
rect -400 7398 13200 7426
rect -400 7342 -286 7398
rect -230 7342 -162 7398
rect -106 7342 -38 7398
rect 18 7342 86 7398
rect 142 7342 210 7398
rect 266 7342 12526 7398
rect 12582 7342 12650 7398
rect 12706 7342 12774 7398
rect 12830 7342 12898 7398
rect 12954 7342 13022 7398
rect 13078 7342 13200 7398
rect -400 7340 13200 7342
rect -400 7284 741 7340
rect 797 7284 883 7340
rect 939 7284 1142 7340
rect 1198 7284 1284 7340
rect 1340 7284 1542 7340
rect 1598 7284 1684 7340
rect 1740 7284 1939 7340
rect 1995 7284 2081 7340
rect 2137 7284 2336 7340
rect 2392 7284 2478 7340
rect 2534 7284 2740 7340
rect 2796 7284 2882 7340
rect 2938 7284 3136 7340
rect 3192 7284 3278 7340
rect 3334 7284 3536 7340
rect 3592 7284 3678 7340
rect 3734 7284 3933 7340
rect 3989 7284 4075 7340
rect 4131 7284 4338 7340
rect 4394 7284 4480 7340
rect 4536 7284 4738 7340
rect 4794 7284 4880 7340
rect 4936 7284 5143 7340
rect 5199 7284 5285 7340
rect 5341 7284 5540 7340
rect 5596 7284 5682 7340
rect 5738 7284 5937 7340
rect 5993 7284 6079 7340
rect 6135 7284 6340 7340
rect 6396 7284 6482 7340
rect 6538 7284 6742 7340
rect 6798 7284 6884 7340
rect 6940 7284 7145 7340
rect 7201 7284 7287 7340
rect 7343 7284 7539 7340
rect 7595 7284 7681 7340
rect 7737 7284 7940 7340
rect 7996 7284 8082 7340
rect 8138 7284 8340 7340
rect 8396 7284 8482 7340
rect 8538 7284 8737 7340
rect 8793 7284 8879 7340
rect 8935 7284 9134 7340
rect 9190 7284 9276 7340
rect 9332 7284 9538 7340
rect 9594 7284 9680 7340
rect 9736 7284 9934 7340
rect 9990 7284 10076 7340
rect 10132 7284 10334 7340
rect 10390 7284 10476 7340
rect 10532 7284 10731 7340
rect 10787 7284 10873 7340
rect 10929 7284 11136 7340
rect 11192 7284 11278 7340
rect 11334 7284 11536 7340
rect 11592 7284 11678 7340
rect 11734 7284 11941 7340
rect 11997 7284 12083 7340
rect 12139 7284 13200 7340
rect -400 7274 13200 7284
rect -400 7218 -286 7274
rect -230 7218 -162 7274
rect -106 7218 -38 7274
rect 18 7218 86 7274
rect 142 7218 210 7274
rect 266 7218 12526 7274
rect 12582 7218 12650 7274
rect 12706 7218 12774 7274
rect 12830 7218 12898 7274
rect 12954 7218 13022 7274
rect 13078 7218 13200 7274
rect -400 7198 13200 7218
rect -400 7150 741 7198
rect -400 7094 -286 7150
rect -230 7094 -162 7150
rect -106 7094 -38 7150
rect 18 7094 86 7150
rect 142 7094 210 7150
rect 266 7142 741 7150
rect 797 7142 883 7198
rect 939 7142 1142 7198
rect 1198 7142 1284 7198
rect 1340 7142 1542 7198
rect 1598 7142 1684 7198
rect 1740 7142 1939 7198
rect 1995 7142 2081 7198
rect 2137 7142 2336 7198
rect 2392 7142 2478 7198
rect 2534 7142 2740 7198
rect 2796 7142 2882 7198
rect 2938 7142 3136 7198
rect 3192 7142 3278 7198
rect 3334 7142 3536 7198
rect 3592 7142 3678 7198
rect 3734 7142 3933 7198
rect 3989 7142 4075 7198
rect 4131 7142 4338 7198
rect 4394 7142 4480 7198
rect 4536 7142 4738 7198
rect 4794 7142 4880 7198
rect 4936 7142 5143 7198
rect 5199 7142 5285 7198
rect 5341 7142 5540 7198
rect 5596 7142 5682 7198
rect 5738 7142 5937 7198
rect 5993 7142 6079 7198
rect 6135 7142 6340 7198
rect 6396 7142 6482 7198
rect 6538 7142 6742 7198
rect 6798 7142 6884 7198
rect 6940 7142 7145 7198
rect 7201 7142 7287 7198
rect 7343 7142 7539 7198
rect 7595 7142 7681 7198
rect 7737 7142 7940 7198
rect 7996 7142 8082 7198
rect 8138 7142 8340 7198
rect 8396 7142 8482 7198
rect 8538 7142 8737 7198
rect 8793 7142 8879 7198
rect 8935 7142 9134 7198
rect 9190 7142 9276 7198
rect 9332 7142 9538 7198
rect 9594 7142 9680 7198
rect 9736 7142 9934 7198
rect 9990 7142 10076 7198
rect 10132 7142 10334 7198
rect 10390 7142 10476 7198
rect 10532 7142 10731 7198
rect 10787 7142 10873 7198
rect 10929 7142 11136 7198
rect 11192 7142 11278 7198
rect 11334 7142 11536 7198
rect 11592 7142 11678 7198
rect 11734 7142 11941 7198
rect 11997 7142 12083 7198
rect 12139 7150 13200 7198
rect 12139 7142 12526 7150
rect 266 7094 12526 7142
rect 12582 7094 12650 7150
rect 12706 7094 12774 7150
rect 12830 7094 12898 7150
rect 12954 7094 13022 7150
rect 13078 7094 13200 7150
rect -400 7056 13200 7094
rect -400 7026 741 7056
rect -400 6970 -286 7026
rect -230 6970 -162 7026
rect -106 6970 -38 7026
rect 18 6970 86 7026
rect 142 6970 210 7026
rect 266 7000 741 7026
rect 797 7000 883 7056
rect 939 7000 1142 7056
rect 1198 7000 1284 7056
rect 1340 7000 1542 7056
rect 1598 7000 1684 7056
rect 1740 7000 1939 7056
rect 1995 7000 2081 7056
rect 2137 7000 2336 7056
rect 2392 7000 2478 7056
rect 2534 7000 2740 7056
rect 2796 7000 2882 7056
rect 2938 7000 3136 7056
rect 3192 7000 3278 7056
rect 3334 7000 3536 7056
rect 3592 7000 3678 7056
rect 3734 7000 3933 7056
rect 3989 7000 4075 7056
rect 4131 7000 4338 7056
rect 4394 7000 4480 7056
rect 4536 7000 4738 7056
rect 4794 7000 4880 7056
rect 4936 7000 5143 7056
rect 5199 7000 5285 7056
rect 5341 7000 5540 7056
rect 5596 7000 5682 7056
rect 5738 7000 5937 7056
rect 5993 7000 6079 7056
rect 6135 7000 6340 7056
rect 6396 7000 6482 7056
rect 6538 7000 6742 7056
rect 6798 7000 6884 7056
rect 6940 7000 7145 7056
rect 7201 7000 7287 7056
rect 7343 7000 7539 7056
rect 7595 7000 7681 7056
rect 7737 7000 7940 7056
rect 7996 7000 8082 7056
rect 8138 7000 8340 7056
rect 8396 7000 8482 7056
rect 8538 7000 8737 7056
rect 8793 7000 8879 7056
rect 8935 7000 9134 7056
rect 9190 7000 9276 7056
rect 9332 7000 9538 7056
rect 9594 7000 9680 7056
rect 9736 7000 9934 7056
rect 9990 7000 10076 7056
rect 10132 7000 10334 7056
rect 10390 7000 10476 7056
rect 10532 7000 10731 7056
rect 10787 7000 10873 7056
rect 10929 7000 11136 7056
rect 11192 7000 11278 7056
rect 11334 7000 11536 7056
rect 11592 7000 11678 7056
rect 11734 7000 11941 7056
rect 11997 7000 12083 7056
rect 12139 7026 13200 7056
rect 12139 7000 12526 7026
rect 266 6970 12526 7000
rect 12582 6970 12650 7026
rect 12706 6970 12774 7026
rect 12830 6970 12898 7026
rect 12954 6970 13022 7026
rect 13078 6970 13200 7026
rect -400 6914 13200 6970
rect -400 6902 741 6914
rect -400 6846 -286 6902
rect -230 6846 -162 6902
rect -106 6846 -38 6902
rect 18 6846 86 6902
rect 142 6846 210 6902
rect 266 6858 741 6902
rect 797 6858 883 6914
rect 939 6858 1142 6914
rect 1198 6858 1284 6914
rect 1340 6858 1542 6914
rect 1598 6858 1684 6914
rect 1740 6858 1939 6914
rect 1995 6858 2081 6914
rect 2137 6858 2336 6914
rect 2392 6858 2478 6914
rect 2534 6858 2740 6914
rect 2796 6858 2882 6914
rect 2938 6858 3136 6914
rect 3192 6858 3278 6914
rect 3334 6858 3536 6914
rect 3592 6858 3678 6914
rect 3734 6858 3933 6914
rect 3989 6858 4075 6914
rect 4131 6858 4338 6914
rect 4394 6858 4480 6914
rect 4536 6858 4738 6914
rect 4794 6858 4880 6914
rect 4936 6858 5143 6914
rect 5199 6858 5285 6914
rect 5341 6858 5540 6914
rect 5596 6858 5682 6914
rect 5738 6858 5937 6914
rect 5993 6858 6079 6914
rect 6135 6858 6340 6914
rect 6396 6858 6482 6914
rect 6538 6858 6742 6914
rect 6798 6858 6884 6914
rect 6940 6858 7145 6914
rect 7201 6858 7287 6914
rect 7343 6858 7539 6914
rect 7595 6858 7681 6914
rect 7737 6858 7940 6914
rect 7996 6858 8082 6914
rect 8138 6858 8340 6914
rect 8396 6858 8482 6914
rect 8538 6858 8737 6914
rect 8793 6858 8879 6914
rect 8935 6858 9134 6914
rect 9190 6858 9276 6914
rect 9332 6858 9538 6914
rect 9594 6858 9680 6914
rect 9736 6858 9934 6914
rect 9990 6858 10076 6914
rect 10132 6858 10334 6914
rect 10390 6858 10476 6914
rect 10532 6858 10731 6914
rect 10787 6858 10873 6914
rect 10929 6858 11136 6914
rect 11192 6858 11278 6914
rect 11334 6858 11536 6914
rect 11592 6858 11678 6914
rect 11734 6858 11941 6914
rect 11997 6858 12083 6914
rect 12139 6902 13200 6914
rect 12139 6858 12526 6902
rect 266 6846 12526 6858
rect 12582 6846 12650 6902
rect 12706 6846 12774 6902
rect 12830 6846 12898 6902
rect 12954 6846 13022 6902
rect 13078 6846 13200 6902
rect -400 6778 13200 6846
rect -400 6722 -286 6778
rect -230 6722 -162 6778
rect -106 6722 -38 6778
rect 18 6722 86 6778
rect 142 6722 210 6778
rect 266 6772 12526 6778
rect 266 6722 741 6772
rect -400 6716 741 6722
rect 797 6716 883 6772
rect 939 6716 1142 6772
rect 1198 6716 1284 6772
rect 1340 6716 1542 6772
rect 1598 6716 1684 6772
rect 1740 6716 1939 6772
rect 1995 6716 2081 6772
rect 2137 6716 2336 6772
rect 2392 6716 2478 6772
rect 2534 6716 2740 6772
rect 2796 6716 2882 6772
rect 2938 6716 3136 6772
rect 3192 6716 3278 6772
rect 3334 6716 3536 6772
rect 3592 6716 3678 6772
rect 3734 6716 3933 6772
rect 3989 6716 4075 6772
rect 4131 6716 4338 6772
rect 4394 6716 4480 6772
rect 4536 6716 4738 6772
rect 4794 6716 4880 6772
rect 4936 6716 5143 6772
rect 5199 6716 5285 6772
rect 5341 6716 5540 6772
rect 5596 6716 5682 6772
rect 5738 6716 5937 6772
rect 5993 6716 6079 6772
rect 6135 6716 6340 6772
rect 6396 6716 6482 6772
rect 6538 6716 6742 6772
rect 6798 6716 6884 6772
rect 6940 6716 7145 6772
rect 7201 6716 7287 6772
rect 7343 6716 7539 6772
rect 7595 6716 7681 6772
rect 7737 6716 7940 6772
rect 7996 6716 8082 6772
rect 8138 6716 8340 6772
rect 8396 6716 8482 6772
rect 8538 6716 8737 6772
rect 8793 6716 8879 6772
rect 8935 6716 9134 6772
rect 9190 6716 9276 6772
rect 9332 6716 9538 6772
rect 9594 6716 9680 6772
rect 9736 6716 9934 6772
rect 9990 6716 10076 6772
rect 10132 6716 10334 6772
rect 10390 6716 10476 6772
rect 10532 6716 10731 6772
rect 10787 6716 10873 6772
rect 10929 6716 11136 6772
rect 11192 6716 11278 6772
rect 11334 6716 11536 6772
rect 11592 6716 11678 6772
rect 11734 6716 11941 6772
rect 11997 6716 12083 6772
rect 12139 6722 12526 6772
rect 12582 6722 12650 6778
rect 12706 6722 12774 6778
rect 12830 6722 12898 6778
rect 12954 6722 13022 6778
rect 13078 6722 13200 6778
rect 12139 6716 13200 6722
rect -400 6654 13200 6716
rect -400 6598 -286 6654
rect -230 6598 -162 6654
rect -106 6598 -38 6654
rect 18 6598 86 6654
rect 142 6598 210 6654
rect 266 6630 12526 6654
rect 266 6598 741 6630
rect -400 6574 741 6598
rect 797 6574 883 6630
rect 939 6574 1142 6630
rect 1198 6574 1284 6630
rect 1340 6574 1542 6630
rect 1598 6574 1684 6630
rect 1740 6574 1939 6630
rect 1995 6574 2081 6630
rect 2137 6574 2336 6630
rect 2392 6574 2478 6630
rect 2534 6574 2740 6630
rect 2796 6574 2882 6630
rect 2938 6574 3136 6630
rect 3192 6574 3278 6630
rect 3334 6574 3536 6630
rect 3592 6574 3678 6630
rect 3734 6574 3933 6630
rect 3989 6574 4075 6630
rect 4131 6574 4338 6630
rect 4394 6574 4480 6630
rect 4536 6574 4738 6630
rect 4794 6574 4880 6630
rect 4936 6574 5143 6630
rect 5199 6574 5285 6630
rect 5341 6574 5540 6630
rect 5596 6574 5682 6630
rect 5738 6574 5937 6630
rect 5993 6574 6079 6630
rect 6135 6574 6340 6630
rect 6396 6574 6482 6630
rect 6538 6574 6742 6630
rect 6798 6574 6884 6630
rect 6940 6574 7145 6630
rect 7201 6574 7287 6630
rect 7343 6574 7539 6630
rect 7595 6574 7681 6630
rect 7737 6574 7940 6630
rect 7996 6574 8082 6630
rect 8138 6574 8340 6630
rect 8396 6574 8482 6630
rect 8538 6574 8737 6630
rect 8793 6574 8879 6630
rect 8935 6574 9134 6630
rect 9190 6574 9276 6630
rect 9332 6574 9538 6630
rect 9594 6574 9680 6630
rect 9736 6574 9934 6630
rect 9990 6574 10076 6630
rect 10132 6574 10334 6630
rect 10390 6574 10476 6630
rect 10532 6574 10731 6630
rect 10787 6574 10873 6630
rect 10929 6574 11136 6630
rect 11192 6574 11278 6630
rect 11334 6574 11536 6630
rect 11592 6574 11678 6630
rect 11734 6574 11941 6630
rect 11997 6574 12083 6630
rect 12139 6598 12526 6630
rect 12582 6598 12650 6654
rect 12706 6598 12774 6654
rect 12830 6598 12898 6654
rect 12954 6598 13022 6654
rect 13078 6598 13200 6654
rect 12139 6574 13200 6598
rect -400 6530 13200 6574
rect -400 6474 -286 6530
rect -230 6474 -162 6530
rect -106 6474 -38 6530
rect 18 6474 86 6530
rect 142 6474 210 6530
rect 266 6488 12526 6530
rect 266 6474 741 6488
rect -400 6432 741 6474
rect 797 6432 883 6488
rect 939 6432 1142 6488
rect 1198 6432 1284 6488
rect 1340 6432 1542 6488
rect 1598 6432 1684 6488
rect 1740 6432 1939 6488
rect 1995 6432 2081 6488
rect 2137 6432 2336 6488
rect 2392 6432 2478 6488
rect 2534 6432 2740 6488
rect 2796 6432 2882 6488
rect 2938 6432 3136 6488
rect 3192 6432 3278 6488
rect 3334 6432 3536 6488
rect 3592 6432 3678 6488
rect 3734 6432 3933 6488
rect 3989 6432 4075 6488
rect 4131 6432 4338 6488
rect 4394 6432 4480 6488
rect 4536 6432 4738 6488
rect 4794 6432 4880 6488
rect 4936 6432 5143 6488
rect 5199 6432 5285 6488
rect 5341 6432 5540 6488
rect 5596 6432 5682 6488
rect 5738 6432 5937 6488
rect 5993 6432 6079 6488
rect 6135 6432 6340 6488
rect 6396 6432 6482 6488
rect 6538 6432 6742 6488
rect 6798 6432 6884 6488
rect 6940 6432 7145 6488
rect 7201 6432 7287 6488
rect 7343 6432 7539 6488
rect 7595 6432 7681 6488
rect 7737 6432 7940 6488
rect 7996 6432 8082 6488
rect 8138 6432 8340 6488
rect 8396 6432 8482 6488
rect 8538 6432 8737 6488
rect 8793 6432 8879 6488
rect 8935 6432 9134 6488
rect 9190 6432 9276 6488
rect 9332 6432 9538 6488
rect 9594 6432 9680 6488
rect 9736 6432 9934 6488
rect 9990 6432 10076 6488
rect 10132 6432 10334 6488
rect 10390 6432 10476 6488
rect 10532 6432 10731 6488
rect 10787 6432 10873 6488
rect 10929 6432 11136 6488
rect 11192 6432 11278 6488
rect 11334 6432 11536 6488
rect 11592 6432 11678 6488
rect 11734 6432 11941 6488
rect 11997 6432 12083 6488
rect 12139 6474 12526 6488
rect 12582 6474 12650 6530
rect 12706 6474 12774 6530
rect 12830 6474 12898 6530
rect 12954 6474 13022 6530
rect 13078 6474 13200 6530
rect 12139 6432 13200 6474
rect -400 6406 13200 6432
rect -400 6350 -286 6406
rect -230 6350 -162 6406
rect -106 6350 -38 6406
rect 18 6350 86 6406
rect 142 6350 210 6406
rect 266 6350 12526 6406
rect 12582 6350 12650 6406
rect 12706 6350 12774 6406
rect 12830 6350 12898 6406
rect 12954 6350 13022 6406
rect 13078 6350 13200 6406
rect -400 6346 13200 6350
rect -400 6290 741 6346
rect 797 6290 883 6346
rect 939 6290 1142 6346
rect 1198 6290 1284 6346
rect 1340 6290 1542 6346
rect 1598 6290 1684 6346
rect 1740 6290 1939 6346
rect 1995 6290 2081 6346
rect 2137 6290 2336 6346
rect 2392 6290 2478 6346
rect 2534 6290 2740 6346
rect 2796 6290 2882 6346
rect 2938 6290 3136 6346
rect 3192 6290 3278 6346
rect 3334 6290 3536 6346
rect 3592 6290 3678 6346
rect 3734 6290 3933 6346
rect 3989 6290 4075 6346
rect 4131 6290 4338 6346
rect 4394 6290 4480 6346
rect 4536 6290 4738 6346
rect 4794 6290 4880 6346
rect 4936 6290 5143 6346
rect 5199 6290 5285 6346
rect 5341 6290 5540 6346
rect 5596 6290 5682 6346
rect 5738 6290 5937 6346
rect 5993 6290 6079 6346
rect 6135 6290 6340 6346
rect 6396 6290 6482 6346
rect 6538 6290 6742 6346
rect 6798 6290 6884 6346
rect 6940 6290 7145 6346
rect 7201 6290 7287 6346
rect 7343 6290 7539 6346
rect 7595 6290 7681 6346
rect 7737 6290 7940 6346
rect 7996 6290 8082 6346
rect 8138 6290 8340 6346
rect 8396 6290 8482 6346
rect 8538 6290 8737 6346
rect 8793 6290 8879 6346
rect 8935 6290 9134 6346
rect 9190 6290 9276 6346
rect 9332 6290 9538 6346
rect 9594 6290 9680 6346
rect 9736 6290 9934 6346
rect 9990 6290 10076 6346
rect 10132 6290 10334 6346
rect 10390 6290 10476 6346
rect 10532 6290 10731 6346
rect 10787 6290 10873 6346
rect 10929 6290 11136 6346
rect 11192 6290 11278 6346
rect 11334 6290 11536 6346
rect 11592 6290 11678 6346
rect 11734 6290 11941 6346
rect 11997 6290 12083 6346
rect 12139 6290 13200 6346
rect -400 6282 13200 6290
rect -400 6226 -286 6282
rect -230 6226 -162 6282
rect -106 6226 -38 6282
rect 18 6226 86 6282
rect 142 6226 210 6282
rect 266 6226 12526 6282
rect 12582 6226 12650 6282
rect 12706 6226 12774 6282
rect 12830 6226 12898 6282
rect 12954 6226 13022 6282
rect 13078 6226 13200 6282
rect -400 6204 13200 6226
rect -400 6158 741 6204
rect -400 6102 -286 6158
rect -230 6102 -162 6158
rect -106 6102 -38 6158
rect 18 6102 86 6158
rect 142 6102 210 6158
rect 266 6148 741 6158
rect 797 6148 883 6204
rect 939 6148 1142 6204
rect 1198 6148 1284 6204
rect 1340 6148 1542 6204
rect 1598 6148 1684 6204
rect 1740 6148 1939 6204
rect 1995 6148 2081 6204
rect 2137 6148 2336 6204
rect 2392 6148 2478 6204
rect 2534 6148 2740 6204
rect 2796 6148 2882 6204
rect 2938 6148 3136 6204
rect 3192 6148 3278 6204
rect 3334 6148 3536 6204
rect 3592 6148 3678 6204
rect 3734 6148 3933 6204
rect 3989 6148 4075 6204
rect 4131 6148 4338 6204
rect 4394 6148 4480 6204
rect 4536 6148 4738 6204
rect 4794 6148 4880 6204
rect 4936 6148 5143 6204
rect 5199 6148 5285 6204
rect 5341 6148 5540 6204
rect 5596 6148 5682 6204
rect 5738 6148 5937 6204
rect 5993 6148 6079 6204
rect 6135 6148 6340 6204
rect 6396 6148 6482 6204
rect 6538 6148 6742 6204
rect 6798 6148 6884 6204
rect 6940 6148 7145 6204
rect 7201 6148 7287 6204
rect 7343 6148 7539 6204
rect 7595 6148 7681 6204
rect 7737 6148 7940 6204
rect 7996 6148 8082 6204
rect 8138 6148 8340 6204
rect 8396 6148 8482 6204
rect 8538 6148 8737 6204
rect 8793 6148 8879 6204
rect 8935 6148 9134 6204
rect 9190 6148 9276 6204
rect 9332 6148 9538 6204
rect 9594 6148 9680 6204
rect 9736 6148 9934 6204
rect 9990 6148 10076 6204
rect 10132 6148 10334 6204
rect 10390 6148 10476 6204
rect 10532 6148 10731 6204
rect 10787 6148 10873 6204
rect 10929 6148 11136 6204
rect 11192 6148 11278 6204
rect 11334 6148 11536 6204
rect 11592 6148 11678 6204
rect 11734 6148 11941 6204
rect 11997 6148 12083 6204
rect 12139 6158 13200 6204
rect 12139 6148 12526 6158
rect 266 6102 12526 6148
rect 12582 6102 12650 6158
rect 12706 6102 12774 6158
rect 12830 6102 12898 6158
rect 12954 6102 13022 6158
rect 13078 6102 13200 6158
rect -400 6062 13200 6102
rect -400 6034 741 6062
rect -400 5978 -286 6034
rect -230 5978 -162 6034
rect -106 5978 -38 6034
rect 18 5978 86 6034
rect 142 5978 210 6034
rect 266 6006 741 6034
rect 797 6006 883 6062
rect 939 6006 1142 6062
rect 1198 6006 1284 6062
rect 1340 6006 1542 6062
rect 1598 6006 1684 6062
rect 1740 6006 1939 6062
rect 1995 6006 2081 6062
rect 2137 6006 2336 6062
rect 2392 6006 2478 6062
rect 2534 6006 2740 6062
rect 2796 6006 2882 6062
rect 2938 6006 3136 6062
rect 3192 6006 3278 6062
rect 3334 6006 3536 6062
rect 3592 6006 3678 6062
rect 3734 6006 3933 6062
rect 3989 6006 4075 6062
rect 4131 6006 4338 6062
rect 4394 6006 4480 6062
rect 4536 6006 4738 6062
rect 4794 6006 4880 6062
rect 4936 6006 5143 6062
rect 5199 6006 5285 6062
rect 5341 6006 5540 6062
rect 5596 6006 5682 6062
rect 5738 6006 5937 6062
rect 5993 6006 6079 6062
rect 6135 6006 6340 6062
rect 6396 6006 6482 6062
rect 6538 6006 6742 6062
rect 6798 6006 6884 6062
rect 6940 6006 7145 6062
rect 7201 6006 7287 6062
rect 7343 6006 7539 6062
rect 7595 6006 7681 6062
rect 7737 6006 7940 6062
rect 7996 6006 8082 6062
rect 8138 6006 8340 6062
rect 8396 6006 8482 6062
rect 8538 6006 8737 6062
rect 8793 6006 8879 6062
rect 8935 6006 9134 6062
rect 9190 6006 9276 6062
rect 9332 6006 9538 6062
rect 9594 6006 9680 6062
rect 9736 6006 9934 6062
rect 9990 6006 10076 6062
rect 10132 6006 10334 6062
rect 10390 6006 10476 6062
rect 10532 6006 10731 6062
rect 10787 6006 10873 6062
rect 10929 6006 11136 6062
rect 11192 6006 11278 6062
rect 11334 6006 11536 6062
rect 11592 6006 11678 6062
rect 11734 6006 11941 6062
rect 11997 6006 12083 6062
rect 12139 6034 13200 6062
rect 12139 6006 12526 6034
rect 266 5978 12526 6006
rect 12582 5978 12650 6034
rect 12706 5978 12774 6034
rect 12830 5978 12898 6034
rect 12954 5978 13022 6034
rect 13078 5978 13200 6034
rect -400 5920 13200 5978
rect -400 5910 741 5920
rect -400 5854 -286 5910
rect -230 5854 -162 5910
rect -106 5854 -38 5910
rect 18 5854 86 5910
rect 142 5854 210 5910
rect 266 5864 741 5910
rect 797 5864 883 5920
rect 939 5864 1142 5920
rect 1198 5864 1284 5920
rect 1340 5864 1542 5920
rect 1598 5864 1684 5920
rect 1740 5864 1939 5920
rect 1995 5864 2081 5920
rect 2137 5864 2336 5920
rect 2392 5864 2478 5920
rect 2534 5864 2740 5920
rect 2796 5864 2882 5920
rect 2938 5864 3136 5920
rect 3192 5864 3278 5920
rect 3334 5864 3536 5920
rect 3592 5864 3678 5920
rect 3734 5864 3933 5920
rect 3989 5864 4075 5920
rect 4131 5864 4338 5920
rect 4394 5864 4480 5920
rect 4536 5864 4738 5920
rect 4794 5864 4880 5920
rect 4936 5864 5143 5920
rect 5199 5864 5285 5920
rect 5341 5864 5540 5920
rect 5596 5864 5682 5920
rect 5738 5864 5937 5920
rect 5993 5864 6079 5920
rect 6135 5864 6340 5920
rect 6396 5864 6482 5920
rect 6538 5864 6742 5920
rect 6798 5864 6884 5920
rect 6940 5864 7145 5920
rect 7201 5864 7287 5920
rect 7343 5864 7539 5920
rect 7595 5864 7681 5920
rect 7737 5864 7940 5920
rect 7996 5864 8082 5920
rect 8138 5864 8340 5920
rect 8396 5864 8482 5920
rect 8538 5864 8737 5920
rect 8793 5864 8879 5920
rect 8935 5864 9134 5920
rect 9190 5864 9276 5920
rect 9332 5864 9538 5920
rect 9594 5864 9680 5920
rect 9736 5864 9934 5920
rect 9990 5864 10076 5920
rect 10132 5864 10334 5920
rect 10390 5864 10476 5920
rect 10532 5864 10731 5920
rect 10787 5864 10873 5920
rect 10929 5864 11136 5920
rect 11192 5864 11278 5920
rect 11334 5864 11536 5920
rect 11592 5864 11678 5920
rect 11734 5864 11941 5920
rect 11997 5864 12083 5920
rect 12139 5910 13200 5920
rect 12139 5864 12526 5910
rect 266 5854 12526 5864
rect 12582 5854 12650 5910
rect 12706 5854 12774 5910
rect 12830 5854 12898 5910
rect 12954 5854 13022 5910
rect 13078 5854 13200 5910
rect -400 5786 13200 5854
rect -400 5730 -286 5786
rect -230 5730 -162 5786
rect -106 5730 -38 5786
rect 18 5730 86 5786
rect 142 5730 210 5786
rect 266 5778 12526 5786
rect 266 5730 741 5778
rect -400 5722 741 5730
rect 797 5722 883 5778
rect 939 5722 1142 5778
rect 1198 5722 1284 5778
rect 1340 5722 1542 5778
rect 1598 5722 1684 5778
rect 1740 5722 1939 5778
rect 1995 5722 2081 5778
rect 2137 5722 2336 5778
rect 2392 5722 2478 5778
rect 2534 5722 2740 5778
rect 2796 5722 2882 5778
rect 2938 5722 3136 5778
rect 3192 5722 3278 5778
rect 3334 5722 3536 5778
rect 3592 5722 3678 5778
rect 3734 5722 3933 5778
rect 3989 5722 4075 5778
rect 4131 5722 4338 5778
rect 4394 5722 4480 5778
rect 4536 5722 4738 5778
rect 4794 5722 4880 5778
rect 4936 5722 5143 5778
rect 5199 5722 5285 5778
rect 5341 5722 5540 5778
rect 5596 5722 5682 5778
rect 5738 5722 5937 5778
rect 5993 5722 6079 5778
rect 6135 5722 6340 5778
rect 6396 5722 6482 5778
rect 6538 5722 6742 5778
rect 6798 5722 6884 5778
rect 6940 5722 7145 5778
rect 7201 5722 7287 5778
rect 7343 5722 7539 5778
rect 7595 5722 7681 5778
rect 7737 5722 7940 5778
rect 7996 5722 8082 5778
rect 8138 5722 8340 5778
rect 8396 5722 8482 5778
rect 8538 5722 8737 5778
rect 8793 5722 8879 5778
rect 8935 5722 9134 5778
rect 9190 5722 9276 5778
rect 9332 5722 9538 5778
rect 9594 5722 9680 5778
rect 9736 5722 9934 5778
rect 9990 5722 10076 5778
rect 10132 5722 10334 5778
rect 10390 5722 10476 5778
rect 10532 5722 10731 5778
rect 10787 5722 10873 5778
rect 10929 5722 11136 5778
rect 11192 5722 11278 5778
rect 11334 5722 11536 5778
rect 11592 5722 11678 5778
rect 11734 5722 11941 5778
rect 11997 5722 12083 5778
rect 12139 5730 12526 5778
rect 12582 5730 12650 5786
rect 12706 5730 12774 5786
rect 12830 5730 12898 5786
rect 12954 5730 13022 5786
rect 13078 5730 13200 5786
rect 12139 5722 13200 5730
rect -400 5662 13200 5722
rect -400 5606 -286 5662
rect -230 5606 -162 5662
rect -106 5606 -38 5662
rect 18 5606 86 5662
rect 142 5606 210 5662
rect 266 5636 12526 5662
rect 266 5606 741 5636
rect -400 5580 741 5606
rect 797 5580 883 5636
rect 939 5580 1142 5636
rect 1198 5580 1284 5636
rect 1340 5580 1542 5636
rect 1598 5580 1684 5636
rect 1740 5580 1939 5636
rect 1995 5580 2081 5636
rect 2137 5580 2336 5636
rect 2392 5580 2478 5636
rect 2534 5580 2740 5636
rect 2796 5580 2882 5636
rect 2938 5580 3136 5636
rect 3192 5580 3278 5636
rect 3334 5580 3536 5636
rect 3592 5580 3678 5636
rect 3734 5580 3933 5636
rect 3989 5580 4075 5636
rect 4131 5580 4338 5636
rect 4394 5580 4480 5636
rect 4536 5580 4738 5636
rect 4794 5580 4880 5636
rect 4936 5580 5143 5636
rect 5199 5580 5285 5636
rect 5341 5580 5540 5636
rect 5596 5580 5682 5636
rect 5738 5580 5937 5636
rect 5993 5580 6079 5636
rect 6135 5580 6340 5636
rect 6396 5580 6482 5636
rect 6538 5580 6742 5636
rect 6798 5580 6884 5636
rect 6940 5580 7145 5636
rect 7201 5580 7287 5636
rect 7343 5580 7539 5636
rect 7595 5580 7681 5636
rect 7737 5580 7940 5636
rect 7996 5580 8082 5636
rect 8138 5580 8340 5636
rect 8396 5580 8482 5636
rect 8538 5580 8737 5636
rect 8793 5580 8879 5636
rect 8935 5580 9134 5636
rect 9190 5580 9276 5636
rect 9332 5580 9538 5636
rect 9594 5580 9680 5636
rect 9736 5580 9934 5636
rect 9990 5580 10076 5636
rect 10132 5580 10334 5636
rect 10390 5580 10476 5636
rect 10532 5580 10731 5636
rect 10787 5580 10873 5636
rect 10929 5580 11136 5636
rect 11192 5580 11278 5636
rect 11334 5580 11536 5636
rect 11592 5580 11678 5636
rect 11734 5580 11941 5636
rect 11997 5580 12083 5636
rect 12139 5606 12526 5636
rect 12582 5606 12650 5662
rect 12706 5606 12774 5662
rect 12830 5606 12898 5662
rect 12954 5606 13022 5662
rect 13078 5606 13200 5662
rect 12139 5580 13200 5606
rect -400 5538 13200 5580
rect -400 5482 -286 5538
rect -230 5482 -162 5538
rect -106 5482 -38 5538
rect 18 5482 86 5538
rect 142 5482 210 5538
rect 266 5494 12526 5538
rect 266 5482 741 5494
rect -400 5438 741 5482
rect 797 5438 883 5494
rect 939 5438 1142 5494
rect 1198 5438 1284 5494
rect 1340 5438 1542 5494
rect 1598 5438 1684 5494
rect 1740 5438 1939 5494
rect 1995 5438 2081 5494
rect 2137 5438 2336 5494
rect 2392 5438 2478 5494
rect 2534 5438 2740 5494
rect 2796 5438 2882 5494
rect 2938 5438 3136 5494
rect 3192 5438 3278 5494
rect 3334 5438 3536 5494
rect 3592 5438 3678 5494
rect 3734 5438 3933 5494
rect 3989 5438 4075 5494
rect 4131 5438 4338 5494
rect 4394 5438 4480 5494
rect 4536 5438 4738 5494
rect 4794 5438 4880 5494
rect 4936 5438 5143 5494
rect 5199 5438 5285 5494
rect 5341 5438 5540 5494
rect 5596 5438 5682 5494
rect 5738 5438 5937 5494
rect 5993 5438 6079 5494
rect 6135 5438 6340 5494
rect 6396 5438 6482 5494
rect 6538 5438 6742 5494
rect 6798 5438 6884 5494
rect 6940 5438 7145 5494
rect 7201 5438 7287 5494
rect 7343 5438 7539 5494
rect 7595 5438 7681 5494
rect 7737 5438 7940 5494
rect 7996 5438 8082 5494
rect 8138 5438 8340 5494
rect 8396 5438 8482 5494
rect 8538 5438 8737 5494
rect 8793 5438 8879 5494
rect 8935 5438 9134 5494
rect 9190 5438 9276 5494
rect 9332 5438 9538 5494
rect 9594 5438 9680 5494
rect 9736 5438 9934 5494
rect 9990 5438 10076 5494
rect 10132 5438 10334 5494
rect 10390 5438 10476 5494
rect 10532 5438 10731 5494
rect 10787 5438 10873 5494
rect 10929 5438 11136 5494
rect 11192 5438 11278 5494
rect 11334 5438 11536 5494
rect 11592 5438 11678 5494
rect 11734 5438 11941 5494
rect 11997 5438 12083 5494
rect 12139 5482 12526 5494
rect 12582 5482 12650 5538
rect 12706 5482 12774 5538
rect 12830 5482 12898 5538
rect 12954 5482 13022 5538
rect 13078 5482 13200 5538
rect 12139 5438 13200 5482
rect -400 5414 13200 5438
rect -400 5358 -286 5414
rect -230 5358 -162 5414
rect -106 5358 -38 5414
rect 18 5358 86 5414
rect 142 5358 210 5414
rect 266 5358 12526 5414
rect 12582 5358 12650 5414
rect 12706 5358 12774 5414
rect 12830 5358 12898 5414
rect 12954 5358 13022 5414
rect 13078 5358 13200 5414
rect -400 5352 13200 5358
rect -400 5296 741 5352
rect 797 5296 883 5352
rect 939 5296 1142 5352
rect 1198 5296 1284 5352
rect 1340 5296 1542 5352
rect 1598 5296 1684 5352
rect 1740 5296 1939 5352
rect 1995 5296 2081 5352
rect 2137 5296 2336 5352
rect 2392 5296 2478 5352
rect 2534 5296 2740 5352
rect 2796 5296 2882 5352
rect 2938 5296 3136 5352
rect 3192 5296 3278 5352
rect 3334 5296 3536 5352
rect 3592 5296 3678 5352
rect 3734 5296 3933 5352
rect 3989 5296 4075 5352
rect 4131 5296 4338 5352
rect 4394 5296 4480 5352
rect 4536 5296 4738 5352
rect 4794 5296 4880 5352
rect 4936 5296 5143 5352
rect 5199 5296 5285 5352
rect 5341 5296 5540 5352
rect 5596 5296 5682 5352
rect 5738 5296 5937 5352
rect 5993 5296 6079 5352
rect 6135 5296 6340 5352
rect 6396 5296 6482 5352
rect 6538 5296 6742 5352
rect 6798 5296 6884 5352
rect 6940 5296 7145 5352
rect 7201 5296 7287 5352
rect 7343 5296 7539 5352
rect 7595 5296 7681 5352
rect 7737 5296 7940 5352
rect 7996 5296 8082 5352
rect 8138 5296 8340 5352
rect 8396 5296 8482 5352
rect 8538 5296 8737 5352
rect 8793 5296 8879 5352
rect 8935 5296 9134 5352
rect 9190 5296 9276 5352
rect 9332 5296 9538 5352
rect 9594 5296 9680 5352
rect 9736 5296 9934 5352
rect 9990 5296 10076 5352
rect 10132 5296 10334 5352
rect 10390 5296 10476 5352
rect 10532 5296 10731 5352
rect 10787 5296 10873 5352
rect 10929 5296 11136 5352
rect 11192 5296 11278 5352
rect 11334 5296 11536 5352
rect 11592 5296 11678 5352
rect 11734 5296 11941 5352
rect 11997 5296 12083 5352
rect 12139 5296 13200 5352
rect -400 5290 13200 5296
rect -400 5234 -286 5290
rect -230 5234 -162 5290
rect -106 5234 -38 5290
rect 18 5234 86 5290
rect 142 5234 210 5290
rect 266 5234 12526 5290
rect 12582 5234 12650 5290
rect 12706 5234 12774 5290
rect 12830 5234 12898 5290
rect 12954 5234 13022 5290
rect 13078 5234 13200 5290
rect -400 5210 13200 5234
rect -400 5166 741 5210
rect -400 5110 -286 5166
rect -230 5110 -162 5166
rect -106 5110 -38 5166
rect 18 5110 86 5166
rect 142 5110 210 5166
rect 266 5154 741 5166
rect 797 5154 883 5210
rect 939 5154 1142 5210
rect 1198 5154 1284 5210
rect 1340 5154 1542 5210
rect 1598 5154 1684 5210
rect 1740 5154 1939 5210
rect 1995 5154 2081 5210
rect 2137 5154 2336 5210
rect 2392 5154 2478 5210
rect 2534 5154 2740 5210
rect 2796 5154 2882 5210
rect 2938 5154 3136 5210
rect 3192 5154 3278 5210
rect 3334 5154 3536 5210
rect 3592 5154 3678 5210
rect 3734 5154 3933 5210
rect 3989 5154 4075 5210
rect 4131 5154 4338 5210
rect 4394 5154 4480 5210
rect 4536 5154 4738 5210
rect 4794 5154 4880 5210
rect 4936 5154 5143 5210
rect 5199 5154 5285 5210
rect 5341 5154 5540 5210
rect 5596 5154 5682 5210
rect 5738 5154 5937 5210
rect 5993 5154 6079 5210
rect 6135 5154 6340 5210
rect 6396 5154 6482 5210
rect 6538 5154 6742 5210
rect 6798 5154 6884 5210
rect 6940 5154 7145 5210
rect 7201 5154 7287 5210
rect 7343 5154 7539 5210
rect 7595 5154 7681 5210
rect 7737 5154 7940 5210
rect 7996 5154 8082 5210
rect 8138 5154 8340 5210
rect 8396 5154 8482 5210
rect 8538 5154 8737 5210
rect 8793 5154 8879 5210
rect 8935 5154 9134 5210
rect 9190 5154 9276 5210
rect 9332 5154 9538 5210
rect 9594 5154 9680 5210
rect 9736 5154 9934 5210
rect 9990 5154 10076 5210
rect 10132 5154 10334 5210
rect 10390 5154 10476 5210
rect 10532 5154 10731 5210
rect 10787 5154 10873 5210
rect 10929 5154 11136 5210
rect 11192 5154 11278 5210
rect 11334 5154 11536 5210
rect 11592 5154 11678 5210
rect 11734 5154 11941 5210
rect 11997 5154 12083 5210
rect 12139 5166 13200 5210
rect 12139 5154 12526 5166
rect 266 5110 12526 5154
rect 12582 5110 12650 5166
rect 12706 5110 12774 5166
rect 12830 5110 12898 5166
rect 12954 5110 13022 5166
rect 13078 5110 13200 5166
rect -400 5068 13200 5110
rect -400 5042 741 5068
rect -400 4986 -286 5042
rect -230 4986 -162 5042
rect -106 4986 -38 5042
rect 18 4986 86 5042
rect 142 4986 210 5042
rect 266 5012 741 5042
rect 797 5012 883 5068
rect 939 5012 1142 5068
rect 1198 5012 1284 5068
rect 1340 5012 1542 5068
rect 1598 5012 1684 5068
rect 1740 5012 1939 5068
rect 1995 5012 2081 5068
rect 2137 5012 2336 5068
rect 2392 5012 2478 5068
rect 2534 5012 2740 5068
rect 2796 5012 2882 5068
rect 2938 5012 3136 5068
rect 3192 5012 3278 5068
rect 3334 5012 3536 5068
rect 3592 5012 3678 5068
rect 3734 5012 3933 5068
rect 3989 5012 4075 5068
rect 4131 5012 4338 5068
rect 4394 5012 4480 5068
rect 4536 5012 4738 5068
rect 4794 5012 4880 5068
rect 4936 5012 5143 5068
rect 5199 5012 5285 5068
rect 5341 5012 5540 5068
rect 5596 5012 5682 5068
rect 5738 5012 5937 5068
rect 5993 5012 6079 5068
rect 6135 5012 6340 5068
rect 6396 5012 6482 5068
rect 6538 5012 6742 5068
rect 6798 5012 6884 5068
rect 6940 5012 7145 5068
rect 7201 5012 7287 5068
rect 7343 5012 7539 5068
rect 7595 5012 7681 5068
rect 7737 5012 7940 5068
rect 7996 5012 8082 5068
rect 8138 5012 8340 5068
rect 8396 5012 8482 5068
rect 8538 5012 8737 5068
rect 8793 5012 8879 5068
rect 8935 5012 9134 5068
rect 9190 5012 9276 5068
rect 9332 5012 9538 5068
rect 9594 5012 9680 5068
rect 9736 5012 9934 5068
rect 9990 5012 10076 5068
rect 10132 5012 10334 5068
rect 10390 5012 10476 5068
rect 10532 5012 10731 5068
rect 10787 5012 10873 5068
rect 10929 5012 11136 5068
rect 11192 5012 11278 5068
rect 11334 5012 11536 5068
rect 11592 5012 11678 5068
rect 11734 5012 11941 5068
rect 11997 5012 12083 5068
rect 12139 5042 13200 5068
rect 12139 5012 12526 5042
rect 266 4986 12526 5012
rect 12582 4986 12650 5042
rect 12706 4986 12774 5042
rect 12830 4986 12898 5042
rect 12954 4986 13022 5042
rect 13078 4986 13200 5042
rect -400 4926 13200 4986
rect -400 4918 741 4926
rect -400 4862 -286 4918
rect -230 4862 -162 4918
rect -106 4862 -38 4918
rect 18 4862 86 4918
rect 142 4862 210 4918
rect 266 4870 741 4918
rect 797 4870 883 4926
rect 939 4870 1142 4926
rect 1198 4870 1284 4926
rect 1340 4870 1542 4926
rect 1598 4870 1684 4926
rect 1740 4870 1939 4926
rect 1995 4870 2081 4926
rect 2137 4870 2336 4926
rect 2392 4870 2478 4926
rect 2534 4870 2740 4926
rect 2796 4870 2882 4926
rect 2938 4870 3136 4926
rect 3192 4870 3278 4926
rect 3334 4870 3536 4926
rect 3592 4870 3678 4926
rect 3734 4870 3933 4926
rect 3989 4870 4075 4926
rect 4131 4870 4338 4926
rect 4394 4870 4480 4926
rect 4536 4870 4738 4926
rect 4794 4870 4880 4926
rect 4936 4870 5143 4926
rect 5199 4870 5285 4926
rect 5341 4870 5540 4926
rect 5596 4870 5682 4926
rect 5738 4870 5937 4926
rect 5993 4870 6079 4926
rect 6135 4870 6340 4926
rect 6396 4870 6482 4926
rect 6538 4870 6742 4926
rect 6798 4870 6884 4926
rect 6940 4870 7145 4926
rect 7201 4870 7287 4926
rect 7343 4870 7539 4926
rect 7595 4870 7681 4926
rect 7737 4870 7940 4926
rect 7996 4870 8082 4926
rect 8138 4870 8340 4926
rect 8396 4870 8482 4926
rect 8538 4870 8737 4926
rect 8793 4870 8879 4926
rect 8935 4870 9134 4926
rect 9190 4870 9276 4926
rect 9332 4870 9538 4926
rect 9594 4870 9680 4926
rect 9736 4870 9934 4926
rect 9990 4870 10076 4926
rect 10132 4870 10334 4926
rect 10390 4870 10476 4926
rect 10532 4870 10731 4926
rect 10787 4870 10873 4926
rect 10929 4870 11136 4926
rect 11192 4870 11278 4926
rect 11334 4870 11536 4926
rect 11592 4870 11678 4926
rect 11734 4870 11941 4926
rect 11997 4870 12083 4926
rect 12139 4918 13200 4926
rect 12139 4870 12526 4918
rect 266 4862 12526 4870
rect 12582 4862 12650 4918
rect 12706 4862 12774 4918
rect 12830 4862 12898 4918
rect 12954 4862 13022 4918
rect 13078 4862 13200 4918
rect -400 4794 13200 4862
rect -400 4738 -286 4794
rect -230 4738 -162 4794
rect -106 4738 -38 4794
rect 18 4738 86 4794
rect 142 4738 210 4794
rect 266 4784 12526 4794
rect 266 4738 741 4784
rect -400 4728 741 4738
rect 797 4728 883 4784
rect 939 4728 1142 4784
rect 1198 4728 1284 4784
rect 1340 4728 1542 4784
rect 1598 4728 1684 4784
rect 1740 4728 1939 4784
rect 1995 4728 2081 4784
rect 2137 4728 2336 4784
rect 2392 4728 2478 4784
rect 2534 4728 2740 4784
rect 2796 4728 2882 4784
rect 2938 4728 3136 4784
rect 3192 4728 3278 4784
rect 3334 4728 3536 4784
rect 3592 4728 3678 4784
rect 3734 4728 3933 4784
rect 3989 4728 4075 4784
rect 4131 4728 4338 4784
rect 4394 4728 4480 4784
rect 4536 4728 4738 4784
rect 4794 4728 4880 4784
rect 4936 4728 5143 4784
rect 5199 4728 5285 4784
rect 5341 4728 5540 4784
rect 5596 4728 5682 4784
rect 5738 4728 5937 4784
rect 5993 4728 6079 4784
rect 6135 4728 6340 4784
rect 6396 4728 6482 4784
rect 6538 4728 6742 4784
rect 6798 4728 6884 4784
rect 6940 4728 7145 4784
rect 7201 4728 7287 4784
rect 7343 4728 7539 4784
rect 7595 4728 7681 4784
rect 7737 4728 7940 4784
rect 7996 4728 8082 4784
rect 8138 4728 8340 4784
rect 8396 4728 8482 4784
rect 8538 4728 8737 4784
rect 8793 4728 8879 4784
rect 8935 4728 9134 4784
rect 9190 4728 9276 4784
rect 9332 4728 9538 4784
rect 9594 4728 9680 4784
rect 9736 4728 9934 4784
rect 9990 4728 10076 4784
rect 10132 4728 10334 4784
rect 10390 4728 10476 4784
rect 10532 4728 10731 4784
rect 10787 4728 10873 4784
rect 10929 4728 11136 4784
rect 11192 4728 11278 4784
rect 11334 4728 11536 4784
rect 11592 4728 11678 4784
rect 11734 4728 11941 4784
rect 11997 4728 12083 4784
rect 12139 4738 12526 4784
rect 12582 4738 12650 4794
rect 12706 4738 12774 4794
rect 12830 4738 12898 4794
rect 12954 4738 13022 4794
rect 13078 4738 13200 4794
rect 12139 4728 13200 4738
rect -400 4670 13200 4728
rect -400 4614 -286 4670
rect -230 4614 -162 4670
rect -106 4614 -38 4670
rect 18 4614 86 4670
rect 142 4614 210 4670
rect 266 4642 12526 4670
rect 266 4614 741 4642
rect -400 4586 741 4614
rect 797 4586 883 4642
rect 939 4586 1142 4642
rect 1198 4586 1284 4642
rect 1340 4586 1542 4642
rect 1598 4586 1684 4642
rect 1740 4586 1939 4642
rect 1995 4586 2081 4642
rect 2137 4586 2336 4642
rect 2392 4586 2478 4642
rect 2534 4586 2740 4642
rect 2796 4586 2882 4642
rect 2938 4586 3136 4642
rect 3192 4586 3278 4642
rect 3334 4586 3536 4642
rect 3592 4586 3678 4642
rect 3734 4586 3933 4642
rect 3989 4586 4075 4642
rect 4131 4586 4338 4642
rect 4394 4586 4480 4642
rect 4536 4586 4738 4642
rect 4794 4586 4880 4642
rect 4936 4586 5143 4642
rect 5199 4586 5285 4642
rect 5341 4586 5540 4642
rect 5596 4586 5682 4642
rect 5738 4586 5937 4642
rect 5993 4586 6079 4642
rect 6135 4586 6340 4642
rect 6396 4586 6482 4642
rect 6538 4586 6742 4642
rect 6798 4586 6884 4642
rect 6940 4586 7145 4642
rect 7201 4586 7287 4642
rect 7343 4586 7539 4642
rect 7595 4586 7681 4642
rect 7737 4586 7940 4642
rect 7996 4586 8082 4642
rect 8138 4586 8340 4642
rect 8396 4586 8482 4642
rect 8538 4586 8737 4642
rect 8793 4586 8879 4642
rect 8935 4586 9134 4642
rect 9190 4586 9276 4642
rect 9332 4586 9538 4642
rect 9594 4586 9680 4642
rect 9736 4586 9934 4642
rect 9990 4586 10076 4642
rect 10132 4586 10334 4642
rect 10390 4586 10476 4642
rect 10532 4586 10731 4642
rect 10787 4586 10873 4642
rect 10929 4586 11136 4642
rect 11192 4586 11278 4642
rect 11334 4586 11536 4642
rect 11592 4586 11678 4642
rect 11734 4586 11941 4642
rect 11997 4586 12083 4642
rect 12139 4614 12526 4642
rect 12582 4614 12650 4670
rect 12706 4614 12774 4670
rect 12830 4614 12898 4670
rect 12954 4614 13022 4670
rect 13078 4614 13200 4670
rect 12139 4586 13200 4614
rect -400 4546 13200 4586
rect -400 4490 -286 4546
rect -230 4490 -162 4546
rect -106 4490 -38 4546
rect 18 4490 86 4546
rect 142 4490 210 4546
rect 266 4500 12526 4546
rect 266 4490 741 4500
rect -400 4444 741 4490
rect 797 4444 883 4500
rect 939 4444 1142 4500
rect 1198 4444 1284 4500
rect 1340 4444 1542 4500
rect 1598 4444 1684 4500
rect 1740 4444 1939 4500
rect 1995 4444 2081 4500
rect 2137 4444 2336 4500
rect 2392 4444 2478 4500
rect 2534 4444 2740 4500
rect 2796 4444 2882 4500
rect 2938 4444 3136 4500
rect 3192 4444 3278 4500
rect 3334 4444 3536 4500
rect 3592 4444 3678 4500
rect 3734 4444 3933 4500
rect 3989 4444 4075 4500
rect 4131 4444 4338 4500
rect 4394 4444 4480 4500
rect 4536 4444 4738 4500
rect 4794 4444 4880 4500
rect 4936 4444 5143 4500
rect 5199 4444 5285 4500
rect 5341 4444 5540 4500
rect 5596 4444 5682 4500
rect 5738 4444 5937 4500
rect 5993 4444 6079 4500
rect 6135 4444 6340 4500
rect 6396 4444 6482 4500
rect 6538 4444 6742 4500
rect 6798 4444 6884 4500
rect 6940 4444 7145 4500
rect 7201 4444 7287 4500
rect 7343 4444 7539 4500
rect 7595 4444 7681 4500
rect 7737 4444 7940 4500
rect 7996 4444 8082 4500
rect 8138 4444 8340 4500
rect 8396 4444 8482 4500
rect 8538 4444 8737 4500
rect 8793 4444 8879 4500
rect 8935 4444 9134 4500
rect 9190 4444 9276 4500
rect 9332 4444 9538 4500
rect 9594 4444 9680 4500
rect 9736 4444 9934 4500
rect 9990 4444 10076 4500
rect 10132 4444 10334 4500
rect 10390 4444 10476 4500
rect 10532 4444 10731 4500
rect 10787 4444 10873 4500
rect 10929 4444 11136 4500
rect 11192 4444 11278 4500
rect 11334 4444 11536 4500
rect 11592 4444 11678 4500
rect 11734 4444 11941 4500
rect 11997 4444 12083 4500
rect 12139 4490 12526 4500
rect 12582 4490 12650 4546
rect 12706 4490 12774 4546
rect 12830 4490 12898 4546
rect 12954 4490 13022 4546
rect 13078 4490 13200 4546
rect 12139 4444 13200 4490
rect -400 4422 13200 4444
rect -400 4366 -286 4422
rect -230 4366 -162 4422
rect -106 4366 -38 4422
rect 18 4366 86 4422
rect 142 4366 210 4422
rect 266 4366 12526 4422
rect 12582 4366 12650 4422
rect 12706 4366 12774 4422
rect 12830 4366 12898 4422
rect 12954 4366 13022 4422
rect 13078 4366 13200 4422
rect -400 4358 13200 4366
rect -400 4302 741 4358
rect 797 4302 883 4358
rect 939 4302 1142 4358
rect 1198 4302 1284 4358
rect 1340 4302 1542 4358
rect 1598 4302 1684 4358
rect 1740 4302 1939 4358
rect 1995 4302 2081 4358
rect 2137 4302 2336 4358
rect 2392 4302 2478 4358
rect 2534 4302 2740 4358
rect 2796 4302 2882 4358
rect 2938 4302 3136 4358
rect 3192 4302 3278 4358
rect 3334 4302 3536 4358
rect 3592 4302 3678 4358
rect 3734 4302 3933 4358
rect 3989 4302 4075 4358
rect 4131 4302 4338 4358
rect 4394 4302 4480 4358
rect 4536 4302 4738 4358
rect 4794 4302 4880 4358
rect 4936 4302 5143 4358
rect 5199 4302 5285 4358
rect 5341 4302 5540 4358
rect 5596 4302 5682 4358
rect 5738 4302 5937 4358
rect 5993 4302 6079 4358
rect 6135 4302 6340 4358
rect 6396 4302 6482 4358
rect 6538 4302 6742 4358
rect 6798 4302 6884 4358
rect 6940 4302 7145 4358
rect 7201 4302 7287 4358
rect 7343 4302 7539 4358
rect 7595 4302 7681 4358
rect 7737 4302 7940 4358
rect 7996 4302 8082 4358
rect 8138 4302 8340 4358
rect 8396 4302 8482 4358
rect 8538 4302 8737 4358
rect 8793 4302 8879 4358
rect 8935 4302 9134 4358
rect 9190 4302 9276 4358
rect 9332 4302 9538 4358
rect 9594 4302 9680 4358
rect 9736 4302 9934 4358
rect 9990 4302 10076 4358
rect 10132 4302 10334 4358
rect 10390 4302 10476 4358
rect 10532 4302 10731 4358
rect 10787 4302 10873 4358
rect 10929 4302 11136 4358
rect 11192 4302 11278 4358
rect 11334 4302 11536 4358
rect 11592 4302 11678 4358
rect 11734 4302 11941 4358
rect 11997 4302 12083 4358
rect 12139 4302 13200 4358
rect -400 4298 13200 4302
rect -400 4242 -286 4298
rect -230 4242 -162 4298
rect -106 4242 -38 4298
rect 18 4242 86 4298
rect 142 4242 210 4298
rect 266 4242 12526 4298
rect 12582 4242 12650 4298
rect 12706 4242 12774 4298
rect 12830 4242 12898 4298
rect 12954 4242 13022 4298
rect 13078 4242 13200 4298
rect -400 4216 13200 4242
rect -400 4174 741 4216
rect -400 4118 -286 4174
rect -230 4118 -162 4174
rect -106 4118 -38 4174
rect 18 4118 86 4174
rect 142 4118 210 4174
rect 266 4160 741 4174
rect 797 4160 883 4216
rect 939 4160 1142 4216
rect 1198 4160 1284 4216
rect 1340 4160 1542 4216
rect 1598 4160 1684 4216
rect 1740 4160 1939 4216
rect 1995 4160 2081 4216
rect 2137 4160 2336 4216
rect 2392 4160 2478 4216
rect 2534 4160 2740 4216
rect 2796 4160 2882 4216
rect 2938 4160 3136 4216
rect 3192 4160 3278 4216
rect 3334 4160 3536 4216
rect 3592 4160 3678 4216
rect 3734 4160 3933 4216
rect 3989 4160 4075 4216
rect 4131 4160 4338 4216
rect 4394 4160 4480 4216
rect 4536 4160 4738 4216
rect 4794 4160 4880 4216
rect 4936 4160 5143 4216
rect 5199 4160 5285 4216
rect 5341 4160 5540 4216
rect 5596 4160 5682 4216
rect 5738 4160 5937 4216
rect 5993 4160 6079 4216
rect 6135 4160 6340 4216
rect 6396 4160 6482 4216
rect 6538 4160 6742 4216
rect 6798 4160 6884 4216
rect 6940 4160 7145 4216
rect 7201 4160 7287 4216
rect 7343 4160 7539 4216
rect 7595 4160 7681 4216
rect 7737 4160 7940 4216
rect 7996 4160 8082 4216
rect 8138 4160 8340 4216
rect 8396 4160 8482 4216
rect 8538 4160 8737 4216
rect 8793 4160 8879 4216
rect 8935 4160 9134 4216
rect 9190 4160 9276 4216
rect 9332 4160 9538 4216
rect 9594 4160 9680 4216
rect 9736 4160 9934 4216
rect 9990 4160 10076 4216
rect 10132 4160 10334 4216
rect 10390 4160 10476 4216
rect 10532 4160 10731 4216
rect 10787 4160 10873 4216
rect 10929 4160 11136 4216
rect 11192 4160 11278 4216
rect 11334 4160 11536 4216
rect 11592 4160 11678 4216
rect 11734 4160 11941 4216
rect 11997 4160 12083 4216
rect 12139 4174 13200 4216
rect 12139 4160 12526 4174
rect 266 4118 12526 4160
rect 12582 4118 12650 4174
rect 12706 4118 12774 4174
rect 12830 4118 12898 4174
rect 12954 4118 13022 4174
rect 13078 4118 13200 4174
rect -400 4074 13200 4118
rect -400 4050 741 4074
rect -400 3994 -286 4050
rect -230 3994 -162 4050
rect -106 3994 -38 4050
rect 18 3994 86 4050
rect 142 3994 210 4050
rect 266 4018 741 4050
rect 797 4018 883 4074
rect 939 4018 1142 4074
rect 1198 4018 1284 4074
rect 1340 4018 1542 4074
rect 1598 4018 1684 4074
rect 1740 4018 1939 4074
rect 1995 4018 2081 4074
rect 2137 4018 2336 4074
rect 2392 4018 2478 4074
rect 2534 4018 2740 4074
rect 2796 4018 2882 4074
rect 2938 4018 3136 4074
rect 3192 4018 3278 4074
rect 3334 4018 3536 4074
rect 3592 4018 3678 4074
rect 3734 4018 3933 4074
rect 3989 4018 4075 4074
rect 4131 4018 4338 4074
rect 4394 4018 4480 4074
rect 4536 4018 4738 4074
rect 4794 4018 4880 4074
rect 4936 4018 5143 4074
rect 5199 4018 5285 4074
rect 5341 4018 5540 4074
rect 5596 4018 5682 4074
rect 5738 4018 5937 4074
rect 5993 4018 6079 4074
rect 6135 4018 6340 4074
rect 6396 4018 6482 4074
rect 6538 4018 6742 4074
rect 6798 4018 6884 4074
rect 6940 4018 7145 4074
rect 7201 4018 7287 4074
rect 7343 4018 7539 4074
rect 7595 4018 7681 4074
rect 7737 4018 7940 4074
rect 7996 4018 8082 4074
rect 8138 4018 8340 4074
rect 8396 4018 8482 4074
rect 8538 4018 8737 4074
rect 8793 4018 8879 4074
rect 8935 4018 9134 4074
rect 9190 4018 9276 4074
rect 9332 4018 9538 4074
rect 9594 4018 9680 4074
rect 9736 4018 9934 4074
rect 9990 4018 10076 4074
rect 10132 4018 10334 4074
rect 10390 4018 10476 4074
rect 10532 4018 10731 4074
rect 10787 4018 10873 4074
rect 10929 4018 11136 4074
rect 11192 4018 11278 4074
rect 11334 4018 11536 4074
rect 11592 4018 11678 4074
rect 11734 4018 11941 4074
rect 11997 4018 12083 4074
rect 12139 4050 13200 4074
rect 12139 4018 12526 4050
rect 266 3994 12526 4018
rect 12582 3994 12650 4050
rect 12706 3994 12774 4050
rect 12830 3994 12898 4050
rect 12954 3994 13022 4050
rect 13078 3994 13200 4050
rect -400 3932 13200 3994
rect -400 3926 741 3932
rect -400 3870 -286 3926
rect -230 3870 -162 3926
rect -106 3870 -38 3926
rect 18 3870 86 3926
rect 142 3870 210 3926
rect 266 3876 741 3926
rect 797 3876 883 3932
rect 939 3876 1142 3932
rect 1198 3876 1284 3932
rect 1340 3876 1542 3932
rect 1598 3876 1684 3932
rect 1740 3876 1939 3932
rect 1995 3876 2081 3932
rect 2137 3876 2336 3932
rect 2392 3876 2478 3932
rect 2534 3876 2740 3932
rect 2796 3876 2882 3932
rect 2938 3876 3136 3932
rect 3192 3876 3278 3932
rect 3334 3876 3536 3932
rect 3592 3876 3678 3932
rect 3734 3876 3933 3932
rect 3989 3876 4075 3932
rect 4131 3876 4338 3932
rect 4394 3876 4480 3932
rect 4536 3876 4738 3932
rect 4794 3876 4880 3932
rect 4936 3876 5143 3932
rect 5199 3876 5285 3932
rect 5341 3876 5540 3932
rect 5596 3876 5682 3932
rect 5738 3876 5937 3932
rect 5993 3876 6079 3932
rect 6135 3876 6340 3932
rect 6396 3876 6482 3932
rect 6538 3876 6742 3932
rect 6798 3876 6884 3932
rect 6940 3876 7145 3932
rect 7201 3876 7287 3932
rect 7343 3876 7539 3932
rect 7595 3876 7681 3932
rect 7737 3876 7940 3932
rect 7996 3876 8082 3932
rect 8138 3876 8340 3932
rect 8396 3876 8482 3932
rect 8538 3876 8737 3932
rect 8793 3876 8879 3932
rect 8935 3876 9134 3932
rect 9190 3876 9276 3932
rect 9332 3876 9538 3932
rect 9594 3876 9680 3932
rect 9736 3876 9934 3932
rect 9990 3876 10076 3932
rect 10132 3876 10334 3932
rect 10390 3876 10476 3932
rect 10532 3876 10731 3932
rect 10787 3876 10873 3932
rect 10929 3876 11136 3932
rect 11192 3876 11278 3932
rect 11334 3876 11536 3932
rect 11592 3876 11678 3932
rect 11734 3876 11941 3932
rect 11997 3876 12083 3932
rect 12139 3926 13200 3932
rect 12139 3876 12526 3926
rect 266 3870 12526 3876
rect 12582 3870 12650 3926
rect 12706 3870 12774 3926
rect 12830 3870 12898 3926
rect 12954 3870 13022 3926
rect 13078 3870 13200 3926
rect -400 3802 13200 3870
rect -400 3746 -286 3802
rect -230 3746 -162 3802
rect -106 3746 -38 3802
rect 18 3746 86 3802
rect 142 3746 210 3802
rect 266 3790 12526 3802
rect 266 3746 741 3790
rect -400 3734 741 3746
rect 797 3734 883 3790
rect 939 3734 1142 3790
rect 1198 3734 1284 3790
rect 1340 3734 1542 3790
rect 1598 3734 1684 3790
rect 1740 3734 1939 3790
rect 1995 3734 2081 3790
rect 2137 3734 2336 3790
rect 2392 3734 2478 3790
rect 2534 3734 2740 3790
rect 2796 3734 2882 3790
rect 2938 3734 3136 3790
rect 3192 3734 3278 3790
rect 3334 3734 3536 3790
rect 3592 3734 3678 3790
rect 3734 3734 3933 3790
rect 3989 3734 4075 3790
rect 4131 3734 4338 3790
rect 4394 3734 4480 3790
rect 4536 3734 4738 3790
rect 4794 3734 4880 3790
rect 4936 3734 5143 3790
rect 5199 3734 5285 3790
rect 5341 3734 5540 3790
rect 5596 3734 5682 3790
rect 5738 3734 5937 3790
rect 5993 3734 6079 3790
rect 6135 3734 6340 3790
rect 6396 3734 6482 3790
rect 6538 3734 6742 3790
rect 6798 3734 6884 3790
rect 6940 3734 7145 3790
rect 7201 3734 7287 3790
rect 7343 3734 7539 3790
rect 7595 3734 7681 3790
rect 7737 3734 7940 3790
rect 7996 3734 8082 3790
rect 8138 3734 8340 3790
rect 8396 3734 8482 3790
rect 8538 3734 8737 3790
rect 8793 3734 8879 3790
rect 8935 3734 9134 3790
rect 9190 3734 9276 3790
rect 9332 3734 9538 3790
rect 9594 3734 9680 3790
rect 9736 3734 9934 3790
rect 9990 3734 10076 3790
rect 10132 3734 10334 3790
rect 10390 3734 10476 3790
rect 10532 3734 10731 3790
rect 10787 3734 10873 3790
rect 10929 3734 11136 3790
rect 11192 3734 11278 3790
rect 11334 3734 11536 3790
rect 11592 3734 11678 3790
rect 11734 3734 11941 3790
rect 11997 3734 12083 3790
rect 12139 3746 12526 3790
rect 12582 3746 12650 3802
rect 12706 3746 12774 3802
rect 12830 3746 12898 3802
rect 12954 3746 13022 3802
rect 13078 3746 13200 3802
rect 12139 3734 13200 3746
rect -400 3678 13200 3734
rect -400 3622 -286 3678
rect -230 3622 -162 3678
rect -106 3622 -38 3678
rect 18 3622 86 3678
rect 142 3622 210 3678
rect 266 3648 12526 3678
rect 266 3622 741 3648
rect -400 3592 741 3622
rect 797 3592 883 3648
rect 939 3592 1142 3648
rect 1198 3592 1284 3648
rect 1340 3592 1542 3648
rect 1598 3592 1684 3648
rect 1740 3592 1939 3648
rect 1995 3592 2081 3648
rect 2137 3592 2336 3648
rect 2392 3592 2478 3648
rect 2534 3592 2740 3648
rect 2796 3592 2882 3648
rect 2938 3592 3136 3648
rect 3192 3592 3278 3648
rect 3334 3592 3536 3648
rect 3592 3592 3678 3648
rect 3734 3592 3933 3648
rect 3989 3592 4075 3648
rect 4131 3592 4338 3648
rect 4394 3592 4480 3648
rect 4536 3592 4738 3648
rect 4794 3592 4880 3648
rect 4936 3592 5143 3648
rect 5199 3592 5285 3648
rect 5341 3592 5540 3648
rect 5596 3592 5682 3648
rect 5738 3592 5937 3648
rect 5993 3592 6079 3648
rect 6135 3592 6340 3648
rect 6396 3592 6482 3648
rect 6538 3592 6742 3648
rect 6798 3592 6884 3648
rect 6940 3592 7145 3648
rect 7201 3592 7287 3648
rect 7343 3592 7539 3648
rect 7595 3592 7681 3648
rect 7737 3592 7940 3648
rect 7996 3592 8082 3648
rect 8138 3592 8340 3648
rect 8396 3592 8482 3648
rect 8538 3592 8737 3648
rect 8793 3592 8879 3648
rect 8935 3592 9134 3648
rect 9190 3592 9276 3648
rect 9332 3592 9538 3648
rect 9594 3592 9680 3648
rect 9736 3592 9934 3648
rect 9990 3592 10076 3648
rect 10132 3592 10334 3648
rect 10390 3592 10476 3648
rect 10532 3592 10731 3648
rect 10787 3592 10873 3648
rect 10929 3592 11136 3648
rect 11192 3592 11278 3648
rect 11334 3592 11536 3648
rect 11592 3592 11678 3648
rect 11734 3592 11941 3648
rect 11997 3592 12083 3648
rect 12139 3622 12526 3648
rect 12582 3622 12650 3678
rect 12706 3622 12774 3678
rect 12830 3622 12898 3678
rect 12954 3622 13022 3678
rect 13078 3622 13200 3678
rect 12139 3592 13200 3622
rect -400 3554 13200 3592
rect -400 3498 -286 3554
rect -230 3498 -162 3554
rect -106 3498 -38 3554
rect 18 3498 86 3554
rect 142 3498 210 3554
rect 266 3506 12526 3554
rect 266 3498 741 3506
rect -400 3450 741 3498
rect 797 3450 883 3506
rect 939 3450 1142 3506
rect 1198 3450 1284 3506
rect 1340 3450 1542 3506
rect 1598 3450 1684 3506
rect 1740 3450 1939 3506
rect 1995 3450 2081 3506
rect 2137 3450 2336 3506
rect 2392 3450 2478 3506
rect 2534 3450 2740 3506
rect 2796 3450 2882 3506
rect 2938 3450 3136 3506
rect 3192 3450 3278 3506
rect 3334 3450 3536 3506
rect 3592 3450 3678 3506
rect 3734 3450 3933 3506
rect 3989 3450 4075 3506
rect 4131 3450 4338 3506
rect 4394 3450 4480 3506
rect 4536 3450 4738 3506
rect 4794 3450 4880 3506
rect 4936 3450 5143 3506
rect 5199 3450 5285 3506
rect 5341 3450 5540 3506
rect 5596 3450 5682 3506
rect 5738 3450 5937 3506
rect 5993 3450 6079 3506
rect 6135 3450 6340 3506
rect 6396 3450 6482 3506
rect 6538 3450 6742 3506
rect 6798 3450 6884 3506
rect 6940 3450 7145 3506
rect 7201 3450 7287 3506
rect 7343 3450 7539 3506
rect 7595 3450 7681 3506
rect 7737 3450 7940 3506
rect 7996 3450 8082 3506
rect 8138 3450 8340 3506
rect 8396 3450 8482 3506
rect 8538 3450 8737 3506
rect 8793 3450 8879 3506
rect 8935 3450 9134 3506
rect 9190 3450 9276 3506
rect 9332 3450 9538 3506
rect 9594 3450 9680 3506
rect 9736 3450 9934 3506
rect 9990 3450 10076 3506
rect 10132 3450 10334 3506
rect 10390 3450 10476 3506
rect 10532 3450 10731 3506
rect 10787 3450 10873 3506
rect 10929 3450 11136 3506
rect 11192 3450 11278 3506
rect 11334 3450 11536 3506
rect 11592 3450 11678 3506
rect 11734 3450 11941 3506
rect 11997 3450 12083 3506
rect 12139 3498 12526 3506
rect 12582 3498 12650 3554
rect 12706 3498 12774 3554
rect 12830 3498 12898 3554
rect 12954 3498 13022 3554
rect 13078 3498 13200 3554
rect 12139 3450 13200 3498
rect -400 3430 13200 3450
rect -400 3374 -286 3430
rect -230 3374 -162 3430
rect -106 3374 -38 3430
rect 18 3374 86 3430
rect 142 3374 210 3430
rect 266 3374 12526 3430
rect 12582 3374 12650 3430
rect 12706 3374 12774 3430
rect 12830 3374 12898 3430
rect 12954 3374 13022 3430
rect 13078 3374 13200 3430
rect -400 3364 13200 3374
rect -400 3308 741 3364
rect 797 3308 883 3364
rect 939 3308 1142 3364
rect 1198 3308 1284 3364
rect 1340 3308 1542 3364
rect 1598 3308 1684 3364
rect 1740 3308 1939 3364
rect 1995 3308 2081 3364
rect 2137 3308 2336 3364
rect 2392 3308 2478 3364
rect 2534 3308 2740 3364
rect 2796 3308 2882 3364
rect 2938 3308 3136 3364
rect 3192 3308 3278 3364
rect 3334 3308 3536 3364
rect 3592 3308 3678 3364
rect 3734 3308 3933 3364
rect 3989 3308 4075 3364
rect 4131 3308 4338 3364
rect 4394 3308 4480 3364
rect 4536 3308 4738 3364
rect 4794 3308 4880 3364
rect 4936 3308 5143 3364
rect 5199 3308 5285 3364
rect 5341 3308 5540 3364
rect 5596 3308 5682 3364
rect 5738 3308 5937 3364
rect 5993 3308 6079 3364
rect 6135 3308 6340 3364
rect 6396 3308 6482 3364
rect 6538 3308 6742 3364
rect 6798 3308 6884 3364
rect 6940 3308 7145 3364
rect 7201 3308 7287 3364
rect 7343 3308 7539 3364
rect 7595 3308 7681 3364
rect 7737 3308 7940 3364
rect 7996 3308 8082 3364
rect 8138 3308 8340 3364
rect 8396 3308 8482 3364
rect 8538 3308 8737 3364
rect 8793 3308 8879 3364
rect 8935 3308 9134 3364
rect 9190 3308 9276 3364
rect 9332 3308 9538 3364
rect 9594 3308 9680 3364
rect 9736 3308 9934 3364
rect 9990 3308 10076 3364
rect 10132 3308 10334 3364
rect 10390 3308 10476 3364
rect 10532 3308 10731 3364
rect 10787 3308 10873 3364
rect 10929 3308 11136 3364
rect 11192 3308 11278 3364
rect 11334 3308 11536 3364
rect 11592 3308 11678 3364
rect 11734 3308 11941 3364
rect 11997 3308 12083 3364
rect 12139 3308 13200 3364
rect -400 3306 13200 3308
rect -400 3250 -286 3306
rect -230 3250 -162 3306
rect -106 3250 -38 3306
rect 18 3250 86 3306
rect 142 3250 210 3306
rect 266 3250 12526 3306
rect 12582 3250 12650 3306
rect 12706 3250 12774 3306
rect 12830 3250 12898 3306
rect 12954 3250 13022 3306
rect 13078 3250 13200 3306
rect -400 3222 13200 3250
rect -400 3182 741 3222
rect -400 3126 -286 3182
rect -230 3126 -162 3182
rect -106 3126 -38 3182
rect 18 3126 86 3182
rect 142 3126 210 3182
rect 266 3166 741 3182
rect 797 3166 883 3222
rect 939 3166 1142 3222
rect 1198 3166 1284 3222
rect 1340 3166 1542 3222
rect 1598 3166 1684 3222
rect 1740 3166 1939 3222
rect 1995 3166 2081 3222
rect 2137 3166 2336 3222
rect 2392 3166 2478 3222
rect 2534 3166 2740 3222
rect 2796 3166 2882 3222
rect 2938 3166 3136 3222
rect 3192 3166 3278 3222
rect 3334 3166 3536 3222
rect 3592 3166 3678 3222
rect 3734 3166 3933 3222
rect 3989 3166 4075 3222
rect 4131 3166 4338 3222
rect 4394 3166 4480 3222
rect 4536 3166 4738 3222
rect 4794 3166 4880 3222
rect 4936 3166 5143 3222
rect 5199 3166 5285 3222
rect 5341 3166 5540 3222
rect 5596 3166 5682 3222
rect 5738 3166 5937 3222
rect 5993 3166 6079 3222
rect 6135 3166 6340 3222
rect 6396 3166 6482 3222
rect 6538 3166 6742 3222
rect 6798 3166 6884 3222
rect 6940 3166 7145 3222
rect 7201 3166 7287 3222
rect 7343 3166 7539 3222
rect 7595 3166 7681 3222
rect 7737 3166 7940 3222
rect 7996 3166 8082 3222
rect 8138 3166 8340 3222
rect 8396 3166 8482 3222
rect 8538 3166 8737 3222
rect 8793 3166 8879 3222
rect 8935 3166 9134 3222
rect 9190 3166 9276 3222
rect 9332 3166 9538 3222
rect 9594 3166 9680 3222
rect 9736 3166 9934 3222
rect 9990 3166 10076 3222
rect 10132 3166 10334 3222
rect 10390 3166 10476 3222
rect 10532 3166 10731 3222
rect 10787 3166 10873 3222
rect 10929 3166 11136 3222
rect 11192 3166 11278 3222
rect 11334 3166 11536 3222
rect 11592 3166 11678 3222
rect 11734 3166 11941 3222
rect 11997 3166 12083 3222
rect 12139 3182 13200 3222
rect 12139 3166 12526 3182
rect 266 3126 12526 3166
rect 12582 3126 12650 3182
rect 12706 3126 12774 3182
rect 12830 3126 12898 3182
rect 12954 3126 13022 3182
rect 13078 3126 13200 3182
rect -400 3080 13200 3126
rect -400 3058 741 3080
rect -400 3002 -286 3058
rect -230 3002 -162 3058
rect -106 3002 -38 3058
rect 18 3002 86 3058
rect 142 3002 210 3058
rect 266 3024 741 3058
rect 797 3024 883 3080
rect 939 3024 1142 3080
rect 1198 3024 1284 3080
rect 1340 3024 1542 3080
rect 1598 3024 1684 3080
rect 1740 3024 1939 3080
rect 1995 3024 2081 3080
rect 2137 3024 2336 3080
rect 2392 3024 2478 3080
rect 2534 3024 2740 3080
rect 2796 3024 2882 3080
rect 2938 3024 3136 3080
rect 3192 3024 3278 3080
rect 3334 3024 3536 3080
rect 3592 3024 3678 3080
rect 3734 3024 3933 3080
rect 3989 3024 4075 3080
rect 4131 3024 4338 3080
rect 4394 3024 4480 3080
rect 4536 3024 4738 3080
rect 4794 3024 4880 3080
rect 4936 3024 5143 3080
rect 5199 3024 5285 3080
rect 5341 3024 5540 3080
rect 5596 3024 5682 3080
rect 5738 3024 5937 3080
rect 5993 3024 6079 3080
rect 6135 3024 6340 3080
rect 6396 3024 6482 3080
rect 6538 3024 6742 3080
rect 6798 3024 6884 3080
rect 6940 3024 7145 3080
rect 7201 3024 7287 3080
rect 7343 3024 7539 3080
rect 7595 3024 7681 3080
rect 7737 3024 7940 3080
rect 7996 3024 8082 3080
rect 8138 3024 8340 3080
rect 8396 3024 8482 3080
rect 8538 3024 8737 3080
rect 8793 3024 8879 3080
rect 8935 3024 9134 3080
rect 9190 3024 9276 3080
rect 9332 3024 9538 3080
rect 9594 3024 9680 3080
rect 9736 3024 9934 3080
rect 9990 3024 10076 3080
rect 10132 3024 10334 3080
rect 10390 3024 10476 3080
rect 10532 3024 10731 3080
rect 10787 3024 10873 3080
rect 10929 3024 11136 3080
rect 11192 3024 11278 3080
rect 11334 3024 11536 3080
rect 11592 3024 11678 3080
rect 11734 3024 11941 3080
rect 11997 3024 12083 3080
rect 12139 3058 13200 3080
rect 12139 3024 12526 3058
rect 266 3002 12526 3024
rect 12582 3002 12650 3058
rect 12706 3002 12774 3058
rect 12830 3002 12898 3058
rect 12954 3002 13022 3058
rect 13078 3002 13200 3058
rect -400 2938 13200 3002
rect -400 2934 741 2938
rect -400 2878 -286 2934
rect -230 2878 -162 2934
rect -106 2878 -38 2934
rect 18 2878 86 2934
rect 142 2878 210 2934
rect 266 2882 741 2934
rect 797 2882 883 2938
rect 939 2882 1142 2938
rect 1198 2882 1284 2938
rect 1340 2882 1542 2938
rect 1598 2882 1684 2938
rect 1740 2882 1939 2938
rect 1995 2882 2081 2938
rect 2137 2882 2336 2938
rect 2392 2882 2478 2938
rect 2534 2882 2740 2938
rect 2796 2882 2882 2938
rect 2938 2882 3136 2938
rect 3192 2882 3278 2938
rect 3334 2882 3536 2938
rect 3592 2882 3678 2938
rect 3734 2882 3933 2938
rect 3989 2882 4075 2938
rect 4131 2882 4338 2938
rect 4394 2882 4480 2938
rect 4536 2882 4738 2938
rect 4794 2882 4880 2938
rect 4936 2882 5143 2938
rect 5199 2882 5285 2938
rect 5341 2882 5540 2938
rect 5596 2882 5682 2938
rect 5738 2882 5937 2938
rect 5993 2882 6079 2938
rect 6135 2882 6340 2938
rect 6396 2882 6482 2938
rect 6538 2882 6742 2938
rect 6798 2882 6884 2938
rect 6940 2882 7145 2938
rect 7201 2882 7287 2938
rect 7343 2882 7539 2938
rect 7595 2882 7681 2938
rect 7737 2882 7940 2938
rect 7996 2882 8082 2938
rect 8138 2882 8340 2938
rect 8396 2882 8482 2938
rect 8538 2882 8737 2938
rect 8793 2882 8879 2938
rect 8935 2882 9134 2938
rect 9190 2882 9276 2938
rect 9332 2882 9538 2938
rect 9594 2882 9680 2938
rect 9736 2882 9934 2938
rect 9990 2882 10076 2938
rect 10132 2882 10334 2938
rect 10390 2882 10476 2938
rect 10532 2882 10731 2938
rect 10787 2882 10873 2938
rect 10929 2882 11136 2938
rect 11192 2882 11278 2938
rect 11334 2882 11536 2938
rect 11592 2882 11678 2938
rect 11734 2882 11941 2938
rect 11997 2882 12083 2938
rect 12139 2934 13200 2938
rect 12139 2882 12526 2934
rect 266 2878 12526 2882
rect 12582 2878 12650 2934
rect 12706 2878 12774 2934
rect 12830 2878 12898 2934
rect 12954 2878 13022 2934
rect 13078 2878 13200 2934
rect -400 2810 13200 2878
rect -400 2754 -286 2810
rect -230 2754 -162 2810
rect -106 2754 -38 2810
rect 18 2754 86 2810
rect 142 2754 210 2810
rect 266 2796 12526 2810
rect 266 2754 741 2796
rect -400 2740 741 2754
rect 797 2740 883 2796
rect 939 2740 1142 2796
rect 1198 2740 1284 2796
rect 1340 2740 1542 2796
rect 1598 2740 1684 2796
rect 1740 2740 1939 2796
rect 1995 2740 2081 2796
rect 2137 2740 2336 2796
rect 2392 2740 2478 2796
rect 2534 2740 2740 2796
rect 2796 2740 2882 2796
rect 2938 2740 3136 2796
rect 3192 2740 3278 2796
rect 3334 2740 3536 2796
rect 3592 2740 3678 2796
rect 3734 2740 3933 2796
rect 3989 2740 4075 2796
rect 4131 2740 4338 2796
rect 4394 2740 4480 2796
rect 4536 2740 4738 2796
rect 4794 2740 4880 2796
rect 4936 2740 5143 2796
rect 5199 2740 5285 2796
rect 5341 2740 5540 2796
rect 5596 2740 5682 2796
rect 5738 2740 5937 2796
rect 5993 2740 6079 2796
rect 6135 2740 6340 2796
rect 6396 2740 6482 2796
rect 6538 2740 6742 2796
rect 6798 2740 6884 2796
rect 6940 2740 7145 2796
rect 7201 2740 7287 2796
rect 7343 2740 7539 2796
rect 7595 2740 7681 2796
rect 7737 2740 7940 2796
rect 7996 2740 8082 2796
rect 8138 2740 8340 2796
rect 8396 2740 8482 2796
rect 8538 2740 8737 2796
rect 8793 2740 8879 2796
rect 8935 2740 9134 2796
rect 9190 2740 9276 2796
rect 9332 2740 9538 2796
rect 9594 2740 9680 2796
rect 9736 2740 9934 2796
rect 9990 2740 10076 2796
rect 10132 2740 10334 2796
rect 10390 2740 10476 2796
rect 10532 2740 10731 2796
rect 10787 2740 10873 2796
rect 10929 2740 11136 2796
rect 11192 2740 11278 2796
rect 11334 2740 11536 2796
rect 11592 2740 11678 2796
rect 11734 2740 11941 2796
rect 11997 2740 12083 2796
rect 12139 2754 12526 2796
rect 12582 2754 12650 2810
rect 12706 2754 12774 2810
rect 12830 2754 12898 2810
rect 12954 2754 13022 2810
rect 13078 2754 13200 2810
rect 12139 2740 13200 2754
rect -400 2686 13200 2740
rect -400 2630 -286 2686
rect -230 2630 -162 2686
rect -106 2630 -38 2686
rect 18 2630 86 2686
rect 142 2630 210 2686
rect 266 2654 12526 2686
rect 266 2630 741 2654
rect -400 2598 741 2630
rect 797 2598 883 2654
rect 939 2598 1142 2654
rect 1198 2598 1284 2654
rect 1340 2598 1542 2654
rect 1598 2598 1684 2654
rect 1740 2598 1939 2654
rect 1995 2598 2081 2654
rect 2137 2598 2336 2654
rect 2392 2598 2478 2654
rect 2534 2598 2740 2654
rect 2796 2598 2882 2654
rect 2938 2598 3136 2654
rect 3192 2598 3278 2654
rect 3334 2598 3536 2654
rect 3592 2598 3678 2654
rect 3734 2598 3933 2654
rect 3989 2598 4075 2654
rect 4131 2598 4338 2654
rect 4394 2598 4480 2654
rect 4536 2598 4738 2654
rect 4794 2598 4880 2654
rect 4936 2598 5143 2654
rect 5199 2598 5285 2654
rect 5341 2598 5540 2654
rect 5596 2598 5682 2654
rect 5738 2598 5937 2654
rect 5993 2598 6079 2654
rect 6135 2598 6340 2654
rect 6396 2598 6482 2654
rect 6538 2598 6742 2654
rect 6798 2598 6884 2654
rect 6940 2598 7145 2654
rect 7201 2598 7287 2654
rect 7343 2598 7539 2654
rect 7595 2598 7681 2654
rect 7737 2598 7940 2654
rect 7996 2598 8082 2654
rect 8138 2598 8340 2654
rect 8396 2598 8482 2654
rect 8538 2598 8737 2654
rect 8793 2598 8879 2654
rect 8935 2598 9134 2654
rect 9190 2598 9276 2654
rect 9332 2598 9538 2654
rect 9594 2598 9680 2654
rect 9736 2598 9934 2654
rect 9990 2598 10076 2654
rect 10132 2598 10334 2654
rect 10390 2598 10476 2654
rect 10532 2598 10731 2654
rect 10787 2598 10873 2654
rect 10929 2598 11136 2654
rect 11192 2598 11278 2654
rect 11334 2598 11536 2654
rect 11592 2598 11678 2654
rect 11734 2598 11941 2654
rect 11997 2598 12083 2654
rect 12139 2630 12526 2654
rect 12582 2630 12650 2686
rect 12706 2630 12774 2686
rect 12830 2630 12898 2686
rect 12954 2630 13022 2686
rect 13078 2630 13200 2686
rect 12139 2598 13200 2630
rect -400 2562 13200 2598
rect -400 2506 -286 2562
rect -230 2506 -162 2562
rect -106 2506 -38 2562
rect 18 2506 86 2562
rect 142 2506 210 2562
rect 266 2512 12526 2562
rect 266 2506 741 2512
rect -400 2456 741 2506
rect 797 2456 883 2512
rect 939 2456 1142 2512
rect 1198 2456 1284 2512
rect 1340 2456 1542 2512
rect 1598 2456 1684 2512
rect 1740 2456 1939 2512
rect 1995 2456 2081 2512
rect 2137 2456 2336 2512
rect 2392 2456 2478 2512
rect 2534 2456 2740 2512
rect 2796 2456 2882 2512
rect 2938 2456 3136 2512
rect 3192 2456 3278 2512
rect 3334 2456 3536 2512
rect 3592 2456 3678 2512
rect 3734 2456 3933 2512
rect 3989 2456 4075 2512
rect 4131 2456 4338 2512
rect 4394 2456 4480 2512
rect 4536 2456 4738 2512
rect 4794 2456 4880 2512
rect 4936 2456 5143 2512
rect 5199 2456 5285 2512
rect 5341 2456 5540 2512
rect 5596 2456 5682 2512
rect 5738 2456 5937 2512
rect 5993 2456 6079 2512
rect 6135 2456 6340 2512
rect 6396 2456 6482 2512
rect 6538 2456 6742 2512
rect 6798 2456 6884 2512
rect 6940 2456 7145 2512
rect 7201 2456 7287 2512
rect 7343 2456 7539 2512
rect 7595 2456 7681 2512
rect 7737 2456 7940 2512
rect 7996 2456 8082 2512
rect 8138 2456 8340 2512
rect 8396 2456 8482 2512
rect 8538 2456 8737 2512
rect 8793 2456 8879 2512
rect 8935 2456 9134 2512
rect 9190 2456 9276 2512
rect 9332 2456 9538 2512
rect 9594 2456 9680 2512
rect 9736 2456 9934 2512
rect 9990 2456 10076 2512
rect 10132 2456 10334 2512
rect 10390 2456 10476 2512
rect 10532 2456 10731 2512
rect 10787 2456 10873 2512
rect 10929 2456 11136 2512
rect 11192 2456 11278 2512
rect 11334 2456 11536 2512
rect 11592 2456 11678 2512
rect 11734 2456 11941 2512
rect 11997 2456 12083 2512
rect 12139 2506 12526 2512
rect 12582 2506 12650 2562
rect 12706 2506 12774 2562
rect 12830 2506 12898 2562
rect 12954 2506 13022 2562
rect 13078 2506 13200 2562
rect 12139 2456 13200 2506
rect -400 2438 13200 2456
rect -400 2382 -286 2438
rect -230 2382 -162 2438
rect -106 2382 -38 2438
rect 18 2382 86 2438
rect 142 2382 210 2438
rect 266 2382 12526 2438
rect 12582 2382 12650 2438
rect 12706 2382 12774 2438
rect 12830 2382 12898 2438
rect 12954 2382 13022 2438
rect 13078 2382 13200 2438
rect -400 2370 13200 2382
rect -400 2314 741 2370
rect 797 2314 883 2370
rect 939 2314 1142 2370
rect 1198 2314 1284 2370
rect 1340 2314 1542 2370
rect 1598 2314 1684 2370
rect 1740 2314 1939 2370
rect 1995 2314 2081 2370
rect 2137 2314 2336 2370
rect 2392 2314 2478 2370
rect 2534 2314 2740 2370
rect 2796 2314 2882 2370
rect 2938 2314 3136 2370
rect 3192 2314 3278 2370
rect 3334 2314 3536 2370
rect 3592 2314 3678 2370
rect 3734 2314 3933 2370
rect 3989 2314 4075 2370
rect 4131 2314 4338 2370
rect 4394 2314 4480 2370
rect 4536 2314 4738 2370
rect 4794 2314 4880 2370
rect 4936 2314 5143 2370
rect 5199 2314 5285 2370
rect 5341 2314 5540 2370
rect 5596 2314 5682 2370
rect 5738 2314 5937 2370
rect 5993 2314 6079 2370
rect 6135 2314 6340 2370
rect 6396 2314 6482 2370
rect 6538 2314 6742 2370
rect 6798 2314 6884 2370
rect 6940 2314 7145 2370
rect 7201 2314 7287 2370
rect 7343 2314 7539 2370
rect 7595 2314 7681 2370
rect 7737 2314 7940 2370
rect 7996 2314 8082 2370
rect 8138 2314 8340 2370
rect 8396 2314 8482 2370
rect 8538 2314 8737 2370
rect 8793 2314 8879 2370
rect 8935 2314 9134 2370
rect 9190 2314 9276 2370
rect 9332 2314 9538 2370
rect 9594 2314 9680 2370
rect 9736 2314 9934 2370
rect 9990 2314 10076 2370
rect 10132 2314 10334 2370
rect 10390 2314 10476 2370
rect 10532 2314 10731 2370
rect 10787 2314 10873 2370
rect 10929 2314 11136 2370
rect 11192 2314 11278 2370
rect 11334 2314 11536 2370
rect 11592 2314 11678 2370
rect 11734 2314 11941 2370
rect 11997 2314 12083 2370
rect 12139 2314 13200 2370
rect -400 2258 -286 2314
rect -230 2258 -162 2314
rect -106 2258 -38 2314
rect 18 2258 86 2314
rect 142 2258 210 2314
rect 266 2258 12526 2314
rect 12582 2258 12650 2314
rect 12706 2258 12774 2314
rect 12830 2258 12898 2314
rect 12954 2258 13022 2314
rect 13078 2258 13200 2314
rect -400 2228 13200 2258
rect -400 2190 741 2228
rect -400 2134 -286 2190
rect -230 2134 -162 2190
rect -106 2134 -38 2190
rect 18 2134 86 2190
rect 142 2134 210 2190
rect 266 2172 741 2190
rect 797 2172 883 2228
rect 939 2172 1142 2228
rect 1198 2172 1284 2228
rect 1340 2172 1542 2228
rect 1598 2172 1684 2228
rect 1740 2172 1939 2228
rect 1995 2172 2081 2228
rect 2137 2172 2336 2228
rect 2392 2172 2478 2228
rect 2534 2172 2740 2228
rect 2796 2172 2882 2228
rect 2938 2172 3136 2228
rect 3192 2172 3278 2228
rect 3334 2172 3536 2228
rect 3592 2172 3678 2228
rect 3734 2172 3933 2228
rect 3989 2172 4075 2228
rect 4131 2172 4338 2228
rect 4394 2172 4480 2228
rect 4536 2172 4738 2228
rect 4794 2172 4880 2228
rect 4936 2172 5143 2228
rect 5199 2172 5285 2228
rect 5341 2172 5540 2228
rect 5596 2172 5682 2228
rect 5738 2172 5937 2228
rect 5993 2172 6079 2228
rect 6135 2172 6340 2228
rect 6396 2172 6482 2228
rect 6538 2172 6742 2228
rect 6798 2172 6884 2228
rect 6940 2172 7145 2228
rect 7201 2172 7287 2228
rect 7343 2172 7539 2228
rect 7595 2172 7681 2228
rect 7737 2172 7940 2228
rect 7996 2172 8082 2228
rect 8138 2172 8340 2228
rect 8396 2172 8482 2228
rect 8538 2172 8737 2228
rect 8793 2172 8879 2228
rect 8935 2172 9134 2228
rect 9190 2172 9276 2228
rect 9332 2172 9538 2228
rect 9594 2172 9680 2228
rect 9736 2172 9934 2228
rect 9990 2172 10076 2228
rect 10132 2172 10334 2228
rect 10390 2172 10476 2228
rect 10532 2172 10731 2228
rect 10787 2172 10873 2228
rect 10929 2172 11136 2228
rect 11192 2172 11278 2228
rect 11334 2172 11536 2228
rect 11592 2172 11678 2228
rect 11734 2172 11941 2228
rect 11997 2172 12083 2228
rect 12139 2190 13200 2228
rect 12139 2172 12526 2190
rect 266 2134 12526 2172
rect 12582 2134 12650 2190
rect 12706 2134 12774 2190
rect 12830 2134 12898 2190
rect 12954 2134 13022 2190
rect 13078 2134 13200 2190
rect -400 2086 13200 2134
rect -400 2066 741 2086
rect -400 2010 -286 2066
rect -230 2010 -162 2066
rect -106 2010 -38 2066
rect 18 2010 86 2066
rect 142 2010 210 2066
rect 266 2030 741 2066
rect 797 2030 883 2086
rect 939 2030 1142 2086
rect 1198 2030 1284 2086
rect 1340 2030 1542 2086
rect 1598 2030 1684 2086
rect 1740 2030 1939 2086
rect 1995 2030 2081 2086
rect 2137 2030 2336 2086
rect 2392 2030 2478 2086
rect 2534 2030 2740 2086
rect 2796 2030 2882 2086
rect 2938 2030 3136 2086
rect 3192 2030 3278 2086
rect 3334 2030 3536 2086
rect 3592 2030 3678 2086
rect 3734 2030 3933 2086
rect 3989 2030 4075 2086
rect 4131 2030 4338 2086
rect 4394 2030 4480 2086
rect 4536 2030 4738 2086
rect 4794 2030 4880 2086
rect 4936 2030 5143 2086
rect 5199 2030 5285 2086
rect 5341 2030 5540 2086
rect 5596 2030 5682 2086
rect 5738 2030 5937 2086
rect 5993 2030 6079 2086
rect 6135 2030 6340 2086
rect 6396 2030 6482 2086
rect 6538 2030 6742 2086
rect 6798 2030 6884 2086
rect 6940 2030 7145 2086
rect 7201 2030 7287 2086
rect 7343 2030 7539 2086
rect 7595 2030 7681 2086
rect 7737 2030 7940 2086
rect 7996 2030 8082 2086
rect 8138 2030 8340 2086
rect 8396 2030 8482 2086
rect 8538 2030 8737 2086
rect 8793 2030 8879 2086
rect 8935 2030 9134 2086
rect 9190 2030 9276 2086
rect 9332 2030 9538 2086
rect 9594 2030 9680 2086
rect 9736 2030 9934 2086
rect 9990 2030 10076 2086
rect 10132 2030 10334 2086
rect 10390 2030 10476 2086
rect 10532 2030 10731 2086
rect 10787 2030 10873 2086
rect 10929 2030 11136 2086
rect 11192 2030 11278 2086
rect 11334 2030 11536 2086
rect 11592 2030 11678 2086
rect 11734 2030 11941 2086
rect 11997 2030 12083 2086
rect 12139 2066 13200 2086
rect 12139 2030 12526 2066
rect 266 2010 12526 2030
rect 12582 2010 12650 2066
rect 12706 2010 12774 2066
rect 12830 2010 12898 2066
rect 12954 2010 13022 2066
rect 13078 2010 13200 2066
rect -400 1944 13200 2010
rect -400 1942 741 1944
rect -400 1886 -286 1942
rect -230 1886 -162 1942
rect -106 1886 -38 1942
rect 18 1886 86 1942
rect 142 1886 210 1942
rect 266 1888 741 1942
rect 797 1888 883 1944
rect 939 1888 1142 1944
rect 1198 1888 1284 1944
rect 1340 1888 1542 1944
rect 1598 1888 1684 1944
rect 1740 1888 1939 1944
rect 1995 1888 2081 1944
rect 2137 1888 2336 1944
rect 2392 1888 2478 1944
rect 2534 1888 2740 1944
rect 2796 1888 2882 1944
rect 2938 1888 3136 1944
rect 3192 1888 3278 1944
rect 3334 1888 3536 1944
rect 3592 1888 3678 1944
rect 3734 1888 3933 1944
rect 3989 1888 4075 1944
rect 4131 1888 4338 1944
rect 4394 1888 4480 1944
rect 4536 1888 4738 1944
rect 4794 1888 4880 1944
rect 4936 1888 5143 1944
rect 5199 1888 5285 1944
rect 5341 1888 5540 1944
rect 5596 1888 5682 1944
rect 5738 1888 5937 1944
rect 5993 1888 6079 1944
rect 6135 1888 6340 1944
rect 6396 1888 6482 1944
rect 6538 1888 6742 1944
rect 6798 1888 6884 1944
rect 6940 1888 7145 1944
rect 7201 1888 7287 1944
rect 7343 1888 7539 1944
rect 7595 1888 7681 1944
rect 7737 1888 7940 1944
rect 7996 1888 8082 1944
rect 8138 1888 8340 1944
rect 8396 1888 8482 1944
rect 8538 1888 8737 1944
rect 8793 1888 8879 1944
rect 8935 1888 9134 1944
rect 9190 1888 9276 1944
rect 9332 1888 9538 1944
rect 9594 1888 9680 1944
rect 9736 1888 9934 1944
rect 9990 1888 10076 1944
rect 10132 1888 10334 1944
rect 10390 1888 10476 1944
rect 10532 1888 10731 1944
rect 10787 1888 10873 1944
rect 10929 1888 11136 1944
rect 11192 1888 11278 1944
rect 11334 1888 11536 1944
rect 11592 1888 11678 1944
rect 11734 1888 11941 1944
rect 11997 1888 12083 1944
rect 12139 1942 13200 1944
rect 12139 1888 12526 1942
rect 266 1886 12526 1888
rect 12582 1886 12650 1942
rect 12706 1886 12774 1942
rect 12830 1886 12898 1942
rect 12954 1886 13022 1942
rect 13078 1886 13200 1942
rect -400 1818 13200 1886
rect -400 1762 -286 1818
rect -230 1762 -162 1818
rect -106 1762 -38 1818
rect 18 1762 86 1818
rect 142 1762 210 1818
rect 266 1802 12526 1818
rect 266 1762 741 1802
rect -400 1746 741 1762
rect 797 1746 883 1802
rect 939 1746 1142 1802
rect 1198 1746 1284 1802
rect 1340 1746 1542 1802
rect 1598 1746 1684 1802
rect 1740 1746 1939 1802
rect 1995 1746 2081 1802
rect 2137 1746 2336 1802
rect 2392 1746 2478 1802
rect 2534 1746 2740 1802
rect 2796 1746 2882 1802
rect 2938 1746 3136 1802
rect 3192 1746 3278 1802
rect 3334 1746 3536 1802
rect 3592 1746 3678 1802
rect 3734 1746 3933 1802
rect 3989 1746 4075 1802
rect 4131 1746 4338 1802
rect 4394 1746 4480 1802
rect 4536 1746 4738 1802
rect 4794 1746 4880 1802
rect 4936 1746 5143 1802
rect 5199 1746 5285 1802
rect 5341 1746 5540 1802
rect 5596 1746 5682 1802
rect 5738 1746 5937 1802
rect 5993 1746 6079 1802
rect 6135 1746 6340 1802
rect 6396 1746 6482 1802
rect 6538 1746 6742 1802
rect 6798 1746 6884 1802
rect 6940 1746 7145 1802
rect 7201 1746 7287 1802
rect 7343 1746 7539 1802
rect 7595 1746 7681 1802
rect 7737 1746 7940 1802
rect 7996 1746 8082 1802
rect 8138 1746 8340 1802
rect 8396 1746 8482 1802
rect 8538 1746 8737 1802
rect 8793 1746 8879 1802
rect 8935 1746 9134 1802
rect 9190 1746 9276 1802
rect 9332 1746 9538 1802
rect 9594 1746 9680 1802
rect 9736 1746 9934 1802
rect 9990 1746 10076 1802
rect 10132 1746 10334 1802
rect 10390 1746 10476 1802
rect 10532 1746 10731 1802
rect 10787 1746 10873 1802
rect 10929 1746 11136 1802
rect 11192 1746 11278 1802
rect 11334 1746 11536 1802
rect 11592 1746 11678 1802
rect 11734 1746 11941 1802
rect 11997 1746 12083 1802
rect 12139 1762 12526 1802
rect 12582 1762 12650 1818
rect 12706 1762 12774 1818
rect 12830 1762 12898 1818
rect 12954 1762 13022 1818
rect 13078 1762 13200 1818
rect 12139 1746 13200 1762
rect -400 1694 13200 1746
rect -400 1638 -286 1694
rect -230 1638 -162 1694
rect -106 1638 -38 1694
rect 18 1638 86 1694
rect 142 1638 210 1694
rect 266 1660 12526 1694
rect 266 1638 741 1660
rect -400 1604 741 1638
rect 797 1604 883 1660
rect 939 1604 1142 1660
rect 1198 1604 1284 1660
rect 1340 1604 1542 1660
rect 1598 1604 1684 1660
rect 1740 1604 1939 1660
rect 1995 1604 2081 1660
rect 2137 1604 2336 1660
rect 2392 1604 2478 1660
rect 2534 1604 2740 1660
rect 2796 1604 2882 1660
rect 2938 1604 3136 1660
rect 3192 1604 3278 1660
rect 3334 1604 3536 1660
rect 3592 1604 3678 1660
rect 3734 1604 3933 1660
rect 3989 1604 4075 1660
rect 4131 1604 4338 1660
rect 4394 1604 4480 1660
rect 4536 1604 4738 1660
rect 4794 1604 4880 1660
rect 4936 1604 5143 1660
rect 5199 1604 5285 1660
rect 5341 1604 5540 1660
rect 5596 1604 5682 1660
rect 5738 1604 5937 1660
rect 5993 1604 6079 1660
rect 6135 1604 6340 1660
rect 6396 1604 6482 1660
rect 6538 1604 6742 1660
rect 6798 1604 6884 1660
rect 6940 1604 7145 1660
rect 7201 1604 7287 1660
rect 7343 1604 7539 1660
rect 7595 1604 7681 1660
rect 7737 1604 7940 1660
rect 7996 1604 8082 1660
rect 8138 1604 8340 1660
rect 8396 1604 8482 1660
rect 8538 1604 8737 1660
rect 8793 1604 8879 1660
rect 8935 1604 9134 1660
rect 9190 1604 9276 1660
rect 9332 1604 9538 1660
rect 9594 1604 9680 1660
rect 9736 1604 9934 1660
rect 9990 1604 10076 1660
rect 10132 1604 10334 1660
rect 10390 1604 10476 1660
rect 10532 1604 10731 1660
rect 10787 1604 10873 1660
rect 10929 1604 11136 1660
rect 11192 1604 11278 1660
rect 11334 1604 11536 1660
rect 11592 1604 11678 1660
rect 11734 1604 11941 1660
rect 11997 1604 12083 1660
rect 12139 1638 12526 1660
rect 12582 1638 12650 1694
rect 12706 1638 12774 1694
rect 12830 1638 12898 1694
rect 12954 1638 13022 1694
rect 13078 1638 13200 1694
rect 12139 1604 13200 1638
rect -400 1570 13200 1604
rect -400 1514 -286 1570
rect -230 1514 -162 1570
rect -106 1514 -38 1570
rect 18 1514 86 1570
rect 142 1514 210 1570
rect 266 1518 12526 1570
rect 266 1514 741 1518
rect -400 1462 741 1514
rect 797 1462 883 1518
rect 939 1462 1142 1518
rect 1198 1462 1284 1518
rect 1340 1462 1542 1518
rect 1598 1462 1684 1518
rect 1740 1462 1939 1518
rect 1995 1462 2081 1518
rect 2137 1462 2336 1518
rect 2392 1462 2478 1518
rect 2534 1462 2740 1518
rect 2796 1462 2882 1518
rect 2938 1462 3136 1518
rect 3192 1462 3278 1518
rect 3334 1462 3536 1518
rect 3592 1462 3678 1518
rect 3734 1462 3933 1518
rect 3989 1462 4075 1518
rect 4131 1462 4338 1518
rect 4394 1462 4480 1518
rect 4536 1462 4738 1518
rect 4794 1462 4880 1518
rect 4936 1462 5143 1518
rect 5199 1462 5285 1518
rect 5341 1462 5540 1518
rect 5596 1462 5682 1518
rect 5738 1462 5937 1518
rect 5993 1462 6079 1518
rect 6135 1462 6340 1518
rect 6396 1462 6482 1518
rect 6538 1462 6742 1518
rect 6798 1462 6884 1518
rect 6940 1462 7145 1518
rect 7201 1462 7287 1518
rect 7343 1462 7539 1518
rect 7595 1462 7681 1518
rect 7737 1462 7940 1518
rect 7996 1462 8082 1518
rect 8138 1462 8340 1518
rect 8396 1462 8482 1518
rect 8538 1462 8737 1518
rect 8793 1462 8879 1518
rect 8935 1462 9134 1518
rect 9190 1462 9276 1518
rect 9332 1462 9538 1518
rect 9594 1462 9680 1518
rect 9736 1462 9934 1518
rect 9990 1462 10076 1518
rect 10132 1462 10334 1518
rect 10390 1462 10476 1518
rect 10532 1462 10731 1518
rect 10787 1462 10873 1518
rect 10929 1462 11136 1518
rect 11192 1462 11278 1518
rect 11334 1462 11536 1518
rect 11592 1462 11678 1518
rect 11734 1462 11941 1518
rect 11997 1462 12083 1518
rect 12139 1514 12526 1518
rect 12582 1514 12650 1570
rect 12706 1514 12774 1570
rect 12830 1514 12898 1570
rect 12954 1514 13022 1570
rect 13078 1514 13200 1570
rect 12139 1462 13200 1514
rect -400 1446 13200 1462
rect -400 1390 -286 1446
rect -230 1390 -162 1446
rect -106 1390 -38 1446
rect 18 1390 86 1446
rect 142 1390 210 1446
rect 266 1390 12526 1446
rect 12582 1390 12650 1446
rect 12706 1390 12774 1446
rect 12830 1390 12898 1446
rect 12954 1390 13022 1446
rect 13078 1390 13200 1446
rect -400 1376 13200 1390
rect -400 1322 741 1376
rect -400 1266 -286 1322
rect -230 1266 -162 1322
rect -106 1266 -38 1322
rect 18 1266 86 1322
rect 142 1266 210 1322
rect 266 1320 741 1322
rect 797 1320 883 1376
rect 939 1320 1142 1376
rect 1198 1320 1284 1376
rect 1340 1320 1542 1376
rect 1598 1320 1684 1376
rect 1740 1320 1939 1376
rect 1995 1320 2081 1376
rect 2137 1320 2336 1376
rect 2392 1320 2478 1376
rect 2534 1320 2740 1376
rect 2796 1320 2882 1376
rect 2938 1320 3136 1376
rect 3192 1320 3278 1376
rect 3334 1320 3536 1376
rect 3592 1320 3678 1376
rect 3734 1320 3933 1376
rect 3989 1320 4075 1376
rect 4131 1320 4338 1376
rect 4394 1320 4480 1376
rect 4536 1320 4738 1376
rect 4794 1320 4880 1376
rect 4936 1320 5143 1376
rect 5199 1320 5285 1376
rect 5341 1320 5540 1376
rect 5596 1320 5682 1376
rect 5738 1320 5937 1376
rect 5993 1320 6079 1376
rect 6135 1320 6340 1376
rect 6396 1320 6482 1376
rect 6538 1320 6742 1376
rect 6798 1320 6884 1376
rect 6940 1320 7145 1376
rect 7201 1320 7287 1376
rect 7343 1320 7539 1376
rect 7595 1320 7681 1376
rect 7737 1320 7940 1376
rect 7996 1320 8082 1376
rect 8138 1320 8340 1376
rect 8396 1320 8482 1376
rect 8538 1320 8737 1376
rect 8793 1320 8879 1376
rect 8935 1320 9134 1376
rect 9190 1320 9276 1376
rect 9332 1320 9538 1376
rect 9594 1320 9680 1376
rect 9736 1320 9934 1376
rect 9990 1320 10076 1376
rect 10132 1320 10334 1376
rect 10390 1320 10476 1376
rect 10532 1320 10731 1376
rect 10787 1320 10873 1376
rect 10929 1320 11136 1376
rect 11192 1320 11278 1376
rect 11334 1320 11536 1376
rect 11592 1320 11678 1376
rect 11734 1320 11941 1376
rect 11997 1320 12083 1376
rect 12139 1322 13200 1376
rect 12139 1320 12526 1322
rect 266 1266 12526 1320
rect 12582 1266 12650 1322
rect 12706 1266 12774 1322
rect 12830 1266 12898 1322
rect 12954 1266 13022 1322
rect 13078 1266 13200 1322
rect -400 1234 13200 1266
rect -400 1198 741 1234
rect -400 1142 -286 1198
rect -230 1142 -162 1198
rect -106 1142 -38 1198
rect 18 1142 86 1198
rect 142 1142 210 1198
rect 266 1178 741 1198
rect 797 1178 883 1234
rect 939 1178 1142 1234
rect 1198 1178 1284 1234
rect 1340 1178 1542 1234
rect 1598 1178 1684 1234
rect 1740 1178 1939 1234
rect 1995 1178 2081 1234
rect 2137 1178 2336 1234
rect 2392 1178 2478 1234
rect 2534 1178 2740 1234
rect 2796 1178 2882 1234
rect 2938 1178 3136 1234
rect 3192 1178 3278 1234
rect 3334 1178 3536 1234
rect 3592 1178 3678 1234
rect 3734 1178 3933 1234
rect 3989 1178 4075 1234
rect 4131 1178 4338 1234
rect 4394 1178 4480 1234
rect 4536 1178 4738 1234
rect 4794 1178 4880 1234
rect 4936 1178 5143 1234
rect 5199 1178 5285 1234
rect 5341 1178 5540 1234
rect 5596 1178 5682 1234
rect 5738 1178 5937 1234
rect 5993 1178 6079 1234
rect 6135 1178 6340 1234
rect 6396 1178 6482 1234
rect 6538 1178 6742 1234
rect 6798 1178 6884 1234
rect 6940 1178 7145 1234
rect 7201 1178 7287 1234
rect 7343 1178 7539 1234
rect 7595 1178 7681 1234
rect 7737 1178 7940 1234
rect 7996 1178 8082 1234
rect 8138 1178 8340 1234
rect 8396 1178 8482 1234
rect 8538 1178 8737 1234
rect 8793 1178 8879 1234
rect 8935 1178 9134 1234
rect 9190 1178 9276 1234
rect 9332 1178 9538 1234
rect 9594 1178 9680 1234
rect 9736 1178 9934 1234
rect 9990 1178 10076 1234
rect 10132 1178 10334 1234
rect 10390 1178 10476 1234
rect 10532 1178 10731 1234
rect 10787 1178 10873 1234
rect 10929 1178 11136 1234
rect 11192 1178 11278 1234
rect 11334 1178 11536 1234
rect 11592 1178 11678 1234
rect 11734 1178 11941 1234
rect 11997 1178 12083 1234
rect 12139 1198 13200 1234
rect 12139 1178 12526 1198
rect 266 1142 12526 1178
rect 12582 1142 12650 1198
rect 12706 1142 12774 1198
rect 12830 1142 12898 1198
rect 12954 1142 13022 1198
rect 13078 1142 13200 1198
rect -400 1092 13200 1142
rect -400 1074 741 1092
rect -400 1018 -286 1074
rect -230 1018 -162 1074
rect -106 1018 -38 1074
rect 18 1018 86 1074
rect 142 1018 210 1074
rect 266 1036 741 1074
rect 797 1036 883 1092
rect 939 1036 1142 1092
rect 1198 1036 1284 1092
rect 1340 1036 1542 1092
rect 1598 1036 1684 1092
rect 1740 1036 1939 1092
rect 1995 1036 2081 1092
rect 2137 1036 2336 1092
rect 2392 1036 2478 1092
rect 2534 1036 2740 1092
rect 2796 1036 2882 1092
rect 2938 1036 3136 1092
rect 3192 1036 3278 1092
rect 3334 1036 3536 1092
rect 3592 1036 3678 1092
rect 3734 1036 3933 1092
rect 3989 1036 4075 1092
rect 4131 1036 4338 1092
rect 4394 1036 4480 1092
rect 4536 1036 4738 1092
rect 4794 1036 4880 1092
rect 4936 1036 5143 1092
rect 5199 1036 5285 1092
rect 5341 1036 5540 1092
rect 5596 1036 5682 1092
rect 5738 1036 5937 1092
rect 5993 1036 6079 1092
rect 6135 1036 6340 1092
rect 6396 1036 6482 1092
rect 6538 1036 6742 1092
rect 6798 1036 6884 1092
rect 6940 1036 7145 1092
rect 7201 1036 7287 1092
rect 7343 1036 7539 1092
rect 7595 1036 7681 1092
rect 7737 1036 7940 1092
rect 7996 1036 8082 1092
rect 8138 1036 8340 1092
rect 8396 1036 8482 1092
rect 8538 1036 8737 1092
rect 8793 1036 8879 1092
rect 8935 1036 9134 1092
rect 9190 1036 9276 1092
rect 9332 1036 9538 1092
rect 9594 1036 9680 1092
rect 9736 1036 9934 1092
rect 9990 1036 10076 1092
rect 10132 1036 10334 1092
rect 10390 1036 10476 1092
rect 10532 1036 10731 1092
rect 10787 1036 10873 1092
rect 10929 1036 11136 1092
rect 11192 1036 11278 1092
rect 11334 1036 11536 1092
rect 11592 1036 11678 1092
rect 11734 1036 11941 1092
rect 11997 1036 12083 1092
rect 12139 1074 13200 1092
rect 12139 1036 12526 1074
rect 266 1018 12526 1036
rect 12582 1018 12650 1074
rect 12706 1018 12774 1074
rect 12830 1018 12898 1074
rect 12954 1018 13022 1074
rect 13078 1018 13200 1074
rect -400 950 13200 1018
rect -400 894 -286 950
rect -230 894 -162 950
rect -106 894 -38 950
rect 18 894 86 950
rect 142 894 210 950
rect 266 894 741 950
rect 797 894 883 950
rect 939 894 1142 950
rect 1198 894 1284 950
rect 1340 894 1542 950
rect 1598 894 1684 950
rect 1740 894 1939 950
rect 1995 894 2081 950
rect 2137 894 2336 950
rect 2392 894 2478 950
rect 2534 894 2740 950
rect 2796 894 2882 950
rect 2938 894 3136 950
rect 3192 894 3278 950
rect 3334 894 3536 950
rect 3592 894 3678 950
rect 3734 894 3933 950
rect 3989 894 4075 950
rect 4131 894 4338 950
rect 4394 894 4480 950
rect 4536 894 4738 950
rect 4794 894 4880 950
rect 4936 894 5143 950
rect 5199 894 5285 950
rect 5341 894 5540 950
rect 5596 894 5682 950
rect 5738 894 5937 950
rect 5993 894 6079 950
rect 6135 894 6340 950
rect 6396 894 6482 950
rect 6538 894 6742 950
rect 6798 894 6884 950
rect 6940 894 7145 950
rect 7201 894 7287 950
rect 7343 894 7539 950
rect 7595 894 7681 950
rect 7737 894 7940 950
rect 7996 894 8082 950
rect 8138 894 8340 950
rect 8396 894 8482 950
rect 8538 894 8737 950
rect 8793 894 8879 950
rect 8935 894 9134 950
rect 9190 894 9276 950
rect 9332 894 9538 950
rect 9594 894 9680 950
rect 9736 894 9934 950
rect 9990 894 10076 950
rect 10132 894 10334 950
rect 10390 894 10476 950
rect 10532 894 10731 950
rect 10787 894 10873 950
rect 10929 894 11136 950
rect 11192 894 11278 950
rect 11334 894 11536 950
rect 11592 894 11678 950
rect 11734 894 11941 950
rect 11997 894 12083 950
rect 12139 894 12526 950
rect 12582 894 12650 950
rect 12706 894 12774 950
rect 12830 894 12898 950
rect 12954 894 13022 950
rect 13078 894 13200 950
rect -400 826 13200 894
rect -400 770 -286 826
rect -230 770 -162 826
rect -106 770 -38 826
rect 18 770 86 826
rect 142 770 210 826
rect 266 808 12526 826
rect 266 770 741 808
rect -400 752 741 770
rect 797 752 883 808
rect 939 752 1142 808
rect 1198 752 1284 808
rect 1340 752 1542 808
rect 1598 752 1684 808
rect 1740 752 1939 808
rect 1995 752 2081 808
rect 2137 752 2336 808
rect 2392 752 2478 808
rect 2534 752 2740 808
rect 2796 752 2882 808
rect 2938 752 3136 808
rect 3192 752 3278 808
rect 3334 752 3536 808
rect 3592 752 3678 808
rect 3734 752 3933 808
rect 3989 752 4075 808
rect 4131 752 4338 808
rect 4394 752 4480 808
rect 4536 752 4738 808
rect 4794 752 4880 808
rect 4936 752 5143 808
rect 5199 752 5285 808
rect 5341 752 5540 808
rect 5596 752 5682 808
rect 5738 752 5937 808
rect 5993 752 6079 808
rect 6135 752 6340 808
rect 6396 752 6482 808
rect 6538 752 6742 808
rect 6798 752 6884 808
rect 6940 752 7145 808
rect 7201 752 7287 808
rect 7343 752 7539 808
rect 7595 752 7681 808
rect 7737 752 7940 808
rect 7996 752 8082 808
rect 8138 752 8340 808
rect 8396 752 8482 808
rect 8538 752 8737 808
rect 8793 752 8879 808
rect 8935 752 9134 808
rect 9190 752 9276 808
rect 9332 752 9538 808
rect 9594 752 9680 808
rect 9736 752 9934 808
rect 9990 752 10076 808
rect 10132 752 10334 808
rect 10390 752 10476 808
rect 10532 752 10731 808
rect 10787 752 10873 808
rect 10929 752 11136 808
rect 11192 752 11278 808
rect 11334 752 11536 808
rect 11592 752 11678 808
rect 11734 752 11941 808
rect 11997 752 12083 808
rect 12139 770 12526 808
rect 12582 770 12650 826
rect 12706 770 12774 826
rect 12830 770 12898 826
rect 12954 770 13022 826
rect 13078 770 13200 826
rect 12139 752 13200 770
rect -400 702 13200 752
rect -400 646 -286 702
rect -230 646 -162 702
rect -106 646 -38 702
rect 18 646 86 702
rect 142 646 210 702
rect 266 666 12526 702
rect 266 646 741 666
rect -400 610 741 646
rect 797 610 883 666
rect 939 610 1142 666
rect 1198 610 1284 666
rect 1340 610 1542 666
rect 1598 610 1684 666
rect 1740 610 1939 666
rect 1995 610 2081 666
rect 2137 610 2336 666
rect 2392 610 2478 666
rect 2534 610 2740 666
rect 2796 610 2882 666
rect 2938 610 3136 666
rect 3192 610 3278 666
rect 3334 610 3536 666
rect 3592 610 3678 666
rect 3734 610 3933 666
rect 3989 610 4075 666
rect 4131 610 4338 666
rect 4394 610 4480 666
rect 4536 610 4738 666
rect 4794 610 4880 666
rect 4936 610 5143 666
rect 5199 610 5285 666
rect 5341 610 5540 666
rect 5596 610 5682 666
rect 5738 610 5937 666
rect 5993 610 6079 666
rect 6135 610 6340 666
rect 6396 610 6482 666
rect 6538 610 6742 666
rect 6798 610 6884 666
rect 6940 610 7145 666
rect 7201 610 7287 666
rect 7343 610 7539 666
rect 7595 610 7681 666
rect 7737 610 7940 666
rect 7996 610 8082 666
rect 8138 610 8340 666
rect 8396 610 8482 666
rect 8538 610 8737 666
rect 8793 610 8879 666
rect 8935 610 9134 666
rect 9190 610 9276 666
rect 9332 610 9538 666
rect 9594 610 9680 666
rect 9736 610 9934 666
rect 9990 610 10076 666
rect 10132 610 10334 666
rect 10390 610 10476 666
rect 10532 610 10731 666
rect 10787 610 10873 666
rect 10929 610 11136 666
rect 11192 610 11278 666
rect 11334 610 11536 666
rect 11592 610 11678 666
rect 11734 610 11941 666
rect 11997 610 12083 666
rect 12139 646 12526 666
rect 12582 646 12650 702
rect 12706 646 12774 702
rect 12830 646 12898 702
rect 12954 646 13022 702
rect 13078 646 13200 702
rect 12139 610 13200 646
rect -400 578 13200 610
rect -400 522 -286 578
rect -230 522 -162 578
rect -106 522 -38 578
rect 18 522 86 578
rect 142 522 210 578
rect 266 524 12526 578
rect 266 522 741 524
rect -400 468 741 522
rect 797 468 883 524
rect 939 468 1142 524
rect 1198 468 1284 524
rect 1340 468 1542 524
rect 1598 468 1684 524
rect 1740 468 1939 524
rect 1995 468 2081 524
rect 2137 468 2336 524
rect 2392 468 2478 524
rect 2534 468 2740 524
rect 2796 468 2882 524
rect 2938 468 3136 524
rect 3192 468 3278 524
rect 3334 468 3536 524
rect 3592 468 3678 524
rect 3734 468 3933 524
rect 3989 468 4075 524
rect 4131 468 4338 524
rect 4394 468 4480 524
rect 4536 468 4738 524
rect 4794 468 4880 524
rect 4936 468 5143 524
rect 5199 468 5285 524
rect 5341 468 5540 524
rect 5596 468 5682 524
rect 5738 468 5937 524
rect 5993 468 6079 524
rect 6135 468 6340 524
rect 6396 468 6482 524
rect 6538 468 6742 524
rect 6798 468 6884 524
rect 6940 468 7145 524
rect 7201 468 7287 524
rect 7343 468 7539 524
rect 7595 468 7681 524
rect 7737 468 7940 524
rect 7996 468 8082 524
rect 8138 468 8340 524
rect 8396 468 8482 524
rect 8538 468 8737 524
rect 8793 468 8879 524
rect 8935 468 9134 524
rect 9190 468 9276 524
rect 9332 468 9538 524
rect 9594 468 9680 524
rect 9736 468 9934 524
rect 9990 468 10076 524
rect 10132 468 10334 524
rect 10390 468 10476 524
rect 10532 468 10731 524
rect 10787 468 10873 524
rect 10929 468 11136 524
rect 11192 468 11278 524
rect 11334 468 11536 524
rect 11592 468 11678 524
rect 11734 468 11941 524
rect 11997 468 12083 524
rect 12139 522 12526 524
rect 12582 522 12650 578
rect 12706 522 12774 578
rect 12830 522 12898 578
rect 12954 522 13022 578
rect 13078 522 13200 578
rect 12139 468 13200 522
rect -400 454 13200 468
rect -400 398 -286 454
rect -230 398 -162 454
rect -106 398 -38 454
rect 18 398 86 454
rect 142 398 210 454
rect 266 398 12526 454
rect 12582 398 12650 454
rect 12706 398 12774 454
rect 12830 398 12898 454
rect 12954 398 13022 454
rect 13078 398 13200 454
rect -400 330 13200 398
rect -400 274 -286 330
rect -230 274 -162 330
rect -106 274 -38 330
rect 18 274 86 330
rect 142 274 210 330
rect 266 302 12526 330
rect 266 274 415 302
rect -400 246 415 274
rect 471 246 557 302
rect 613 246 699 302
rect 755 246 841 302
rect 897 246 983 302
rect 1039 246 1125 302
rect 1181 246 1267 302
rect 1323 246 1409 302
rect 1465 246 1551 302
rect 1607 246 1693 302
rect 1749 246 1835 302
rect 1891 246 1977 302
rect 2033 246 2119 302
rect 2175 246 2261 302
rect 2317 246 2403 302
rect 2459 246 2545 302
rect 2601 246 2687 302
rect 2743 246 2829 302
rect 2885 246 2971 302
rect 3027 246 3113 302
rect 3169 246 3255 302
rect 3311 246 3397 302
rect 3453 246 3539 302
rect 3595 246 3681 302
rect 3737 246 3823 302
rect 3879 246 3965 302
rect 4021 246 4107 302
rect 4163 246 4249 302
rect 4305 246 4391 302
rect 4447 246 4533 302
rect 4589 246 4675 302
rect 4731 246 4817 302
rect 4873 246 4959 302
rect 5015 246 5101 302
rect 5157 246 5243 302
rect 5299 246 5385 302
rect 5441 246 5527 302
rect 5583 246 5669 302
rect 5725 246 5811 302
rect 5867 246 5953 302
rect 6009 246 6095 302
rect 6151 246 6237 302
rect 6293 246 6379 302
rect 6435 246 6521 302
rect 6577 246 6663 302
rect 6719 246 6805 302
rect 6861 246 6947 302
rect 7003 246 7089 302
rect 7145 246 7231 302
rect 7287 246 7373 302
rect 7429 246 7515 302
rect 7571 246 7657 302
rect 7713 246 7799 302
rect 7855 246 7941 302
rect 7997 246 8083 302
rect 8139 246 8225 302
rect 8281 246 8367 302
rect 8423 246 8509 302
rect 8565 246 8651 302
rect 8707 246 8793 302
rect 8849 246 8935 302
rect 8991 246 9077 302
rect 9133 246 9219 302
rect 9275 246 9361 302
rect 9417 246 9503 302
rect 9559 246 9645 302
rect 9701 246 9787 302
rect 9843 246 9929 302
rect 9985 246 10071 302
rect 10127 246 10213 302
rect 10269 246 10355 302
rect 10411 246 10497 302
rect 10553 246 10639 302
rect 10695 246 10781 302
rect 10837 246 10923 302
rect 10979 246 11065 302
rect 11121 246 11207 302
rect 11263 246 11349 302
rect 11405 246 11491 302
rect 11547 246 11633 302
rect 11689 246 11775 302
rect 11831 246 11917 302
rect 11973 246 12059 302
rect 12115 246 12201 302
rect 12257 246 12343 302
rect 12399 274 12526 302
rect 12582 274 12650 330
rect 12706 274 12774 330
rect 12830 274 12898 330
rect 12954 274 13022 330
rect 13078 274 13200 330
rect 12399 246 13200 274
rect -400 206 13200 246
rect -400 150 -286 206
rect -230 150 -162 206
rect -106 150 -38 206
rect 18 150 86 206
rect 142 150 210 206
rect 266 160 12526 206
rect 266 150 415 160
rect -400 104 415 150
rect 471 104 557 160
rect 613 104 699 160
rect 755 104 841 160
rect 897 104 983 160
rect 1039 104 1125 160
rect 1181 104 1267 160
rect 1323 104 1409 160
rect 1465 104 1551 160
rect 1607 104 1693 160
rect 1749 104 1835 160
rect 1891 104 1977 160
rect 2033 104 2119 160
rect 2175 104 2261 160
rect 2317 104 2403 160
rect 2459 104 2545 160
rect 2601 104 2687 160
rect 2743 104 2829 160
rect 2885 104 2971 160
rect 3027 104 3113 160
rect 3169 104 3255 160
rect 3311 104 3397 160
rect 3453 104 3539 160
rect 3595 104 3681 160
rect 3737 104 3823 160
rect 3879 104 3965 160
rect 4021 104 4107 160
rect 4163 104 4249 160
rect 4305 104 4391 160
rect 4447 104 4533 160
rect 4589 104 4675 160
rect 4731 104 4817 160
rect 4873 104 4959 160
rect 5015 104 5101 160
rect 5157 104 5243 160
rect 5299 104 5385 160
rect 5441 104 5527 160
rect 5583 104 5669 160
rect 5725 104 5811 160
rect 5867 104 5953 160
rect 6009 104 6095 160
rect 6151 104 6237 160
rect 6293 104 6379 160
rect 6435 104 6521 160
rect 6577 104 6663 160
rect 6719 104 6805 160
rect 6861 104 6947 160
rect 7003 104 7089 160
rect 7145 104 7231 160
rect 7287 104 7373 160
rect 7429 104 7515 160
rect 7571 104 7657 160
rect 7713 104 7799 160
rect 7855 104 7941 160
rect 7997 104 8083 160
rect 8139 104 8225 160
rect 8281 104 8367 160
rect 8423 104 8509 160
rect 8565 104 8651 160
rect 8707 104 8793 160
rect 8849 104 8935 160
rect 8991 104 9077 160
rect 9133 104 9219 160
rect 9275 104 9361 160
rect 9417 104 9503 160
rect 9559 104 9645 160
rect 9701 104 9787 160
rect 9843 104 9929 160
rect 9985 104 10071 160
rect 10127 104 10213 160
rect 10269 104 10355 160
rect 10411 104 10497 160
rect 10553 104 10639 160
rect 10695 104 10781 160
rect 10837 104 10923 160
rect 10979 104 11065 160
rect 11121 104 11207 160
rect 11263 104 11349 160
rect 11405 104 11491 160
rect 11547 104 11633 160
rect 11689 104 11775 160
rect 11831 104 11917 160
rect 11973 104 12059 160
rect 12115 104 12201 160
rect 12257 104 12343 160
rect 12399 150 12526 160
rect 12582 150 12650 206
rect 12706 150 12774 206
rect 12830 150 12898 206
rect 12954 150 13022 206
rect 13078 150 13200 206
rect 12399 104 13200 150
rect -400 0 13200 104
<< glass >>
rect 400 400 12400 12400
use M3_M2_CDNS_40661954729333  M3_M2_CDNS_40661954729333_0
timestamp 1698431365
transform 0 -1 -10 1 0 6254
box 0 0 1 1
use M3_M2_CDNS_40661954729333  M3_M2_CDNS_40661954729333_1
timestamp 1698431365
transform 0 -1 12802 1 0 6254
box 0 0 1 1
use M3_M2_CDNS_40661954729334  M3_M2_CDNS_40661954729334_0
timestamp 1698431365
transform 1 0 6407 0 1 203
box 0 0 1 1
use M3_M2_CDNS_40661954729335  M3_M2_CDNS_40661954729335_0
timestamp 1698431365
transform 1 0 6408 0 1 12735
box 0 0 1 1
use M3_M2_CDNS_40661954729336  M3_M2_CDNS_40661954729336_0
timestamp 1698431365
transform 0 -1 12040 1 0 6389
box 0 0 1 1
use M3_M2_CDNS_40661954729336  M3_M2_CDNS_40661954729336_1
timestamp 1698431365
transform 0 -1 11635 1 0 6389
box 0 0 1 1
use M3_M2_CDNS_40661954729336  M3_M2_CDNS_40661954729336_2
timestamp 1698431365
transform 0 -1 11235 1 0 6389
box 0 0 1 1
use M3_M2_CDNS_40661954729336  M3_M2_CDNS_40661954729336_3
timestamp 1698431365
transform 0 -1 10830 1 0 6389
box 0 0 1 1
use M3_M2_CDNS_40661954729336  M3_M2_CDNS_40661954729336_4
timestamp 1698431365
transform 0 -1 10433 1 0 6389
box 0 0 1 1
use M3_M2_CDNS_40661954729336  M3_M2_CDNS_40661954729336_5
timestamp 1698431365
transform 0 -1 10033 1 0 6389
box 0 0 1 1
use M3_M2_CDNS_40661954729336  M3_M2_CDNS_40661954729336_6
timestamp 1698431365
transform 0 -1 9637 1 0 6389
box 0 0 1 1
use M3_M2_CDNS_40661954729336  M3_M2_CDNS_40661954729336_7
timestamp 1698431365
transform 0 -1 9233 1 0 6389
box 0 0 1 1
use M3_M2_CDNS_40661954729336  M3_M2_CDNS_40661954729336_8
timestamp 1698431365
transform 0 -1 8836 1 0 6389
box 0 0 1 1
use M3_M2_CDNS_40661954729336  M3_M2_CDNS_40661954729336_9
timestamp 1698431365
transform 0 -1 8439 1 0 6389
box 0 0 1 1
use M3_M2_CDNS_40661954729336  M3_M2_CDNS_40661954729336_10
timestamp 1698431365
transform 0 -1 8039 1 0 6389
box 0 0 1 1
use M3_M2_CDNS_40661954729336  M3_M2_CDNS_40661954729336_11
timestamp 1698431365
transform 0 -1 7638 1 0 6389
box 0 0 1 1
use M3_M2_CDNS_40661954729336  M3_M2_CDNS_40661954729336_12
timestamp 1698431365
transform 0 -1 2435 1 0 6389
box 0 0 1 1
use M3_M2_CDNS_40661954729336  M3_M2_CDNS_40661954729336_13
timestamp 1698431365
transform 0 -1 2038 1 0 6389
box 0 0 1 1
use M3_M2_CDNS_40661954729336  M3_M2_CDNS_40661954729336_14
timestamp 1698431365
transform 0 -1 840 1 0 6389
box 0 0 1 1
use M3_M2_CDNS_40661954729336  M3_M2_CDNS_40661954729336_15
timestamp 1698431365
transform 0 -1 1641 1 0 6389
box 0 0 1 1
use M3_M2_CDNS_40661954729336  M3_M2_CDNS_40661954729336_16
timestamp 1698431365
transform 0 -1 1241 1 0 6389
box 0 0 1 1
use M3_M2_CDNS_40661954729336  M3_M2_CDNS_40661954729336_17
timestamp 1698431365
transform 0 -1 2839 1 0 6389
box 0 0 1 1
use M3_M2_CDNS_40661954729336  M3_M2_CDNS_40661954729336_18
timestamp 1698431365
transform 0 -1 3235 1 0 6389
box 0 0 1 1
use M3_M2_CDNS_40661954729336  M3_M2_CDNS_40661954729336_19
timestamp 1698431365
transform 0 -1 7244 1 0 6389
box 0 0 1 1
use M3_M2_CDNS_40661954729336  M3_M2_CDNS_40661954729336_20
timestamp 1698431365
transform 0 -1 4032 1 0 6389
box 0 0 1 1
use M3_M2_CDNS_40661954729336  M3_M2_CDNS_40661954729336_21
timestamp 1698431365
transform 0 -1 4437 1 0 6389
box 0 0 1 1
use M3_M2_CDNS_40661954729336  M3_M2_CDNS_40661954729336_22
timestamp 1698431365
transform 0 -1 4837 1 0 6389
box 0 0 1 1
use M3_M2_CDNS_40661954729336  M3_M2_CDNS_40661954729336_23
timestamp 1698431365
transform 0 -1 5242 1 0 6389
box 0 0 1 1
use M3_M2_CDNS_40661954729336  M3_M2_CDNS_40661954729336_24
timestamp 1698431365
transform 0 -1 5639 1 0 6389
box 0 0 1 1
use M3_M2_CDNS_40661954729336  M3_M2_CDNS_40661954729336_25
timestamp 1698431365
transform 0 -1 6036 1 0 6389
box 0 0 1 1
use M3_M2_CDNS_40661954729336  M3_M2_CDNS_40661954729336_26
timestamp 1698431365
transform 0 -1 6439 1 0 6389
box 0 0 1 1
use M3_M2_CDNS_40661954729336  M3_M2_CDNS_40661954729336_27
timestamp 1698431365
transform 0 -1 6841 1 0 6389
box 0 0 1 1
use M3_M2_CDNS_40661954729336  M3_M2_CDNS_40661954729336_28
timestamp 1698431365
transform 0 -1 3635 1 0 6389
box 0 0 1 1
use M4_M3_CDNS_40661954729337  M4_M3_CDNS_40661954729337_0
timestamp 1698431365
transform 0 -1 12802 1 0 6254
box 0 0 1 1
use M4_M3_CDNS_40661954729337  M4_M3_CDNS_40661954729337_1
timestamp 1698431365
transform 0 -1 -10 1 0 6254
box 0 0 1 1
use M4_M3_CDNS_40661954729338  M4_M3_CDNS_40661954729338_0
timestamp 1698431365
transform 1 0 6408 0 1 12735
box 0 0 1 1
use M4_M3_CDNS_40661954729339  M4_M3_CDNS_40661954729339_0
timestamp 1698431365
transform 1 0 6407 0 1 203
box 0 0 1 1
use M4_M3_CDNS_40661954729340  M4_M3_CDNS_40661954729340_0
timestamp 1698431365
transform 0 -1 11635 1 0 6389
box 0 0 1 1
use M4_M3_CDNS_40661954729340  M4_M3_CDNS_40661954729340_1
timestamp 1698431365
transform 0 -1 11235 1 0 6389
box 0 0 1 1
use M4_M3_CDNS_40661954729340  M4_M3_CDNS_40661954729340_2
timestamp 1698431365
transform 0 -1 10830 1 0 6389
box 0 0 1 1
use M4_M3_CDNS_40661954729340  M4_M3_CDNS_40661954729340_3
timestamp 1698431365
transform 0 -1 10433 1 0 6389
box 0 0 1 1
use M4_M3_CDNS_40661954729340  M4_M3_CDNS_40661954729340_4
timestamp 1698431365
transform 0 -1 10033 1 0 6389
box 0 0 1 1
use M4_M3_CDNS_40661954729340  M4_M3_CDNS_40661954729340_5
timestamp 1698431365
transform 0 -1 9637 1 0 6389
box 0 0 1 1
use M4_M3_CDNS_40661954729340  M4_M3_CDNS_40661954729340_6
timestamp 1698431365
transform 0 -1 9233 1 0 6389
box 0 0 1 1
use M4_M3_CDNS_40661954729340  M4_M3_CDNS_40661954729340_7
timestamp 1698431365
transform 0 -1 8836 1 0 6389
box 0 0 1 1
use M4_M3_CDNS_40661954729340  M4_M3_CDNS_40661954729340_8
timestamp 1698431365
transform 0 -1 8439 1 0 6389
box 0 0 1 1
use M4_M3_CDNS_40661954729340  M4_M3_CDNS_40661954729340_9
timestamp 1698431365
transform 0 -1 8039 1 0 6389
box 0 0 1 1
use M4_M3_CDNS_40661954729340  M4_M3_CDNS_40661954729340_10
timestamp 1698431365
transform 0 -1 7638 1 0 6389
box 0 0 1 1
use M4_M3_CDNS_40661954729340  M4_M3_CDNS_40661954729340_11
timestamp 1698431365
transform 0 -1 7244 1 0 6389
box 0 0 1 1
use M4_M3_CDNS_40661954729340  M4_M3_CDNS_40661954729340_12
timestamp 1698431365
transform 0 -1 6841 1 0 6389
box 0 0 1 1
use M4_M3_CDNS_40661954729340  M4_M3_CDNS_40661954729340_13
timestamp 1698431365
transform 0 -1 6439 1 0 6389
box 0 0 1 1
use M4_M3_CDNS_40661954729340  M4_M3_CDNS_40661954729340_14
timestamp 1698431365
transform 0 -1 6036 1 0 6389
box 0 0 1 1
use M4_M3_CDNS_40661954729340  M4_M3_CDNS_40661954729340_15
timestamp 1698431365
transform 0 -1 12040 1 0 6389
box 0 0 1 1
use M4_M3_CDNS_40661954729340  M4_M3_CDNS_40661954729340_16
timestamp 1698431365
transform 0 -1 840 1 0 6389
box 0 0 1 1
use M4_M3_CDNS_40661954729340  M4_M3_CDNS_40661954729340_17
timestamp 1698431365
transform 0 -1 1241 1 0 6389
box 0 0 1 1
use M4_M3_CDNS_40661954729340  M4_M3_CDNS_40661954729340_18
timestamp 1698431365
transform 0 -1 1641 1 0 6389
box 0 0 1 1
use M4_M3_CDNS_40661954729340  M4_M3_CDNS_40661954729340_19
timestamp 1698431365
transform 0 -1 2038 1 0 6389
box 0 0 1 1
use M4_M3_CDNS_40661954729340  M4_M3_CDNS_40661954729340_20
timestamp 1698431365
transform 0 -1 2435 1 0 6389
box 0 0 1 1
use M4_M3_CDNS_40661954729340  M4_M3_CDNS_40661954729340_21
timestamp 1698431365
transform 0 -1 2839 1 0 6389
box 0 0 1 1
use M4_M3_CDNS_40661954729340  M4_M3_CDNS_40661954729340_22
timestamp 1698431365
transform 0 -1 3235 1 0 6389
box 0 0 1 1
use M4_M3_CDNS_40661954729340  M4_M3_CDNS_40661954729340_23
timestamp 1698431365
transform 0 -1 3635 1 0 6389
box 0 0 1 1
use M4_M3_CDNS_40661954729340  M4_M3_CDNS_40661954729340_24
timestamp 1698431365
transform 0 -1 4032 1 0 6389
box 0 0 1 1
use M4_M3_CDNS_40661954729340  M4_M3_CDNS_40661954729340_25
timestamp 1698431365
transform 0 -1 4437 1 0 6389
box 0 0 1 1
use M4_M3_CDNS_40661954729340  M4_M3_CDNS_40661954729340_26
timestamp 1698431365
transform 0 -1 4837 1 0 6389
box 0 0 1 1
use M4_M3_CDNS_40661954729340  M4_M3_CDNS_40661954729340_27
timestamp 1698431365
transform 0 -1 5639 1 0 6389
box 0 0 1 1
use M4_M3_CDNS_40661954729340  M4_M3_CDNS_40661954729340_28
timestamp 1698431365
transform 0 -1 5242 1 0 6389
box 0 0 1 1
<< properties >>
string GDS_END 506756
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 498266
string path 5.000 311.025 5.000 6.350 
<< end >>
