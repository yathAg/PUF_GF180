magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 377 3670 870
rect -86 352 2919 377
rect 3171 352 3670 377
<< pwell >>
rect 2919 352 3171 377
rect -86 -86 3670 352
<< mvnmos >>
rect 124 68 244 232
rect 308 68 428 232
rect 532 68 652 232
rect 716 68 836 232
rect 940 68 1060 232
rect 1124 68 1244 232
rect 1348 68 1468 232
rect 1532 68 1652 232
rect 1828 68 1948 232
rect 2012 68 2132 232
rect 2236 68 2356 232
rect 2420 68 2540 232
rect 2644 68 2764 232
rect 2828 68 2948 232
rect 3140 68 3260 232
rect 3324 68 3444 232
<< mvpmos >>
rect 124 497 224 716
rect 328 497 428 716
rect 532 497 632 716
rect 736 497 836 716
rect 940 497 1040 716
rect 1144 497 1244 716
rect 1348 497 1448 716
rect 1552 497 1652 716
rect 1828 497 1928 716
rect 2032 497 2132 716
rect 2236 497 2336 716
rect 2440 497 2540 716
rect 2644 497 2744 716
rect 2848 497 2948 716
rect 3140 497 3240 716
rect 3344 497 3444 716
<< mvndiff >>
rect 3008 244 3080 257
rect 3008 232 3021 244
rect 36 128 124 232
rect 36 82 49 128
rect 95 82 124 128
rect 36 68 124 82
rect 244 68 308 232
rect 428 160 532 232
rect 428 114 457 160
rect 503 114 532 160
rect 428 68 532 114
rect 652 68 716 232
rect 836 127 940 232
rect 836 81 865 127
rect 911 81 940 127
rect 836 68 940 81
rect 1060 68 1124 232
rect 1244 171 1348 232
rect 1244 125 1273 171
rect 1319 125 1348 171
rect 1244 68 1348 125
rect 1468 68 1532 232
rect 1652 127 1828 232
rect 1652 81 1681 127
rect 1727 81 1828 127
rect 1652 68 1828 81
rect 1948 68 2012 232
rect 2132 178 2236 232
rect 2132 132 2161 178
rect 2207 132 2236 178
rect 2132 68 2236 132
rect 2356 68 2420 232
rect 2540 135 2644 232
rect 2540 89 2569 135
rect 2615 89 2644 135
rect 2540 68 2644 89
rect 2764 68 2828 232
rect 2948 198 3021 232
rect 3067 232 3080 244
rect 3067 198 3140 232
rect 2948 68 3140 198
rect 3260 68 3324 232
rect 3444 135 3532 232
rect 3444 89 3473 135
rect 3519 89 3532 135
rect 3444 68 3532 89
<< mvpdiff >>
rect 36 659 124 716
rect 36 519 49 659
rect 95 519 124 659
rect 36 497 124 519
rect 224 659 328 716
rect 224 613 253 659
rect 299 613 328 659
rect 224 497 328 613
rect 428 659 532 716
rect 428 519 457 659
rect 503 519 532 659
rect 428 497 532 519
rect 632 659 736 716
rect 632 613 661 659
rect 707 613 736 659
rect 632 497 736 613
rect 836 659 940 716
rect 836 519 865 659
rect 911 519 940 659
rect 836 497 940 519
rect 1040 659 1144 716
rect 1040 613 1069 659
rect 1115 613 1144 659
rect 1040 497 1144 613
rect 1244 659 1348 716
rect 1244 519 1273 659
rect 1319 519 1348 659
rect 1244 497 1348 519
rect 1448 659 1552 716
rect 1448 613 1477 659
rect 1523 613 1552 659
rect 1448 497 1552 613
rect 1652 659 1828 716
rect 1652 519 1681 659
rect 1727 519 1828 659
rect 1652 497 1828 519
rect 1928 581 2032 716
rect 1928 535 1957 581
rect 2003 535 2032 581
rect 1928 497 2032 535
rect 2132 678 2236 716
rect 2132 632 2161 678
rect 2207 632 2236 678
rect 2132 497 2236 632
rect 2336 581 2440 716
rect 2336 535 2365 581
rect 2411 535 2440 581
rect 2336 497 2440 535
rect 2540 678 2644 716
rect 2540 632 2569 678
rect 2615 632 2644 678
rect 2540 497 2644 632
rect 2744 581 2848 716
rect 2744 535 2773 581
rect 2819 535 2848 581
rect 2744 497 2848 535
rect 2948 678 3140 716
rect 2948 632 3065 678
rect 3111 632 3140 678
rect 2948 497 3140 632
rect 3240 581 3344 716
rect 3240 535 3269 581
rect 3315 535 3344 581
rect 3240 497 3344 535
rect 3444 659 3532 716
rect 3444 519 3473 659
rect 3519 519 3532 659
rect 3444 497 3532 519
<< mvndiffc >>
rect 49 82 95 128
rect 457 114 503 160
rect 865 81 911 127
rect 1273 125 1319 171
rect 1681 81 1727 127
rect 2161 132 2207 178
rect 2569 89 2615 135
rect 3021 198 3067 244
rect 3473 89 3519 135
<< mvpdiffc >>
rect 49 519 95 659
rect 253 613 299 659
rect 457 519 503 659
rect 661 613 707 659
rect 865 519 911 659
rect 1069 613 1115 659
rect 1273 519 1319 659
rect 1477 613 1523 659
rect 1681 519 1727 659
rect 1957 535 2003 581
rect 2161 632 2207 678
rect 2365 535 2411 581
rect 2569 632 2615 678
rect 2773 535 2819 581
rect 3065 632 3111 678
rect 3269 535 3315 581
rect 3473 519 3519 659
<< polysilicon >>
rect 124 716 224 760
rect 328 716 428 760
rect 532 716 632 760
rect 736 716 836 760
rect 940 716 1040 760
rect 1144 716 1244 760
rect 1348 716 1448 760
rect 1552 716 1652 760
rect 1828 716 1928 760
rect 2032 716 2132 760
rect 2236 716 2336 760
rect 2440 716 2540 760
rect 2644 716 2744 760
rect 2848 716 2948 760
rect 3140 716 3240 760
rect 3344 716 3444 760
rect 124 394 224 497
rect 124 348 137 394
rect 183 348 224 394
rect 124 288 224 348
rect 328 415 428 497
rect 328 369 359 415
rect 405 394 428 415
rect 532 415 632 497
rect 532 394 565 415
rect 405 369 565 394
rect 611 369 632 415
rect 328 348 632 369
rect 328 288 428 348
rect 124 232 244 288
rect 308 232 428 288
rect 532 288 632 348
rect 736 394 836 497
rect 940 394 1040 497
rect 736 348 1040 394
rect 736 311 836 348
rect 736 288 761 311
rect 532 232 652 288
rect 716 265 761 288
rect 807 265 836 311
rect 716 232 836 265
rect 940 311 1040 348
rect 940 265 969 311
rect 1015 288 1040 311
rect 1144 415 1244 497
rect 1144 369 1170 415
rect 1216 394 1244 415
rect 1348 415 1448 497
rect 1348 394 1377 415
rect 1216 369 1377 394
rect 1423 369 1448 415
rect 1144 348 1448 369
rect 1144 288 1244 348
rect 1015 265 1060 288
rect 940 232 1060 265
rect 1124 232 1244 288
rect 1348 288 1448 348
rect 1552 324 1652 497
rect 1532 311 1652 324
rect 1348 232 1468 288
rect 1532 265 1567 311
rect 1613 265 1652 311
rect 1532 232 1652 265
rect 1828 412 1928 497
rect 1828 399 1948 412
rect 1828 353 1889 399
rect 1935 353 1948 399
rect 1828 232 1948 353
rect 2032 394 2132 497
rect 2236 415 2336 497
rect 2236 394 2272 415
rect 2032 369 2272 394
rect 2318 369 2336 415
rect 2032 348 2336 369
rect 2032 288 2132 348
rect 2012 232 2132 288
rect 2236 288 2336 348
rect 2440 365 2540 497
rect 2644 365 2744 497
rect 2440 312 2744 365
rect 2440 288 2464 312
rect 2236 232 2356 288
rect 2420 266 2464 288
rect 2510 292 2673 312
rect 2510 266 2540 292
rect 2420 232 2540 266
rect 2644 266 2673 292
rect 2719 288 2744 312
rect 2848 415 2948 497
rect 2848 369 2872 415
rect 2918 369 2948 415
rect 2848 358 2948 369
rect 3140 358 3240 497
rect 3344 428 3444 497
rect 3344 407 3364 428
rect 2848 318 3240 358
rect 2848 288 2948 318
rect 2719 266 2764 288
rect 2644 232 2764 266
rect 2828 232 2948 288
rect 3140 288 3240 318
rect 3324 288 3364 407
rect 3410 288 3444 428
rect 3140 232 3260 288
rect 3324 232 3444 288
rect 124 24 244 68
rect 308 24 428 68
rect 532 24 652 68
rect 716 24 836 68
rect 940 24 1060 68
rect 1124 24 1244 68
rect 1348 24 1468 68
rect 1532 24 1652 68
rect 1828 24 1948 68
rect 2012 24 2132 68
rect 2236 24 2356 68
rect 2420 24 2540 68
rect 2644 24 2764 68
rect 2828 24 2948 68
rect 3140 24 3260 68
rect 3324 24 3444 68
<< polycontact >>
rect 137 348 183 394
rect 359 369 405 415
rect 565 369 611 415
rect 761 265 807 311
rect 969 265 1015 311
rect 1170 369 1216 415
rect 1377 369 1423 415
rect 1567 265 1613 311
rect 1889 353 1935 399
rect 2272 369 2318 415
rect 2464 266 2510 312
rect 2673 266 2719 312
rect 2872 369 2918 415
rect 3364 288 3410 428
<< metal1 >>
rect 0 724 3584 844
rect 38 659 106 678
rect 38 519 49 659
rect 95 543 106 659
rect 242 659 310 724
rect 242 613 253 659
rect 299 613 310 659
rect 242 602 310 613
rect 446 659 514 678
rect 446 543 457 659
rect 95 519 457 543
rect 503 543 514 659
rect 650 659 718 724
rect 650 613 661 659
rect 707 613 718 659
rect 650 602 718 613
rect 854 659 922 678
rect 854 543 865 659
rect 503 519 865 543
rect 911 543 922 659
rect 1058 659 1126 724
rect 1058 613 1069 659
rect 1115 613 1126 659
rect 1058 602 1126 613
rect 1262 659 1330 678
rect 1262 543 1273 659
rect 911 519 1273 543
rect 1319 543 1330 659
rect 1466 659 1534 724
rect 1466 613 1477 659
rect 1523 613 1534 659
rect 1466 602 1534 613
rect 1670 659 2161 678
rect 1670 543 1681 659
rect 1319 519 1681 543
rect 1727 632 2161 659
rect 2207 632 2569 678
rect 2615 632 3065 678
rect 3111 659 3530 678
rect 3111 632 3473 659
rect 1727 519 1738 632
rect 38 497 1738 519
rect 1797 581 3334 582
rect 1797 535 1957 581
rect 2003 535 2365 581
rect 2411 535 2773 581
rect 2819 535 3269 581
rect 3315 535 3334 581
rect 1797 534 3334 535
rect 124 394 204 445
rect 124 348 137 394
rect 183 348 204 394
rect 328 415 1448 426
rect 328 369 359 415
rect 405 369 565 415
rect 611 369 1170 415
rect 1216 369 1377 415
rect 1423 369 1448 415
rect 328 360 1448 369
rect 124 312 204 348
rect 124 311 1624 312
rect 124 265 761 311
rect 807 265 969 311
rect 1015 265 1567 311
rect 1613 265 1624 311
rect 124 246 675 265
rect 1797 219 1843 534
rect 1889 399 2104 428
rect 1935 353 2104 399
rect 2236 415 2946 424
rect 2236 369 2272 415
rect 2318 369 2872 415
rect 2918 369 2946 415
rect 2236 360 2946 369
rect 1889 342 2104 353
rect 2032 312 2104 342
rect 2032 266 2464 312
rect 2510 266 2673 312
rect 2719 266 2802 312
rect 2032 248 2802 266
rect 753 200 1843 219
rect 753 178 2236 200
rect 753 173 2161 178
rect 753 160 799 173
rect 49 128 95 139
rect 445 114 457 160
rect 503 114 799 160
rect 1273 171 1319 173
rect 49 60 95 82
rect 854 81 865 127
rect 911 81 922 127
rect 1797 132 2161 173
rect 2207 132 2236 178
rect 2756 152 2802 248
rect 3010 244 3116 534
rect 3462 519 3473 632
rect 3519 519 3530 659
rect 3462 497 3530 519
rect 3010 198 3021 244
rect 3067 198 3116 244
rect 3364 428 3410 447
rect 3364 152 3410 288
rect 1273 114 1319 125
rect 854 60 922 81
rect 1670 81 1681 127
rect 1727 81 1738 127
rect 1797 106 2236 132
rect 2569 135 2615 146
rect 1670 60 1738 81
rect 2756 106 3410 152
rect 3473 135 3519 146
rect 2569 60 2615 89
rect 3473 60 3519 89
rect 0 -60 3584 60
<< labels >>
flabel metal1 s 3364 428 3410 447 0 FreeSans 600 0 0 0 A2
port 2 nsew default input
flabel metal1 s 328 360 1448 426 0 FreeSans 600 0 0 0 B1
port 3 nsew default input
flabel metal1 s 124 312 204 445 0 FreeSans 600 0 0 0 B2
port 4 nsew default input
flabel metal1 s 0 724 3584 844 0 FreeSans 600 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 3473 139 3519 146 0 FreeSans 600 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel metal1 s 1797 534 3334 582 0 FreeSans 600 0 0 0 ZN
port 5 nsew default output
flabel metal1 s 2236 360 2946 424 0 FreeSans 600 0 0 0 A1
port 1 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 7 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 8 nsew ground bidirectional
rlabel metal1 s 3364 342 3410 428 1 A2
port 2 nsew default input
rlabel metal1 s 1889 342 2104 428 1 A2
port 2 nsew default input
rlabel metal1 s 3364 312 3410 342 1 A2
port 2 nsew default input
rlabel metal1 s 2032 312 2104 342 1 A2
port 2 nsew default input
rlabel metal1 s 3364 248 3410 312 1 A2
port 2 nsew default input
rlabel metal1 s 2032 248 2802 312 1 A2
port 2 nsew default input
rlabel metal1 s 3364 152 3410 248 1 A2
port 2 nsew default input
rlabel metal1 s 2756 152 2802 248 1 A2
port 2 nsew default input
rlabel metal1 s 2756 106 3410 152 1 A2
port 2 nsew default input
rlabel metal1 s 124 265 1624 312 1 B2
port 4 nsew default input
rlabel metal1 s 124 246 675 265 1 B2
port 4 nsew default input
rlabel metal1 s 3010 219 3116 534 1 ZN
port 5 nsew default output
rlabel metal1 s 1797 219 1843 534 1 ZN
port 5 nsew default output
rlabel metal1 s 3010 200 3116 219 1 ZN
port 5 nsew default output
rlabel metal1 s 753 200 1843 219 1 ZN
port 5 nsew default output
rlabel metal1 s 3010 198 3116 200 1 ZN
port 5 nsew default output
rlabel metal1 s 753 198 2236 200 1 ZN
port 5 nsew default output
rlabel metal1 s 753 173 2236 198 1 ZN
port 5 nsew default output
rlabel metal1 s 1797 160 2236 173 1 ZN
port 5 nsew default output
rlabel metal1 s 1273 160 1319 173 1 ZN
port 5 nsew default output
rlabel metal1 s 753 160 799 173 1 ZN
port 5 nsew default output
rlabel metal1 s 1797 114 2236 160 1 ZN
port 5 nsew default output
rlabel metal1 s 1273 114 1319 160 1 ZN
port 5 nsew default output
rlabel metal1 s 445 114 799 160 1 ZN
port 5 nsew default output
rlabel metal1 s 1797 106 2236 114 1 ZN
port 5 nsew default output
rlabel metal1 s 1466 602 1534 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1058 602 1126 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 650 602 718 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 242 602 310 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2569 139 2615 146 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3473 127 3519 139 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2569 127 2615 139 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 49 127 95 139 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3473 60 3519 127 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2569 60 2615 127 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1670 60 1738 127 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 854 60 922 127 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 127 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3584 60 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3584 784
string GDS_END 1276460
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1269310
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
