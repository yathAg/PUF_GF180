magic
tech gf180mcuA
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 453 1990 1094
<< pwell >>
rect -86 -86 1990 453
<< mvnmos >>
rect 124 69 244 333
rect 348 69 468 333
rect 572 69 692 333
rect 796 69 916 333
rect 1026 69 1146 333
rect 1220 69 1340 333
rect 1444 69 1564 333
rect 1628 69 1748 333
<< mvpmos >>
rect 144 573 244 939
rect 358 573 458 939
rect 582 573 682 939
rect 796 573 896 939
rect 1036 647 1136 939
rect 1240 647 1340 939
rect 1444 647 1544 939
rect 1648 647 1748 939
<< mvndiff >>
rect 36 305 124 333
rect 36 165 49 305
rect 95 165 124 305
rect 36 69 124 165
rect 244 285 348 333
rect 244 239 273 285
rect 319 239 348 285
rect 244 69 348 239
rect 468 211 572 333
rect 468 165 497 211
rect 543 165 572 211
rect 468 69 572 165
rect 692 314 796 333
rect 692 268 721 314
rect 767 268 796 314
rect 692 69 796 268
rect 916 305 1026 333
rect 916 165 945 305
rect 991 165 1026 305
rect 916 69 1026 165
rect 1146 69 1220 333
rect 1340 294 1444 333
rect 1340 154 1369 294
rect 1415 154 1444 294
rect 1340 69 1444 154
rect 1564 69 1628 333
rect 1748 305 1836 333
rect 1748 165 1777 305
rect 1823 165 1836 305
rect 1748 69 1836 165
<< mvpdiff >>
rect 56 923 144 939
rect 56 783 69 923
rect 115 783 144 923
rect 56 573 144 783
rect 244 573 358 939
rect 458 861 582 939
rect 458 721 487 861
rect 533 721 582 861
rect 458 573 582 721
rect 682 573 796 939
rect 896 923 1036 939
rect 896 783 925 923
rect 971 783 1036 923
rect 896 647 1036 783
rect 1136 861 1240 939
rect 1136 721 1165 861
rect 1211 721 1240 861
rect 1136 647 1240 721
rect 1340 923 1444 939
rect 1340 783 1369 923
rect 1415 783 1444 923
rect 1340 647 1444 783
rect 1544 861 1648 939
rect 1544 721 1573 861
rect 1619 721 1648 861
rect 1544 647 1648 721
rect 1748 923 1836 939
rect 1748 783 1777 923
rect 1823 783 1836 923
rect 1748 647 1836 783
rect 896 573 976 647
<< mvndiffc >>
rect 49 165 95 305
rect 273 239 319 285
rect 497 165 543 211
rect 721 268 767 314
rect 945 165 991 305
rect 1369 154 1415 294
rect 1777 165 1823 305
<< mvpdiffc >>
rect 69 783 115 923
rect 487 721 533 861
rect 925 783 971 923
rect 1165 721 1211 861
rect 1369 783 1415 923
rect 1573 721 1619 861
rect 1777 783 1823 923
<< polysilicon >>
rect 144 939 244 983
rect 358 939 458 983
rect 582 939 682 983
rect 796 939 896 983
rect 1036 939 1136 983
rect 1240 939 1340 983
rect 1444 939 1544 983
rect 1648 939 1748 983
rect 144 513 244 573
rect 358 513 458 573
rect 582 513 682 573
rect 144 500 310 513
rect 144 454 251 500
rect 297 454 310 500
rect 144 441 310 454
rect 358 500 682 513
rect 358 454 371 500
rect 417 454 682 500
rect 358 441 682 454
rect 144 377 244 441
rect 358 377 468 441
rect 124 333 244 377
rect 348 333 468 377
rect 572 377 682 441
rect 796 500 896 573
rect 796 454 809 500
rect 855 454 896 500
rect 796 377 896 454
rect 1036 500 1136 647
rect 1036 454 1077 500
rect 1123 454 1136 500
rect 1036 377 1136 454
rect 1240 513 1340 647
rect 1444 513 1544 647
rect 1240 500 1544 513
rect 1240 454 1257 500
rect 1303 454 1544 500
rect 1240 441 1544 454
rect 1240 377 1340 441
rect 572 333 692 377
rect 796 333 916 377
rect 1026 333 1146 377
rect 1220 333 1340 377
rect 1444 377 1544 441
rect 1648 500 1748 647
rect 1648 454 1661 500
rect 1707 454 1748 500
rect 1648 377 1748 454
rect 1444 333 1564 377
rect 1628 333 1748 377
rect 124 25 244 69
rect 348 25 468 69
rect 572 25 692 69
rect 796 25 916 69
rect 1026 25 1146 69
rect 1220 25 1340 69
rect 1444 25 1564 69
rect 1628 25 1748 69
<< polycontact >>
rect 251 454 297 500
rect 371 454 417 500
rect 809 454 855 500
rect 1077 454 1123 500
rect 1257 454 1303 500
rect 1661 454 1707 500
<< metal1 >>
rect 0 923 1904 1098
rect 0 918 69 923
rect 115 918 925 923
rect 69 772 115 783
rect 173 861 533 872
rect 173 814 487 861
rect 173 716 219 814
rect 148 675 219 716
rect 971 918 1369 923
rect 925 772 971 783
rect 1165 861 1211 872
rect 533 721 1165 726
rect 1415 918 1777 923
rect 1369 772 1415 783
rect 1573 861 1619 872
rect 1211 721 1573 726
rect 1823 918 1904 923
rect 1777 772 1823 783
rect 487 680 1619 721
rect 49 305 95 316
rect 148 314 194 675
rect 240 588 524 634
rect 240 500 308 588
rect 478 542 524 588
rect 1066 588 1707 634
rect 240 454 251 500
rect 297 454 308 500
rect 359 500 418 542
rect 359 454 371 500
rect 417 454 418 500
rect 478 500 866 542
rect 478 454 809 500
rect 855 454 866 500
rect 1066 500 1134 588
rect 1066 454 1077 500
rect 1123 454 1134 500
rect 1246 500 1314 542
rect 1246 454 1257 500
rect 1303 454 1314 500
rect 1374 500 1707 588
rect 1374 454 1661 500
rect 359 443 418 454
rect 1374 443 1707 454
rect 945 351 1823 397
rect 148 285 721 314
rect 148 239 273 285
rect 319 268 721 285
rect 767 268 778 314
rect 945 305 991 351
rect 1777 305 1823 351
rect 148 228 319 239
rect 497 211 945 222
rect 95 165 497 182
rect 543 165 945 211
rect 49 136 991 165
rect 1369 294 1415 305
rect 1777 154 1823 165
rect 1369 90 1415 154
rect 0 -90 1904 90
<< labels >>
flabel metal1 s 359 443 418 542 0 FreeSans 200 0 0 0 A1
port 1 nsew default input
flabel metal1 s 240 588 524 634 0 FreeSans 200 0 0 0 A2
port 2 nsew default input
flabel metal1 s 1066 588 1707 634 0 FreeSans 200 0 0 0 B
port 3 nsew default input
flabel metal1 s 1246 454 1314 542 0 FreeSans 200 0 0 0 C
port 4 nsew default input
flabel metal1 s 0 918 1904 1098 0 FreeSans 200 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 1369 90 1415 305 0 FreeSans 200 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel metal1 s 1573 814 1619 872 0 FreeSans 200 0 0 0 ZN
port 5 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 7 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 8 nsew ground bidirectional
rlabel metal1 s 478 542 524 588 1 A2
port 2 nsew default input
rlabel metal1 s 240 542 308 588 1 A2
port 2 nsew default input
rlabel metal1 s 478 454 866 542 1 A2
port 2 nsew default input
rlabel metal1 s 240 454 308 542 1 A2
port 2 nsew default input
rlabel metal1 s 1374 454 1707 588 1 B
port 3 nsew default input
rlabel metal1 s 1066 454 1134 588 1 B
port 3 nsew default input
rlabel metal1 s 1374 443 1707 454 1 B
port 3 nsew default input
rlabel metal1 s 1165 814 1211 872 1 ZN
port 5 nsew default output
rlabel metal1 s 173 814 533 872 1 ZN
port 5 nsew default output
rlabel metal1 s 1573 726 1619 814 1 ZN
port 5 nsew default output
rlabel metal1 s 1165 726 1211 814 1 ZN
port 5 nsew default output
rlabel metal1 s 487 726 533 814 1 ZN
port 5 nsew default output
rlabel metal1 s 173 726 219 814 1 ZN
port 5 nsew default output
rlabel metal1 s 487 716 1619 726 1 ZN
port 5 nsew default output
rlabel metal1 s 173 716 219 726 1 ZN
port 5 nsew default output
rlabel metal1 s 487 680 1619 716 1 ZN
port 5 nsew default output
rlabel metal1 s 148 680 219 716 1 ZN
port 5 nsew default output
rlabel metal1 s 148 675 219 680 1 ZN
port 5 nsew default output
rlabel metal1 s 148 314 194 675 1 ZN
port 5 nsew default output
rlabel metal1 s 148 268 778 314 1 ZN
port 5 nsew default output
rlabel metal1 s 148 228 319 268 1 ZN
port 5 nsew default output
rlabel metal1 s 1777 772 1823 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1369 772 1415 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 925 772 971 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 69 772 115 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 -90 1904 90 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1904 1008
string GDS_END 212564
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 207412
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
