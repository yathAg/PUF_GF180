************************************************************************
* auCdl Netlist:
* 
* Library Name:  TCG_Library
* Top Cell Name: nplus_u
* View Name:     schematic
* Netlisted on:  Nov 24 09:29:33 2021
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM

*.GLOBAL gnd!

*.PIN gnd!

************************************************************************
* Library Name: TCG_Library
* Cell Name:    nplus_u
* View Name:    schematic
************************************************************************

.SUBCKT nplus_u I1_0_0_0_0_0_R0_MINUS I1_0_0_0_0_0_R0_PLUS 
+ I1_0_0_0_1_0_R0_MINUS I1_0_0_0_1_0_R0_PLUS I1_0_0_1_0_0_R0_MINUS 
+ I1_0_0_1_0_0_R0_PLUS I1_0_0_1_1_0_R0_MINUS I1_0_0_1_1_0_R0_PLUS 
+ I1_0_0_2_0_0_R0_MINUS I1_0_0_2_0_0_R0_PLUS I1_0_0_2_1_0_R0_MINUS 
+ I1_0_0_2_1_0_R0_PLUS I1_0_1_0_0_0_R0_MINUS I1_0_1_0_0_0_R0_PLUS 
+ I1_0_1_0_1_0_R0_MINUS I1_0_1_0_1_0_R0_PLUS I1_0_1_1_0_0_R0_MINUS 
+ I1_0_1_1_0_0_R0_PLUS I1_0_1_1_1_0_R0_MINUS I1_0_1_1_1_0_R0_PLUS 
+ I1_0_1_2_0_0_R0_MINUS I1_0_1_2_0_0_R0_PLUS I1_0_1_2_1_0_R0_MINUS 
+ I1_0_1_2_1_0_R0_PLUS I1_0_2_0_0_0_R0_MINUS I1_0_2_0_0_0_R0_PLUS 
+ I1_0_2_0_1_0_R0_MINUS I1_0_2_0_1_0_R0_PLUS I1_0_2_1_0_0_R0_MINUS 
+ I1_0_2_1_0_0_R0_PLUS I1_0_2_1_1_0_R0_MINUS I1_0_2_1_1_0_R0_PLUS 
+ I1_0_2_2_0_0_R0_MINUS I1_0_2_2_0_0_R0_PLUS I1_0_2_2_1_0_R0_MINUS 
+ I1_0_2_2_1_0_R0_PLUS I1_1_0_0_0_0_R0_MINUS I1_1_0_0_0_0_R0_PLUS 
+ I1_1_0_0_1_0_R0_MINUS I1_1_0_0_1_0_R0_PLUS I1_1_0_1_0_0_R0_MINUS 
+ I1_1_0_1_0_0_R0_PLUS I1_1_0_1_1_0_R0_MINUS I1_1_0_1_1_0_R0_PLUS 
+ I1_1_0_2_0_0_R0_MINUS I1_1_0_2_0_0_R0_PLUS I1_1_0_2_1_0_R0_MINUS 
+ I1_1_0_2_1_0_R0_PLUS I1_1_1_0_0_0_R0_MINUS I1_1_1_0_0_0_R0_PLUS 
+ I1_1_1_0_1_0_R0_MINUS I1_1_1_0_1_0_R0_PLUS I1_1_1_1_0_0_R0_MINUS 
+ I1_1_1_1_0_0_R0_PLUS I1_1_1_1_1_0_R0_MINUS I1_1_1_1_1_0_R0_PLUS 
+ I1_1_1_2_0_0_R0_MINUS I1_1_1_2_0_0_R0_PLUS I1_1_1_2_1_0_R0_MINUS 
+ I1_1_1_2_1_0_R0_PLUS I1_1_2_0_0_0_R0_MINUS I1_1_2_0_0_0_R0_PLUS 
+ I1_1_2_0_1_0_R0_MINUS I1_1_2_0_1_0_R0_PLUS I1_1_2_1_0_0_R0_MINUS 
+ I1_1_2_1_0_0_R0_PLUS I1_1_2_1_1_0_R0_MINUS I1_1_2_1_1_0_R0_PLUS 
+ I1_1_2_2_0_0_R0_MINUS I1_1_2_2_0_0_R0_PLUS I1_1_2_2_1_0_R0_MINUS 
+ I1_1_2_2_1_0_R0_PLUS I1_2_0_0_0_0_R0_MINUS I1_2_0_0_0_0_R0_PLUS 
+ I1_2_0_0_1_0_R0_MINUS I1_2_0_0_1_0_R0_PLUS I1_2_0_1_0_0_R0_MINUS 
+ I1_2_0_1_0_0_R0_PLUS I1_2_0_1_1_0_R0_MINUS I1_2_0_1_1_0_R0_PLUS 
+ I1_2_0_2_0_0_R0_MINUS I1_2_0_2_0_0_R0_PLUS I1_2_0_2_1_0_R0_MINUS 
+ I1_2_0_2_1_0_R0_PLUS I1_2_1_0_0_0_R0_MINUS I1_2_1_0_0_0_R0_PLUS 
+ I1_2_1_0_1_0_R0_MINUS I1_2_1_0_1_0_R0_PLUS I1_2_1_1_0_0_R0_MINUS 
+ I1_2_1_1_0_0_R0_PLUS I1_2_1_1_1_0_R0_MINUS I1_2_1_1_1_0_R0_PLUS 
+ I1_2_1_2_0_0_R0_MINUS I1_2_1_2_0_0_R0_PLUS I1_2_1_2_1_0_R0_MINUS 
+ I1_2_1_2_1_0_R0_PLUS I1_2_2_0_0_0_R0_MINUS I1_2_2_0_0_0_R0_PLUS 
+ I1_2_2_0_1_0_R0_MINUS I1_2_2_0_1_0_R0_PLUS I1_2_2_1_0_0_R0_MINUS 
+ I1_2_2_1_0_0_R0_PLUS I1_2_2_1_1_0_R0_MINUS I1_2_2_1_1_0_R0_PLUS 
+ I1_2_2_2_0_0_R0_MINUS I1_2_2_2_0_0_R0_PLUS I1_2_2_2_1_0_R0_MINUS 
+ I1_2_2_2_1_0_R0_PLUS I1_default_MINUS I1_default_PLUS gnd!
*.PININFO I1_0_0_0_0_0_R0_MINUS:I I1_0_0_0_0_0_R0_PLUS:I 
*.PININFO I1_0_0_0_1_0_R0_MINUS:I I1_0_0_0_1_0_R0_PLUS:I 
*.PININFO I1_0_0_1_0_0_R0_MINUS:I I1_0_0_1_0_0_R0_PLUS:I 
*.PININFO I1_0_0_1_1_0_R0_MINUS:I I1_0_0_1_1_0_R0_PLUS:I 
*.PININFO I1_0_0_2_0_0_R0_MINUS:I I1_0_0_2_0_0_R0_PLUS:I 
*.PININFO I1_0_0_2_1_0_R0_MINUS:I I1_0_0_2_1_0_R0_PLUS:I 
*.PININFO I1_0_1_0_0_0_R0_MINUS:I I1_0_1_0_0_0_R0_PLUS:I 
*.PININFO I1_0_1_0_1_0_R0_MINUS:I I1_0_1_0_1_0_R0_PLUS:I 
*.PININFO I1_0_1_1_0_0_R0_MINUS:I I1_0_1_1_0_0_R0_PLUS:I 
*.PININFO I1_0_1_1_1_0_R0_MINUS:I I1_0_1_1_1_0_R0_PLUS:I 
*.PININFO I1_0_1_2_0_0_R0_MINUS:I I1_0_1_2_0_0_R0_PLUS:I 
*.PININFO I1_0_1_2_1_0_R0_MINUS:I I1_0_1_2_1_0_R0_PLUS:I 
*.PININFO I1_0_2_0_0_0_R0_MINUS:I I1_0_2_0_0_0_R0_PLUS:I 
*.PININFO I1_0_2_0_1_0_R0_MINUS:I I1_0_2_0_1_0_R0_PLUS:I 
*.PININFO I1_0_2_1_0_0_R0_MINUS:I I1_0_2_1_0_0_R0_PLUS:I 
*.PININFO I1_0_2_1_1_0_R0_MINUS:I I1_0_2_1_1_0_R0_PLUS:I 
*.PININFO I1_0_2_2_0_0_R0_MINUS:I I1_0_2_2_0_0_R0_PLUS:I 
*.PININFO I1_0_2_2_1_0_R0_MINUS:I I1_0_2_2_1_0_R0_PLUS:I 
*.PININFO I1_1_0_0_0_0_R0_MINUS:I I1_1_0_0_0_0_R0_PLUS:I 
*.PININFO I1_1_0_0_1_0_R0_MINUS:I I1_1_0_0_1_0_R0_PLUS:I 
*.PININFO I1_1_0_1_0_0_R0_MINUS:I I1_1_0_1_0_0_R0_PLUS:I 
*.PININFO I1_1_0_1_1_0_R0_MINUS:I I1_1_0_1_1_0_R0_PLUS:I 
*.PININFO I1_1_0_2_0_0_R0_MINUS:I I1_1_0_2_0_0_R0_PLUS:I 
*.PININFO I1_1_0_2_1_0_R0_MINUS:I I1_1_0_2_1_0_R0_PLUS:I 
*.PININFO I1_1_1_0_0_0_R0_MINUS:I I1_1_1_0_0_0_R0_PLUS:I 
*.PININFO I1_1_1_0_1_0_R0_MINUS:I I1_1_1_0_1_0_R0_PLUS:I 
*.PININFO I1_1_1_1_0_0_R0_MINUS:I I1_1_1_1_0_0_R0_PLUS:I 
*.PININFO I1_1_1_1_1_0_R0_MINUS:I I1_1_1_1_1_0_R0_PLUS:I 
*.PININFO I1_1_1_2_0_0_R0_MINUS:I I1_1_1_2_0_0_R0_PLUS:I 
*.PININFO I1_1_1_2_1_0_R0_MINUS:I I1_1_1_2_1_0_R0_PLUS:I 
*.PININFO I1_1_2_0_0_0_R0_MINUS:I I1_1_2_0_0_0_R0_PLUS:I 
*.PININFO I1_1_2_0_1_0_R0_MINUS:I I1_1_2_0_1_0_R0_PLUS:I 
*.PININFO I1_1_2_1_0_0_R0_MINUS:I I1_1_2_1_0_0_R0_PLUS:I 
*.PININFO I1_1_2_1_1_0_R0_MINUS:I I1_1_2_1_1_0_R0_PLUS:I 
*.PININFO I1_1_2_2_0_0_R0_MINUS:I I1_1_2_2_0_0_R0_PLUS:I 
*.PININFO I1_1_2_2_1_0_R0_MINUS:I I1_1_2_2_1_0_R0_PLUS:I 
*.PININFO I1_2_0_0_0_0_R0_MINUS:I I1_2_0_0_0_0_R0_PLUS:I 
*.PININFO I1_2_0_0_1_0_R0_MINUS:I I1_2_0_0_1_0_R0_PLUS:I 
*.PININFO I1_2_0_1_0_0_R0_MINUS:I I1_2_0_1_0_0_R0_PLUS:I 
*.PININFO I1_2_0_1_1_0_R0_MINUS:I I1_2_0_1_1_0_R0_PLUS:I 
*.PININFO I1_2_0_2_0_0_R0_MINUS:I I1_2_0_2_0_0_R0_PLUS:I 
*.PININFO I1_2_0_2_1_0_R0_MINUS:I I1_2_0_2_1_0_R0_PLUS:I 
*.PININFO I1_2_1_0_0_0_R0_MINUS:I I1_2_1_0_0_0_R0_PLUS:I 
*.PININFO I1_2_1_0_1_0_R0_MINUS:I I1_2_1_0_1_0_R0_PLUS:I 
*.PININFO I1_2_1_1_0_0_R0_MINUS:I I1_2_1_1_0_0_R0_PLUS:I 
*.PININFO I1_2_1_1_1_0_R0_MINUS:I I1_2_1_1_1_0_R0_PLUS:I 
*.PININFO I1_2_1_2_0_0_R0_MINUS:I I1_2_1_2_0_0_R0_PLUS:I 
*.PININFO I1_2_1_2_1_0_R0_MINUS:I I1_2_1_2_1_0_R0_PLUS:I 
*.PININFO I1_2_2_0_0_0_R0_MINUS:I I1_2_2_0_0_0_R0_PLUS:I 
*.PININFO I1_2_2_0_1_0_R0_MINUS:I I1_2_2_0_1_0_R0_PLUS:I 
*.PININFO I1_2_2_1_0_0_R0_MINUS:I I1_2_2_1_0_0_R0_PLUS:I 
*.PININFO I1_2_2_1_1_0_R0_MINUS:I I1_2_2_1_1_0_R0_PLUS:I 
*.PININFO I1_2_2_2_0_0_R0_MINUS:I I1_2_2_2_0_0_R0_PLUS:I 
*.PININFO I1_2_2_2_1_0_R0_MINUS:I I1_2_2_2_1_0_R0_PLUS:I I1_default_MINUS:I 
*.PININFO I1_default_PLUS:I gnd!:I
RI1_2_2_2_1_0_R0 I1_2_2_2_1_0_R0_PLUS I1_2_2_2_1_0_R0_MINUS gnd! 
+ nplus_u m=8.0 l=50u w=50u r=60.6187 par=8.0 s=1
RI1_2_2_2_0_0_R0 I1_2_2_2_0_0_R0_PLUS I1_2_2_2_0_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=50u w=50u r=60.6187 par=1.0 s=8
RI1_2_2_1_1_0_R0 I1_2_2_1_1_0_R0_PLUS I1_2_2_1_1_0_R0_MINUS gnd! 
+ nplus_u m=3.0 l=50u w=50u r=60.6187 par=3.0 s=1
RI1_2_2_1_0_0_R0 I1_2_2_1_0_0_R0_PLUS I1_2_2_1_0_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=50u w=50u r=60.6187 par=1.0 s=3
RI1_2_2_0_1_0_R0 I1_2_2_0_1_0_R0_PLUS I1_2_2_0_1_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=50u w=50u r=60.6187 par=1.0 s=1
RI1_2_2_0_0_0_R0 I1_2_2_0_0_0_R0_PLUS I1_2_2_0_0_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=50u w=50u r=60.6187 par=1.0 s=1
RI1_2_1_2_1_0_R0 I1_2_1_2_1_0_R0_PLUS I1_2_1_2_1_0_R0_MINUS gnd! 
+ nplus_u m=8.0 l=7.6u w=50u r=9.84027 par=8.0 s=1
RI1_2_1_2_0_0_R0 I1_2_1_2_0_0_R0_PLUS I1_2_1_2_0_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=7.6u w=50u r=9.84027 par=1.0 s=8
RI1_2_1_1_1_0_R0 I1_2_1_1_1_0_R0_PLUS I1_2_1_1_1_0_R0_MINUS gnd! 
+ nplus_u m=3.0 l=7.6u w=50u r=9.84027 par=3.0 s=1
RI1_2_1_1_0_0_R0 I1_2_1_1_0_0_R0_PLUS I1_2_1_1_0_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=7.6u w=50u r=9.84027 par=1.0 s=3
RI1_2_1_0_1_0_R0 I1_2_1_0_1_0_R0_PLUS I1_2_1_0_1_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=7.6u w=50u r=9.84027 par=1.0 s=1
RI1_2_1_0_0_0_R0 I1_2_1_0_0_0_R0_PLUS I1_2_1_0_0_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=7.6u w=50u r=9.84027 par=1.0 s=1
RI1_2_0_2_1_0_R0 I1_2_0_2_1_0_R0_PLUS I1_2_0_2_1_0_R0_MINUS gnd! 
+ nplus_u m=8.0 l=1.6u w=50u r=2.65464 par=8.0 s=1
RI1_2_0_2_0_0_R0 I1_2_0_2_0_0_R0_PLUS I1_2_0_2_0_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=1.6u w=50u r=2.65464 par=1.0 s=8
RI1_2_0_1_1_0_R0 I1_2_0_1_1_0_R0_PLUS I1_2_0_1_1_0_R0_MINUS gnd! 
+ nplus_u m=3.0 l=1.6u w=50u r=2.65464 par=3.0 s=1
RI1_2_0_1_0_0_R0 I1_2_0_1_0_0_R0_PLUS I1_2_0_1_0_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=1.6u w=50u r=2.65464 par=1.0 s=3
RI1_2_0_0_1_0_R0 I1_2_0_0_1_0_R0_PLUS I1_2_0_0_1_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=1.6u w=50u r=2.65464 par=1.0 s=1
RI1_2_0_0_0_0_R0 I1_2_0_0_0_0_R0_PLUS I1_2_0_0_0_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=1.6u w=50u r=2.65464 par=1.0 s=1
RI1_1_2_2_1_0_R0 I1_1_2_2_1_0_R0_PLUS I1_1_2_2_1_0_R0_MINUS gnd! 
+ nplus_u m=8.0 l=50u w=3.62u r=816.397 par=8.0 s=1
RI1_1_2_2_0_0_R0 I1_1_2_2_0_0_R0_PLUS I1_1_2_2_0_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=50u w=3.62u r=816.397 par=1.0 s=8
RI1_1_2_1_1_0_R0 I1_1_2_1_1_0_R0_PLUS I1_1_2_1_1_0_R0_MINUS gnd! 
+ nplus_u m=3.0 l=50u w=3.62u r=816.397 par=3.0 s=1
RI1_1_2_1_0_0_R0 I1_1_2_1_0_0_R0_PLUS I1_1_2_1_0_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=50u w=3.62u r=816.397 par=1.0 s=3
RI1_1_2_0_1_0_R0 I1_1_2_0_1_0_R0_PLUS I1_1_2_0_1_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=50u w=3.62u r=816.397 par=1.0 s=1
RI1_1_2_0_0_0_R0 I1_1_2_0_0_0_R0_PLUS I1_1_2_0_0_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=50u w=3.62u r=816.397 par=1.0 s=1
RI1_1_1_2_1_0_R0 I1_1_1_2_1_0_R0_PLUS I1_1_1_2_1_0_R0_MINUS gnd! 
+ nplus_u m=8.0 l=7.6u w=3.62u r=132.526 par=8.0 s=1
RI1_1_1_2_0_0_R0 I1_1_1_2_0_0_R0_PLUS I1_1_1_2_0_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=7.6u w=3.62u r=132.526 par=1.0 s=8
RI1_1_1_1_1_0_R0 I1_1_1_1_1_0_R0_PLUS I1_1_1_1_1_0_R0_MINUS gnd! 
+ nplus_u m=3.0 l=7.6u w=3.62u r=132.526 par=3.0 s=1
RI1_1_1_1_0_0_R0 I1_1_1_1_0_0_R0_PLUS I1_1_1_1_0_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=7.6u w=3.62u r=132.526 par=1.0 s=3
RI1_1_1_0_1_0_R0 I1_1_1_0_1_0_R0_PLUS I1_1_1_0_1_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=7.6u w=3.62u r=132.526 par=1.0 s=1
RI1_1_1_0_0_0_R0 I1_1_1_0_0_0_R0_PLUS I1_1_1_0_0_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=7.6u w=3.62u r=132.526 par=1.0 s=1
RI1_1_0_2_1_0_R0 I1_1_0_2_1_0_R0_PLUS I1_1_0_2_1_0_R0_MINUS gnd! 
+ nplus_u m=8.0 l=1.6u w=3.62u r=35.752 par=8.0 s=1
RI1_1_0_2_0_0_R0 I1_1_0_2_0_0_R0_PLUS I1_1_0_2_0_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=1.6u w=3.62u r=35.752 par=1.0 s=8
RI1_1_0_1_1_0_R0 I1_1_0_1_1_0_R0_PLUS I1_1_0_1_1_0_R0_MINUS gnd! 
+ nplus_u m=3.0 l=1.6u w=3.62u r=35.752 par=3.0 s=1
RI1_1_0_1_0_0_R0 I1_1_0_1_0_0_R0_PLUS I1_1_0_1_0_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=1.6u w=3.62u r=35.752 par=1.0 s=3
RI1_1_0_0_1_0_R0 I1_1_0_0_1_0_R0_PLUS I1_1_0_0_1_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=1.6u w=3.62u r=35.752 par=1.0 s=1
RI1_1_0_0_0_0_R0 I1_1_0_0_0_0_R0_PLUS I1_1_0_0_0_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=1.6u w=3.62u r=35.752 par=1.0 s=1
RI1_0_2_2_1_0_R0 I1_0_2_2_1_0_R0_PLUS I1_0_2_2_1_0_R0_MINUS gnd! 
+ nplus_u m=8.0 l=50u w=800n r=3.37444K par=8.0 s=1
RI1_0_2_2_0_0_R0 I1_0_2_2_0_0_R0_PLUS I1_0_2_2_0_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=50u w=800n r=3.37444K par=1.0 s=8
RI1_0_2_1_1_0_R0 I1_0_2_1_1_0_R0_PLUS I1_0_2_1_1_0_R0_MINUS gnd! 
+ nplus_u m=3.0 l=50u w=800n r=3.37444K par=3.0 s=1
RI1_0_2_1_0_0_R0 I1_0_2_1_0_0_R0_PLUS I1_0_2_1_0_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=50u w=800n r=3.37444K par=1.0 s=3
RI1_0_2_0_1_0_R0 I1_0_2_0_1_0_R0_PLUS I1_0_2_0_1_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=50u w=800n r=3.37444K par=1.0 s=1
RI1_0_2_0_0_0_R0 I1_0_2_0_0_0_R0_PLUS I1_0_2_0_0_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=50u w=800n r=3.37444K par=1.0 s=1
RI1_0_1_2_1_0_R0 I1_0_1_2_1_0_R0_PLUS I1_0_1_2_1_0_R0_MINUS gnd! 
+ nplus_u m=8.0 l=7.6u w=800n r=547.775 par=8.0 s=1
RI1_0_1_2_0_0_R0 I1_0_1_2_0_0_R0_PLUS I1_0_1_2_0_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=7.6u w=800n r=547.775 par=1.0 s=8
RI1_0_1_1_1_0_R0 I1_0_1_1_1_0_R0_PLUS I1_0_1_1_1_0_R0_MINUS gnd! 
+ nplus_u m=3.0 l=7.6u w=800n r=547.775 par=3.0 s=1
RI1_0_1_1_0_0_R0 I1_0_1_1_0_0_R0_PLUS I1_0_1_1_0_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=7.6u w=800n r=547.775 par=1.0 s=3
RI1_0_1_0_1_0_R0 I1_0_1_0_1_0_R0_PLUS I1_0_1_0_1_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=7.6u w=800n r=547.775 par=1.0 s=1
RI1_0_1_0_0_0_R0 I1_0_1_0_0_0_R0_PLUS I1_0_1_0_0_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=7.6u w=800n r=547.775 par=1.0 s=1
RI1_0_0_2_1_0_R0 I1_0_0_2_1_0_R0_PLUS I1_0_0_2_1_0_R0_MINUS gnd! 
+ nplus_u m=8.0 l=1.6u w=800n r=147.775 par=8.0 s=1
RI1_0_0_2_0_0_R0 I1_0_0_2_0_0_R0_PLUS I1_0_0_2_0_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=1.6u w=800n r=147.775 par=1.0 s=8
RI1_0_0_1_1_0_R0 I1_0_0_1_1_0_R0_PLUS I1_0_0_1_1_0_R0_MINUS gnd! 
+ nplus_u m=3.0 l=1.6u w=800n r=147.775 par=3.0 s=1
RI1_0_0_1_0_0_R0 I1_0_0_1_0_0_R0_PLUS I1_0_0_1_0_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=1.6u w=800n r=147.775 par=1.0 s=3
RI1_0_0_0_1_0_R0 I1_0_0_0_1_0_R0_PLUS I1_0_0_0_1_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=1.6u w=800n r=147.775 par=1.0 s=1
RI1_0_0_0_0_0_R0 I1_0_0_0_0_0_R0_PLUS I1_0_0_0_0_0_R0_MINUS gnd! 
+ nplus_u m=1.0 l=1.6u w=800n r=147.775 par=1.0 s=1
RI1_default I1_default_PLUS I1_default_MINUS gnd! nplus_u m=1.0 l=2u 
+ w=1u r=142.7251 par=1.0 s=1
.ENDS

