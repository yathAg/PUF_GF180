magic
tech gf180mcuA
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -51 24849 13013 25405
rect -51 505 505 24849
rect 12457 505 13013 24849
rect -51 -51 13013 505
<< mvnmos >>
rect 1481 23733 11481 23873
rect 1481 23489 11481 23629
rect 1481 23245 11481 23385
rect 1481 23001 11481 23141
rect 1481 22757 11481 22897
rect 1481 22513 11481 22653
rect 1481 22269 11481 22409
rect 1481 22025 11481 22165
rect 1481 21781 11481 21921
rect 1481 21537 11481 21677
rect 1481 21293 11481 21433
rect 1481 21049 11481 21189
rect 1481 20805 11481 20945
rect 1481 20561 11481 20701
rect 1481 20317 11481 20457
rect 1481 20073 11481 20213
rect 1481 19829 11481 19969
rect 1481 19585 11481 19725
rect 1481 19341 11481 19481
rect 1481 19097 11481 19237
rect 1481 17861 11481 18001
rect 1481 17617 11481 17757
rect 1481 17373 11481 17513
rect 1481 17129 11481 17269
rect 1481 16885 11481 17025
rect 1481 16641 11481 16781
rect 1481 16397 11481 16537
rect 1481 16153 11481 16293
rect 1481 15909 11481 16049
rect 1481 15665 11481 15805
rect 1481 15421 11481 15561
rect 1481 15177 11481 15317
rect 1481 14933 11481 15073
rect 1481 14689 11481 14829
rect 1481 14445 11481 14585
rect 1481 14201 11481 14341
rect 1481 13957 11481 14097
rect 1481 13713 11481 13853
rect 1481 13469 11481 13609
rect 1481 13225 11481 13365
rect 1481 11989 11481 12129
rect 1481 11745 11481 11885
rect 1481 11501 11481 11641
rect 1481 11257 11481 11397
rect 1481 11013 11481 11153
rect 1481 10769 11481 10909
rect 1481 10525 11481 10665
rect 1481 10281 11481 10421
rect 1481 10037 11481 10177
rect 1481 9793 11481 9933
rect 1481 9549 11481 9689
rect 1481 9305 11481 9445
rect 1481 9061 11481 9201
rect 1481 8817 11481 8957
rect 1481 8573 11481 8713
rect 1481 8329 11481 8469
rect 1481 8085 11481 8225
rect 1481 7841 11481 7981
rect 1481 7597 11481 7737
rect 1481 7353 11481 7493
rect 1481 6117 11481 6257
rect 1481 5873 11481 6013
rect 1481 5629 11481 5769
rect 1481 5385 11481 5525
rect 1481 5141 11481 5281
rect 1481 4897 11481 5037
rect 1481 4653 11481 4793
rect 1481 4409 11481 4549
rect 1481 4165 11481 4305
rect 1481 3921 11481 4061
rect 1481 3677 11481 3817
rect 1481 3433 11481 3573
rect 1481 3189 11481 3329
rect 1481 2945 11481 3085
rect 1481 2701 11481 2841
rect 1481 2457 11481 2597
rect 1481 2213 11481 2353
rect 1481 1969 11481 2109
rect 1481 1725 11481 1865
rect 1481 1481 11481 1621
<< mvndiff >>
rect 1481 23948 11481 23961
rect 1481 23902 1494 23948
rect 11468 23902 11481 23948
rect 1481 23873 11481 23902
rect 1481 23704 11481 23733
rect 1481 23658 1494 23704
rect 11468 23658 11481 23704
rect 1481 23629 11481 23658
rect 1481 23460 11481 23489
rect 1481 23414 1494 23460
rect 11468 23414 11481 23460
rect 1481 23385 11481 23414
rect 1481 23216 11481 23245
rect 1481 23170 1494 23216
rect 11468 23170 11481 23216
rect 1481 23141 11481 23170
rect 1481 22972 11481 23001
rect 1481 22926 1494 22972
rect 11468 22926 11481 22972
rect 1481 22897 11481 22926
rect 1481 22728 11481 22757
rect 1481 22682 1494 22728
rect 11468 22682 11481 22728
rect 1481 22653 11481 22682
rect 1481 22484 11481 22513
rect 1481 22438 1494 22484
rect 11468 22438 11481 22484
rect 1481 22409 11481 22438
rect 1481 22240 11481 22269
rect 1481 22194 1494 22240
rect 11468 22194 11481 22240
rect 1481 22165 11481 22194
rect 1481 21996 11481 22025
rect 1481 21950 1494 21996
rect 11468 21950 11481 21996
rect 1481 21921 11481 21950
rect 1481 21752 11481 21781
rect 1481 21706 1494 21752
rect 11468 21706 11481 21752
rect 1481 21677 11481 21706
rect 1481 21508 11481 21537
rect 1481 21462 1494 21508
rect 11468 21462 11481 21508
rect 1481 21433 11481 21462
rect 1481 21264 11481 21293
rect 1481 21218 1494 21264
rect 11468 21218 11481 21264
rect 1481 21189 11481 21218
rect 1481 21020 11481 21049
rect 1481 20974 1494 21020
rect 11468 20974 11481 21020
rect 1481 20945 11481 20974
rect 1481 20776 11481 20805
rect 1481 20730 1494 20776
rect 11468 20730 11481 20776
rect 1481 20701 11481 20730
rect 1481 20532 11481 20561
rect 1481 20486 1494 20532
rect 11468 20486 11481 20532
rect 1481 20457 11481 20486
rect 1481 20288 11481 20317
rect 1481 20242 1494 20288
rect 11468 20242 11481 20288
rect 1481 20213 11481 20242
rect 1481 20044 11481 20073
rect 1481 19998 1494 20044
rect 11468 19998 11481 20044
rect 1481 19969 11481 19998
rect 1481 19800 11481 19829
rect 1481 19754 1494 19800
rect 11468 19754 11481 19800
rect 1481 19725 11481 19754
rect 1481 19556 11481 19585
rect 1481 19510 1494 19556
rect 11468 19510 11481 19556
rect 1481 19481 11481 19510
rect 1481 19312 11481 19341
rect 1481 19266 1494 19312
rect 11468 19266 11481 19312
rect 1481 19237 11481 19266
rect 1481 19068 11481 19097
rect 1481 19022 1494 19068
rect 11468 19022 11481 19068
rect 1481 19009 11481 19022
rect 1481 18076 11481 18089
rect 1481 18030 1494 18076
rect 11468 18030 11481 18076
rect 1481 18001 11481 18030
rect 1481 17832 11481 17861
rect 1481 17786 1494 17832
rect 11468 17786 11481 17832
rect 1481 17757 11481 17786
rect 1481 17588 11481 17617
rect 1481 17542 1494 17588
rect 11468 17542 11481 17588
rect 1481 17513 11481 17542
rect 1481 17344 11481 17373
rect 1481 17298 1494 17344
rect 11468 17298 11481 17344
rect 1481 17269 11481 17298
rect 1481 17100 11481 17129
rect 1481 17054 1494 17100
rect 11468 17054 11481 17100
rect 1481 17025 11481 17054
rect 1481 16856 11481 16885
rect 1481 16810 1494 16856
rect 11468 16810 11481 16856
rect 1481 16781 11481 16810
rect 1481 16612 11481 16641
rect 1481 16566 1494 16612
rect 11468 16566 11481 16612
rect 1481 16537 11481 16566
rect 1481 16368 11481 16397
rect 1481 16322 1494 16368
rect 11468 16322 11481 16368
rect 1481 16293 11481 16322
rect 1481 16124 11481 16153
rect 1481 16078 1494 16124
rect 11468 16078 11481 16124
rect 1481 16049 11481 16078
rect 1481 15880 11481 15909
rect 1481 15834 1494 15880
rect 11468 15834 11481 15880
rect 1481 15805 11481 15834
rect 1481 15636 11481 15665
rect 1481 15590 1494 15636
rect 11468 15590 11481 15636
rect 1481 15561 11481 15590
rect 1481 15392 11481 15421
rect 1481 15346 1494 15392
rect 11468 15346 11481 15392
rect 1481 15317 11481 15346
rect 1481 15148 11481 15177
rect 1481 15102 1494 15148
rect 11468 15102 11481 15148
rect 1481 15073 11481 15102
rect 1481 14904 11481 14933
rect 1481 14858 1494 14904
rect 11468 14858 11481 14904
rect 1481 14829 11481 14858
rect 1481 14660 11481 14689
rect 1481 14614 1494 14660
rect 11468 14614 11481 14660
rect 1481 14585 11481 14614
rect 1481 14416 11481 14445
rect 1481 14370 1494 14416
rect 11468 14370 11481 14416
rect 1481 14341 11481 14370
rect 1481 14172 11481 14201
rect 1481 14126 1494 14172
rect 11468 14126 11481 14172
rect 1481 14097 11481 14126
rect 1481 13928 11481 13957
rect 1481 13882 1494 13928
rect 11468 13882 11481 13928
rect 1481 13853 11481 13882
rect 1481 13684 11481 13713
rect 1481 13638 1494 13684
rect 11468 13638 11481 13684
rect 1481 13609 11481 13638
rect 1481 13440 11481 13469
rect 1481 13394 1494 13440
rect 11468 13394 11481 13440
rect 1481 13365 11481 13394
rect 1481 13196 11481 13225
rect 1481 13150 1494 13196
rect 11468 13150 11481 13196
rect 1481 13137 11481 13150
rect 1481 12204 11481 12217
rect 1481 12158 1494 12204
rect 11468 12158 11481 12204
rect 1481 12129 11481 12158
rect 1481 11960 11481 11989
rect 1481 11914 1494 11960
rect 11468 11914 11481 11960
rect 1481 11885 11481 11914
rect 1481 11716 11481 11745
rect 1481 11670 1494 11716
rect 11468 11670 11481 11716
rect 1481 11641 11481 11670
rect 1481 11472 11481 11501
rect 1481 11426 1494 11472
rect 11468 11426 11481 11472
rect 1481 11397 11481 11426
rect 1481 11228 11481 11257
rect 1481 11182 1494 11228
rect 11468 11182 11481 11228
rect 1481 11153 11481 11182
rect 1481 10984 11481 11013
rect 1481 10938 1494 10984
rect 11468 10938 11481 10984
rect 1481 10909 11481 10938
rect 1481 10740 11481 10769
rect 1481 10694 1494 10740
rect 11468 10694 11481 10740
rect 1481 10665 11481 10694
rect 1481 10496 11481 10525
rect 1481 10450 1494 10496
rect 11468 10450 11481 10496
rect 1481 10421 11481 10450
rect 1481 10252 11481 10281
rect 1481 10206 1494 10252
rect 11468 10206 11481 10252
rect 1481 10177 11481 10206
rect 1481 10008 11481 10037
rect 1481 9962 1494 10008
rect 11468 9962 11481 10008
rect 1481 9933 11481 9962
rect 1481 9764 11481 9793
rect 1481 9718 1494 9764
rect 11468 9718 11481 9764
rect 1481 9689 11481 9718
rect 1481 9520 11481 9549
rect 1481 9474 1494 9520
rect 11468 9474 11481 9520
rect 1481 9445 11481 9474
rect 1481 9276 11481 9305
rect 1481 9230 1494 9276
rect 11468 9230 11481 9276
rect 1481 9201 11481 9230
rect 1481 9032 11481 9061
rect 1481 8986 1494 9032
rect 11468 8986 11481 9032
rect 1481 8957 11481 8986
rect 1481 8788 11481 8817
rect 1481 8742 1494 8788
rect 11468 8742 11481 8788
rect 1481 8713 11481 8742
rect 1481 8544 11481 8573
rect 1481 8498 1494 8544
rect 11468 8498 11481 8544
rect 1481 8469 11481 8498
rect 1481 8300 11481 8329
rect 1481 8254 1494 8300
rect 11468 8254 11481 8300
rect 1481 8225 11481 8254
rect 1481 8056 11481 8085
rect 1481 8010 1494 8056
rect 11468 8010 11481 8056
rect 1481 7981 11481 8010
rect 1481 7812 11481 7841
rect 1481 7766 1494 7812
rect 11468 7766 11481 7812
rect 1481 7737 11481 7766
rect 1481 7568 11481 7597
rect 1481 7522 1494 7568
rect 11468 7522 11481 7568
rect 1481 7493 11481 7522
rect 1481 7324 11481 7353
rect 1481 7278 1494 7324
rect 11468 7278 11481 7324
rect 1481 7265 11481 7278
rect 1481 6332 11481 6345
rect 1481 6286 1494 6332
rect 11468 6286 11481 6332
rect 1481 6257 11481 6286
rect 1481 6088 11481 6117
rect 1481 6042 1494 6088
rect 11468 6042 11481 6088
rect 1481 6013 11481 6042
rect 1481 5844 11481 5873
rect 1481 5798 1494 5844
rect 11468 5798 11481 5844
rect 1481 5769 11481 5798
rect 1481 5600 11481 5629
rect 1481 5554 1494 5600
rect 11468 5554 11481 5600
rect 1481 5525 11481 5554
rect 1481 5356 11481 5385
rect 1481 5310 1494 5356
rect 11468 5310 11481 5356
rect 1481 5281 11481 5310
rect 1481 5112 11481 5141
rect 1481 5066 1494 5112
rect 11468 5066 11481 5112
rect 1481 5037 11481 5066
rect 1481 4868 11481 4897
rect 1481 4822 1494 4868
rect 11468 4822 11481 4868
rect 1481 4793 11481 4822
rect 1481 4624 11481 4653
rect 1481 4578 1494 4624
rect 11468 4578 11481 4624
rect 1481 4549 11481 4578
rect 1481 4380 11481 4409
rect 1481 4334 1494 4380
rect 11468 4334 11481 4380
rect 1481 4305 11481 4334
rect 1481 4136 11481 4165
rect 1481 4090 1494 4136
rect 11468 4090 11481 4136
rect 1481 4061 11481 4090
rect 1481 3892 11481 3921
rect 1481 3846 1494 3892
rect 11468 3846 11481 3892
rect 1481 3817 11481 3846
rect 1481 3648 11481 3677
rect 1481 3602 1494 3648
rect 11468 3602 11481 3648
rect 1481 3573 11481 3602
rect 1481 3404 11481 3433
rect 1481 3358 1494 3404
rect 11468 3358 11481 3404
rect 1481 3329 11481 3358
rect 1481 3160 11481 3189
rect 1481 3114 1494 3160
rect 11468 3114 11481 3160
rect 1481 3085 11481 3114
rect 1481 2916 11481 2945
rect 1481 2870 1494 2916
rect 11468 2870 11481 2916
rect 1481 2841 11481 2870
rect 1481 2672 11481 2701
rect 1481 2626 1494 2672
rect 11468 2626 11481 2672
rect 1481 2597 11481 2626
rect 1481 2428 11481 2457
rect 1481 2382 1494 2428
rect 11468 2382 11481 2428
rect 1481 2353 11481 2382
rect 1481 2184 11481 2213
rect 1481 2138 1494 2184
rect 11468 2138 11481 2184
rect 1481 2109 11481 2138
rect 1481 1940 11481 1969
rect 1481 1894 1494 1940
rect 11468 1894 11481 1940
rect 1481 1865 11481 1894
rect 1481 1696 11481 1725
rect 1481 1650 1494 1696
rect 11468 1650 11481 1696
rect 1481 1621 11481 1650
rect 1481 1452 11481 1481
rect 1481 1406 1494 1452
rect 11468 1406 11481 1452
rect 1481 1393 11481 1406
<< mvndiffc >>
rect 1494 23902 11468 23948
rect 1494 23658 11468 23704
rect 1494 23414 11468 23460
rect 1494 23170 11468 23216
rect 1494 22926 11468 22972
rect 1494 22682 11468 22728
rect 1494 22438 11468 22484
rect 1494 22194 11468 22240
rect 1494 21950 11468 21996
rect 1494 21706 11468 21752
rect 1494 21462 11468 21508
rect 1494 21218 11468 21264
rect 1494 20974 11468 21020
rect 1494 20730 11468 20776
rect 1494 20486 11468 20532
rect 1494 20242 11468 20288
rect 1494 19998 11468 20044
rect 1494 19754 11468 19800
rect 1494 19510 11468 19556
rect 1494 19266 11468 19312
rect 1494 19022 11468 19068
rect 1494 18030 11468 18076
rect 1494 17786 11468 17832
rect 1494 17542 11468 17588
rect 1494 17298 11468 17344
rect 1494 17054 11468 17100
rect 1494 16810 11468 16856
rect 1494 16566 11468 16612
rect 1494 16322 11468 16368
rect 1494 16078 11468 16124
rect 1494 15834 11468 15880
rect 1494 15590 11468 15636
rect 1494 15346 11468 15392
rect 1494 15102 11468 15148
rect 1494 14858 11468 14904
rect 1494 14614 11468 14660
rect 1494 14370 11468 14416
rect 1494 14126 11468 14172
rect 1494 13882 11468 13928
rect 1494 13638 11468 13684
rect 1494 13394 11468 13440
rect 1494 13150 11468 13196
rect 1494 12158 11468 12204
rect 1494 11914 11468 11960
rect 1494 11670 11468 11716
rect 1494 11426 11468 11472
rect 1494 11182 11468 11228
rect 1494 10938 11468 10984
rect 1494 10694 11468 10740
rect 1494 10450 11468 10496
rect 1494 10206 11468 10252
rect 1494 9962 11468 10008
rect 1494 9718 11468 9764
rect 1494 9474 11468 9520
rect 1494 9230 11468 9276
rect 1494 8986 11468 9032
rect 1494 8742 11468 8788
rect 1494 8498 11468 8544
rect 1494 8254 11468 8300
rect 1494 8010 11468 8056
rect 1494 7766 11468 7812
rect 1494 7522 11468 7568
rect 1494 7278 11468 7324
rect 1494 6286 11468 6332
rect 1494 6042 11468 6088
rect 1494 5798 11468 5844
rect 1494 5554 11468 5600
rect 1494 5310 11468 5356
rect 1494 5066 11468 5112
rect 1494 4822 11468 4868
rect 1494 4578 11468 4624
rect 1494 4334 11468 4380
rect 1494 4090 11468 4136
rect 1494 3846 11468 3892
rect 1494 3602 11468 3648
rect 1494 3358 11468 3404
rect 1494 3114 11468 3160
rect 1494 2870 11468 2916
rect 1494 2626 11468 2672
rect 1494 2382 11468 2428
rect 1494 2138 11468 2184
rect 1494 1894 11468 1940
rect 1494 1650 11468 1696
rect 1494 1406 11468 1452
<< psubdiff >>
rect 582 24700 12380 24722
rect 582 654 604 24700
rect 950 24354 1058 24700
rect 11904 24354 12012 24700
rect 950 24332 12012 24354
rect 950 18644 972 24332
rect 11990 18644 12012 24332
rect 950 18622 12012 18644
rect 950 18476 1058 18622
rect 11904 18476 12012 18622
rect 950 18454 12012 18476
rect 950 12772 972 18454
rect 11990 12772 12012 18454
rect 950 12750 12012 12772
rect 950 12604 1058 12750
rect 11904 12604 12012 12750
rect 950 12582 12012 12604
rect 950 6900 972 12582
rect 11990 6900 12012 12582
rect 950 6878 12012 6900
rect 950 6732 1058 6878
rect 11904 6732 12012 6878
rect 950 6710 12012 6732
rect 950 1022 972 6710
rect 11990 1022 12012 6710
rect 950 1000 12012 1022
rect 950 654 1058 1000
rect 11904 654 12012 1000
rect 12358 654 12380 24700
rect 582 632 12380 654
<< nsubdiff >>
rect 32 25300 12930 25322
rect 32 54 54 25300
rect 400 24954 508 25300
rect 12454 24954 12562 25300
rect 400 24932 12562 24954
rect 400 422 422 24932
rect 12540 422 12562 24932
rect 400 400 12562 422
rect 400 54 508 400
rect 12454 54 12562 400
rect 12908 54 12930 25300
rect 32 32 12930 54
<< psubdiffcont >>
rect 604 654 950 24700
rect 1058 24354 11904 24700
rect 1058 18476 11904 18622
rect 1058 12604 11904 12750
rect 1058 6732 11904 6878
rect 1058 654 11904 1000
rect 12012 654 12358 24700
<< nsubdiffcont >>
rect 54 54 400 25300
rect 508 24954 12454 25300
rect 508 54 12454 400
rect 12562 54 12908 25300
<< polysilicon >>
rect 1237 23808 1481 23873
rect 1237 19162 1256 23808
rect 1402 23733 1481 23808
rect 11481 23808 11725 23873
rect 11481 23733 11560 23808
rect 1402 23629 1421 23733
rect 11541 23629 11560 23733
rect 1402 23489 1481 23629
rect 11481 23489 11560 23629
rect 1402 23385 1421 23489
rect 11541 23385 11560 23489
rect 1402 23245 1481 23385
rect 11481 23245 11560 23385
rect 1402 23141 1421 23245
rect 11541 23141 11560 23245
rect 1402 23001 1481 23141
rect 11481 23001 11560 23141
rect 1402 22897 1421 23001
rect 11541 22897 11560 23001
rect 1402 22757 1481 22897
rect 11481 22757 11560 22897
rect 1402 22653 1421 22757
rect 11541 22653 11560 22757
rect 1402 22513 1481 22653
rect 11481 22513 11560 22653
rect 1402 22409 1421 22513
rect 11541 22409 11560 22513
rect 1402 22269 1481 22409
rect 11481 22269 11560 22409
rect 1402 22165 1421 22269
rect 11541 22165 11560 22269
rect 1402 22025 1481 22165
rect 11481 22025 11560 22165
rect 1402 21921 1421 22025
rect 11541 21921 11560 22025
rect 1402 21781 1481 21921
rect 11481 21781 11560 21921
rect 1402 21677 1421 21781
rect 11541 21677 11560 21781
rect 1402 21537 1481 21677
rect 11481 21537 11560 21677
rect 1402 21433 1421 21537
rect 11541 21433 11560 21537
rect 1402 21293 1481 21433
rect 11481 21293 11560 21433
rect 1402 21189 1421 21293
rect 11541 21189 11560 21293
rect 1402 21049 1481 21189
rect 11481 21049 11560 21189
rect 1402 20945 1421 21049
rect 11541 20945 11560 21049
rect 1402 20805 1481 20945
rect 11481 20805 11560 20945
rect 1402 20701 1421 20805
rect 11541 20701 11560 20805
rect 1402 20561 1481 20701
rect 11481 20561 11560 20701
rect 1402 20457 1421 20561
rect 11541 20457 11560 20561
rect 1402 20317 1481 20457
rect 11481 20317 11560 20457
rect 1402 20213 1421 20317
rect 11541 20213 11560 20317
rect 1402 20073 1481 20213
rect 11481 20073 11560 20213
rect 1402 19969 1421 20073
rect 11541 19969 11560 20073
rect 1402 19829 1481 19969
rect 11481 19829 11560 19969
rect 1402 19725 1421 19829
rect 11541 19725 11560 19829
rect 1402 19585 1481 19725
rect 11481 19585 11560 19725
rect 1402 19481 1421 19585
rect 11541 19481 11560 19585
rect 1402 19341 1481 19481
rect 11481 19341 11560 19481
rect 1402 19237 1421 19341
rect 11541 19237 11560 19341
rect 1402 19162 1481 19237
rect 1237 19097 1481 19162
rect 11481 19162 11560 19237
rect 11706 19162 11725 23808
rect 11481 19097 11725 19162
rect 1237 17936 1481 18001
rect 1237 13290 1256 17936
rect 1402 17861 1481 17936
rect 11481 17936 11725 18001
rect 11481 17861 11560 17936
rect 1402 17757 1421 17861
rect 11541 17757 11560 17861
rect 1402 17617 1481 17757
rect 11481 17617 11560 17757
rect 1402 17513 1421 17617
rect 11541 17513 11560 17617
rect 1402 17373 1481 17513
rect 11481 17373 11560 17513
rect 1402 17269 1421 17373
rect 11541 17269 11560 17373
rect 1402 17129 1481 17269
rect 11481 17129 11560 17269
rect 1402 17025 1421 17129
rect 11541 17025 11560 17129
rect 1402 16885 1481 17025
rect 11481 16885 11560 17025
rect 1402 16781 1421 16885
rect 11541 16781 11560 16885
rect 1402 16641 1481 16781
rect 11481 16641 11560 16781
rect 1402 16537 1421 16641
rect 11541 16537 11560 16641
rect 1402 16397 1481 16537
rect 11481 16397 11560 16537
rect 1402 16293 1421 16397
rect 11541 16293 11560 16397
rect 1402 16153 1481 16293
rect 11481 16153 11560 16293
rect 1402 16049 1421 16153
rect 11541 16049 11560 16153
rect 1402 15909 1481 16049
rect 11481 15909 11560 16049
rect 1402 15805 1421 15909
rect 11541 15805 11560 15909
rect 1402 15665 1481 15805
rect 11481 15665 11560 15805
rect 1402 15561 1421 15665
rect 11541 15561 11560 15665
rect 1402 15421 1481 15561
rect 11481 15421 11560 15561
rect 1402 15317 1421 15421
rect 11541 15317 11560 15421
rect 1402 15177 1481 15317
rect 11481 15177 11560 15317
rect 1402 15073 1421 15177
rect 11541 15073 11560 15177
rect 1402 14933 1481 15073
rect 11481 14933 11560 15073
rect 1402 14829 1421 14933
rect 11541 14829 11560 14933
rect 1402 14689 1481 14829
rect 11481 14689 11560 14829
rect 1402 14585 1421 14689
rect 11541 14585 11560 14689
rect 1402 14445 1481 14585
rect 11481 14445 11560 14585
rect 1402 14341 1421 14445
rect 11541 14341 11560 14445
rect 1402 14201 1481 14341
rect 11481 14201 11560 14341
rect 1402 14097 1421 14201
rect 11541 14097 11560 14201
rect 1402 13957 1481 14097
rect 11481 13957 11560 14097
rect 1402 13853 1421 13957
rect 11541 13853 11560 13957
rect 1402 13713 1481 13853
rect 11481 13713 11560 13853
rect 1402 13609 1421 13713
rect 11541 13609 11560 13713
rect 1402 13469 1481 13609
rect 11481 13469 11560 13609
rect 1402 13365 1421 13469
rect 11541 13365 11560 13469
rect 1402 13290 1481 13365
rect 1237 13225 1481 13290
rect 11481 13290 11560 13365
rect 11706 13290 11725 17936
rect 11481 13225 11725 13290
rect 1237 12064 1481 12129
rect 1237 7418 1256 12064
rect 1402 11989 1481 12064
rect 11481 12064 11725 12129
rect 11481 11989 11560 12064
rect 1402 11885 1421 11989
rect 11541 11885 11560 11989
rect 1402 11745 1481 11885
rect 11481 11745 11560 11885
rect 1402 11641 1421 11745
rect 11541 11641 11560 11745
rect 1402 11501 1481 11641
rect 11481 11501 11560 11641
rect 1402 11397 1421 11501
rect 11541 11397 11560 11501
rect 1402 11257 1481 11397
rect 11481 11257 11560 11397
rect 1402 11153 1421 11257
rect 11541 11153 11560 11257
rect 1402 11013 1481 11153
rect 11481 11013 11560 11153
rect 1402 10909 1421 11013
rect 11541 10909 11560 11013
rect 1402 10769 1481 10909
rect 11481 10769 11560 10909
rect 1402 10665 1421 10769
rect 11541 10665 11560 10769
rect 1402 10525 1481 10665
rect 11481 10525 11560 10665
rect 1402 10421 1421 10525
rect 11541 10421 11560 10525
rect 1402 10281 1481 10421
rect 11481 10281 11560 10421
rect 1402 10177 1421 10281
rect 11541 10177 11560 10281
rect 1402 10037 1481 10177
rect 11481 10037 11560 10177
rect 1402 9933 1421 10037
rect 11541 9933 11560 10037
rect 1402 9793 1481 9933
rect 11481 9793 11560 9933
rect 1402 9689 1421 9793
rect 11541 9689 11560 9793
rect 1402 9549 1481 9689
rect 11481 9549 11560 9689
rect 1402 9445 1421 9549
rect 11541 9445 11560 9549
rect 1402 9305 1481 9445
rect 11481 9305 11560 9445
rect 1402 9201 1421 9305
rect 11541 9201 11560 9305
rect 1402 9061 1481 9201
rect 11481 9061 11560 9201
rect 1402 8957 1421 9061
rect 11541 8957 11560 9061
rect 1402 8817 1481 8957
rect 11481 8817 11560 8957
rect 1402 8713 1421 8817
rect 11541 8713 11560 8817
rect 1402 8573 1481 8713
rect 11481 8573 11560 8713
rect 1402 8469 1421 8573
rect 11541 8469 11560 8573
rect 1402 8329 1481 8469
rect 11481 8329 11560 8469
rect 1402 8225 1421 8329
rect 11541 8225 11560 8329
rect 1402 8085 1481 8225
rect 11481 8085 11560 8225
rect 1402 7981 1421 8085
rect 11541 7981 11560 8085
rect 1402 7841 1481 7981
rect 11481 7841 11560 7981
rect 1402 7737 1421 7841
rect 11541 7737 11560 7841
rect 1402 7597 1481 7737
rect 11481 7597 11560 7737
rect 1402 7493 1421 7597
rect 11541 7493 11560 7597
rect 1402 7418 1481 7493
rect 1237 7353 1481 7418
rect 11481 7418 11560 7493
rect 11706 7418 11725 12064
rect 11481 7353 11725 7418
rect 1237 6192 1481 6257
rect 1237 1546 1256 6192
rect 1402 6117 1481 6192
rect 11481 6192 11725 6257
rect 11481 6117 11560 6192
rect 1402 6013 1421 6117
rect 11541 6013 11560 6117
rect 1402 5873 1481 6013
rect 11481 5873 11560 6013
rect 1402 5769 1421 5873
rect 11541 5769 11560 5873
rect 1402 5629 1481 5769
rect 11481 5629 11560 5769
rect 1402 5525 1421 5629
rect 11541 5525 11560 5629
rect 1402 5385 1481 5525
rect 11481 5385 11560 5525
rect 1402 5281 1421 5385
rect 11541 5281 11560 5385
rect 1402 5141 1481 5281
rect 11481 5141 11560 5281
rect 1402 5037 1421 5141
rect 11541 5037 11560 5141
rect 1402 4897 1481 5037
rect 11481 4897 11560 5037
rect 1402 4793 1421 4897
rect 11541 4793 11560 4897
rect 1402 4653 1481 4793
rect 11481 4653 11560 4793
rect 1402 4549 1421 4653
rect 11541 4549 11560 4653
rect 1402 4409 1481 4549
rect 11481 4409 11560 4549
rect 1402 4305 1421 4409
rect 11541 4305 11560 4409
rect 1402 4165 1481 4305
rect 11481 4165 11560 4305
rect 1402 4061 1421 4165
rect 11541 4061 11560 4165
rect 1402 3921 1481 4061
rect 11481 3921 11560 4061
rect 1402 3817 1421 3921
rect 11541 3817 11560 3921
rect 1402 3677 1481 3817
rect 11481 3677 11560 3817
rect 1402 3573 1421 3677
rect 11541 3573 11560 3677
rect 1402 3433 1481 3573
rect 11481 3433 11560 3573
rect 1402 3329 1421 3433
rect 11541 3329 11560 3433
rect 1402 3189 1481 3329
rect 11481 3189 11560 3329
rect 1402 3085 1421 3189
rect 11541 3085 11560 3189
rect 1402 2945 1481 3085
rect 11481 2945 11560 3085
rect 1402 2841 1421 2945
rect 11541 2841 11560 2945
rect 1402 2701 1481 2841
rect 11481 2701 11560 2841
rect 1402 2597 1421 2701
rect 11541 2597 11560 2701
rect 1402 2457 1481 2597
rect 11481 2457 11560 2597
rect 1402 2353 1421 2457
rect 11541 2353 11560 2457
rect 1402 2213 1481 2353
rect 11481 2213 11560 2353
rect 1402 2109 1421 2213
rect 11541 2109 11560 2213
rect 1402 1969 1481 2109
rect 11481 1969 11560 2109
rect 1402 1865 1421 1969
rect 11541 1865 11560 1969
rect 1402 1725 1481 1865
rect 11481 1725 11560 1865
rect 1402 1621 1421 1725
rect 11541 1621 11560 1725
rect 1402 1546 1481 1621
rect 1237 1481 1481 1546
rect 11481 1546 11560 1621
rect 11706 1546 11725 6192
rect 11481 1481 11725 1546
<< polycontact >>
rect 1256 19162 1402 23808
rect 11560 19162 11706 23808
rect 1256 13290 1402 17936
rect 11560 13290 11706 17936
rect 1256 7418 1402 12064
rect 11560 7418 11706 12064
rect 1256 1546 1402 6192
rect 11560 1546 11706 6192
<< metal1 >>
rect 43 25300 12919 25311
rect 43 54 54 25300
rect 400 25261 508 25300
rect 400 25209 406 25261
rect 458 25209 508 25261
rect 400 25153 508 25209
rect 400 25101 406 25153
rect 458 25101 508 25153
rect 400 25045 508 25101
rect 400 24993 406 25045
rect 458 24993 508 25045
rect 400 24954 508 24993
rect 12454 24954 12562 25300
rect 400 24943 12562 24954
rect 400 411 411 24943
rect 593 24700 12369 24711
rect 593 654 604 24700
rect 950 24354 1058 24700
rect 11904 24354 12012 24700
rect 950 24343 12012 24354
rect 950 18641 961 24343
rect 1213 24053 11749 24253
rect 1213 23887 1413 24053
rect 1481 23951 11481 23963
rect 1481 23948 3433 23951
rect 3485 23948 3541 23951
rect 3593 23948 3649 23951
rect 3701 23948 3757 23951
rect 3809 23948 3865 23951
rect 3917 23948 3973 23951
rect 4025 23948 4081 23951
rect 4133 23948 4189 23951
rect 4241 23948 4297 23951
rect 4349 23948 4405 23951
rect 4457 23948 4513 23951
rect 4565 23948 4621 23951
rect 4673 23948 4729 23951
rect 4781 23948 4837 23951
rect 4889 23948 4945 23951
rect 4997 23948 5053 23951
rect 5105 23948 5161 23951
rect 5213 23948 6566 23951
rect 6618 23948 6674 23951
rect 6726 23948 6782 23951
rect 6834 23948 6890 23951
rect 6942 23948 6998 23951
rect 7050 23948 7106 23951
rect 7158 23948 7214 23951
rect 7266 23948 7322 23951
rect 7374 23948 7430 23951
rect 7482 23948 7538 23951
rect 7590 23948 9677 23951
rect 9729 23948 9785 23951
rect 9837 23948 9893 23951
rect 9945 23948 10001 23951
rect 10053 23948 10109 23951
rect 10161 23948 10217 23951
rect 10269 23948 10325 23951
rect 10377 23948 10433 23951
rect 10485 23948 10541 23951
rect 10593 23948 10649 23951
rect 10701 23948 10757 23951
rect 10809 23948 10865 23951
rect 10917 23948 10973 23951
rect 11025 23948 11081 23951
rect 11133 23948 11189 23951
rect 11241 23948 11297 23951
rect 11349 23948 11405 23951
rect 11457 23948 11481 23951
rect 1481 23902 1494 23948
rect 11468 23902 11481 23948
rect 1481 23899 3433 23902
rect 3485 23899 3541 23902
rect 3593 23899 3649 23902
rect 3701 23899 3757 23902
rect 3809 23899 3865 23902
rect 3917 23899 3973 23902
rect 4025 23899 4081 23902
rect 4133 23899 4189 23902
rect 4241 23899 4297 23902
rect 4349 23899 4405 23902
rect 4457 23899 4513 23902
rect 4565 23899 4621 23902
rect 4673 23899 4729 23902
rect 4781 23899 4837 23902
rect 4889 23899 4945 23902
rect 4997 23899 5053 23902
rect 5105 23899 5161 23902
rect 5213 23899 6566 23902
rect 6618 23899 6674 23902
rect 6726 23899 6782 23902
rect 6834 23899 6890 23902
rect 6942 23899 6998 23902
rect 7050 23899 7106 23902
rect 7158 23899 7214 23902
rect 7266 23899 7322 23902
rect 7374 23899 7430 23902
rect 7482 23899 7538 23902
rect 7590 23899 9677 23902
rect 9729 23899 9785 23902
rect 9837 23899 9893 23902
rect 9945 23899 10001 23902
rect 10053 23899 10109 23902
rect 10161 23899 10217 23902
rect 10269 23899 10325 23902
rect 10377 23899 10433 23902
rect 10485 23899 10541 23902
rect 10593 23899 10649 23902
rect 10701 23899 10757 23902
rect 10809 23899 10865 23902
rect 10917 23899 10973 23902
rect 11025 23899 11081 23902
rect 11133 23899 11189 23902
rect 11241 23899 11297 23902
rect 11349 23899 11405 23902
rect 11457 23899 11481 23902
rect 1481 23887 11481 23899
rect 11549 23887 11749 24053
rect 1213 23835 1233 23887
rect 1285 23835 1341 23887
rect 1393 23835 1413 23887
rect 1213 23808 1413 23835
rect 1213 23779 1256 23808
rect 1213 23727 1233 23779
rect 1213 23671 1256 23727
rect 1213 23619 1233 23671
rect 1213 23563 1256 23619
rect 1213 23511 1233 23563
rect 1213 23455 1256 23511
rect 1213 23403 1233 23455
rect 1213 23347 1256 23403
rect 1213 23295 1233 23347
rect 1213 23239 1256 23295
rect 1213 23187 1233 23239
rect 1213 23131 1256 23187
rect 1213 23079 1233 23131
rect 1213 23023 1256 23079
rect 1213 22971 1233 23023
rect 1213 22915 1256 22971
rect 1213 22863 1233 22915
rect 1213 22807 1256 22863
rect 1213 22755 1233 22807
rect 1213 22699 1256 22755
rect 1213 22647 1233 22699
rect 1213 22591 1256 22647
rect 1213 22539 1233 22591
rect 1213 22483 1256 22539
rect 1213 22431 1233 22483
rect 1213 22375 1256 22431
rect 1213 22323 1233 22375
rect 1213 22267 1256 22323
rect 1213 22215 1233 22267
rect 1213 22159 1256 22215
rect 1213 22107 1233 22159
rect 1213 22051 1256 22107
rect 1213 21999 1233 22051
rect 1213 21943 1256 21999
rect 1213 21891 1233 21943
rect 1213 21835 1256 21891
rect 1213 21783 1233 21835
rect 1213 21727 1256 21783
rect 1213 21675 1233 21727
rect 1213 21619 1256 21675
rect 1213 21567 1233 21619
rect 1213 21511 1256 21567
rect 1213 21459 1233 21511
rect 1213 21403 1256 21459
rect 1213 21351 1233 21403
rect 1213 21295 1256 21351
rect 1213 21243 1233 21295
rect 1213 21187 1256 21243
rect 1213 21135 1233 21187
rect 1213 21079 1256 21135
rect 1213 21027 1233 21079
rect 1213 20971 1256 21027
rect 1213 20919 1233 20971
rect 1213 20863 1256 20919
rect 1213 20811 1233 20863
rect 1213 20755 1256 20811
rect 1213 20703 1233 20755
rect 1213 20647 1256 20703
rect 1213 20595 1233 20647
rect 1213 20539 1256 20595
rect 1213 20487 1233 20539
rect 1213 20431 1256 20487
rect 1213 20379 1233 20431
rect 1213 20323 1256 20379
rect 1213 20271 1233 20323
rect 1213 20215 1256 20271
rect 1213 20163 1233 20215
rect 1213 20107 1256 20163
rect 1213 20055 1233 20107
rect 1213 19999 1256 20055
rect 1213 19947 1233 19999
rect 1213 19891 1256 19947
rect 1213 19839 1233 19891
rect 1213 19783 1256 19839
rect 1213 19731 1233 19783
rect 1213 19675 1256 19731
rect 1213 19623 1233 19675
rect 1213 19567 1256 19623
rect 1213 19515 1233 19567
rect 1213 19459 1256 19515
rect 1213 19407 1233 19459
rect 1213 19351 1256 19407
rect 1213 19299 1233 19351
rect 1213 19243 1256 19299
rect 1213 19191 1233 19243
rect 1213 19162 1256 19191
rect 1402 19162 1413 23808
rect 11549 23835 11569 23887
rect 11621 23835 11677 23887
rect 11729 23835 11749 23887
rect 11549 23808 11749 23835
rect 1481 23707 11481 23719
rect 1481 23704 1505 23707
rect 1557 23704 1613 23707
rect 1665 23704 1721 23707
rect 1773 23704 1829 23707
rect 1881 23704 1937 23707
rect 1989 23704 2045 23707
rect 2097 23704 2153 23707
rect 2205 23704 2261 23707
rect 2313 23704 2369 23707
rect 2421 23704 2477 23707
rect 2529 23704 2585 23707
rect 2637 23704 2693 23707
rect 2745 23704 2801 23707
rect 2853 23704 2909 23707
rect 2961 23704 3017 23707
rect 3069 23704 3125 23707
rect 3177 23704 3233 23707
rect 3285 23704 5372 23707
rect 5424 23704 5480 23707
rect 5532 23704 5588 23707
rect 5640 23704 5696 23707
rect 5748 23704 5804 23707
rect 5856 23704 5912 23707
rect 5964 23704 6020 23707
rect 6072 23704 6128 23707
rect 6180 23704 6236 23707
rect 6288 23704 6344 23707
rect 6396 23704 7749 23707
rect 7801 23704 7857 23707
rect 7909 23704 7965 23707
rect 8017 23704 8073 23707
rect 8125 23704 8181 23707
rect 8233 23704 8289 23707
rect 8341 23704 8397 23707
rect 8449 23704 8505 23707
rect 8557 23704 8613 23707
rect 8665 23704 8721 23707
rect 8773 23704 8829 23707
rect 8881 23704 8937 23707
rect 8989 23704 9045 23707
rect 9097 23704 9153 23707
rect 9205 23704 9261 23707
rect 9313 23704 9369 23707
rect 9421 23704 9477 23707
rect 9529 23704 11481 23707
rect 1481 23658 1494 23704
rect 11468 23658 11481 23704
rect 1481 23655 1505 23658
rect 1557 23655 1613 23658
rect 1665 23655 1721 23658
rect 1773 23655 1829 23658
rect 1881 23655 1937 23658
rect 1989 23655 2045 23658
rect 2097 23655 2153 23658
rect 2205 23655 2261 23658
rect 2313 23655 2369 23658
rect 2421 23655 2477 23658
rect 2529 23655 2585 23658
rect 2637 23655 2693 23658
rect 2745 23655 2801 23658
rect 2853 23655 2909 23658
rect 2961 23655 3017 23658
rect 3069 23655 3125 23658
rect 3177 23655 3233 23658
rect 3285 23655 5372 23658
rect 5424 23655 5480 23658
rect 5532 23655 5588 23658
rect 5640 23655 5696 23658
rect 5748 23655 5804 23658
rect 5856 23655 5912 23658
rect 5964 23655 6020 23658
rect 6072 23655 6128 23658
rect 6180 23655 6236 23658
rect 6288 23655 6344 23658
rect 6396 23655 7749 23658
rect 7801 23655 7857 23658
rect 7909 23655 7965 23658
rect 8017 23655 8073 23658
rect 8125 23655 8181 23658
rect 8233 23655 8289 23658
rect 8341 23655 8397 23658
rect 8449 23655 8505 23658
rect 8557 23655 8613 23658
rect 8665 23655 8721 23658
rect 8773 23655 8829 23658
rect 8881 23655 8937 23658
rect 8989 23655 9045 23658
rect 9097 23655 9153 23658
rect 9205 23655 9261 23658
rect 9313 23655 9369 23658
rect 9421 23655 9477 23658
rect 9529 23655 11481 23658
rect 1481 23643 11481 23655
rect 1481 23463 11481 23475
rect 1481 23460 3433 23463
rect 3485 23460 3541 23463
rect 3593 23460 3649 23463
rect 3701 23460 3757 23463
rect 3809 23460 3865 23463
rect 3917 23460 3973 23463
rect 4025 23460 4081 23463
rect 4133 23460 4189 23463
rect 4241 23460 4297 23463
rect 4349 23460 4405 23463
rect 4457 23460 4513 23463
rect 4565 23460 4621 23463
rect 4673 23460 4729 23463
rect 4781 23460 4837 23463
rect 4889 23460 4945 23463
rect 4997 23460 5053 23463
rect 5105 23460 5161 23463
rect 5213 23460 6566 23463
rect 6618 23460 6674 23463
rect 6726 23460 6782 23463
rect 6834 23460 6890 23463
rect 6942 23460 6998 23463
rect 7050 23460 7106 23463
rect 7158 23460 7214 23463
rect 7266 23460 7322 23463
rect 7374 23460 7430 23463
rect 7482 23460 7538 23463
rect 7590 23460 9677 23463
rect 9729 23460 9785 23463
rect 9837 23460 9893 23463
rect 9945 23460 10001 23463
rect 10053 23460 10109 23463
rect 10161 23460 10217 23463
rect 10269 23460 10325 23463
rect 10377 23460 10433 23463
rect 10485 23460 10541 23463
rect 10593 23460 10649 23463
rect 10701 23460 10757 23463
rect 10809 23460 10865 23463
rect 10917 23460 10973 23463
rect 11025 23460 11081 23463
rect 11133 23460 11189 23463
rect 11241 23460 11297 23463
rect 11349 23460 11405 23463
rect 11457 23460 11481 23463
rect 1481 23414 1494 23460
rect 11468 23414 11481 23460
rect 1481 23411 3433 23414
rect 3485 23411 3541 23414
rect 3593 23411 3649 23414
rect 3701 23411 3757 23414
rect 3809 23411 3865 23414
rect 3917 23411 3973 23414
rect 4025 23411 4081 23414
rect 4133 23411 4189 23414
rect 4241 23411 4297 23414
rect 4349 23411 4405 23414
rect 4457 23411 4513 23414
rect 4565 23411 4621 23414
rect 4673 23411 4729 23414
rect 4781 23411 4837 23414
rect 4889 23411 4945 23414
rect 4997 23411 5053 23414
rect 5105 23411 5161 23414
rect 5213 23411 6566 23414
rect 6618 23411 6674 23414
rect 6726 23411 6782 23414
rect 6834 23411 6890 23414
rect 6942 23411 6998 23414
rect 7050 23411 7106 23414
rect 7158 23411 7214 23414
rect 7266 23411 7322 23414
rect 7374 23411 7430 23414
rect 7482 23411 7538 23414
rect 7590 23411 9677 23414
rect 9729 23411 9785 23414
rect 9837 23411 9893 23414
rect 9945 23411 10001 23414
rect 10053 23411 10109 23414
rect 10161 23411 10217 23414
rect 10269 23411 10325 23414
rect 10377 23411 10433 23414
rect 10485 23411 10541 23414
rect 10593 23411 10649 23414
rect 10701 23411 10757 23414
rect 10809 23411 10865 23414
rect 10917 23411 10973 23414
rect 11025 23411 11081 23414
rect 11133 23411 11189 23414
rect 11241 23411 11297 23414
rect 11349 23411 11405 23414
rect 11457 23411 11481 23414
rect 1481 23399 11481 23411
rect 1481 23219 11481 23231
rect 1481 23216 1505 23219
rect 1557 23216 1613 23219
rect 1665 23216 1721 23219
rect 1773 23216 1829 23219
rect 1881 23216 1937 23219
rect 1989 23216 2045 23219
rect 2097 23216 2153 23219
rect 2205 23216 2261 23219
rect 2313 23216 2369 23219
rect 2421 23216 2477 23219
rect 2529 23216 2585 23219
rect 2637 23216 2693 23219
rect 2745 23216 2801 23219
rect 2853 23216 2909 23219
rect 2961 23216 3017 23219
rect 3069 23216 3125 23219
rect 3177 23216 3233 23219
rect 3285 23216 5372 23219
rect 5424 23216 5480 23219
rect 5532 23216 5588 23219
rect 5640 23216 5696 23219
rect 5748 23216 5804 23219
rect 5856 23216 5912 23219
rect 5964 23216 6020 23219
rect 6072 23216 6128 23219
rect 6180 23216 6236 23219
rect 6288 23216 6344 23219
rect 6396 23216 7749 23219
rect 7801 23216 7857 23219
rect 7909 23216 7965 23219
rect 8017 23216 8073 23219
rect 8125 23216 8181 23219
rect 8233 23216 8289 23219
rect 8341 23216 8397 23219
rect 8449 23216 8505 23219
rect 8557 23216 8613 23219
rect 8665 23216 8721 23219
rect 8773 23216 8829 23219
rect 8881 23216 8937 23219
rect 8989 23216 9045 23219
rect 9097 23216 9153 23219
rect 9205 23216 9261 23219
rect 9313 23216 9369 23219
rect 9421 23216 9477 23219
rect 9529 23216 11481 23219
rect 1481 23170 1494 23216
rect 11468 23170 11481 23216
rect 1481 23167 1505 23170
rect 1557 23167 1613 23170
rect 1665 23167 1721 23170
rect 1773 23167 1829 23170
rect 1881 23167 1937 23170
rect 1989 23167 2045 23170
rect 2097 23167 2153 23170
rect 2205 23167 2261 23170
rect 2313 23167 2369 23170
rect 2421 23167 2477 23170
rect 2529 23167 2585 23170
rect 2637 23167 2693 23170
rect 2745 23167 2801 23170
rect 2853 23167 2909 23170
rect 2961 23167 3017 23170
rect 3069 23167 3125 23170
rect 3177 23167 3233 23170
rect 3285 23167 5372 23170
rect 5424 23167 5480 23170
rect 5532 23167 5588 23170
rect 5640 23167 5696 23170
rect 5748 23167 5804 23170
rect 5856 23167 5912 23170
rect 5964 23167 6020 23170
rect 6072 23167 6128 23170
rect 6180 23167 6236 23170
rect 6288 23167 6344 23170
rect 6396 23167 7749 23170
rect 7801 23167 7857 23170
rect 7909 23167 7965 23170
rect 8017 23167 8073 23170
rect 8125 23167 8181 23170
rect 8233 23167 8289 23170
rect 8341 23167 8397 23170
rect 8449 23167 8505 23170
rect 8557 23167 8613 23170
rect 8665 23167 8721 23170
rect 8773 23167 8829 23170
rect 8881 23167 8937 23170
rect 8989 23167 9045 23170
rect 9097 23167 9153 23170
rect 9205 23167 9261 23170
rect 9313 23167 9369 23170
rect 9421 23167 9477 23170
rect 9529 23167 11481 23170
rect 1481 23155 11481 23167
rect 1481 22975 11481 22987
rect 1481 22972 3433 22975
rect 3485 22972 3541 22975
rect 3593 22972 3649 22975
rect 3701 22972 3757 22975
rect 3809 22972 3865 22975
rect 3917 22972 3973 22975
rect 4025 22972 4081 22975
rect 4133 22972 4189 22975
rect 4241 22972 4297 22975
rect 4349 22972 4405 22975
rect 4457 22972 4513 22975
rect 4565 22972 4621 22975
rect 4673 22972 4729 22975
rect 4781 22972 4837 22975
rect 4889 22972 4945 22975
rect 4997 22972 5053 22975
rect 5105 22972 5161 22975
rect 5213 22972 6566 22975
rect 6618 22972 6674 22975
rect 6726 22972 6782 22975
rect 6834 22972 6890 22975
rect 6942 22972 6998 22975
rect 7050 22972 7106 22975
rect 7158 22972 7214 22975
rect 7266 22972 7322 22975
rect 7374 22972 7430 22975
rect 7482 22972 7538 22975
rect 7590 22972 9677 22975
rect 9729 22972 9785 22975
rect 9837 22972 9893 22975
rect 9945 22972 10001 22975
rect 10053 22972 10109 22975
rect 10161 22972 10217 22975
rect 10269 22972 10325 22975
rect 10377 22972 10433 22975
rect 10485 22972 10541 22975
rect 10593 22972 10649 22975
rect 10701 22972 10757 22975
rect 10809 22972 10865 22975
rect 10917 22972 10973 22975
rect 11025 22972 11081 22975
rect 11133 22972 11189 22975
rect 11241 22972 11297 22975
rect 11349 22972 11405 22975
rect 11457 22972 11481 22975
rect 1481 22926 1494 22972
rect 11468 22926 11481 22972
rect 1481 22923 3433 22926
rect 3485 22923 3541 22926
rect 3593 22923 3649 22926
rect 3701 22923 3757 22926
rect 3809 22923 3865 22926
rect 3917 22923 3973 22926
rect 4025 22923 4081 22926
rect 4133 22923 4189 22926
rect 4241 22923 4297 22926
rect 4349 22923 4405 22926
rect 4457 22923 4513 22926
rect 4565 22923 4621 22926
rect 4673 22923 4729 22926
rect 4781 22923 4837 22926
rect 4889 22923 4945 22926
rect 4997 22923 5053 22926
rect 5105 22923 5161 22926
rect 5213 22923 6566 22926
rect 6618 22923 6674 22926
rect 6726 22923 6782 22926
rect 6834 22923 6890 22926
rect 6942 22923 6998 22926
rect 7050 22923 7106 22926
rect 7158 22923 7214 22926
rect 7266 22923 7322 22926
rect 7374 22923 7430 22926
rect 7482 22923 7538 22926
rect 7590 22923 9677 22926
rect 9729 22923 9785 22926
rect 9837 22923 9893 22926
rect 9945 22923 10001 22926
rect 10053 22923 10109 22926
rect 10161 22923 10217 22926
rect 10269 22923 10325 22926
rect 10377 22923 10433 22926
rect 10485 22923 10541 22926
rect 10593 22923 10649 22926
rect 10701 22923 10757 22926
rect 10809 22923 10865 22926
rect 10917 22923 10973 22926
rect 11025 22923 11081 22926
rect 11133 22923 11189 22926
rect 11241 22923 11297 22926
rect 11349 22923 11405 22926
rect 11457 22923 11481 22926
rect 1481 22911 11481 22923
rect 1481 22731 11481 22743
rect 1481 22728 1505 22731
rect 1557 22728 1613 22731
rect 1665 22728 1721 22731
rect 1773 22728 1829 22731
rect 1881 22728 1937 22731
rect 1989 22728 2045 22731
rect 2097 22728 2153 22731
rect 2205 22728 2261 22731
rect 2313 22728 2369 22731
rect 2421 22728 2477 22731
rect 2529 22728 2585 22731
rect 2637 22728 2693 22731
rect 2745 22728 2801 22731
rect 2853 22728 2909 22731
rect 2961 22728 3017 22731
rect 3069 22728 3125 22731
rect 3177 22728 3233 22731
rect 3285 22728 5372 22731
rect 5424 22728 5480 22731
rect 5532 22728 5588 22731
rect 5640 22728 5696 22731
rect 5748 22728 5804 22731
rect 5856 22728 5912 22731
rect 5964 22728 6020 22731
rect 6072 22728 6128 22731
rect 6180 22728 6236 22731
rect 6288 22728 6344 22731
rect 6396 22728 7749 22731
rect 7801 22728 7857 22731
rect 7909 22728 7965 22731
rect 8017 22728 8073 22731
rect 8125 22728 8181 22731
rect 8233 22728 8289 22731
rect 8341 22728 8397 22731
rect 8449 22728 8505 22731
rect 8557 22728 8613 22731
rect 8665 22728 8721 22731
rect 8773 22728 8829 22731
rect 8881 22728 8937 22731
rect 8989 22728 9045 22731
rect 9097 22728 9153 22731
rect 9205 22728 9261 22731
rect 9313 22728 9369 22731
rect 9421 22728 9477 22731
rect 9529 22728 11481 22731
rect 1481 22682 1494 22728
rect 11468 22682 11481 22728
rect 1481 22679 1505 22682
rect 1557 22679 1613 22682
rect 1665 22679 1721 22682
rect 1773 22679 1829 22682
rect 1881 22679 1937 22682
rect 1989 22679 2045 22682
rect 2097 22679 2153 22682
rect 2205 22679 2261 22682
rect 2313 22679 2369 22682
rect 2421 22679 2477 22682
rect 2529 22679 2585 22682
rect 2637 22679 2693 22682
rect 2745 22679 2801 22682
rect 2853 22679 2909 22682
rect 2961 22679 3017 22682
rect 3069 22679 3125 22682
rect 3177 22679 3233 22682
rect 3285 22679 5372 22682
rect 5424 22679 5480 22682
rect 5532 22679 5588 22682
rect 5640 22679 5696 22682
rect 5748 22679 5804 22682
rect 5856 22679 5912 22682
rect 5964 22679 6020 22682
rect 6072 22679 6128 22682
rect 6180 22679 6236 22682
rect 6288 22679 6344 22682
rect 6396 22679 7749 22682
rect 7801 22679 7857 22682
rect 7909 22679 7965 22682
rect 8017 22679 8073 22682
rect 8125 22679 8181 22682
rect 8233 22679 8289 22682
rect 8341 22679 8397 22682
rect 8449 22679 8505 22682
rect 8557 22679 8613 22682
rect 8665 22679 8721 22682
rect 8773 22679 8829 22682
rect 8881 22679 8937 22682
rect 8989 22679 9045 22682
rect 9097 22679 9153 22682
rect 9205 22679 9261 22682
rect 9313 22679 9369 22682
rect 9421 22679 9477 22682
rect 9529 22679 11481 22682
rect 1481 22667 11481 22679
rect 1481 22487 11481 22499
rect 1481 22484 3433 22487
rect 3485 22484 3541 22487
rect 3593 22484 3649 22487
rect 3701 22484 3757 22487
rect 3809 22484 3865 22487
rect 3917 22484 3973 22487
rect 4025 22484 4081 22487
rect 4133 22484 4189 22487
rect 4241 22484 4297 22487
rect 4349 22484 4405 22487
rect 4457 22484 4513 22487
rect 4565 22484 4621 22487
rect 4673 22484 4729 22487
rect 4781 22484 4837 22487
rect 4889 22484 4945 22487
rect 4997 22484 5053 22487
rect 5105 22484 5161 22487
rect 5213 22484 6566 22487
rect 6618 22484 6674 22487
rect 6726 22484 6782 22487
rect 6834 22484 6890 22487
rect 6942 22484 6998 22487
rect 7050 22484 7106 22487
rect 7158 22484 7214 22487
rect 7266 22484 7322 22487
rect 7374 22484 7430 22487
rect 7482 22484 7538 22487
rect 7590 22484 9677 22487
rect 9729 22484 9785 22487
rect 9837 22484 9893 22487
rect 9945 22484 10001 22487
rect 10053 22484 10109 22487
rect 10161 22484 10217 22487
rect 10269 22484 10325 22487
rect 10377 22484 10433 22487
rect 10485 22484 10541 22487
rect 10593 22484 10649 22487
rect 10701 22484 10757 22487
rect 10809 22484 10865 22487
rect 10917 22484 10973 22487
rect 11025 22484 11081 22487
rect 11133 22484 11189 22487
rect 11241 22484 11297 22487
rect 11349 22484 11405 22487
rect 11457 22484 11481 22487
rect 1481 22438 1494 22484
rect 11468 22438 11481 22484
rect 1481 22435 3433 22438
rect 3485 22435 3541 22438
rect 3593 22435 3649 22438
rect 3701 22435 3757 22438
rect 3809 22435 3865 22438
rect 3917 22435 3973 22438
rect 4025 22435 4081 22438
rect 4133 22435 4189 22438
rect 4241 22435 4297 22438
rect 4349 22435 4405 22438
rect 4457 22435 4513 22438
rect 4565 22435 4621 22438
rect 4673 22435 4729 22438
rect 4781 22435 4837 22438
rect 4889 22435 4945 22438
rect 4997 22435 5053 22438
rect 5105 22435 5161 22438
rect 5213 22435 6566 22438
rect 6618 22435 6674 22438
rect 6726 22435 6782 22438
rect 6834 22435 6890 22438
rect 6942 22435 6998 22438
rect 7050 22435 7106 22438
rect 7158 22435 7214 22438
rect 7266 22435 7322 22438
rect 7374 22435 7430 22438
rect 7482 22435 7538 22438
rect 7590 22435 9677 22438
rect 9729 22435 9785 22438
rect 9837 22435 9893 22438
rect 9945 22435 10001 22438
rect 10053 22435 10109 22438
rect 10161 22435 10217 22438
rect 10269 22435 10325 22438
rect 10377 22435 10433 22438
rect 10485 22435 10541 22438
rect 10593 22435 10649 22438
rect 10701 22435 10757 22438
rect 10809 22435 10865 22438
rect 10917 22435 10973 22438
rect 11025 22435 11081 22438
rect 11133 22435 11189 22438
rect 11241 22435 11297 22438
rect 11349 22435 11405 22438
rect 11457 22435 11481 22438
rect 1481 22423 11481 22435
rect 1481 22243 11481 22255
rect 1481 22240 1505 22243
rect 1557 22240 1613 22243
rect 1665 22240 1721 22243
rect 1773 22240 1829 22243
rect 1881 22240 1937 22243
rect 1989 22240 2045 22243
rect 2097 22240 2153 22243
rect 2205 22240 2261 22243
rect 2313 22240 2369 22243
rect 2421 22240 2477 22243
rect 2529 22240 2585 22243
rect 2637 22240 2693 22243
rect 2745 22240 2801 22243
rect 2853 22240 2909 22243
rect 2961 22240 3017 22243
rect 3069 22240 3125 22243
rect 3177 22240 3233 22243
rect 3285 22240 5372 22243
rect 5424 22240 5480 22243
rect 5532 22240 5588 22243
rect 5640 22240 5696 22243
rect 5748 22240 5804 22243
rect 5856 22240 5912 22243
rect 5964 22240 6020 22243
rect 6072 22240 6128 22243
rect 6180 22240 6236 22243
rect 6288 22240 6344 22243
rect 6396 22240 7749 22243
rect 7801 22240 7857 22243
rect 7909 22240 7965 22243
rect 8017 22240 8073 22243
rect 8125 22240 8181 22243
rect 8233 22240 8289 22243
rect 8341 22240 8397 22243
rect 8449 22240 8505 22243
rect 8557 22240 8613 22243
rect 8665 22240 8721 22243
rect 8773 22240 8829 22243
rect 8881 22240 8937 22243
rect 8989 22240 9045 22243
rect 9097 22240 9153 22243
rect 9205 22240 9261 22243
rect 9313 22240 9369 22243
rect 9421 22240 9477 22243
rect 9529 22240 11481 22243
rect 1481 22194 1494 22240
rect 11468 22194 11481 22240
rect 1481 22191 1505 22194
rect 1557 22191 1613 22194
rect 1665 22191 1721 22194
rect 1773 22191 1829 22194
rect 1881 22191 1937 22194
rect 1989 22191 2045 22194
rect 2097 22191 2153 22194
rect 2205 22191 2261 22194
rect 2313 22191 2369 22194
rect 2421 22191 2477 22194
rect 2529 22191 2585 22194
rect 2637 22191 2693 22194
rect 2745 22191 2801 22194
rect 2853 22191 2909 22194
rect 2961 22191 3017 22194
rect 3069 22191 3125 22194
rect 3177 22191 3233 22194
rect 3285 22191 5372 22194
rect 5424 22191 5480 22194
rect 5532 22191 5588 22194
rect 5640 22191 5696 22194
rect 5748 22191 5804 22194
rect 5856 22191 5912 22194
rect 5964 22191 6020 22194
rect 6072 22191 6128 22194
rect 6180 22191 6236 22194
rect 6288 22191 6344 22194
rect 6396 22191 7749 22194
rect 7801 22191 7857 22194
rect 7909 22191 7965 22194
rect 8017 22191 8073 22194
rect 8125 22191 8181 22194
rect 8233 22191 8289 22194
rect 8341 22191 8397 22194
rect 8449 22191 8505 22194
rect 8557 22191 8613 22194
rect 8665 22191 8721 22194
rect 8773 22191 8829 22194
rect 8881 22191 8937 22194
rect 8989 22191 9045 22194
rect 9097 22191 9153 22194
rect 9205 22191 9261 22194
rect 9313 22191 9369 22194
rect 9421 22191 9477 22194
rect 9529 22191 11481 22194
rect 1481 22179 11481 22191
rect 1481 21999 11481 22011
rect 1481 21996 3433 21999
rect 3485 21996 3541 21999
rect 3593 21996 3649 21999
rect 3701 21996 3757 21999
rect 3809 21996 3865 21999
rect 3917 21996 3973 21999
rect 4025 21996 4081 21999
rect 4133 21996 4189 21999
rect 4241 21996 4297 21999
rect 4349 21996 4405 21999
rect 4457 21996 4513 21999
rect 4565 21996 4621 21999
rect 4673 21996 4729 21999
rect 4781 21996 4837 21999
rect 4889 21996 4945 21999
rect 4997 21996 5053 21999
rect 5105 21996 5161 21999
rect 5213 21996 6566 21999
rect 6618 21996 6674 21999
rect 6726 21996 6782 21999
rect 6834 21996 6890 21999
rect 6942 21996 6998 21999
rect 7050 21996 7106 21999
rect 7158 21996 7214 21999
rect 7266 21996 7322 21999
rect 7374 21996 7430 21999
rect 7482 21996 7538 21999
rect 7590 21996 9677 21999
rect 9729 21996 9785 21999
rect 9837 21996 9893 21999
rect 9945 21996 10001 21999
rect 10053 21996 10109 21999
rect 10161 21996 10217 21999
rect 10269 21996 10325 21999
rect 10377 21996 10433 21999
rect 10485 21996 10541 21999
rect 10593 21996 10649 21999
rect 10701 21996 10757 21999
rect 10809 21996 10865 21999
rect 10917 21996 10973 21999
rect 11025 21996 11081 21999
rect 11133 21996 11189 21999
rect 11241 21996 11297 21999
rect 11349 21996 11405 21999
rect 11457 21996 11481 21999
rect 1481 21950 1494 21996
rect 11468 21950 11481 21996
rect 1481 21947 3433 21950
rect 3485 21947 3541 21950
rect 3593 21947 3649 21950
rect 3701 21947 3757 21950
rect 3809 21947 3865 21950
rect 3917 21947 3973 21950
rect 4025 21947 4081 21950
rect 4133 21947 4189 21950
rect 4241 21947 4297 21950
rect 4349 21947 4405 21950
rect 4457 21947 4513 21950
rect 4565 21947 4621 21950
rect 4673 21947 4729 21950
rect 4781 21947 4837 21950
rect 4889 21947 4945 21950
rect 4997 21947 5053 21950
rect 5105 21947 5161 21950
rect 5213 21947 6566 21950
rect 6618 21947 6674 21950
rect 6726 21947 6782 21950
rect 6834 21947 6890 21950
rect 6942 21947 6998 21950
rect 7050 21947 7106 21950
rect 7158 21947 7214 21950
rect 7266 21947 7322 21950
rect 7374 21947 7430 21950
rect 7482 21947 7538 21950
rect 7590 21947 9677 21950
rect 9729 21947 9785 21950
rect 9837 21947 9893 21950
rect 9945 21947 10001 21950
rect 10053 21947 10109 21950
rect 10161 21947 10217 21950
rect 10269 21947 10325 21950
rect 10377 21947 10433 21950
rect 10485 21947 10541 21950
rect 10593 21947 10649 21950
rect 10701 21947 10757 21950
rect 10809 21947 10865 21950
rect 10917 21947 10973 21950
rect 11025 21947 11081 21950
rect 11133 21947 11189 21950
rect 11241 21947 11297 21950
rect 11349 21947 11405 21950
rect 11457 21947 11481 21950
rect 1481 21935 11481 21947
rect 1481 21755 11481 21767
rect 1481 21752 1505 21755
rect 1557 21752 1613 21755
rect 1665 21752 1721 21755
rect 1773 21752 1829 21755
rect 1881 21752 1937 21755
rect 1989 21752 2045 21755
rect 2097 21752 2153 21755
rect 2205 21752 2261 21755
rect 2313 21752 2369 21755
rect 2421 21752 2477 21755
rect 2529 21752 2585 21755
rect 2637 21752 2693 21755
rect 2745 21752 2801 21755
rect 2853 21752 2909 21755
rect 2961 21752 3017 21755
rect 3069 21752 3125 21755
rect 3177 21752 3233 21755
rect 3285 21752 5372 21755
rect 5424 21752 5480 21755
rect 5532 21752 5588 21755
rect 5640 21752 5696 21755
rect 5748 21752 5804 21755
rect 5856 21752 5912 21755
rect 5964 21752 6020 21755
rect 6072 21752 6128 21755
rect 6180 21752 6236 21755
rect 6288 21752 6344 21755
rect 6396 21752 7749 21755
rect 7801 21752 7857 21755
rect 7909 21752 7965 21755
rect 8017 21752 8073 21755
rect 8125 21752 8181 21755
rect 8233 21752 8289 21755
rect 8341 21752 8397 21755
rect 8449 21752 8505 21755
rect 8557 21752 8613 21755
rect 8665 21752 8721 21755
rect 8773 21752 8829 21755
rect 8881 21752 8937 21755
rect 8989 21752 9045 21755
rect 9097 21752 9153 21755
rect 9205 21752 9261 21755
rect 9313 21752 9369 21755
rect 9421 21752 9477 21755
rect 9529 21752 11481 21755
rect 1481 21706 1494 21752
rect 11468 21706 11481 21752
rect 1481 21703 1505 21706
rect 1557 21703 1613 21706
rect 1665 21703 1721 21706
rect 1773 21703 1829 21706
rect 1881 21703 1937 21706
rect 1989 21703 2045 21706
rect 2097 21703 2153 21706
rect 2205 21703 2261 21706
rect 2313 21703 2369 21706
rect 2421 21703 2477 21706
rect 2529 21703 2585 21706
rect 2637 21703 2693 21706
rect 2745 21703 2801 21706
rect 2853 21703 2909 21706
rect 2961 21703 3017 21706
rect 3069 21703 3125 21706
rect 3177 21703 3233 21706
rect 3285 21703 5372 21706
rect 5424 21703 5480 21706
rect 5532 21703 5588 21706
rect 5640 21703 5696 21706
rect 5748 21703 5804 21706
rect 5856 21703 5912 21706
rect 5964 21703 6020 21706
rect 6072 21703 6128 21706
rect 6180 21703 6236 21706
rect 6288 21703 6344 21706
rect 6396 21703 7749 21706
rect 7801 21703 7857 21706
rect 7909 21703 7965 21706
rect 8017 21703 8073 21706
rect 8125 21703 8181 21706
rect 8233 21703 8289 21706
rect 8341 21703 8397 21706
rect 8449 21703 8505 21706
rect 8557 21703 8613 21706
rect 8665 21703 8721 21706
rect 8773 21703 8829 21706
rect 8881 21703 8937 21706
rect 8989 21703 9045 21706
rect 9097 21703 9153 21706
rect 9205 21703 9261 21706
rect 9313 21703 9369 21706
rect 9421 21703 9477 21706
rect 9529 21703 11481 21706
rect 1481 21691 11481 21703
rect 1481 21511 11481 21523
rect 1481 21508 3433 21511
rect 3485 21508 3541 21511
rect 3593 21508 3649 21511
rect 3701 21508 3757 21511
rect 3809 21508 3865 21511
rect 3917 21508 3973 21511
rect 4025 21508 4081 21511
rect 4133 21508 4189 21511
rect 4241 21508 4297 21511
rect 4349 21508 4405 21511
rect 4457 21508 4513 21511
rect 4565 21508 4621 21511
rect 4673 21508 4729 21511
rect 4781 21508 4837 21511
rect 4889 21508 4945 21511
rect 4997 21508 5053 21511
rect 5105 21508 5161 21511
rect 5213 21508 6566 21511
rect 6618 21508 6674 21511
rect 6726 21508 6782 21511
rect 6834 21508 6890 21511
rect 6942 21508 6998 21511
rect 7050 21508 7106 21511
rect 7158 21508 7214 21511
rect 7266 21508 7322 21511
rect 7374 21508 7430 21511
rect 7482 21508 7538 21511
rect 7590 21508 9677 21511
rect 9729 21508 9785 21511
rect 9837 21508 9893 21511
rect 9945 21508 10001 21511
rect 10053 21508 10109 21511
rect 10161 21508 10217 21511
rect 10269 21508 10325 21511
rect 10377 21508 10433 21511
rect 10485 21508 10541 21511
rect 10593 21508 10649 21511
rect 10701 21508 10757 21511
rect 10809 21508 10865 21511
rect 10917 21508 10973 21511
rect 11025 21508 11081 21511
rect 11133 21508 11189 21511
rect 11241 21508 11297 21511
rect 11349 21508 11405 21511
rect 11457 21508 11481 21511
rect 1481 21462 1494 21508
rect 11468 21462 11481 21508
rect 1481 21459 3433 21462
rect 3485 21459 3541 21462
rect 3593 21459 3649 21462
rect 3701 21459 3757 21462
rect 3809 21459 3865 21462
rect 3917 21459 3973 21462
rect 4025 21459 4081 21462
rect 4133 21459 4189 21462
rect 4241 21459 4297 21462
rect 4349 21459 4405 21462
rect 4457 21459 4513 21462
rect 4565 21459 4621 21462
rect 4673 21459 4729 21462
rect 4781 21459 4837 21462
rect 4889 21459 4945 21462
rect 4997 21459 5053 21462
rect 5105 21459 5161 21462
rect 5213 21459 6566 21462
rect 6618 21459 6674 21462
rect 6726 21459 6782 21462
rect 6834 21459 6890 21462
rect 6942 21459 6998 21462
rect 7050 21459 7106 21462
rect 7158 21459 7214 21462
rect 7266 21459 7322 21462
rect 7374 21459 7430 21462
rect 7482 21459 7538 21462
rect 7590 21459 9677 21462
rect 9729 21459 9785 21462
rect 9837 21459 9893 21462
rect 9945 21459 10001 21462
rect 10053 21459 10109 21462
rect 10161 21459 10217 21462
rect 10269 21459 10325 21462
rect 10377 21459 10433 21462
rect 10485 21459 10541 21462
rect 10593 21459 10649 21462
rect 10701 21459 10757 21462
rect 10809 21459 10865 21462
rect 10917 21459 10973 21462
rect 11025 21459 11081 21462
rect 11133 21459 11189 21462
rect 11241 21459 11297 21462
rect 11349 21459 11405 21462
rect 11457 21459 11481 21462
rect 1481 21447 11481 21459
rect 1481 21267 11481 21279
rect 1481 21264 1505 21267
rect 1557 21264 1613 21267
rect 1665 21264 1721 21267
rect 1773 21264 1829 21267
rect 1881 21264 1937 21267
rect 1989 21264 2045 21267
rect 2097 21264 2153 21267
rect 2205 21264 2261 21267
rect 2313 21264 2369 21267
rect 2421 21264 2477 21267
rect 2529 21264 2585 21267
rect 2637 21264 2693 21267
rect 2745 21264 2801 21267
rect 2853 21264 2909 21267
rect 2961 21264 3017 21267
rect 3069 21264 3125 21267
rect 3177 21264 3233 21267
rect 3285 21264 5372 21267
rect 5424 21264 5480 21267
rect 5532 21264 5588 21267
rect 5640 21264 5696 21267
rect 5748 21264 5804 21267
rect 5856 21264 5912 21267
rect 5964 21264 6020 21267
rect 6072 21264 6128 21267
rect 6180 21264 6236 21267
rect 6288 21264 6344 21267
rect 6396 21264 7749 21267
rect 7801 21264 7857 21267
rect 7909 21264 7965 21267
rect 8017 21264 8073 21267
rect 8125 21264 8181 21267
rect 8233 21264 8289 21267
rect 8341 21264 8397 21267
rect 8449 21264 8505 21267
rect 8557 21264 8613 21267
rect 8665 21264 8721 21267
rect 8773 21264 8829 21267
rect 8881 21264 8937 21267
rect 8989 21264 9045 21267
rect 9097 21264 9153 21267
rect 9205 21264 9261 21267
rect 9313 21264 9369 21267
rect 9421 21264 9477 21267
rect 9529 21264 11481 21267
rect 1481 21218 1494 21264
rect 11468 21218 11481 21264
rect 1481 21215 1505 21218
rect 1557 21215 1613 21218
rect 1665 21215 1721 21218
rect 1773 21215 1829 21218
rect 1881 21215 1937 21218
rect 1989 21215 2045 21218
rect 2097 21215 2153 21218
rect 2205 21215 2261 21218
rect 2313 21215 2369 21218
rect 2421 21215 2477 21218
rect 2529 21215 2585 21218
rect 2637 21215 2693 21218
rect 2745 21215 2801 21218
rect 2853 21215 2909 21218
rect 2961 21215 3017 21218
rect 3069 21215 3125 21218
rect 3177 21215 3233 21218
rect 3285 21215 5372 21218
rect 5424 21215 5480 21218
rect 5532 21215 5588 21218
rect 5640 21215 5696 21218
rect 5748 21215 5804 21218
rect 5856 21215 5912 21218
rect 5964 21215 6020 21218
rect 6072 21215 6128 21218
rect 6180 21215 6236 21218
rect 6288 21215 6344 21218
rect 6396 21215 7749 21218
rect 7801 21215 7857 21218
rect 7909 21215 7965 21218
rect 8017 21215 8073 21218
rect 8125 21215 8181 21218
rect 8233 21215 8289 21218
rect 8341 21215 8397 21218
rect 8449 21215 8505 21218
rect 8557 21215 8613 21218
rect 8665 21215 8721 21218
rect 8773 21215 8829 21218
rect 8881 21215 8937 21218
rect 8989 21215 9045 21218
rect 9097 21215 9153 21218
rect 9205 21215 9261 21218
rect 9313 21215 9369 21218
rect 9421 21215 9477 21218
rect 9529 21215 11481 21218
rect 1481 21203 11481 21215
rect 1481 21023 11481 21035
rect 1481 21020 3433 21023
rect 3485 21020 3541 21023
rect 3593 21020 3649 21023
rect 3701 21020 3757 21023
rect 3809 21020 3865 21023
rect 3917 21020 3973 21023
rect 4025 21020 4081 21023
rect 4133 21020 4189 21023
rect 4241 21020 4297 21023
rect 4349 21020 4405 21023
rect 4457 21020 4513 21023
rect 4565 21020 4621 21023
rect 4673 21020 4729 21023
rect 4781 21020 4837 21023
rect 4889 21020 4945 21023
rect 4997 21020 5053 21023
rect 5105 21020 5161 21023
rect 5213 21020 6566 21023
rect 6618 21020 6674 21023
rect 6726 21020 6782 21023
rect 6834 21020 6890 21023
rect 6942 21020 6998 21023
rect 7050 21020 7106 21023
rect 7158 21020 7214 21023
rect 7266 21020 7322 21023
rect 7374 21020 7430 21023
rect 7482 21020 7538 21023
rect 7590 21020 9677 21023
rect 9729 21020 9785 21023
rect 9837 21020 9893 21023
rect 9945 21020 10001 21023
rect 10053 21020 10109 21023
rect 10161 21020 10217 21023
rect 10269 21020 10325 21023
rect 10377 21020 10433 21023
rect 10485 21020 10541 21023
rect 10593 21020 10649 21023
rect 10701 21020 10757 21023
rect 10809 21020 10865 21023
rect 10917 21020 10973 21023
rect 11025 21020 11081 21023
rect 11133 21020 11189 21023
rect 11241 21020 11297 21023
rect 11349 21020 11405 21023
rect 11457 21020 11481 21023
rect 1481 20974 1494 21020
rect 11468 20974 11481 21020
rect 1481 20971 3433 20974
rect 3485 20971 3541 20974
rect 3593 20971 3649 20974
rect 3701 20971 3757 20974
rect 3809 20971 3865 20974
rect 3917 20971 3973 20974
rect 4025 20971 4081 20974
rect 4133 20971 4189 20974
rect 4241 20971 4297 20974
rect 4349 20971 4405 20974
rect 4457 20971 4513 20974
rect 4565 20971 4621 20974
rect 4673 20971 4729 20974
rect 4781 20971 4837 20974
rect 4889 20971 4945 20974
rect 4997 20971 5053 20974
rect 5105 20971 5161 20974
rect 5213 20971 6566 20974
rect 6618 20971 6674 20974
rect 6726 20971 6782 20974
rect 6834 20971 6890 20974
rect 6942 20971 6998 20974
rect 7050 20971 7106 20974
rect 7158 20971 7214 20974
rect 7266 20971 7322 20974
rect 7374 20971 7430 20974
rect 7482 20971 7538 20974
rect 7590 20971 9677 20974
rect 9729 20971 9785 20974
rect 9837 20971 9893 20974
rect 9945 20971 10001 20974
rect 10053 20971 10109 20974
rect 10161 20971 10217 20974
rect 10269 20971 10325 20974
rect 10377 20971 10433 20974
rect 10485 20971 10541 20974
rect 10593 20971 10649 20974
rect 10701 20971 10757 20974
rect 10809 20971 10865 20974
rect 10917 20971 10973 20974
rect 11025 20971 11081 20974
rect 11133 20971 11189 20974
rect 11241 20971 11297 20974
rect 11349 20971 11405 20974
rect 11457 20971 11481 20974
rect 1481 20959 11481 20971
rect 1481 20779 11481 20791
rect 1481 20776 1505 20779
rect 1557 20776 1613 20779
rect 1665 20776 1721 20779
rect 1773 20776 1829 20779
rect 1881 20776 1937 20779
rect 1989 20776 2045 20779
rect 2097 20776 2153 20779
rect 2205 20776 2261 20779
rect 2313 20776 2369 20779
rect 2421 20776 2477 20779
rect 2529 20776 2585 20779
rect 2637 20776 2693 20779
rect 2745 20776 2801 20779
rect 2853 20776 2909 20779
rect 2961 20776 3017 20779
rect 3069 20776 3125 20779
rect 3177 20776 3233 20779
rect 3285 20776 5372 20779
rect 5424 20776 5480 20779
rect 5532 20776 5588 20779
rect 5640 20776 5696 20779
rect 5748 20776 5804 20779
rect 5856 20776 5912 20779
rect 5964 20776 6020 20779
rect 6072 20776 6128 20779
rect 6180 20776 6236 20779
rect 6288 20776 6344 20779
rect 6396 20776 7749 20779
rect 7801 20776 7857 20779
rect 7909 20776 7965 20779
rect 8017 20776 8073 20779
rect 8125 20776 8181 20779
rect 8233 20776 8289 20779
rect 8341 20776 8397 20779
rect 8449 20776 8505 20779
rect 8557 20776 8613 20779
rect 8665 20776 8721 20779
rect 8773 20776 8829 20779
rect 8881 20776 8937 20779
rect 8989 20776 9045 20779
rect 9097 20776 9153 20779
rect 9205 20776 9261 20779
rect 9313 20776 9369 20779
rect 9421 20776 9477 20779
rect 9529 20776 11481 20779
rect 1481 20730 1494 20776
rect 11468 20730 11481 20776
rect 1481 20727 1505 20730
rect 1557 20727 1613 20730
rect 1665 20727 1721 20730
rect 1773 20727 1829 20730
rect 1881 20727 1937 20730
rect 1989 20727 2045 20730
rect 2097 20727 2153 20730
rect 2205 20727 2261 20730
rect 2313 20727 2369 20730
rect 2421 20727 2477 20730
rect 2529 20727 2585 20730
rect 2637 20727 2693 20730
rect 2745 20727 2801 20730
rect 2853 20727 2909 20730
rect 2961 20727 3017 20730
rect 3069 20727 3125 20730
rect 3177 20727 3233 20730
rect 3285 20727 5372 20730
rect 5424 20727 5480 20730
rect 5532 20727 5588 20730
rect 5640 20727 5696 20730
rect 5748 20727 5804 20730
rect 5856 20727 5912 20730
rect 5964 20727 6020 20730
rect 6072 20727 6128 20730
rect 6180 20727 6236 20730
rect 6288 20727 6344 20730
rect 6396 20727 7749 20730
rect 7801 20727 7857 20730
rect 7909 20727 7965 20730
rect 8017 20727 8073 20730
rect 8125 20727 8181 20730
rect 8233 20727 8289 20730
rect 8341 20727 8397 20730
rect 8449 20727 8505 20730
rect 8557 20727 8613 20730
rect 8665 20727 8721 20730
rect 8773 20727 8829 20730
rect 8881 20727 8937 20730
rect 8989 20727 9045 20730
rect 9097 20727 9153 20730
rect 9205 20727 9261 20730
rect 9313 20727 9369 20730
rect 9421 20727 9477 20730
rect 9529 20727 11481 20730
rect 1481 20715 11481 20727
rect 1481 20535 11481 20547
rect 1481 20532 3433 20535
rect 3485 20532 3541 20535
rect 3593 20532 3649 20535
rect 3701 20532 3757 20535
rect 3809 20532 3865 20535
rect 3917 20532 3973 20535
rect 4025 20532 4081 20535
rect 4133 20532 4189 20535
rect 4241 20532 4297 20535
rect 4349 20532 4405 20535
rect 4457 20532 4513 20535
rect 4565 20532 4621 20535
rect 4673 20532 4729 20535
rect 4781 20532 4837 20535
rect 4889 20532 4945 20535
rect 4997 20532 5053 20535
rect 5105 20532 5161 20535
rect 5213 20532 6566 20535
rect 6618 20532 6674 20535
rect 6726 20532 6782 20535
rect 6834 20532 6890 20535
rect 6942 20532 6998 20535
rect 7050 20532 7106 20535
rect 7158 20532 7214 20535
rect 7266 20532 7322 20535
rect 7374 20532 7430 20535
rect 7482 20532 7538 20535
rect 7590 20532 9677 20535
rect 9729 20532 9785 20535
rect 9837 20532 9893 20535
rect 9945 20532 10001 20535
rect 10053 20532 10109 20535
rect 10161 20532 10217 20535
rect 10269 20532 10325 20535
rect 10377 20532 10433 20535
rect 10485 20532 10541 20535
rect 10593 20532 10649 20535
rect 10701 20532 10757 20535
rect 10809 20532 10865 20535
rect 10917 20532 10973 20535
rect 11025 20532 11081 20535
rect 11133 20532 11189 20535
rect 11241 20532 11297 20535
rect 11349 20532 11405 20535
rect 11457 20532 11481 20535
rect 1481 20486 1494 20532
rect 11468 20486 11481 20532
rect 1481 20483 3433 20486
rect 3485 20483 3541 20486
rect 3593 20483 3649 20486
rect 3701 20483 3757 20486
rect 3809 20483 3865 20486
rect 3917 20483 3973 20486
rect 4025 20483 4081 20486
rect 4133 20483 4189 20486
rect 4241 20483 4297 20486
rect 4349 20483 4405 20486
rect 4457 20483 4513 20486
rect 4565 20483 4621 20486
rect 4673 20483 4729 20486
rect 4781 20483 4837 20486
rect 4889 20483 4945 20486
rect 4997 20483 5053 20486
rect 5105 20483 5161 20486
rect 5213 20483 6566 20486
rect 6618 20483 6674 20486
rect 6726 20483 6782 20486
rect 6834 20483 6890 20486
rect 6942 20483 6998 20486
rect 7050 20483 7106 20486
rect 7158 20483 7214 20486
rect 7266 20483 7322 20486
rect 7374 20483 7430 20486
rect 7482 20483 7538 20486
rect 7590 20483 9677 20486
rect 9729 20483 9785 20486
rect 9837 20483 9893 20486
rect 9945 20483 10001 20486
rect 10053 20483 10109 20486
rect 10161 20483 10217 20486
rect 10269 20483 10325 20486
rect 10377 20483 10433 20486
rect 10485 20483 10541 20486
rect 10593 20483 10649 20486
rect 10701 20483 10757 20486
rect 10809 20483 10865 20486
rect 10917 20483 10973 20486
rect 11025 20483 11081 20486
rect 11133 20483 11189 20486
rect 11241 20483 11297 20486
rect 11349 20483 11405 20486
rect 11457 20483 11481 20486
rect 1481 20471 11481 20483
rect 1481 20291 11481 20303
rect 1481 20288 1505 20291
rect 1557 20288 1613 20291
rect 1665 20288 1721 20291
rect 1773 20288 1829 20291
rect 1881 20288 1937 20291
rect 1989 20288 2045 20291
rect 2097 20288 2153 20291
rect 2205 20288 2261 20291
rect 2313 20288 2369 20291
rect 2421 20288 2477 20291
rect 2529 20288 2585 20291
rect 2637 20288 2693 20291
rect 2745 20288 2801 20291
rect 2853 20288 2909 20291
rect 2961 20288 3017 20291
rect 3069 20288 3125 20291
rect 3177 20288 3233 20291
rect 3285 20288 5372 20291
rect 5424 20288 5480 20291
rect 5532 20288 5588 20291
rect 5640 20288 5696 20291
rect 5748 20288 5804 20291
rect 5856 20288 5912 20291
rect 5964 20288 6020 20291
rect 6072 20288 6128 20291
rect 6180 20288 6236 20291
rect 6288 20288 6344 20291
rect 6396 20288 7749 20291
rect 7801 20288 7857 20291
rect 7909 20288 7965 20291
rect 8017 20288 8073 20291
rect 8125 20288 8181 20291
rect 8233 20288 8289 20291
rect 8341 20288 8397 20291
rect 8449 20288 8505 20291
rect 8557 20288 8613 20291
rect 8665 20288 8721 20291
rect 8773 20288 8829 20291
rect 8881 20288 8937 20291
rect 8989 20288 9045 20291
rect 9097 20288 9153 20291
rect 9205 20288 9261 20291
rect 9313 20288 9369 20291
rect 9421 20288 9477 20291
rect 9529 20288 11481 20291
rect 1481 20242 1494 20288
rect 11468 20242 11481 20288
rect 1481 20239 1505 20242
rect 1557 20239 1613 20242
rect 1665 20239 1721 20242
rect 1773 20239 1829 20242
rect 1881 20239 1937 20242
rect 1989 20239 2045 20242
rect 2097 20239 2153 20242
rect 2205 20239 2261 20242
rect 2313 20239 2369 20242
rect 2421 20239 2477 20242
rect 2529 20239 2585 20242
rect 2637 20239 2693 20242
rect 2745 20239 2801 20242
rect 2853 20239 2909 20242
rect 2961 20239 3017 20242
rect 3069 20239 3125 20242
rect 3177 20239 3233 20242
rect 3285 20239 5372 20242
rect 5424 20239 5480 20242
rect 5532 20239 5588 20242
rect 5640 20239 5696 20242
rect 5748 20239 5804 20242
rect 5856 20239 5912 20242
rect 5964 20239 6020 20242
rect 6072 20239 6128 20242
rect 6180 20239 6236 20242
rect 6288 20239 6344 20242
rect 6396 20239 7749 20242
rect 7801 20239 7857 20242
rect 7909 20239 7965 20242
rect 8017 20239 8073 20242
rect 8125 20239 8181 20242
rect 8233 20239 8289 20242
rect 8341 20239 8397 20242
rect 8449 20239 8505 20242
rect 8557 20239 8613 20242
rect 8665 20239 8721 20242
rect 8773 20239 8829 20242
rect 8881 20239 8937 20242
rect 8989 20239 9045 20242
rect 9097 20239 9153 20242
rect 9205 20239 9261 20242
rect 9313 20239 9369 20242
rect 9421 20239 9477 20242
rect 9529 20239 11481 20242
rect 1481 20227 11481 20239
rect 1481 20047 11481 20059
rect 1481 20044 3433 20047
rect 3485 20044 3541 20047
rect 3593 20044 3649 20047
rect 3701 20044 3757 20047
rect 3809 20044 3865 20047
rect 3917 20044 3973 20047
rect 4025 20044 4081 20047
rect 4133 20044 4189 20047
rect 4241 20044 4297 20047
rect 4349 20044 4405 20047
rect 4457 20044 4513 20047
rect 4565 20044 4621 20047
rect 4673 20044 4729 20047
rect 4781 20044 4837 20047
rect 4889 20044 4945 20047
rect 4997 20044 5053 20047
rect 5105 20044 5161 20047
rect 5213 20044 6566 20047
rect 6618 20044 6674 20047
rect 6726 20044 6782 20047
rect 6834 20044 6890 20047
rect 6942 20044 6998 20047
rect 7050 20044 7106 20047
rect 7158 20044 7214 20047
rect 7266 20044 7322 20047
rect 7374 20044 7430 20047
rect 7482 20044 7538 20047
rect 7590 20044 9677 20047
rect 9729 20044 9785 20047
rect 9837 20044 9893 20047
rect 9945 20044 10001 20047
rect 10053 20044 10109 20047
rect 10161 20044 10217 20047
rect 10269 20044 10325 20047
rect 10377 20044 10433 20047
rect 10485 20044 10541 20047
rect 10593 20044 10649 20047
rect 10701 20044 10757 20047
rect 10809 20044 10865 20047
rect 10917 20044 10973 20047
rect 11025 20044 11081 20047
rect 11133 20044 11189 20047
rect 11241 20044 11297 20047
rect 11349 20044 11405 20047
rect 11457 20044 11481 20047
rect 1481 19998 1494 20044
rect 11468 19998 11481 20044
rect 1481 19995 3433 19998
rect 3485 19995 3541 19998
rect 3593 19995 3649 19998
rect 3701 19995 3757 19998
rect 3809 19995 3865 19998
rect 3917 19995 3973 19998
rect 4025 19995 4081 19998
rect 4133 19995 4189 19998
rect 4241 19995 4297 19998
rect 4349 19995 4405 19998
rect 4457 19995 4513 19998
rect 4565 19995 4621 19998
rect 4673 19995 4729 19998
rect 4781 19995 4837 19998
rect 4889 19995 4945 19998
rect 4997 19995 5053 19998
rect 5105 19995 5161 19998
rect 5213 19995 6566 19998
rect 6618 19995 6674 19998
rect 6726 19995 6782 19998
rect 6834 19995 6890 19998
rect 6942 19995 6998 19998
rect 7050 19995 7106 19998
rect 7158 19995 7214 19998
rect 7266 19995 7322 19998
rect 7374 19995 7430 19998
rect 7482 19995 7538 19998
rect 7590 19995 9677 19998
rect 9729 19995 9785 19998
rect 9837 19995 9893 19998
rect 9945 19995 10001 19998
rect 10053 19995 10109 19998
rect 10161 19995 10217 19998
rect 10269 19995 10325 19998
rect 10377 19995 10433 19998
rect 10485 19995 10541 19998
rect 10593 19995 10649 19998
rect 10701 19995 10757 19998
rect 10809 19995 10865 19998
rect 10917 19995 10973 19998
rect 11025 19995 11081 19998
rect 11133 19995 11189 19998
rect 11241 19995 11297 19998
rect 11349 19995 11405 19998
rect 11457 19995 11481 19998
rect 1481 19983 11481 19995
rect 1481 19803 11481 19815
rect 1481 19800 1505 19803
rect 1557 19800 1613 19803
rect 1665 19800 1721 19803
rect 1773 19800 1829 19803
rect 1881 19800 1937 19803
rect 1989 19800 2045 19803
rect 2097 19800 2153 19803
rect 2205 19800 2261 19803
rect 2313 19800 2369 19803
rect 2421 19800 2477 19803
rect 2529 19800 2585 19803
rect 2637 19800 2693 19803
rect 2745 19800 2801 19803
rect 2853 19800 2909 19803
rect 2961 19800 3017 19803
rect 3069 19800 3125 19803
rect 3177 19800 3233 19803
rect 3285 19800 5372 19803
rect 5424 19800 5480 19803
rect 5532 19800 5588 19803
rect 5640 19800 5696 19803
rect 5748 19800 5804 19803
rect 5856 19800 5912 19803
rect 5964 19800 6020 19803
rect 6072 19800 6128 19803
rect 6180 19800 6236 19803
rect 6288 19800 6344 19803
rect 6396 19800 7749 19803
rect 7801 19800 7857 19803
rect 7909 19800 7965 19803
rect 8017 19800 8073 19803
rect 8125 19800 8181 19803
rect 8233 19800 8289 19803
rect 8341 19800 8397 19803
rect 8449 19800 8505 19803
rect 8557 19800 8613 19803
rect 8665 19800 8721 19803
rect 8773 19800 8829 19803
rect 8881 19800 8937 19803
rect 8989 19800 9045 19803
rect 9097 19800 9153 19803
rect 9205 19800 9261 19803
rect 9313 19800 9369 19803
rect 9421 19800 9477 19803
rect 9529 19800 11481 19803
rect 1481 19754 1494 19800
rect 11468 19754 11481 19800
rect 1481 19751 1505 19754
rect 1557 19751 1613 19754
rect 1665 19751 1721 19754
rect 1773 19751 1829 19754
rect 1881 19751 1937 19754
rect 1989 19751 2045 19754
rect 2097 19751 2153 19754
rect 2205 19751 2261 19754
rect 2313 19751 2369 19754
rect 2421 19751 2477 19754
rect 2529 19751 2585 19754
rect 2637 19751 2693 19754
rect 2745 19751 2801 19754
rect 2853 19751 2909 19754
rect 2961 19751 3017 19754
rect 3069 19751 3125 19754
rect 3177 19751 3233 19754
rect 3285 19751 5372 19754
rect 5424 19751 5480 19754
rect 5532 19751 5588 19754
rect 5640 19751 5696 19754
rect 5748 19751 5804 19754
rect 5856 19751 5912 19754
rect 5964 19751 6020 19754
rect 6072 19751 6128 19754
rect 6180 19751 6236 19754
rect 6288 19751 6344 19754
rect 6396 19751 7749 19754
rect 7801 19751 7857 19754
rect 7909 19751 7965 19754
rect 8017 19751 8073 19754
rect 8125 19751 8181 19754
rect 8233 19751 8289 19754
rect 8341 19751 8397 19754
rect 8449 19751 8505 19754
rect 8557 19751 8613 19754
rect 8665 19751 8721 19754
rect 8773 19751 8829 19754
rect 8881 19751 8937 19754
rect 8989 19751 9045 19754
rect 9097 19751 9153 19754
rect 9205 19751 9261 19754
rect 9313 19751 9369 19754
rect 9421 19751 9477 19754
rect 9529 19751 11481 19754
rect 1481 19739 11481 19751
rect 1481 19559 11481 19571
rect 1481 19556 3433 19559
rect 3485 19556 3541 19559
rect 3593 19556 3649 19559
rect 3701 19556 3757 19559
rect 3809 19556 3865 19559
rect 3917 19556 3973 19559
rect 4025 19556 4081 19559
rect 4133 19556 4189 19559
rect 4241 19556 4297 19559
rect 4349 19556 4405 19559
rect 4457 19556 4513 19559
rect 4565 19556 4621 19559
rect 4673 19556 4729 19559
rect 4781 19556 4837 19559
rect 4889 19556 4945 19559
rect 4997 19556 5053 19559
rect 5105 19556 5161 19559
rect 5213 19556 6566 19559
rect 6618 19556 6674 19559
rect 6726 19556 6782 19559
rect 6834 19556 6890 19559
rect 6942 19556 6998 19559
rect 7050 19556 7106 19559
rect 7158 19556 7214 19559
rect 7266 19556 7322 19559
rect 7374 19556 7430 19559
rect 7482 19556 7538 19559
rect 7590 19556 9677 19559
rect 9729 19556 9785 19559
rect 9837 19556 9893 19559
rect 9945 19556 10001 19559
rect 10053 19556 10109 19559
rect 10161 19556 10217 19559
rect 10269 19556 10325 19559
rect 10377 19556 10433 19559
rect 10485 19556 10541 19559
rect 10593 19556 10649 19559
rect 10701 19556 10757 19559
rect 10809 19556 10865 19559
rect 10917 19556 10973 19559
rect 11025 19556 11081 19559
rect 11133 19556 11189 19559
rect 11241 19556 11297 19559
rect 11349 19556 11405 19559
rect 11457 19556 11481 19559
rect 1481 19510 1494 19556
rect 11468 19510 11481 19556
rect 1481 19507 3433 19510
rect 3485 19507 3541 19510
rect 3593 19507 3649 19510
rect 3701 19507 3757 19510
rect 3809 19507 3865 19510
rect 3917 19507 3973 19510
rect 4025 19507 4081 19510
rect 4133 19507 4189 19510
rect 4241 19507 4297 19510
rect 4349 19507 4405 19510
rect 4457 19507 4513 19510
rect 4565 19507 4621 19510
rect 4673 19507 4729 19510
rect 4781 19507 4837 19510
rect 4889 19507 4945 19510
rect 4997 19507 5053 19510
rect 5105 19507 5161 19510
rect 5213 19507 6566 19510
rect 6618 19507 6674 19510
rect 6726 19507 6782 19510
rect 6834 19507 6890 19510
rect 6942 19507 6998 19510
rect 7050 19507 7106 19510
rect 7158 19507 7214 19510
rect 7266 19507 7322 19510
rect 7374 19507 7430 19510
rect 7482 19507 7538 19510
rect 7590 19507 9677 19510
rect 9729 19507 9785 19510
rect 9837 19507 9893 19510
rect 9945 19507 10001 19510
rect 10053 19507 10109 19510
rect 10161 19507 10217 19510
rect 10269 19507 10325 19510
rect 10377 19507 10433 19510
rect 10485 19507 10541 19510
rect 10593 19507 10649 19510
rect 10701 19507 10757 19510
rect 10809 19507 10865 19510
rect 10917 19507 10973 19510
rect 11025 19507 11081 19510
rect 11133 19507 11189 19510
rect 11241 19507 11297 19510
rect 11349 19507 11405 19510
rect 11457 19507 11481 19510
rect 1481 19495 11481 19507
rect 1481 19315 11481 19327
rect 1481 19312 1505 19315
rect 1557 19312 1613 19315
rect 1665 19312 1721 19315
rect 1773 19312 1829 19315
rect 1881 19312 1937 19315
rect 1989 19312 2045 19315
rect 2097 19312 2153 19315
rect 2205 19312 2261 19315
rect 2313 19312 2369 19315
rect 2421 19312 2477 19315
rect 2529 19312 2585 19315
rect 2637 19312 2693 19315
rect 2745 19312 2801 19315
rect 2853 19312 2909 19315
rect 2961 19312 3017 19315
rect 3069 19312 3125 19315
rect 3177 19312 3233 19315
rect 3285 19312 5372 19315
rect 5424 19312 5480 19315
rect 5532 19312 5588 19315
rect 5640 19312 5696 19315
rect 5748 19312 5804 19315
rect 5856 19312 5912 19315
rect 5964 19312 6020 19315
rect 6072 19312 6128 19315
rect 6180 19312 6236 19315
rect 6288 19312 6344 19315
rect 6396 19312 7749 19315
rect 7801 19312 7857 19315
rect 7909 19312 7965 19315
rect 8017 19312 8073 19315
rect 8125 19312 8181 19315
rect 8233 19312 8289 19315
rect 8341 19312 8397 19315
rect 8449 19312 8505 19315
rect 8557 19312 8613 19315
rect 8665 19312 8721 19315
rect 8773 19312 8829 19315
rect 8881 19312 8937 19315
rect 8989 19312 9045 19315
rect 9097 19312 9153 19315
rect 9205 19312 9261 19315
rect 9313 19312 9369 19315
rect 9421 19312 9477 19315
rect 9529 19312 11481 19315
rect 1481 19266 1494 19312
rect 11468 19266 11481 19312
rect 1481 19263 1505 19266
rect 1557 19263 1613 19266
rect 1665 19263 1721 19266
rect 1773 19263 1829 19266
rect 1881 19263 1937 19266
rect 1989 19263 2045 19266
rect 2097 19263 2153 19266
rect 2205 19263 2261 19266
rect 2313 19263 2369 19266
rect 2421 19263 2477 19266
rect 2529 19263 2585 19266
rect 2637 19263 2693 19266
rect 2745 19263 2801 19266
rect 2853 19263 2909 19266
rect 2961 19263 3017 19266
rect 3069 19263 3125 19266
rect 3177 19263 3233 19266
rect 3285 19263 5372 19266
rect 5424 19263 5480 19266
rect 5532 19263 5588 19266
rect 5640 19263 5696 19266
rect 5748 19263 5804 19266
rect 5856 19263 5912 19266
rect 5964 19263 6020 19266
rect 6072 19263 6128 19266
rect 6180 19263 6236 19266
rect 6288 19263 6344 19266
rect 6396 19263 7749 19266
rect 7801 19263 7857 19266
rect 7909 19263 7965 19266
rect 8017 19263 8073 19266
rect 8125 19263 8181 19266
rect 8233 19263 8289 19266
rect 8341 19263 8397 19266
rect 8449 19263 8505 19266
rect 8557 19263 8613 19266
rect 8665 19263 8721 19266
rect 8773 19263 8829 19266
rect 8881 19263 8937 19266
rect 8989 19263 9045 19266
rect 9097 19263 9153 19266
rect 9205 19263 9261 19266
rect 9313 19263 9369 19266
rect 9421 19263 9477 19266
rect 9529 19263 11481 19266
rect 1481 19251 11481 19263
rect 1213 19135 1413 19162
rect 1213 19083 1233 19135
rect 1285 19083 1341 19135
rect 1393 19083 1413 19135
rect 11549 19162 11560 23808
rect 11706 23779 11749 23808
rect 11729 23727 11749 23779
rect 11706 23671 11749 23727
rect 11729 23619 11749 23671
rect 11706 23563 11749 23619
rect 11729 23511 11749 23563
rect 11706 23455 11749 23511
rect 11729 23403 11749 23455
rect 11706 23347 11749 23403
rect 11729 23295 11749 23347
rect 11706 23239 11749 23295
rect 11729 23187 11749 23239
rect 11706 23131 11749 23187
rect 11729 23079 11749 23131
rect 11706 23023 11749 23079
rect 11729 22971 11749 23023
rect 11706 22915 11749 22971
rect 11729 22863 11749 22915
rect 11706 22807 11749 22863
rect 11729 22755 11749 22807
rect 11706 22699 11749 22755
rect 11729 22647 11749 22699
rect 11706 22591 11749 22647
rect 11729 22539 11749 22591
rect 11706 22483 11749 22539
rect 11729 22431 11749 22483
rect 11706 22375 11749 22431
rect 11729 22323 11749 22375
rect 11706 22267 11749 22323
rect 11729 22215 11749 22267
rect 11706 22159 11749 22215
rect 11729 22107 11749 22159
rect 11706 22051 11749 22107
rect 11729 21999 11749 22051
rect 11706 21943 11749 21999
rect 11729 21891 11749 21943
rect 11706 21835 11749 21891
rect 11729 21783 11749 21835
rect 11706 21727 11749 21783
rect 11729 21675 11749 21727
rect 11706 21619 11749 21675
rect 11729 21567 11749 21619
rect 11706 21511 11749 21567
rect 11729 21459 11749 21511
rect 11706 21403 11749 21459
rect 11729 21351 11749 21403
rect 11706 21295 11749 21351
rect 11729 21243 11749 21295
rect 11706 21187 11749 21243
rect 11729 21135 11749 21187
rect 11706 21079 11749 21135
rect 11729 21027 11749 21079
rect 11706 20971 11749 21027
rect 11729 20919 11749 20971
rect 11706 20863 11749 20919
rect 11729 20811 11749 20863
rect 11706 20755 11749 20811
rect 11729 20703 11749 20755
rect 11706 20647 11749 20703
rect 11729 20595 11749 20647
rect 11706 20539 11749 20595
rect 11729 20487 11749 20539
rect 11706 20431 11749 20487
rect 11729 20379 11749 20431
rect 11706 20323 11749 20379
rect 11729 20271 11749 20323
rect 11706 20215 11749 20271
rect 11729 20163 11749 20215
rect 11706 20107 11749 20163
rect 11729 20055 11749 20107
rect 11706 19999 11749 20055
rect 11729 19947 11749 19999
rect 11706 19891 11749 19947
rect 11729 19839 11749 19891
rect 11706 19783 11749 19839
rect 11729 19731 11749 19783
rect 11706 19675 11749 19731
rect 11729 19623 11749 19675
rect 11706 19567 11749 19623
rect 11729 19515 11749 19567
rect 11706 19459 11749 19515
rect 11729 19407 11749 19459
rect 11706 19351 11749 19407
rect 11729 19299 11749 19351
rect 11706 19243 11749 19299
rect 11729 19191 11749 19243
rect 11706 19162 11749 19191
rect 11549 19135 11749 19162
rect 11549 19083 11569 19135
rect 11621 19083 11677 19135
rect 11729 19083 11749 19135
rect 1213 18920 1413 19083
rect 1481 19071 11481 19083
rect 1481 19068 3433 19071
rect 3485 19068 3541 19071
rect 3593 19068 3649 19071
rect 3701 19068 3757 19071
rect 3809 19068 3865 19071
rect 3917 19068 3973 19071
rect 4025 19068 4081 19071
rect 4133 19068 4189 19071
rect 4241 19068 4297 19071
rect 4349 19068 4405 19071
rect 4457 19068 4513 19071
rect 4565 19068 4621 19071
rect 4673 19068 4729 19071
rect 4781 19068 4837 19071
rect 4889 19068 4945 19071
rect 4997 19068 5053 19071
rect 5105 19068 5161 19071
rect 5213 19068 6566 19071
rect 6618 19068 6674 19071
rect 6726 19068 6782 19071
rect 6834 19068 6890 19071
rect 6942 19068 6998 19071
rect 7050 19068 7106 19071
rect 7158 19068 7214 19071
rect 7266 19068 7322 19071
rect 7374 19068 7430 19071
rect 7482 19068 7538 19071
rect 7590 19068 9677 19071
rect 9729 19068 9785 19071
rect 9837 19068 9893 19071
rect 9945 19068 10001 19071
rect 10053 19068 10109 19071
rect 10161 19068 10217 19071
rect 10269 19068 10325 19071
rect 10377 19068 10433 19071
rect 10485 19068 10541 19071
rect 10593 19068 10649 19071
rect 10701 19068 10757 19071
rect 10809 19068 10865 19071
rect 10917 19068 10973 19071
rect 11025 19068 11081 19071
rect 11133 19068 11189 19071
rect 11241 19068 11297 19071
rect 11349 19068 11405 19071
rect 11457 19068 11481 19071
rect 1481 19022 1494 19068
rect 11468 19022 11481 19068
rect 1481 19019 3433 19022
rect 3485 19019 3541 19022
rect 3593 19019 3649 19022
rect 3701 19019 3757 19022
rect 3809 19019 3865 19022
rect 3917 19019 3973 19022
rect 4025 19019 4081 19022
rect 4133 19019 4189 19022
rect 4241 19019 4297 19022
rect 4349 19019 4405 19022
rect 4457 19019 4513 19022
rect 4565 19019 4621 19022
rect 4673 19019 4729 19022
rect 4781 19019 4837 19022
rect 4889 19019 4945 19022
rect 4997 19019 5053 19022
rect 5105 19019 5161 19022
rect 5213 19019 6566 19022
rect 6618 19019 6674 19022
rect 6726 19019 6782 19022
rect 6834 19019 6890 19022
rect 6942 19019 6998 19022
rect 7050 19019 7106 19022
rect 7158 19019 7214 19022
rect 7266 19019 7322 19022
rect 7374 19019 7430 19022
rect 7482 19019 7538 19022
rect 7590 19019 9677 19022
rect 9729 19019 9785 19022
rect 9837 19019 9893 19022
rect 9945 19019 10001 19022
rect 10053 19019 10109 19022
rect 10161 19019 10217 19022
rect 10269 19019 10325 19022
rect 10377 19019 10433 19022
rect 10485 19019 10541 19022
rect 10593 19019 10649 19022
rect 10701 19019 10757 19022
rect 10809 19019 10865 19022
rect 10917 19019 10973 19022
rect 11025 19019 11081 19022
rect 11133 19019 11189 19022
rect 11241 19019 11297 19022
rect 11349 19019 11405 19022
rect 11457 19019 11481 19022
rect 1481 19007 11481 19019
rect 11549 18920 11749 19083
rect 1213 18720 11749 18920
rect 12001 18641 12012 24343
rect 950 18629 12012 18641
rect 950 18622 1505 18629
rect 1557 18622 1613 18629
rect 1665 18622 1721 18629
rect 1773 18622 1829 18629
rect 1881 18622 1937 18629
rect 1989 18622 2045 18629
rect 2097 18622 2153 18629
rect 2205 18622 2261 18629
rect 2313 18622 2369 18629
rect 2421 18622 2477 18629
rect 2529 18622 2585 18629
rect 2637 18622 2693 18629
rect 2745 18622 2801 18629
rect 2853 18622 2909 18629
rect 2961 18622 3017 18629
rect 3069 18622 3125 18629
rect 3177 18622 3233 18629
rect 3285 18622 5372 18629
rect 5424 18622 5480 18629
rect 5532 18622 5588 18629
rect 5640 18622 5696 18629
rect 5748 18622 5804 18629
rect 5856 18622 5912 18629
rect 5964 18622 6020 18629
rect 6072 18622 6128 18629
rect 6180 18622 6236 18629
rect 6288 18622 6344 18629
rect 6396 18622 7749 18629
rect 7801 18622 7857 18629
rect 7909 18622 7965 18629
rect 8017 18622 8073 18629
rect 8125 18622 8181 18629
rect 8233 18622 8289 18629
rect 8341 18622 8397 18629
rect 8449 18622 8505 18629
rect 8557 18622 8613 18629
rect 8665 18622 8721 18629
rect 8773 18622 8829 18629
rect 8881 18622 8937 18629
rect 8989 18622 9045 18629
rect 9097 18622 9153 18629
rect 9205 18622 9261 18629
rect 9313 18622 9369 18629
rect 9421 18622 9477 18629
rect 9529 18622 12012 18629
rect 950 18476 1058 18622
rect 11904 18476 12012 18622
rect 950 18469 1505 18476
rect 1557 18469 1613 18476
rect 1665 18469 1721 18476
rect 1773 18469 1829 18476
rect 1881 18469 1937 18476
rect 1989 18469 2045 18476
rect 2097 18469 2153 18476
rect 2205 18469 2261 18476
rect 2313 18469 2369 18476
rect 2421 18469 2477 18476
rect 2529 18469 2585 18476
rect 2637 18469 2693 18476
rect 2745 18469 2801 18476
rect 2853 18469 2909 18476
rect 2961 18469 3017 18476
rect 3069 18469 3125 18476
rect 3177 18469 3233 18476
rect 3285 18469 5372 18476
rect 5424 18469 5480 18476
rect 5532 18469 5588 18476
rect 5640 18469 5696 18476
rect 5748 18469 5804 18476
rect 5856 18469 5912 18476
rect 5964 18469 6020 18476
rect 6072 18469 6128 18476
rect 6180 18469 6236 18476
rect 6288 18469 6344 18476
rect 6396 18469 7749 18476
rect 7801 18469 7857 18476
rect 7909 18469 7965 18476
rect 8017 18469 8073 18476
rect 8125 18469 8181 18476
rect 8233 18469 8289 18476
rect 8341 18469 8397 18476
rect 8449 18469 8505 18476
rect 8557 18469 8613 18476
rect 8665 18469 8721 18476
rect 8773 18469 8829 18476
rect 8881 18469 8937 18476
rect 8989 18469 9045 18476
rect 9097 18469 9153 18476
rect 9205 18469 9261 18476
rect 9313 18469 9369 18476
rect 9421 18469 9477 18476
rect 9529 18469 12012 18476
rect 950 18457 12012 18469
rect 950 12769 961 18457
rect 1213 18178 11749 18378
rect 1213 18015 1413 18178
rect 1481 18079 11481 18091
rect 1481 18076 3433 18079
rect 3485 18076 3541 18079
rect 3593 18076 3649 18079
rect 3701 18076 3757 18079
rect 3809 18076 3865 18079
rect 3917 18076 3973 18079
rect 4025 18076 4081 18079
rect 4133 18076 4189 18079
rect 4241 18076 4297 18079
rect 4349 18076 4405 18079
rect 4457 18076 4513 18079
rect 4565 18076 4621 18079
rect 4673 18076 4729 18079
rect 4781 18076 4837 18079
rect 4889 18076 4945 18079
rect 4997 18076 5053 18079
rect 5105 18076 5161 18079
rect 5213 18076 6566 18079
rect 6618 18076 6674 18079
rect 6726 18076 6782 18079
rect 6834 18076 6890 18079
rect 6942 18076 6998 18079
rect 7050 18076 7106 18079
rect 7158 18076 7214 18079
rect 7266 18076 7322 18079
rect 7374 18076 7430 18079
rect 7482 18076 7538 18079
rect 7590 18076 9677 18079
rect 9729 18076 9785 18079
rect 9837 18076 9893 18079
rect 9945 18076 10001 18079
rect 10053 18076 10109 18079
rect 10161 18076 10217 18079
rect 10269 18076 10325 18079
rect 10377 18076 10433 18079
rect 10485 18076 10541 18079
rect 10593 18076 10649 18079
rect 10701 18076 10757 18079
rect 10809 18076 10865 18079
rect 10917 18076 10973 18079
rect 11025 18076 11081 18079
rect 11133 18076 11189 18079
rect 11241 18076 11297 18079
rect 11349 18076 11405 18079
rect 11457 18076 11481 18079
rect 1481 18030 1494 18076
rect 11468 18030 11481 18076
rect 1481 18027 3433 18030
rect 3485 18027 3541 18030
rect 3593 18027 3649 18030
rect 3701 18027 3757 18030
rect 3809 18027 3865 18030
rect 3917 18027 3973 18030
rect 4025 18027 4081 18030
rect 4133 18027 4189 18030
rect 4241 18027 4297 18030
rect 4349 18027 4405 18030
rect 4457 18027 4513 18030
rect 4565 18027 4621 18030
rect 4673 18027 4729 18030
rect 4781 18027 4837 18030
rect 4889 18027 4945 18030
rect 4997 18027 5053 18030
rect 5105 18027 5161 18030
rect 5213 18027 6566 18030
rect 6618 18027 6674 18030
rect 6726 18027 6782 18030
rect 6834 18027 6890 18030
rect 6942 18027 6998 18030
rect 7050 18027 7106 18030
rect 7158 18027 7214 18030
rect 7266 18027 7322 18030
rect 7374 18027 7430 18030
rect 7482 18027 7538 18030
rect 7590 18027 9677 18030
rect 9729 18027 9785 18030
rect 9837 18027 9893 18030
rect 9945 18027 10001 18030
rect 10053 18027 10109 18030
rect 10161 18027 10217 18030
rect 10269 18027 10325 18030
rect 10377 18027 10433 18030
rect 10485 18027 10541 18030
rect 10593 18027 10649 18030
rect 10701 18027 10757 18030
rect 10809 18027 10865 18030
rect 10917 18027 10973 18030
rect 11025 18027 11081 18030
rect 11133 18027 11189 18030
rect 11241 18027 11297 18030
rect 11349 18027 11405 18030
rect 11457 18027 11481 18030
rect 1481 18015 11481 18027
rect 11549 18015 11749 18178
rect 1213 17963 1233 18015
rect 1285 17963 1341 18015
rect 1393 17963 1413 18015
rect 1213 17936 1413 17963
rect 1213 17907 1256 17936
rect 1213 17855 1233 17907
rect 1213 17799 1256 17855
rect 1213 17747 1233 17799
rect 1213 17691 1256 17747
rect 1213 17639 1233 17691
rect 1213 17583 1256 17639
rect 1213 17531 1233 17583
rect 1213 17475 1256 17531
rect 1213 17423 1233 17475
rect 1213 17367 1256 17423
rect 1213 17315 1233 17367
rect 1213 17259 1256 17315
rect 1213 17207 1233 17259
rect 1213 17151 1256 17207
rect 1213 17099 1233 17151
rect 1213 17043 1256 17099
rect 1213 16991 1233 17043
rect 1213 16935 1256 16991
rect 1213 16883 1233 16935
rect 1213 16827 1256 16883
rect 1213 16775 1233 16827
rect 1213 16719 1256 16775
rect 1213 16667 1233 16719
rect 1213 16611 1256 16667
rect 1213 16559 1233 16611
rect 1213 16503 1256 16559
rect 1213 16451 1233 16503
rect 1213 16395 1256 16451
rect 1213 16343 1233 16395
rect 1213 16287 1256 16343
rect 1213 16235 1233 16287
rect 1213 16179 1256 16235
rect 1213 16127 1233 16179
rect 1213 16071 1256 16127
rect 1213 16019 1233 16071
rect 1213 15963 1256 16019
rect 1213 15911 1233 15963
rect 1213 15855 1256 15911
rect 1213 15803 1233 15855
rect 1213 15747 1256 15803
rect 1213 15695 1233 15747
rect 1213 15639 1256 15695
rect 1213 15587 1233 15639
rect 1213 15531 1256 15587
rect 1213 15479 1233 15531
rect 1213 15423 1256 15479
rect 1213 15371 1233 15423
rect 1213 15315 1256 15371
rect 1213 15263 1233 15315
rect 1213 15207 1256 15263
rect 1213 15155 1233 15207
rect 1213 15099 1256 15155
rect 1213 15047 1233 15099
rect 1213 14991 1256 15047
rect 1213 14939 1233 14991
rect 1213 14883 1256 14939
rect 1213 14831 1233 14883
rect 1213 14775 1256 14831
rect 1213 14723 1233 14775
rect 1213 14667 1256 14723
rect 1213 14615 1233 14667
rect 1213 14559 1256 14615
rect 1213 14507 1233 14559
rect 1213 14451 1256 14507
rect 1213 14399 1233 14451
rect 1213 14343 1256 14399
rect 1213 14291 1233 14343
rect 1213 14235 1256 14291
rect 1213 14183 1233 14235
rect 1213 14127 1256 14183
rect 1213 14075 1233 14127
rect 1213 14019 1256 14075
rect 1213 13967 1233 14019
rect 1213 13911 1256 13967
rect 1213 13859 1233 13911
rect 1213 13803 1256 13859
rect 1213 13751 1233 13803
rect 1213 13695 1256 13751
rect 1213 13643 1233 13695
rect 1213 13587 1256 13643
rect 1213 13535 1233 13587
rect 1213 13479 1256 13535
rect 1213 13427 1233 13479
rect 1213 13371 1256 13427
rect 1213 13319 1233 13371
rect 1213 13290 1256 13319
rect 1402 13290 1413 17936
rect 11549 17963 11569 18015
rect 11621 17963 11677 18015
rect 11729 17963 11749 18015
rect 11549 17936 11749 17963
rect 1481 17835 11481 17847
rect 1481 17832 1505 17835
rect 1557 17832 1613 17835
rect 1665 17832 1721 17835
rect 1773 17832 1829 17835
rect 1881 17832 1937 17835
rect 1989 17832 2045 17835
rect 2097 17832 2153 17835
rect 2205 17832 2261 17835
rect 2313 17832 2369 17835
rect 2421 17832 2477 17835
rect 2529 17832 2585 17835
rect 2637 17832 2693 17835
rect 2745 17832 2801 17835
rect 2853 17832 2909 17835
rect 2961 17832 3017 17835
rect 3069 17832 3125 17835
rect 3177 17832 3233 17835
rect 3285 17832 5372 17835
rect 5424 17832 5480 17835
rect 5532 17832 5588 17835
rect 5640 17832 5696 17835
rect 5748 17832 5804 17835
rect 5856 17832 5912 17835
rect 5964 17832 6020 17835
rect 6072 17832 6128 17835
rect 6180 17832 6236 17835
rect 6288 17832 6344 17835
rect 6396 17832 7749 17835
rect 7801 17832 7857 17835
rect 7909 17832 7965 17835
rect 8017 17832 8073 17835
rect 8125 17832 8181 17835
rect 8233 17832 8289 17835
rect 8341 17832 8397 17835
rect 8449 17832 8505 17835
rect 8557 17832 8613 17835
rect 8665 17832 8721 17835
rect 8773 17832 8829 17835
rect 8881 17832 8937 17835
rect 8989 17832 9045 17835
rect 9097 17832 9153 17835
rect 9205 17832 9261 17835
rect 9313 17832 9369 17835
rect 9421 17832 9477 17835
rect 9529 17832 11481 17835
rect 1481 17786 1494 17832
rect 11468 17786 11481 17832
rect 1481 17783 1505 17786
rect 1557 17783 1613 17786
rect 1665 17783 1721 17786
rect 1773 17783 1829 17786
rect 1881 17783 1937 17786
rect 1989 17783 2045 17786
rect 2097 17783 2153 17786
rect 2205 17783 2261 17786
rect 2313 17783 2369 17786
rect 2421 17783 2477 17786
rect 2529 17783 2585 17786
rect 2637 17783 2693 17786
rect 2745 17783 2801 17786
rect 2853 17783 2909 17786
rect 2961 17783 3017 17786
rect 3069 17783 3125 17786
rect 3177 17783 3233 17786
rect 3285 17783 5372 17786
rect 5424 17783 5480 17786
rect 5532 17783 5588 17786
rect 5640 17783 5696 17786
rect 5748 17783 5804 17786
rect 5856 17783 5912 17786
rect 5964 17783 6020 17786
rect 6072 17783 6128 17786
rect 6180 17783 6236 17786
rect 6288 17783 6344 17786
rect 6396 17783 7749 17786
rect 7801 17783 7857 17786
rect 7909 17783 7965 17786
rect 8017 17783 8073 17786
rect 8125 17783 8181 17786
rect 8233 17783 8289 17786
rect 8341 17783 8397 17786
rect 8449 17783 8505 17786
rect 8557 17783 8613 17786
rect 8665 17783 8721 17786
rect 8773 17783 8829 17786
rect 8881 17783 8937 17786
rect 8989 17783 9045 17786
rect 9097 17783 9153 17786
rect 9205 17783 9261 17786
rect 9313 17783 9369 17786
rect 9421 17783 9477 17786
rect 9529 17783 11481 17786
rect 1481 17771 11481 17783
rect 1481 17591 11481 17603
rect 1481 17588 3433 17591
rect 3485 17588 3541 17591
rect 3593 17588 3649 17591
rect 3701 17588 3757 17591
rect 3809 17588 3865 17591
rect 3917 17588 3973 17591
rect 4025 17588 4081 17591
rect 4133 17588 4189 17591
rect 4241 17588 4297 17591
rect 4349 17588 4405 17591
rect 4457 17588 4513 17591
rect 4565 17588 4621 17591
rect 4673 17588 4729 17591
rect 4781 17588 4837 17591
rect 4889 17588 4945 17591
rect 4997 17588 5053 17591
rect 5105 17588 5161 17591
rect 5213 17588 6566 17591
rect 6618 17588 6674 17591
rect 6726 17588 6782 17591
rect 6834 17588 6890 17591
rect 6942 17588 6998 17591
rect 7050 17588 7106 17591
rect 7158 17588 7214 17591
rect 7266 17588 7322 17591
rect 7374 17588 7430 17591
rect 7482 17588 7538 17591
rect 7590 17588 9677 17591
rect 9729 17588 9785 17591
rect 9837 17588 9893 17591
rect 9945 17588 10001 17591
rect 10053 17588 10109 17591
rect 10161 17588 10217 17591
rect 10269 17588 10325 17591
rect 10377 17588 10433 17591
rect 10485 17588 10541 17591
rect 10593 17588 10649 17591
rect 10701 17588 10757 17591
rect 10809 17588 10865 17591
rect 10917 17588 10973 17591
rect 11025 17588 11081 17591
rect 11133 17588 11189 17591
rect 11241 17588 11297 17591
rect 11349 17588 11405 17591
rect 11457 17588 11481 17591
rect 1481 17542 1494 17588
rect 11468 17542 11481 17588
rect 1481 17539 3433 17542
rect 3485 17539 3541 17542
rect 3593 17539 3649 17542
rect 3701 17539 3757 17542
rect 3809 17539 3865 17542
rect 3917 17539 3973 17542
rect 4025 17539 4081 17542
rect 4133 17539 4189 17542
rect 4241 17539 4297 17542
rect 4349 17539 4405 17542
rect 4457 17539 4513 17542
rect 4565 17539 4621 17542
rect 4673 17539 4729 17542
rect 4781 17539 4837 17542
rect 4889 17539 4945 17542
rect 4997 17539 5053 17542
rect 5105 17539 5161 17542
rect 5213 17539 6566 17542
rect 6618 17539 6674 17542
rect 6726 17539 6782 17542
rect 6834 17539 6890 17542
rect 6942 17539 6998 17542
rect 7050 17539 7106 17542
rect 7158 17539 7214 17542
rect 7266 17539 7322 17542
rect 7374 17539 7430 17542
rect 7482 17539 7538 17542
rect 7590 17539 9677 17542
rect 9729 17539 9785 17542
rect 9837 17539 9893 17542
rect 9945 17539 10001 17542
rect 10053 17539 10109 17542
rect 10161 17539 10217 17542
rect 10269 17539 10325 17542
rect 10377 17539 10433 17542
rect 10485 17539 10541 17542
rect 10593 17539 10649 17542
rect 10701 17539 10757 17542
rect 10809 17539 10865 17542
rect 10917 17539 10973 17542
rect 11025 17539 11081 17542
rect 11133 17539 11189 17542
rect 11241 17539 11297 17542
rect 11349 17539 11405 17542
rect 11457 17539 11481 17542
rect 1481 17527 11481 17539
rect 1481 17347 11481 17359
rect 1481 17344 1505 17347
rect 1557 17344 1613 17347
rect 1665 17344 1721 17347
rect 1773 17344 1829 17347
rect 1881 17344 1937 17347
rect 1989 17344 2045 17347
rect 2097 17344 2153 17347
rect 2205 17344 2261 17347
rect 2313 17344 2369 17347
rect 2421 17344 2477 17347
rect 2529 17344 2585 17347
rect 2637 17344 2693 17347
rect 2745 17344 2801 17347
rect 2853 17344 2909 17347
rect 2961 17344 3017 17347
rect 3069 17344 3125 17347
rect 3177 17344 3233 17347
rect 3285 17344 5372 17347
rect 5424 17344 5480 17347
rect 5532 17344 5588 17347
rect 5640 17344 5696 17347
rect 5748 17344 5804 17347
rect 5856 17344 5912 17347
rect 5964 17344 6020 17347
rect 6072 17344 6128 17347
rect 6180 17344 6236 17347
rect 6288 17344 6344 17347
rect 6396 17344 7749 17347
rect 7801 17344 7857 17347
rect 7909 17344 7965 17347
rect 8017 17344 8073 17347
rect 8125 17344 8181 17347
rect 8233 17344 8289 17347
rect 8341 17344 8397 17347
rect 8449 17344 8505 17347
rect 8557 17344 8613 17347
rect 8665 17344 8721 17347
rect 8773 17344 8829 17347
rect 8881 17344 8937 17347
rect 8989 17344 9045 17347
rect 9097 17344 9153 17347
rect 9205 17344 9261 17347
rect 9313 17344 9369 17347
rect 9421 17344 9477 17347
rect 9529 17344 11481 17347
rect 1481 17298 1494 17344
rect 11468 17298 11481 17344
rect 1481 17295 1505 17298
rect 1557 17295 1613 17298
rect 1665 17295 1721 17298
rect 1773 17295 1829 17298
rect 1881 17295 1937 17298
rect 1989 17295 2045 17298
rect 2097 17295 2153 17298
rect 2205 17295 2261 17298
rect 2313 17295 2369 17298
rect 2421 17295 2477 17298
rect 2529 17295 2585 17298
rect 2637 17295 2693 17298
rect 2745 17295 2801 17298
rect 2853 17295 2909 17298
rect 2961 17295 3017 17298
rect 3069 17295 3125 17298
rect 3177 17295 3233 17298
rect 3285 17295 5372 17298
rect 5424 17295 5480 17298
rect 5532 17295 5588 17298
rect 5640 17295 5696 17298
rect 5748 17295 5804 17298
rect 5856 17295 5912 17298
rect 5964 17295 6020 17298
rect 6072 17295 6128 17298
rect 6180 17295 6236 17298
rect 6288 17295 6344 17298
rect 6396 17295 7749 17298
rect 7801 17295 7857 17298
rect 7909 17295 7965 17298
rect 8017 17295 8073 17298
rect 8125 17295 8181 17298
rect 8233 17295 8289 17298
rect 8341 17295 8397 17298
rect 8449 17295 8505 17298
rect 8557 17295 8613 17298
rect 8665 17295 8721 17298
rect 8773 17295 8829 17298
rect 8881 17295 8937 17298
rect 8989 17295 9045 17298
rect 9097 17295 9153 17298
rect 9205 17295 9261 17298
rect 9313 17295 9369 17298
rect 9421 17295 9477 17298
rect 9529 17295 11481 17298
rect 1481 17283 11481 17295
rect 1481 17103 11481 17115
rect 1481 17100 3433 17103
rect 3485 17100 3541 17103
rect 3593 17100 3649 17103
rect 3701 17100 3757 17103
rect 3809 17100 3865 17103
rect 3917 17100 3973 17103
rect 4025 17100 4081 17103
rect 4133 17100 4189 17103
rect 4241 17100 4297 17103
rect 4349 17100 4405 17103
rect 4457 17100 4513 17103
rect 4565 17100 4621 17103
rect 4673 17100 4729 17103
rect 4781 17100 4837 17103
rect 4889 17100 4945 17103
rect 4997 17100 5053 17103
rect 5105 17100 5161 17103
rect 5213 17100 6566 17103
rect 6618 17100 6674 17103
rect 6726 17100 6782 17103
rect 6834 17100 6890 17103
rect 6942 17100 6998 17103
rect 7050 17100 7106 17103
rect 7158 17100 7214 17103
rect 7266 17100 7322 17103
rect 7374 17100 7430 17103
rect 7482 17100 7538 17103
rect 7590 17100 9677 17103
rect 9729 17100 9785 17103
rect 9837 17100 9893 17103
rect 9945 17100 10001 17103
rect 10053 17100 10109 17103
rect 10161 17100 10217 17103
rect 10269 17100 10325 17103
rect 10377 17100 10433 17103
rect 10485 17100 10541 17103
rect 10593 17100 10649 17103
rect 10701 17100 10757 17103
rect 10809 17100 10865 17103
rect 10917 17100 10973 17103
rect 11025 17100 11081 17103
rect 11133 17100 11189 17103
rect 11241 17100 11297 17103
rect 11349 17100 11405 17103
rect 11457 17100 11481 17103
rect 1481 17054 1494 17100
rect 11468 17054 11481 17100
rect 1481 17051 3433 17054
rect 3485 17051 3541 17054
rect 3593 17051 3649 17054
rect 3701 17051 3757 17054
rect 3809 17051 3865 17054
rect 3917 17051 3973 17054
rect 4025 17051 4081 17054
rect 4133 17051 4189 17054
rect 4241 17051 4297 17054
rect 4349 17051 4405 17054
rect 4457 17051 4513 17054
rect 4565 17051 4621 17054
rect 4673 17051 4729 17054
rect 4781 17051 4837 17054
rect 4889 17051 4945 17054
rect 4997 17051 5053 17054
rect 5105 17051 5161 17054
rect 5213 17051 6566 17054
rect 6618 17051 6674 17054
rect 6726 17051 6782 17054
rect 6834 17051 6890 17054
rect 6942 17051 6998 17054
rect 7050 17051 7106 17054
rect 7158 17051 7214 17054
rect 7266 17051 7322 17054
rect 7374 17051 7430 17054
rect 7482 17051 7538 17054
rect 7590 17051 9677 17054
rect 9729 17051 9785 17054
rect 9837 17051 9893 17054
rect 9945 17051 10001 17054
rect 10053 17051 10109 17054
rect 10161 17051 10217 17054
rect 10269 17051 10325 17054
rect 10377 17051 10433 17054
rect 10485 17051 10541 17054
rect 10593 17051 10649 17054
rect 10701 17051 10757 17054
rect 10809 17051 10865 17054
rect 10917 17051 10973 17054
rect 11025 17051 11081 17054
rect 11133 17051 11189 17054
rect 11241 17051 11297 17054
rect 11349 17051 11405 17054
rect 11457 17051 11481 17054
rect 1481 17039 11481 17051
rect 1481 16859 11481 16871
rect 1481 16856 1505 16859
rect 1557 16856 1613 16859
rect 1665 16856 1721 16859
rect 1773 16856 1829 16859
rect 1881 16856 1937 16859
rect 1989 16856 2045 16859
rect 2097 16856 2153 16859
rect 2205 16856 2261 16859
rect 2313 16856 2369 16859
rect 2421 16856 2477 16859
rect 2529 16856 2585 16859
rect 2637 16856 2693 16859
rect 2745 16856 2801 16859
rect 2853 16856 2909 16859
rect 2961 16856 3017 16859
rect 3069 16856 3125 16859
rect 3177 16856 3233 16859
rect 3285 16856 5372 16859
rect 5424 16856 5480 16859
rect 5532 16856 5588 16859
rect 5640 16856 5696 16859
rect 5748 16856 5804 16859
rect 5856 16856 5912 16859
rect 5964 16856 6020 16859
rect 6072 16856 6128 16859
rect 6180 16856 6236 16859
rect 6288 16856 6344 16859
rect 6396 16856 7749 16859
rect 7801 16856 7857 16859
rect 7909 16856 7965 16859
rect 8017 16856 8073 16859
rect 8125 16856 8181 16859
rect 8233 16856 8289 16859
rect 8341 16856 8397 16859
rect 8449 16856 8505 16859
rect 8557 16856 8613 16859
rect 8665 16856 8721 16859
rect 8773 16856 8829 16859
rect 8881 16856 8937 16859
rect 8989 16856 9045 16859
rect 9097 16856 9153 16859
rect 9205 16856 9261 16859
rect 9313 16856 9369 16859
rect 9421 16856 9477 16859
rect 9529 16856 11481 16859
rect 1481 16810 1494 16856
rect 11468 16810 11481 16856
rect 1481 16807 1505 16810
rect 1557 16807 1613 16810
rect 1665 16807 1721 16810
rect 1773 16807 1829 16810
rect 1881 16807 1937 16810
rect 1989 16807 2045 16810
rect 2097 16807 2153 16810
rect 2205 16807 2261 16810
rect 2313 16807 2369 16810
rect 2421 16807 2477 16810
rect 2529 16807 2585 16810
rect 2637 16807 2693 16810
rect 2745 16807 2801 16810
rect 2853 16807 2909 16810
rect 2961 16807 3017 16810
rect 3069 16807 3125 16810
rect 3177 16807 3233 16810
rect 3285 16807 5372 16810
rect 5424 16807 5480 16810
rect 5532 16807 5588 16810
rect 5640 16807 5696 16810
rect 5748 16807 5804 16810
rect 5856 16807 5912 16810
rect 5964 16807 6020 16810
rect 6072 16807 6128 16810
rect 6180 16807 6236 16810
rect 6288 16807 6344 16810
rect 6396 16807 7749 16810
rect 7801 16807 7857 16810
rect 7909 16807 7965 16810
rect 8017 16807 8073 16810
rect 8125 16807 8181 16810
rect 8233 16807 8289 16810
rect 8341 16807 8397 16810
rect 8449 16807 8505 16810
rect 8557 16807 8613 16810
rect 8665 16807 8721 16810
rect 8773 16807 8829 16810
rect 8881 16807 8937 16810
rect 8989 16807 9045 16810
rect 9097 16807 9153 16810
rect 9205 16807 9261 16810
rect 9313 16807 9369 16810
rect 9421 16807 9477 16810
rect 9529 16807 11481 16810
rect 1481 16795 11481 16807
rect 1481 16615 11481 16627
rect 1481 16612 3433 16615
rect 3485 16612 3541 16615
rect 3593 16612 3649 16615
rect 3701 16612 3757 16615
rect 3809 16612 3865 16615
rect 3917 16612 3973 16615
rect 4025 16612 4081 16615
rect 4133 16612 4189 16615
rect 4241 16612 4297 16615
rect 4349 16612 4405 16615
rect 4457 16612 4513 16615
rect 4565 16612 4621 16615
rect 4673 16612 4729 16615
rect 4781 16612 4837 16615
rect 4889 16612 4945 16615
rect 4997 16612 5053 16615
rect 5105 16612 5161 16615
rect 5213 16612 6566 16615
rect 6618 16612 6674 16615
rect 6726 16612 6782 16615
rect 6834 16612 6890 16615
rect 6942 16612 6998 16615
rect 7050 16612 7106 16615
rect 7158 16612 7214 16615
rect 7266 16612 7322 16615
rect 7374 16612 7430 16615
rect 7482 16612 7538 16615
rect 7590 16612 9677 16615
rect 9729 16612 9785 16615
rect 9837 16612 9893 16615
rect 9945 16612 10001 16615
rect 10053 16612 10109 16615
rect 10161 16612 10217 16615
rect 10269 16612 10325 16615
rect 10377 16612 10433 16615
rect 10485 16612 10541 16615
rect 10593 16612 10649 16615
rect 10701 16612 10757 16615
rect 10809 16612 10865 16615
rect 10917 16612 10973 16615
rect 11025 16612 11081 16615
rect 11133 16612 11189 16615
rect 11241 16612 11297 16615
rect 11349 16612 11405 16615
rect 11457 16612 11481 16615
rect 1481 16566 1494 16612
rect 11468 16566 11481 16612
rect 1481 16563 3433 16566
rect 3485 16563 3541 16566
rect 3593 16563 3649 16566
rect 3701 16563 3757 16566
rect 3809 16563 3865 16566
rect 3917 16563 3973 16566
rect 4025 16563 4081 16566
rect 4133 16563 4189 16566
rect 4241 16563 4297 16566
rect 4349 16563 4405 16566
rect 4457 16563 4513 16566
rect 4565 16563 4621 16566
rect 4673 16563 4729 16566
rect 4781 16563 4837 16566
rect 4889 16563 4945 16566
rect 4997 16563 5053 16566
rect 5105 16563 5161 16566
rect 5213 16563 6566 16566
rect 6618 16563 6674 16566
rect 6726 16563 6782 16566
rect 6834 16563 6890 16566
rect 6942 16563 6998 16566
rect 7050 16563 7106 16566
rect 7158 16563 7214 16566
rect 7266 16563 7322 16566
rect 7374 16563 7430 16566
rect 7482 16563 7538 16566
rect 7590 16563 9677 16566
rect 9729 16563 9785 16566
rect 9837 16563 9893 16566
rect 9945 16563 10001 16566
rect 10053 16563 10109 16566
rect 10161 16563 10217 16566
rect 10269 16563 10325 16566
rect 10377 16563 10433 16566
rect 10485 16563 10541 16566
rect 10593 16563 10649 16566
rect 10701 16563 10757 16566
rect 10809 16563 10865 16566
rect 10917 16563 10973 16566
rect 11025 16563 11081 16566
rect 11133 16563 11189 16566
rect 11241 16563 11297 16566
rect 11349 16563 11405 16566
rect 11457 16563 11481 16566
rect 1481 16551 11481 16563
rect 1481 16371 11481 16383
rect 1481 16368 1505 16371
rect 1557 16368 1613 16371
rect 1665 16368 1721 16371
rect 1773 16368 1829 16371
rect 1881 16368 1937 16371
rect 1989 16368 2045 16371
rect 2097 16368 2153 16371
rect 2205 16368 2261 16371
rect 2313 16368 2369 16371
rect 2421 16368 2477 16371
rect 2529 16368 2585 16371
rect 2637 16368 2693 16371
rect 2745 16368 2801 16371
rect 2853 16368 2909 16371
rect 2961 16368 3017 16371
rect 3069 16368 3125 16371
rect 3177 16368 3233 16371
rect 3285 16368 5372 16371
rect 5424 16368 5480 16371
rect 5532 16368 5588 16371
rect 5640 16368 5696 16371
rect 5748 16368 5804 16371
rect 5856 16368 5912 16371
rect 5964 16368 6020 16371
rect 6072 16368 6128 16371
rect 6180 16368 6236 16371
rect 6288 16368 6344 16371
rect 6396 16368 7749 16371
rect 7801 16368 7857 16371
rect 7909 16368 7965 16371
rect 8017 16368 8073 16371
rect 8125 16368 8181 16371
rect 8233 16368 8289 16371
rect 8341 16368 8397 16371
rect 8449 16368 8505 16371
rect 8557 16368 8613 16371
rect 8665 16368 8721 16371
rect 8773 16368 8829 16371
rect 8881 16368 8937 16371
rect 8989 16368 9045 16371
rect 9097 16368 9153 16371
rect 9205 16368 9261 16371
rect 9313 16368 9369 16371
rect 9421 16368 9477 16371
rect 9529 16368 11481 16371
rect 1481 16322 1494 16368
rect 11468 16322 11481 16368
rect 1481 16319 1505 16322
rect 1557 16319 1613 16322
rect 1665 16319 1721 16322
rect 1773 16319 1829 16322
rect 1881 16319 1937 16322
rect 1989 16319 2045 16322
rect 2097 16319 2153 16322
rect 2205 16319 2261 16322
rect 2313 16319 2369 16322
rect 2421 16319 2477 16322
rect 2529 16319 2585 16322
rect 2637 16319 2693 16322
rect 2745 16319 2801 16322
rect 2853 16319 2909 16322
rect 2961 16319 3017 16322
rect 3069 16319 3125 16322
rect 3177 16319 3233 16322
rect 3285 16319 5372 16322
rect 5424 16319 5480 16322
rect 5532 16319 5588 16322
rect 5640 16319 5696 16322
rect 5748 16319 5804 16322
rect 5856 16319 5912 16322
rect 5964 16319 6020 16322
rect 6072 16319 6128 16322
rect 6180 16319 6236 16322
rect 6288 16319 6344 16322
rect 6396 16319 7749 16322
rect 7801 16319 7857 16322
rect 7909 16319 7965 16322
rect 8017 16319 8073 16322
rect 8125 16319 8181 16322
rect 8233 16319 8289 16322
rect 8341 16319 8397 16322
rect 8449 16319 8505 16322
rect 8557 16319 8613 16322
rect 8665 16319 8721 16322
rect 8773 16319 8829 16322
rect 8881 16319 8937 16322
rect 8989 16319 9045 16322
rect 9097 16319 9153 16322
rect 9205 16319 9261 16322
rect 9313 16319 9369 16322
rect 9421 16319 9477 16322
rect 9529 16319 11481 16322
rect 1481 16307 11481 16319
rect 1481 16127 11481 16139
rect 1481 16124 3433 16127
rect 3485 16124 3541 16127
rect 3593 16124 3649 16127
rect 3701 16124 3757 16127
rect 3809 16124 3865 16127
rect 3917 16124 3973 16127
rect 4025 16124 4081 16127
rect 4133 16124 4189 16127
rect 4241 16124 4297 16127
rect 4349 16124 4405 16127
rect 4457 16124 4513 16127
rect 4565 16124 4621 16127
rect 4673 16124 4729 16127
rect 4781 16124 4837 16127
rect 4889 16124 4945 16127
rect 4997 16124 5053 16127
rect 5105 16124 5161 16127
rect 5213 16124 6566 16127
rect 6618 16124 6674 16127
rect 6726 16124 6782 16127
rect 6834 16124 6890 16127
rect 6942 16124 6998 16127
rect 7050 16124 7106 16127
rect 7158 16124 7214 16127
rect 7266 16124 7322 16127
rect 7374 16124 7430 16127
rect 7482 16124 7538 16127
rect 7590 16124 9677 16127
rect 9729 16124 9785 16127
rect 9837 16124 9893 16127
rect 9945 16124 10001 16127
rect 10053 16124 10109 16127
rect 10161 16124 10217 16127
rect 10269 16124 10325 16127
rect 10377 16124 10433 16127
rect 10485 16124 10541 16127
rect 10593 16124 10649 16127
rect 10701 16124 10757 16127
rect 10809 16124 10865 16127
rect 10917 16124 10973 16127
rect 11025 16124 11081 16127
rect 11133 16124 11189 16127
rect 11241 16124 11297 16127
rect 11349 16124 11405 16127
rect 11457 16124 11481 16127
rect 1481 16078 1494 16124
rect 11468 16078 11481 16124
rect 1481 16075 3433 16078
rect 3485 16075 3541 16078
rect 3593 16075 3649 16078
rect 3701 16075 3757 16078
rect 3809 16075 3865 16078
rect 3917 16075 3973 16078
rect 4025 16075 4081 16078
rect 4133 16075 4189 16078
rect 4241 16075 4297 16078
rect 4349 16075 4405 16078
rect 4457 16075 4513 16078
rect 4565 16075 4621 16078
rect 4673 16075 4729 16078
rect 4781 16075 4837 16078
rect 4889 16075 4945 16078
rect 4997 16075 5053 16078
rect 5105 16075 5161 16078
rect 5213 16075 6566 16078
rect 6618 16075 6674 16078
rect 6726 16075 6782 16078
rect 6834 16075 6890 16078
rect 6942 16075 6998 16078
rect 7050 16075 7106 16078
rect 7158 16075 7214 16078
rect 7266 16075 7322 16078
rect 7374 16075 7430 16078
rect 7482 16075 7538 16078
rect 7590 16075 9677 16078
rect 9729 16075 9785 16078
rect 9837 16075 9893 16078
rect 9945 16075 10001 16078
rect 10053 16075 10109 16078
rect 10161 16075 10217 16078
rect 10269 16075 10325 16078
rect 10377 16075 10433 16078
rect 10485 16075 10541 16078
rect 10593 16075 10649 16078
rect 10701 16075 10757 16078
rect 10809 16075 10865 16078
rect 10917 16075 10973 16078
rect 11025 16075 11081 16078
rect 11133 16075 11189 16078
rect 11241 16075 11297 16078
rect 11349 16075 11405 16078
rect 11457 16075 11481 16078
rect 1481 16063 11481 16075
rect 1481 15883 11481 15895
rect 1481 15880 1505 15883
rect 1557 15880 1613 15883
rect 1665 15880 1721 15883
rect 1773 15880 1829 15883
rect 1881 15880 1937 15883
rect 1989 15880 2045 15883
rect 2097 15880 2153 15883
rect 2205 15880 2261 15883
rect 2313 15880 2369 15883
rect 2421 15880 2477 15883
rect 2529 15880 2585 15883
rect 2637 15880 2693 15883
rect 2745 15880 2801 15883
rect 2853 15880 2909 15883
rect 2961 15880 3017 15883
rect 3069 15880 3125 15883
rect 3177 15880 3233 15883
rect 3285 15880 5372 15883
rect 5424 15880 5480 15883
rect 5532 15880 5588 15883
rect 5640 15880 5696 15883
rect 5748 15880 5804 15883
rect 5856 15880 5912 15883
rect 5964 15880 6020 15883
rect 6072 15880 6128 15883
rect 6180 15880 6236 15883
rect 6288 15880 6344 15883
rect 6396 15880 7749 15883
rect 7801 15880 7857 15883
rect 7909 15880 7965 15883
rect 8017 15880 8073 15883
rect 8125 15880 8181 15883
rect 8233 15880 8289 15883
rect 8341 15880 8397 15883
rect 8449 15880 8505 15883
rect 8557 15880 8613 15883
rect 8665 15880 8721 15883
rect 8773 15880 8829 15883
rect 8881 15880 8937 15883
rect 8989 15880 9045 15883
rect 9097 15880 9153 15883
rect 9205 15880 9261 15883
rect 9313 15880 9369 15883
rect 9421 15880 9477 15883
rect 9529 15880 11481 15883
rect 1481 15834 1494 15880
rect 11468 15834 11481 15880
rect 1481 15831 1505 15834
rect 1557 15831 1613 15834
rect 1665 15831 1721 15834
rect 1773 15831 1829 15834
rect 1881 15831 1937 15834
rect 1989 15831 2045 15834
rect 2097 15831 2153 15834
rect 2205 15831 2261 15834
rect 2313 15831 2369 15834
rect 2421 15831 2477 15834
rect 2529 15831 2585 15834
rect 2637 15831 2693 15834
rect 2745 15831 2801 15834
rect 2853 15831 2909 15834
rect 2961 15831 3017 15834
rect 3069 15831 3125 15834
rect 3177 15831 3233 15834
rect 3285 15831 5372 15834
rect 5424 15831 5480 15834
rect 5532 15831 5588 15834
rect 5640 15831 5696 15834
rect 5748 15831 5804 15834
rect 5856 15831 5912 15834
rect 5964 15831 6020 15834
rect 6072 15831 6128 15834
rect 6180 15831 6236 15834
rect 6288 15831 6344 15834
rect 6396 15831 7749 15834
rect 7801 15831 7857 15834
rect 7909 15831 7965 15834
rect 8017 15831 8073 15834
rect 8125 15831 8181 15834
rect 8233 15831 8289 15834
rect 8341 15831 8397 15834
rect 8449 15831 8505 15834
rect 8557 15831 8613 15834
rect 8665 15831 8721 15834
rect 8773 15831 8829 15834
rect 8881 15831 8937 15834
rect 8989 15831 9045 15834
rect 9097 15831 9153 15834
rect 9205 15831 9261 15834
rect 9313 15831 9369 15834
rect 9421 15831 9477 15834
rect 9529 15831 11481 15834
rect 1481 15819 11481 15831
rect 1481 15639 11481 15651
rect 1481 15636 3433 15639
rect 3485 15636 3541 15639
rect 3593 15636 3649 15639
rect 3701 15636 3757 15639
rect 3809 15636 3865 15639
rect 3917 15636 3973 15639
rect 4025 15636 4081 15639
rect 4133 15636 4189 15639
rect 4241 15636 4297 15639
rect 4349 15636 4405 15639
rect 4457 15636 4513 15639
rect 4565 15636 4621 15639
rect 4673 15636 4729 15639
rect 4781 15636 4837 15639
rect 4889 15636 4945 15639
rect 4997 15636 5053 15639
rect 5105 15636 5161 15639
rect 5213 15636 6566 15639
rect 6618 15636 6674 15639
rect 6726 15636 6782 15639
rect 6834 15636 6890 15639
rect 6942 15636 6998 15639
rect 7050 15636 7106 15639
rect 7158 15636 7214 15639
rect 7266 15636 7322 15639
rect 7374 15636 7430 15639
rect 7482 15636 7538 15639
rect 7590 15636 9677 15639
rect 9729 15636 9785 15639
rect 9837 15636 9893 15639
rect 9945 15636 10001 15639
rect 10053 15636 10109 15639
rect 10161 15636 10217 15639
rect 10269 15636 10325 15639
rect 10377 15636 10433 15639
rect 10485 15636 10541 15639
rect 10593 15636 10649 15639
rect 10701 15636 10757 15639
rect 10809 15636 10865 15639
rect 10917 15636 10973 15639
rect 11025 15636 11081 15639
rect 11133 15636 11189 15639
rect 11241 15636 11297 15639
rect 11349 15636 11405 15639
rect 11457 15636 11481 15639
rect 1481 15590 1494 15636
rect 11468 15590 11481 15636
rect 1481 15587 3433 15590
rect 3485 15587 3541 15590
rect 3593 15587 3649 15590
rect 3701 15587 3757 15590
rect 3809 15587 3865 15590
rect 3917 15587 3973 15590
rect 4025 15587 4081 15590
rect 4133 15587 4189 15590
rect 4241 15587 4297 15590
rect 4349 15587 4405 15590
rect 4457 15587 4513 15590
rect 4565 15587 4621 15590
rect 4673 15587 4729 15590
rect 4781 15587 4837 15590
rect 4889 15587 4945 15590
rect 4997 15587 5053 15590
rect 5105 15587 5161 15590
rect 5213 15587 6566 15590
rect 6618 15587 6674 15590
rect 6726 15587 6782 15590
rect 6834 15587 6890 15590
rect 6942 15587 6998 15590
rect 7050 15587 7106 15590
rect 7158 15587 7214 15590
rect 7266 15587 7322 15590
rect 7374 15587 7430 15590
rect 7482 15587 7538 15590
rect 7590 15587 9677 15590
rect 9729 15587 9785 15590
rect 9837 15587 9893 15590
rect 9945 15587 10001 15590
rect 10053 15587 10109 15590
rect 10161 15587 10217 15590
rect 10269 15587 10325 15590
rect 10377 15587 10433 15590
rect 10485 15587 10541 15590
rect 10593 15587 10649 15590
rect 10701 15587 10757 15590
rect 10809 15587 10865 15590
rect 10917 15587 10973 15590
rect 11025 15587 11081 15590
rect 11133 15587 11189 15590
rect 11241 15587 11297 15590
rect 11349 15587 11405 15590
rect 11457 15587 11481 15590
rect 1481 15575 11481 15587
rect 1481 15395 11481 15407
rect 1481 15392 1505 15395
rect 1557 15392 1613 15395
rect 1665 15392 1721 15395
rect 1773 15392 1829 15395
rect 1881 15392 1937 15395
rect 1989 15392 2045 15395
rect 2097 15392 2153 15395
rect 2205 15392 2261 15395
rect 2313 15392 2369 15395
rect 2421 15392 2477 15395
rect 2529 15392 2585 15395
rect 2637 15392 2693 15395
rect 2745 15392 2801 15395
rect 2853 15392 2909 15395
rect 2961 15392 3017 15395
rect 3069 15392 3125 15395
rect 3177 15392 3233 15395
rect 3285 15392 5372 15395
rect 5424 15392 5480 15395
rect 5532 15392 5588 15395
rect 5640 15392 5696 15395
rect 5748 15392 5804 15395
rect 5856 15392 5912 15395
rect 5964 15392 6020 15395
rect 6072 15392 6128 15395
rect 6180 15392 6236 15395
rect 6288 15392 6344 15395
rect 6396 15392 7749 15395
rect 7801 15392 7857 15395
rect 7909 15392 7965 15395
rect 8017 15392 8073 15395
rect 8125 15392 8181 15395
rect 8233 15392 8289 15395
rect 8341 15392 8397 15395
rect 8449 15392 8505 15395
rect 8557 15392 8613 15395
rect 8665 15392 8721 15395
rect 8773 15392 8829 15395
rect 8881 15392 8937 15395
rect 8989 15392 9045 15395
rect 9097 15392 9153 15395
rect 9205 15392 9261 15395
rect 9313 15392 9369 15395
rect 9421 15392 9477 15395
rect 9529 15392 11481 15395
rect 1481 15346 1494 15392
rect 11468 15346 11481 15392
rect 1481 15343 1505 15346
rect 1557 15343 1613 15346
rect 1665 15343 1721 15346
rect 1773 15343 1829 15346
rect 1881 15343 1937 15346
rect 1989 15343 2045 15346
rect 2097 15343 2153 15346
rect 2205 15343 2261 15346
rect 2313 15343 2369 15346
rect 2421 15343 2477 15346
rect 2529 15343 2585 15346
rect 2637 15343 2693 15346
rect 2745 15343 2801 15346
rect 2853 15343 2909 15346
rect 2961 15343 3017 15346
rect 3069 15343 3125 15346
rect 3177 15343 3233 15346
rect 3285 15343 5372 15346
rect 5424 15343 5480 15346
rect 5532 15343 5588 15346
rect 5640 15343 5696 15346
rect 5748 15343 5804 15346
rect 5856 15343 5912 15346
rect 5964 15343 6020 15346
rect 6072 15343 6128 15346
rect 6180 15343 6236 15346
rect 6288 15343 6344 15346
rect 6396 15343 7749 15346
rect 7801 15343 7857 15346
rect 7909 15343 7965 15346
rect 8017 15343 8073 15346
rect 8125 15343 8181 15346
rect 8233 15343 8289 15346
rect 8341 15343 8397 15346
rect 8449 15343 8505 15346
rect 8557 15343 8613 15346
rect 8665 15343 8721 15346
rect 8773 15343 8829 15346
rect 8881 15343 8937 15346
rect 8989 15343 9045 15346
rect 9097 15343 9153 15346
rect 9205 15343 9261 15346
rect 9313 15343 9369 15346
rect 9421 15343 9477 15346
rect 9529 15343 11481 15346
rect 1481 15331 11481 15343
rect 1481 15151 11481 15163
rect 1481 15148 3433 15151
rect 3485 15148 3541 15151
rect 3593 15148 3649 15151
rect 3701 15148 3757 15151
rect 3809 15148 3865 15151
rect 3917 15148 3973 15151
rect 4025 15148 4081 15151
rect 4133 15148 4189 15151
rect 4241 15148 4297 15151
rect 4349 15148 4405 15151
rect 4457 15148 4513 15151
rect 4565 15148 4621 15151
rect 4673 15148 4729 15151
rect 4781 15148 4837 15151
rect 4889 15148 4945 15151
rect 4997 15148 5053 15151
rect 5105 15148 5161 15151
rect 5213 15148 6566 15151
rect 6618 15148 6674 15151
rect 6726 15148 6782 15151
rect 6834 15148 6890 15151
rect 6942 15148 6998 15151
rect 7050 15148 7106 15151
rect 7158 15148 7214 15151
rect 7266 15148 7322 15151
rect 7374 15148 7430 15151
rect 7482 15148 7538 15151
rect 7590 15148 9677 15151
rect 9729 15148 9785 15151
rect 9837 15148 9893 15151
rect 9945 15148 10001 15151
rect 10053 15148 10109 15151
rect 10161 15148 10217 15151
rect 10269 15148 10325 15151
rect 10377 15148 10433 15151
rect 10485 15148 10541 15151
rect 10593 15148 10649 15151
rect 10701 15148 10757 15151
rect 10809 15148 10865 15151
rect 10917 15148 10973 15151
rect 11025 15148 11081 15151
rect 11133 15148 11189 15151
rect 11241 15148 11297 15151
rect 11349 15148 11405 15151
rect 11457 15148 11481 15151
rect 1481 15102 1494 15148
rect 11468 15102 11481 15148
rect 1481 15099 3433 15102
rect 3485 15099 3541 15102
rect 3593 15099 3649 15102
rect 3701 15099 3757 15102
rect 3809 15099 3865 15102
rect 3917 15099 3973 15102
rect 4025 15099 4081 15102
rect 4133 15099 4189 15102
rect 4241 15099 4297 15102
rect 4349 15099 4405 15102
rect 4457 15099 4513 15102
rect 4565 15099 4621 15102
rect 4673 15099 4729 15102
rect 4781 15099 4837 15102
rect 4889 15099 4945 15102
rect 4997 15099 5053 15102
rect 5105 15099 5161 15102
rect 5213 15099 6566 15102
rect 6618 15099 6674 15102
rect 6726 15099 6782 15102
rect 6834 15099 6890 15102
rect 6942 15099 6998 15102
rect 7050 15099 7106 15102
rect 7158 15099 7214 15102
rect 7266 15099 7322 15102
rect 7374 15099 7430 15102
rect 7482 15099 7538 15102
rect 7590 15099 9677 15102
rect 9729 15099 9785 15102
rect 9837 15099 9893 15102
rect 9945 15099 10001 15102
rect 10053 15099 10109 15102
rect 10161 15099 10217 15102
rect 10269 15099 10325 15102
rect 10377 15099 10433 15102
rect 10485 15099 10541 15102
rect 10593 15099 10649 15102
rect 10701 15099 10757 15102
rect 10809 15099 10865 15102
rect 10917 15099 10973 15102
rect 11025 15099 11081 15102
rect 11133 15099 11189 15102
rect 11241 15099 11297 15102
rect 11349 15099 11405 15102
rect 11457 15099 11481 15102
rect 1481 15087 11481 15099
rect 1481 14907 11481 14919
rect 1481 14904 1505 14907
rect 1557 14904 1613 14907
rect 1665 14904 1721 14907
rect 1773 14904 1829 14907
rect 1881 14904 1937 14907
rect 1989 14904 2045 14907
rect 2097 14904 2153 14907
rect 2205 14904 2261 14907
rect 2313 14904 2369 14907
rect 2421 14904 2477 14907
rect 2529 14904 2585 14907
rect 2637 14904 2693 14907
rect 2745 14904 2801 14907
rect 2853 14904 2909 14907
rect 2961 14904 3017 14907
rect 3069 14904 3125 14907
rect 3177 14904 3233 14907
rect 3285 14904 5372 14907
rect 5424 14904 5480 14907
rect 5532 14904 5588 14907
rect 5640 14904 5696 14907
rect 5748 14904 5804 14907
rect 5856 14904 5912 14907
rect 5964 14904 6020 14907
rect 6072 14904 6128 14907
rect 6180 14904 6236 14907
rect 6288 14904 6344 14907
rect 6396 14904 7749 14907
rect 7801 14904 7857 14907
rect 7909 14904 7965 14907
rect 8017 14904 8073 14907
rect 8125 14904 8181 14907
rect 8233 14904 8289 14907
rect 8341 14904 8397 14907
rect 8449 14904 8505 14907
rect 8557 14904 8613 14907
rect 8665 14904 8721 14907
rect 8773 14904 8829 14907
rect 8881 14904 8937 14907
rect 8989 14904 9045 14907
rect 9097 14904 9153 14907
rect 9205 14904 9261 14907
rect 9313 14904 9369 14907
rect 9421 14904 9477 14907
rect 9529 14904 11481 14907
rect 1481 14858 1494 14904
rect 11468 14858 11481 14904
rect 1481 14855 1505 14858
rect 1557 14855 1613 14858
rect 1665 14855 1721 14858
rect 1773 14855 1829 14858
rect 1881 14855 1937 14858
rect 1989 14855 2045 14858
rect 2097 14855 2153 14858
rect 2205 14855 2261 14858
rect 2313 14855 2369 14858
rect 2421 14855 2477 14858
rect 2529 14855 2585 14858
rect 2637 14855 2693 14858
rect 2745 14855 2801 14858
rect 2853 14855 2909 14858
rect 2961 14855 3017 14858
rect 3069 14855 3125 14858
rect 3177 14855 3233 14858
rect 3285 14855 5372 14858
rect 5424 14855 5480 14858
rect 5532 14855 5588 14858
rect 5640 14855 5696 14858
rect 5748 14855 5804 14858
rect 5856 14855 5912 14858
rect 5964 14855 6020 14858
rect 6072 14855 6128 14858
rect 6180 14855 6236 14858
rect 6288 14855 6344 14858
rect 6396 14855 7749 14858
rect 7801 14855 7857 14858
rect 7909 14855 7965 14858
rect 8017 14855 8073 14858
rect 8125 14855 8181 14858
rect 8233 14855 8289 14858
rect 8341 14855 8397 14858
rect 8449 14855 8505 14858
rect 8557 14855 8613 14858
rect 8665 14855 8721 14858
rect 8773 14855 8829 14858
rect 8881 14855 8937 14858
rect 8989 14855 9045 14858
rect 9097 14855 9153 14858
rect 9205 14855 9261 14858
rect 9313 14855 9369 14858
rect 9421 14855 9477 14858
rect 9529 14855 11481 14858
rect 1481 14843 11481 14855
rect 1481 14663 11481 14675
rect 1481 14660 3433 14663
rect 3485 14660 3541 14663
rect 3593 14660 3649 14663
rect 3701 14660 3757 14663
rect 3809 14660 3865 14663
rect 3917 14660 3973 14663
rect 4025 14660 4081 14663
rect 4133 14660 4189 14663
rect 4241 14660 4297 14663
rect 4349 14660 4405 14663
rect 4457 14660 4513 14663
rect 4565 14660 4621 14663
rect 4673 14660 4729 14663
rect 4781 14660 4837 14663
rect 4889 14660 4945 14663
rect 4997 14660 5053 14663
rect 5105 14660 5161 14663
rect 5213 14660 6566 14663
rect 6618 14660 6674 14663
rect 6726 14660 6782 14663
rect 6834 14660 6890 14663
rect 6942 14660 6998 14663
rect 7050 14660 7106 14663
rect 7158 14660 7214 14663
rect 7266 14660 7322 14663
rect 7374 14660 7430 14663
rect 7482 14660 7538 14663
rect 7590 14660 9677 14663
rect 9729 14660 9785 14663
rect 9837 14660 9893 14663
rect 9945 14660 10001 14663
rect 10053 14660 10109 14663
rect 10161 14660 10217 14663
rect 10269 14660 10325 14663
rect 10377 14660 10433 14663
rect 10485 14660 10541 14663
rect 10593 14660 10649 14663
rect 10701 14660 10757 14663
rect 10809 14660 10865 14663
rect 10917 14660 10973 14663
rect 11025 14660 11081 14663
rect 11133 14660 11189 14663
rect 11241 14660 11297 14663
rect 11349 14660 11405 14663
rect 11457 14660 11481 14663
rect 1481 14614 1494 14660
rect 11468 14614 11481 14660
rect 1481 14611 3433 14614
rect 3485 14611 3541 14614
rect 3593 14611 3649 14614
rect 3701 14611 3757 14614
rect 3809 14611 3865 14614
rect 3917 14611 3973 14614
rect 4025 14611 4081 14614
rect 4133 14611 4189 14614
rect 4241 14611 4297 14614
rect 4349 14611 4405 14614
rect 4457 14611 4513 14614
rect 4565 14611 4621 14614
rect 4673 14611 4729 14614
rect 4781 14611 4837 14614
rect 4889 14611 4945 14614
rect 4997 14611 5053 14614
rect 5105 14611 5161 14614
rect 5213 14611 6566 14614
rect 6618 14611 6674 14614
rect 6726 14611 6782 14614
rect 6834 14611 6890 14614
rect 6942 14611 6998 14614
rect 7050 14611 7106 14614
rect 7158 14611 7214 14614
rect 7266 14611 7322 14614
rect 7374 14611 7430 14614
rect 7482 14611 7538 14614
rect 7590 14611 9677 14614
rect 9729 14611 9785 14614
rect 9837 14611 9893 14614
rect 9945 14611 10001 14614
rect 10053 14611 10109 14614
rect 10161 14611 10217 14614
rect 10269 14611 10325 14614
rect 10377 14611 10433 14614
rect 10485 14611 10541 14614
rect 10593 14611 10649 14614
rect 10701 14611 10757 14614
rect 10809 14611 10865 14614
rect 10917 14611 10973 14614
rect 11025 14611 11081 14614
rect 11133 14611 11189 14614
rect 11241 14611 11297 14614
rect 11349 14611 11405 14614
rect 11457 14611 11481 14614
rect 1481 14599 11481 14611
rect 1481 14419 11481 14431
rect 1481 14416 1505 14419
rect 1557 14416 1613 14419
rect 1665 14416 1721 14419
rect 1773 14416 1829 14419
rect 1881 14416 1937 14419
rect 1989 14416 2045 14419
rect 2097 14416 2153 14419
rect 2205 14416 2261 14419
rect 2313 14416 2369 14419
rect 2421 14416 2477 14419
rect 2529 14416 2585 14419
rect 2637 14416 2693 14419
rect 2745 14416 2801 14419
rect 2853 14416 2909 14419
rect 2961 14416 3017 14419
rect 3069 14416 3125 14419
rect 3177 14416 3233 14419
rect 3285 14416 5372 14419
rect 5424 14416 5480 14419
rect 5532 14416 5588 14419
rect 5640 14416 5696 14419
rect 5748 14416 5804 14419
rect 5856 14416 5912 14419
rect 5964 14416 6020 14419
rect 6072 14416 6128 14419
rect 6180 14416 6236 14419
rect 6288 14416 6344 14419
rect 6396 14416 7749 14419
rect 7801 14416 7857 14419
rect 7909 14416 7965 14419
rect 8017 14416 8073 14419
rect 8125 14416 8181 14419
rect 8233 14416 8289 14419
rect 8341 14416 8397 14419
rect 8449 14416 8505 14419
rect 8557 14416 8613 14419
rect 8665 14416 8721 14419
rect 8773 14416 8829 14419
rect 8881 14416 8937 14419
rect 8989 14416 9045 14419
rect 9097 14416 9153 14419
rect 9205 14416 9261 14419
rect 9313 14416 9369 14419
rect 9421 14416 9477 14419
rect 9529 14416 11481 14419
rect 1481 14370 1494 14416
rect 11468 14370 11481 14416
rect 1481 14367 1505 14370
rect 1557 14367 1613 14370
rect 1665 14367 1721 14370
rect 1773 14367 1829 14370
rect 1881 14367 1937 14370
rect 1989 14367 2045 14370
rect 2097 14367 2153 14370
rect 2205 14367 2261 14370
rect 2313 14367 2369 14370
rect 2421 14367 2477 14370
rect 2529 14367 2585 14370
rect 2637 14367 2693 14370
rect 2745 14367 2801 14370
rect 2853 14367 2909 14370
rect 2961 14367 3017 14370
rect 3069 14367 3125 14370
rect 3177 14367 3233 14370
rect 3285 14367 5372 14370
rect 5424 14367 5480 14370
rect 5532 14367 5588 14370
rect 5640 14367 5696 14370
rect 5748 14367 5804 14370
rect 5856 14367 5912 14370
rect 5964 14367 6020 14370
rect 6072 14367 6128 14370
rect 6180 14367 6236 14370
rect 6288 14367 6344 14370
rect 6396 14367 7749 14370
rect 7801 14367 7857 14370
rect 7909 14367 7965 14370
rect 8017 14367 8073 14370
rect 8125 14367 8181 14370
rect 8233 14367 8289 14370
rect 8341 14367 8397 14370
rect 8449 14367 8505 14370
rect 8557 14367 8613 14370
rect 8665 14367 8721 14370
rect 8773 14367 8829 14370
rect 8881 14367 8937 14370
rect 8989 14367 9045 14370
rect 9097 14367 9153 14370
rect 9205 14367 9261 14370
rect 9313 14367 9369 14370
rect 9421 14367 9477 14370
rect 9529 14367 11481 14370
rect 1481 14355 11481 14367
rect 1481 14175 11481 14187
rect 1481 14172 3433 14175
rect 3485 14172 3541 14175
rect 3593 14172 3649 14175
rect 3701 14172 3757 14175
rect 3809 14172 3865 14175
rect 3917 14172 3973 14175
rect 4025 14172 4081 14175
rect 4133 14172 4189 14175
rect 4241 14172 4297 14175
rect 4349 14172 4405 14175
rect 4457 14172 4513 14175
rect 4565 14172 4621 14175
rect 4673 14172 4729 14175
rect 4781 14172 4837 14175
rect 4889 14172 4945 14175
rect 4997 14172 5053 14175
rect 5105 14172 5161 14175
rect 5213 14172 6566 14175
rect 6618 14172 6674 14175
rect 6726 14172 6782 14175
rect 6834 14172 6890 14175
rect 6942 14172 6998 14175
rect 7050 14172 7106 14175
rect 7158 14172 7214 14175
rect 7266 14172 7322 14175
rect 7374 14172 7430 14175
rect 7482 14172 7538 14175
rect 7590 14172 9677 14175
rect 9729 14172 9785 14175
rect 9837 14172 9893 14175
rect 9945 14172 10001 14175
rect 10053 14172 10109 14175
rect 10161 14172 10217 14175
rect 10269 14172 10325 14175
rect 10377 14172 10433 14175
rect 10485 14172 10541 14175
rect 10593 14172 10649 14175
rect 10701 14172 10757 14175
rect 10809 14172 10865 14175
rect 10917 14172 10973 14175
rect 11025 14172 11081 14175
rect 11133 14172 11189 14175
rect 11241 14172 11297 14175
rect 11349 14172 11405 14175
rect 11457 14172 11481 14175
rect 1481 14126 1494 14172
rect 11468 14126 11481 14172
rect 1481 14123 3433 14126
rect 3485 14123 3541 14126
rect 3593 14123 3649 14126
rect 3701 14123 3757 14126
rect 3809 14123 3865 14126
rect 3917 14123 3973 14126
rect 4025 14123 4081 14126
rect 4133 14123 4189 14126
rect 4241 14123 4297 14126
rect 4349 14123 4405 14126
rect 4457 14123 4513 14126
rect 4565 14123 4621 14126
rect 4673 14123 4729 14126
rect 4781 14123 4837 14126
rect 4889 14123 4945 14126
rect 4997 14123 5053 14126
rect 5105 14123 5161 14126
rect 5213 14123 6566 14126
rect 6618 14123 6674 14126
rect 6726 14123 6782 14126
rect 6834 14123 6890 14126
rect 6942 14123 6998 14126
rect 7050 14123 7106 14126
rect 7158 14123 7214 14126
rect 7266 14123 7322 14126
rect 7374 14123 7430 14126
rect 7482 14123 7538 14126
rect 7590 14123 9677 14126
rect 9729 14123 9785 14126
rect 9837 14123 9893 14126
rect 9945 14123 10001 14126
rect 10053 14123 10109 14126
rect 10161 14123 10217 14126
rect 10269 14123 10325 14126
rect 10377 14123 10433 14126
rect 10485 14123 10541 14126
rect 10593 14123 10649 14126
rect 10701 14123 10757 14126
rect 10809 14123 10865 14126
rect 10917 14123 10973 14126
rect 11025 14123 11081 14126
rect 11133 14123 11189 14126
rect 11241 14123 11297 14126
rect 11349 14123 11405 14126
rect 11457 14123 11481 14126
rect 1481 14111 11481 14123
rect 1481 13931 11481 13943
rect 1481 13928 1505 13931
rect 1557 13928 1613 13931
rect 1665 13928 1721 13931
rect 1773 13928 1829 13931
rect 1881 13928 1937 13931
rect 1989 13928 2045 13931
rect 2097 13928 2153 13931
rect 2205 13928 2261 13931
rect 2313 13928 2369 13931
rect 2421 13928 2477 13931
rect 2529 13928 2585 13931
rect 2637 13928 2693 13931
rect 2745 13928 2801 13931
rect 2853 13928 2909 13931
rect 2961 13928 3017 13931
rect 3069 13928 3125 13931
rect 3177 13928 3233 13931
rect 3285 13928 5372 13931
rect 5424 13928 5480 13931
rect 5532 13928 5588 13931
rect 5640 13928 5696 13931
rect 5748 13928 5804 13931
rect 5856 13928 5912 13931
rect 5964 13928 6020 13931
rect 6072 13928 6128 13931
rect 6180 13928 6236 13931
rect 6288 13928 6344 13931
rect 6396 13928 7749 13931
rect 7801 13928 7857 13931
rect 7909 13928 7965 13931
rect 8017 13928 8073 13931
rect 8125 13928 8181 13931
rect 8233 13928 8289 13931
rect 8341 13928 8397 13931
rect 8449 13928 8505 13931
rect 8557 13928 8613 13931
rect 8665 13928 8721 13931
rect 8773 13928 8829 13931
rect 8881 13928 8937 13931
rect 8989 13928 9045 13931
rect 9097 13928 9153 13931
rect 9205 13928 9261 13931
rect 9313 13928 9369 13931
rect 9421 13928 9477 13931
rect 9529 13928 11481 13931
rect 1481 13882 1494 13928
rect 11468 13882 11481 13928
rect 1481 13879 1505 13882
rect 1557 13879 1613 13882
rect 1665 13879 1721 13882
rect 1773 13879 1829 13882
rect 1881 13879 1937 13882
rect 1989 13879 2045 13882
rect 2097 13879 2153 13882
rect 2205 13879 2261 13882
rect 2313 13879 2369 13882
rect 2421 13879 2477 13882
rect 2529 13879 2585 13882
rect 2637 13879 2693 13882
rect 2745 13879 2801 13882
rect 2853 13879 2909 13882
rect 2961 13879 3017 13882
rect 3069 13879 3125 13882
rect 3177 13879 3233 13882
rect 3285 13879 5372 13882
rect 5424 13879 5480 13882
rect 5532 13879 5588 13882
rect 5640 13879 5696 13882
rect 5748 13879 5804 13882
rect 5856 13879 5912 13882
rect 5964 13879 6020 13882
rect 6072 13879 6128 13882
rect 6180 13879 6236 13882
rect 6288 13879 6344 13882
rect 6396 13879 7749 13882
rect 7801 13879 7857 13882
rect 7909 13879 7965 13882
rect 8017 13879 8073 13882
rect 8125 13879 8181 13882
rect 8233 13879 8289 13882
rect 8341 13879 8397 13882
rect 8449 13879 8505 13882
rect 8557 13879 8613 13882
rect 8665 13879 8721 13882
rect 8773 13879 8829 13882
rect 8881 13879 8937 13882
rect 8989 13879 9045 13882
rect 9097 13879 9153 13882
rect 9205 13879 9261 13882
rect 9313 13879 9369 13882
rect 9421 13879 9477 13882
rect 9529 13879 11481 13882
rect 1481 13867 11481 13879
rect 1481 13687 11481 13699
rect 1481 13684 3433 13687
rect 3485 13684 3541 13687
rect 3593 13684 3649 13687
rect 3701 13684 3757 13687
rect 3809 13684 3865 13687
rect 3917 13684 3973 13687
rect 4025 13684 4081 13687
rect 4133 13684 4189 13687
rect 4241 13684 4297 13687
rect 4349 13684 4405 13687
rect 4457 13684 4513 13687
rect 4565 13684 4621 13687
rect 4673 13684 4729 13687
rect 4781 13684 4837 13687
rect 4889 13684 4945 13687
rect 4997 13684 5053 13687
rect 5105 13684 5161 13687
rect 5213 13684 6566 13687
rect 6618 13684 6674 13687
rect 6726 13684 6782 13687
rect 6834 13684 6890 13687
rect 6942 13684 6998 13687
rect 7050 13684 7106 13687
rect 7158 13684 7214 13687
rect 7266 13684 7322 13687
rect 7374 13684 7430 13687
rect 7482 13684 7538 13687
rect 7590 13684 9677 13687
rect 9729 13684 9785 13687
rect 9837 13684 9893 13687
rect 9945 13684 10001 13687
rect 10053 13684 10109 13687
rect 10161 13684 10217 13687
rect 10269 13684 10325 13687
rect 10377 13684 10433 13687
rect 10485 13684 10541 13687
rect 10593 13684 10649 13687
rect 10701 13684 10757 13687
rect 10809 13684 10865 13687
rect 10917 13684 10973 13687
rect 11025 13684 11081 13687
rect 11133 13684 11189 13687
rect 11241 13684 11297 13687
rect 11349 13684 11405 13687
rect 11457 13684 11481 13687
rect 1481 13638 1494 13684
rect 11468 13638 11481 13684
rect 1481 13635 3433 13638
rect 3485 13635 3541 13638
rect 3593 13635 3649 13638
rect 3701 13635 3757 13638
rect 3809 13635 3865 13638
rect 3917 13635 3973 13638
rect 4025 13635 4081 13638
rect 4133 13635 4189 13638
rect 4241 13635 4297 13638
rect 4349 13635 4405 13638
rect 4457 13635 4513 13638
rect 4565 13635 4621 13638
rect 4673 13635 4729 13638
rect 4781 13635 4837 13638
rect 4889 13635 4945 13638
rect 4997 13635 5053 13638
rect 5105 13635 5161 13638
rect 5213 13635 6566 13638
rect 6618 13635 6674 13638
rect 6726 13635 6782 13638
rect 6834 13635 6890 13638
rect 6942 13635 6998 13638
rect 7050 13635 7106 13638
rect 7158 13635 7214 13638
rect 7266 13635 7322 13638
rect 7374 13635 7430 13638
rect 7482 13635 7538 13638
rect 7590 13635 9677 13638
rect 9729 13635 9785 13638
rect 9837 13635 9893 13638
rect 9945 13635 10001 13638
rect 10053 13635 10109 13638
rect 10161 13635 10217 13638
rect 10269 13635 10325 13638
rect 10377 13635 10433 13638
rect 10485 13635 10541 13638
rect 10593 13635 10649 13638
rect 10701 13635 10757 13638
rect 10809 13635 10865 13638
rect 10917 13635 10973 13638
rect 11025 13635 11081 13638
rect 11133 13635 11189 13638
rect 11241 13635 11297 13638
rect 11349 13635 11405 13638
rect 11457 13635 11481 13638
rect 1481 13623 11481 13635
rect 1481 13443 11481 13455
rect 1481 13440 1505 13443
rect 1557 13440 1613 13443
rect 1665 13440 1721 13443
rect 1773 13440 1829 13443
rect 1881 13440 1937 13443
rect 1989 13440 2045 13443
rect 2097 13440 2153 13443
rect 2205 13440 2261 13443
rect 2313 13440 2369 13443
rect 2421 13440 2477 13443
rect 2529 13440 2585 13443
rect 2637 13440 2693 13443
rect 2745 13440 2801 13443
rect 2853 13440 2909 13443
rect 2961 13440 3017 13443
rect 3069 13440 3125 13443
rect 3177 13440 3233 13443
rect 3285 13440 5372 13443
rect 5424 13440 5480 13443
rect 5532 13440 5588 13443
rect 5640 13440 5696 13443
rect 5748 13440 5804 13443
rect 5856 13440 5912 13443
rect 5964 13440 6020 13443
rect 6072 13440 6128 13443
rect 6180 13440 6236 13443
rect 6288 13440 6344 13443
rect 6396 13440 7749 13443
rect 7801 13440 7857 13443
rect 7909 13440 7965 13443
rect 8017 13440 8073 13443
rect 8125 13440 8181 13443
rect 8233 13440 8289 13443
rect 8341 13440 8397 13443
rect 8449 13440 8505 13443
rect 8557 13440 8613 13443
rect 8665 13440 8721 13443
rect 8773 13440 8829 13443
rect 8881 13440 8937 13443
rect 8989 13440 9045 13443
rect 9097 13440 9153 13443
rect 9205 13440 9261 13443
rect 9313 13440 9369 13443
rect 9421 13440 9477 13443
rect 9529 13440 11481 13443
rect 1481 13394 1494 13440
rect 11468 13394 11481 13440
rect 1481 13391 1505 13394
rect 1557 13391 1613 13394
rect 1665 13391 1721 13394
rect 1773 13391 1829 13394
rect 1881 13391 1937 13394
rect 1989 13391 2045 13394
rect 2097 13391 2153 13394
rect 2205 13391 2261 13394
rect 2313 13391 2369 13394
rect 2421 13391 2477 13394
rect 2529 13391 2585 13394
rect 2637 13391 2693 13394
rect 2745 13391 2801 13394
rect 2853 13391 2909 13394
rect 2961 13391 3017 13394
rect 3069 13391 3125 13394
rect 3177 13391 3233 13394
rect 3285 13391 5372 13394
rect 5424 13391 5480 13394
rect 5532 13391 5588 13394
rect 5640 13391 5696 13394
rect 5748 13391 5804 13394
rect 5856 13391 5912 13394
rect 5964 13391 6020 13394
rect 6072 13391 6128 13394
rect 6180 13391 6236 13394
rect 6288 13391 6344 13394
rect 6396 13391 7749 13394
rect 7801 13391 7857 13394
rect 7909 13391 7965 13394
rect 8017 13391 8073 13394
rect 8125 13391 8181 13394
rect 8233 13391 8289 13394
rect 8341 13391 8397 13394
rect 8449 13391 8505 13394
rect 8557 13391 8613 13394
rect 8665 13391 8721 13394
rect 8773 13391 8829 13394
rect 8881 13391 8937 13394
rect 8989 13391 9045 13394
rect 9097 13391 9153 13394
rect 9205 13391 9261 13394
rect 9313 13391 9369 13394
rect 9421 13391 9477 13394
rect 9529 13391 11481 13394
rect 1481 13379 11481 13391
rect 1213 13263 1413 13290
rect 1213 13211 1233 13263
rect 1285 13211 1341 13263
rect 1393 13211 1413 13263
rect 11549 13290 11560 17936
rect 11706 17907 11749 17936
rect 11729 17855 11749 17907
rect 11706 17799 11749 17855
rect 11729 17747 11749 17799
rect 11706 17691 11749 17747
rect 11729 17639 11749 17691
rect 11706 17583 11749 17639
rect 11729 17531 11749 17583
rect 11706 17475 11749 17531
rect 11729 17423 11749 17475
rect 11706 17367 11749 17423
rect 11729 17315 11749 17367
rect 11706 17259 11749 17315
rect 11729 17207 11749 17259
rect 11706 17151 11749 17207
rect 11729 17099 11749 17151
rect 11706 17043 11749 17099
rect 11729 16991 11749 17043
rect 11706 16935 11749 16991
rect 11729 16883 11749 16935
rect 11706 16827 11749 16883
rect 11729 16775 11749 16827
rect 11706 16719 11749 16775
rect 11729 16667 11749 16719
rect 11706 16611 11749 16667
rect 11729 16559 11749 16611
rect 11706 16503 11749 16559
rect 11729 16451 11749 16503
rect 11706 16395 11749 16451
rect 11729 16343 11749 16395
rect 11706 16287 11749 16343
rect 11729 16235 11749 16287
rect 11706 16179 11749 16235
rect 11729 16127 11749 16179
rect 11706 16071 11749 16127
rect 11729 16019 11749 16071
rect 11706 15963 11749 16019
rect 11729 15911 11749 15963
rect 11706 15855 11749 15911
rect 11729 15803 11749 15855
rect 11706 15747 11749 15803
rect 11729 15695 11749 15747
rect 11706 15639 11749 15695
rect 11729 15587 11749 15639
rect 11706 15531 11749 15587
rect 11729 15479 11749 15531
rect 11706 15423 11749 15479
rect 11729 15371 11749 15423
rect 11706 15315 11749 15371
rect 11729 15263 11749 15315
rect 11706 15207 11749 15263
rect 11729 15155 11749 15207
rect 11706 15099 11749 15155
rect 11729 15047 11749 15099
rect 11706 14991 11749 15047
rect 11729 14939 11749 14991
rect 11706 14883 11749 14939
rect 11729 14831 11749 14883
rect 11706 14775 11749 14831
rect 11729 14723 11749 14775
rect 11706 14667 11749 14723
rect 11729 14615 11749 14667
rect 11706 14559 11749 14615
rect 11729 14507 11749 14559
rect 11706 14451 11749 14507
rect 11729 14399 11749 14451
rect 11706 14343 11749 14399
rect 11729 14291 11749 14343
rect 11706 14235 11749 14291
rect 11729 14183 11749 14235
rect 11706 14127 11749 14183
rect 11729 14075 11749 14127
rect 11706 14019 11749 14075
rect 11729 13967 11749 14019
rect 11706 13911 11749 13967
rect 11729 13859 11749 13911
rect 11706 13803 11749 13859
rect 11729 13751 11749 13803
rect 11706 13695 11749 13751
rect 11729 13643 11749 13695
rect 11706 13587 11749 13643
rect 11729 13535 11749 13587
rect 11706 13479 11749 13535
rect 11729 13427 11749 13479
rect 11706 13371 11749 13427
rect 11729 13319 11749 13371
rect 11706 13290 11749 13319
rect 11549 13263 11749 13290
rect 11549 13211 11569 13263
rect 11621 13211 11677 13263
rect 11729 13211 11749 13263
rect 1213 13048 1413 13211
rect 1481 13199 11481 13211
rect 1481 13196 3433 13199
rect 3485 13196 3541 13199
rect 3593 13196 3649 13199
rect 3701 13196 3757 13199
rect 3809 13196 3865 13199
rect 3917 13196 3973 13199
rect 4025 13196 4081 13199
rect 4133 13196 4189 13199
rect 4241 13196 4297 13199
rect 4349 13196 4405 13199
rect 4457 13196 4513 13199
rect 4565 13196 4621 13199
rect 4673 13196 4729 13199
rect 4781 13196 4837 13199
rect 4889 13196 4945 13199
rect 4997 13196 5053 13199
rect 5105 13196 5161 13199
rect 5213 13196 6566 13199
rect 6618 13196 6674 13199
rect 6726 13196 6782 13199
rect 6834 13196 6890 13199
rect 6942 13196 6998 13199
rect 7050 13196 7106 13199
rect 7158 13196 7214 13199
rect 7266 13196 7322 13199
rect 7374 13196 7430 13199
rect 7482 13196 7538 13199
rect 7590 13196 9677 13199
rect 9729 13196 9785 13199
rect 9837 13196 9893 13199
rect 9945 13196 10001 13199
rect 10053 13196 10109 13199
rect 10161 13196 10217 13199
rect 10269 13196 10325 13199
rect 10377 13196 10433 13199
rect 10485 13196 10541 13199
rect 10593 13196 10649 13199
rect 10701 13196 10757 13199
rect 10809 13196 10865 13199
rect 10917 13196 10973 13199
rect 11025 13196 11081 13199
rect 11133 13196 11189 13199
rect 11241 13196 11297 13199
rect 11349 13196 11405 13199
rect 11457 13196 11481 13199
rect 1481 13150 1494 13196
rect 11468 13150 11481 13196
rect 1481 13147 3433 13150
rect 3485 13147 3541 13150
rect 3593 13147 3649 13150
rect 3701 13147 3757 13150
rect 3809 13147 3865 13150
rect 3917 13147 3973 13150
rect 4025 13147 4081 13150
rect 4133 13147 4189 13150
rect 4241 13147 4297 13150
rect 4349 13147 4405 13150
rect 4457 13147 4513 13150
rect 4565 13147 4621 13150
rect 4673 13147 4729 13150
rect 4781 13147 4837 13150
rect 4889 13147 4945 13150
rect 4997 13147 5053 13150
rect 5105 13147 5161 13150
rect 5213 13147 6566 13150
rect 6618 13147 6674 13150
rect 6726 13147 6782 13150
rect 6834 13147 6890 13150
rect 6942 13147 6998 13150
rect 7050 13147 7106 13150
rect 7158 13147 7214 13150
rect 7266 13147 7322 13150
rect 7374 13147 7430 13150
rect 7482 13147 7538 13150
rect 7590 13147 9677 13150
rect 9729 13147 9785 13150
rect 9837 13147 9893 13150
rect 9945 13147 10001 13150
rect 10053 13147 10109 13150
rect 10161 13147 10217 13150
rect 10269 13147 10325 13150
rect 10377 13147 10433 13150
rect 10485 13147 10541 13150
rect 10593 13147 10649 13150
rect 10701 13147 10757 13150
rect 10809 13147 10865 13150
rect 10917 13147 10973 13150
rect 11025 13147 11081 13150
rect 11133 13147 11189 13150
rect 11241 13147 11297 13150
rect 11349 13147 11405 13150
rect 11457 13147 11481 13150
rect 1481 13135 11481 13147
rect 11549 13048 11749 13211
rect 1213 12848 11749 13048
rect 12001 12769 12012 18457
rect 950 12757 12012 12769
rect 950 12750 1505 12757
rect 1557 12750 1613 12757
rect 1665 12750 1721 12757
rect 1773 12750 1829 12757
rect 1881 12750 1937 12757
rect 1989 12750 2045 12757
rect 2097 12750 2153 12757
rect 2205 12750 2261 12757
rect 2313 12750 2369 12757
rect 2421 12750 2477 12757
rect 2529 12750 2585 12757
rect 2637 12750 2693 12757
rect 2745 12750 2801 12757
rect 2853 12750 2909 12757
rect 2961 12750 3017 12757
rect 3069 12750 3125 12757
rect 3177 12750 3233 12757
rect 3285 12750 5372 12757
rect 5424 12750 5480 12757
rect 5532 12750 5588 12757
rect 5640 12750 5696 12757
rect 5748 12750 5804 12757
rect 5856 12750 5912 12757
rect 5964 12750 6020 12757
rect 6072 12750 6128 12757
rect 6180 12750 6236 12757
rect 6288 12750 6344 12757
rect 6396 12750 7749 12757
rect 7801 12750 7857 12757
rect 7909 12750 7965 12757
rect 8017 12750 8073 12757
rect 8125 12750 8181 12757
rect 8233 12750 8289 12757
rect 8341 12750 8397 12757
rect 8449 12750 8505 12757
rect 8557 12750 8613 12757
rect 8665 12750 8721 12757
rect 8773 12750 8829 12757
rect 8881 12750 8937 12757
rect 8989 12750 9045 12757
rect 9097 12750 9153 12757
rect 9205 12750 9261 12757
rect 9313 12750 9369 12757
rect 9421 12750 9477 12757
rect 9529 12750 12012 12757
rect 950 12604 1058 12750
rect 11904 12604 12012 12750
rect 950 12597 1505 12604
rect 1557 12597 1613 12604
rect 1665 12597 1721 12604
rect 1773 12597 1829 12604
rect 1881 12597 1937 12604
rect 1989 12597 2045 12604
rect 2097 12597 2153 12604
rect 2205 12597 2261 12604
rect 2313 12597 2369 12604
rect 2421 12597 2477 12604
rect 2529 12597 2585 12604
rect 2637 12597 2693 12604
rect 2745 12597 2801 12604
rect 2853 12597 2909 12604
rect 2961 12597 3017 12604
rect 3069 12597 3125 12604
rect 3177 12597 3233 12604
rect 3285 12597 5372 12604
rect 5424 12597 5480 12604
rect 5532 12597 5588 12604
rect 5640 12597 5696 12604
rect 5748 12597 5804 12604
rect 5856 12597 5912 12604
rect 5964 12597 6020 12604
rect 6072 12597 6128 12604
rect 6180 12597 6236 12604
rect 6288 12597 6344 12604
rect 6396 12597 7749 12604
rect 7801 12597 7857 12604
rect 7909 12597 7965 12604
rect 8017 12597 8073 12604
rect 8125 12597 8181 12604
rect 8233 12597 8289 12604
rect 8341 12597 8397 12604
rect 8449 12597 8505 12604
rect 8557 12597 8613 12604
rect 8665 12597 8721 12604
rect 8773 12597 8829 12604
rect 8881 12597 8937 12604
rect 8989 12597 9045 12604
rect 9097 12597 9153 12604
rect 9205 12597 9261 12604
rect 9313 12597 9369 12604
rect 9421 12597 9477 12604
rect 9529 12597 12012 12604
rect 950 12585 12012 12597
rect 950 6897 961 12585
rect 1213 12306 11749 12506
rect 1213 12143 1413 12306
rect 1481 12207 11481 12219
rect 1481 12204 3433 12207
rect 3485 12204 3541 12207
rect 3593 12204 3649 12207
rect 3701 12204 3757 12207
rect 3809 12204 3865 12207
rect 3917 12204 3973 12207
rect 4025 12204 4081 12207
rect 4133 12204 4189 12207
rect 4241 12204 4297 12207
rect 4349 12204 4405 12207
rect 4457 12204 4513 12207
rect 4565 12204 4621 12207
rect 4673 12204 4729 12207
rect 4781 12204 4837 12207
rect 4889 12204 4945 12207
rect 4997 12204 5053 12207
rect 5105 12204 5161 12207
rect 5213 12204 6566 12207
rect 6618 12204 6674 12207
rect 6726 12204 6782 12207
rect 6834 12204 6890 12207
rect 6942 12204 6998 12207
rect 7050 12204 7106 12207
rect 7158 12204 7214 12207
rect 7266 12204 7322 12207
rect 7374 12204 7430 12207
rect 7482 12204 7538 12207
rect 7590 12204 9677 12207
rect 9729 12204 9785 12207
rect 9837 12204 9893 12207
rect 9945 12204 10001 12207
rect 10053 12204 10109 12207
rect 10161 12204 10217 12207
rect 10269 12204 10325 12207
rect 10377 12204 10433 12207
rect 10485 12204 10541 12207
rect 10593 12204 10649 12207
rect 10701 12204 10757 12207
rect 10809 12204 10865 12207
rect 10917 12204 10973 12207
rect 11025 12204 11081 12207
rect 11133 12204 11189 12207
rect 11241 12204 11297 12207
rect 11349 12204 11405 12207
rect 11457 12204 11481 12207
rect 1481 12158 1494 12204
rect 11468 12158 11481 12204
rect 1481 12155 3433 12158
rect 3485 12155 3541 12158
rect 3593 12155 3649 12158
rect 3701 12155 3757 12158
rect 3809 12155 3865 12158
rect 3917 12155 3973 12158
rect 4025 12155 4081 12158
rect 4133 12155 4189 12158
rect 4241 12155 4297 12158
rect 4349 12155 4405 12158
rect 4457 12155 4513 12158
rect 4565 12155 4621 12158
rect 4673 12155 4729 12158
rect 4781 12155 4837 12158
rect 4889 12155 4945 12158
rect 4997 12155 5053 12158
rect 5105 12155 5161 12158
rect 5213 12155 6566 12158
rect 6618 12155 6674 12158
rect 6726 12155 6782 12158
rect 6834 12155 6890 12158
rect 6942 12155 6998 12158
rect 7050 12155 7106 12158
rect 7158 12155 7214 12158
rect 7266 12155 7322 12158
rect 7374 12155 7430 12158
rect 7482 12155 7538 12158
rect 7590 12155 9677 12158
rect 9729 12155 9785 12158
rect 9837 12155 9893 12158
rect 9945 12155 10001 12158
rect 10053 12155 10109 12158
rect 10161 12155 10217 12158
rect 10269 12155 10325 12158
rect 10377 12155 10433 12158
rect 10485 12155 10541 12158
rect 10593 12155 10649 12158
rect 10701 12155 10757 12158
rect 10809 12155 10865 12158
rect 10917 12155 10973 12158
rect 11025 12155 11081 12158
rect 11133 12155 11189 12158
rect 11241 12155 11297 12158
rect 11349 12155 11405 12158
rect 11457 12155 11481 12158
rect 1481 12143 11481 12155
rect 11549 12143 11749 12306
rect 1213 12091 1233 12143
rect 1285 12091 1341 12143
rect 1393 12091 1413 12143
rect 1213 12064 1413 12091
rect 1213 12035 1256 12064
rect 1213 11983 1233 12035
rect 1213 11927 1256 11983
rect 1213 11875 1233 11927
rect 1213 11819 1256 11875
rect 1213 11767 1233 11819
rect 1213 11711 1256 11767
rect 1213 11659 1233 11711
rect 1213 11603 1256 11659
rect 1213 11551 1233 11603
rect 1213 11495 1256 11551
rect 1213 11443 1233 11495
rect 1213 11387 1256 11443
rect 1213 11335 1233 11387
rect 1213 11279 1256 11335
rect 1213 11227 1233 11279
rect 1213 11171 1256 11227
rect 1213 11119 1233 11171
rect 1213 11063 1256 11119
rect 1213 11011 1233 11063
rect 1213 10955 1256 11011
rect 1213 10903 1233 10955
rect 1213 10847 1256 10903
rect 1213 10795 1233 10847
rect 1213 10739 1256 10795
rect 1213 10687 1233 10739
rect 1213 10631 1256 10687
rect 1213 10579 1233 10631
rect 1213 10523 1256 10579
rect 1213 10471 1233 10523
rect 1213 10415 1256 10471
rect 1213 10363 1233 10415
rect 1213 10307 1256 10363
rect 1213 10255 1233 10307
rect 1213 10199 1256 10255
rect 1213 10147 1233 10199
rect 1213 10091 1256 10147
rect 1213 10039 1233 10091
rect 1213 9983 1256 10039
rect 1213 9931 1233 9983
rect 1213 9875 1256 9931
rect 1213 9823 1233 9875
rect 1213 9767 1256 9823
rect 1213 9715 1233 9767
rect 1213 9659 1256 9715
rect 1213 9607 1233 9659
rect 1213 9551 1256 9607
rect 1213 9499 1233 9551
rect 1213 9443 1256 9499
rect 1213 9391 1233 9443
rect 1213 9335 1256 9391
rect 1213 9283 1233 9335
rect 1213 9227 1256 9283
rect 1213 9175 1233 9227
rect 1213 9119 1256 9175
rect 1213 9067 1233 9119
rect 1213 9011 1256 9067
rect 1213 8959 1233 9011
rect 1213 8903 1256 8959
rect 1213 8851 1233 8903
rect 1213 8795 1256 8851
rect 1213 8743 1233 8795
rect 1213 8687 1256 8743
rect 1213 8635 1233 8687
rect 1213 8579 1256 8635
rect 1213 8527 1233 8579
rect 1213 8471 1256 8527
rect 1213 8419 1233 8471
rect 1213 8363 1256 8419
rect 1213 8311 1233 8363
rect 1213 8255 1256 8311
rect 1213 8203 1233 8255
rect 1213 8147 1256 8203
rect 1213 8095 1233 8147
rect 1213 8039 1256 8095
rect 1213 7987 1233 8039
rect 1213 7931 1256 7987
rect 1213 7879 1233 7931
rect 1213 7823 1256 7879
rect 1213 7771 1233 7823
rect 1213 7715 1256 7771
rect 1213 7663 1233 7715
rect 1213 7607 1256 7663
rect 1213 7555 1233 7607
rect 1213 7499 1256 7555
rect 1213 7447 1233 7499
rect 1213 7418 1256 7447
rect 1402 7418 1413 12064
rect 11549 12091 11569 12143
rect 11621 12091 11677 12143
rect 11729 12091 11749 12143
rect 11549 12064 11749 12091
rect 1481 11963 11481 11975
rect 1481 11960 1505 11963
rect 1557 11960 1613 11963
rect 1665 11960 1721 11963
rect 1773 11960 1829 11963
rect 1881 11960 1937 11963
rect 1989 11960 2045 11963
rect 2097 11960 2153 11963
rect 2205 11960 2261 11963
rect 2313 11960 2369 11963
rect 2421 11960 2477 11963
rect 2529 11960 2585 11963
rect 2637 11960 2693 11963
rect 2745 11960 2801 11963
rect 2853 11960 2909 11963
rect 2961 11960 3017 11963
rect 3069 11960 3125 11963
rect 3177 11960 3233 11963
rect 3285 11960 5372 11963
rect 5424 11960 5480 11963
rect 5532 11960 5588 11963
rect 5640 11960 5696 11963
rect 5748 11960 5804 11963
rect 5856 11960 5912 11963
rect 5964 11960 6020 11963
rect 6072 11960 6128 11963
rect 6180 11960 6236 11963
rect 6288 11960 6344 11963
rect 6396 11960 7749 11963
rect 7801 11960 7857 11963
rect 7909 11960 7965 11963
rect 8017 11960 8073 11963
rect 8125 11960 8181 11963
rect 8233 11960 8289 11963
rect 8341 11960 8397 11963
rect 8449 11960 8505 11963
rect 8557 11960 8613 11963
rect 8665 11960 8721 11963
rect 8773 11960 8829 11963
rect 8881 11960 8937 11963
rect 8989 11960 9045 11963
rect 9097 11960 9153 11963
rect 9205 11960 9261 11963
rect 9313 11960 9369 11963
rect 9421 11960 9477 11963
rect 9529 11960 11481 11963
rect 1481 11914 1494 11960
rect 11468 11914 11481 11960
rect 1481 11911 1505 11914
rect 1557 11911 1613 11914
rect 1665 11911 1721 11914
rect 1773 11911 1829 11914
rect 1881 11911 1937 11914
rect 1989 11911 2045 11914
rect 2097 11911 2153 11914
rect 2205 11911 2261 11914
rect 2313 11911 2369 11914
rect 2421 11911 2477 11914
rect 2529 11911 2585 11914
rect 2637 11911 2693 11914
rect 2745 11911 2801 11914
rect 2853 11911 2909 11914
rect 2961 11911 3017 11914
rect 3069 11911 3125 11914
rect 3177 11911 3233 11914
rect 3285 11911 5372 11914
rect 5424 11911 5480 11914
rect 5532 11911 5588 11914
rect 5640 11911 5696 11914
rect 5748 11911 5804 11914
rect 5856 11911 5912 11914
rect 5964 11911 6020 11914
rect 6072 11911 6128 11914
rect 6180 11911 6236 11914
rect 6288 11911 6344 11914
rect 6396 11911 7749 11914
rect 7801 11911 7857 11914
rect 7909 11911 7965 11914
rect 8017 11911 8073 11914
rect 8125 11911 8181 11914
rect 8233 11911 8289 11914
rect 8341 11911 8397 11914
rect 8449 11911 8505 11914
rect 8557 11911 8613 11914
rect 8665 11911 8721 11914
rect 8773 11911 8829 11914
rect 8881 11911 8937 11914
rect 8989 11911 9045 11914
rect 9097 11911 9153 11914
rect 9205 11911 9261 11914
rect 9313 11911 9369 11914
rect 9421 11911 9477 11914
rect 9529 11911 11481 11914
rect 1481 11899 11481 11911
rect 1481 11719 11481 11731
rect 1481 11716 3433 11719
rect 3485 11716 3541 11719
rect 3593 11716 3649 11719
rect 3701 11716 3757 11719
rect 3809 11716 3865 11719
rect 3917 11716 3973 11719
rect 4025 11716 4081 11719
rect 4133 11716 4189 11719
rect 4241 11716 4297 11719
rect 4349 11716 4405 11719
rect 4457 11716 4513 11719
rect 4565 11716 4621 11719
rect 4673 11716 4729 11719
rect 4781 11716 4837 11719
rect 4889 11716 4945 11719
rect 4997 11716 5053 11719
rect 5105 11716 5161 11719
rect 5213 11716 6566 11719
rect 6618 11716 6674 11719
rect 6726 11716 6782 11719
rect 6834 11716 6890 11719
rect 6942 11716 6998 11719
rect 7050 11716 7106 11719
rect 7158 11716 7214 11719
rect 7266 11716 7322 11719
rect 7374 11716 7430 11719
rect 7482 11716 7538 11719
rect 7590 11716 9677 11719
rect 9729 11716 9785 11719
rect 9837 11716 9893 11719
rect 9945 11716 10001 11719
rect 10053 11716 10109 11719
rect 10161 11716 10217 11719
rect 10269 11716 10325 11719
rect 10377 11716 10433 11719
rect 10485 11716 10541 11719
rect 10593 11716 10649 11719
rect 10701 11716 10757 11719
rect 10809 11716 10865 11719
rect 10917 11716 10973 11719
rect 11025 11716 11081 11719
rect 11133 11716 11189 11719
rect 11241 11716 11297 11719
rect 11349 11716 11405 11719
rect 11457 11716 11481 11719
rect 1481 11670 1494 11716
rect 11468 11670 11481 11716
rect 1481 11667 3433 11670
rect 3485 11667 3541 11670
rect 3593 11667 3649 11670
rect 3701 11667 3757 11670
rect 3809 11667 3865 11670
rect 3917 11667 3973 11670
rect 4025 11667 4081 11670
rect 4133 11667 4189 11670
rect 4241 11667 4297 11670
rect 4349 11667 4405 11670
rect 4457 11667 4513 11670
rect 4565 11667 4621 11670
rect 4673 11667 4729 11670
rect 4781 11667 4837 11670
rect 4889 11667 4945 11670
rect 4997 11667 5053 11670
rect 5105 11667 5161 11670
rect 5213 11667 6566 11670
rect 6618 11667 6674 11670
rect 6726 11667 6782 11670
rect 6834 11667 6890 11670
rect 6942 11667 6998 11670
rect 7050 11667 7106 11670
rect 7158 11667 7214 11670
rect 7266 11667 7322 11670
rect 7374 11667 7430 11670
rect 7482 11667 7538 11670
rect 7590 11667 9677 11670
rect 9729 11667 9785 11670
rect 9837 11667 9893 11670
rect 9945 11667 10001 11670
rect 10053 11667 10109 11670
rect 10161 11667 10217 11670
rect 10269 11667 10325 11670
rect 10377 11667 10433 11670
rect 10485 11667 10541 11670
rect 10593 11667 10649 11670
rect 10701 11667 10757 11670
rect 10809 11667 10865 11670
rect 10917 11667 10973 11670
rect 11025 11667 11081 11670
rect 11133 11667 11189 11670
rect 11241 11667 11297 11670
rect 11349 11667 11405 11670
rect 11457 11667 11481 11670
rect 1481 11655 11481 11667
rect 1481 11475 11481 11487
rect 1481 11472 1505 11475
rect 1557 11472 1613 11475
rect 1665 11472 1721 11475
rect 1773 11472 1829 11475
rect 1881 11472 1937 11475
rect 1989 11472 2045 11475
rect 2097 11472 2153 11475
rect 2205 11472 2261 11475
rect 2313 11472 2369 11475
rect 2421 11472 2477 11475
rect 2529 11472 2585 11475
rect 2637 11472 2693 11475
rect 2745 11472 2801 11475
rect 2853 11472 2909 11475
rect 2961 11472 3017 11475
rect 3069 11472 3125 11475
rect 3177 11472 3233 11475
rect 3285 11472 5372 11475
rect 5424 11472 5480 11475
rect 5532 11472 5588 11475
rect 5640 11472 5696 11475
rect 5748 11472 5804 11475
rect 5856 11472 5912 11475
rect 5964 11472 6020 11475
rect 6072 11472 6128 11475
rect 6180 11472 6236 11475
rect 6288 11472 6344 11475
rect 6396 11472 7749 11475
rect 7801 11472 7857 11475
rect 7909 11472 7965 11475
rect 8017 11472 8073 11475
rect 8125 11472 8181 11475
rect 8233 11472 8289 11475
rect 8341 11472 8397 11475
rect 8449 11472 8505 11475
rect 8557 11472 8613 11475
rect 8665 11472 8721 11475
rect 8773 11472 8829 11475
rect 8881 11472 8937 11475
rect 8989 11472 9045 11475
rect 9097 11472 9153 11475
rect 9205 11472 9261 11475
rect 9313 11472 9369 11475
rect 9421 11472 9477 11475
rect 9529 11472 11481 11475
rect 1481 11426 1494 11472
rect 11468 11426 11481 11472
rect 1481 11423 1505 11426
rect 1557 11423 1613 11426
rect 1665 11423 1721 11426
rect 1773 11423 1829 11426
rect 1881 11423 1937 11426
rect 1989 11423 2045 11426
rect 2097 11423 2153 11426
rect 2205 11423 2261 11426
rect 2313 11423 2369 11426
rect 2421 11423 2477 11426
rect 2529 11423 2585 11426
rect 2637 11423 2693 11426
rect 2745 11423 2801 11426
rect 2853 11423 2909 11426
rect 2961 11423 3017 11426
rect 3069 11423 3125 11426
rect 3177 11423 3233 11426
rect 3285 11423 5372 11426
rect 5424 11423 5480 11426
rect 5532 11423 5588 11426
rect 5640 11423 5696 11426
rect 5748 11423 5804 11426
rect 5856 11423 5912 11426
rect 5964 11423 6020 11426
rect 6072 11423 6128 11426
rect 6180 11423 6236 11426
rect 6288 11423 6344 11426
rect 6396 11423 7749 11426
rect 7801 11423 7857 11426
rect 7909 11423 7965 11426
rect 8017 11423 8073 11426
rect 8125 11423 8181 11426
rect 8233 11423 8289 11426
rect 8341 11423 8397 11426
rect 8449 11423 8505 11426
rect 8557 11423 8613 11426
rect 8665 11423 8721 11426
rect 8773 11423 8829 11426
rect 8881 11423 8937 11426
rect 8989 11423 9045 11426
rect 9097 11423 9153 11426
rect 9205 11423 9261 11426
rect 9313 11423 9369 11426
rect 9421 11423 9477 11426
rect 9529 11423 11481 11426
rect 1481 11411 11481 11423
rect 1481 11231 11481 11243
rect 1481 11228 3433 11231
rect 3485 11228 3541 11231
rect 3593 11228 3649 11231
rect 3701 11228 3757 11231
rect 3809 11228 3865 11231
rect 3917 11228 3973 11231
rect 4025 11228 4081 11231
rect 4133 11228 4189 11231
rect 4241 11228 4297 11231
rect 4349 11228 4405 11231
rect 4457 11228 4513 11231
rect 4565 11228 4621 11231
rect 4673 11228 4729 11231
rect 4781 11228 4837 11231
rect 4889 11228 4945 11231
rect 4997 11228 5053 11231
rect 5105 11228 5161 11231
rect 5213 11228 6566 11231
rect 6618 11228 6674 11231
rect 6726 11228 6782 11231
rect 6834 11228 6890 11231
rect 6942 11228 6998 11231
rect 7050 11228 7106 11231
rect 7158 11228 7214 11231
rect 7266 11228 7322 11231
rect 7374 11228 7430 11231
rect 7482 11228 7538 11231
rect 7590 11228 9677 11231
rect 9729 11228 9785 11231
rect 9837 11228 9893 11231
rect 9945 11228 10001 11231
rect 10053 11228 10109 11231
rect 10161 11228 10217 11231
rect 10269 11228 10325 11231
rect 10377 11228 10433 11231
rect 10485 11228 10541 11231
rect 10593 11228 10649 11231
rect 10701 11228 10757 11231
rect 10809 11228 10865 11231
rect 10917 11228 10973 11231
rect 11025 11228 11081 11231
rect 11133 11228 11189 11231
rect 11241 11228 11297 11231
rect 11349 11228 11405 11231
rect 11457 11228 11481 11231
rect 1481 11182 1494 11228
rect 11468 11182 11481 11228
rect 1481 11179 3433 11182
rect 3485 11179 3541 11182
rect 3593 11179 3649 11182
rect 3701 11179 3757 11182
rect 3809 11179 3865 11182
rect 3917 11179 3973 11182
rect 4025 11179 4081 11182
rect 4133 11179 4189 11182
rect 4241 11179 4297 11182
rect 4349 11179 4405 11182
rect 4457 11179 4513 11182
rect 4565 11179 4621 11182
rect 4673 11179 4729 11182
rect 4781 11179 4837 11182
rect 4889 11179 4945 11182
rect 4997 11179 5053 11182
rect 5105 11179 5161 11182
rect 5213 11179 6566 11182
rect 6618 11179 6674 11182
rect 6726 11179 6782 11182
rect 6834 11179 6890 11182
rect 6942 11179 6998 11182
rect 7050 11179 7106 11182
rect 7158 11179 7214 11182
rect 7266 11179 7322 11182
rect 7374 11179 7430 11182
rect 7482 11179 7538 11182
rect 7590 11179 9677 11182
rect 9729 11179 9785 11182
rect 9837 11179 9893 11182
rect 9945 11179 10001 11182
rect 10053 11179 10109 11182
rect 10161 11179 10217 11182
rect 10269 11179 10325 11182
rect 10377 11179 10433 11182
rect 10485 11179 10541 11182
rect 10593 11179 10649 11182
rect 10701 11179 10757 11182
rect 10809 11179 10865 11182
rect 10917 11179 10973 11182
rect 11025 11179 11081 11182
rect 11133 11179 11189 11182
rect 11241 11179 11297 11182
rect 11349 11179 11405 11182
rect 11457 11179 11481 11182
rect 1481 11167 11481 11179
rect 1481 10987 11481 10999
rect 1481 10984 1505 10987
rect 1557 10984 1613 10987
rect 1665 10984 1721 10987
rect 1773 10984 1829 10987
rect 1881 10984 1937 10987
rect 1989 10984 2045 10987
rect 2097 10984 2153 10987
rect 2205 10984 2261 10987
rect 2313 10984 2369 10987
rect 2421 10984 2477 10987
rect 2529 10984 2585 10987
rect 2637 10984 2693 10987
rect 2745 10984 2801 10987
rect 2853 10984 2909 10987
rect 2961 10984 3017 10987
rect 3069 10984 3125 10987
rect 3177 10984 3233 10987
rect 3285 10984 5372 10987
rect 5424 10984 5480 10987
rect 5532 10984 5588 10987
rect 5640 10984 5696 10987
rect 5748 10984 5804 10987
rect 5856 10984 5912 10987
rect 5964 10984 6020 10987
rect 6072 10984 6128 10987
rect 6180 10984 6236 10987
rect 6288 10984 6344 10987
rect 6396 10984 7749 10987
rect 7801 10984 7857 10987
rect 7909 10984 7965 10987
rect 8017 10984 8073 10987
rect 8125 10984 8181 10987
rect 8233 10984 8289 10987
rect 8341 10984 8397 10987
rect 8449 10984 8505 10987
rect 8557 10984 8613 10987
rect 8665 10984 8721 10987
rect 8773 10984 8829 10987
rect 8881 10984 8937 10987
rect 8989 10984 9045 10987
rect 9097 10984 9153 10987
rect 9205 10984 9261 10987
rect 9313 10984 9369 10987
rect 9421 10984 9477 10987
rect 9529 10984 11481 10987
rect 1481 10938 1494 10984
rect 11468 10938 11481 10984
rect 1481 10935 1505 10938
rect 1557 10935 1613 10938
rect 1665 10935 1721 10938
rect 1773 10935 1829 10938
rect 1881 10935 1937 10938
rect 1989 10935 2045 10938
rect 2097 10935 2153 10938
rect 2205 10935 2261 10938
rect 2313 10935 2369 10938
rect 2421 10935 2477 10938
rect 2529 10935 2585 10938
rect 2637 10935 2693 10938
rect 2745 10935 2801 10938
rect 2853 10935 2909 10938
rect 2961 10935 3017 10938
rect 3069 10935 3125 10938
rect 3177 10935 3233 10938
rect 3285 10935 5372 10938
rect 5424 10935 5480 10938
rect 5532 10935 5588 10938
rect 5640 10935 5696 10938
rect 5748 10935 5804 10938
rect 5856 10935 5912 10938
rect 5964 10935 6020 10938
rect 6072 10935 6128 10938
rect 6180 10935 6236 10938
rect 6288 10935 6344 10938
rect 6396 10935 7749 10938
rect 7801 10935 7857 10938
rect 7909 10935 7965 10938
rect 8017 10935 8073 10938
rect 8125 10935 8181 10938
rect 8233 10935 8289 10938
rect 8341 10935 8397 10938
rect 8449 10935 8505 10938
rect 8557 10935 8613 10938
rect 8665 10935 8721 10938
rect 8773 10935 8829 10938
rect 8881 10935 8937 10938
rect 8989 10935 9045 10938
rect 9097 10935 9153 10938
rect 9205 10935 9261 10938
rect 9313 10935 9369 10938
rect 9421 10935 9477 10938
rect 9529 10935 11481 10938
rect 1481 10923 11481 10935
rect 1481 10743 11481 10755
rect 1481 10740 3433 10743
rect 3485 10740 3541 10743
rect 3593 10740 3649 10743
rect 3701 10740 3757 10743
rect 3809 10740 3865 10743
rect 3917 10740 3973 10743
rect 4025 10740 4081 10743
rect 4133 10740 4189 10743
rect 4241 10740 4297 10743
rect 4349 10740 4405 10743
rect 4457 10740 4513 10743
rect 4565 10740 4621 10743
rect 4673 10740 4729 10743
rect 4781 10740 4837 10743
rect 4889 10740 4945 10743
rect 4997 10740 5053 10743
rect 5105 10740 5161 10743
rect 5213 10740 6566 10743
rect 6618 10740 6674 10743
rect 6726 10740 6782 10743
rect 6834 10740 6890 10743
rect 6942 10740 6998 10743
rect 7050 10740 7106 10743
rect 7158 10740 7214 10743
rect 7266 10740 7322 10743
rect 7374 10740 7430 10743
rect 7482 10740 7538 10743
rect 7590 10740 9677 10743
rect 9729 10740 9785 10743
rect 9837 10740 9893 10743
rect 9945 10740 10001 10743
rect 10053 10740 10109 10743
rect 10161 10740 10217 10743
rect 10269 10740 10325 10743
rect 10377 10740 10433 10743
rect 10485 10740 10541 10743
rect 10593 10740 10649 10743
rect 10701 10740 10757 10743
rect 10809 10740 10865 10743
rect 10917 10740 10973 10743
rect 11025 10740 11081 10743
rect 11133 10740 11189 10743
rect 11241 10740 11297 10743
rect 11349 10740 11405 10743
rect 11457 10740 11481 10743
rect 1481 10694 1494 10740
rect 11468 10694 11481 10740
rect 1481 10691 3433 10694
rect 3485 10691 3541 10694
rect 3593 10691 3649 10694
rect 3701 10691 3757 10694
rect 3809 10691 3865 10694
rect 3917 10691 3973 10694
rect 4025 10691 4081 10694
rect 4133 10691 4189 10694
rect 4241 10691 4297 10694
rect 4349 10691 4405 10694
rect 4457 10691 4513 10694
rect 4565 10691 4621 10694
rect 4673 10691 4729 10694
rect 4781 10691 4837 10694
rect 4889 10691 4945 10694
rect 4997 10691 5053 10694
rect 5105 10691 5161 10694
rect 5213 10691 6566 10694
rect 6618 10691 6674 10694
rect 6726 10691 6782 10694
rect 6834 10691 6890 10694
rect 6942 10691 6998 10694
rect 7050 10691 7106 10694
rect 7158 10691 7214 10694
rect 7266 10691 7322 10694
rect 7374 10691 7430 10694
rect 7482 10691 7538 10694
rect 7590 10691 9677 10694
rect 9729 10691 9785 10694
rect 9837 10691 9893 10694
rect 9945 10691 10001 10694
rect 10053 10691 10109 10694
rect 10161 10691 10217 10694
rect 10269 10691 10325 10694
rect 10377 10691 10433 10694
rect 10485 10691 10541 10694
rect 10593 10691 10649 10694
rect 10701 10691 10757 10694
rect 10809 10691 10865 10694
rect 10917 10691 10973 10694
rect 11025 10691 11081 10694
rect 11133 10691 11189 10694
rect 11241 10691 11297 10694
rect 11349 10691 11405 10694
rect 11457 10691 11481 10694
rect 1481 10679 11481 10691
rect 1481 10499 11481 10511
rect 1481 10496 1505 10499
rect 1557 10496 1613 10499
rect 1665 10496 1721 10499
rect 1773 10496 1829 10499
rect 1881 10496 1937 10499
rect 1989 10496 2045 10499
rect 2097 10496 2153 10499
rect 2205 10496 2261 10499
rect 2313 10496 2369 10499
rect 2421 10496 2477 10499
rect 2529 10496 2585 10499
rect 2637 10496 2693 10499
rect 2745 10496 2801 10499
rect 2853 10496 2909 10499
rect 2961 10496 3017 10499
rect 3069 10496 3125 10499
rect 3177 10496 3233 10499
rect 3285 10496 5372 10499
rect 5424 10496 5480 10499
rect 5532 10496 5588 10499
rect 5640 10496 5696 10499
rect 5748 10496 5804 10499
rect 5856 10496 5912 10499
rect 5964 10496 6020 10499
rect 6072 10496 6128 10499
rect 6180 10496 6236 10499
rect 6288 10496 6344 10499
rect 6396 10496 7749 10499
rect 7801 10496 7857 10499
rect 7909 10496 7965 10499
rect 8017 10496 8073 10499
rect 8125 10496 8181 10499
rect 8233 10496 8289 10499
rect 8341 10496 8397 10499
rect 8449 10496 8505 10499
rect 8557 10496 8613 10499
rect 8665 10496 8721 10499
rect 8773 10496 8829 10499
rect 8881 10496 8937 10499
rect 8989 10496 9045 10499
rect 9097 10496 9153 10499
rect 9205 10496 9261 10499
rect 9313 10496 9369 10499
rect 9421 10496 9477 10499
rect 9529 10496 11481 10499
rect 1481 10450 1494 10496
rect 11468 10450 11481 10496
rect 1481 10447 1505 10450
rect 1557 10447 1613 10450
rect 1665 10447 1721 10450
rect 1773 10447 1829 10450
rect 1881 10447 1937 10450
rect 1989 10447 2045 10450
rect 2097 10447 2153 10450
rect 2205 10447 2261 10450
rect 2313 10447 2369 10450
rect 2421 10447 2477 10450
rect 2529 10447 2585 10450
rect 2637 10447 2693 10450
rect 2745 10447 2801 10450
rect 2853 10447 2909 10450
rect 2961 10447 3017 10450
rect 3069 10447 3125 10450
rect 3177 10447 3233 10450
rect 3285 10447 5372 10450
rect 5424 10447 5480 10450
rect 5532 10447 5588 10450
rect 5640 10447 5696 10450
rect 5748 10447 5804 10450
rect 5856 10447 5912 10450
rect 5964 10447 6020 10450
rect 6072 10447 6128 10450
rect 6180 10447 6236 10450
rect 6288 10447 6344 10450
rect 6396 10447 7749 10450
rect 7801 10447 7857 10450
rect 7909 10447 7965 10450
rect 8017 10447 8073 10450
rect 8125 10447 8181 10450
rect 8233 10447 8289 10450
rect 8341 10447 8397 10450
rect 8449 10447 8505 10450
rect 8557 10447 8613 10450
rect 8665 10447 8721 10450
rect 8773 10447 8829 10450
rect 8881 10447 8937 10450
rect 8989 10447 9045 10450
rect 9097 10447 9153 10450
rect 9205 10447 9261 10450
rect 9313 10447 9369 10450
rect 9421 10447 9477 10450
rect 9529 10447 11481 10450
rect 1481 10435 11481 10447
rect 1481 10255 11481 10267
rect 1481 10252 3433 10255
rect 3485 10252 3541 10255
rect 3593 10252 3649 10255
rect 3701 10252 3757 10255
rect 3809 10252 3865 10255
rect 3917 10252 3973 10255
rect 4025 10252 4081 10255
rect 4133 10252 4189 10255
rect 4241 10252 4297 10255
rect 4349 10252 4405 10255
rect 4457 10252 4513 10255
rect 4565 10252 4621 10255
rect 4673 10252 4729 10255
rect 4781 10252 4837 10255
rect 4889 10252 4945 10255
rect 4997 10252 5053 10255
rect 5105 10252 5161 10255
rect 5213 10252 6566 10255
rect 6618 10252 6674 10255
rect 6726 10252 6782 10255
rect 6834 10252 6890 10255
rect 6942 10252 6998 10255
rect 7050 10252 7106 10255
rect 7158 10252 7214 10255
rect 7266 10252 7322 10255
rect 7374 10252 7430 10255
rect 7482 10252 7538 10255
rect 7590 10252 9677 10255
rect 9729 10252 9785 10255
rect 9837 10252 9893 10255
rect 9945 10252 10001 10255
rect 10053 10252 10109 10255
rect 10161 10252 10217 10255
rect 10269 10252 10325 10255
rect 10377 10252 10433 10255
rect 10485 10252 10541 10255
rect 10593 10252 10649 10255
rect 10701 10252 10757 10255
rect 10809 10252 10865 10255
rect 10917 10252 10973 10255
rect 11025 10252 11081 10255
rect 11133 10252 11189 10255
rect 11241 10252 11297 10255
rect 11349 10252 11405 10255
rect 11457 10252 11481 10255
rect 1481 10206 1494 10252
rect 11468 10206 11481 10252
rect 1481 10203 3433 10206
rect 3485 10203 3541 10206
rect 3593 10203 3649 10206
rect 3701 10203 3757 10206
rect 3809 10203 3865 10206
rect 3917 10203 3973 10206
rect 4025 10203 4081 10206
rect 4133 10203 4189 10206
rect 4241 10203 4297 10206
rect 4349 10203 4405 10206
rect 4457 10203 4513 10206
rect 4565 10203 4621 10206
rect 4673 10203 4729 10206
rect 4781 10203 4837 10206
rect 4889 10203 4945 10206
rect 4997 10203 5053 10206
rect 5105 10203 5161 10206
rect 5213 10203 6566 10206
rect 6618 10203 6674 10206
rect 6726 10203 6782 10206
rect 6834 10203 6890 10206
rect 6942 10203 6998 10206
rect 7050 10203 7106 10206
rect 7158 10203 7214 10206
rect 7266 10203 7322 10206
rect 7374 10203 7430 10206
rect 7482 10203 7538 10206
rect 7590 10203 9677 10206
rect 9729 10203 9785 10206
rect 9837 10203 9893 10206
rect 9945 10203 10001 10206
rect 10053 10203 10109 10206
rect 10161 10203 10217 10206
rect 10269 10203 10325 10206
rect 10377 10203 10433 10206
rect 10485 10203 10541 10206
rect 10593 10203 10649 10206
rect 10701 10203 10757 10206
rect 10809 10203 10865 10206
rect 10917 10203 10973 10206
rect 11025 10203 11081 10206
rect 11133 10203 11189 10206
rect 11241 10203 11297 10206
rect 11349 10203 11405 10206
rect 11457 10203 11481 10206
rect 1481 10191 11481 10203
rect 1481 10011 11481 10023
rect 1481 10008 1505 10011
rect 1557 10008 1613 10011
rect 1665 10008 1721 10011
rect 1773 10008 1829 10011
rect 1881 10008 1937 10011
rect 1989 10008 2045 10011
rect 2097 10008 2153 10011
rect 2205 10008 2261 10011
rect 2313 10008 2369 10011
rect 2421 10008 2477 10011
rect 2529 10008 2585 10011
rect 2637 10008 2693 10011
rect 2745 10008 2801 10011
rect 2853 10008 2909 10011
rect 2961 10008 3017 10011
rect 3069 10008 3125 10011
rect 3177 10008 3233 10011
rect 3285 10008 5372 10011
rect 5424 10008 5480 10011
rect 5532 10008 5588 10011
rect 5640 10008 5696 10011
rect 5748 10008 5804 10011
rect 5856 10008 5912 10011
rect 5964 10008 6020 10011
rect 6072 10008 6128 10011
rect 6180 10008 6236 10011
rect 6288 10008 6344 10011
rect 6396 10008 7749 10011
rect 7801 10008 7857 10011
rect 7909 10008 7965 10011
rect 8017 10008 8073 10011
rect 8125 10008 8181 10011
rect 8233 10008 8289 10011
rect 8341 10008 8397 10011
rect 8449 10008 8505 10011
rect 8557 10008 8613 10011
rect 8665 10008 8721 10011
rect 8773 10008 8829 10011
rect 8881 10008 8937 10011
rect 8989 10008 9045 10011
rect 9097 10008 9153 10011
rect 9205 10008 9261 10011
rect 9313 10008 9369 10011
rect 9421 10008 9477 10011
rect 9529 10008 11481 10011
rect 1481 9962 1494 10008
rect 11468 9962 11481 10008
rect 1481 9959 1505 9962
rect 1557 9959 1613 9962
rect 1665 9959 1721 9962
rect 1773 9959 1829 9962
rect 1881 9959 1937 9962
rect 1989 9959 2045 9962
rect 2097 9959 2153 9962
rect 2205 9959 2261 9962
rect 2313 9959 2369 9962
rect 2421 9959 2477 9962
rect 2529 9959 2585 9962
rect 2637 9959 2693 9962
rect 2745 9959 2801 9962
rect 2853 9959 2909 9962
rect 2961 9959 3017 9962
rect 3069 9959 3125 9962
rect 3177 9959 3233 9962
rect 3285 9959 5372 9962
rect 5424 9959 5480 9962
rect 5532 9959 5588 9962
rect 5640 9959 5696 9962
rect 5748 9959 5804 9962
rect 5856 9959 5912 9962
rect 5964 9959 6020 9962
rect 6072 9959 6128 9962
rect 6180 9959 6236 9962
rect 6288 9959 6344 9962
rect 6396 9959 7749 9962
rect 7801 9959 7857 9962
rect 7909 9959 7965 9962
rect 8017 9959 8073 9962
rect 8125 9959 8181 9962
rect 8233 9959 8289 9962
rect 8341 9959 8397 9962
rect 8449 9959 8505 9962
rect 8557 9959 8613 9962
rect 8665 9959 8721 9962
rect 8773 9959 8829 9962
rect 8881 9959 8937 9962
rect 8989 9959 9045 9962
rect 9097 9959 9153 9962
rect 9205 9959 9261 9962
rect 9313 9959 9369 9962
rect 9421 9959 9477 9962
rect 9529 9959 11481 9962
rect 1481 9947 11481 9959
rect 1481 9767 11481 9779
rect 1481 9764 3433 9767
rect 3485 9764 3541 9767
rect 3593 9764 3649 9767
rect 3701 9764 3757 9767
rect 3809 9764 3865 9767
rect 3917 9764 3973 9767
rect 4025 9764 4081 9767
rect 4133 9764 4189 9767
rect 4241 9764 4297 9767
rect 4349 9764 4405 9767
rect 4457 9764 4513 9767
rect 4565 9764 4621 9767
rect 4673 9764 4729 9767
rect 4781 9764 4837 9767
rect 4889 9764 4945 9767
rect 4997 9764 5053 9767
rect 5105 9764 5161 9767
rect 5213 9764 6566 9767
rect 6618 9764 6674 9767
rect 6726 9764 6782 9767
rect 6834 9764 6890 9767
rect 6942 9764 6998 9767
rect 7050 9764 7106 9767
rect 7158 9764 7214 9767
rect 7266 9764 7322 9767
rect 7374 9764 7430 9767
rect 7482 9764 7538 9767
rect 7590 9764 9677 9767
rect 9729 9764 9785 9767
rect 9837 9764 9893 9767
rect 9945 9764 10001 9767
rect 10053 9764 10109 9767
rect 10161 9764 10217 9767
rect 10269 9764 10325 9767
rect 10377 9764 10433 9767
rect 10485 9764 10541 9767
rect 10593 9764 10649 9767
rect 10701 9764 10757 9767
rect 10809 9764 10865 9767
rect 10917 9764 10973 9767
rect 11025 9764 11081 9767
rect 11133 9764 11189 9767
rect 11241 9764 11297 9767
rect 11349 9764 11405 9767
rect 11457 9764 11481 9767
rect 1481 9718 1494 9764
rect 11468 9718 11481 9764
rect 1481 9715 3433 9718
rect 3485 9715 3541 9718
rect 3593 9715 3649 9718
rect 3701 9715 3757 9718
rect 3809 9715 3865 9718
rect 3917 9715 3973 9718
rect 4025 9715 4081 9718
rect 4133 9715 4189 9718
rect 4241 9715 4297 9718
rect 4349 9715 4405 9718
rect 4457 9715 4513 9718
rect 4565 9715 4621 9718
rect 4673 9715 4729 9718
rect 4781 9715 4837 9718
rect 4889 9715 4945 9718
rect 4997 9715 5053 9718
rect 5105 9715 5161 9718
rect 5213 9715 6566 9718
rect 6618 9715 6674 9718
rect 6726 9715 6782 9718
rect 6834 9715 6890 9718
rect 6942 9715 6998 9718
rect 7050 9715 7106 9718
rect 7158 9715 7214 9718
rect 7266 9715 7322 9718
rect 7374 9715 7430 9718
rect 7482 9715 7538 9718
rect 7590 9715 9677 9718
rect 9729 9715 9785 9718
rect 9837 9715 9893 9718
rect 9945 9715 10001 9718
rect 10053 9715 10109 9718
rect 10161 9715 10217 9718
rect 10269 9715 10325 9718
rect 10377 9715 10433 9718
rect 10485 9715 10541 9718
rect 10593 9715 10649 9718
rect 10701 9715 10757 9718
rect 10809 9715 10865 9718
rect 10917 9715 10973 9718
rect 11025 9715 11081 9718
rect 11133 9715 11189 9718
rect 11241 9715 11297 9718
rect 11349 9715 11405 9718
rect 11457 9715 11481 9718
rect 1481 9703 11481 9715
rect 1481 9523 11481 9535
rect 1481 9520 1505 9523
rect 1557 9520 1613 9523
rect 1665 9520 1721 9523
rect 1773 9520 1829 9523
rect 1881 9520 1937 9523
rect 1989 9520 2045 9523
rect 2097 9520 2153 9523
rect 2205 9520 2261 9523
rect 2313 9520 2369 9523
rect 2421 9520 2477 9523
rect 2529 9520 2585 9523
rect 2637 9520 2693 9523
rect 2745 9520 2801 9523
rect 2853 9520 2909 9523
rect 2961 9520 3017 9523
rect 3069 9520 3125 9523
rect 3177 9520 3233 9523
rect 3285 9520 5372 9523
rect 5424 9520 5480 9523
rect 5532 9520 5588 9523
rect 5640 9520 5696 9523
rect 5748 9520 5804 9523
rect 5856 9520 5912 9523
rect 5964 9520 6020 9523
rect 6072 9520 6128 9523
rect 6180 9520 6236 9523
rect 6288 9520 6344 9523
rect 6396 9520 7749 9523
rect 7801 9520 7857 9523
rect 7909 9520 7965 9523
rect 8017 9520 8073 9523
rect 8125 9520 8181 9523
rect 8233 9520 8289 9523
rect 8341 9520 8397 9523
rect 8449 9520 8505 9523
rect 8557 9520 8613 9523
rect 8665 9520 8721 9523
rect 8773 9520 8829 9523
rect 8881 9520 8937 9523
rect 8989 9520 9045 9523
rect 9097 9520 9153 9523
rect 9205 9520 9261 9523
rect 9313 9520 9369 9523
rect 9421 9520 9477 9523
rect 9529 9520 11481 9523
rect 1481 9474 1494 9520
rect 11468 9474 11481 9520
rect 1481 9471 1505 9474
rect 1557 9471 1613 9474
rect 1665 9471 1721 9474
rect 1773 9471 1829 9474
rect 1881 9471 1937 9474
rect 1989 9471 2045 9474
rect 2097 9471 2153 9474
rect 2205 9471 2261 9474
rect 2313 9471 2369 9474
rect 2421 9471 2477 9474
rect 2529 9471 2585 9474
rect 2637 9471 2693 9474
rect 2745 9471 2801 9474
rect 2853 9471 2909 9474
rect 2961 9471 3017 9474
rect 3069 9471 3125 9474
rect 3177 9471 3233 9474
rect 3285 9471 5372 9474
rect 5424 9471 5480 9474
rect 5532 9471 5588 9474
rect 5640 9471 5696 9474
rect 5748 9471 5804 9474
rect 5856 9471 5912 9474
rect 5964 9471 6020 9474
rect 6072 9471 6128 9474
rect 6180 9471 6236 9474
rect 6288 9471 6344 9474
rect 6396 9471 7749 9474
rect 7801 9471 7857 9474
rect 7909 9471 7965 9474
rect 8017 9471 8073 9474
rect 8125 9471 8181 9474
rect 8233 9471 8289 9474
rect 8341 9471 8397 9474
rect 8449 9471 8505 9474
rect 8557 9471 8613 9474
rect 8665 9471 8721 9474
rect 8773 9471 8829 9474
rect 8881 9471 8937 9474
rect 8989 9471 9045 9474
rect 9097 9471 9153 9474
rect 9205 9471 9261 9474
rect 9313 9471 9369 9474
rect 9421 9471 9477 9474
rect 9529 9471 11481 9474
rect 1481 9459 11481 9471
rect 1481 9279 11481 9291
rect 1481 9276 3433 9279
rect 3485 9276 3541 9279
rect 3593 9276 3649 9279
rect 3701 9276 3757 9279
rect 3809 9276 3865 9279
rect 3917 9276 3973 9279
rect 4025 9276 4081 9279
rect 4133 9276 4189 9279
rect 4241 9276 4297 9279
rect 4349 9276 4405 9279
rect 4457 9276 4513 9279
rect 4565 9276 4621 9279
rect 4673 9276 4729 9279
rect 4781 9276 4837 9279
rect 4889 9276 4945 9279
rect 4997 9276 5053 9279
rect 5105 9276 5161 9279
rect 5213 9276 6566 9279
rect 6618 9276 6674 9279
rect 6726 9276 6782 9279
rect 6834 9276 6890 9279
rect 6942 9276 6998 9279
rect 7050 9276 7106 9279
rect 7158 9276 7214 9279
rect 7266 9276 7322 9279
rect 7374 9276 7430 9279
rect 7482 9276 7538 9279
rect 7590 9276 9677 9279
rect 9729 9276 9785 9279
rect 9837 9276 9893 9279
rect 9945 9276 10001 9279
rect 10053 9276 10109 9279
rect 10161 9276 10217 9279
rect 10269 9276 10325 9279
rect 10377 9276 10433 9279
rect 10485 9276 10541 9279
rect 10593 9276 10649 9279
rect 10701 9276 10757 9279
rect 10809 9276 10865 9279
rect 10917 9276 10973 9279
rect 11025 9276 11081 9279
rect 11133 9276 11189 9279
rect 11241 9276 11297 9279
rect 11349 9276 11405 9279
rect 11457 9276 11481 9279
rect 1481 9230 1494 9276
rect 11468 9230 11481 9276
rect 1481 9227 3433 9230
rect 3485 9227 3541 9230
rect 3593 9227 3649 9230
rect 3701 9227 3757 9230
rect 3809 9227 3865 9230
rect 3917 9227 3973 9230
rect 4025 9227 4081 9230
rect 4133 9227 4189 9230
rect 4241 9227 4297 9230
rect 4349 9227 4405 9230
rect 4457 9227 4513 9230
rect 4565 9227 4621 9230
rect 4673 9227 4729 9230
rect 4781 9227 4837 9230
rect 4889 9227 4945 9230
rect 4997 9227 5053 9230
rect 5105 9227 5161 9230
rect 5213 9227 6566 9230
rect 6618 9227 6674 9230
rect 6726 9227 6782 9230
rect 6834 9227 6890 9230
rect 6942 9227 6998 9230
rect 7050 9227 7106 9230
rect 7158 9227 7214 9230
rect 7266 9227 7322 9230
rect 7374 9227 7430 9230
rect 7482 9227 7538 9230
rect 7590 9227 9677 9230
rect 9729 9227 9785 9230
rect 9837 9227 9893 9230
rect 9945 9227 10001 9230
rect 10053 9227 10109 9230
rect 10161 9227 10217 9230
rect 10269 9227 10325 9230
rect 10377 9227 10433 9230
rect 10485 9227 10541 9230
rect 10593 9227 10649 9230
rect 10701 9227 10757 9230
rect 10809 9227 10865 9230
rect 10917 9227 10973 9230
rect 11025 9227 11081 9230
rect 11133 9227 11189 9230
rect 11241 9227 11297 9230
rect 11349 9227 11405 9230
rect 11457 9227 11481 9230
rect 1481 9215 11481 9227
rect 1481 9035 11481 9047
rect 1481 9032 1505 9035
rect 1557 9032 1613 9035
rect 1665 9032 1721 9035
rect 1773 9032 1829 9035
rect 1881 9032 1937 9035
rect 1989 9032 2045 9035
rect 2097 9032 2153 9035
rect 2205 9032 2261 9035
rect 2313 9032 2369 9035
rect 2421 9032 2477 9035
rect 2529 9032 2585 9035
rect 2637 9032 2693 9035
rect 2745 9032 2801 9035
rect 2853 9032 2909 9035
rect 2961 9032 3017 9035
rect 3069 9032 3125 9035
rect 3177 9032 3233 9035
rect 3285 9032 5372 9035
rect 5424 9032 5480 9035
rect 5532 9032 5588 9035
rect 5640 9032 5696 9035
rect 5748 9032 5804 9035
rect 5856 9032 5912 9035
rect 5964 9032 6020 9035
rect 6072 9032 6128 9035
rect 6180 9032 6236 9035
rect 6288 9032 6344 9035
rect 6396 9032 7749 9035
rect 7801 9032 7857 9035
rect 7909 9032 7965 9035
rect 8017 9032 8073 9035
rect 8125 9032 8181 9035
rect 8233 9032 8289 9035
rect 8341 9032 8397 9035
rect 8449 9032 8505 9035
rect 8557 9032 8613 9035
rect 8665 9032 8721 9035
rect 8773 9032 8829 9035
rect 8881 9032 8937 9035
rect 8989 9032 9045 9035
rect 9097 9032 9153 9035
rect 9205 9032 9261 9035
rect 9313 9032 9369 9035
rect 9421 9032 9477 9035
rect 9529 9032 11481 9035
rect 1481 8986 1494 9032
rect 11468 8986 11481 9032
rect 1481 8983 1505 8986
rect 1557 8983 1613 8986
rect 1665 8983 1721 8986
rect 1773 8983 1829 8986
rect 1881 8983 1937 8986
rect 1989 8983 2045 8986
rect 2097 8983 2153 8986
rect 2205 8983 2261 8986
rect 2313 8983 2369 8986
rect 2421 8983 2477 8986
rect 2529 8983 2585 8986
rect 2637 8983 2693 8986
rect 2745 8983 2801 8986
rect 2853 8983 2909 8986
rect 2961 8983 3017 8986
rect 3069 8983 3125 8986
rect 3177 8983 3233 8986
rect 3285 8983 5372 8986
rect 5424 8983 5480 8986
rect 5532 8983 5588 8986
rect 5640 8983 5696 8986
rect 5748 8983 5804 8986
rect 5856 8983 5912 8986
rect 5964 8983 6020 8986
rect 6072 8983 6128 8986
rect 6180 8983 6236 8986
rect 6288 8983 6344 8986
rect 6396 8983 7749 8986
rect 7801 8983 7857 8986
rect 7909 8983 7965 8986
rect 8017 8983 8073 8986
rect 8125 8983 8181 8986
rect 8233 8983 8289 8986
rect 8341 8983 8397 8986
rect 8449 8983 8505 8986
rect 8557 8983 8613 8986
rect 8665 8983 8721 8986
rect 8773 8983 8829 8986
rect 8881 8983 8937 8986
rect 8989 8983 9045 8986
rect 9097 8983 9153 8986
rect 9205 8983 9261 8986
rect 9313 8983 9369 8986
rect 9421 8983 9477 8986
rect 9529 8983 11481 8986
rect 1481 8971 11481 8983
rect 1481 8791 11481 8803
rect 1481 8788 3433 8791
rect 3485 8788 3541 8791
rect 3593 8788 3649 8791
rect 3701 8788 3757 8791
rect 3809 8788 3865 8791
rect 3917 8788 3973 8791
rect 4025 8788 4081 8791
rect 4133 8788 4189 8791
rect 4241 8788 4297 8791
rect 4349 8788 4405 8791
rect 4457 8788 4513 8791
rect 4565 8788 4621 8791
rect 4673 8788 4729 8791
rect 4781 8788 4837 8791
rect 4889 8788 4945 8791
rect 4997 8788 5053 8791
rect 5105 8788 5161 8791
rect 5213 8788 6566 8791
rect 6618 8788 6674 8791
rect 6726 8788 6782 8791
rect 6834 8788 6890 8791
rect 6942 8788 6998 8791
rect 7050 8788 7106 8791
rect 7158 8788 7214 8791
rect 7266 8788 7322 8791
rect 7374 8788 7430 8791
rect 7482 8788 7538 8791
rect 7590 8788 9677 8791
rect 9729 8788 9785 8791
rect 9837 8788 9893 8791
rect 9945 8788 10001 8791
rect 10053 8788 10109 8791
rect 10161 8788 10217 8791
rect 10269 8788 10325 8791
rect 10377 8788 10433 8791
rect 10485 8788 10541 8791
rect 10593 8788 10649 8791
rect 10701 8788 10757 8791
rect 10809 8788 10865 8791
rect 10917 8788 10973 8791
rect 11025 8788 11081 8791
rect 11133 8788 11189 8791
rect 11241 8788 11297 8791
rect 11349 8788 11405 8791
rect 11457 8788 11481 8791
rect 1481 8742 1494 8788
rect 11468 8742 11481 8788
rect 1481 8739 3433 8742
rect 3485 8739 3541 8742
rect 3593 8739 3649 8742
rect 3701 8739 3757 8742
rect 3809 8739 3865 8742
rect 3917 8739 3973 8742
rect 4025 8739 4081 8742
rect 4133 8739 4189 8742
rect 4241 8739 4297 8742
rect 4349 8739 4405 8742
rect 4457 8739 4513 8742
rect 4565 8739 4621 8742
rect 4673 8739 4729 8742
rect 4781 8739 4837 8742
rect 4889 8739 4945 8742
rect 4997 8739 5053 8742
rect 5105 8739 5161 8742
rect 5213 8739 6566 8742
rect 6618 8739 6674 8742
rect 6726 8739 6782 8742
rect 6834 8739 6890 8742
rect 6942 8739 6998 8742
rect 7050 8739 7106 8742
rect 7158 8739 7214 8742
rect 7266 8739 7322 8742
rect 7374 8739 7430 8742
rect 7482 8739 7538 8742
rect 7590 8739 9677 8742
rect 9729 8739 9785 8742
rect 9837 8739 9893 8742
rect 9945 8739 10001 8742
rect 10053 8739 10109 8742
rect 10161 8739 10217 8742
rect 10269 8739 10325 8742
rect 10377 8739 10433 8742
rect 10485 8739 10541 8742
rect 10593 8739 10649 8742
rect 10701 8739 10757 8742
rect 10809 8739 10865 8742
rect 10917 8739 10973 8742
rect 11025 8739 11081 8742
rect 11133 8739 11189 8742
rect 11241 8739 11297 8742
rect 11349 8739 11405 8742
rect 11457 8739 11481 8742
rect 1481 8727 11481 8739
rect 1481 8547 11481 8559
rect 1481 8544 1505 8547
rect 1557 8544 1613 8547
rect 1665 8544 1721 8547
rect 1773 8544 1829 8547
rect 1881 8544 1937 8547
rect 1989 8544 2045 8547
rect 2097 8544 2153 8547
rect 2205 8544 2261 8547
rect 2313 8544 2369 8547
rect 2421 8544 2477 8547
rect 2529 8544 2585 8547
rect 2637 8544 2693 8547
rect 2745 8544 2801 8547
rect 2853 8544 2909 8547
rect 2961 8544 3017 8547
rect 3069 8544 3125 8547
rect 3177 8544 3233 8547
rect 3285 8544 5372 8547
rect 5424 8544 5480 8547
rect 5532 8544 5588 8547
rect 5640 8544 5696 8547
rect 5748 8544 5804 8547
rect 5856 8544 5912 8547
rect 5964 8544 6020 8547
rect 6072 8544 6128 8547
rect 6180 8544 6236 8547
rect 6288 8544 6344 8547
rect 6396 8544 7749 8547
rect 7801 8544 7857 8547
rect 7909 8544 7965 8547
rect 8017 8544 8073 8547
rect 8125 8544 8181 8547
rect 8233 8544 8289 8547
rect 8341 8544 8397 8547
rect 8449 8544 8505 8547
rect 8557 8544 8613 8547
rect 8665 8544 8721 8547
rect 8773 8544 8829 8547
rect 8881 8544 8937 8547
rect 8989 8544 9045 8547
rect 9097 8544 9153 8547
rect 9205 8544 9261 8547
rect 9313 8544 9369 8547
rect 9421 8544 9477 8547
rect 9529 8544 11481 8547
rect 1481 8498 1494 8544
rect 11468 8498 11481 8544
rect 1481 8495 1505 8498
rect 1557 8495 1613 8498
rect 1665 8495 1721 8498
rect 1773 8495 1829 8498
rect 1881 8495 1937 8498
rect 1989 8495 2045 8498
rect 2097 8495 2153 8498
rect 2205 8495 2261 8498
rect 2313 8495 2369 8498
rect 2421 8495 2477 8498
rect 2529 8495 2585 8498
rect 2637 8495 2693 8498
rect 2745 8495 2801 8498
rect 2853 8495 2909 8498
rect 2961 8495 3017 8498
rect 3069 8495 3125 8498
rect 3177 8495 3233 8498
rect 3285 8495 5372 8498
rect 5424 8495 5480 8498
rect 5532 8495 5588 8498
rect 5640 8495 5696 8498
rect 5748 8495 5804 8498
rect 5856 8495 5912 8498
rect 5964 8495 6020 8498
rect 6072 8495 6128 8498
rect 6180 8495 6236 8498
rect 6288 8495 6344 8498
rect 6396 8495 7749 8498
rect 7801 8495 7857 8498
rect 7909 8495 7965 8498
rect 8017 8495 8073 8498
rect 8125 8495 8181 8498
rect 8233 8495 8289 8498
rect 8341 8495 8397 8498
rect 8449 8495 8505 8498
rect 8557 8495 8613 8498
rect 8665 8495 8721 8498
rect 8773 8495 8829 8498
rect 8881 8495 8937 8498
rect 8989 8495 9045 8498
rect 9097 8495 9153 8498
rect 9205 8495 9261 8498
rect 9313 8495 9369 8498
rect 9421 8495 9477 8498
rect 9529 8495 11481 8498
rect 1481 8483 11481 8495
rect 1481 8303 11481 8315
rect 1481 8300 3433 8303
rect 3485 8300 3541 8303
rect 3593 8300 3649 8303
rect 3701 8300 3757 8303
rect 3809 8300 3865 8303
rect 3917 8300 3973 8303
rect 4025 8300 4081 8303
rect 4133 8300 4189 8303
rect 4241 8300 4297 8303
rect 4349 8300 4405 8303
rect 4457 8300 4513 8303
rect 4565 8300 4621 8303
rect 4673 8300 4729 8303
rect 4781 8300 4837 8303
rect 4889 8300 4945 8303
rect 4997 8300 5053 8303
rect 5105 8300 5161 8303
rect 5213 8300 6566 8303
rect 6618 8300 6674 8303
rect 6726 8300 6782 8303
rect 6834 8300 6890 8303
rect 6942 8300 6998 8303
rect 7050 8300 7106 8303
rect 7158 8300 7214 8303
rect 7266 8300 7322 8303
rect 7374 8300 7430 8303
rect 7482 8300 7538 8303
rect 7590 8300 9677 8303
rect 9729 8300 9785 8303
rect 9837 8300 9893 8303
rect 9945 8300 10001 8303
rect 10053 8300 10109 8303
rect 10161 8300 10217 8303
rect 10269 8300 10325 8303
rect 10377 8300 10433 8303
rect 10485 8300 10541 8303
rect 10593 8300 10649 8303
rect 10701 8300 10757 8303
rect 10809 8300 10865 8303
rect 10917 8300 10973 8303
rect 11025 8300 11081 8303
rect 11133 8300 11189 8303
rect 11241 8300 11297 8303
rect 11349 8300 11405 8303
rect 11457 8300 11481 8303
rect 1481 8254 1494 8300
rect 11468 8254 11481 8300
rect 1481 8251 3433 8254
rect 3485 8251 3541 8254
rect 3593 8251 3649 8254
rect 3701 8251 3757 8254
rect 3809 8251 3865 8254
rect 3917 8251 3973 8254
rect 4025 8251 4081 8254
rect 4133 8251 4189 8254
rect 4241 8251 4297 8254
rect 4349 8251 4405 8254
rect 4457 8251 4513 8254
rect 4565 8251 4621 8254
rect 4673 8251 4729 8254
rect 4781 8251 4837 8254
rect 4889 8251 4945 8254
rect 4997 8251 5053 8254
rect 5105 8251 5161 8254
rect 5213 8251 6566 8254
rect 6618 8251 6674 8254
rect 6726 8251 6782 8254
rect 6834 8251 6890 8254
rect 6942 8251 6998 8254
rect 7050 8251 7106 8254
rect 7158 8251 7214 8254
rect 7266 8251 7322 8254
rect 7374 8251 7430 8254
rect 7482 8251 7538 8254
rect 7590 8251 9677 8254
rect 9729 8251 9785 8254
rect 9837 8251 9893 8254
rect 9945 8251 10001 8254
rect 10053 8251 10109 8254
rect 10161 8251 10217 8254
rect 10269 8251 10325 8254
rect 10377 8251 10433 8254
rect 10485 8251 10541 8254
rect 10593 8251 10649 8254
rect 10701 8251 10757 8254
rect 10809 8251 10865 8254
rect 10917 8251 10973 8254
rect 11025 8251 11081 8254
rect 11133 8251 11189 8254
rect 11241 8251 11297 8254
rect 11349 8251 11405 8254
rect 11457 8251 11481 8254
rect 1481 8239 11481 8251
rect 1481 8059 11481 8071
rect 1481 8056 1505 8059
rect 1557 8056 1613 8059
rect 1665 8056 1721 8059
rect 1773 8056 1829 8059
rect 1881 8056 1937 8059
rect 1989 8056 2045 8059
rect 2097 8056 2153 8059
rect 2205 8056 2261 8059
rect 2313 8056 2369 8059
rect 2421 8056 2477 8059
rect 2529 8056 2585 8059
rect 2637 8056 2693 8059
rect 2745 8056 2801 8059
rect 2853 8056 2909 8059
rect 2961 8056 3017 8059
rect 3069 8056 3125 8059
rect 3177 8056 3233 8059
rect 3285 8056 5372 8059
rect 5424 8056 5480 8059
rect 5532 8056 5588 8059
rect 5640 8056 5696 8059
rect 5748 8056 5804 8059
rect 5856 8056 5912 8059
rect 5964 8056 6020 8059
rect 6072 8056 6128 8059
rect 6180 8056 6236 8059
rect 6288 8056 6344 8059
rect 6396 8056 7749 8059
rect 7801 8056 7857 8059
rect 7909 8056 7965 8059
rect 8017 8056 8073 8059
rect 8125 8056 8181 8059
rect 8233 8056 8289 8059
rect 8341 8056 8397 8059
rect 8449 8056 8505 8059
rect 8557 8056 8613 8059
rect 8665 8056 8721 8059
rect 8773 8056 8829 8059
rect 8881 8056 8937 8059
rect 8989 8056 9045 8059
rect 9097 8056 9153 8059
rect 9205 8056 9261 8059
rect 9313 8056 9369 8059
rect 9421 8056 9477 8059
rect 9529 8056 11481 8059
rect 1481 8010 1494 8056
rect 11468 8010 11481 8056
rect 1481 8007 1505 8010
rect 1557 8007 1613 8010
rect 1665 8007 1721 8010
rect 1773 8007 1829 8010
rect 1881 8007 1937 8010
rect 1989 8007 2045 8010
rect 2097 8007 2153 8010
rect 2205 8007 2261 8010
rect 2313 8007 2369 8010
rect 2421 8007 2477 8010
rect 2529 8007 2585 8010
rect 2637 8007 2693 8010
rect 2745 8007 2801 8010
rect 2853 8007 2909 8010
rect 2961 8007 3017 8010
rect 3069 8007 3125 8010
rect 3177 8007 3233 8010
rect 3285 8007 5372 8010
rect 5424 8007 5480 8010
rect 5532 8007 5588 8010
rect 5640 8007 5696 8010
rect 5748 8007 5804 8010
rect 5856 8007 5912 8010
rect 5964 8007 6020 8010
rect 6072 8007 6128 8010
rect 6180 8007 6236 8010
rect 6288 8007 6344 8010
rect 6396 8007 7749 8010
rect 7801 8007 7857 8010
rect 7909 8007 7965 8010
rect 8017 8007 8073 8010
rect 8125 8007 8181 8010
rect 8233 8007 8289 8010
rect 8341 8007 8397 8010
rect 8449 8007 8505 8010
rect 8557 8007 8613 8010
rect 8665 8007 8721 8010
rect 8773 8007 8829 8010
rect 8881 8007 8937 8010
rect 8989 8007 9045 8010
rect 9097 8007 9153 8010
rect 9205 8007 9261 8010
rect 9313 8007 9369 8010
rect 9421 8007 9477 8010
rect 9529 8007 11481 8010
rect 1481 7995 11481 8007
rect 1481 7815 11481 7827
rect 1481 7812 3433 7815
rect 3485 7812 3541 7815
rect 3593 7812 3649 7815
rect 3701 7812 3757 7815
rect 3809 7812 3865 7815
rect 3917 7812 3973 7815
rect 4025 7812 4081 7815
rect 4133 7812 4189 7815
rect 4241 7812 4297 7815
rect 4349 7812 4405 7815
rect 4457 7812 4513 7815
rect 4565 7812 4621 7815
rect 4673 7812 4729 7815
rect 4781 7812 4837 7815
rect 4889 7812 4945 7815
rect 4997 7812 5053 7815
rect 5105 7812 5161 7815
rect 5213 7812 6566 7815
rect 6618 7812 6674 7815
rect 6726 7812 6782 7815
rect 6834 7812 6890 7815
rect 6942 7812 6998 7815
rect 7050 7812 7106 7815
rect 7158 7812 7214 7815
rect 7266 7812 7322 7815
rect 7374 7812 7430 7815
rect 7482 7812 7538 7815
rect 7590 7812 9677 7815
rect 9729 7812 9785 7815
rect 9837 7812 9893 7815
rect 9945 7812 10001 7815
rect 10053 7812 10109 7815
rect 10161 7812 10217 7815
rect 10269 7812 10325 7815
rect 10377 7812 10433 7815
rect 10485 7812 10541 7815
rect 10593 7812 10649 7815
rect 10701 7812 10757 7815
rect 10809 7812 10865 7815
rect 10917 7812 10973 7815
rect 11025 7812 11081 7815
rect 11133 7812 11189 7815
rect 11241 7812 11297 7815
rect 11349 7812 11405 7815
rect 11457 7812 11481 7815
rect 1481 7766 1494 7812
rect 11468 7766 11481 7812
rect 1481 7763 3433 7766
rect 3485 7763 3541 7766
rect 3593 7763 3649 7766
rect 3701 7763 3757 7766
rect 3809 7763 3865 7766
rect 3917 7763 3973 7766
rect 4025 7763 4081 7766
rect 4133 7763 4189 7766
rect 4241 7763 4297 7766
rect 4349 7763 4405 7766
rect 4457 7763 4513 7766
rect 4565 7763 4621 7766
rect 4673 7763 4729 7766
rect 4781 7763 4837 7766
rect 4889 7763 4945 7766
rect 4997 7763 5053 7766
rect 5105 7763 5161 7766
rect 5213 7763 6566 7766
rect 6618 7763 6674 7766
rect 6726 7763 6782 7766
rect 6834 7763 6890 7766
rect 6942 7763 6998 7766
rect 7050 7763 7106 7766
rect 7158 7763 7214 7766
rect 7266 7763 7322 7766
rect 7374 7763 7430 7766
rect 7482 7763 7538 7766
rect 7590 7763 9677 7766
rect 9729 7763 9785 7766
rect 9837 7763 9893 7766
rect 9945 7763 10001 7766
rect 10053 7763 10109 7766
rect 10161 7763 10217 7766
rect 10269 7763 10325 7766
rect 10377 7763 10433 7766
rect 10485 7763 10541 7766
rect 10593 7763 10649 7766
rect 10701 7763 10757 7766
rect 10809 7763 10865 7766
rect 10917 7763 10973 7766
rect 11025 7763 11081 7766
rect 11133 7763 11189 7766
rect 11241 7763 11297 7766
rect 11349 7763 11405 7766
rect 11457 7763 11481 7766
rect 1481 7751 11481 7763
rect 1481 7571 11481 7583
rect 1481 7568 1505 7571
rect 1557 7568 1613 7571
rect 1665 7568 1721 7571
rect 1773 7568 1829 7571
rect 1881 7568 1937 7571
rect 1989 7568 2045 7571
rect 2097 7568 2153 7571
rect 2205 7568 2261 7571
rect 2313 7568 2369 7571
rect 2421 7568 2477 7571
rect 2529 7568 2585 7571
rect 2637 7568 2693 7571
rect 2745 7568 2801 7571
rect 2853 7568 2909 7571
rect 2961 7568 3017 7571
rect 3069 7568 3125 7571
rect 3177 7568 3233 7571
rect 3285 7568 5372 7571
rect 5424 7568 5480 7571
rect 5532 7568 5588 7571
rect 5640 7568 5696 7571
rect 5748 7568 5804 7571
rect 5856 7568 5912 7571
rect 5964 7568 6020 7571
rect 6072 7568 6128 7571
rect 6180 7568 6236 7571
rect 6288 7568 6344 7571
rect 6396 7568 7749 7571
rect 7801 7568 7857 7571
rect 7909 7568 7965 7571
rect 8017 7568 8073 7571
rect 8125 7568 8181 7571
rect 8233 7568 8289 7571
rect 8341 7568 8397 7571
rect 8449 7568 8505 7571
rect 8557 7568 8613 7571
rect 8665 7568 8721 7571
rect 8773 7568 8829 7571
rect 8881 7568 8937 7571
rect 8989 7568 9045 7571
rect 9097 7568 9153 7571
rect 9205 7568 9261 7571
rect 9313 7568 9369 7571
rect 9421 7568 9477 7571
rect 9529 7568 11481 7571
rect 1481 7522 1494 7568
rect 11468 7522 11481 7568
rect 1481 7519 1505 7522
rect 1557 7519 1613 7522
rect 1665 7519 1721 7522
rect 1773 7519 1829 7522
rect 1881 7519 1937 7522
rect 1989 7519 2045 7522
rect 2097 7519 2153 7522
rect 2205 7519 2261 7522
rect 2313 7519 2369 7522
rect 2421 7519 2477 7522
rect 2529 7519 2585 7522
rect 2637 7519 2693 7522
rect 2745 7519 2801 7522
rect 2853 7519 2909 7522
rect 2961 7519 3017 7522
rect 3069 7519 3125 7522
rect 3177 7519 3233 7522
rect 3285 7519 5372 7522
rect 5424 7519 5480 7522
rect 5532 7519 5588 7522
rect 5640 7519 5696 7522
rect 5748 7519 5804 7522
rect 5856 7519 5912 7522
rect 5964 7519 6020 7522
rect 6072 7519 6128 7522
rect 6180 7519 6236 7522
rect 6288 7519 6344 7522
rect 6396 7519 7749 7522
rect 7801 7519 7857 7522
rect 7909 7519 7965 7522
rect 8017 7519 8073 7522
rect 8125 7519 8181 7522
rect 8233 7519 8289 7522
rect 8341 7519 8397 7522
rect 8449 7519 8505 7522
rect 8557 7519 8613 7522
rect 8665 7519 8721 7522
rect 8773 7519 8829 7522
rect 8881 7519 8937 7522
rect 8989 7519 9045 7522
rect 9097 7519 9153 7522
rect 9205 7519 9261 7522
rect 9313 7519 9369 7522
rect 9421 7519 9477 7522
rect 9529 7519 11481 7522
rect 1481 7507 11481 7519
rect 1213 7391 1413 7418
rect 1213 7339 1233 7391
rect 1285 7339 1341 7391
rect 1393 7339 1413 7391
rect 11549 7418 11560 12064
rect 11706 12035 11749 12064
rect 11729 11983 11749 12035
rect 11706 11927 11749 11983
rect 11729 11875 11749 11927
rect 11706 11819 11749 11875
rect 11729 11767 11749 11819
rect 11706 11711 11749 11767
rect 11729 11659 11749 11711
rect 11706 11603 11749 11659
rect 11729 11551 11749 11603
rect 11706 11495 11749 11551
rect 11729 11443 11749 11495
rect 11706 11387 11749 11443
rect 11729 11335 11749 11387
rect 11706 11279 11749 11335
rect 11729 11227 11749 11279
rect 11706 11171 11749 11227
rect 11729 11119 11749 11171
rect 11706 11063 11749 11119
rect 11729 11011 11749 11063
rect 11706 10955 11749 11011
rect 11729 10903 11749 10955
rect 11706 10847 11749 10903
rect 11729 10795 11749 10847
rect 11706 10739 11749 10795
rect 11729 10687 11749 10739
rect 11706 10631 11749 10687
rect 11729 10579 11749 10631
rect 11706 10523 11749 10579
rect 11729 10471 11749 10523
rect 11706 10415 11749 10471
rect 11729 10363 11749 10415
rect 11706 10307 11749 10363
rect 11729 10255 11749 10307
rect 11706 10199 11749 10255
rect 11729 10147 11749 10199
rect 11706 10091 11749 10147
rect 11729 10039 11749 10091
rect 11706 9983 11749 10039
rect 11729 9931 11749 9983
rect 11706 9875 11749 9931
rect 11729 9823 11749 9875
rect 11706 9767 11749 9823
rect 11729 9715 11749 9767
rect 11706 9659 11749 9715
rect 11729 9607 11749 9659
rect 11706 9551 11749 9607
rect 11729 9499 11749 9551
rect 11706 9443 11749 9499
rect 11729 9391 11749 9443
rect 11706 9335 11749 9391
rect 11729 9283 11749 9335
rect 11706 9227 11749 9283
rect 11729 9175 11749 9227
rect 11706 9119 11749 9175
rect 11729 9067 11749 9119
rect 11706 9011 11749 9067
rect 11729 8959 11749 9011
rect 11706 8903 11749 8959
rect 11729 8851 11749 8903
rect 11706 8795 11749 8851
rect 11729 8743 11749 8795
rect 11706 8687 11749 8743
rect 11729 8635 11749 8687
rect 11706 8579 11749 8635
rect 11729 8527 11749 8579
rect 11706 8471 11749 8527
rect 11729 8419 11749 8471
rect 11706 8363 11749 8419
rect 11729 8311 11749 8363
rect 11706 8255 11749 8311
rect 11729 8203 11749 8255
rect 11706 8147 11749 8203
rect 11729 8095 11749 8147
rect 11706 8039 11749 8095
rect 11729 7987 11749 8039
rect 11706 7931 11749 7987
rect 11729 7879 11749 7931
rect 11706 7823 11749 7879
rect 11729 7771 11749 7823
rect 11706 7715 11749 7771
rect 11729 7663 11749 7715
rect 11706 7607 11749 7663
rect 11729 7555 11749 7607
rect 11706 7499 11749 7555
rect 11729 7447 11749 7499
rect 11706 7418 11749 7447
rect 11549 7391 11749 7418
rect 11549 7339 11569 7391
rect 11621 7339 11677 7391
rect 11729 7339 11749 7391
rect 1213 7176 1413 7339
rect 1481 7327 11481 7339
rect 1481 7324 3433 7327
rect 3485 7324 3541 7327
rect 3593 7324 3649 7327
rect 3701 7324 3757 7327
rect 3809 7324 3865 7327
rect 3917 7324 3973 7327
rect 4025 7324 4081 7327
rect 4133 7324 4189 7327
rect 4241 7324 4297 7327
rect 4349 7324 4405 7327
rect 4457 7324 4513 7327
rect 4565 7324 4621 7327
rect 4673 7324 4729 7327
rect 4781 7324 4837 7327
rect 4889 7324 4945 7327
rect 4997 7324 5053 7327
rect 5105 7324 5161 7327
rect 5213 7324 6566 7327
rect 6618 7324 6674 7327
rect 6726 7324 6782 7327
rect 6834 7324 6890 7327
rect 6942 7324 6998 7327
rect 7050 7324 7106 7327
rect 7158 7324 7214 7327
rect 7266 7324 7322 7327
rect 7374 7324 7430 7327
rect 7482 7324 7538 7327
rect 7590 7324 9677 7327
rect 9729 7324 9785 7327
rect 9837 7324 9893 7327
rect 9945 7324 10001 7327
rect 10053 7324 10109 7327
rect 10161 7324 10217 7327
rect 10269 7324 10325 7327
rect 10377 7324 10433 7327
rect 10485 7324 10541 7327
rect 10593 7324 10649 7327
rect 10701 7324 10757 7327
rect 10809 7324 10865 7327
rect 10917 7324 10973 7327
rect 11025 7324 11081 7327
rect 11133 7324 11189 7327
rect 11241 7324 11297 7327
rect 11349 7324 11405 7327
rect 11457 7324 11481 7327
rect 1481 7278 1494 7324
rect 11468 7278 11481 7324
rect 1481 7275 3433 7278
rect 3485 7275 3541 7278
rect 3593 7275 3649 7278
rect 3701 7275 3757 7278
rect 3809 7275 3865 7278
rect 3917 7275 3973 7278
rect 4025 7275 4081 7278
rect 4133 7275 4189 7278
rect 4241 7275 4297 7278
rect 4349 7275 4405 7278
rect 4457 7275 4513 7278
rect 4565 7275 4621 7278
rect 4673 7275 4729 7278
rect 4781 7275 4837 7278
rect 4889 7275 4945 7278
rect 4997 7275 5053 7278
rect 5105 7275 5161 7278
rect 5213 7275 6566 7278
rect 6618 7275 6674 7278
rect 6726 7275 6782 7278
rect 6834 7275 6890 7278
rect 6942 7275 6998 7278
rect 7050 7275 7106 7278
rect 7158 7275 7214 7278
rect 7266 7275 7322 7278
rect 7374 7275 7430 7278
rect 7482 7275 7538 7278
rect 7590 7275 9677 7278
rect 9729 7275 9785 7278
rect 9837 7275 9893 7278
rect 9945 7275 10001 7278
rect 10053 7275 10109 7278
rect 10161 7275 10217 7278
rect 10269 7275 10325 7278
rect 10377 7275 10433 7278
rect 10485 7275 10541 7278
rect 10593 7275 10649 7278
rect 10701 7275 10757 7278
rect 10809 7275 10865 7278
rect 10917 7275 10973 7278
rect 11025 7275 11081 7278
rect 11133 7275 11189 7278
rect 11241 7275 11297 7278
rect 11349 7275 11405 7278
rect 11457 7275 11481 7278
rect 1481 7263 11481 7275
rect 11549 7176 11749 7339
rect 1213 6976 11749 7176
rect 12001 6897 12012 12585
rect 950 6885 12012 6897
rect 950 6878 1505 6885
rect 1557 6878 1613 6885
rect 1665 6878 1721 6885
rect 1773 6878 1829 6885
rect 1881 6878 1937 6885
rect 1989 6878 2045 6885
rect 2097 6878 2153 6885
rect 2205 6878 2261 6885
rect 2313 6878 2369 6885
rect 2421 6878 2477 6885
rect 2529 6878 2585 6885
rect 2637 6878 2693 6885
rect 2745 6878 2801 6885
rect 2853 6878 2909 6885
rect 2961 6878 3017 6885
rect 3069 6878 3125 6885
rect 3177 6878 3233 6885
rect 3285 6878 5372 6885
rect 5424 6878 5480 6885
rect 5532 6878 5588 6885
rect 5640 6878 5696 6885
rect 5748 6878 5804 6885
rect 5856 6878 5912 6885
rect 5964 6878 6020 6885
rect 6072 6878 6128 6885
rect 6180 6878 6236 6885
rect 6288 6878 6344 6885
rect 6396 6878 7749 6885
rect 7801 6878 7857 6885
rect 7909 6878 7965 6885
rect 8017 6878 8073 6885
rect 8125 6878 8181 6885
rect 8233 6878 8289 6885
rect 8341 6878 8397 6885
rect 8449 6878 8505 6885
rect 8557 6878 8613 6885
rect 8665 6878 8721 6885
rect 8773 6878 8829 6885
rect 8881 6878 8937 6885
rect 8989 6878 9045 6885
rect 9097 6878 9153 6885
rect 9205 6878 9261 6885
rect 9313 6878 9369 6885
rect 9421 6878 9477 6885
rect 9529 6878 12012 6885
rect 950 6732 1058 6878
rect 11904 6732 12012 6878
rect 950 6725 1505 6732
rect 1557 6725 1613 6732
rect 1665 6725 1721 6732
rect 1773 6725 1829 6732
rect 1881 6725 1937 6732
rect 1989 6725 2045 6732
rect 2097 6725 2153 6732
rect 2205 6725 2261 6732
rect 2313 6725 2369 6732
rect 2421 6725 2477 6732
rect 2529 6725 2585 6732
rect 2637 6725 2693 6732
rect 2745 6725 2801 6732
rect 2853 6725 2909 6732
rect 2961 6725 3017 6732
rect 3069 6725 3125 6732
rect 3177 6725 3233 6732
rect 3285 6725 5372 6732
rect 5424 6725 5480 6732
rect 5532 6725 5588 6732
rect 5640 6725 5696 6732
rect 5748 6725 5804 6732
rect 5856 6725 5912 6732
rect 5964 6725 6020 6732
rect 6072 6725 6128 6732
rect 6180 6725 6236 6732
rect 6288 6725 6344 6732
rect 6396 6725 7749 6732
rect 7801 6725 7857 6732
rect 7909 6725 7965 6732
rect 8017 6725 8073 6732
rect 8125 6725 8181 6732
rect 8233 6725 8289 6732
rect 8341 6725 8397 6732
rect 8449 6725 8505 6732
rect 8557 6725 8613 6732
rect 8665 6725 8721 6732
rect 8773 6725 8829 6732
rect 8881 6725 8937 6732
rect 8989 6725 9045 6732
rect 9097 6725 9153 6732
rect 9205 6725 9261 6732
rect 9313 6725 9369 6732
rect 9421 6725 9477 6732
rect 9529 6725 12012 6732
rect 950 6713 12012 6725
rect 950 1011 961 6713
rect 1213 6434 11749 6634
rect 1213 6271 1413 6434
rect 1481 6335 11481 6347
rect 1481 6332 3433 6335
rect 3485 6332 3541 6335
rect 3593 6332 3649 6335
rect 3701 6332 3757 6335
rect 3809 6332 3865 6335
rect 3917 6332 3973 6335
rect 4025 6332 4081 6335
rect 4133 6332 4189 6335
rect 4241 6332 4297 6335
rect 4349 6332 4405 6335
rect 4457 6332 4513 6335
rect 4565 6332 4621 6335
rect 4673 6332 4729 6335
rect 4781 6332 4837 6335
rect 4889 6332 4945 6335
rect 4997 6332 5053 6335
rect 5105 6332 5161 6335
rect 5213 6332 6566 6335
rect 6618 6332 6674 6335
rect 6726 6332 6782 6335
rect 6834 6332 6890 6335
rect 6942 6332 6998 6335
rect 7050 6332 7106 6335
rect 7158 6332 7214 6335
rect 7266 6332 7322 6335
rect 7374 6332 7430 6335
rect 7482 6332 7538 6335
rect 7590 6332 9677 6335
rect 9729 6332 9785 6335
rect 9837 6332 9893 6335
rect 9945 6332 10001 6335
rect 10053 6332 10109 6335
rect 10161 6332 10217 6335
rect 10269 6332 10325 6335
rect 10377 6332 10433 6335
rect 10485 6332 10541 6335
rect 10593 6332 10649 6335
rect 10701 6332 10757 6335
rect 10809 6332 10865 6335
rect 10917 6332 10973 6335
rect 11025 6332 11081 6335
rect 11133 6332 11189 6335
rect 11241 6332 11297 6335
rect 11349 6332 11405 6335
rect 11457 6332 11481 6335
rect 1481 6286 1494 6332
rect 11468 6286 11481 6332
rect 1481 6283 3433 6286
rect 3485 6283 3541 6286
rect 3593 6283 3649 6286
rect 3701 6283 3757 6286
rect 3809 6283 3865 6286
rect 3917 6283 3973 6286
rect 4025 6283 4081 6286
rect 4133 6283 4189 6286
rect 4241 6283 4297 6286
rect 4349 6283 4405 6286
rect 4457 6283 4513 6286
rect 4565 6283 4621 6286
rect 4673 6283 4729 6286
rect 4781 6283 4837 6286
rect 4889 6283 4945 6286
rect 4997 6283 5053 6286
rect 5105 6283 5161 6286
rect 5213 6283 6566 6286
rect 6618 6283 6674 6286
rect 6726 6283 6782 6286
rect 6834 6283 6890 6286
rect 6942 6283 6998 6286
rect 7050 6283 7106 6286
rect 7158 6283 7214 6286
rect 7266 6283 7322 6286
rect 7374 6283 7430 6286
rect 7482 6283 7538 6286
rect 7590 6283 9677 6286
rect 9729 6283 9785 6286
rect 9837 6283 9893 6286
rect 9945 6283 10001 6286
rect 10053 6283 10109 6286
rect 10161 6283 10217 6286
rect 10269 6283 10325 6286
rect 10377 6283 10433 6286
rect 10485 6283 10541 6286
rect 10593 6283 10649 6286
rect 10701 6283 10757 6286
rect 10809 6283 10865 6286
rect 10917 6283 10973 6286
rect 11025 6283 11081 6286
rect 11133 6283 11189 6286
rect 11241 6283 11297 6286
rect 11349 6283 11405 6286
rect 11457 6283 11481 6286
rect 1481 6271 11481 6283
rect 11549 6271 11749 6434
rect 1213 6219 1233 6271
rect 1285 6219 1341 6271
rect 1393 6219 1413 6271
rect 1213 6192 1413 6219
rect 1213 6163 1256 6192
rect 1213 6111 1233 6163
rect 1213 6055 1256 6111
rect 1213 6003 1233 6055
rect 1213 5947 1256 6003
rect 1213 5895 1233 5947
rect 1213 5839 1256 5895
rect 1213 5787 1233 5839
rect 1213 5731 1256 5787
rect 1213 5679 1233 5731
rect 1213 5623 1256 5679
rect 1213 5571 1233 5623
rect 1213 5515 1256 5571
rect 1213 5463 1233 5515
rect 1213 5407 1256 5463
rect 1213 5355 1233 5407
rect 1213 5299 1256 5355
rect 1213 5247 1233 5299
rect 1213 5191 1256 5247
rect 1213 5139 1233 5191
rect 1213 5083 1256 5139
rect 1213 5031 1233 5083
rect 1213 4975 1256 5031
rect 1213 4923 1233 4975
rect 1213 4867 1256 4923
rect 1213 4815 1233 4867
rect 1213 4759 1256 4815
rect 1213 4707 1233 4759
rect 1213 4651 1256 4707
rect 1213 4599 1233 4651
rect 1213 4543 1256 4599
rect 1213 4491 1233 4543
rect 1213 4435 1256 4491
rect 1213 4383 1233 4435
rect 1213 4327 1256 4383
rect 1213 4275 1233 4327
rect 1213 4219 1256 4275
rect 1213 4167 1233 4219
rect 1213 4111 1256 4167
rect 1213 4059 1233 4111
rect 1213 4003 1256 4059
rect 1213 3951 1233 4003
rect 1213 3895 1256 3951
rect 1213 3843 1233 3895
rect 1213 3787 1256 3843
rect 1213 3735 1233 3787
rect 1213 3679 1256 3735
rect 1213 3627 1233 3679
rect 1213 3571 1256 3627
rect 1213 3519 1233 3571
rect 1213 3463 1256 3519
rect 1213 3411 1233 3463
rect 1213 3355 1256 3411
rect 1213 3303 1233 3355
rect 1213 3247 1256 3303
rect 1213 3195 1233 3247
rect 1213 3139 1256 3195
rect 1213 3087 1233 3139
rect 1213 3031 1256 3087
rect 1213 2979 1233 3031
rect 1213 2923 1256 2979
rect 1213 2871 1233 2923
rect 1213 2815 1256 2871
rect 1213 2763 1233 2815
rect 1213 2707 1256 2763
rect 1213 2655 1233 2707
rect 1213 2599 1256 2655
rect 1213 2547 1233 2599
rect 1213 2491 1256 2547
rect 1213 2439 1233 2491
rect 1213 2383 1256 2439
rect 1213 2331 1233 2383
rect 1213 2275 1256 2331
rect 1213 2223 1233 2275
rect 1213 2167 1256 2223
rect 1213 2115 1233 2167
rect 1213 2059 1256 2115
rect 1213 2007 1233 2059
rect 1213 1951 1256 2007
rect 1213 1899 1233 1951
rect 1213 1843 1256 1899
rect 1213 1791 1233 1843
rect 1213 1735 1256 1791
rect 1213 1683 1233 1735
rect 1213 1627 1256 1683
rect 1213 1575 1233 1627
rect 1213 1546 1256 1575
rect 1402 1546 1413 6192
rect 11549 6219 11569 6271
rect 11621 6219 11677 6271
rect 11729 6219 11749 6271
rect 11549 6192 11749 6219
rect 1481 6091 11481 6103
rect 1481 6088 1505 6091
rect 1557 6088 1613 6091
rect 1665 6088 1721 6091
rect 1773 6088 1829 6091
rect 1881 6088 1937 6091
rect 1989 6088 2045 6091
rect 2097 6088 2153 6091
rect 2205 6088 2261 6091
rect 2313 6088 2369 6091
rect 2421 6088 2477 6091
rect 2529 6088 2585 6091
rect 2637 6088 2693 6091
rect 2745 6088 2801 6091
rect 2853 6088 2909 6091
rect 2961 6088 3017 6091
rect 3069 6088 3125 6091
rect 3177 6088 3233 6091
rect 3285 6088 5372 6091
rect 5424 6088 5480 6091
rect 5532 6088 5588 6091
rect 5640 6088 5696 6091
rect 5748 6088 5804 6091
rect 5856 6088 5912 6091
rect 5964 6088 6020 6091
rect 6072 6088 6128 6091
rect 6180 6088 6236 6091
rect 6288 6088 6344 6091
rect 6396 6088 7749 6091
rect 7801 6088 7857 6091
rect 7909 6088 7965 6091
rect 8017 6088 8073 6091
rect 8125 6088 8181 6091
rect 8233 6088 8289 6091
rect 8341 6088 8397 6091
rect 8449 6088 8505 6091
rect 8557 6088 8613 6091
rect 8665 6088 8721 6091
rect 8773 6088 8829 6091
rect 8881 6088 8937 6091
rect 8989 6088 9045 6091
rect 9097 6088 9153 6091
rect 9205 6088 9261 6091
rect 9313 6088 9369 6091
rect 9421 6088 9477 6091
rect 9529 6088 11481 6091
rect 1481 6042 1494 6088
rect 11468 6042 11481 6088
rect 1481 6039 1505 6042
rect 1557 6039 1613 6042
rect 1665 6039 1721 6042
rect 1773 6039 1829 6042
rect 1881 6039 1937 6042
rect 1989 6039 2045 6042
rect 2097 6039 2153 6042
rect 2205 6039 2261 6042
rect 2313 6039 2369 6042
rect 2421 6039 2477 6042
rect 2529 6039 2585 6042
rect 2637 6039 2693 6042
rect 2745 6039 2801 6042
rect 2853 6039 2909 6042
rect 2961 6039 3017 6042
rect 3069 6039 3125 6042
rect 3177 6039 3233 6042
rect 3285 6039 5372 6042
rect 5424 6039 5480 6042
rect 5532 6039 5588 6042
rect 5640 6039 5696 6042
rect 5748 6039 5804 6042
rect 5856 6039 5912 6042
rect 5964 6039 6020 6042
rect 6072 6039 6128 6042
rect 6180 6039 6236 6042
rect 6288 6039 6344 6042
rect 6396 6039 7749 6042
rect 7801 6039 7857 6042
rect 7909 6039 7965 6042
rect 8017 6039 8073 6042
rect 8125 6039 8181 6042
rect 8233 6039 8289 6042
rect 8341 6039 8397 6042
rect 8449 6039 8505 6042
rect 8557 6039 8613 6042
rect 8665 6039 8721 6042
rect 8773 6039 8829 6042
rect 8881 6039 8937 6042
rect 8989 6039 9045 6042
rect 9097 6039 9153 6042
rect 9205 6039 9261 6042
rect 9313 6039 9369 6042
rect 9421 6039 9477 6042
rect 9529 6039 11481 6042
rect 1481 6027 11481 6039
rect 1481 5847 11481 5859
rect 1481 5844 3433 5847
rect 3485 5844 3541 5847
rect 3593 5844 3649 5847
rect 3701 5844 3757 5847
rect 3809 5844 3865 5847
rect 3917 5844 3973 5847
rect 4025 5844 4081 5847
rect 4133 5844 4189 5847
rect 4241 5844 4297 5847
rect 4349 5844 4405 5847
rect 4457 5844 4513 5847
rect 4565 5844 4621 5847
rect 4673 5844 4729 5847
rect 4781 5844 4837 5847
rect 4889 5844 4945 5847
rect 4997 5844 5053 5847
rect 5105 5844 5161 5847
rect 5213 5844 6566 5847
rect 6618 5844 6674 5847
rect 6726 5844 6782 5847
rect 6834 5844 6890 5847
rect 6942 5844 6998 5847
rect 7050 5844 7106 5847
rect 7158 5844 7214 5847
rect 7266 5844 7322 5847
rect 7374 5844 7430 5847
rect 7482 5844 7538 5847
rect 7590 5844 9677 5847
rect 9729 5844 9785 5847
rect 9837 5844 9893 5847
rect 9945 5844 10001 5847
rect 10053 5844 10109 5847
rect 10161 5844 10217 5847
rect 10269 5844 10325 5847
rect 10377 5844 10433 5847
rect 10485 5844 10541 5847
rect 10593 5844 10649 5847
rect 10701 5844 10757 5847
rect 10809 5844 10865 5847
rect 10917 5844 10973 5847
rect 11025 5844 11081 5847
rect 11133 5844 11189 5847
rect 11241 5844 11297 5847
rect 11349 5844 11405 5847
rect 11457 5844 11481 5847
rect 1481 5798 1494 5844
rect 11468 5798 11481 5844
rect 1481 5795 3433 5798
rect 3485 5795 3541 5798
rect 3593 5795 3649 5798
rect 3701 5795 3757 5798
rect 3809 5795 3865 5798
rect 3917 5795 3973 5798
rect 4025 5795 4081 5798
rect 4133 5795 4189 5798
rect 4241 5795 4297 5798
rect 4349 5795 4405 5798
rect 4457 5795 4513 5798
rect 4565 5795 4621 5798
rect 4673 5795 4729 5798
rect 4781 5795 4837 5798
rect 4889 5795 4945 5798
rect 4997 5795 5053 5798
rect 5105 5795 5161 5798
rect 5213 5795 6566 5798
rect 6618 5795 6674 5798
rect 6726 5795 6782 5798
rect 6834 5795 6890 5798
rect 6942 5795 6998 5798
rect 7050 5795 7106 5798
rect 7158 5795 7214 5798
rect 7266 5795 7322 5798
rect 7374 5795 7430 5798
rect 7482 5795 7538 5798
rect 7590 5795 9677 5798
rect 9729 5795 9785 5798
rect 9837 5795 9893 5798
rect 9945 5795 10001 5798
rect 10053 5795 10109 5798
rect 10161 5795 10217 5798
rect 10269 5795 10325 5798
rect 10377 5795 10433 5798
rect 10485 5795 10541 5798
rect 10593 5795 10649 5798
rect 10701 5795 10757 5798
rect 10809 5795 10865 5798
rect 10917 5795 10973 5798
rect 11025 5795 11081 5798
rect 11133 5795 11189 5798
rect 11241 5795 11297 5798
rect 11349 5795 11405 5798
rect 11457 5795 11481 5798
rect 1481 5783 11481 5795
rect 1481 5603 11481 5615
rect 1481 5600 1505 5603
rect 1557 5600 1613 5603
rect 1665 5600 1721 5603
rect 1773 5600 1829 5603
rect 1881 5600 1937 5603
rect 1989 5600 2045 5603
rect 2097 5600 2153 5603
rect 2205 5600 2261 5603
rect 2313 5600 2369 5603
rect 2421 5600 2477 5603
rect 2529 5600 2585 5603
rect 2637 5600 2693 5603
rect 2745 5600 2801 5603
rect 2853 5600 2909 5603
rect 2961 5600 3017 5603
rect 3069 5600 3125 5603
rect 3177 5600 3233 5603
rect 3285 5600 5372 5603
rect 5424 5600 5480 5603
rect 5532 5600 5588 5603
rect 5640 5600 5696 5603
rect 5748 5600 5804 5603
rect 5856 5600 5912 5603
rect 5964 5600 6020 5603
rect 6072 5600 6128 5603
rect 6180 5600 6236 5603
rect 6288 5600 6344 5603
rect 6396 5600 7749 5603
rect 7801 5600 7857 5603
rect 7909 5600 7965 5603
rect 8017 5600 8073 5603
rect 8125 5600 8181 5603
rect 8233 5600 8289 5603
rect 8341 5600 8397 5603
rect 8449 5600 8505 5603
rect 8557 5600 8613 5603
rect 8665 5600 8721 5603
rect 8773 5600 8829 5603
rect 8881 5600 8937 5603
rect 8989 5600 9045 5603
rect 9097 5600 9153 5603
rect 9205 5600 9261 5603
rect 9313 5600 9369 5603
rect 9421 5600 9477 5603
rect 9529 5600 11481 5603
rect 1481 5554 1494 5600
rect 11468 5554 11481 5600
rect 1481 5551 1505 5554
rect 1557 5551 1613 5554
rect 1665 5551 1721 5554
rect 1773 5551 1829 5554
rect 1881 5551 1937 5554
rect 1989 5551 2045 5554
rect 2097 5551 2153 5554
rect 2205 5551 2261 5554
rect 2313 5551 2369 5554
rect 2421 5551 2477 5554
rect 2529 5551 2585 5554
rect 2637 5551 2693 5554
rect 2745 5551 2801 5554
rect 2853 5551 2909 5554
rect 2961 5551 3017 5554
rect 3069 5551 3125 5554
rect 3177 5551 3233 5554
rect 3285 5551 5372 5554
rect 5424 5551 5480 5554
rect 5532 5551 5588 5554
rect 5640 5551 5696 5554
rect 5748 5551 5804 5554
rect 5856 5551 5912 5554
rect 5964 5551 6020 5554
rect 6072 5551 6128 5554
rect 6180 5551 6236 5554
rect 6288 5551 6344 5554
rect 6396 5551 7749 5554
rect 7801 5551 7857 5554
rect 7909 5551 7965 5554
rect 8017 5551 8073 5554
rect 8125 5551 8181 5554
rect 8233 5551 8289 5554
rect 8341 5551 8397 5554
rect 8449 5551 8505 5554
rect 8557 5551 8613 5554
rect 8665 5551 8721 5554
rect 8773 5551 8829 5554
rect 8881 5551 8937 5554
rect 8989 5551 9045 5554
rect 9097 5551 9153 5554
rect 9205 5551 9261 5554
rect 9313 5551 9369 5554
rect 9421 5551 9477 5554
rect 9529 5551 11481 5554
rect 1481 5539 11481 5551
rect 1481 5359 11481 5371
rect 1481 5356 3433 5359
rect 3485 5356 3541 5359
rect 3593 5356 3649 5359
rect 3701 5356 3757 5359
rect 3809 5356 3865 5359
rect 3917 5356 3973 5359
rect 4025 5356 4081 5359
rect 4133 5356 4189 5359
rect 4241 5356 4297 5359
rect 4349 5356 4405 5359
rect 4457 5356 4513 5359
rect 4565 5356 4621 5359
rect 4673 5356 4729 5359
rect 4781 5356 4837 5359
rect 4889 5356 4945 5359
rect 4997 5356 5053 5359
rect 5105 5356 5161 5359
rect 5213 5356 6566 5359
rect 6618 5356 6674 5359
rect 6726 5356 6782 5359
rect 6834 5356 6890 5359
rect 6942 5356 6998 5359
rect 7050 5356 7106 5359
rect 7158 5356 7214 5359
rect 7266 5356 7322 5359
rect 7374 5356 7430 5359
rect 7482 5356 7538 5359
rect 7590 5356 9677 5359
rect 9729 5356 9785 5359
rect 9837 5356 9893 5359
rect 9945 5356 10001 5359
rect 10053 5356 10109 5359
rect 10161 5356 10217 5359
rect 10269 5356 10325 5359
rect 10377 5356 10433 5359
rect 10485 5356 10541 5359
rect 10593 5356 10649 5359
rect 10701 5356 10757 5359
rect 10809 5356 10865 5359
rect 10917 5356 10973 5359
rect 11025 5356 11081 5359
rect 11133 5356 11189 5359
rect 11241 5356 11297 5359
rect 11349 5356 11405 5359
rect 11457 5356 11481 5359
rect 1481 5310 1494 5356
rect 11468 5310 11481 5356
rect 1481 5307 3433 5310
rect 3485 5307 3541 5310
rect 3593 5307 3649 5310
rect 3701 5307 3757 5310
rect 3809 5307 3865 5310
rect 3917 5307 3973 5310
rect 4025 5307 4081 5310
rect 4133 5307 4189 5310
rect 4241 5307 4297 5310
rect 4349 5307 4405 5310
rect 4457 5307 4513 5310
rect 4565 5307 4621 5310
rect 4673 5307 4729 5310
rect 4781 5307 4837 5310
rect 4889 5307 4945 5310
rect 4997 5307 5053 5310
rect 5105 5307 5161 5310
rect 5213 5307 6566 5310
rect 6618 5307 6674 5310
rect 6726 5307 6782 5310
rect 6834 5307 6890 5310
rect 6942 5307 6998 5310
rect 7050 5307 7106 5310
rect 7158 5307 7214 5310
rect 7266 5307 7322 5310
rect 7374 5307 7430 5310
rect 7482 5307 7538 5310
rect 7590 5307 9677 5310
rect 9729 5307 9785 5310
rect 9837 5307 9893 5310
rect 9945 5307 10001 5310
rect 10053 5307 10109 5310
rect 10161 5307 10217 5310
rect 10269 5307 10325 5310
rect 10377 5307 10433 5310
rect 10485 5307 10541 5310
rect 10593 5307 10649 5310
rect 10701 5307 10757 5310
rect 10809 5307 10865 5310
rect 10917 5307 10973 5310
rect 11025 5307 11081 5310
rect 11133 5307 11189 5310
rect 11241 5307 11297 5310
rect 11349 5307 11405 5310
rect 11457 5307 11481 5310
rect 1481 5295 11481 5307
rect 1481 5115 11481 5127
rect 1481 5112 1505 5115
rect 1557 5112 1613 5115
rect 1665 5112 1721 5115
rect 1773 5112 1829 5115
rect 1881 5112 1937 5115
rect 1989 5112 2045 5115
rect 2097 5112 2153 5115
rect 2205 5112 2261 5115
rect 2313 5112 2369 5115
rect 2421 5112 2477 5115
rect 2529 5112 2585 5115
rect 2637 5112 2693 5115
rect 2745 5112 2801 5115
rect 2853 5112 2909 5115
rect 2961 5112 3017 5115
rect 3069 5112 3125 5115
rect 3177 5112 3233 5115
rect 3285 5112 5372 5115
rect 5424 5112 5480 5115
rect 5532 5112 5588 5115
rect 5640 5112 5696 5115
rect 5748 5112 5804 5115
rect 5856 5112 5912 5115
rect 5964 5112 6020 5115
rect 6072 5112 6128 5115
rect 6180 5112 6236 5115
rect 6288 5112 6344 5115
rect 6396 5112 7749 5115
rect 7801 5112 7857 5115
rect 7909 5112 7965 5115
rect 8017 5112 8073 5115
rect 8125 5112 8181 5115
rect 8233 5112 8289 5115
rect 8341 5112 8397 5115
rect 8449 5112 8505 5115
rect 8557 5112 8613 5115
rect 8665 5112 8721 5115
rect 8773 5112 8829 5115
rect 8881 5112 8937 5115
rect 8989 5112 9045 5115
rect 9097 5112 9153 5115
rect 9205 5112 9261 5115
rect 9313 5112 9369 5115
rect 9421 5112 9477 5115
rect 9529 5112 11481 5115
rect 1481 5066 1494 5112
rect 11468 5066 11481 5112
rect 1481 5063 1505 5066
rect 1557 5063 1613 5066
rect 1665 5063 1721 5066
rect 1773 5063 1829 5066
rect 1881 5063 1937 5066
rect 1989 5063 2045 5066
rect 2097 5063 2153 5066
rect 2205 5063 2261 5066
rect 2313 5063 2369 5066
rect 2421 5063 2477 5066
rect 2529 5063 2585 5066
rect 2637 5063 2693 5066
rect 2745 5063 2801 5066
rect 2853 5063 2909 5066
rect 2961 5063 3017 5066
rect 3069 5063 3125 5066
rect 3177 5063 3233 5066
rect 3285 5063 5372 5066
rect 5424 5063 5480 5066
rect 5532 5063 5588 5066
rect 5640 5063 5696 5066
rect 5748 5063 5804 5066
rect 5856 5063 5912 5066
rect 5964 5063 6020 5066
rect 6072 5063 6128 5066
rect 6180 5063 6236 5066
rect 6288 5063 6344 5066
rect 6396 5063 7749 5066
rect 7801 5063 7857 5066
rect 7909 5063 7965 5066
rect 8017 5063 8073 5066
rect 8125 5063 8181 5066
rect 8233 5063 8289 5066
rect 8341 5063 8397 5066
rect 8449 5063 8505 5066
rect 8557 5063 8613 5066
rect 8665 5063 8721 5066
rect 8773 5063 8829 5066
rect 8881 5063 8937 5066
rect 8989 5063 9045 5066
rect 9097 5063 9153 5066
rect 9205 5063 9261 5066
rect 9313 5063 9369 5066
rect 9421 5063 9477 5066
rect 9529 5063 11481 5066
rect 1481 5051 11481 5063
rect 1481 4871 11481 4883
rect 1481 4868 3433 4871
rect 3485 4868 3541 4871
rect 3593 4868 3649 4871
rect 3701 4868 3757 4871
rect 3809 4868 3865 4871
rect 3917 4868 3973 4871
rect 4025 4868 4081 4871
rect 4133 4868 4189 4871
rect 4241 4868 4297 4871
rect 4349 4868 4405 4871
rect 4457 4868 4513 4871
rect 4565 4868 4621 4871
rect 4673 4868 4729 4871
rect 4781 4868 4837 4871
rect 4889 4868 4945 4871
rect 4997 4868 5053 4871
rect 5105 4868 5161 4871
rect 5213 4868 6566 4871
rect 6618 4868 6674 4871
rect 6726 4868 6782 4871
rect 6834 4868 6890 4871
rect 6942 4868 6998 4871
rect 7050 4868 7106 4871
rect 7158 4868 7214 4871
rect 7266 4868 7322 4871
rect 7374 4868 7430 4871
rect 7482 4868 7538 4871
rect 7590 4868 9677 4871
rect 9729 4868 9785 4871
rect 9837 4868 9893 4871
rect 9945 4868 10001 4871
rect 10053 4868 10109 4871
rect 10161 4868 10217 4871
rect 10269 4868 10325 4871
rect 10377 4868 10433 4871
rect 10485 4868 10541 4871
rect 10593 4868 10649 4871
rect 10701 4868 10757 4871
rect 10809 4868 10865 4871
rect 10917 4868 10973 4871
rect 11025 4868 11081 4871
rect 11133 4868 11189 4871
rect 11241 4868 11297 4871
rect 11349 4868 11405 4871
rect 11457 4868 11481 4871
rect 1481 4822 1494 4868
rect 11468 4822 11481 4868
rect 1481 4819 3433 4822
rect 3485 4819 3541 4822
rect 3593 4819 3649 4822
rect 3701 4819 3757 4822
rect 3809 4819 3865 4822
rect 3917 4819 3973 4822
rect 4025 4819 4081 4822
rect 4133 4819 4189 4822
rect 4241 4819 4297 4822
rect 4349 4819 4405 4822
rect 4457 4819 4513 4822
rect 4565 4819 4621 4822
rect 4673 4819 4729 4822
rect 4781 4819 4837 4822
rect 4889 4819 4945 4822
rect 4997 4819 5053 4822
rect 5105 4819 5161 4822
rect 5213 4819 6566 4822
rect 6618 4819 6674 4822
rect 6726 4819 6782 4822
rect 6834 4819 6890 4822
rect 6942 4819 6998 4822
rect 7050 4819 7106 4822
rect 7158 4819 7214 4822
rect 7266 4819 7322 4822
rect 7374 4819 7430 4822
rect 7482 4819 7538 4822
rect 7590 4819 9677 4822
rect 9729 4819 9785 4822
rect 9837 4819 9893 4822
rect 9945 4819 10001 4822
rect 10053 4819 10109 4822
rect 10161 4819 10217 4822
rect 10269 4819 10325 4822
rect 10377 4819 10433 4822
rect 10485 4819 10541 4822
rect 10593 4819 10649 4822
rect 10701 4819 10757 4822
rect 10809 4819 10865 4822
rect 10917 4819 10973 4822
rect 11025 4819 11081 4822
rect 11133 4819 11189 4822
rect 11241 4819 11297 4822
rect 11349 4819 11405 4822
rect 11457 4819 11481 4822
rect 1481 4807 11481 4819
rect 1481 4627 11481 4639
rect 1481 4624 1505 4627
rect 1557 4624 1613 4627
rect 1665 4624 1721 4627
rect 1773 4624 1829 4627
rect 1881 4624 1937 4627
rect 1989 4624 2045 4627
rect 2097 4624 2153 4627
rect 2205 4624 2261 4627
rect 2313 4624 2369 4627
rect 2421 4624 2477 4627
rect 2529 4624 2585 4627
rect 2637 4624 2693 4627
rect 2745 4624 2801 4627
rect 2853 4624 2909 4627
rect 2961 4624 3017 4627
rect 3069 4624 3125 4627
rect 3177 4624 3233 4627
rect 3285 4624 5372 4627
rect 5424 4624 5480 4627
rect 5532 4624 5588 4627
rect 5640 4624 5696 4627
rect 5748 4624 5804 4627
rect 5856 4624 5912 4627
rect 5964 4624 6020 4627
rect 6072 4624 6128 4627
rect 6180 4624 6236 4627
rect 6288 4624 6344 4627
rect 6396 4624 7749 4627
rect 7801 4624 7857 4627
rect 7909 4624 7965 4627
rect 8017 4624 8073 4627
rect 8125 4624 8181 4627
rect 8233 4624 8289 4627
rect 8341 4624 8397 4627
rect 8449 4624 8505 4627
rect 8557 4624 8613 4627
rect 8665 4624 8721 4627
rect 8773 4624 8829 4627
rect 8881 4624 8937 4627
rect 8989 4624 9045 4627
rect 9097 4624 9153 4627
rect 9205 4624 9261 4627
rect 9313 4624 9369 4627
rect 9421 4624 9477 4627
rect 9529 4624 11481 4627
rect 1481 4578 1494 4624
rect 11468 4578 11481 4624
rect 1481 4575 1505 4578
rect 1557 4575 1613 4578
rect 1665 4575 1721 4578
rect 1773 4575 1829 4578
rect 1881 4575 1937 4578
rect 1989 4575 2045 4578
rect 2097 4575 2153 4578
rect 2205 4575 2261 4578
rect 2313 4575 2369 4578
rect 2421 4575 2477 4578
rect 2529 4575 2585 4578
rect 2637 4575 2693 4578
rect 2745 4575 2801 4578
rect 2853 4575 2909 4578
rect 2961 4575 3017 4578
rect 3069 4575 3125 4578
rect 3177 4575 3233 4578
rect 3285 4575 5372 4578
rect 5424 4575 5480 4578
rect 5532 4575 5588 4578
rect 5640 4575 5696 4578
rect 5748 4575 5804 4578
rect 5856 4575 5912 4578
rect 5964 4575 6020 4578
rect 6072 4575 6128 4578
rect 6180 4575 6236 4578
rect 6288 4575 6344 4578
rect 6396 4575 7749 4578
rect 7801 4575 7857 4578
rect 7909 4575 7965 4578
rect 8017 4575 8073 4578
rect 8125 4575 8181 4578
rect 8233 4575 8289 4578
rect 8341 4575 8397 4578
rect 8449 4575 8505 4578
rect 8557 4575 8613 4578
rect 8665 4575 8721 4578
rect 8773 4575 8829 4578
rect 8881 4575 8937 4578
rect 8989 4575 9045 4578
rect 9097 4575 9153 4578
rect 9205 4575 9261 4578
rect 9313 4575 9369 4578
rect 9421 4575 9477 4578
rect 9529 4575 11481 4578
rect 1481 4563 11481 4575
rect 1481 4383 11481 4395
rect 1481 4380 3433 4383
rect 3485 4380 3541 4383
rect 3593 4380 3649 4383
rect 3701 4380 3757 4383
rect 3809 4380 3865 4383
rect 3917 4380 3973 4383
rect 4025 4380 4081 4383
rect 4133 4380 4189 4383
rect 4241 4380 4297 4383
rect 4349 4380 4405 4383
rect 4457 4380 4513 4383
rect 4565 4380 4621 4383
rect 4673 4380 4729 4383
rect 4781 4380 4837 4383
rect 4889 4380 4945 4383
rect 4997 4380 5053 4383
rect 5105 4380 5161 4383
rect 5213 4380 6566 4383
rect 6618 4380 6674 4383
rect 6726 4380 6782 4383
rect 6834 4380 6890 4383
rect 6942 4380 6998 4383
rect 7050 4380 7106 4383
rect 7158 4380 7214 4383
rect 7266 4380 7322 4383
rect 7374 4380 7430 4383
rect 7482 4380 7538 4383
rect 7590 4380 9677 4383
rect 9729 4380 9785 4383
rect 9837 4380 9893 4383
rect 9945 4380 10001 4383
rect 10053 4380 10109 4383
rect 10161 4380 10217 4383
rect 10269 4380 10325 4383
rect 10377 4380 10433 4383
rect 10485 4380 10541 4383
rect 10593 4380 10649 4383
rect 10701 4380 10757 4383
rect 10809 4380 10865 4383
rect 10917 4380 10973 4383
rect 11025 4380 11081 4383
rect 11133 4380 11189 4383
rect 11241 4380 11297 4383
rect 11349 4380 11405 4383
rect 11457 4380 11481 4383
rect 1481 4334 1494 4380
rect 11468 4334 11481 4380
rect 1481 4331 3433 4334
rect 3485 4331 3541 4334
rect 3593 4331 3649 4334
rect 3701 4331 3757 4334
rect 3809 4331 3865 4334
rect 3917 4331 3973 4334
rect 4025 4331 4081 4334
rect 4133 4331 4189 4334
rect 4241 4331 4297 4334
rect 4349 4331 4405 4334
rect 4457 4331 4513 4334
rect 4565 4331 4621 4334
rect 4673 4331 4729 4334
rect 4781 4331 4837 4334
rect 4889 4331 4945 4334
rect 4997 4331 5053 4334
rect 5105 4331 5161 4334
rect 5213 4331 6566 4334
rect 6618 4331 6674 4334
rect 6726 4331 6782 4334
rect 6834 4331 6890 4334
rect 6942 4331 6998 4334
rect 7050 4331 7106 4334
rect 7158 4331 7214 4334
rect 7266 4331 7322 4334
rect 7374 4331 7430 4334
rect 7482 4331 7538 4334
rect 7590 4331 9677 4334
rect 9729 4331 9785 4334
rect 9837 4331 9893 4334
rect 9945 4331 10001 4334
rect 10053 4331 10109 4334
rect 10161 4331 10217 4334
rect 10269 4331 10325 4334
rect 10377 4331 10433 4334
rect 10485 4331 10541 4334
rect 10593 4331 10649 4334
rect 10701 4331 10757 4334
rect 10809 4331 10865 4334
rect 10917 4331 10973 4334
rect 11025 4331 11081 4334
rect 11133 4331 11189 4334
rect 11241 4331 11297 4334
rect 11349 4331 11405 4334
rect 11457 4331 11481 4334
rect 1481 4319 11481 4331
rect 1481 4139 11481 4151
rect 1481 4136 1505 4139
rect 1557 4136 1613 4139
rect 1665 4136 1721 4139
rect 1773 4136 1829 4139
rect 1881 4136 1937 4139
rect 1989 4136 2045 4139
rect 2097 4136 2153 4139
rect 2205 4136 2261 4139
rect 2313 4136 2369 4139
rect 2421 4136 2477 4139
rect 2529 4136 2585 4139
rect 2637 4136 2693 4139
rect 2745 4136 2801 4139
rect 2853 4136 2909 4139
rect 2961 4136 3017 4139
rect 3069 4136 3125 4139
rect 3177 4136 3233 4139
rect 3285 4136 5372 4139
rect 5424 4136 5480 4139
rect 5532 4136 5588 4139
rect 5640 4136 5696 4139
rect 5748 4136 5804 4139
rect 5856 4136 5912 4139
rect 5964 4136 6020 4139
rect 6072 4136 6128 4139
rect 6180 4136 6236 4139
rect 6288 4136 6344 4139
rect 6396 4136 7749 4139
rect 7801 4136 7857 4139
rect 7909 4136 7965 4139
rect 8017 4136 8073 4139
rect 8125 4136 8181 4139
rect 8233 4136 8289 4139
rect 8341 4136 8397 4139
rect 8449 4136 8505 4139
rect 8557 4136 8613 4139
rect 8665 4136 8721 4139
rect 8773 4136 8829 4139
rect 8881 4136 8937 4139
rect 8989 4136 9045 4139
rect 9097 4136 9153 4139
rect 9205 4136 9261 4139
rect 9313 4136 9369 4139
rect 9421 4136 9477 4139
rect 9529 4136 11481 4139
rect 1481 4090 1494 4136
rect 11468 4090 11481 4136
rect 1481 4087 1505 4090
rect 1557 4087 1613 4090
rect 1665 4087 1721 4090
rect 1773 4087 1829 4090
rect 1881 4087 1937 4090
rect 1989 4087 2045 4090
rect 2097 4087 2153 4090
rect 2205 4087 2261 4090
rect 2313 4087 2369 4090
rect 2421 4087 2477 4090
rect 2529 4087 2585 4090
rect 2637 4087 2693 4090
rect 2745 4087 2801 4090
rect 2853 4087 2909 4090
rect 2961 4087 3017 4090
rect 3069 4087 3125 4090
rect 3177 4087 3233 4090
rect 3285 4087 5372 4090
rect 5424 4087 5480 4090
rect 5532 4087 5588 4090
rect 5640 4087 5696 4090
rect 5748 4087 5804 4090
rect 5856 4087 5912 4090
rect 5964 4087 6020 4090
rect 6072 4087 6128 4090
rect 6180 4087 6236 4090
rect 6288 4087 6344 4090
rect 6396 4087 7749 4090
rect 7801 4087 7857 4090
rect 7909 4087 7965 4090
rect 8017 4087 8073 4090
rect 8125 4087 8181 4090
rect 8233 4087 8289 4090
rect 8341 4087 8397 4090
rect 8449 4087 8505 4090
rect 8557 4087 8613 4090
rect 8665 4087 8721 4090
rect 8773 4087 8829 4090
rect 8881 4087 8937 4090
rect 8989 4087 9045 4090
rect 9097 4087 9153 4090
rect 9205 4087 9261 4090
rect 9313 4087 9369 4090
rect 9421 4087 9477 4090
rect 9529 4087 11481 4090
rect 1481 4075 11481 4087
rect 1481 3895 11481 3907
rect 1481 3892 3433 3895
rect 3485 3892 3541 3895
rect 3593 3892 3649 3895
rect 3701 3892 3757 3895
rect 3809 3892 3865 3895
rect 3917 3892 3973 3895
rect 4025 3892 4081 3895
rect 4133 3892 4189 3895
rect 4241 3892 4297 3895
rect 4349 3892 4405 3895
rect 4457 3892 4513 3895
rect 4565 3892 4621 3895
rect 4673 3892 4729 3895
rect 4781 3892 4837 3895
rect 4889 3892 4945 3895
rect 4997 3892 5053 3895
rect 5105 3892 5161 3895
rect 5213 3892 6566 3895
rect 6618 3892 6674 3895
rect 6726 3892 6782 3895
rect 6834 3892 6890 3895
rect 6942 3892 6998 3895
rect 7050 3892 7106 3895
rect 7158 3892 7214 3895
rect 7266 3892 7322 3895
rect 7374 3892 7430 3895
rect 7482 3892 7538 3895
rect 7590 3892 9677 3895
rect 9729 3892 9785 3895
rect 9837 3892 9893 3895
rect 9945 3892 10001 3895
rect 10053 3892 10109 3895
rect 10161 3892 10217 3895
rect 10269 3892 10325 3895
rect 10377 3892 10433 3895
rect 10485 3892 10541 3895
rect 10593 3892 10649 3895
rect 10701 3892 10757 3895
rect 10809 3892 10865 3895
rect 10917 3892 10973 3895
rect 11025 3892 11081 3895
rect 11133 3892 11189 3895
rect 11241 3892 11297 3895
rect 11349 3892 11405 3895
rect 11457 3892 11481 3895
rect 1481 3846 1494 3892
rect 11468 3846 11481 3892
rect 1481 3843 3433 3846
rect 3485 3843 3541 3846
rect 3593 3843 3649 3846
rect 3701 3843 3757 3846
rect 3809 3843 3865 3846
rect 3917 3843 3973 3846
rect 4025 3843 4081 3846
rect 4133 3843 4189 3846
rect 4241 3843 4297 3846
rect 4349 3843 4405 3846
rect 4457 3843 4513 3846
rect 4565 3843 4621 3846
rect 4673 3843 4729 3846
rect 4781 3843 4837 3846
rect 4889 3843 4945 3846
rect 4997 3843 5053 3846
rect 5105 3843 5161 3846
rect 5213 3843 6566 3846
rect 6618 3843 6674 3846
rect 6726 3843 6782 3846
rect 6834 3843 6890 3846
rect 6942 3843 6998 3846
rect 7050 3843 7106 3846
rect 7158 3843 7214 3846
rect 7266 3843 7322 3846
rect 7374 3843 7430 3846
rect 7482 3843 7538 3846
rect 7590 3843 9677 3846
rect 9729 3843 9785 3846
rect 9837 3843 9893 3846
rect 9945 3843 10001 3846
rect 10053 3843 10109 3846
rect 10161 3843 10217 3846
rect 10269 3843 10325 3846
rect 10377 3843 10433 3846
rect 10485 3843 10541 3846
rect 10593 3843 10649 3846
rect 10701 3843 10757 3846
rect 10809 3843 10865 3846
rect 10917 3843 10973 3846
rect 11025 3843 11081 3846
rect 11133 3843 11189 3846
rect 11241 3843 11297 3846
rect 11349 3843 11405 3846
rect 11457 3843 11481 3846
rect 1481 3831 11481 3843
rect 1481 3651 11481 3663
rect 1481 3648 1505 3651
rect 1557 3648 1613 3651
rect 1665 3648 1721 3651
rect 1773 3648 1829 3651
rect 1881 3648 1937 3651
rect 1989 3648 2045 3651
rect 2097 3648 2153 3651
rect 2205 3648 2261 3651
rect 2313 3648 2369 3651
rect 2421 3648 2477 3651
rect 2529 3648 2585 3651
rect 2637 3648 2693 3651
rect 2745 3648 2801 3651
rect 2853 3648 2909 3651
rect 2961 3648 3017 3651
rect 3069 3648 3125 3651
rect 3177 3648 3233 3651
rect 3285 3648 5372 3651
rect 5424 3648 5480 3651
rect 5532 3648 5588 3651
rect 5640 3648 5696 3651
rect 5748 3648 5804 3651
rect 5856 3648 5912 3651
rect 5964 3648 6020 3651
rect 6072 3648 6128 3651
rect 6180 3648 6236 3651
rect 6288 3648 6344 3651
rect 6396 3648 7749 3651
rect 7801 3648 7857 3651
rect 7909 3648 7965 3651
rect 8017 3648 8073 3651
rect 8125 3648 8181 3651
rect 8233 3648 8289 3651
rect 8341 3648 8397 3651
rect 8449 3648 8505 3651
rect 8557 3648 8613 3651
rect 8665 3648 8721 3651
rect 8773 3648 8829 3651
rect 8881 3648 8937 3651
rect 8989 3648 9045 3651
rect 9097 3648 9153 3651
rect 9205 3648 9261 3651
rect 9313 3648 9369 3651
rect 9421 3648 9477 3651
rect 9529 3648 11481 3651
rect 1481 3602 1494 3648
rect 11468 3602 11481 3648
rect 1481 3599 1505 3602
rect 1557 3599 1613 3602
rect 1665 3599 1721 3602
rect 1773 3599 1829 3602
rect 1881 3599 1937 3602
rect 1989 3599 2045 3602
rect 2097 3599 2153 3602
rect 2205 3599 2261 3602
rect 2313 3599 2369 3602
rect 2421 3599 2477 3602
rect 2529 3599 2585 3602
rect 2637 3599 2693 3602
rect 2745 3599 2801 3602
rect 2853 3599 2909 3602
rect 2961 3599 3017 3602
rect 3069 3599 3125 3602
rect 3177 3599 3233 3602
rect 3285 3599 5372 3602
rect 5424 3599 5480 3602
rect 5532 3599 5588 3602
rect 5640 3599 5696 3602
rect 5748 3599 5804 3602
rect 5856 3599 5912 3602
rect 5964 3599 6020 3602
rect 6072 3599 6128 3602
rect 6180 3599 6236 3602
rect 6288 3599 6344 3602
rect 6396 3599 7749 3602
rect 7801 3599 7857 3602
rect 7909 3599 7965 3602
rect 8017 3599 8073 3602
rect 8125 3599 8181 3602
rect 8233 3599 8289 3602
rect 8341 3599 8397 3602
rect 8449 3599 8505 3602
rect 8557 3599 8613 3602
rect 8665 3599 8721 3602
rect 8773 3599 8829 3602
rect 8881 3599 8937 3602
rect 8989 3599 9045 3602
rect 9097 3599 9153 3602
rect 9205 3599 9261 3602
rect 9313 3599 9369 3602
rect 9421 3599 9477 3602
rect 9529 3599 11481 3602
rect 1481 3587 11481 3599
rect 1481 3407 11481 3419
rect 1481 3404 3433 3407
rect 3485 3404 3541 3407
rect 3593 3404 3649 3407
rect 3701 3404 3757 3407
rect 3809 3404 3865 3407
rect 3917 3404 3973 3407
rect 4025 3404 4081 3407
rect 4133 3404 4189 3407
rect 4241 3404 4297 3407
rect 4349 3404 4405 3407
rect 4457 3404 4513 3407
rect 4565 3404 4621 3407
rect 4673 3404 4729 3407
rect 4781 3404 4837 3407
rect 4889 3404 4945 3407
rect 4997 3404 5053 3407
rect 5105 3404 5161 3407
rect 5213 3404 6566 3407
rect 6618 3404 6674 3407
rect 6726 3404 6782 3407
rect 6834 3404 6890 3407
rect 6942 3404 6998 3407
rect 7050 3404 7106 3407
rect 7158 3404 7214 3407
rect 7266 3404 7322 3407
rect 7374 3404 7430 3407
rect 7482 3404 7538 3407
rect 7590 3404 9677 3407
rect 9729 3404 9785 3407
rect 9837 3404 9893 3407
rect 9945 3404 10001 3407
rect 10053 3404 10109 3407
rect 10161 3404 10217 3407
rect 10269 3404 10325 3407
rect 10377 3404 10433 3407
rect 10485 3404 10541 3407
rect 10593 3404 10649 3407
rect 10701 3404 10757 3407
rect 10809 3404 10865 3407
rect 10917 3404 10973 3407
rect 11025 3404 11081 3407
rect 11133 3404 11189 3407
rect 11241 3404 11297 3407
rect 11349 3404 11405 3407
rect 11457 3404 11481 3407
rect 1481 3358 1494 3404
rect 11468 3358 11481 3404
rect 1481 3355 3433 3358
rect 3485 3355 3541 3358
rect 3593 3355 3649 3358
rect 3701 3355 3757 3358
rect 3809 3355 3865 3358
rect 3917 3355 3973 3358
rect 4025 3355 4081 3358
rect 4133 3355 4189 3358
rect 4241 3355 4297 3358
rect 4349 3355 4405 3358
rect 4457 3355 4513 3358
rect 4565 3355 4621 3358
rect 4673 3355 4729 3358
rect 4781 3355 4837 3358
rect 4889 3355 4945 3358
rect 4997 3355 5053 3358
rect 5105 3355 5161 3358
rect 5213 3355 6566 3358
rect 6618 3355 6674 3358
rect 6726 3355 6782 3358
rect 6834 3355 6890 3358
rect 6942 3355 6998 3358
rect 7050 3355 7106 3358
rect 7158 3355 7214 3358
rect 7266 3355 7322 3358
rect 7374 3355 7430 3358
rect 7482 3355 7538 3358
rect 7590 3355 9677 3358
rect 9729 3355 9785 3358
rect 9837 3355 9893 3358
rect 9945 3355 10001 3358
rect 10053 3355 10109 3358
rect 10161 3355 10217 3358
rect 10269 3355 10325 3358
rect 10377 3355 10433 3358
rect 10485 3355 10541 3358
rect 10593 3355 10649 3358
rect 10701 3355 10757 3358
rect 10809 3355 10865 3358
rect 10917 3355 10973 3358
rect 11025 3355 11081 3358
rect 11133 3355 11189 3358
rect 11241 3355 11297 3358
rect 11349 3355 11405 3358
rect 11457 3355 11481 3358
rect 1481 3343 11481 3355
rect 1481 3163 11481 3175
rect 1481 3160 1505 3163
rect 1557 3160 1613 3163
rect 1665 3160 1721 3163
rect 1773 3160 1829 3163
rect 1881 3160 1937 3163
rect 1989 3160 2045 3163
rect 2097 3160 2153 3163
rect 2205 3160 2261 3163
rect 2313 3160 2369 3163
rect 2421 3160 2477 3163
rect 2529 3160 2585 3163
rect 2637 3160 2693 3163
rect 2745 3160 2801 3163
rect 2853 3160 2909 3163
rect 2961 3160 3017 3163
rect 3069 3160 3125 3163
rect 3177 3160 3233 3163
rect 3285 3160 5372 3163
rect 5424 3160 5480 3163
rect 5532 3160 5588 3163
rect 5640 3160 5696 3163
rect 5748 3160 5804 3163
rect 5856 3160 5912 3163
rect 5964 3160 6020 3163
rect 6072 3160 6128 3163
rect 6180 3160 6236 3163
rect 6288 3160 6344 3163
rect 6396 3160 7749 3163
rect 7801 3160 7857 3163
rect 7909 3160 7965 3163
rect 8017 3160 8073 3163
rect 8125 3160 8181 3163
rect 8233 3160 8289 3163
rect 8341 3160 8397 3163
rect 8449 3160 8505 3163
rect 8557 3160 8613 3163
rect 8665 3160 8721 3163
rect 8773 3160 8829 3163
rect 8881 3160 8937 3163
rect 8989 3160 9045 3163
rect 9097 3160 9153 3163
rect 9205 3160 9261 3163
rect 9313 3160 9369 3163
rect 9421 3160 9477 3163
rect 9529 3160 11481 3163
rect 1481 3114 1494 3160
rect 11468 3114 11481 3160
rect 1481 3111 1505 3114
rect 1557 3111 1613 3114
rect 1665 3111 1721 3114
rect 1773 3111 1829 3114
rect 1881 3111 1937 3114
rect 1989 3111 2045 3114
rect 2097 3111 2153 3114
rect 2205 3111 2261 3114
rect 2313 3111 2369 3114
rect 2421 3111 2477 3114
rect 2529 3111 2585 3114
rect 2637 3111 2693 3114
rect 2745 3111 2801 3114
rect 2853 3111 2909 3114
rect 2961 3111 3017 3114
rect 3069 3111 3125 3114
rect 3177 3111 3233 3114
rect 3285 3111 5372 3114
rect 5424 3111 5480 3114
rect 5532 3111 5588 3114
rect 5640 3111 5696 3114
rect 5748 3111 5804 3114
rect 5856 3111 5912 3114
rect 5964 3111 6020 3114
rect 6072 3111 6128 3114
rect 6180 3111 6236 3114
rect 6288 3111 6344 3114
rect 6396 3111 7749 3114
rect 7801 3111 7857 3114
rect 7909 3111 7965 3114
rect 8017 3111 8073 3114
rect 8125 3111 8181 3114
rect 8233 3111 8289 3114
rect 8341 3111 8397 3114
rect 8449 3111 8505 3114
rect 8557 3111 8613 3114
rect 8665 3111 8721 3114
rect 8773 3111 8829 3114
rect 8881 3111 8937 3114
rect 8989 3111 9045 3114
rect 9097 3111 9153 3114
rect 9205 3111 9261 3114
rect 9313 3111 9369 3114
rect 9421 3111 9477 3114
rect 9529 3111 11481 3114
rect 1481 3099 11481 3111
rect 1481 2919 11481 2931
rect 1481 2916 3433 2919
rect 3485 2916 3541 2919
rect 3593 2916 3649 2919
rect 3701 2916 3757 2919
rect 3809 2916 3865 2919
rect 3917 2916 3973 2919
rect 4025 2916 4081 2919
rect 4133 2916 4189 2919
rect 4241 2916 4297 2919
rect 4349 2916 4405 2919
rect 4457 2916 4513 2919
rect 4565 2916 4621 2919
rect 4673 2916 4729 2919
rect 4781 2916 4837 2919
rect 4889 2916 4945 2919
rect 4997 2916 5053 2919
rect 5105 2916 5161 2919
rect 5213 2916 6566 2919
rect 6618 2916 6674 2919
rect 6726 2916 6782 2919
rect 6834 2916 6890 2919
rect 6942 2916 6998 2919
rect 7050 2916 7106 2919
rect 7158 2916 7214 2919
rect 7266 2916 7322 2919
rect 7374 2916 7430 2919
rect 7482 2916 7538 2919
rect 7590 2916 9677 2919
rect 9729 2916 9785 2919
rect 9837 2916 9893 2919
rect 9945 2916 10001 2919
rect 10053 2916 10109 2919
rect 10161 2916 10217 2919
rect 10269 2916 10325 2919
rect 10377 2916 10433 2919
rect 10485 2916 10541 2919
rect 10593 2916 10649 2919
rect 10701 2916 10757 2919
rect 10809 2916 10865 2919
rect 10917 2916 10973 2919
rect 11025 2916 11081 2919
rect 11133 2916 11189 2919
rect 11241 2916 11297 2919
rect 11349 2916 11405 2919
rect 11457 2916 11481 2919
rect 1481 2870 1494 2916
rect 11468 2870 11481 2916
rect 1481 2867 3433 2870
rect 3485 2867 3541 2870
rect 3593 2867 3649 2870
rect 3701 2867 3757 2870
rect 3809 2867 3865 2870
rect 3917 2867 3973 2870
rect 4025 2867 4081 2870
rect 4133 2867 4189 2870
rect 4241 2867 4297 2870
rect 4349 2867 4405 2870
rect 4457 2867 4513 2870
rect 4565 2867 4621 2870
rect 4673 2867 4729 2870
rect 4781 2867 4837 2870
rect 4889 2867 4945 2870
rect 4997 2867 5053 2870
rect 5105 2867 5161 2870
rect 5213 2867 6566 2870
rect 6618 2867 6674 2870
rect 6726 2867 6782 2870
rect 6834 2867 6890 2870
rect 6942 2867 6998 2870
rect 7050 2867 7106 2870
rect 7158 2867 7214 2870
rect 7266 2867 7322 2870
rect 7374 2867 7430 2870
rect 7482 2867 7538 2870
rect 7590 2867 9677 2870
rect 9729 2867 9785 2870
rect 9837 2867 9893 2870
rect 9945 2867 10001 2870
rect 10053 2867 10109 2870
rect 10161 2867 10217 2870
rect 10269 2867 10325 2870
rect 10377 2867 10433 2870
rect 10485 2867 10541 2870
rect 10593 2867 10649 2870
rect 10701 2867 10757 2870
rect 10809 2867 10865 2870
rect 10917 2867 10973 2870
rect 11025 2867 11081 2870
rect 11133 2867 11189 2870
rect 11241 2867 11297 2870
rect 11349 2867 11405 2870
rect 11457 2867 11481 2870
rect 1481 2855 11481 2867
rect 1481 2675 11481 2687
rect 1481 2672 1505 2675
rect 1557 2672 1613 2675
rect 1665 2672 1721 2675
rect 1773 2672 1829 2675
rect 1881 2672 1937 2675
rect 1989 2672 2045 2675
rect 2097 2672 2153 2675
rect 2205 2672 2261 2675
rect 2313 2672 2369 2675
rect 2421 2672 2477 2675
rect 2529 2672 2585 2675
rect 2637 2672 2693 2675
rect 2745 2672 2801 2675
rect 2853 2672 2909 2675
rect 2961 2672 3017 2675
rect 3069 2672 3125 2675
rect 3177 2672 3233 2675
rect 3285 2672 5372 2675
rect 5424 2672 5480 2675
rect 5532 2672 5588 2675
rect 5640 2672 5696 2675
rect 5748 2672 5804 2675
rect 5856 2672 5912 2675
rect 5964 2672 6020 2675
rect 6072 2672 6128 2675
rect 6180 2672 6236 2675
rect 6288 2672 6344 2675
rect 6396 2672 7749 2675
rect 7801 2672 7857 2675
rect 7909 2672 7965 2675
rect 8017 2672 8073 2675
rect 8125 2672 8181 2675
rect 8233 2672 8289 2675
rect 8341 2672 8397 2675
rect 8449 2672 8505 2675
rect 8557 2672 8613 2675
rect 8665 2672 8721 2675
rect 8773 2672 8829 2675
rect 8881 2672 8937 2675
rect 8989 2672 9045 2675
rect 9097 2672 9153 2675
rect 9205 2672 9261 2675
rect 9313 2672 9369 2675
rect 9421 2672 9477 2675
rect 9529 2672 11481 2675
rect 1481 2626 1494 2672
rect 11468 2626 11481 2672
rect 1481 2623 1505 2626
rect 1557 2623 1613 2626
rect 1665 2623 1721 2626
rect 1773 2623 1829 2626
rect 1881 2623 1937 2626
rect 1989 2623 2045 2626
rect 2097 2623 2153 2626
rect 2205 2623 2261 2626
rect 2313 2623 2369 2626
rect 2421 2623 2477 2626
rect 2529 2623 2585 2626
rect 2637 2623 2693 2626
rect 2745 2623 2801 2626
rect 2853 2623 2909 2626
rect 2961 2623 3017 2626
rect 3069 2623 3125 2626
rect 3177 2623 3233 2626
rect 3285 2623 5372 2626
rect 5424 2623 5480 2626
rect 5532 2623 5588 2626
rect 5640 2623 5696 2626
rect 5748 2623 5804 2626
rect 5856 2623 5912 2626
rect 5964 2623 6020 2626
rect 6072 2623 6128 2626
rect 6180 2623 6236 2626
rect 6288 2623 6344 2626
rect 6396 2623 7749 2626
rect 7801 2623 7857 2626
rect 7909 2623 7965 2626
rect 8017 2623 8073 2626
rect 8125 2623 8181 2626
rect 8233 2623 8289 2626
rect 8341 2623 8397 2626
rect 8449 2623 8505 2626
rect 8557 2623 8613 2626
rect 8665 2623 8721 2626
rect 8773 2623 8829 2626
rect 8881 2623 8937 2626
rect 8989 2623 9045 2626
rect 9097 2623 9153 2626
rect 9205 2623 9261 2626
rect 9313 2623 9369 2626
rect 9421 2623 9477 2626
rect 9529 2623 11481 2626
rect 1481 2611 11481 2623
rect 1481 2431 11481 2443
rect 1481 2428 3433 2431
rect 3485 2428 3541 2431
rect 3593 2428 3649 2431
rect 3701 2428 3757 2431
rect 3809 2428 3865 2431
rect 3917 2428 3973 2431
rect 4025 2428 4081 2431
rect 4133 2428 4189 2431
rect 4241 2428 4297 2431
rect 4349 2428 4405 2431
rect 4457 2428 4513 2431
rect 4565 2428 4621 2431
rect 4673 2428 4729 2431
rect 4781 2428 4837 2431
rect 4889 2428 4945 2431
rect 4997 2428 5053 2431
rect 5105 2428 5161 2431
rect 5213 2428 6566 2431
rect 6618 2428 6674 2431
rect 6726 2428 6782 2431
rect 6834 2428 6890 2431
rect 6942 2428 6998 2431
rect 7050 2428 7106 2431
rect 7158 2428 7214 2431
rect 7266 2428 7322 2431
rect 7374 2428 7430 2431
rect 7482 2428 7538 2431
rect 7590 2428 9677 2431
rect 9729 2428 9785 2431
rect 9837 2428 9893 2431
rect 9945 2428 10001 2431
rect 10053 2428 10109 2431
rect 10161 2428 10217 2431
rect 10269 2428 10325 2431
rect 10377 2428 10433 2431
rect 10485 2428 10541 2431
rect 10593 2428 10649 2431
rect 10701 2428 10757 2431
rect 10809 2428 10865 2431
rect 10917 2428 10973 2431
rect 11025 2428 11081 2431
rect 11133 2428 11189 2431
rect 11241 2428 11297 2431
rect 11349 2428 11405 2431
rect 11457 2428 11481 2431
rect 1481 2382 1494 2428
rect 11468 2382 11481 2428
rect 1481 2379 3433 2382
rect 3485 2379 3541 2382
rect 3593 2379 3649 2382
rect 3701 2379 3757 2382
rect 3809 2379 3865 2382
rect 3917 2379 3973 2382
rect 4025 2379 4081 2382
rect 4133 2379 4189 2382
rect 4241 2379 4297 2382
rect 4349 2379 4405 2382
rect 4457 2379 4513 2382
rect 4565 2379 4621 2382
rect 4673 2379 4729 2382
rect 4781 2379 4837 2382
rect 4889 2379 4945 2382
rect 4997 2379 5053 2382
rect 5105 2379 5161 2382
rect 5213 2379 6566 2382
rect 6618 2379 6674 2382
rect 6726 2379 6782 2382
rect 6834 2379 6890 2382
rect 6942 2379 6998 2382
rect 7050 2379 7106 2382
rect 7158 2379 7214 2382
rect 7266 2379 7322 2382
rect 7374 2379 7430 2382
rect 7482 2379 7538 2382
rect 7590 2379 9677 2382
rect 9729 2379 9785 2382
rect 9837 2379 9893 2382
rect 9945 2379 10001 2382
rect 10053 2379 10109 2382
rect 10161 2379 10217 2382
rect 10269 2379 10325 2382
rect 10377 2379 10433 2382
rect 10485 2379 10541 2382
rect 10593 2379 10649 2382
rect 10701 2379 10757 2382
rect 10809 2379 10865 2382
rect 10917 2379 10973 2382
rect 11025 2379 11081 2382
rect 11133 2379 11189 2382
rect 11241 2379 11297 2382
rect 11349 2379 11405 2382
rect 11457 2379 11481 2382
rect 1481 2367 11481 2379
rect 1481 2187 11481 2199
rect 1481 2184 1505 2187
rect 1557 2184 1613 2187
rect 1665 2184 1721 2187
rect 1773 2184 1829 2187
rect 1881 2184 1937 2187
rect 1989 2184 2045 2187
rect 2097 2184 2153 2187
rect 2205 2184 2261 2187
rect 2313 2184 2369 2187
rect 2421 2184 2477 2187
rect 2529 2184 2585 2187
rect 2637 2184 2693 2187
rect 2745 2184 2801 2187
rect 2853 2184 2909 2187
rect 2961 2184 3017 2187
rect 3069 2184 3125 2187
rect 3177 2184 3233 2187
rect 3285 2184 5372 2187
rect 5424 2184 5480 2187
rect 5532 2184 5588 2187
rect 5640 2184 5696 2187
rect 5748 2184 5804 2187
rect 5856 2184 5912 2187
rect 5964 2184 6020 2187
rect 6072 2184 6128 2187
rect 6180 2184 6236 2187
rect 6288 2184 6344 2187
rect 6396 2184 7749 2187
rect 7801 2184 7857 2187
rect 7909 2184 7965 2187
rect 8017 2184 8073 2187
rect 8125 2184 8181 2187
rect 8233 2184 8289 2187
rect 8341 2184 8397 2187
rect 8449 2184 8505 2187
rect 8557 2184 8613 2187
rect 8665 2184 8721 2187
rect 8773 2184 8829 2187
rect 8881 2184 8937 2187
rect 8989 2184 9045 2187
rect 9097 2184 9153 2187
rect 9205 2184 9261 2187
rect 9313 2184 9369 2187
rect 9421 2184 9477 2187
rect 9529 2184 11481 2187
rect 1481 2138 1494 2184
rect 11468 2138 11481 2184
rect 1481 2135 1505 2138
rect 1557 2135 1613 2138
rect 1665 2135 1721 2138
rect 1773 2135 1829 2138
rect 1881 2135 1937 2138
rect 1989 2135 2045 2138
rect 2097 2135 2153 2138
rect 2205 2135 2261 2138
rect 2313 2135 2369 2138
rect 2421 2135 2477 2138
rect 2529 2135 2585 2138
rect 2637 2135 2693 2138
rect 2745 2135 2801 2138
rect 2853 2135 2909 2138
rect 2961 2135 3017 2138
rect 3069 2135 3125 2138
rect 3177 2135 3233 2138
rect 3285 2135 5372 2138
rect 5424 2135 5480 2138
rect 5532 2135 5588 2138
rect 5640 2135 5696 2138
rect 5748 2135 5804 2138
rect 5856 2135 5912 2138
rect 5964 2135 6020 2138
rect 6072 2135 6128 2138
rect 6180 2135 6236 2138
rect 6288 2135 6344 2138
rect 6396 2135 7749 2138
rect 7801 2135 7857 2138
rect 7909 2135 7965 2138
rect 8017 2135 8073 2138
rect 8125 2135 8181 2138
rect 8233 2135 8289 2138
rect 8341 2135 8397 2138
rect 8449 2135 8505 2138
rect 8557 2135 8613 2138
rect 8665 2135 8721 2138
rect 8773 2135 8829 2138
rect 8881 2135 8937 2138
rect 8989 2135 9045 2138
rect 9097 2135 9153 2138
rect 9205 2135 9261 2138
rect 9313 2135 9369 2138
rect 9421 2135 9477 2138
rect 9529 2135 11481 2138
rect 1481 2123 11481 2135
rect 1481 1943 11481 1955
rect 1481 1940 3433 1943
rect 3485 1940 3541 1943
rect 3593 1940 3649 1943
rect 3701 1940 3757 1943
rect 3809 1940 3865 1943
rect 3917 1940 3973 1943
rect 4025 1940 4081 1943
rect 4133 1940 4189 1943
rect 4241 1940 4297 1943
rect 4349 1940 4405 1943
rect 4457 1940 4513 1943
rect 4565 1940 4621 1943
rect 4673 1940 4729 1943
rect 4781 1940 4837 1943
rect 4889 1940 4945 1943
rect 4997 1940 5053 1943
rect 5105 1940 5161 1943
rect 5213 1940 6566 1943
rect 6618 1940 6674 1943
rect 6726 1940 6782 1943
rect 6834 1940 6890 1943
rect 6942 1940 6998 1943
rect 7050 1940 7106 1943
rect 7158 1940 7214 1943
rect 7266 1940 7322 1943
rect 7374 1940 7430 1943
rect 7482 1940 7538 1943
rect 7590 1940 9677 1943
rect 9729 1940 9785 1943
rect 9837 1940 9893 1943
rect 9945 1940 10001 1943
rect 10053 1940 10109 1943
rect 10161 1940 10217 1943
rect 10269 1940 10325 1943
rect 10377 1940 10433 1943
rect 10485 1940 10541 1943
rect 10593 1940 10649 1943
rect 10701 1940 10757 1943
rect 10809 1940 10865 1943
rect 10917 1940 10973 1943
rect 11025 1940 11081 1943
rect 11133 1940 11189 1943
rect 11241 1940 11297 1943
rect 11349 1940 11405 1943
rect 11457 1940 11481 1943
rect 1481 1894 1494 1940
rect 11468 1894 11481 1940
rect 1481 1891 3433 1894
rect 3485 1891 3541 1894
rect 3593 1891 3649 1894
rect 3701 1891 3757 1894
rect 3809 1891 3865 1894
rect 3917 1891 3973 1894
rect 4025 1891 4081 1894
rect 4133 1891 4189 1894
rect 4241 1891 4297 1894
rect 4349 1891 4405 1894
rect 4457 1891 4513 1894
rect 4565 1891 4621 1894
rect 4673 1891 4729 1894
rect 4781 1891 4837 1894
rect 4889 1891 4945 1894
rect 4997 1891 5053 1894
rect 5105 1891 5161 1894
rect 5213 1891 6566 1894
rect 6618 1891 6674 1894
rect 6726 1891 6782 1894
rect 6834 1891 6890 1894
rect 6942 1891 6998 1894
rect 7050 1891 7106 1894
rect 7158 1891 7214 1894
rect 7266 1891 7322 1894
rect 7374 1891 7430 1894
rect 7482 1891 7538 1894
rect 7590 1891 9677 1894
rect 9729 1891 9785 1894
rect 9837 1891 9893 1894
rect 9945 1891 10001 1894
rect 10053 1891 10109 1894
rect 10161 1891 10217 1894
rect 10269 1891 10325 1894
rect 10377 1891 10433 1894
rect 10485 1891 10541 1894
rect 10593 1891 10649 1894
rect 10701 1891 10757 1894
rect 10809 1891 10865 1894
rect 10917 1891 10973 1894
rect 11025 1891 11081 1894
rect 11133 1891 11189 1894
rect 11241 1891 11297 1894
rect 11349 1891 11405 1894
rect 11457 1891 11481 1894
rect 1481 1879 11481 1891
rect 1481 1699 11481 1711
rect 1481 1696 1505 1699
rect 1557 1696 1613 1699
rect 1665 1696 1721 1699
rect 1773 1696 1829 1699
rect 1881 1696 1937 1699
rect 1989 1696 2045 1699
rect 2097 1696 2153 1699
rect 2205 1696 2261 1699
rect 2313 1696 2369 1699
rect 2421 1696 2477 1699
rect 2529 1696 2585 1699
rect 2637 1696 2693 1699
rect 2745 1696 2801 1699
rect 2853 1696 2909 1699
rect 2961 1696 3017 1699
rect 3069 1696 3125 1699
rect 3177 1696 3233 1699
rect 3285 1696 5372 1699
rect 5424 1696 5480 1699
rect 5532 1696 5588 1699
rect 5640 1696 5696 1699
rect 5748 1696 5804 1699
rect 5856 1696 5912 1699
rect 5964 1696 6020 1699
rect 6072 1696 6128 1699
rect 6180 1696 6236 1699
rect 6288 1696 6344 1699
rect 6396 1696 7749 1699
rect 7801 1696 7857 1699
rect 7909 1696 7965 1699
rect 8017 1696 8073 1699
rect 8125 1696 8181 1699
rect 8233 1696 8289 1699
rect 8341 1696 8397 1699
rect 8449 1696 8505 1699
rect 8557 1696 8613 1699
rect 8665 1696 8721 1699
rect 8773 1696 8829 1699
rect 8881 1696 8937 1699
rect 8989 1696 9045 1699
rect 9097 1696 9153 1699
rect 9205 1696 9261 1699
rect 9313 1696 9369 1699
rect 9421 1696 9477 1699
rect 9529 1696 11481 1699
rect 1481 1650 1494 1696
rect 11468 1650 11481 1696
rect 1481 1647 1505 1650
rect 1557 1647 1613 1650
rect 1665 1647 1721 1650
rect 1773 1647 1829 1650
rect 1881 1647 1937 1650
rect 1989 1647 2045 1650
rect 2097 1647 2153 1650
rect 2205 1647 2261 1650
rect 2313 1647 2369 1650
rect 2421 1647 2477 1650
rect 2529 1647 2585 1650
rect 2637 1647 2693 1650
rect 2745 1647 2801 1650
rect 2853 1647 2909 1650
rect 2961 1647 3017 1650
rect 3069 1647 3125 1650
rect 3177 1647 3233 1650
rect 3285 1647 5372 1650
rect 5424 1647 5480 1650
rect 5532 1647 5588 1650
rect 5640 1647 5696 1650
rect 5748 1647 5804 1650
rect 5856 1647 5912 1650
rect 5964 1647 6020 1650
rect 6072 1647 6128 1650
rect 6180 1647 6236 1650
rect 6288 1647 6344 1650
rect 6396 1647 7749 1650
rect 7801 1647 7857 1650
rect 7909 1647 7965 1650
rect 8017 1647 8073 1650
rect 8125 1647 8181 1650
rect 8233 1647 8289 1650
rect 8341 1647 8397 1650
rect 8449 1647 8505 1650
rect 8557 1647 8613 1650
rect 8665 1647 8721 1650
rect 8773 1647 8829 1650
rect 8881 1647 8937 1650
rect 8989 1647 9045 1650
rect 9097 1647 9153 1650
rect 9205 1647 9261 1650
rect 9313 1647 9369 1650
rect 9421 1647 9477 1650
rect 9529 1647 11481 1650
rect 1481 1635 11481 1647
rect 1213 1519 1413 1546
rect 1213 1467 1233 1519
rect 1285 1467 1341 1519
rect 1393 1467 1413 1519
rect 11549 1546 11560 6192
rect 11706 6163 11749 6192
rect 11729 6111 11749 6163
rect 11706 6055 11749 6111
rect 11729 6003 11749 6055
rect 11706 5947 11749 6003
rect 11729 5895 11749 5947
rect 11706 5839 11749 5895
rect 11729 5787 11749 5839
rect 11706 5731 11749 5787
rect 11729 5679 11749 5731
rect 11706 5623 11749 5679
rect 11729 5571 11749 5623
rect 11706 5515 11749 5571
rect 11729 5463 11749 5515
rect 11706 5407 11749 5463
rect 11729 5355 11749 5407
rect 11706 5299 11749 5355
rect 11729 5247 11749 5299
rect 11706 5191 11749 5247
rect 11729 5139 11749 5191
rect 11706 5083 11749 5139
rect 11729 5031 11749 5083
rect 11706 4975 11749 5031
rect 11729 4923 11749 4975
rect 11706 4867 11749 4923
rect 11729 4815 11749 4867
rect 11706 4759 11749 4815
rect 11729 4707 11749 4759
rect 11706 4651 11749 4707
rect 11729 4599 11749 4651
rect 11706 4543 11749 4599
rect 11729 4491 11749 4543
rect 11706 4435 11749 4491
rect 11729 4383 11749 4435
rect 11706 4327 11749 4383
rect 11729 4275 11749 4327
rect 11706 4219 11749 4275
rect 11729 4167 11749 4219
rect 11706 4111 11749 4167
rect 11729 4059 11749 4111
rect 11706 4003 11749 4059
rect 11729 3951 11749 4003
rect 11706 3895 11749 3951
rect 11729 3843 11749 3895
rect 11706 3787 11749 3843
rect 11729 3735 11749 3787
rect 11706 3679 11749 3735
rect 11729 3627 11749 3679
rect 11706 3571 11749 3627
rect 11729 3519 11749 3571
rect 11706 3463 11749 3519
rect 11729 3411 11749 3463
rect 11706 3355 11749 3411
rect 11729 3303 11749 3355
rect 11706 3247 11749 3303
rect 11729 3195 11749 3247
rect 11706 3139 11749 3195
rect 11729 3087 11749 3139
rect 11706 3031 11749 3087
rect 11729 2979 11749 3031
rect 11706 2923 11749 2979
rect 11729 2871 11749 2923
rect 11706 2815 11749 2871
rect 11729 2763 11749 2815
rect 11706 2707 11749 2763
rect 11729 2655 11749 2707
rect 11706 2599 11749 2655
rect 11729 2547 11749 2599
rect 11706 2491 11749 2547
rect 11729 2439 11749 2491
rect 11706 2383 11749 2439
rect 11729 2331 11749 2383
rect 11706 2275 11749 2331
rect 11729 2223 11749 2275
rect 11706 2167 11749 2223
rect 11729 2115 11749 2167
rect 11706 2059 11749 2115
rect 11729 2007 11749 2059
rect 11706 1951 11749 2007
rect 11729 1899 11749 1951
rect 11706 1843 11749 1899
rect 11729 1791 11749 1843
rect 11706 1735 11749 1791
rect 11729 1683 11749 1735
rect 11706 1627 11749 1683
rect 11729 1575 11749 1627
rect 11706 1546 11749 1575
rect 11549 1519 11749 1546
rect 11549 1467 11569 1519
rect 11621 1467 11677 1519
rect 11729 1467 11749 1519
rect 1213 1298 1413 1467
rect 1481 1455 11481 1467
rect 1481 1452 3433 1455
rect 3485 1452 3541 1455
rect 3593 1452 3649 1455
rect 3701 1452 3757 1455
rect 3809 1452 3865 1455
rect 3917 1452 3973 1455
rect 4025 1452 4081 1455
rect 4133 1452 4189 1455
rect 4241 1452 4297 1455
rect 4349 1452 4405 1455
rect 4457 1452 4513 1455
rect 4565 1452 4621 1455
rect 4673 1452 4729 1455
rect 4781 1452 4837 1455
rect 4889 1452 4945 1455
rect 4997 1452 5053 1455
rect 5105 1452 5161 1455
rect 5213 1452 6566 1455
rect 6618 1452 6674 1455
rect 6726 1452 6782 1455
rect 6834 1452 6890 1455
rect 6942 1452 6998 1455
rect 7050 1452 7106 1455
rect 7158 1452 7214 1455
rect 7266 1452 7322 1455
rect 7374 1452 7430 1455
rect 7482 1452 7538 1455
rect 7590 1452 9677 1455
rect 9729 1452 9785 1455
rect 9837 1452 9893 1455
rect 9945 1452 10001 1455
rect 10053 1452 10109 1455
rect 10161 1452 10217 1455
rect 10269 1452 10325 1455
rect 10377 1452 10433 1455
rect 10485 1452 10541 1455
rect 10593 1452 10649 1455
rect 10701 1452 10757 1455
rect 10809 1452 10865 1455
rect 10917 1452 10973 1455
rect 11025 1452 11081 1455
rect 11133 1452 11189 1455
rect 11241 1452 11297 1455
rect 11349 1452 11405 1455
rect 11457 1452 11481 1455
rect 1481 1406 1494 1452
rect 11468 1406 11481 1452
rect 1481 1403 3433 1406
rect 3485 1403 3541 1406
rect 3593 1403 3649 1406
rect 3701 1403 3757 1406
rect 3809 1403 3865 1406
rect 3917 1403 3973 1406
rect 4025 1403 4081 1406
rect 4133 1403 4189 1406
rect 4241 1403 4297 1406
rect 4349 1403 4405 1406
rect 4457 1403 4513 1406
rect 4565 1403 4621 1406
rect 4673 1403 4729 1406
rect 4781 1403 4837 1406
rect 4889 1403 4945 1406
rect 4997 1403 5053 1406
rect 5105 1403 5161 1406
rect 5213 1403 6566 1406
rect 6618 1403 6674 1406
rect 6726 1403 6782 1406
rect 6834 1403 6890 1406
rect 6942 1403 6998 1406
rect 7050 1403 7106 1406
rect 7158 1403 7214 1406
rect 7266 1403 7322 1406
rect 7374 1403 7430 1406
rect 7482 1403 7538 1406
rect 7590 1403 9677 1406
rect 9729 1403 9785 1406
rect 9837 1403 9893 1406
rect 9945 1403 10001 1406
rect 10053 1403 10109 1406
rect 10161 1403 10217 1406
rect 10269 1403 10325 1406
rect 10377 1403 10433 1406
rect 10485 1403 10541 1406
rect 10593 1403 10649 1406
rect 10701 1403 10757 1406
rect 10809 1403 10865 1406
rect 10917 1403 10973 1406
rect 11025 1403 11081 1406
rect 11133 1403 11189 1406
rect 11241 1403 11297 1406
rect 11349 1403 11405 1406
rect 11457 1403 11481 1406
rect 1481 1391 11481 1403
rect 11549 1298 11749 1467
rect 1213 1098 11749 1298
rect 12001 1011 12012 6713
rect 950 1000 12012 1011
rect 950 654 1058 1000
rect 11904 654 12012 1000
rect 12358 654 12369 24700
rect 593 643 12369 654
rect 12551 411 12562 24943
rect 400 400 12562 411
rect 400 361 508 400
rect 400 309 406 361
rect 458 309 508 361
rect 400 253 508 309
rect 400 201 406 253
rect 458 201 508 253
rect 400 145 508 201
rect 400 93 406 145
rect 458 93 508 145
rect 400 54 508 93
rect 12454 54 12562 400
rect 12908 54 12919 25300
rect 43 43 12919 54
<< via1 >>
rect 82 25209 134 25261
rect 190 25209 242 25261
rect 298 25209 350 25261
rect 406 25209 458 25261
rect 514 25209 566 25261
rect 622 25209 674 25261
rect 730 25209 782 25261
rect 838 25209 890 25261
rect 946 25209 998 25261
rect 1054 25209 1106 25261
rect 3433 25209 3485 25261
rect 3541 25209 3593 25261
rect 3649 25209 3701 25261
rect 3757 25209 3809 25261
rect 3865 25209 3917 25261
rect 3973 25209 4025 25261
rect 4081 25209 4133 25261
rect 4189 25209 4241 25261
rect 4297 25209 4349 25261
rect 4405 25209 4457 25261
rect 4513 25209 4565 25261
rect 4621 25209 4673 25261
rect 4729 25209 4781 25261
rect 4837 25209 4889 25261
rect 4945 25209 4997 25261
rect 5053 25209 5105 25261
rect 5161 25209 5213 25261
rect 6566 25209 6618 25261
rect 6674 25209 6726 25261
rect 6782 25209 6834 25261
rect 6890 25209 6942 25261
rect 6998 25209 7050 25261
rect 7106 25209 7158 25261
rect 7214 25209 7266 25261
rect 7322 25209 7374 25261
rect 7430 25209 7482 25261
rect 7538 25209 7590 25261
rect 9677 25209 9729 25261
rect 9785 25209 9837 25261
rect 9893 25209 9945 25261
rect 10001 25209 10053 25261
rect 10109 25209 10161 25261
rect 10217 25209 10269 25261
rect 10325 25209 10377 25261
rect 10433 25209 10485 25261
rect 10541 25209 10593 25261
rect 10649 25209 10701 25261
rect 10757 25209 10809 25261
rect 10865 25209 10917 25261
rect 10973 25209 11025 25261
rect 11081 25209 11133 25261
rect 11189 25209 11241 25261
rect 11297 25209 11349 25261
rect 11405 25209 11457 25261
rect 82 25101 134 25153
rect 190 25101 242 25153
rect 298 25101 350 25153
rect 406 25101 458 25153
rect 514 25101 566 25153
rect 622 25101 674 25153
rect 730 25101 782 25153
rect 838 25101 890 25153
rect 946 25101 998 25153
rect 1054 25101 1106 25153
rect 3433 25101 3485 25153
rect 3541 25101 3593 25153
rect 3649 25101 3701 25153
rect 3757 25101 3809 25153
rect 3865 25101 3917 25153
rect 3973 25101 4025 25153
rect 4081 25101 4133 25153
rect 4189 25101 4241 25153
rect 4297 25101 4349 25153
rect 4405 25101 4457 25153
rect 4513 25101 4565 25153
rect 4621 25101 4673 25153
rect 4729 25101 4781 25153
rect 4837 25101 4889 25153
rect 4945 25101 4997 25153
rect 5053 25101 5105 25153
rect 5161 25101 5213 25153
rect 6566 25101 6618 25153
rect 6674 25101 6726 25153
rect 6782 25101 6834 25153
rect 6890 25101 6942 25153
rect 6998 25101 7050 25153
rect 7106 25101 7158 25153
rect 7214 25101 7266 25153
rect 7322 25101 7374 25153
rect 7430 25101 7482 25153
rect 7538 25101 7590 25153
rect 9677 25101 9729 25153
rect 9785 25101 9837 25153
rect 9893 25101 9945 25153
rect 10001 25101 10053 25153
rect 10109 25101 10161 25153
rect 10217 25101 10269 25153
rect 10325 25101 10377 25153
rect 10433 25101 10485 25153
rect 10541 25101 10593 25153
rect 10649 25101 10701 25153
rect 10757 25101 10809 25153
rect 10865 25101 10917 25153
rect 10973 25101 11025 25153
rect 11081 25101 11133 25153
rect 11189 25101 11241 25153
rect 11297 25101 11349 25153
rect 11405 25101 11457 25153
rect 82 24993 134 25045
rect 190 24993 242 25045
rect 298 24993 350 25045
rect 406 24993 458 25045
rect 514 24993 566 25045
rect 622 24993 674 25045
rect 730 24993 782 25045
rect 838 24993 890 25045
rect 946 24993 998 25045
rect 1054 24993 1106 25045
rect 3433 24993 3485 25045
rect 3541 24993 3593 25045
rect 3649 24993 3701 25045
rect 3757 24993 3809 25045
rect 3865 24993 3917 25045
rect 3973 24993 4025 25045
rect 4081 24993 4133 25045
rect 4189 24993 4241 25045
rect 4297 24993 4349 25045
rect 4405 24993 4457 25045
rect 4513 24993 4565 25045
rect 4621 24993 4673 25045
rect 4729 24993 4781 25045
rect 4837 24993 4889 25045
rect 4945 24993 4997 25045
rect 5053 24993 5105 25045
rect 5161 24993 5213 25045
rect 6566 24993 6618 25045
rect 6674 24993 6726 25045
rect 6782 24993 6834 25045
rect 6890 24993 6942 25045
rect 6998 24993 7050 25045
rect 7106 24993 7158 25045
rect 7214 24993 7266 25045
rect 7322 24993 7374 25045
rect 7430 24993 7482 25045
rect 7538 24993 7590 25045
rect 9677 24993 9729 25045
rect 9785 24993 9837 25045
rect 9893 24993 9945 25045
rect 10001 24993 10053 25045
rect 10109 24993 10161 25045
rect 10217 24993 10269 25045
rect 10325 24993 10377 25045
rect 10433 24993 10485 25045
rect 10541 24993 10593 25045
rect 10649 24993 10701 25045
rect 10757 24993 10809 25045
rect 10865 24993 10917 25045
rect 10973 24993 11025 25045
rect 11081 24993 11133 25045
rect 11189 24993 11241 25045
rect 11297 24993 11349 25045
rect 11405 24993 11457 25045
rect 93 24801 145 24853
rect 201 24801 253 24853
rect 309 24801 361 24853
rect 93 24693 145 24745
rect 201 24693 253 24745
rect 309 24693 361 24745
rect 93 24585 145 24637
rect 201 24585 253 24637
rect 309 24585 361 24637
rect 93 24477 145 24529
rect 201 24477 253 24529
rect 309 24477 361 24529
rect 93 24369 145 24421
rect 201 24369 253 24421
rect 309 24369 361 24421
rect 93 24261 145 24313
rect 201 24261 253 24313
rect 309 24261 361 24313
rect 93 24153 145 24205
rect 201 24153 253 24205
rect 309 24153 361 24205
rect 93 24045 145 24097
rect 201 24045 253 24097
rect 309 24045 361 24097
rect 93 23937 145 23989
rect 201 23937 253 23989
rect 309 23937 361 23989
rect 93 23829 145 23881
rect 201 23829 253 23881
rect 309 23829 361 23881
rect 93 23721 145 23773
rect 201 23721 253 23773
rect 309 23721 361 23773
rect 93 23613 145 23665
rect 201 23613 253 23665
rect 309 23613 361 23665
rect 93 23505 145 23557
rect 201 23505 253 23557
rect 309 23505 361 23557
rect 93 23397 145 23449
rect 201 23397 253 23449
rect 309 23397 361 23449
rect 93 23289 145 23341
rect 201 23289 253 23341
rect 309 23289 361 23341
rect 93 23181 145 23233
rect 201 23181 253 23233
rect 309 23181 361 23233
rect 93 23073 145 23125
rect 201 23073 253 23125
rect 309 23073 361 23125
rect 93 22965 145 23017
rect 201 22965 253 23017
rect 309 22965 361 23017
rect 93 22857 145 22909
rect 201 22857 253 22909
rect 309 22857 361 22909
rect 93 22749 145 22801
rect 201 22749 253 22801
rect 309 22749 361 22801
rect 93 22641 145 22693
rect 201 22641 253 22693
rect 309 22641 361 22693
rect 93 22533 145 22585
rect 201 22533 253 22585
rect 309 22533 361 22585
rect 93 22425 145 22477
rect 201 22425 253 22477
rect 309 22425 361 22477
rect 93 22317 145 22369
rect 201 22317 253 22369
rect 309 22317 361 22369
rect 93 22209 145 22261
rect 201 22209 253 22261
rect 309 22209 361 22261
rect 93 22101 145 22153
rect 201 22101 253 22153
rect 309 22101 361 22153
rect 93 21993 145 22045
rect 201 21993 253 22045
rect 309 21993 361 22045
rect 93 21885 145 21937
rect 201 21885 253 21937
rect 309 21885 361 21937
rect 93 21777 145 21829
rect 201 21777 253 21829
rect 309 21777 361 21829
rect 93 21669 145 21721
rect 201 21669 253 21721
rect 309 21669 361 21721
rect 93 21561 145 21613
rect 201 21561 253 21613
rect 309 21561 361 21613
rect 93 21453 145 21505
rect 201 21453 253 21505
rect 309 21453 361 21505
rect 93 21345 145 21397
rect 201 21345 253 21397
rect 309 21345 361 21397
rect 93 21237 145 21289
rect 201 21237 253 21289
rect 309 21237 361 21289
rect 93 21129 145 21181
rect 201 21129 253 21181
rect 309 21129 361 21181
rect 93 21021 145 21073
rect 201 21021 253 21073
rect 309 21021 361 21073
rect 93 20913 145 20965
rect 201 20913 253 20965
rect 309 20913 361 20965
rect 93 20805 145 20857
rect 201 20805 253 20857
rect 309 20805 361 20857
rect 93 20697 145 20749
rect 201 20697 253 20749
rect 309 20697 361 20749
rect 93 20589 145 20641
rect 201 20589 253 20641
rect 309 20589 361 20641
rect 93 20481 145 20533
rect 201 20481 253 20533
rect 309 20481 361 20533
rect 93 20373 145 20425
rect 201 20373 253 20425
rect 309 20373 361 20425
rect 93 20265 145 20317
rect 201 20265 253 20317
rect 309 20265 361 20317
rect 93 20157 145 20209
rect 201 20157 253 20209
rect 309 20157 361 20209
rect 93 20049 145 20101
rect 201 20049 253 20101
rect 309 20049 361 20101
rect 93 19941 145 19993
rect 201 19941 253 19993
rect 309 19941 361 19993
rect 93 19833 145 19885
rect 201 19833 253 19885
rect 309 19833 361 19885
rect 93 19725 145 19777
rect 201 19725 253 19777
rect 309 19725 361 19777
rect 93 19617 145 19669
rect 201 19617 253 19669
rect 309 19617 361 19669
rect 93 19509 145 19561
rect 201 19509 253 19561
rect 309 19509 361 19561
rect 93 19401 145 19453
rect 201 19401 253 19453
rect 309 19401 361 19453
rect 93 19293 145 19345
rect 201 19293 253 19345
rect 309 19293 361 19345
rect 93 19185 145 19237
rect 201 19185 253 19237
rect 309 19185 361 19237
rect 93 19077 145 19129
rect 201 19077 253 19129
rect 309 19077 361 19129
rect 93 18969 145 19021
rect 201 18969 253 19021
rect 309 18969 361 19021
rect 93 18861 145 18913
rect 201 18861 253 18913
rect 309 18861 361 18913
rect 93 18753 145 18805
rect 201 18753 253 18805
rect 309 18753 361 18805
rect 93 18645 145 18697
rect 201 18645 253 18697
rect 309 18645 361 18697
rect 93 18537 145 18589
rect 201 18537 253 18589
rect 309 18537 361 18589
rect 93 18429 145 18481
rect 201 18429 253 18481
rect 309 18429 361 18481
rect 93 18321 145 18373
rect 201 18321 253 18373
rect 309 18321 361 18373
rect 93 18213 145 18265
rect 201 18213 253 18265
rect 309 18213 361 18265
rect 93 18105 145 18157
rect 201 18105 253 18157
rect 309 18105 361 18157
rect 93 17997 145 18049
rect 201 17997 253 18049
rect 309 17997 361 18049
rect 93 17889 145 17941
rect 201 17889 253 17941
rect 309 17889 361 17941
rect 93 17781 145 17833
rect 201 17781 253 17833
rect 309 17781 361 17833
rect 93 17673 145 17725
rect 201 17673 253 17725
rect 309 17673 361 17725
rect 93 17565 145 17617
rect 201 17565 253 17617
rect 309 17565 361 17617
rect 93 17457 145 17509
rect 201 17457 253 17509
rect 309 17457 361 17509
rect 93 17349 145 17401
rect 201 17349 253 17401
rect 309 17349 361 17401
rect 93 17241 145 17293
rect 201 17241 253 17293
rect 309 17241 361 17293
rect 93 17133 145 17185
rect 201 17133 253 17185
rect 309 17133 361 17185
rect 93 17025 145 17077
rect 201 17025 253 17077
rect 309 17025 361 17077
rect 93 16917 145 16969
rect 201 16917 253 16969
rect 309 16917 361 16969
rect 93 16809 145 16861
rect 201 16809 253 16861
rect 309 16809 361 16861
rect 93 16701 145 16753
rect 201 16701 253 16753
rect 309 16701 361 16753
rect 93 16593 145 16645
rect 201 16593 253 16645
rect 309 16593 361 16645
rect 93 16485 145 16537
rect 201 16485 253 16537
rect 309 16485 361 16537
rect 93 16377 145 16429
rect 201 16377 253 16429
rect 309 16377 361 16429
rect 93 16269 145 16321
rect 201 16269 253 16321
rect 309 16269 361 16321
rect 93 16161 145 16213
rect 201 16161 253 16213
rect 309 16161 361 16213
rect 93 16053 145 16105
rect 201 16053 253 16105
rect 309 16053 361 16105
rect 93 15945 145 15997
rect 201 15945 253 15997
rect 309 15945 361 15997
rect 93 15837 145 15889
rect 201 15837 253 15889
rect 309 15837 361 15889
rect 93 15729 145 15781
rect 201 15729 253 15781
rect 309 15729 361 15781
rect 93 15621 145 15673
rect 201 15621 253 15673
rect 309 15621 361 15673
rect 93 15513 145 15565
rect 201 15513 253 15565
rect 309 15513 361 15565
rect 93 15405 145 15457
rect 201 15405 253 15457
rect 309 15405 361 15457
rect 93 15297 145 15349
rect 201 15297 253 15349
rect 309 15297 361 15349
rect 93 15189 145 15241
rect 201 15189 253 15241
rect 309 15189 361 15241
rect 93 15081 145 15133
rect 201 15081 253 15133
rect 309 15081 361 15133
rect 93 14973 145 15025
rect 201 14973 253 15025
rect 309 14973 361 15025
rect 93 14865 145 14917
rect 201 14865 253 14917
rect 309 14865 361 14917
rect 93 14757 145 14809
rect 201 14757 253 14809
rect 309 14757 361 14809
rect 93 14649 145 14701
rect 201 14649 253 14701
rect 309 14649 361 14701
rect 93 14541 145 14593
rect 201 14541 253 14593
rect 309 14541 361 14593
rect 93 14433 145 14485
rect 201 14433 253 14485
rect 309 14433 361 14485
rect 93 14325 145 14377
rect 201 14325 253 14377
rect 309 14325 361 14377
rect 93 14217 145 14269
rect 201 14217 253 14269
rect 309 14217 361 14269
rect 93 14109 145 14161
rect 201 14109 253 14161
rect 309 14109 361 14161
rect 93 14001 145 14053
rect 201 14001 253 14053
rect 309 14001 361 14053
rect 93 13893 145 13945
rect 201 13893 253 13945
rect 309 13893 361 13945
rect 93 13785 145 13837
rect 201 13785 253 13837
rect 309 13785 361 13837
rect 93 13677 145 13729
rect 201 13677 253 13729
rect 309 13677 361 13729
rect 93 13569 145 13621
rect 201 13569 253 13621
rect 309 13569 361 13621
rect 93 13461 145 13513
rect 201 13461 253 13513
rect 309 13461 361 13513
rect 93 13353 145 13405
rect 201 13353 253 13405
rect 309 13353 361 13405
rect 93 13245 145 13297
rect 201 13245 253 13297
rect 309 13245 361 13297
rect 93 13137 145 13189
rect 201 13137 253 13189
rect 309 13137 361 13189
rect 93 13029 145 13081
rect 201 13029 253 13081
rect 309 13029 361 13081
rect 93 12921 145 12973
rect 201 12921 253 12973
rect 309 12921 361 12973
rect 93 12813 145 12865
rect 201 12813 253 12865
rect 309 12813 361 12865
rect 93 12705 145 12757
rect 201 12705 253 12757
rect 309 12705 361 12757
rect 93 12597 145 12649
rect 201 12597 253 12649
rect 309 12597 361 12649
rect 93 12489 145 12541
rect 201 12489 253 12541
rect 309 12489 361 12541
rect 93 12381 145 12433
rect 201 12381 253 12433
rect 309 12381 361 12433
rect 93 12273 145 12325
rect 201 12273 253 12325
rect 309 12273 361 12325
rect 93 12165 145 12217
rect 201 12165 253 12217
rect 309 12165 361 12217
rect 93 12057 145 12109
rect 201 12057 253 12109
rect 309 12057 361 12109
rect 93 11949 145 12001
rect 201 11949 253 12001
rect 309 11949 361 12001
rect 93 11841 145 11893
rect 201 11841 253 11893
rect 309 11841 361 11893
rect 93 11733 145 11785
rect 201 11733 253 11785
rect 309 11733 361 11785
rect 93 11625 145 11677
rect 201 11625 253 11677
rect 309 11625 361 11677
rect 93 11517 145 11569
rect 201 11517 253 11569
rect 309 11517 361 11569
rect 93 11409 145 11461
rect 201 11409 253 11461
rect 309 11409 361 11461
rect 93 11301 145 11353
rect 201 11301 253 11353
rect 309 11301 361 11353
rect 93 11193 145 11245
rect 201 11193 253 11245
rect 309 11193 361 11245
rect 93 11085 145 11137
rect 201 11085 253 11137
rect 309 11085 361 11137
rect 93 10977 145 11029
rect 201 10977 253 11029
rect 309 10977 361 11029
rect 93 10869 145 10921
rect 201 10869 253 10921
rect 309 10869 361 10921
rect 93 10761 145 10813
rect 201 10761 253 10813
rect 309 10761 361 10813
rect 93 10653 145 10705
rect 201 10653 253 10705
rect 309 10653 361 10705
rect 93 10545 145 10597
rect 201 10545 253 10597
rect 309 10545 361 10597
rect 93 10437 145 10489
rect 201 10437 253 10489
rect 309 10437 361 10489
rect 93 10329 145 10381
rect 201 10329 253 10381
rect 309 10329 361 10381
rect 93 10221 145 10273
rect 201 10221 253 10273
rect 309 10221 361 10273
rect 93 10113 145 10165
rect 201 10113 253 10165
rect 309 10113 361 10165
rect 93 10005 145 10057
rect 201 10005 253 10057
rect 309 10005 361 10057
rect 93 9897 145 9949
rect 201 9897 253 9949
rect 309 9897 361 9949
rect 93 9789 145 9841
rect 201 9789 253 9841
rect 309 9789 361 9841
rect 93 9681 145 9733
rect 201 9681 253 9733
rect 309 9681 361 9733
rect 93 9573 145 9625
rect 201 9573 253 9625
rect 309 9573 361 9625
rect 93 9465 145 9517
rect 201 9465 253 9517
rect 309 9465 361 9517
rect 93 9357 145 9409
rect 201 9357 253 9409
rect 309 9357 361 9409
rect 93 9249 145 9301
rect 201 9249 253 9301
rect 309 9249 361 9301
rect 93 9141 145 9193
rect 201 9141 253 9193
rect 309 9141 361 9193
rect 93 9033 145 9085
rect 201 9033 253 9085
rect 309 9033 361 9085
rect 93 8925 145 8977
rect 201 8925 253 8977
rect 309 8925 361 8977
rect 93 8817 145 8869
rect 201 8817 253 8869
rect 309 8817 361 8869
rect 93 8709 145 8761
rect 201 8709 253 8761
rect 309 8709 361 8761
rect 93 8601 145 8653
rect 201 8601 253 8653
rect 309 8601 361 8653
rect 93 8493 145 8545
rect 201 8493 253 8545
rect 309 8493 361 8545
rect 93 8385 145 8437
rect 201 8385 253 8437
rect 309 8385 361 8437
rect 93 8277 145 8329
rect 201 8277 253 8329
rect 309 8277 361 8329
rect 93 8169 145 8221
rect 201 8169 253 8221
rect 309 8169 361 8221
rect 93 8061 145 8113
rect 201 8061 253 8113
rect 309 8061 361 8113
rect 93 7953 145 8005
rect 201 7953 253 8005
rect 309 7953 361 8005
rect 93 7845 145 7897
rect 201 7845 253 7897
rect 309 7845 361 7897
rect 93 7737 145 7789
rect 201 7737 253 7789
rect 309 7737 361 7789
rect 93 7629 145 7681
rect 201 7629 253 7681
rect 309 7629 361 7681
rect 93 7521 145 7573
rect 201 7521 253 7573
rect 309 7521 361 7573
rect 93 7413 145 7465
rect 201 7413 253 7465
rect 309 7413 361 7465
rect 93 7305 145 7357
rect 201 7305 253 7357
rect 309 7305 361 7357
rect 93 7197 145 7249
rect 201 7197 253 7249
rect 309 7197 361 7249
rect 93 7089 145 7141
rect 201 7089 253 7141
rect 309 7089 361 7141
rect 93 6981 145 7033
rect 201 6981 253 7033
rect 309 6981 361 7033
rect 93 6873 145 6925
rect 201 6873 253 6925
rect 309 6873 361 6925
rect 93 6765 145 6817
rect 201 6765 253 6817
rect 309 6765 361 6817
rect 93 6657 145 6709
rect 201 6657 253 6709
rect 309 6657 361 6709
rect 93 6549 145 6601
rect 201 6549 253 6601
rect 309 6549 361 6601
rect 93 6441 145 6493
rect 201 6441 253 6493
rect 309 6441 361 6493
rect 93 6333 145 6385
rect 201 6333 253 6385
rect 309 6333 361 6385
rect 93 6225 145 6277
rect 201 6225 253 6277
rect 309 6225 361 6277
rect 93 6117 145 6169
rect 201 6117 253 6169
rect 309 6117 361 6169
rect 93 6009 145 6061
rect 201 6009 253 6061
rect 309 6009 361 6061
rect 93 5901 145 5953
rect 201 5901 253 5953
rect 309 5901 361 5953
rect 93 5793 145 5845
rect 201 5793 253 5845
rect 309 5793 361 5845
rect 93 5685 145 5737
rect 201 5685 253 5737
rect 309 5685 361 5737
rect 93 5577 145 5629
rect 201 5577 253 5629
rect 309 5577 361 5629
rect 93 5469 145 5521
rect 201 5469 253 5521
rect 309 5469 361 5521
rect 93 5361 145 5413
rect 201 5361 253 5413
rect 309 5361 361 5413
rect 93 5253 145 5305
rect 201 5253 253 5305
rect 309 5253 361 5305
rect 93 5145 145 5197
rect 201 5145 253 5197
rect 309 5145 361 5197
rect 93 5037 145 5089
rect 201 5037 253 5089
rect 309 5037 361 5089
rect 93 4929 145 4981
rect 201 4929 253 4981
rect 309 4929 361 4981
rect 93 4821 145 4873
rect 201 4821 253 4873
rect 309 4821 361 4873
rect 93 4713 145 4765
rect 201 4713 253 4765
rect 309 4713 361 4765
rect 93 4605 145 4657
rect 201 4605 253 4657
rect 309 4605 361 4657
rect 93 4497 145 4549
rect 201 4497 253 4549
rect 309 4497 361 4549
rect 93 4389 145 4441
rect 201 4389 253 4441
rect 309 4389 361 4441
rect 93 4281 145 4333
rect 201 4281 253 4333
rect 309 4281 361 4333
rect 93 4173 145 4225
rect 201 4173 253 4225
rect 309 4173 361 4225
rect 93 4065 145 4117
rect 201 4065 253 4117
rect 309 4065 361 4117
rect 93 3957 145 4009
rect 201 3957 253 4009
rect 309 3957 361 4009
rect 93 3849 145 3901
rect 201 3849 253 3901
rect 309 3849 361 3901
rect 93 3741 145 3793
rect 201 3741 253 3793
rect 309 3741 361 3793
rect 93 3633 145 3685
rect 201 3633 253 3685
rect 309 3633 361 3685
rect 93 3525 145 3577
rect 201 3525 253 3577
rect 309 3525 361 3577
rect 93 3417 145 3469
rect 201 3417 253 3469
rect 309 3417 361 3469
rect 93 3309 145 3361
rect 201 3309 253 3361
rect 309 3309 361 3361
rect 93 3201 145 3253
rect 201 3201 253 3253
rect 309 3201 361 3253
rect 93 3093 145 3145
rect 201 3093 253 3145
rect 309 3093 361 3145
rect 93 2985 145 3037
rect 201 2985 253 3037
rect 309 2985 361 3037
rect 93 2877 145 2929
rect 201 2877 253 2929
rect 309 2877 361 2929
rect 93 2769 145 2821
rect 201 2769 253 2821
rect 309 2769 361 2821
rect 93 2661 145 2713
rect 201 2661 253 2713
rect 309 2661 361 2713
rect 93 2553 145 2605
rect 201 2553 253 2605
rect 309 2553 361 2605
rect 93 2445 145 2497
rect 201 2445 253 2497
rect 309 2445 361 2497
rect 93 2337 145 2389
rect 201 2337 253 2389
rect 309 2337 361 2389
rect 93 2229 145 2281
rect 201 2229 253 2281
rect 309 2229 361 2281
rect 93 2121 145 2173
rect 201 2121 253 2173
rect 309 2121 361 2173
rect 93 2013 145 2065
rect 201 2013 253 2065
rect 309 2013 361 2065
rect 93 1905 145 1957
rect 201 1905 253 1957
rect 309 1905 361 1957
rect 93 1797 145 1849
rect 201 1797 253 1849
rect 309 1797 361 1849
rect 93 1689 145 1741
rect 201 1689 253 1741
rect 309 1689 361 1741
rect 93 1581 145 1633
rect 201 1581 253 1633
rect 309 1581 361 1633
rect 93 1473 145 1525
rect 201 1473 253 1525
rect 309 1473 361 1525
rect 93 1365 145 1417
rect 201 1365 253 1417
rect 309 1365 361 1417
rect 93 1257 145 1309
rect 201 1257 253 1309
rect 309 1257 361 1309
rect 93 1149 145 1201
rect 201 1149 253 1201
rect 309 1149 361 1201
rect 93 1041 145 1093
rect 201 1041 253 1093
rect 309 1041 361 1093
rect 93 933 145 985
rect 201 933 253 985
rect 309 933 361 985
rect 93 825 145 877
rect 201 825 253 877
rect 309 825 361 877
rect 93 717 145 769
rect 201 717 253 769
rect 309 717 361 769
rect 93 609 145 661
rect 201 609 253 661
rect 309 609 361 661
rect 93 501 145 553
rect 201 501 253 553
rect 309 501 361 553
rect 1505 24609 1557 24661
rect 1613 24609 1665 24661
rect 1721 24609 1773 24661
rect 1829 24609 1881 24661
rect 1937 24609 1989 24661
rect 2045 24609 2097 24661
rect 2153 24609 2205 24661
rect 2261 24609 2313 24661
rect 2369 24609 2421 24661
rect 2477 24609 2529 24661
rect 2585 24609 2637 24661
rect 2693 24609 2745 24661
rect 2801 24609 2853 24661
rect 2909 24609 2961 24661
rect 3017 24609 3069 24661
rect 3125 24609 3177 24661
rect 3233 24609 3285 24661
rect 5372 24609 5424 24661
rect 5480 24609 5532 24661
rect 5588 24609 5640 24661
rect 5696 24609 5748 24661
rect 5804 24609 5856 24661
rect 5912 24609 5964 24661
rect 6020 24609 6072 24661
rect 6128 24609 6180 24661
rect 6236 24609 6288 24661
rect 6344 24609 6396 24661
rect 7749 24609 7801 24661
rect 7857 24609 7909 24661
rect 7965 24609 8017 24661
rect 8073 24609 8125 24661
rect 8181 24609 8233 24661
rect 8289 24609 8341 24661
rect 8397 24609 8449 24661
rect 8505 24609 8557 24661
rect 8613 24609 8665 24661
rect 8721 24609 8773 24661
rect 8829 24609 8881 24661
rect 8937 24609 8989 24661
rect 9045 24609 9097 24661
rect 9153 24609 9205 24661
rect 9261 24609 9313 24661
rect 9369 24609 9421 24661
rect 9477 24609 9529 24661
rect 1505 24501 1557 24553
rect 1613 24501 1665 24553
rect 1721 24501 1773 24553
rect 1829 24501 1881 24553
rect 1937 24501 1989 24553
rect 2045 24501 2097 24553
rect 2153 24501 2205 24553
rect 2261 24501 2313 24553
rect 2369 24501 2421 24553
rect 2477 24501 2529 24553
rect 2585 24501 2637 24553
rect 2693 24501 2745 24553
rect 2801 24501 2853 24553
rect 2909 24501 2961 24553
rect 3017 24501 3069 24553
rect 3125 24501 3177 24553
rect 3233 24501 3285 24553
rect 5372 24501 5424 24553
rect 5480 24501 5532 24553
rect 5588 24501 5640 24553
rect 5696 24501 5748 24553
rect 5804 24501 5856 24553
rect 5912 24501 5964 24553
rect 6020 24501 6072 24553
rect 6128 24501 6180 24553
rect 6236 24501 6288 24553
rect 6344 24501 6396 24553
rect 7749 24501 7801 24553
rect 7857 24501 7909 24553
rect 7965 24501 8017 24553
rect 8073 24501 8125 24553
rect 8181 24501 8233 24553
rect 8289 24501 8341 24553
rect 8397 24501 8449 24553
rect 8505 24501 8557 24553
rect 8613 24501 8665 24553
rect 8721 24501 8773 24553
rect 8829 24501 8881 24553
rect 8937 24501 8989 24553
rect 9045 24501 9097 24553
rect 9153 24501 9205 24553
rect 9261 24501 9313 24553
rect 9369 24501 9421 24553
rect 9477 24501 9529 24553
rect 1505 24393 1557 24445
rect 1613 24393 1665 24445
rect 1721 24393 1773 24445
rect 1829 24393 1881 24445
rect 1937 24393 1989 24445
rect 2045 24393 2097 24445
rect 2153 24393 2205 24445
rect 2261 24393 2313 24445
rect 2369 24393 2421 24445
rect 2477 24393 2529 24445
rect 2585 24393 2637 24445
rect 2693 24393 2745 24445
rect 2801 24393 2853 24445
rect 2909 24393 2961 24445
rect 3017 24393 3069 24445
rect 3125 24393 3177 24445
rect 3233 24393 3285 24445
rect 5372 24393 5424 24445
rect 5480 24393 5532 24445
rect 5588 24393 5640 24445
rect 5696 24393 5748 24445
rect 5804 24393 5856 24445
rect 5912 24393 5964 24445
rect 6020 24393 6072 24445
rect 6128 24393 6180 24445
rect 6236 24393 6288 24445
rect 6344 24393 6396 24445
rect 7749 24393 7801 24445
rect 7857 24393 7909 24445
rect 7965 24393 8017 24445
rect 8073 24393 8125 24445
rect 8181 24393 8233 24445
rect 8289 24393 8341 24445
rect 8397 24393 8449 24445
rect 8505 24393 8557 24445
rect 8613 24393 8665 24445
rect 8721 24393 8773 24445
rect 8829 24393 8881 24445
rect 8937 24393 8989 24445
rect 9045 24393 9097 24445
rect 9153 24393 9205 24445
rect 9261 24393 9313 24445
rect 9369 24393 9421 24445
rect 9477 24393 9529 24445
rect 12051 24585 12103 24637
rect 12159 24585 12211 24637
rect 12267 24585 12319 24637
rect 12051 24477 12103 24529
rect 12159 24477 12211 24529
rect 12267 24477 12319 24529
rect 12051 24369 12103 24421
rect 12159 24369 12211 24421
rect 12267 24369 12319 24421
rect 3433 23948 3485 23951
rect 3541 23948 3593 23951
rect 3649 23948 3701 23951
rect 3757 23948 3809 23951
rect 3865 23948 3917 23951
rect 3973 23948 4025 23951
rect 4081 23948 4133 23951
rect 4189 23948 4241 23951
rect 4297 23948 4349 23951
rect 4405 23948 4457 23951
rect 4513 23948 4565 23951
rect 4621 23948 4673 23951
rect 4729 23948 4781 23951
rect 4837 23948 4889 23951
rect 4945 23948 4997 23951
rect 5053 23948 5105 23951
rect 5161 23948 5213 23951
rect 6566 23948 6618 23951
rect 6674 23948 6726 23951
rect 6782 23948 6834 23951
rect 6890 23948 6942 23951
rect 6998 23948 7050 23951
rect 7106 23948 7158 23951
rect 7214 23948 7266 23951
rect 7322 23948 7374 23951
rect 7430 23948 7482 23951
rect 7538 23948 7590 23951
rect 9677 23948 9729 23951
rect 9785 23948 9837 23951
rect 9893 23948 9945 23951
rect 10001 23948 10053 23951
rect 10109 23948 10161 23951
rect 10217 23948 10269 23951
rect 10325 23948 10377 23951
rect 10433 23948 10485 23951
rect 10541 23948 10593 23951
rect 10649 23948 10701 23951
rect 10757 23948 10809 23951
rect 10865 23948 10917 23951
rect 10973 23948 11025 23951
rect 11081 23948 11133 23951
rect 11189 23948 11241 23951
rect 11297 23948 11349 23951
rect 11405 23948 11457 23951
rect 3433 23902 3485 23948
rect 3541 23902 3593 23948
rect 3649 23902 3701 23948
rect 3757 23902 3809 23948
rect 3865 23902 3917 23948
rect 3973 23902 4025 23948
rect 4081 23902 4133 23948
rect 4189 23902 4241 23948
rect 4297 23902 4349 23948
rect 4405 23902 4457 23948
rect 4513 23902 4565 23948
rect 4621 23902 4673 23948
rect 4729 23902 4781 23948
rect 4837 23902 4889 23948
rect 4945 23902 4997 23948
rect 5053 23902 5105 23948
rect 5161 23902 5213 23948
rect 6566 23902 6618 23948
rect 6674 23902 6726 23948
rect 6782 23902 6834 23948
rect 6890 23902 6942 23948
rect 6998 23902 7050 23948
rect 7106 23902 7158 23948
rect 7214 23902 7266 23948
rect 7322 23902 7374 23948
rect 7430 23902 7482 23948
rect 7538 23902 7590 23948
rect 9677 23902 9729 23948
rect 9785 23902 9837 23948
rect 9893 23902 9945 23948
rect 10001 23902 10053 23948
rect 10109 23902 10161 23948
rect 10217 23902 10269 23948
rect 10325 23902 10377 23948
rect 10433 23902 10485 23948
rect 10541 23902 10593 23948
rect 10649 23902 10701 23948
rect 10757 23902 10809 23948
rect 10865 23902 10917 23948
rect 10973 23902 11025 23948
rect 11081 23902 11133 23948
rect 11189 23902 11241 23948
rect 11297 23902 11349 23948
rect 11405 23902 11457 23948
rect 3433 23899 3485 23902
rect 3541 23899 3593 23902
rect 3649 23899 3701 23902
rect 3757 23899 3809 23902
rect 3865 23899 3917 23902
rect 3973 23899 4025 23902
rect 4081 23899 4133 23902
rect 4189 23899 4241 23902
rect 4297 23899 4349 23902
rect 4405 23899 4457 23902
rect 4513 23899 4565 23902
rect 4621 23899 4673 23902
rect 4729 23899 4781 23902
rect 4837 23899 4889 23902
rect 4945 23899 4997 23902
rect 5053 23899 5105 23902
rect 5161 23899 5213 23902
rect 6566 23899 6618 23902
rect 6674 23899 6726 23902
rect 6782 23899 6834 23902
rect 6890 23899 6942 23902
rect 6998 23899 7050 23902
rect 7106 23899 7158 23902
rect 7214 23899 7266 23902
rect 7322 23899 7374 23902
rect 7430 23899 7482 23902
rect 7538 23899 7590 23902
rect 9677 23899 9729 23902
rect 9785 23899 9837 23902
rect 9893 23899 9945 23902
rect 10001 23899 10053 23902
rect 10109 23899 10161 23902
rect 10217 23899 10269 23902
rect 10325 23899 10377 23902
rect 10433 23899 10485 23902
rect 10541 23899 10593 23902
rect 10649 23899 10701 23902
rect 10757 23899 10809 23902
rect 10865 23899 10917 23902
rect 10973 23899 11025 23902
rect 11081 23899 11133 23902
rect 11189 23899 11241 23902
rect 11297 23899 11349 23902
rect 11405 23899 11457 23902
rect 1233 23835 1285 23887
rect 1341 23835 1393 23887
rect 1233 23727 1256 23779
rect 1256 23727 1285 23779
rect 1341 23727 1393 23779
rect 1233 23619 1256 23671
rect 1256 23619 1285 23671
rect 1341 23619 1393 23671
rect 1233 23511 1256 23563
rect 1256 23511 1285 23563
rect 1341 23511 1393 23563
rect 1233 23403 1256 23455
rect 1256 23403 1285 23455
rect 1341 23403 1393 23455
rect 1233 23295 1256 23347
rect 1256 23295 1285 23347
rect 1341 23295 1393 23347
rect 1233 23187 1256 23239
rect 1256 23187 1285 23239
rect 1341 23187 1393 23239
rect 1233 23079 1256 23131
rect 1256 23079 1285 23131
rect 1341 23079 1393 23131
rect 1233 22971 1256 23023
rect 1256 22971 1285 23023
rect 1341 22971 1393 23023
rect 1233 22863 1256 22915
rect 1256 22863 1285 22915
rect 1341 22863 1393 22915
rect 1233 22755 1256 22807
rect 1256 22755 1285 22807
rect 1341 22755 1393 22807
rect 1233 22647 1256 22699
rect 1256 22647 1285 22699
rect 1341 22647 1393 22699
rect 1233 22539 1256 22591
rect 1256 22539 1285 22591
rect 1341 22539 1393 22591
rect 1233 22431 1256 22483
rect 1256 22431 1285 22483
rect 1341 22431 1393 22483
rect 1233 22323 1256 22375
rect 1256 22323 1285 22375
rect 1341 22323 1393 22375
rect 1233 22215 1256 22267
rect 1256 22215 1285 22267
rect 1341 22215 1393 22267
rect 1233 22107 1256 22159
rect 1256 22107 1285 22159
rect 1341 22107 1393 22159
rect 1233 21999 1256 22051
rect 1256 21999 1285 22051
rect 1341 21999 1393 22051
rect 1233 21891 1256 21943
rect 1256 21891 1285 21943
rect 1341 21891 1393 21943
rect 1233 21783 1256 21835
rect 1256 21783 1285 21835
rect 1341 21783 1393 21835
rect 1233 21675 1256 21727
rect 1256 21675 1285 21727
rect 1341 21675 1393 21727
rect 1233 21567 1256 21619
rect 1256 21567 1285 21619
rect 1341 21567 1393 21619
rect 1233 21459 1256 21511
rect 1256 21459 1285 21511
rect 1341 21459 1393 21511
rect 1233 21351 1256 21403
rect 1256 21351 1285 21403
rect 1341 21351 1393 21403
rect 1233 21243 1256 21295
rect 1256 21243 1285 21295
rect 1341 21243 1393 21295
rect 1233 21135 1256 21187
rect 1256 21135 1285 21187
rect 1341 21135 1393 21187
rect 1233 21027 1256 21079
rect 1256 21027 1285 21079
rect 1341 21027 1393 21079
rect 1233 20919 1256 20971
rect 1256 20919 1285 20971
rect 1341 20919 1393 20971
rect 1233 20811 1256 20863
rect 1256 20811 1285 20863
rect 1341 20811 1393 20863
rect 1233 20703 1256 20755
rect 1256 20703 1285 20755
rect 1341 20703 1393 20755
rect 1233 20595 1256 20647
rect 1256 20595 1285 20647
rect 1341 20595 1393 20647
rect 1233 20487 1256 20539
rect 1256 20487 1285 20539
rect 1341 20487 1393 20539
rect 1233 20379 1256 20431
rect 1256 20379 1285 20431
rect 1341 20379 1393 20431
rect 1233 20271 1256 20323
rect 1256 20271 1285 20323
rect 1341 20271 1393 20323
rect 1233 20163 1256 20215
rect 1256 20163 1285 20215
rect 1341 20163 1393 20215
rect 1233 20055 1256 20107
rect 1256 20055 1285 20107
rect 1341 20055 1393 20107
rect 1233 19947 1256 19999
rect 1256 19947 1285 19999
rect 1341 19947 1393 19999
rect 1233 19839 1256 19891
rect 1256 19839 1285 19891
rect 1341 19839 1393 19891
rect 1233 19731 1256 19783
rect 1256 19731 1285 19783
rect 1341 19731 1393 19783
rect 1233 19623 1256 19675
rect 1256 19623 1285 19675
rect 1341 19623 1393 19675
rect 1233 19515 1256 19567
rect 1256 19515 1285 19567
rect 1341 19515 1393 19567
rect 1233 19407 1256 19459
rect 1256 19407 1285 19459
rect 1341 19407 1393 19459
rect 1233 19299 1256 19351
rect 1256 19299 1285 19351
rect 1341 19299 1393 19351
rect 1233 19191 1256 19243
rect 1256 19191 1285 19243
rect 1341 19191 1393 19243
rect 11569 23835 11621 23887
rect 11677 23835 11729 23887
rect 1505 23704 1557 23707
rect 1613 23704 1665 23707
rect 1721 23704 1773 23707
rect 1829 23704 1881 23707
rect 1937 23704 1989 23707
rect 2045 23704 2097 23707
rect 2153 23704 2205 23707
rect 2261 23704 2313 23707
rect 2369 23704 2421 23707
rect 2477 23704 2529 23707
rect 2585 23704 2637 23707
rect 2693 23704 2745 23707
rect 2801 23704 2853 23707
rect 2909 23704 2961 23707
rect 3017 23704 3069 23707
rect 3125 23704 3177 23707
rect 3233 23704 3285 23707
rect 5372 23704 5424 23707
rect 5480 23704 5532 23707
rect 5588 23704 5640 23707
rect 5696 23704 5748 23707
rect 5804 23704 5856 23707
rect 5912 23704 5964 23707
rect 6020 23704 6072 23707
rect 6128 23704 6180 23707
rect 6236 23704 6288 23707
rect 6344 23704 6396 23707
rect 7749 23704 7801 23707
rect 7857 23704 7909 23707
rect 7965 23704 8017 23707
rect 8073 23704 8125 23707
rect 8181 23704 8233 23707
rect 8289 23704 8341 23707
rect 8397 23704 8449 23707
rect 8505 23704 8557 23707
rect 8613 23704 8665 23707
rect 8721 23704 8773 23707
rect 8829 23704 8881 23707
rect 8937 23704 8989 23707
rect 9045 23704 9097 23707
rect 9153 23704 9205 23707
rect 9261 23704 9313 23707
rect 9369 23704 9421 23707
rect 9477 23704 9529 23707
rect 1505 23658 1557 23704
rect 1613 23658 1665 23704
rect 1721 23658 1773 23704
rect 1829 23658 1881 23704
rect 1937 23658 1989 23704
rect 2045 23658 2097 23704
rect 2153 23658 2205 23704
rect 2261 23658 2313 23704
rect 2369 23658 2421 23704
rect 2477 23658 2529 23704
rect 2585 23658 2637 23704
rect 2693 23658 2745 23704
rect 2801 23658 2853 23704
rect 2909 23658 2961 23704
rect 3017 23658 3069 23704
rect 3125 23658 3177 23704
rect 3233 23658 3285 23704
rect 5372 23658 5424 23704
rect 5480 23658 5532 23704
rect 5588 23658 5640 23704
rect 5696 23658 5748 23704
rect 5804 23658 5856 23704
rect 5912 23658 5964 23704
rect 6020 23658 6072 23704
rect 6128 23658 6180 23704
rect 6236 23658 6288 23704
rect 6344 23658 6396 23704
rect 7749 23658 7801 23704
rect 7857 23658 7909 23704
rect 7965 23658 8017 23704
rect 8073 23658 8125 23704
rect 8181 23658 8233 23704
rect 8289 23658 8341 23704
rect 8397 23658 8449 23704
rect 8505 23658 8557 23704
rect 8613 23658 8665 23704
rect 8721 23658 8773 23704
rect 8829 23658 8881 23704
rect 8937 23658 8989 23704
rect 9045 23658 9097 23704
rect 9153 23658 9205 23704
rect 9261 23658 9313 23704
rect 9369 23658 9421 23704
rect 9477 23658 9529 23704
rect 1505 23655 1557 23658
rect 1613 23655 1665 23658
rect 1721 23655 1773 23658
rect 1829 23655 1881 23658
rect 1937 23655 1989 23658
rect 2045 23655 2097 23658
rect 2153 23655 2205 23658
rect 2261 23655 2313 23658
rect 2369 23655 2421 23658
rect 2477 23655 2529 23658
rect 2585 23655 2637 23658
rect 2693 23655 2745 23658
rect 2801 23655 2853 23658
rect 2909 23655 2961 23658
rect 3017 23655 3069 23658
rect 3125 23655 3177 23658
rect 3233 23655 3285 23658
rect 5372 23655 5424 23658
rect 5480 23655 5532 23658
rect 5588 23655 5640 23658
rect 5696 23655 5748 23658
rect 5804 23655 5856 23658
rect 5912 23655 5964 23658
rect 6020 23655 6072 23658
rect 6128 23655 6180 23658
rect 6236 23655 6288 23658
rect 6344 23655 6396 23658
rect 7749 23655 7801 23658
rect 7857 23655 7909 23658
rect 7965 23655 8017 23658
rect 8073 23655 8125 23658
rect 8181 23655 8233 23658
rect 8289 23655 8341 23658
rect 8397 23655 8449 23658
rect 8505 23655 8557 23658
rect 8613 23655 8665 23658
rect 8721 23655 8773 23658
rect 8829 23655 8881 23658
rect 8937 23655 8989 23658
rect 9045 23655 9097 23658
rect 9153 23655 9205 23658
rect 9261 23655 9313 23658
rect 9369 23655 9421 23658
rect 9477 23655 9529 23658
rect 3433 23460 3485 23463
rect 3541 23460 3593 23463
rect 3649 23460 3701 23463
rect 3757 23460 3809 23463
rect 3865 23460 3917 23463
rect 3973 23460 4025 23463
rect 4081 23460 4133 23463
rect 4189 23460 4241 23463
rect 4297 23460 4349 23463
rect 4405 23460 4457 23463
rect 4513 23460 4565 23463
rect 4621 23460 4673 23463
rect 4729 23460 4781 23463
rect 4837 23460 4889 23463
rect 4945 23460 4997 23463
rect 5053 23460 5105 23463
rect 5161 23460 5213 23463
rect 6566 23460 6618 23463
rect 6674 23460 6726 23463
rect 6782 23460 6834 23463
rect 6890 23460 6942 23463
rect 6998 23460 7050 23463
rect 7106 23460 7158 23463
rect 7214 23460 7266 23463
rect 7322 23460 7374 23463
rect 7430 23460 7482 23463
rect 7538 23460 7590 23463
rect 9677 23460 9729 23463
rect 9785 23460 9837 23463
rect 9893 23460 9945 23463
rect 10001 23460 10053 23463
rect 10109 23460 10161 23463
rect 10217 23460 10269 23463
rect 10325 23460 10377 23463
rect 10433 23460 10485 23463
rect 10541 23460 10593 23463
rect 10649 23460 10701 23463
rect 10757 23460 10809 23463
rect 10865 23460 10917 23463
rect 10973 23460 11025 23463
rect 11081 23460 11133 23463
rect 11189 23460 11241 23463
rect 11297 23460 11349 23463
rect 11405 23460 11457 23463
rect 3433 23414 3485 23460
rect 3541 23414 3593 23460
rect 3649 23414 3701 23460
rect 3757 23414 3809 23460
rect 3865 23414 3917 23460
rect 3973 23414 4025 23460
rect 4081 23414 4133 23460
rect 4189 23414 4241 23460
rect 4297 23414 4349 23460
rect 4405 23414 4457 23460
rect 4513 23414 4565 23460
rect 4621 23414 4673 23460
rect 4729 23414 4781 23460
rect 4837 23414 4889 23460
rect 4945 23414 4997 23460
rect 5053 23414 5105 23460
rect 5161 23414 5213 23460
rect 6566 23414 6618 23460
rect 6674 23414 6726 23460
rect 6782 23414 6834 23460
rect 6890 23414 6942 23460
rect 6998 23414 7050 23460
rect 7106 23414 7158 23460
rect 7214 23414 7266 23460
rect 7322 23414 7374 23460
rect 7430 23414 7482 23460
rect 7538 23414 7590 23460
rect 9677 23414 9729 23460
rect 9785 23414 9837 23460
rect 9893 23414 9945 23460
rect 10001 23414 10053 23460
rect 10109 23414 10161 23460
rect 10217 23414 10269 23460
rect 10325 23414 10377 23460
rect 10433 23414 10485 23460
rect 10541 23414 10593 23460
rect 10649 23414 10701 23460
rect 10757 23414 10809 23460
rect 10865 23414 10917 23460
rect 10973 23414 11025 23460
rect 11081 23414 11133 23460
rect 11189 23414 11241 23460
rect 11297 23414 11349 23460
rect 11405 23414 11457 23460
rect 3433 23411 3485 23414
rect 3541 23411 3593 23414
rect 3649 23411 3701 23414
rect 3757 23411 3809 23414
rect 3865 23411 3917 23414
rect 3973 23411 4025 23414
rect 4081 23411 4133 23414
rect 4189 23411 4241 23414
rect 4297 23411 4349 23414
rect 4405 23411 4457 23414
rect 4513 23411 4565 23414
rect 4621 23411 4673 23414
rect 4729 23411 4781 23414
rect 4837 23411 4889 23414
rect 4945 23411 4997 23414
rect 5053 23411 5105 23414
rect 5161 23411 5213 23414
rect 6566 23411 6618 23414
rect 6674 23411 6726 23414
rect 6782 23411 6834 23414
rect 6890 23411 6942 23414
rect 6998 23411 7050 23414
rect 7106 23411 7158 23414
rect 7214 23411 7266 23414
rect 7322 23411 7374 23414
rect 7430 23411 7482 23414
rect 7538 23411 7590 23414
rect 9677 23411 9729 23414
rect 9785 23411 9837 23414
rect 9893 23411 9945 23414
rect 10001 23411 10053 23414
rect 10109 23411 10161 23414
rect 10217 23411 10269 23414
rect 10325 23411 10377 23414
rect 10433 23411 10485 23414
rect 10541 23411 10593 23414
rect 10649 23411 10701 23414
rect 10757 23411 10809 23414
rect 10865 23411 10917 23414
rect 10973 23411 11025 23414
rect 11081 23411 11133 23414
rect 11189 23411 11241 23414
rect 11297 23411 11349 23414
rect 11405 23411 11457 23414
rect 1505 23216 1557 23219
rect 1613 23216 1665 23219
rect 1721 23216 1773 23219
rect 1829 23216 1881 23219
rect 1937 23216 1989 23219
rect 2045 23216 2097 23219
rect 2153 23216 2205 23219
rect 2261 23216 2313 23219
rect 2369 23216 2421 23219
rect 2477 23216 2529 23219
rect 2585 23216 2637 23219
rect 2693 23216 2745 23219
rect 2801 23216 2853 23219
rect 2909 23216 2961 23219
rect 3017 23216 3069 23219
rect 3125 23216 3177 23219
rect 3233 23216 3285 23219
rect 5372 23216 5424 23219
rect 5480 23216 5532 23219
rect 5588 23216 5640 23219
rect 5696 23216 5748 23219
rect 5804 23216 5856 23219
rect 5912 23216 5964 23219
rect 6020 23216 6072 23219
rect 6128 23216 6180 23219
rect 6236 23216 6288 23219
rect 6344 23216 6396 23219
rect 7749 23216 7801 23219
rect 7857 23216 7909 23219
rect 7965 23216 8017 23219
rect 8073 23216 8125 23219
rect 8181 23216 8233 23219
rect 8289 23216 8341 23219
rect 8397 23216 8449 23219
rect 8505 23216 8557 23219
rect 8613 23216 8665 23219
rect 8721 23216 8773 23219
rect 8829 23216 8881 23219
rect 8937 23216 8989 23219
rect 9045 23216 9097 23219
rect 9153 23216 9205 23219
rect 9261 23216 9313 23219
rect 9369 23216 9421 23219
rect 9477 23216 9529 23219
rect 1505 23170 1557 23216
rect 1613 23170 1665 23216
rect 1721 23170 1773 23216
rect 1829 23170 1881 23216
rect 1937 23170 1989 23216
rect 2045 23170 2097 23216
rect 2153 23170 2205 23216
rect 2261 23170 2313 23216
rect 2369 23170 2421 23216
rect 2477 23170 2529 23216
rect 2585 23170 2637 23216
rect 2693 23170 2745 23216
rect 2801 23170 2853 23216
rect 2909 23170 2961 23216
rect 3017 23170 3069 23216
rect 3125 23170 3177 23216
rect 3233 23170 3285 23216
rect 5372 23170 5424 23216
rect 5480 23170 5532 23216
rect 5588 23170 5640 23216
rect 5696 23170 5748 23216
rect 5804 23170 5856 23216
rect 5912 23170 5964 23216
rect 6020 23170 6072 23216
rect 6128 23170 6180 23216
rect 6236 23170 6288 23216
rect 6344 23170 6396 23216
rect 7749 23170 7801 23216
rect 7857 23170 7909 23216
rect 7965 23170 8017 23216
rect 8073 23170 8125 23216
rect 8181 23170 8233 23216
rect 8289 23170 8341 23216
rect 8397 23170 8449 23216
rect 8505 23170 8557 23216
rect 8613 23170 8665 23216
rect 8721 23170 8773 23216
rect 8829 23170 8881 23216
rect 8937 23170 8989 23216
rect 9045 23170 9097 23216
rect 9153 23170 9205 23216
rect 9261 23170 9313 23216
rect 9369 23170 9421 23216
rect 9477 23170 9529 23216
rect 1505 23167 1557 23170
rect 1613 23167 1665 23170
rect 1721 23167 1773 23170
rect 1829 23167 1881 23170
rect 1937 23167 1989 23170
rect 2045 23167 2097 23170
rect 2153 23167 2205 23170
rect 2261 23167 2313 23170
rect 2369 23167 2421 23170
rect 2477 23167 2529 23170
rect 2585 23167 2637 23170
rect 2693 23167 2745 23170
rect 2801 23167 2853 23170
rect 2909 23167 2961 23170
rect 3017 23167 3069 23170
rect 3125 23167 3177 23170
rect 3233 23167 3285 23170
rect 5372 23167 5424 23170
rect 5480 23167 5532 23170
rect 5588 23167 5640 23170
rect 5696 23167 5748 23170
rect 5804 23167 5856 23170
rect 5912 23167 5964 23170
rect 6020 23167 6072 23170
rect 6128 23167 6180 23170
rect 6236 23167 6288 23170
rect 6344 23167 6396 23170
rect 7749 23167 7801 23170
rect 7857 23167 7909 23170
rect 7965 23167 8017 23170
rect 8073 23167 8125 23170
rect 8181 23167 8233 23170
rect 8289 23167 8341 23170
rect 8397 23167 8449 23170
rect 8505 23167 8557 23170
rect 8613 23167 8665 23170
rect 8721 23167 8773 23170
rect 8829 23167 8881 23170
rect 8937 23167 8989 23170
rect 9045 23167 9097 23170
rect 9153 23167 9205 23170
rect 9261 23167 9313 23170
rect 9369 23167 9421 23170
rect 9477 23167 9529 23170
rect 3433 22972 3485 22975
rect 3541 22972 3593 22975
rect 3649 22972 3701 22975
rect 3757 22972 3809 22975
rect 3865 22972 3917 22975
rect 3973 22972 4025 22975
rect 4081 22972 4133 22975
rect 4189 22972 4241 22975
rect 4297 22972 4349 22975
rect 4405 22972 4457 22975
rect 4513 22972 4565 22975
rect 4621 22972 4673 22975
rect 4729 22972 4781 22975
rect 4837 22972 4889 22975
rect 4945 22972 4997 22975
rect 5053 22972 5105 22975
rect 5161 22972 5213 22975
rect 6566 22972 6618 22975
rect 6674 22972 6726 22975
rect 6782 22972 6834 22975
rect 6890 22972 6942 22975
rect 6998 22972 7050 22975
rect 7106 22972 7158 22975
rect 7214 22972 7266 22975
rect 7322 22972 7374 22975
rect 7430 22972 7482 22975
rect 7538 22972 7590 22975
rect 9677 22972 9729 22975
rect 9785 22972 9837 22975
rect 9893 22972 9945 22975
rect 10001 22972 10053 22975
rect 10109 22972 10161 22975
rect 10217 22972 10269 22975
rect 10325 22972 10377 22975
rect 10433 22972 10485 22975
rect 10541 22972 10593 22975
rect 10649 22972 10701 22975
rect 10757 22972 10809 22975
rect 10865 22972 10917 22975
rect 10973 22972 11025 22975
rect 11081 22972 11133 22975
rect 11189 22972 11241 22975
rect 11297 22972 11349 22975
rect 11405 22972 11457 22975
rect 3433 22926 3485 22972
rect 3541 22926 3593 22972
rect 3649 22926 3701 22972
rect 3757 22926 3809 22972
rect 3865 22926 3917 22972
rect 3973 22926 4025 22972
rect 4081 22926 4133 22972
rect 4189 22926 4241 22972
rect 4297 22926 4349 22972
rect 4405 22926 4457 22972
rect 4513 22926 4565 22972
rect 4621 22926 4673 22972
rect 4729 22926 4781 22972
rect 4837 22926 4889 22972
rect 4945 22926 4997 22972
rect 5053 22926 5105 22972
rect 5161 22926 5213 22972
rect 6566 22926 6618 22972
rect 6674 22926 6726 22972
rect 6782 22926 6834 22972
rect 6890 22926 6942 22972
rect 6998 22926 7050 22972
rect 7106 22926 7158 22972
rect 7214 22926 7266 22972
rect 7322 22926 7374 22972
rect 7430 22926 7482 22972
rect 7538 22926 7590 22972
rect 9677 22926 9729 22972
rect 9785 22926 9837 22972
rect 9893 22926 9945 22972
rect 10001 22926 10053 22972
rect 10109 22926 10161 22972
rect 10217 22926 10269 22972
rect 10325 22926 10377 22972
rect 10433 22926 10485 22972
rect 10541 22926 10593 22972
rect 10649 22926 10701 22972
rect 10757 22926 10809 22972
rect 10865 22926 10917 22972
rect 10973 22926 11025 22972
rect 11081 22926 11133 22972
rect 11189 22926 11241 22972
rect 11297 22926 11349 22972
rect 11405 22926 11457 22972
rect 3433 22923 3485 22926
rect 3541 22923 3593 22926
rect 3649 22923 3701 22926
rect 3757 22923 3809 22926
rect 3865 22923 3917 22926
rect 3973 22923 4025 22926
rect 4081 22923 4133 22926
rect 4189 22923 4241 22926
rect 4297 22923 4349 22926
rect 4405 22923 4457 22926
rect 4513 22923 4565 22926
rect 4621 22923 4673 22926
rect 4729 22923 4781 22926
rect 4837 22923 4889 22926
rect 4945 22923 4997 22926
rect 5053 22923 5105 22926
rect 5161 22923 5213 22926
rect 6566 22923 6618 22926
rect 6674 22923 6726 22926
rect 6782 22923 6834 22926
rect 6890 22923 6942 22926
rect 6998 22923 7050 22926
rect 7106 22923 7158 22926
rect 7214 22923 7266 22926
rect 7322 22923 7374 22926
rect 7430 22923 7482 22926
rect 7538 22923 7590 22926
rect 9677 22923 9729 22926
rect 9785 22923 9837 22926
rect 9893 22923 9945 22926
rect 10001 22923 10053 22926
rect 10109 22923 10161 22926
rect 10217 22923 10269 22926
rect 10325 22923 10377 22926
rect 10433 22923 10485 22926
rect 10541 22923 10593 22926
rect 10649 22923 10701 22926
rect 10757 22923 10809 22926
rect 10865 22923 10917 22926
rect 10973 22923 11025 22926
rect 11081 22923 11133 22926
rect 11189 22923 11241 22926
rect 11297 22923 11349 22926
rect 11405 22923 11457 22926
rect 1505 22728 1557 22731
rect 1613 22728 1665 22731
rect 1721 22728 1773 22731
rect 1829 22728 1881 22731
rect 1937 22728 1989 22731
rect 2045 22728 2097 22731
rect 2153 22728 2205 22731
rect 2261 22728 2313 22731
rect 2369 22728 2421 22731
rect 2477 22728 2529 22731
rect 2585 22728 2637 22731
rect 2693 22728 2745 22731
rect 2801 22728 2853 22731
rect 2909 22728 2961 22731
rect 3017 22728 3069 22731
rect 3125 22728 3177 22731
rect 3233 22728 3285 22731
rect 5372 22728 5424 22731
rect 5480 22728 5532 22731
rect 5588 22728 5640 22731
rect 5696 22728 5748 22731
rect 5804 22728 5856 22731
rect 5912 22728 5964 22731
rect 6020 22728 6072 22731
rect 6128 22728 6180 22731
rect 6236 22728 6288 22731
rect 6344 22728 6396 22731
rect 7749 22728 7801 22731
rect 7857 22728 7909 22731
rect 7965 22728 8017 22731
rect 8073 22728 8125 22731
rect 8181 22728 8233 22731
rect 8289 22728 8341 22731
rect 8397 22728 8449 22731
rect 8505 22728 8557 22731
rect 8613 22728 8665 22731
rect 8721 22728 8773 22731
rect 8829 22728 8881 22731
rect 8937 22728 8989 22731
rect 9045 22728 9097 22731
rect 9153 22728 9205 22731
rect 9261 22728 9313 22731
rect 9369 22728 9421 22731
rect 9477 22728 9529 22731
rect 1505 22682 1557 22728
rect 1613 22682 1665 22728
rect 1721 22682 1773 22728
rect 1829 22682 1881 22728
rect 1937 22682 1989 22728
rect 2045 22682 2097 22728
rect 2153 22682 2205 22728
rect 2261 22682 2313 22728
rect 2369 22682 2421 22728
rect 2477 22682 2529 22728
rect 2585 22682 2637 22728
rect 2693 22682 2745 22728
rect 2801 22682 2853 22728
rect 2909 22682 2961 22728
rect 3017 22682 3069 22728
rect 3125 22682 3177 22728
rect 3233 22682 3285 22728
rect 5372 22682 5424 22728
rect 5480 22682 5532 22728
rect 5588 22682 5640 22728
rect 5696 22682 5748 22728
rect 5804 22682 5856 22728
rect 5912 22682 5964 22728
rect 6020 22682 6072 22728
rect 6128 22682 6180 22728
rect 6236 22682 6288 22728
rect 6344 22682 6396 22728
rect 7749 22682 7801 22728
rect 7857 22682 7909 22728
rect 7965 22682 8017 22728
rect 8073 22682 8125 22728
rect 8181 22682 8233 22728
rect 8289 22682 8341 22728
rect 8397 22682 8449 22728
rect 8505 22682 8557 22728
rect 8613 22682 8665 22728
rect 8721 22682 8773 22728
rect 8829 22682 8881 22728
rect 8937 22682 8989 22728
rect 9045 22682 9097 22728
rect 9153 22682 9205 22728
rect 9261 22682 9313 22728
rect 9369 22682 9421 22728
rect 9477 22682 9529 22728
rect 1505 22679 1557 22682
rect 1613 22679 1665 22682
rect 1721 22679 1773 22682
rect 1829 22679 1881 22682
rect 1937 22679 1989 22682
rect 2045 22679 2097 22682
rect 2153 22679 2205 22682
rect 2261 22679 2313 22682
rect 2369 22679 2421 22682
rect 2477 22679 2529 22682
rect 2585 22679 2637 22682
rect 2693 22679 2745 22682
rect 2801 22679 2853 22682
rect 2909 22679 2961 22682
rect 3017 22679 3069 22682
rect 3125 22679 3177 22682
rect 3233 22679 3285 22682
rect 5372 22679 5424 22682
rect 5480 22679 5532 22682
rect 5588 22679 5640 22682
rect 5696 22679 5748 22682
rect 5804 22679 5856 22682
rect 5912 22679 5964 22682
rect 6020 22679 6072 22682
rect 6128 22679 6180 22682
rect 6236 22679 6288 22682
rect 6344 22679 6396 22682
rect 7749 22679 7801 22682
rect 7857 22679 7909 22682
rect 7965 22679 8017 22682
rect 8073 22679 8125 22682
rect 8181 22679 8233 22682
rect 8289 22679 8341 22682
rect 8397 22679 8449 22682
rect 8505 22679 8557 22682
rect 8613 22679 8665 22682
rect 8721 22679 8773 22682
rect 8829 22679 8881 22682
rect 8937 22679 8989 22682
rect 9045 22679 9097 22682
rect 9153 22679 9205 22682
rect 9261 22679 9313 22682
rect 9369 22679 9421 22682
rect 9477 22679 9529 22682
rect 3433 22484 3485 22487
rect 3541 22484 3593 22487
rect 3649 22484 3701 22487
rect 3757 22484 3809 22487
rect 3865 22484 3917 22487
rect 3973 22484 4025 22487
rect 4081 22484 4133 22487
rect 4189 22484 4241 22487
rect 4297 22484 4349 22487
rect 4405 22484 4457 22487
rect 4513 22484 4565 22487
rect 4621 22484 4673 22487
rect 4729 22484 4781 22487
rect 4837 22484 4889 22487
rect 4945 22484 4997 22487
rect 5053 22484 5105 22487
rect 5161 22484 5213 22487
rect 6566 22484 6618 22487
rect 6674 22484 6726 22487
rect 6782 22484 6834 22487
rect 6890 22484 6942 22487
rect 6998 22484 7050 22487
rect 7106 22484 7158 22487
rect 7214 22484 7266 22487
rect 7322 22484 7374 22487
rect 7430 22484 7482 22487
rect 7538 22484 7590 22487
rect 9677 22484 9729 22487
rect 9785 22484 9837 22487
rect 9893 22484 9945 22487
rect 10001 22484 10053 22487
rect 10109 22484 10161 22487
rect 10217 22484 10269 22487
rect 10325 22484 10377 22487
rect 10433 22484 10485 22487
rect 10541 22484 10593 22487
rect 10649 22484 10701 22487
rect 10757 22484 10809 22487
rect 10865 22484 10917 22487
rect 10973 22484 11025 22487
rect 11081 22484 11133 22487
rect 11189 22484 11241 22487
rect 11297 22484 11349 22487
rect 11405 22484 11457 22487
rect 3433 22438 3485 22484
rect 3541 22438 3593 22484
rect 3649 22438 3701 22484
rect 3757 22438 3809 22484
rect 3865 22438 3917 22484
rect 3973 22438 4025 22484
rect 4081 22438 4133 22484
rect 4189 22438 4241 22484
rect 4297 22438 4349 22484
rect 4405 22438 4457 22484
rect 4513 22438 4565 22484
rect 4621 22438 4673 22484
rect 4729 22438 4781 22484
rect 4837 22438 4889 22484
rect 4945 22438 4997 22484
rect 5053 22438 5105 22484
rect 5161 22438 5213 22484
rect 6566 22438 6618 22484
rect 6674 22438 6726 22484
rect 6782 22438 6834 22484
rect 6890 22438 6942 22484
rect 6998 22438 7050 22484
rect 7106 22438 7158 22484
rect 7214 22438 7266 22484
rect 7322 22438 7374 22484
rect 7430 22438 7482 22484
rect 7538 22438 7590 22484
rect 9677 22438 9729 22484
rect 9785 22438 9837 22484
rect 9893 22438 9945 22484
rect 10001 22438 10053 22484
rect 10109 22438 10161 22484
rect 10217 22438 10269 22484
rect 10325 22438 10377 22484
rect 10433 22438 10485 22484
rect 10541 22438 10593 22484
rect 10649 22438 10701 22484
rect 10757 22438 10809 22484
rect 10865 22438 10917 22484
rect 10973 22438 11025 22484
rect 11081 22438 11133 22484
rect 11189 22438 11241 22484
rect 11297 22438 11349 22484
rect 11405 22438 11457 22484
rect 3433 22435 3485 22438
rect 3541 22435 3593 22438
rect 3649 22435 3701 22438
rect 3757 22435 3809 22438
rect 3865 22435 3917 22438
rect 3973 22435 4025 22438
rect 4081 22435 4133 22438
rect 4189 22435 4241 22438
rect 4297 22435 4349 22438
rect 4405 22435 4457 22438
rect 4513 22435 4565 22438
rect 4621 22435 4673 22438
rect 4729 22435 4781 22438
rect 4837 22435 4889 22438
rect 4945 22435 4997 22438
rect 5053 22435 5105 22438
rect 5161 22435 5213 22438
rect 6566 22435 6618 22438
rect 6674 22435 6726 22438
rect 6782 22435 6834 22438
rect 6890 22435 6942 22438
rect 6998 22435 7050 22438
rect 7106 22435 7158 22438
rect 7214 22435 7266 22438
rect 7322 22435 7374 22438
rect 7430 22435 7482 22438
rect 7538 22435 7590 22438
rect 9677 22435 9729 22438
rect 9785 22435 9837 22438
rect 9893 22435 9945 22438
rect 10001 22435 10053 22438
rect 10109 22435 10161 22438
rect 10217 22435 10269 22438
rect 10325 22435 10377 22438
rect 10433 22435 10485 22438
rect 10541 22435 10593 22438
rect 10649 22435 10701 22438
rect 10757 22435 10809 22438
rect 10865 22435 10917 22438
rect 10973 22435 11025 22438
rect 11081 22435 11133 22438
rect 11189 22435 11241 22438
rect 11297 22435 11349 22438
rect 11405 22435 11457 22438
rect 1505 22240 1557 22243
rect 1613 22240 1665 22243
rect 1721 22240 1773 22243
rect 1829 22240 1881 22243
rect 1937 22240 1989 22243
rect 2045 22240 2097 22243
rect 2153 22240 2205 22243
rect 2261 22240 2313 22243
rect 2369 22240 2421 22243
rect 2477 22240 2529 22243
rect 2585 22240 2637 22243
rect 2693 22240 2745 22243
rect 2801 22240 2853 22243
rect 2909 22240 2961 22243
rect 3017 22240 3069 22243
rect 3125 22240 3177 22243
rect 3233 22240 3285 22243
rect 5372 22240 5424 22243
rect 5480 22240 5532 22243
rect 5588 22240 5640 22243
rect 5696 22240 5748 22243
rect 5804 22240 5856 22243
rect 5912 22240 5964 22243
rect 6020 22240 6072 22243
rect 6128 22240 6180 22243
rect 6236 22240 6288 22243
rect 6344 22240 6396 22243
rect 7749 22240 7801 22243
rect 7857 22240 7909 22243
rect 7965 22240 8017 22243
rect 8073 22240 8125 22243
rect 8181 22240 8233 22243
rect 8289 22240 8341 22243
rect 8397 22240 8449 22243
rect 8505 22240 8557 22243
rect 8613 22240 8665 22243
rect 8721 22240 8773 22243
rect 8829 22240 8881 22243
rect 8937 22240 8989 22243
rect 9045 22240 9097 22243
rect 9153 22240 9205 22243
rect 9261 22240 9313 22243
rect 9369 22240 9421 22243
rect 9477 22240 9529 22243
rect 1505 22194 1557 22240
rect 1613 22194 1665 22240
rect 1721 22194 1773 22240
rect 1829 22194 1881 22240
rect 1937 22194 1989 22240
rect 2045 22194 2097 22240
rect 2153 22194 2205 22240
rect 2261 22194 2313 22240
rect 2369 22194 2421 22240
rect 2477 22194 2529 22240
rect 2585 22194 2637 22240
rect 2693 22194 2745 22240
rect 2801 22194 2853 22240
rect 2909 22194 2961 22240
rect 3017 22194 3069 22240
rect 3125 22194 3177 22240
rect 3233 22194 3285 22240
rect 5372 22194 5424 22240
rect 5480 22194 5532 22240
rect 5588 22194 5640 22240
rect 5696 22194 5748 22240
rect 5804 22194 5856 22240
rect 5912 22194 5964 22240
rect 6020 22194 6072 22240
rect 6128 22194 6180 22240
rect 6236 22194 6288 22240
rect 6344 22194 6396 22240
rect 7749 22194 7801 22240
rect 7857 22194 7909 22240
rect 7965 22194 8017 22240
rect 8073 22194 8125 22240
rect 8181 22194 8233 22240
rect 8289 22194 8341 22240
rect 8397 22194 8449 22240
rect 8505 22194 8557 22240
rect 8613 22194 8665 22240
rect 8721 22194 8773 22240
rect 8829 22194 8881 22240
rect 8937 22194 8989 22240
rect 9045 22194 9097 22240
rect 9153 22194 9205 22240
rect 9261 22194 9313 22240
rect 9369 22194 9421 22240
rect 9477 22194 9529 22240
rect 1505 22191 1557 22194
rect 1613 22191 1665 22194
rect 1721 22191 1773 22194
rect 1829 22191 1881 22194
rect 1937 22191 1989 22194
rect 2045 22191 2097 22194
rect 2153 22191 2205 22194
rect 2261 22191 2313 22194
rect 2369 22191 2421 22194
rect 2477 22191 2529 22194
rect 2585 22191 2637 22194
rect 2693 22191 2745 22194
rect 2801 22191 2853 22194
rect 2909 22191 2961 22194
rect 3017 22191 3069 22194
rect 3125 22191 3177 22194
rect 3233 22191 3285 22194
rect 5372 22191 5424 22194
rect 5480 22191 5532 22194
rect 5588 22191 5640 22194
rect 5696 22191 5748 22194
rect 5804 22191 5856 22194
rect 5912 22191 5964 22194
rect 6020 22191 6072 22194
rect 6128 22191 6180 22194
rect 6236 22191 6288 22194
rect 6344 22191 6396 22194
rect 7749 22191 7801 22194
rect 7857 22191 7909 22194
rect 7965 22191 8017 22194
rect 8073 22191 8125 22194
rect 8181 22191 8233 22194
rect 8289 22191 8341 22194
rect 8397 22191 8449 22194
rect 8505 22191 8557 22194
rect 8613 22191 8665 22194
rect 8721 22191 8773 22194
rect 8829 22191 8881 22194
rect 8937 22191 8989 22194
rect 9045 22191 9097 22194
rect 9153 22191 9205 22194
rect 9261 22191 9313 22194
rect 9369 22191 9421 22194
rect 9477 22191 9529 22194
rect 3433 21996 3485 21999
rect 3541 21996 3593 21999
rect 3649 21996 3701 21999
rect 3757 21996 3809 21999
rect 3865 21996 3917 21999
rect 3973 21996 4025 21999
rect 4081 21996 4133 21999
rect 4189 21996 4241 21999
rect 4297 21996 4349 21999
rect 4405 21996 4457 21999
rect 4513 21996 4565 21999
rect 4621 21996 4673 21999
rect 4729 21996 4781 21999
rect 4837 21996 4889 21999
rect 4945 21996 4997 21999
rect 5053 21996 5105 21999
rect 5161 21996 5213 21999
rect 6566 21996 6618 21999
rect 6674 21996 6726 21999
rect 6782 21996 6834 21999
rect 6890 21996 6942 21999
rect 6998 21996 7050 21999
rect 7106 21996 7158 21999
rect 7214 21996 7266 21999
rect 7322 21996 7374 21999
rect 7430 21996 7482 21999
rect 7538 21996 7590 21999
rect 9677 21996 9729 21999
rect 9785 21996 9837 21999
rect 9893 21996 9945 21999
rect 10001 21996 10053 21999
rect 10109 21996 10161 21999
rect 10217 21996 10269 21999
rect 10325 21996 10377 21999
rect 10433 21996 10485 21999
rect 10541 21996 10593 21999
rect 10649 21996 10701 21999
rect 10757 21996 10809 21999
rect 10865 21996 10917 21999
rect 10973 21996 11025 21999
rect 11081 21996 11133 21999
rect 11189 21996 11241 21999
rect 11297 21996 11349 21999
rect 11405 21996 11457 21999
rect 3433 21950 3485 21996
rect 3541 21950 3593 21996
rect 3649 21950 3701 21996
rect 3757 21950 3809 21996
rect 3865 21950 3917 21996
rect 3973 21950 4025 21996
rect 4081 21950 4133 21996
rect 4189 21950 4241 21996
rect 4297 21950 4349 21996
rect 4405 21950 4457 21996
rect 4513 21950 4565 21996
rect 4621 21950 4673 21996
rect 4729 21950 4781 21996
rect 4837 21950 4889 21996
rect 4945 21950 4997 21996
rect 5053 21950 5105 21996
rect 5161 21950 5213 21996
rect 6566 21950 6618 21996
rect 6674 21950 6726 21996
rect 6782 21950 6834 21996
rect 6890 21950 6942 21996
rect 6998 21950 7050 21996
rect 7106 21950 7158 21996
rect 7214 21950 7266 21996
rect 7322 21950 7374 21996
rect 7430 21950 7482 21996
rect 7538 21950 7590 21996
rect 9677 21950 9729 21996
rect 9785 21950 9837 21996
rect 9893 21950 9945 21996
rect 10001 21950 10053 21996
rect 10109 21950 10161 21996
rect 10217 21950 10269 21996
rect 10325 21950 10377 21996
rect 10433 21950 10485 21996
rect 10541 21950 10593 21996
rect 10649 21950 10701 21996
rect 10757 21950 10809 21996
rect 10865 21950 10917 21996
rect 10973 21950 11025 21996
rect 11081 21950 11133 21996
rect 11189 21950 11241 21996
rect 11297 21950 11349 21996
rect 11405 21950 11457 21996
rect 3433 21947 3485 21950
rect 3541 21947 3593 21950
rect 3649 21947 3701 21950
rect 3757 21947 3809 21950
rect 3865 21947 3917 21950
rect 3973 21947 4025 21950
rect 4081 21947 4133 21950
rect 4189 21947 4241 21950
rect 4297 21947 4349 21950
rect 4405 21947 4457 21950
rect 4513 21947 4565 21950
rect 4621 21947 4673 21950
rect 4729 21947 4781 21950
rect 4837 21947 4889 21950
rect 4945 21947 4997 21950
rect 5053 21947 5105 21950
rect 5161 21947 5213 21950
rect 6566 21947 6618 21950
rect 6674 21947 6726 21950
rect 6782 21947 6834 21950
rect 6890 21947 6942 21950
rect 6998 21947 7050 21950
rect 7106 21947 7158 21950
rect 7214 21947 7266 21950
rect 7322 21947 7374 21950
rect 7430 21947 7482 21950
rect 7538 21947 7590 21950
rect 9677 21947 9729 21950
rect 9785 21947 9837 21950
rect 9893 21947 9945 21950
rect 10001 21947 10053 21950
rect 10109 21947 10161 21950
rect 10217 21947 10269 21950
rect 10325 21947 10377 21950
rect 10433 21947 10485 21950
rect 10541 21947 10593 21950
rect 10649 21947 10701 21950
rect 10757 21947 10809 21950
rect 10865 21947 10917 21950
rect 10973 21947 11025 21950
rect 11081 21947 11133 21950
rect 11189 21947 11241 21950
rect 11297 21947 11349 21950
rect 11405 21947 11457 21950
rect 1505 21752 1557 21755
rect 1613 21752 1665 21755
rect 1721 21752 1773 21755
rect 1829 21752 1881 21755
rect 1937 21752 1989 21755
rect 2045 21752 2097 21755
rect 2153 21752 2205 21755
rect 2261 21752 2313 21755
rect 2369 21752 2421 21755
rect 2477 21752 2529 21755
rect 2585 21752 2637 21755
rect 2693 21752 2745 21755
rect 2801 21752 2853 21755
rect 2909 21752 2961 21755
rect 3017 21752 3069 21755
rect 3125 21752 3177 21755
rect 3233 21752 3285 21755
rect 5372 21752 5424 21755
rect 5480 21752 5532 21755
rect 5588 21752 5640 21755
rect 5696 21752 5748 21755
rect 5804 21752 5856 21755
rect 5912 21752 5964 21755
rect 6020 21752 6072 21755
rect 6128 21752 6180 21755
rect 6236 21752 6288 21755
rect 6344 21752 6396 21755
rect 7749 21752 7801 21755
rect 7857 21752 7909 21755
rect 7965 21752 8017 21755
rect 8073 21752 8125 21755
rect 8181 21752 8233 21755
rect 8289 21752 8341 21755
rect 8397 21752 8449 21755
rect 8505 21752 8557 21755
rect 8613 21752 8665 21755
rect 8721 21752 8773 21755
rect 8829 21752 8881 21755
rect 8937 21752 8989 21755
rect 9045 21752 9097 21755
rect 9153 21752 9205 21755
rect 9261 21752 9313 21755
rect 9369 21752 9421 21755
rect 9477 21752 9529 21755
rect 1505 21706 1557 21752
rect 1613 21706 1665 21752
rect 1721 21706 1773 21752
rect 1829 21706 1881 21752
rect 1937 21706 1989 21752
rect 2045 21706 2097 21752
rect 2153 21706 2205 21752
rect 2261 21706 2313 21752
rect 2369 21706 2421 21752
rect 2477 21706 2529 21752
rect 2585 21706 2637 21752
rect 2693 21706 2745 21752
rect 2801 21706 2853 21752
rect 2909 21706 2961 21752
rect 3017 21706 3069 21752
rect 3125 21706 3177 21752
rect 3233 21706 3285 21752
rect 5372 21706 5424 21752
rect 5480 21706 5532 21752
rect 5588 21706 5640 21752
rect 5696 21706 5748 21752
rect 5804 21706 5856 21752
rect 5912 21706 5964 21752
rect 6020 21706 6072 21752
rect 6128 21706 6180 21752
rect 6236 21706 6288 21752
rect 6344 21706 6396 21752
rect 7749 21706 7801 21752
rect 7857 21706 7909 21752
rect 7965 21706 8017 21752
rect 8073 21706 8125 21752
rect 8181 21706 8233 21752
rect 8289 21706 8341 21752
rect 8397 21706 8449 21752
rect 8505 21706 8557 21752
rect 8613 21706 8665 21752
rect 8721 21706 8773 21752
rect 8829 21706 8881 21752
rect 8937 21706 8989 21752
rect 9045 21706 9097 21752
rect 9153 21706 9205 21752
rect 9261 21706 9313 21752
rect 9369 21706 9421 21752
rect 9477 21706 9529 21752
rect 1505 21703 1557 21706
rect 1613 21703 1665 21706
rect 1721 21703 1773 21706
rect 1829 21703 1881 21706
rect 1937 21703 1989 21706
rect 2045 21703 2097 21706
rect 2153 21703 2205 21706
rect 2261 21703 2313 21706
rect 2369 21703 2421 21706
rect 2477 21703 2529 21706
rect 2585 21703 2637 21706
rect 2693 21703 2745 21706
rect 2801 21703 2853 21706
rect 2909 21703 2961 21706
rect 3017 21703 3069 21706
rect 3125 21703 3177 21706
rect 3233 21703 3285 21706
rect 5372 21703 5424 21706
rect 5480 21703 5532 21706
rect 5588 21703 5640 21706
rect 5696 21703 5748 21706
rect 5804 21703 5856 21706
rect 5912 21703 5964 21706
rect 6020 21703 6072 21706
rect 6128 21703 6180 21706
rect 6236 21703 6288 21706
rect 6344 21703 6396 21706
rect 7749 21703 7801 21706
rect 7857 21703 7909 21706
rect 7965 21703 8017 21706
rect 8073 21703 8125 21706
rect 8181 21703 8233 21706
rect 8289 21703 8341 21706
rect 8397 21703 8449 21706
rect 8505 21703 8557 21706
rect 8613 21703 8665 21706
rect 8721 21703 8773 21706
rect 8829 21703 8881 21706
rect 8937 21703 8989 21706
rect 9045 21703 9097 21706
rect 9153 21703 9205 21706
rect 9261 21703 9313 21706
rect 9369 21703 9421 21706
rect 9477 21703 9529 21706
rect 3433 21508 3485 21511
rect 3541 21508 3593 21511
rect 3649 21508 3701 21511
rect 3757 21508 3809 21511
rect 3865 21508 3917 21511
rect 3973 21508 4025 21511
rect 4081 21508 4133 21511
rect 4189 21508 4241 21511
rect 4297 21508 4349 21511
rect 4405 21508 4457 21511
rect 4513 21508 4565 21511
rect 4621 21508 4673 21511
rect 4729 21508 4781 21511
rect 4837 21508 4889 21511
rect 4945 21508 4997 21511
rect 5053 21508 5105 21511
rect 5161 21508 5213 21511
rect 6566 21508 6618 21511
rect 6674 21508 6726 21511
rect 6782 21508 6834 21511
rect 6890 21508 6942 21511
rect 6998 21508 7050 21511
rect 7106 21508 7158 21511
rect 7214 21508 7266 21511
rect 7322 21508 7374 21511
rect 7430 21508 7482 21511
rect 7538 21508 7590 21511
rect 9677 21508 9729 21511
rect 9785 21508 9837 21511
rect 9893 21508 9945 21511
rect 10001 21508 10053 21511
rect 10109 21508 10161 21511
rect 10217 21508 10269 21511
rect 10325 21508 10377 21511
rect 10433 21508 10485 21511
rect 10541 21508 10593 21511
rect 10649 21508 10701 21511
rect 10757 21508 10809 21511
rect 10865 21508 10917 21511
rect 10973 21508 11025 21511
rect 11081 21508 11133 21511
rect 11189 21508 11241 21511
rect 11297 21508 11349 21511
rect 11405 21508 11457 21511
rect 3433 21462 3485 21508
rect 3541 21462 3593 21508
rect 3649 21462 3701 21508
rect 3757 21462 3809 21508
rect 3865 21462 3917 21508
rect 3973 21462 4025 21508
rect 4081 21462 4133 21508
rect 4189 21462 4241 21508
rect 4297 21462 4349 21508
rect 4405 21462 4457 21508
rect 4513 21462 4565 21508
rect 4621 21462 4673 21508
rect 4729 21462 4781 21508
rect 4837 21462 4889 21508
rect 4945 21462 4997 21508
rect 5053 21462 5105 21508
rect 5161 21462 5213 21508
rect 6566 21462 6618 21508
rect 6674 21462 6726 21508
rect 6782 21462 6834 21508
rect 6890 21462 6942 21508
rect 6998 21462 7050 21508
rect 7106 21462 7158 21508
rect 7214 21462 7266 21508
rect 7322 21462 7374 21508
rect 7430 21462 7482 21508
rect 7538 21462 7590 21508
rect 9677 21462 9729 21508
rect 9785 21462 9837 21508
rect 9893 21462 9945 21508
rect 10001 21462 10053 21508
rect 10109 21462 10161 21508
rect 10217 21462 10269 21508
rect 10325 21462 10377 21508
rect 10433 21462 10485 21508
rect 10541 21462 10593 21508
rect 10649 21462 10701 21508
rect 10757 21462 10809 21508
rect 10865 21462 10917 21508
rect 10973 21462 11025 21508
rect 11081 21462 11133 21508
rect 11189 21462 11241 21508
rect 11297 21462 11349 21508
rect 11405 21462 11457 21508
rect 3433 21459 3485 21462
rect 3541 21459 3593 21462
rect 3649 21459 3701 21462
rect 3757 21459 3809 21462
rect 3865 21459 3917 21462
rect 3973 21459 4025 21462
rect 4081 21459 4133 21462
rect 4189 21459 4241 21462
rect 4297 21459 4349 21462
rect 4405 21459 4457 21462
rect 4513 21459 4565 21462
rect 4621 21459 4673 21462
rect 4729 21459 4781 21462
rect 4837 21459 4889 21462
rect 4945 21459 4997 21462
rect 5053 21459 5105 21462
rect 5161 21459 5213 21462
rect 6566 21459 6618 21462
rect 6674 21459 6726 21462
rect 6782 21459 6834 21462
rect 6890 21459 6942 21462
rect 6998 21459 7050 21462
rect 7106 21459 7158 21462
rect 7214 21459 7266 21462
rect 7322 21459 7374 21462
rect 7430 21459 7482 21462
rect 7538 21459 7590 21462
rect 9677 21459 9729 21462
rect 9785 21459 9837 21462
rect 9893 21459 9945 21462
rect 10001 21459 10053 21462
rect 10109 21459 10161 21462
rect 10217 21459 10269 21462
rect 10325 21459 10377 21462
rect 10433 21459 10485 21462
rect 10541 21459 10593 21462
rect 10649 21459 10701 21462
rect 10757 21459 10809 21462
rect 10865 21459 10917 21462
rect 10973 21459 11025 21462
rect 11081 21459 11133 21462
rect 11189 21459 11241 21462
rect 11297 21459 11349 21462
rect 11405 21459 11457 21462
rect 1505 21264 1557 21267
rect 1613 21264 1665 21267
rect 1721 21264 1773 21267
rect 1829 21264 1881 21267
rect 1937 21264 1989 21267
rect 2045 21264 2097 21267
rect 2153 21264 2205 21267
rect 2261 21264 2313 21267
rect 2369 21264 2421 21267
rect 2477 21264 2529 21267
rect 2585 21264 2637 21267
rect 2693 21264 2745 21267
rect 2801 21264 2853 21267
rect 2909 21264 2961 21267
rect 3017 21264 3069 21267
rect 3125 21264 3177 21267
rect 3233 21264 3285 21267
rect 5372 21264 5424 21267
rect 5480 21264 5532 21267
rect 5588 21264 5640 21267
rect 5696 21264 5748 21267
rect 5804 21264 5856 21267
rect 5912 21264 5964 21267
rect 6020 21264 6072 21267
rect 6128 21264 6180 21267
rect 6236 21264 6288 21267
rect 6344 21264 6396 21267
rect 7749 21264 7801 21267
rect 7857 21264 7909 21267
rect 7965 21264 8017 21267
rect 8073 21264 8125 21267
rect 8181 21264 8233 21267
rect 8289 21264 8341 21267
rect 8397 21264 8449 21267
rect 8505 21264 8557 21267
rect 8613 21264 8665 21267
rect 8721 21264 8773 21267
rect 8829 21264 8881 21267
rect 8937 21264 8989 21267
rect 9045 21264 9097 21267
rect 9153 21264 9205 21267
rect 9261 21264 9313 21267
rect 9369 21264 9421 21267
rect 9477 21264 9529 21267
rect 1505 21218 1557 21264
rect 1613 21218 1665 21264
rect 1721 21218 1773 21264
rect 1829 21218 1881 21264
rect 1937 21218 1989 21264
rect 2045 21218 2097 21264
rect 2153 21218 2205 21264
rect 2261 21218 2313 21264
rect 2369 21218 2421 21264
rect 2477 21218 2529 21264
rect 2585 21218 2637 21264
rect 2693 21218 2745 21264
rect 2801 21218 2853 21264
rect 2909 21218 2961 21264
rect 3017 21218 3069 21264
rect 3125 21218 3177 21264
rect 3233 21218 3285 21264
rect 5372 21218 5424 21264
rect 5480 21218 5532 21264
rect 5588 21218 5640 21264
rect 5696 21218 5748 21264
rect 5804 21218 5856 21264
rect 5912 21218 5964 21264
rect 6020 21218 6072 21264
rect 6128 21218 6180 21264
rect 6236 21218 6288 21264
rect 6344 21218 6396 21264
rect 7749 21218 7801 21264
rect 7857 21218 7909 21264
rect 7965 21218 8017 21264
rect 8073 21218 8125 21264
rect 8181 21218 8233 21264
rect 8289 21218 8341 21264
rect 8397 21218 8449 21264
rect 8505 21218 8557 21264
rect 8613 21218 8665 21264
rect 8721 21218 8773 21264
rect 8829 21218 8881 21264
rect 8937 21218 8989 21264
rect 9045 21218 9097 21264
rect 9153 21218 9205 21264
rect 9261 21218 9313 21264
rect 9369 21218 9421 21264
rect 9477 21218 9529 21264
rect 1505 21215 1557 21218
rect 1613 21215 1665 21218
rect 1721 21215 1773 21218
rect 1829 21215 1881 21218
rect 1937 21215 1989 21218
rect 2045 21215 2097 21218
rect 2153 21215 2205 21218
rect 2261 21215 2313 21218
rect 2369 21215 2421 21218
rect 2477 21215 2529 21218
rect 2585 21215 2637 21218
rect 2693 21215 2745 21218
rect 2801 21215 2853 21218
rect 2909 21215 2961 21218
rect 3017 21215 3069 21218
rect 3125 21215 3177 21218
rect 3233 21215 3285 21218
rect 5372 21215 5424 21218
rect 5480 21215 5532 21218
rect 5588 21215 5640 21218
rect 5696 21215 5748 21218
rect 5804 21215 5856 21218
rect 5912 21215 5964 21218
rect 6020 21215 6072 21218
rect 6128 21215 6180 21218
rect 6236 21215 6288 21218
rect 6344 21215 6396 21218
rect 7749 21215 7801 21218
rect 7857 21215 7909 21218
rect 7965 21215 8017 21218
rect 8073 21215 8125 21218
rect 8181 21215 8233 21218
rect 8289 21215 8341 21218
rect 8397 21215 8449 21218
rect 8505 21215 8557 21218
rect 8613 21215 8665 21218
rect 8721 21215 8773 21218
rect 8829 21215 8881 21218
rect 8937 21215 8989 21218
rect 9045 21215 9097 21218
rect 9153 21215 9205 21218
rect 9261 21215 9313 21218
rect 9369 21215 9421 21218
rect 9477 21215 9529 21218
rect 3433 21020 3485 21023
rect 3541 21020 3593 21023
rect 3649 21020 3701 21023
rect 3757 21020 3809 21023
rect 3865 21020 3917 21023
rect 3973 21020 4025 21023
rect 4081 21020 4133 21023
rect 4189 21020 4241 21023
rect 4297 21020 4349 21023
rect 4405 21020 4457 21023
rect 4513 21020 4565 21023
rect 4621 21020 4673 21023
rect 4729 21020 4781 21023
rect 4837 21020 4889 21023
rect 4945 21020 4997 21023
rect 5053 21020 5105 21023
rect 5161 21020 5213 21023
rect 6566 21020 6618 21023
rect 6674 21020 6726 21023
rect 6782 21020 6834 21023
rect 6890 21020 6942 21023
rect 6998 21020 7050 21023
rect 7106 21020 7158 21023
rect 7214 21020 7266 21023
rect 7322 21020 7374 21023
rect 7430 21020 7482 21023
rect 7538 21020 7590 21023
rect 9677 21020 9729 21023
rect 9785 21020 9837 21023
rect 9893 21020 9945 21023
rect 10001 21020 10053 21023
rect 10109 21020 10161 21023
rect 10217 21020 10269 21023
rect 10325 21020 10377 21023
rect 10433 21020 10485 21023
rect 10541 21020 10593 21023
rect 10649 21020 10701 21023
rect 10757 21020 10809 21023
rect 10865 21020 10917 21023
rect 10973 21020 11025 21023
rect 11081 21020 11133 21023
rect 11189 21020 11241 21023
rect 11297 21020 11349 21023
rect 11405 21020 11457 21023
rect 3433 20974 3485 21020
rect 3541 20974 3593 21020
rect 3649 20974 3701 21020
rect 3757 20974 3809 21020
rect 3865 20974 3917 21020
rect 3973 20974 4025 21020
rect 4081 20974 4133 21020
rect 4189 20974 4241 21020
rect 4297 20974 4349 21020
rect 4405 20974 4457 21020
rect 4513 20974 4565 21020
rect 4621 20974 4673 21020
rect 4729 20974 4781 21020
rect 4837 20974 4889 21020
rect 4945 20974 4997 21020
rect 5053 20974 5105 21020
rect 5161 20974 5213 21020
rect 6566 20974 6618 21020
rect 6674 20974 6726 21020
rect 6782 20974 6834 21020
rect 6890 20974 6942 21020
rect 6998 20974 7050 21020
rect 7106 20974 7158 21020
rect 7214 20974 7266 21020
rect 7322 20974 7374 21020
rect 7430 20974 7482 21020
rect 7538 20974 7590 21020
rect 9677 20974 9729 21020
rect 9785 20974 9837 21020
rect 9893 20974 9945 21020
rect 10001 20974 10053 21020
rect 10109 20974 10161 21020
rect 10217 20974 10269 21020
rect 10325 20974 10377 21020
rect 10433 20974 10485 21020
rect 10541 20974 10593 21020
rect 10649 20974 10701 21020
rect 10757 20974 10809 21020
rect 10865 20974 10917 21020
rect 10973 20974 11025 21020
rect 11081 20974 11133 21020
rect 11189 20974 11241 21020
rect 11297 20974 11349 21020
rect 11405 20974 11457 21020
rect 3433 20971 3485 20974
rect 3541 20971 3593 20974
rect 3649 20971 3701 20974
rect 3757 20971 3809 20974
rect 3865 20971 3917 20974
rect 3973 20971 4025 20974
rect 4081 20971 4133 20974
rect 4189 20971 4241 20974
rect 4297 20971 4349 20974
rect 4405 20971 4457 20974
rect 4513 20971 4565 20974
rect 4621 20971 4673 20974
rect 4729 20971 4781 20974
rect 4837 20971 4889 20974
rect 4945 20971 4997 20974
rect 5053 20971 5105 20974
rect 5161 20971 5213 20974
rect 6566 20971 6618 20974
rect 6674 20971 6726 20974
rect 6782 20971 6834 20974
rect 6890 20971 6942 20974
rect 6998 20971 7050 20974
rect 7106 20971 7158 20974
rect 7214 20971 7266 20974
rect 7322 20971 7374 20974
rect 7430 20971 7482 20974
rect 7538 20971 7590 20974
rect 9677 20971 9729 20974
rect 9785 20971 9837 20974
rect 9893 20971 9945 20974
rect 10001 20971 10053 20974
rect 10109 20971 10161 20974
rect 10217 20971 10269 20974
rect 10325 20971 10377 20974
rect 10433 20971 10485 20974
rect 10541 20971 10593 20974
rect 10649 20971 10701 20974
rect 10757 20971 10809 20974
rect 10865 20971 10917 20974
rect 10973 20971 11025 20974
rect 11081 20971 11133 20974
rect 11189 20971 11241 20974
rect 11297 20971 11349 20974
rect 11405 20971 11457 20974
rect 1505 20776 1557 20779
rect 1613 20776 1665 20779
rect 1721 20776 1773 20779
rect 1829 20776 1881 20779
rect 1937 20776 1989 20779
rect 2045 20776 2097 20779
rect 2153 20776 2205 20779
rect 2261 20776 2313 20779
rect 2369 20776 2421 20779
rect 2477 20776 2529 20779
rect 2585 20776 2637 20779
rect 2693 20776 2745 20779
rect 2801 20776 2853 20779
rect 2909 20776 2961 20779
rect 3017 20776 3069 20779
rect 3125 20776 3177 20779
rect 3233 20776 3285 20779
rect 5372 20776 5424 20779
rect 5480 20776 5532 20779
rect 5588 20776 5640 20779
rect 5696 20776 5748 20779
rect 5804 20776 5856 20779
rect 5912 20776 5964 20779
rect 6020 20776 6072 20779
rect 6128 20776 6180 20779
rect 6236 20776 6288 20779
rect 6344 20776 6396 20779
rect 7749 20776 7801 20779
rect 7857 20776 7909 20779
rect 7965 20776 8017 20779
rect 8073 20776 8125 20779
rect 8181 20776 8233 20779
rect 8289 20776 8341 20779
rect 8397 20776 8449 20779
rect 8505 20776 8557 20779
rect 8613 20776 8665 20779
rect 8721 20776 8773 20779
rect 8829 20776 8881 20779
rect 8937 20776 8989 20779
rect 9045 20776 9097 20779
rect 9153 20776 9205 20779
rect 9261 20776 9313 20779
rect 9369 20776 9421 20779
rect 9477 20776 9529 20779
rect 1505 20730 1557 20776
rect 1613 20730 1665 20776
rect 1721 20730 1773 20776
rect 1829 20730 1881 20776
rect 1937 20730 1989 20776
rect 2045 20730 2097 20776
rect 2153 20730 2205 20776
rect 2261 20730 2313 20776
rect 2369 20730 2421 20776
rect 2477 20730 2529 20776
rect 2585 20730 2637 20776
rect 2693 20730 2745 20776
rect 2801 20730 2853 20776
rect 2909 20730 2961 20776
rect 3017 20730 3069 20776
rect 3125 20730 3177 20776
rect 3233 20730 3285 20776
rect 5372 20730 5424 20776
rect 5480 20730 5532 20776
rect 5588 20730 5640 20776
rect 5696 20730 5748 20776
rect 5804 20730 5856 20776
rect 5912 20730 5964 20776
rect 6020 20730 6072 20776
rect 6128 20730 6180 20776
rect 6236 20730 6288 20776
rect 6344 20730 6396 20776
rect 7749 20730 7801 20776
rect 7857 20730 7909 20776
rect 7965 20730 8017 20776
rect 8073 20730 8125 20776
rect 8181 20730 8233 20776
rect 8289 20730 8341 20776
rect 8397 20730 8449 20776
rect 8505 20730 8557 20776
rect 8613 20730 8665 20776
rect 8721 20730 8773 20776
rect 8829 20730 8881 20776
rect 8937 20730 8989 20776
rect 9045 20730 9097 20776
rect 9153 20730 9205 20776
rect 9261 20730 9313 20776
rect 9369 20730 9421 20776
rect 9477 20730 9529 20776
rect 1505 20727 1557 20730
rect 1613 20727 1665 20730
rect 1721 20727 1773 20730
rect 1829 20727 1881 20730
rect 1937 20727 1989 20730
rect 2045 20727 2097 20730
rect 2153 20727 2205 20730
rect 2261 20727 2313 20730
rect 2369 20727 2421 20730
rect 2477 20727 2529 20730
rect 2585 20727 2637 20730
rect 2693 20727 2745 20730
rect 2801 20727 2853 20730
rect 2909 20727 2961 20730
rect 3017 20727 3069 20730
rect 3125 20727 3177 20730
rect 3233 20727 3285 20730
rect 5372 20727 5424 20730
rect 5480 20727 5532 20730
rect 5588 20727 5640 20730
rect 5696 20727 5748 20730
rect 5804 20727 5856 20730
rect 5912 20727 5964 20730
rect 6020 20727 6072 20730
rect 6128 20727 6180 20730
rect 6236 20727 6288 20730
rect 6344 20727 6396 20730
rect 7749 20727 7801 20730
rect 7857 20727 7909 20730
rect 7965 20727 8017 20730
rect 8073 20727 8125 20730
rect 8181 20727 8233 20730
rect 8289 20727 8341 20730
rect 8397 20727 8449 20730
rect 8505 20727 8557 20730
rect 8613 20727 8665 20730
rect 8721 20727 8773 20730
rect 8829 20727 8881 20730
rect 8937 20727 8989 20730
rect 9045 20727 9097 20730
rect 9153 20727 9205 20730
rect 9261 20727 9313 20730
rect 9369 20727 9421 20730
rect 9477 20727 9529 20730
rect 3433 20532 3485 20535
rect 3541 20532 3593 20535
rect 3649 20532 3701 20535
rect 3757 20532 3809 20535
rect 3865 20532 3917 20535
rect 3973 20532 4025 20535
rect 4081 20532 4133 20535
rect 4189 20532 4241 20535
rect 4297 20532 4349 20535
rect 4405 20532 4457 20535
rect 4513 20532 4565 20535
rect 4621 20532 4673 20535
rect 4729 20532 4781 20535
rect 4837 20532 4889 20535
rect 4945 20532 4997 20535
rect 5053 20532 5105 20535
rect 5161 20532 5213 20535
rect 6566 20532 6618 20535
rect 6674 20532 6726 20535
rect 6782 20532 6834 20535
rect 6890 20532 6942 20535
rect 6998 20532 7050 20535
rect 7106 20532 7158 20535
rect 7214 20532 7266 20535
rect 7322 20532 7374 20535
rect 7430 20532 7482 20535
rect 7538 20532 7590 20535
rect 9677 20532 9729 20535
rect 9785 20532 9837 20535
rect 9893 20532 9945 20535
rect 10001 20532 10053 20535
rect 10109 20532 10161 20535
rect 10217 20532 10269 20535
rect 10325 20532 10377 20535
rect 10433 20532 10485 20535
rect 10541 20532 10593 20535
rect 10649 20532 10701 20535
rect 10757 20532 10809 20535
rect 10865 20532 10917 20535
rect 10973 20532 11025 20535
rect 11081 20532 11133 20535
rect 11189 20532 11241 20535
rect 11297 20532 11349 20535
rect 11405 20532 11457 20535
rect 3433 20486 3485 20532
rect 3541 20486 3593 20532
rect 3649 20486 3701 20532
rect 3757 20486 3809 20532
rect 3865 20486 3917 20532
rect 3973 20486 4025 20532
rect 4081 20486 4133 20532
rect 4189 20486 4241 20532
rect 4297 20486 4349 20532
rect 4405 20486 4457 20532
rect 4513 20486 4565 20532
rect 4621 20486 4673 20532
rect 4729 20486 4781 20532
rect 4837 20486 4889 20532
rect 4945 20486 4997 20532
rect 5053 20486 5105 20532
rect 5161 20486 5213 20532
rect 6566 20486 6618 20532
rect 6674 20486 6726 20532
rect 6782 20486 6834 20532
rect 6890 20486 6942 20532
rect 6998 20486 7050 20532
rect 7106 20486 7158 20532
rect 7214 20486 7266 20532
rect 7322 20486 7374 20532
rect 7430 20486 7482 20532
rect 7538 20486 7590 20532
rect 9677 20486 9729 20532
rect 9785 20486 9837 20532
rect 9893 20486 9945 20532
rect 10001 20486 10053 20532
rect 10109 20486 10161 20532
rect 10217 20486 10269 20532
rect 10325 20486 10377 20532
rect 10433 20486 10485 20532
rect 10541 20486 10593 20532
rect 10649 20486 10701 20532
rect 10757 20486 10809 20532
rect 10865 20486 10917 20532
rect 10973 20486 11025 20532
rect 11081 20486 11133 20532
rect 11189 20486 11241 20532
rect 11297 20486 11349 20532
rect 11405 20486 11457 20532
rect 3433 20483 3485 20486
rect 3541 20483 3593 20486
rect 3649 20483 3701 20486
rect 3757 20483 3809 20486
rect 3865 20483 3917 20486
rect 3973 20483 4025 20486
rect 4081 20483 4133 20486
rect 4189 20483 4241 20486
rect 4297 20483 4349 20486
rect 4405 20483 4457 20486
rect 4513 20483 4565 20486
rect 4621 20483 4673 20486
rect 4729 20483 4781 20486
rect 4837 20483 4889 20486
rect 4945 20483 4997 20486
rect 5053 20483 5105 20486
rect 5161 20483 5213 20486
rect 6566 20483 6618 20486
rect 6674 20483 6726 20486
rect 6782 20483 6834 20486
rect 6890 20483 6942 20486
rect 6998 20483 7050 20486
rect 7106 20483 7158 20486
rect 7214 20483 7266 20486
rect 7322 20483 7374 20486
rect 7430 20483 7482 20486
rect 7538 20483 7590 20486
rect 9677 20483 9729 20486
rect 9785 20483 9837 20486
rect 9893 20483 9945 20486
rect 10001 20483 10053 20486
rect 10109 20483 10161 20486
rect 10217 20483 10269 20486
rect 10325 20483 10377 20486
rect 10433 20483 10485 20486
rect 10541 20483 10593 20486
rect 10649 20483 10701 20486
rect 10757 20483 10809 20486
rect 10865 20483 10917 20486
rect 10973 20483 11025 20486
rect 11081 20483 11133 20486
rect 11189 20483 11241 20486
rect 11297 20483 11349 20486
rect 11405 20483 11457 20486
rect 1505 20288 1557 20291
rect 1613 20288 1665 20291
rect 1721 20288 1773 20291
rect 1829 20288 1881 20291
rect 1937 20288 1989 20291
rect 2045 20288 2097 20291
rect 2153 20288 2205 20291
rect 2261 20288 2313 20291
rect 2369 20288 2421 20291
rect 2477 20288 2529 20291
rect 2585 20288 2637 20291
rect 2693 20288 2745 20291
rect 2801 20288 2853 20291
rect 2909 20288 2961 20291
rect 3017 20288 3069 20291
rect 3125 20288 3177 20291
rect 3233 20288 3285 20291
rect 5372 20288 5424 20291
rect 5480 20288 5532 20291
rect 5588 20288 5640 20291
rect 5696 20288 5748 20291
rect 5804 20288 5856 20291
rect 5912 20288 5964 20291
rect 6020 20288 6072 20291
rect 6128 20288 6180 20291
rect 6236 20288 6288 20291
rect 6344 20288 6396 20291
rect 7749 20288 7801 20291
rect 7857 20288 7909 20291
rect 7965 20288 8017 20291
rect 8073 20288 8125 20291
rect 8181 20288 8233 20291
rect 8289 20288 8341 20291
rect 8397 20288 8449 20291
rect 8505 20288 8557 20291
rect 8613 20288 8665 20291
rect 8721 20288 8773 20291
rect 8829 20288 8881 20291
rect 8937 20288 8989 20291
rect 9045 20288 9097 20291
rect 9153 20288 9205 20291
rect 9261 20288 9313 20291
rect 9369 20288 9421 20291
rect 9477 20288 9529 20291
rect 1505 20242 1557 20288
rect 1613 20242 1665 20288
rect 1721 20242 1773 20288
rect 1829 20242 1881 20288
rect 1937 20242 1989 20288
rect 2045 20242 2097 20288
rect 2153 20242 2205 20288
rect 2261 20242 2313 20288
rect 2369 20242 2421 20288
rect 2477 20242 2529 20288
rect 2585 20242 2637 20288
rect 2693 20242 2745 20288
rect 2801 20242 2853 20288
rect 2909 20242 2961 20288
rect 3017 20242 3069 20288
rect 3125 20242 3177 20288
rect 3233 20242 3285 20288
rect 5372 20242 5424 20288
rect 5480 20242 5532 20288
rect 5588 20242 5640 20288
rect 5696 20242 5748 20288
rect 5804 20242 5856 20288
rect 5912 20242 5964 20288
rect 6020 20242 6072 20288
rect 6128 20242 6180 20288
rect 6236 20242 6288 20288
rect 6344 20242 6396 20288
rect 7749 20242 7801 20288
rect 7857 20242 7909 20288
rect 7965 20242 8017 20288
rect 8073 20242 8125 20288
rect 8181 20242 8233 20288
rect 8289 20242 8341 20288
rect 8397 20242 8449 20288
rect 8505 20242 8557 20288
rect 8613 20242 8665 20288
rect 8721 20242 8773 20288
rect 8829 20242 8881 20288
rect 8937 20242 8989 20288
rect 9045 20242 9097 20288
rect 9153 20242 9205 20288
rect 9261 20242 9313 20288
rect 9369 20242 9421 20288
rect 9477 20242 9529 20288
rect 1505 20239 1557 20242
rect 1613 20239 1665 20242
rect 1721 20239 1773 20242
rect 1829 20239 1881 20242
rect 1937 20239 1989 20242
rect 2045 20239 2097 20242
rect 2153 20239 2205 20242
rect 2261 20239 2313 20242
rect 2369 20239 2421 20242
rect 2477 20239 2529 20242
rect 2585 20239 2637 20242
rect 2693 20239 2745 20242
rect 2801 20239 2853 20242
rect 2909 20239 2961 20242
rect 3017 20239 3069 20242
rect 3125 20239 3177 20242
rect 3233 20239 3285 20242
rect 5372 20239 5424 20242
rect 5480 20239 5532 20242
rect 5588 20239 5640 20242
rect 5696 20239 5748 20242
rect 5804 20239 5856 20242
rect 5912 20239 5964 20242
rect 6020 20239 6072 20242
rect 6128 20239 6180 20242
rect 6236 20239 6288 20242
rect 6344 20239 6396 20242
rect 7749 20239 7801 20242
rect 7857 20239 7909 20242
rect 7965 20239 8017 20242
rect 8073 20239 8125 20242
rect 8181 20239 8233 20242
rect 8289 20239 8341 20242
rect 8397 20239 8449 20242
rect 8505 20239 8557 20242
rect 8613 20239 8665 20242
rect 8721 20239 8773 20242
rect 8829 20239 8881 20242
rect 8937 20239 8989 20242
rect 9045 20239 9097 20242
rect 9153 20239 9205 20242
rect 9261 20239 9313 20242
rect 9369 20239 9421 20242
rect 9477 20239 9529 20242
rect 3433 20044 3485 20047
rect 3541 20044 3593 20047
rect 3649 20044 3701 20047
rect 3757 20044 3809 20047
rect 3865 20044 3917 20047
rect 3973 20044 4025 20047
rect 4081 20044 4133 20047
rect 4189 20044 4241 20047
rect 4297 20044 4349 20047
rect 4405 20044 4457 20047
rect 4513 20044 4565 20047
rect 4621 20044 4673 20047
rect 4729 20044 4781 20047
rect 4837 20044 4889 20047
rect 4945 20044 4997 20047
rect 5053 20044 5105 20047
rect 5161 20044 5213 20047
rect 6566 20044 6618 20047
rect 6674 20044 6726 20047
rect 6782 20044 6834 20047
rect 6890 20044 6942 20047
rect 6998 20044 7050 20047
rect 7106 20044 7158 20047
rect 7214 20044 7266 20047
rect 7322 20044 7374 20047
rect 7430 20044 7482 20047
rect 7538 20044 7590 20047
rect 9677 20044 9729 20047
rect 9785 20044 9837 20047
rect 9893 20044 9945 20047
rect 10001 20044 10053 20047
rect 10109 20044 10161 20047
rect 10217 20044 10269 20047
rect 10325 20044 10377 20047
rect 10433 20044 10485 20047
rect 10541 20044 10593 20047
rect 10649 20044 10701 20047
rect 10757 20044 10809 20047
rect 10865 20044 10917 20047
rect 10973 20044 11025 20047
rect 11081 20044 11133 20047
rect 11189 20044 11241 20047
rect 11297 20044 11349 20047
rect 11405 20044 11457 20047
rect 3433 19998 3485 20044
rect 3541 19998 3593 20044
rect 3649 19998 3701 20044
rect 3757 19998 3809 20044
rect 3865 19998 3917 20044
rect 3973 19998 4025 20044
rect 4081 19998 4133 20044
rect 4189 19998 4241 20044
rect 4297 19998 4349 20044
rect 4405 19998 4457 20044
rect 4513 19998 4565 20044
rect 4621 19998 4673 20044
rect 4729 19998 4781 20044
rect 4837 19998 4889 20044
rect 4945 19998 4997 20044
rect 5053 19998 5105 20044
rect 5161 19998 5213 20044
rect 6566 19998 6618 20044
rect 6674 19998 6726 20044
rect 6782 19998 6834 20044
rect 6890 19998 6942 20044
rect 6998 19998 7050 20044
rect 7106 19998 7158 20044
rect 7214 19998 7266 20044
rect 7322 19998 7374 20044
rect 7430 19998 7482 20044
rect 7538 19998 7590 20044
rect 9677 19998 9729 20044
rect 9785 19998 9837 20044
rect 9893 19998 9945 20044
rect 10001 19998 10053 20044
rect 10109 19998 10161 20044
rect 10217 19998 10269 20044
rect 10325 19998 10377 20044
rect 10433 19998 10485 20044
rect 10541 19998 10593 20044
rect 10649 19998 10701 20044
rect 10757 19998 10809 20044
rect 10865 19998 10917 20044
rect 10973 19998 11025 20044
rect 11081 19998 11133 20044
rect 11189 19998 11241 20044
rect 11297 19998 11349 20044
rect 11405 19998 11457 20044
rect 3433 19995 3485 19998
rect 3541 19995 3593 19998
rect 3649 19995 3701 19998
rect 3757 19995 3809 19998
rect 3865 19995 3917 19998
rect 3973 19995 4025 19998
rect 4081 19995 4133 19998
rect 4189 19995 4241 19998
rect 4297 19995 4349 19998
rect 4405 19995 4457 19998
rect 4513 19995 4565 19998
rect 4621 19995 4673 19998
rect 4729 19995 4781 19998
rect 4837 19995 4889 19998
rect 4945 19995 4997 19998
rect 5053 19995 5105 19998
rect 5161 19995 5213 19998
rect 6566 19995 6618 19998
rect 6674 19995 6726 19998
rect 6782 19995 6834 19998
rect 6890 19995 6942 19998
rect 6998 19995 7050 19998
rect 7106 19995 7158 19998
rect 7214 19995 7266 19998
rect 7322 19995 7374 19998
rect 7430 19995 7482 19998
rect 7538 19995 7590 19998
rect 9677 19995 9729 19998
rect 9785 19995 9837 19998
rect 9893 19995 9945 19998
rect 10001 19995 10053 19998
rect 10109 19995 10161 19998
rect 10217 19995 10269 19998
rect 10325 19995 10377 19998
rect 10433 19995 10485 19998
rect 10541 19995 10593 19998
rect 10649 19995 10701 19998
rect 10757 19995 10809 19998
rect 10865 19995 10917 19998
rect 10973 19995 11025 19998
rect 11081 19995 11133 19998
rect 11189 19995 11241 19998
rect 11297 19995 11349 19998
rect 11405 19995 11457 19998
rect 1505 19800 1557 19803
rect 1613 19800 1665 19803
rect 1721 19800 1773 19803
rect 1829 19800 1881 19803
rect 1937 19800 1989 19803
rect 2045 19800 2097 19803
rect 2153 19800 2205 19803
rect 2261 19800 2313 19803
rect 2369 19800 2421 19803
rect 2477 19800 2529 19803
rect 2585 19800 2637 19803
rect 2693 19800 2745 19803
rect 2801 19800 2853 19803
rect 2909 19800 2961 19803
rect 3017 19800 3069 19803
rect 3125 19800 3177 19803
rect 3233 19800 3285 19803
rect 5372 19800 5424 19803
rect 5480 19800 5532 19803
rect 5588 19800 5640 19803
rect 5696 19800 5748 19803
rect 5804 19800 5856 19803
rect 5912 19800 5964 19803
rect 6020 19800 6072 19803
rect 6128 19800 6180 19803
rect 6236 19800 6288 19803
rect 6344 19800 6396 19803
rect 7749 19800 7801 19803
rect 7857 19800 7909 19803
rect 7965 19800 8017 19803
rect 8073 19800 8125 19803
rect 8181 19800 8233 19803
rect 8289 19800 8341 19803
rect 8397 19800 8449 19803
rect 8505 19800 8557 19803
rect 8613 19800 8665 19803
rect 8721 19800 8773 19803
rect 8829 19800 8881 19803
rect 8937 19800 8989 19803
rect 9045 19800 9097 19803
rect 9153 19800 9205 19803
rect 9261 19800 9313 19803
rect 9369 19800 9421 19803
rect 9477 19800 9529 19803
rect 1505 19754 1557 19800
rect 1613 19754 1665 19800
rect 1721 19754 1773 19800
rect 1829 19754 1881 19800
rect 1937 19754 1989 19800
rect 2045 19754 2097 19800
rect 2153 19754 2205 19800
rect 2261 19754 2313 19800
rect 2369 19754 2421 19800
rect 2477 19754 2529 19800
rect 2585 19754 2637 19800
rect 2693 19754 2745 19800
rect 2801 19754 2853 19800
rect 2909 19754 2961 19800
rect 3017 19754 3069 19800
rect 3125 19754 3177 19800
rect 3233 19754 3285 19800
rect 5372 19754 5424 19800
rect 5480 19754 5532 19800
rect 5588 19754 5640 19800
rect 5696 19754 5748 19800
rect 5804 19754 5856 19800
rect 5912 19754 5964 19800
rect 6020 19754 6072 19800
rect 6128 19754 6180 19800
rect 6236 19754 6288 19800
rect 6344 19754 6396 19800
rect 7749 19754 7801 19800
rect 7857 19754 7909 19800
rect 7965 19754 8017 19800
rect 8073 19754 8125 19800
rect 8181 19754 8233 19800
rect 8289 19754 8341 19800
rect 8397 19754 8449 19800
rect 8505 19754 8557 19800
rect 8613 19754 8665 19800
rect 8721 19754 8773 19800
rect 8829 19754 8881 19800
rect 8937 19754 8989 19800
rect 9045 19754 9097 19800
rect 9153 19754 9205 19800
rect 9261 19754 9313 19800
rect 9369 19754 9421 19800
rect 9477 19754 9529 19800
rect 1505 19751 1557 19754
rect 1613 19751 1665 19754
rect 1721 19751 1773 19754
rect 1829 19751 1881 19754
rect 1937 19751 1989 19754
rect 2045 19751 2097 19754
rect 2153 19751 2205 19754
rect 2261 19751 2313 19754
rect 2369 19751 2421 19754
rect 2477 19751 2529 19754
rect 2585 19751 2637 19754
rect 2693 19751 2745 19754
rect 2801 19751 2853 19754
rect 2909 19751 2961 19754
rect 3017 19751 3069 19754
rect 3125 19751 3177 19754
rect 3233 19751 3285 19754
rect 5372 19751 5424 19754
rect 5480 19751 5532 19754
rect 5588 19751 5640 19754
rect 5696 19751 5748 19754
rect 5804 19751 5856 19754
rect 5912 19751 5964 19754
rect 6020 19751 6072 19754
rect 6128 19751 6180 19754
rect 6236 19751 6288 19754
rect 6344 19751 6396 19754
rect 7749 19751 7801 19754
rect 7857 19751 7909 19754
rect 7965 19751 8017 19754
rect 8073 19751 8125 19754
rect 8181 19751 8233 19754
rect 8289 19751 8341 19754
rect 8397 19751 8449 19754
rect 8505 19751 8557 19754
rect 8613 19751 8665 19754
rect 8721 19751 8773 19754
rect 8829 19751 8881 19754
rect 8937 19751 8989 19754
rect 9045 19751 9097 19754
rect 9153 19751 9205 19754
rect 9261 19751 9313 19754
rect 9369 19751 9421 19754
rect 9477 19751 9529 19754
rect 3433 19556 3485 19559
rect 3541 19556 3593 19559
rect 3649 19556 3701 19559
rect 3757 19556 3809 19559
rect 3865 19556 3917 19559
rect 3973 19556 4025 19559
rect 4081 19556 4133 19559
rect 4189 19556 4241 19559
rect 4297 19556 4349 19559
rect 4405 19556 4457 19559
rect 4513 19556 4565 19559
rect 4621 19556 4673 19559
rect 4729 19556 4781 19559
rect 4837 19556 4889 19559
rect 4945 19556 4997 19559
rect 5053 19556 5105 19559
rect 5161 19556 5213 19559
rect 6566 19556 6618 19559
rect 6674 19556 6726 19559
rect 6782 19556 6834 19559
rect 6890 19556 6942 19559
rect 6998 19556 7050 19559
rect 7106 19556 7158 19559
rect 7214 19556 7266 19559
rect 7322 19556 7374 19559
rect 7430 19556 7482 19559
rect 7538 19556 7590 19559
rect 9677 19556 9729 19559
rect 9785 19556 9837 19559
rect 9893 19556 9945 19559
rect 10001 19556 10053 19559
rect 10109 19556 10161 19559
rect 10217 19556 10269 19559
rect 10325 19556 10377 19559
rect 10433 19556 10485 19559
rect 10541 19556 10593 19559
rect 10649 19556 10701 19559
rect 10757 19556 10809 19559
rect 10865 19556 10917 19559
rect 10973 19556 11025 19559
rect 11081 19556 11133 19559
rect 11189 19556 11241 19559
rect 11297 19556 11349 19559
rect 11405 19556 11457 19559
rect 3433 19510 3485 19556
rect 3541 19510 3593 19556
rect 3649 19510 3701 19556
rect 3757 19510 3809 19556
rect 3865 19510 3917 19556
rect 3973 19510 4025 19556
rect 4081 19510 4133 19556
rect 4189 19510 4241 19556
rect 4297 19510 4349 19556
rect 4405 19510 4457 19556
rect 4513 19510 4565 19556
rect 4621 19510 4673 19556
rect 4729 19510 4781 19556
rect 4837 19510 4889 19556
rect 4945 19510 4997 19556
rect 5053 19510 5105 19556
rect 5161 19510 5213 19556
rect 6566 19510 6618 19556
rect 6674 19510 6726 19556
rect 6782 19510 6834 19556
rect 6890 19510 6942 19556
rect 6998 19510 7050 19556
rect 7106 19510 7158 19556
rect 7214 19510 7266 19556
rect 7322 19510 7374 19556
rect 7430 19510 7482 19556
rect 7538 19510 7590 19556
rect 9677 19510 9729 19556
rect 9785 19510 9837 19556
rect 9893 19510 9945 19556
rect 10001 19510 10053 19556
rect 10109 19510 10161 19556
rect 10217 19510 10269 19556
rect 10325 19510 10377 19556
rect 10433 19510 10485 19556
rect 10541 19510 10593 19556
rect 10649 19510 10701 19556
rect 10757 19510 10809 19556
rect 10865 19510 10917 19556
rect 10973 19510 11025 19556
rect 11081 19510 11133 19556
rect 11189 19510 11241 19556
rect 11297 19510 11349 19556
rect 11405 19510 11457 19556
rect 3433 19507 3485 19510
rect 3541 19507 3593 19510
rect 3649 19507 3701 19510
rect 3757 19507 3809 19510
rect 3865 19507 3917 19510
rect 3973 19507 4025 19510
rect 4081 19507 4133 19510
rect 4189 19507 4241 19510
rect 4297 19507 4349 19510
rect 4405 19507 4457 19510
rect 4513 19507 4565 19510
rect 4621 19507 4673 19510
rect 4729 19507 4781 19510
rect 4837 19507 4889 19510
rect 4945 19507 4997 19510
rect 5053 19507 5105 19510
rect 5161 19507 5213 19510
rect 6566 19507 6618 19510
rect 6674 19507 6726 19510
rect 6782 19507 6834 19510
rect 6890 19507 6942 19510
rect 6998 19507 7050 19510
rect 7106 19507 7158 19510
rect 7214 19507 7266 19510
rect 7322 19507 7374 19510
rect 7430 19507 7482 19510
rect 7538 19507 7590 19510
rect 9677 19507 9729 19510
rect 9785 19507 9837 19510
rect 9893 19507 9945 19510
rect 10001 19507 10053 19510
rect 10109 19507 10161 19510
rect 10217 19507 10269 19510
rect 10325 19507 10377 19510
rect 10433 19507 10485 19510
rect 10541 19507 10593 19510
rect 10649 19507 10701 19510
rect 10757 19507 10809 19510
rect 10865 19507 10917 19510
rect 10973 19507 11025 19510
rect 11081 19507 11133 19510
rect 11189 19507 11241 19510
rect 11297 19507 11349 19510
rect 11405 19507 11457 19510
rect 1505 19312 1557 19315
rect 1613 19312 1665 19315
rect 1721 19312 1773 19315
rect 1829 19312 1881 19315
rect 1937 19312 1989 19315
rect 2045 19312 2097 19315
rect 2153 19312 2205 19315
rect 2261 19312 2313 19315
rect 2369 19312 2421 19315
rect 2477 19312 2529 19315
rect 2585 19312 2637 19315
rect 2693 19312 2745 19315
rect 2801 19312 2853 19315
rect 2909 19312 2961 19315
rect 3017 19312 3069 19315
rect 3125 19312 3177 19315
rect 3233 19312 3285 19315
rect 5372 19312 5424 19315
rect 5480 19312 5532 19315
rect 5588 19312 5640 19315
rect 5696 19312 5748 19315
rect 5804 19312 5856 19315
rect 5912 19312 5964 19315
rect 6020 19312 6072 19315
rect 6128 19312 6180 19315
rect 6236 19312 6288 19315
rect 6344 19312 6396 19315
rect 7749 19312 7801 19315
rect 7857 19312 7909 19315
rect 7965 19312 8017 19315
rect 8073 19312 8125 19315
rect 8181 19312 8233 19315
rect 8289 19312 8341 19315
rect 8397 19312 8449 19315
rect 8505 19312 8557 19315
rect 8613 19312 8665 19315
rect 8721 19312 8773 19315
rect 8829 19312 8881 19315
rect 8937 19312 8989 19315
rect 9045 19312 9097 19315
rect 9153 19312 9205 19315
rect 9261 19312 9313 19315
rect 9369 19312 9421 19315
rect 9477 19312 9529 19315
rect 1505 19266 1557 19312
rect 1613 19266 1665 19312
rect 1721 19266 1773 19312
rect 1829 19266 1881 19312
rect 1937 19266 1989 19312
rect 2045 19266 2097 19312
rect 2153 19266 2205 19312
rect 2261 19266 2313 19312
rect 2369 19266 2421 19312
rect 2477 19266 2529 19312
rect 2585 19266 2637 19312
rect 2693 19266 2745 19312
rect 2801 19266 2853 19312
rect 2909 19266 2961 19312
rect 3017 19266 3069 19312
rect 3125 19266 3177 19312
rect 3233 19266 3285 19312
rect 5372 19266 5424 19312
rect 5480 19266 5532 19312
rect 5588 19266 5640 19312
rect 5696 19266 5748 19312
rect 5804 19266 5856 19312
rect 5912 19266 5964 19312
rect 6020 19266 6072 19312
rect 6128 19266 6180 19312
rect 6236 19266 6288 19312
rect 6344 19266 6396 19312
rect 7749 19266 7801 19312
rect 7857 19266 7909 19312
rect 7965 19266 8017 19312
rect 8073 19266 8125 19312
rect 8181 19266 8233 19312
rect 8289 19266 8341 19312
rect 8397 19266 8449 19312
rect 8505 19266 8557 19312
rect 8613 19266 8665 19312
rect 8721 19266 8773 19312
rect 8829 19266 8881 19312
rect 8937 19266 8989 19312
rect 9045 19266 9097 19312
rect 9153 19266 9205 19312
rect 9261 19266 9313 19312
rect 9369 19266 9421 19312
rect 9477 19266 9529 19312
rect 1505 19263 1557 19266
rect 1613 19263 1665 19266
rect 1721 19263 1773 19266
rect 1829 19263 1881 19266
rect 1937 19263 1989 19266
rect 2045 19263 2097 19266
rect 2153 19263 2205 19266
rect 2261 19263 2313 19266
rect 2369 19263 2421 19266
rect 2477 19263 2529 19266
rect 2585 19263 2637 19266
rect 2693 19263 2745 19266
rect 2801 19263 2853 19266
rect 2909 19263 2961 19266
rect 3017 19263 3069 19266
rect 3125 19263 3177 19266
rect 3233 19263 3285 19266
rect 5372 19263 5424 19266
rect 5480 19263 5532 19266
rect 5588 19263 5640 19266
rect 5696 19263 5748 19266
rect 5804 19263 5856 19266
rect 5912 19263 5964 19266
rect 6020 19263 6072 19266
rect 6128 19263 6180 19266
rect 6236 19263 6288 19266
rect 6344 19263 6396 19266
rect 7749 19263 7801 19266
rect 7857 19263 7909 19266
rect 7965 19263 8017 19266
rect 8073 19263 8125 19266
rect 8181 19263 8233 19266
rect 8289 19263 8341 19266
rect 8397 19263 8449 19266
rect 8505 19263 8557 19266
rect 8613 19263 8665 19266
rect 8721 19263 8773 19266
rect 8829 19263 8881 19266
rect 8937 19263 8989 19266
rect 9045 19263 9097 19266
rect 9153 19263 9205 19266
rect 9261 19263 9313 19266
rect 9369 19263 9421 19266
rect 9477 19263 9529 19266
rect 1233 19083 1285 19135
rect 1341 19083 1393 19135
rect 11569 23727 11621 23779
rect 11677 23727 11706 23779
rect 11706 23727 11729 23779
rect 11569 23619 11621 23671
rect 11677 23619 11706 23671
rect 11706 23619 11729 23671
rect 11569 23511 11621 23563
rect 11677 23511 11706 23563
rect 11706 23511 11729 23563
rect 11569 23403 11621 23455
rect 11677 23403 11706 23455
rect 11706 23403 11729 23455
rect 11569 23295 11621 23347
rect 11677 23295 11706 23347
rect 11706 23295 11729 23347
rect 11569 23187 11621 23239
rect 11677 23187 11706 23239
rect 11706 23187 11729 23239
rect 11569 23079 11621 23131
rect 11677 23079 11706 23131
rect 11706 23079 11729 23131
rect 11569 22971 11621 23023
rect 11677 22971 11706 23023
rect 11706 22971 11729 23023
rect 11569 22863 11621 22915
rect 11677 22863 11706 22915
rect 11706 22863 11729 22915
rect 11569 22755 11621 22807
rect 11677 22755 11706 22807
rect 11706 22755 11729 22807
rect 11569 22647 11621 22699
rect 11677 22647 11706 22699
rect 11706 22647 11729 22699
rect 11569 22539 11621 22591
rect 11677 22539 11706 22591
rect 11706 22539 11729 22591
rect 11569 22431 11621 22483
rect 11677 22431 11706 22483
rect 11706 22431 11729 22483
rect 11569 22323 11621 22375
rect 11677 22323 11706 22375
rect 11706 22323 11729 22375
rect 11569 22215 11621 22267
rect 11677 22215 11706 22267
rect 11706 22215 11729 22267
rect 11569 22107 11621 22159
rect 11677 22107 11706 22159
rect 11706 22107 11729 22159
rect 11569 21999 11621 22051
rect 11677 21999 11706 22051
rect 11706 21999 11729 22051
rect 11569 21891 11621 21943
rect 11677 21891 11706 21943
rect 11706 21891 11729 21943
rect 11569 21783 11621 21835
rect 11677 21783 11706 21835
rect 11706 21783 11729 21835
rect 11569 21675 11621 21727
rect 11677 21675 11706 21727
rect 11706 21675 11729 21727
rect 11569 21567 11621 21619
rect 11677 21567 11706 21619
rect 11706 21567 11729 21619
rect 11569 21459 11621 21511
rect 11677 21459 11706 21511
rect 11706 21459 11729 21511
rect 11569 21351 11621 21403
rect 11677 21351 11706 21403
rect 11706 21351 11729 21403
rect 11569 21243 11621 21295
rect 11677 21243 11706 21295
rect 11706 21243 11729 21295
rect 11569 21135 11621 21187
rect 11677 21135 11706 21187
rect 11706 21135 11729 21187
rect 11569 21027 11621 21079
rect 11677 21027 11706 21079
rect 11706 21027 11729 21079
rect 11569 20919 11621 20971
rect 11677 20919 11706 20971
rect 11706 20919 11729 20971
rect 11569 20811 11621 20863
rect 11677 20811 11706 20863
rect 11706 20811 11729 20863
rect 11569 20703 11621 20755
rect 11677 20703 11706 20755
rect 11706 20703 11729 20755
rect 11569 20595 11621 20647
rect 11677 20595 11706 20647
rect 11706 20595 11729 20647
rect 11569 20487 11621 20539
rect 11677 20487 11706 20539
rect 11706 20487 11729 20539
rect 11569 20379 11621 20431
rect 11677 20379 11706 20431
rect 11706 20379 11729 20431
rect 11569 20271 11621 20323
rect 11677 20271 11706 20323
rect 11706 20271 11729 20323
rect 11569 20163 11621 20215
rect 11677 20163 11706 20215
rect 11706 20163 11729 20215
rect 11569 20055 11621 20107
rect 11677 20055 11706 20107
rect 11706 20055 11729 20107
rect 11569 19947 11621 19999
rect 11677 19947 11706 19999
rect 11706 19947 11729 19999
rect 11569 19839 11621 19891
rect 11677 19839 11706 19891
rect 11706 19839 11729 19891
rect 11569 19731 11621 19783
rect 11677 19731 11706 19783
rect 11706 19731 11729 19783
rect 11569 19623 11621 19675
rect 11677 19623 11706 19675
rect 11706 19623 11729 19675
rect 11569 19515 11621 19567
rect 11677 19515 11706 19567
rect 11706 19515 11729 19567
rect 11569 19407 11621 19459
rect 11677 19407 11706 19459
rect 11706 19407 11729 19459
rect 11569 19299 11621 19351
rect 11677 19299 11706 19351
rect 11706 19299 11729 19351
rect 11569 19191 11621 19243
rect 11677 19191 11706 19243
rect 11706 19191 11729 19243
rect 11569 19083 11621 19135
rect 11677 19083 11729 19135
rect 3433 19068 3485 19071
rect 3541 19068 3593 19071
rect 3649 19068 3701 19071
rect 3757 19068 3809 19071
rect 3865 19068 3917 19071
rect 3973 19068 4025 19071
rect 4081 19068 4133 19071
rect 4189 19068 4241 19071
rect 4297 19068 4349 19071
rect 4405 19068 4457 19071
rect 4513 19068 4565 19071
rect 4621 19068 4673 19071
rect 4729 19068 4781 19071
rect 4837 19068 4889 19071
rect 4945 19068 4997 19071
rect 5053 19068 5105 19071
rect 5161 19068 5213 19071
rect 6566 19068 6618 19071
rect 6674 19068 6726 19071
rect 6782 19068 6834 19071
rect 6890 19068 6942 19071
rect 6998 19068 7050 19071
rect 7106 19068 7158 19071
rect 7214 19068 7266 19071
rect 7322 19068 7374 19071
rect 7430 19068 7482 19071
rect 7538 19068 7590 19071
rect 9677 19068 9729 19071
rect 9785 19068 9837 19071
rect 9893 19068 9945 19071
rect 10001 19068 10053 19071
rect 10109 19068 10161 19071
rect 10217 19068 10269 19071
rect 10325 19068 10377 19071
rect 10433 19068 10485 19071
rect 10541 19068 10593 19071
rect 10649 19068 10701 19071
rect 10757 19068 10809 19071
rect 10865 19068 10917 19071
rect 10973 19068 11025 19071
rect 11081 19068 11133 19071
rect 11189 19068 11241 19071
rect 11297 19068 11349 19071
rect 11405 19068 11457 19071
rect 3433 19022 3485 19068
rect 3541 19022 3593 19068
rect 3649 19022 3701 19068
rect 3757 19022 3809 19068
rect 3865 19022 3917 19068
rect 3973 19022 4025 19068
rect 4081 19022 4133 19068
rect 4189 19022 4241 19068
rect 4297 19022 4349 19068
rect 4405 19022 4457 19068
rect 4513 19022 4565 19068
rect 4621 19022 4673 19068
rect 4729 19022 4781 19068
rect 4837 19022 4889 19068
rect 4945 19022 4997 19068
rect 5053 19022 5105 19068
rect 5161 19022 5213 19068
rect 6566 19022 6618 19068
rect 6674 19022 6726 19068
rect 6782 19022 6834 19068
rect 6890 19022 6942 19068
rect 6998 19022 7050 19068
rect 7106 19022 7158 19068
rect 7214 19022 7266 19068
rect 7322 19022 7374 19068
rect 7430 19022 7482 19068
rect 7538 19022 7590 19068
rect 9677 19022 9729 19068
rect 9785 19022 9837 19068
rect 9893 19022 9945 19068
rect 10001 19022 10053 19068
rect 10109 19022 10161 19068
rect 10217 19022 10269 19068
rect 10325 19022 10377 19068
rect 10433 19022 10485 19068
rect 10541 19022 10593 19068
rect 10649 19022 10701 19068
rect 10757 19022 10809 19068
rect 10865 19022 10917 19068
rect 10973 19022 11025 19068
rect 11081 19022 11133 19068
rect 11189 19022 11241 19068
rect 11297 19022 11349 19068
rect 11405 19022 11457 19068
rect 3433 19019 3485 19022
rect 3541 19019 3593 19022
rect 3649 19019 3701 19022
rect 3757 19019 3809 19022
rect 3865 19019 3917 19022
rect 3973 19019 4025 19022
rect 4081 19019 4133 19022
rect 4189 19019 4241 19022
rect 4297 19019 4349 19022
rect 4405 19019 4457 19022
rect 4513 19019 4565 19022
rect 4621 19019 4673 19022
rect 4729 19019 4781 19022
rect 4837 19019 4889 19022
rect 4945 19019 4997 19022
rect 5053 19019 5105 19022
rect 5161 19019 5213 19022
rect 6566 19019 6618 19022
rect 6674 19019 6726 19022
rect 6782 19019 6834 19022
rect 6890 19019 6942 19022
rect 6998 19019 7050 19022
rect 7106 19019 7158 19022
rect 7214 19019 7266 19022
rect 7322 19019 7374 19022
rect 7430 19019 7482 19022
rect 7538 19019 7590 19022
rect 9677 19019 9729 19022
rect 9785 19019 9837 19022
rect 9893 19019 9945 19022
rect 10001 19019 10053 19022
rect 10109 19019 10161 19022
rect 10217 19019 10269 19022
rect 10325 19019 10377 19022
rect 10433 19019 10485 19022
rect 10541 19019 10593 19022
rect 10649 19019 10701 19022
rect 10757 19019 10809 19022
rect 10865 19019 10917 19022
rect 10973 19019 11025 19022
rect 11081 19019 11133 19022
rect 11189 19019 11241 19022
rect 11297 19019 11349 19022
rect 11405 19019 11457 19022
rect 12051 24261 12103 24313
rect 12159 24261 12211 24313
rect 12267 24261 12319 24313
rect 12051 24153 12103 24205
rect 12159 24153 12211 24205
rect 12267 24153 12319 24205
rect 12051 24045 12103 24097
rect 12159 24045 12211 24097
rect 12267 24045 12319 24097
rect 12051 23937 12103 23989
rect 12159 23937 12211 23989
rect 12267 23937 12319 23989
rect 12051 23829 12103 23881
rect 12159 23829 12211 23881
rect 12267 23829 12319 23881
rect 12051 23721 12103 23773
rect 12159 23721 12211 23773
rect 12267 23721 12319 23773
rect 12051 23613 12103 23665
rect 12159 23613 12211 23665
rect 12267 23613 12319 23665
rect 12051 23505 12103 23557
rect 12159 23505 12211 23557
rect 12267 23505 12319 23557
rect 12051 23397 12103 23449
rect 12159 23397 12211 23449
rect 12267 23397 12319 23449
rect 12051 23289 12103 23341
rect 12159 23289 12211 23341
rect 12267 23289 12319 23341
rect 12051 23181 12103 23233
rect 12159 23181 12211 23233
rect 12267 23181 12319 23233
rect 12051 23073 12103 23125
rect 12159 23073 12211 23125
rect 12267 23073 12319 23125
rect 12051 22965 12103 23017
rect 12159 22965 12211 23017
rect 12267 22965 12319 23017
rect 12051 22857 12103 22909
rect 12159 22857 12211 22909
rect 12267 22857 12319 22909
rect 12051 22749 12103 22801
rect 12159 22749 12211 22801
rect 12267 22749 12319 22801
rect 12051 22641 12103 22693
rect 12159 22641 12211 22693
rect 12267 22641 12319 22693
rect 12051 22533 12103 22585
rect 12159 22533 12211 22585
rect 12267 22533 12319 22585
rect 12051 22425 12103 22477
rect 12159 22425 12211 22477
rect 12267 22425 12319 22477
rect 12051 22317 12103 22369
rect 12159 22317 12211 22369
rect 12267 22317 12319 22369
rect 12051 22209 12103 22261
rect 12159 22209 12211 22261
rect 12267 22209 12319 22261
rect 12051 22101 12103 22153
rect 12159 22101 12211 22153
rect 12267 22101 12319 22153
rect 12051 21993 12103 22045
rect 12159 21993 12211 22045
rect 12267 21993 12319 22045
rect 12051 21885 12103 21937
rect 12159 21885 12211 21937
rect 12267 21885 12319 21937
rect 12051 21777 12103 21829
rect 12159 21777 12211 21829
rect 12267 21777 12319 21829
rect 12051 21669 12103 21721
rect 12159 21669 12211 21721
rect 12267 21669 12319 21721
rect 12051 21561 12103 21613
rect 12159 21561 12211 21613
rect 12267 21561 12319 21613
rect 12051 21453 12103 21505
rect 12159 21453 12211 21505
rect 12267 21453 12319 21505
rect 12051 21345 12103 21397
rect 12159 21345 12211 21397
rect 12267 21345 12319 21397
rect 12051 21237 12103 21289
rect 12159 21237 12211 21289
rect 12267 21237 12319 21289
rect 12051 21129 12103 21181
rect 12159 21129 12211 21181
rect 12267 21129 12319 21181
rect 12051 21021 12103 21073
rect 12159 21021 12211 21073
rect 12267 21021 12319 21073
rect 12051 20913 12103 20965
rect 12159 20913 12211 20965
rect 12267 20913 12319 20965
rect 12051 20805 12103 20857
rect 12159 20805 12211 20857
rect 12267 20805 12319 20857
rect 12051 20697 12103 20749
rect 12159 20697 12211 20749
rect 12267 20697 12319 20749
rect 12051 20589 12103 20641
rect 12159 20589 12211 20641
rect 12267 20589 12319 20641
rect 12051 20481 12103 20533
rect 12159 20481 12211 20533
rect 12267 20481 12319 20533
rect 12051 20373 12103 20425
rect 12159 20373 12211 20425
rect 12267 20373 12319 20425
rect 12051 20265 12103 20317
rect 12159 20265 12211 20317
rect 12267 20265 12319 20317
rect 12051 20157 12103 20209
rect 12159 20157 12211 20209
rect 12267 20157 12319 20209
rect 12051 20049 12103 20101
rect 12159 20049 12211 20101
rect 12267 20049 12319 20101
rect 12051 19941 12103 19993
rect 12159 19941 12211 19993
rect 12267 19941 12319 19993
rect 12051 19833 12103 19885
rect 12159 19833 12211 19885
rect 12267 19833 12319 19885
rect 12051 19725 12103 19777
rect 12159 19725 12211 19777
rect 12267 19725 12319 19777
rect 12051 19617 12103 19669
rect 12159 19617 12211 19669
rect 12267 19617 12319 19669
rect 12051 19509 12103 19561
rect 12159 19509 12211 19561
rect 12267 19509 12319 19561
rect 12051 19401 12103 19453
rect 12159 19401 12211 19453
rect 12267 19401 12319 19453
rect 12051 19293 12103 19345
rect 12159 19293 12211 19345
rect 12267 19293 12319 19345
rect 12051 19185 12103 19237
rect 12159 19185 12211 19237
rect 12267 19185 12319 19237
rect 12051 19077 12103 19129
rect 12159 19077 12211 19129
rect 12267 19077 12319 19129
rect 12051 18969 12103 19021
rect 12159 18969 12211 19021
rect 12267 18969 12319 19021
rect 12051 18861 12103 18913
rect 12159 18861 12211 18913
rect 12267 18861 12319 18913
rect 12051 18753 12103 18805
rect 12159 18753 12211 18805
rect 12267 18753 12319 18805
rect 12051 18645 12103 18697
rect 12159 18645 12211 18697
rect 12267 18645 12319 18697
rect 1505 18622 1557 18629
rect 1613 18622 1665 18629
rect 1721 18622 1773 18629
rect 1829 18622 1881 18629
rect 1937 18622 1989 18629
rect 2045 18622 2097 18629
rect 2153 18622 2205 18629
rect 2261 18622 2313 18629
rect 2369 18622 2421 18629
rect 2477 18622 2529 18629
rect 2585 18622 2637 18629
rect 2693 18622 2745 18629
rect 2801 18622 2853 18629
rect 2909 18622 2961 18629
rect 3017 18622 3069 18629
rect 3125 18622 3177 18629
rect 3233 18622 3285 18629
rect 5372 18622 5424 18629
rect 5480 18622 5532 18629
rect 5588 18622 5640 18629
rect 5696 18622 5748 18629
rect 5804 18622 5856 18629
rect 5912 18622 5964 18629
rect 6020 18622 6072 18629
rect 6128 18622 6180 18629
rect 6236 18622 6288 18629
rect 6344 18622 6396 18629
rect 7749 18622 7801 18629
rect 7857 18622 7909 18629
rect 7965 18622 8017 18629
rect 8073 18622 8125 18629
rect 8181 18622 8233 18629
rect 8289 18622 8341 18629
rect 8397 18622 8449 18629
rect 8505 18622 8557 18629
rect 8613 18622 8665 18629
rect 8721 18622 8773 18629
rect 8829 18622 8881 18629
rect 8937 18622 8989 18629
rect 9045 18622 9097 18629
rect 9153 18622 9205 18629
rect 9261 18622 9313 18629
rect 9369 18622 9421 18629
rect 9477 18622 9529 18629
rect 1505 18577 1557 18622
rect 1613 18577 1665 18622
rect 1721 18577 1773 18622
rect 1829 18577 1881 18622
rect 1937 18577 1989 18622
rect 2045 18577 2097 18622
rect 2153 18577 2205 18622
rect 2261 18577 2313 18622
rect 2369 18577 2421 18622
rect 2477 18577 2529 18622
rect 2585 18577 2637 18622
rect 2693 18577 2745 18622
rect 2801 18577 2853 18622
rect 2909 18577 2961 18622
rect 3017 18577 3069 18622
rect 3125 18577 3177 18622
rect 3233 18577 3285 18622
rect 5372 18577 5424 18622
rect 5480 18577 5532 18622
rect 5588 18577 5640 18622
rect 5696 18577 5748 18622
rect 5804 18577 5856 18622
rect 5912 18577 5964 18622
rect 6020 18577 6072 18622
rect 6128 18577 6180 18622
rect 6236 18577 6288 18622
rect 6344 18577 6396 18622
rect 7749 18577 7801 18622
rect 7857 18577 7909 18622
rect 7965 18577 8017 18622
rect 8073 18577 8125 18622
rect 8181 18577 8233 18622
rect 8289 18577 8341 18622
rect 8397 18577 8449 18622
rect 8505 18577 8557 18622
rect 8613 18577 8665 18622
rect 8721 18577 8773 18622
rect 8829 18577 8881 18622
rect 8937 18577 8989 18622
rect 9045 18577 9097 18622
rect 9153 18577 9205 18622
rect 9261 18577 9313 18622
rect 9369 18577 9421 18622
rect 9477 18577 9529 18622
rect 1505 18476 1557 18521
rect 1613 18476 1665 18521
rect 1721 18476 1773 18521
rect 1829 18476 1881 18521
rect 1937 18476 1989 18521
rect 2045 18476 2097 18521
rect 2153 18476 2205 18521
rect 2261 18476 2313 18521
rect 2369 18476 2421 18521
rect 2477 18476 2529 18521
rect 2585 18476 2637 18521
rect 2693 18476 2745 18521
rect 2801 18476 2853 18521
rect 2909 18476 2961 18521
rect 3017 18476 3069 18521
rect 3125 18476 3177 18521
rect 3233 18476 3285 18521
rect 5372 18476 5424 18521
rect 5480 18476 5532 18521
rect 5588 18476 5640 18521
rect 5696 18476 5748 18521
rect 5804 18476 5856 18521
rect 5912 18476 5964 18521
rect 6020 18476 6072 18521
rect 6128 18476 6180 18521
rect 6236 18476 6288 18521
rect 6344 18476 6396 18521
rect 7749 18476 7801 18521
rect 7857 18476 7909 18521
rect 7965 18476 8017 18521
rect 8073 18476 8125 18521
rect 8181 18476 8233 18521
rect 8289 18476 8341 18521
rect 8397 18476 8449 18521
rect 8505 18476 8557 18521
rect 8613 18476 8665 18521
rect 8721 18476 8773 18521
rect 8829 18476 8881 18521
rect 8937 18476 8989 18521
rect 9045 18476 9097 18521
rect 9153 18476 9205 18521
rect 9261 18476 9313 18521
rect 9369 18476 9421 18521
rect 9477 18476 9529 18521
rect 12051 18537 12103 18589
rect 12159 18537 12211 18589
rect 12267 18537 12319 18589
rect 1505 18469 1557 18476
rect 1613 18469 1665 18476
rect 1721 18469 1773 18476
rect 1829 18469 1881 18476
rect 1937 18469 1989 18476
rect 2045 18469 2097 18476
rect 2153 18469 2205 18476
rect 2261 18469 2313 18476
rect 2369 18469 2421 18476
rect 2477 18469 2529 18476
rect 2585 18469 2637 18476
rect 2693 18469 2745 18476
rect 2801 18469 2853 18476
rect 2909 18469 2961 18476
rect 3017 18469 3069 18476
rect 3125 18469 3177 18476
rect 3233 18469 3285 18476
rect 5372 18469 5424 18476
rect 5480 18469 5532 18476
rect 5588 18469 5640 18476
rect 5696 18469 5748 18476
rect 5804 18469 5856 18476
rect 5912 18469 5964 18476
rect 6020 18469 6072 18476
rect 6128 18469 6180 18476
rect 6236 18469 6288 18476
rect 6344 18469 6396 18476
rect 7749 18469 7801 18476
rect 7857 18469 7909 18476
rect 7965 18469 8017 18476
rect 8073 18469 8125 18476
rect 8181 18469 8233 18476
rect 8289 18469 8341 18476
rect 8397 18469 8449 18476
rect 8505 18469 8557 18476
rect 8613 18469 8665 18476
rect 8721 18469 8773 18476
rect 8829 18469 8881 18476
rect 8937 18469 8989 18476
rect 9045 18469 9097 18476
rect 9153 18469 9205 18476
rect 9261 18469 9313 18476
rect 9369 18469 9421 18476
rect 9477 18469 9529 18476
rect 3433 18076 3485 18079
rect 3541 18076 3593 18079
rect 3649 18076 3701 18079
rect 3757 18076 3809 18079
rect 3865 18076 3917 18079
rect 3973 18076 4025 18079
rect 4081 18076 4133 18079
rect 4189 18076 4241 18079
rect 4297 18076 4349 18079
rect 4405 18076 4457 18079
rect 4513 18076 4565 18079
rect 4621 18076 4673 18079
rect 4729 18076 4781 18079
rect 4837 18076 4889 18079
rect 4945 18076 4997 18079
rect 5053 18076 5105 18079
rect 5161 18076 5213 18079
rect 6566 18076 6618 18079
rect 6674 18076 6726 18079
rect 6782 18076 6834 18079
rect 6890 18076 6942 18079
rect 6998 18076 7050 18079
rect 7106 18076 7158 18079
rect 7214 18076 7266 18079
rect 7322 18076 7374 18079
rect 7430 18076 7482 18079
rect 7538 18076 7590 18079
rect 9677 18076 9729 18079
rect 9785 18076 9837 18079
rect 9893 18076 9945 18079
rect 10001 18076 10053 18079
rect 10109 18076 10161 18079
rect 10217 18076 10269 18079
rect 10325 18076 10377 18079
rect 10433 18076 10485 18079
rect 10541 18076 10593 18079
rect 10649 18076 10701 18079
rect 10757 18076 10809 18079
rect 10865 18076 10917 18079
rect 10973 18076 11025 18079
rect 11081 18076 11133 18079
rect 11189 18076 11241 18079
rect 11297 18076 11349 18079
rect 11405 18076 11457 18079
rect 3433 18030 3485 18076
rect 3541 18030 3593 18076
rect 3649 18030 3701 18076
rect 3757 18030 3809 18076
rect 3865 18030 3917 18076
rect 3973 18030 4025 18076
rect 4081 18030 4133 18076
rect 4189 18030 4241 18076
rect 4297 18030 4349 18076
rect 4405 18030 4457 18076
rect 4513 18030 4565 18076
rect 4621 18030 4673 18076
rect 4729 18030 4781 18076
rect 4837 18030 4889 18076
rect 4945 18030 4997 18076
rect 5053 18030 5105 18076
rect 5161 18030 5213 18076
rect 6566 18030 6618 18076
rect 6674 18030 6726 18076
rect 6782 18030 6834 18076
rect 6890 18030 6942 18076
rect 6998 18030 7050 18076
rect 7106 18030 7158 18076
rect 7214 18030 7266 18076
rect 7322 18030 7374 18076
rect 7430 18030 7482 18076
rect 7538 18030 7590 18076
rect 9677 18030 9729 18076
rect 9785 18030 9837 18076
rect 9893 18030 9945 18076
rect 10001 18030 10053 18076
rect 10109 18030 10161 18076
rect 10217 18030 10269 18076
rect 10325 18030 10377 18076
rect 10433 18030 10485 18076
rect 10541 18030 10593 18076
rect 10649 18030 10701 18076
rect 10757 18030 10809 18076
rect 10865 18030 10917 18076
rect 10973 18030 11025 18076
rect 11081 18030 11133 18076
rect 11189 18030 11241 18076
rect 11297 18030 11349 18076
rect 11405 18030 11457 18076
rect 3433 18027 3485 18030
rect 3541 18027 3593 18030
rect 3649 18027 3701 18030
rect 3757 18027 3809 18030
rect 3865 18027 3917 18030
rect 3973 18027 4025 18030
rect 4081 18027 4133 18030
rect 4189 18027 4241 18030
rect 4297 18027 4349 18030
rect 4405 18027 4457 18030
rect 4513 18027 4565 18030
rect 4621 18027 4673 18030
rect 4729 18027 4781 18030
rect 4837 18027 4889 18030
rect 4945 18027 4997 18030
rect 5053 18027 5105 18030
rect 5161 18027 5213 18030
rect 6566 18027 6618 18030
rect 6674 18027 6726 18030
rect 6782 18027 6834 18030
rect 6890 18027 6942 18030
rect 6998 18027 7050 18030
rect 7106 18027 7158 18030
rect 7214 18027 7266 18030
rect 7322 18027 7374 18030
rect 7430 18027 7482 18030
rect 7538 18027 7590 18030
rect 9677 18027 9729 18030
rect 9785 18027 9837 18030
rect 9893 18027 9945 18030
rect 10001 18027 10053 18030
rect 10109 18027 10161 18030
rect 10217 18027 10269 18030
rect 10325 18027 10377 18030
rect 10433 18027 10485 18030
rect 10541 18027 10593 18030
rect 10649 18027 10701 18030
rect 10757 18027 10809 18030
rect 10865 18027 10917 18030
rect 10973 18027 11025 18030
rect 11081 18027 11133 18030
rect 11189 18027 11241 18030
rect 11297 18027 11349 18030
rect 11405 18027 11457 18030
rect 1233 17963 1285 18015
rect 1341 17963 1393 18015
rect 1233 17855 1256 17907
rect 1256 17855 1285 17907
rect 1341 17855 1393 17907
rect 1233 17747 1256 17799
rect 1256 17747 1285 17799
rect 1341 17747 1393 17799
rect 1233 17639 1256 17691
rect 1256 17639 1285 17691
rect 1341 17639 1393 17691
rect 1233 17531 1256 17583
rect 1256 17531 1285 17583
rect 1341 17531 1393 17583
rect 1233 17423 1256 17475
rect 1256 17423 1285 17475
rect 1341 17423 1393 17475
rect 1233 17315 1256 17367
rect 1256 17315 1285 17367
rect 1341 17315 1393 17367
rect 1233 17207 1256 17259
rect 1256 17207 1285 17259
rect 1341 17207 1393 17259
rect 1233 17099 1256 17151
rect 1256 17099 1285 17151
rect 1341 17099 1393 17151
rect 1233 16991 1256 17043
rect 1256 16991 1285 17043
rect 1341 16991 1393 17043
rect 1233 16883 1256 16935
rect 1256 16883 1285 16935
rect 1341 16883 1393 16935
rect 1233 16775 1256 16827
rect 1256 16775 1285 16827
rect 1341 16775 1393 16827
rect 1233 16667 1256 16719
rect 1256 16667 1285 16719
rect 1341 16667 1393 16719
rect 1233 16559 1256 16611
rect 1256 16559 1285 16611
rect 1341 16559 1393 16611
rect 1233 16451 1256 16503
rect 1256 16451 1285 16503
rect 1341 16451 1393 16503
rect 1233 16343 1256 16395
rect 1256 16343 1285 16395
rect 1341 16343 1393 16395
rect 1233 16235 1256 16287
rect 1256 16235 1285 16287
rect 1341 16235 1393 16287
rect 1233 16127 1256 16179
rect 1256 16127 1285 16179
rect 1341 16127 1393 16179
rect 1233 16019 1256 16071
rect 1256 16019 1285 16071
rect 1341 16019 1393 16071
rect 1233 15911 1256 15963
rect 1256 15911 1285 15963
rect 1341 15911 1393 15963
rect 1233 15803 1256 15855
rect 1256 15803 1285 15855
rect 1341 15803 1393 15855
rect 1233 15695 1256 15747
rect 1256 15695 1285 15747
rect 1341 15695 1393 15747
rect 1233 15587 1256 15639
rect 1256 15587 1285 15639
rect 1341 15587 1393 15639
rect 1233 15479 1256 15531
rect 1256 15479 1285 15531
rect 1341 15479 1393 15531
rect 1233 15371 1256 15423
rect 1256 15371 1285 15423
rect 1341 15371 1393 15423
rect 1233 15263 1256 15315
rect 1256 15263 1285 15315
rect 1341 15263 1393 15315
rect 1233 15155 1256 15207
rect 1256 15155 1285 15207
rect 1341 15155 1393 15207
rect 1233 15047 1256 15099
rect 1256 15047 1285 15099
rect 1341 15047 1393 15099
rect 1233 14939 1256 14991
rect 1256 14939 1285 14991
rect 1341 14939 1393 14991
rect 1233 14831 1256 14883
rect 1256 14831 1285 14883
rect 1341 14831 1393 14883
rect 1233 14723 1256 14775
rect 1256 14723 1285 14775
rect 1341 14723 1393 14775
rect 1233 14615 1256 14667
rect 1256 14615 1285 14667
rect 1341 14615 1393 14667
rect 1233 14507 1256 14559
rect 1256 14507 1285 14559
rect 1341 14507 1393 14559
rect 1233 14399 1256 14451
rect 1256 14399 1285 14451
rect 1341 14399 1393 14451
rect 1233 14291 1256 14343
rect 1256 14291 1285 14343
rect 1341 14291 1393 14343
rect 1233 14183 1256 14235
rect 1256 14183 1285 14235
rect 1341 14183 1393 14235
rect 1233 14075 1256 14127
rect 1256 14075 1285 14127
rect 1341 14075 1393 14127
rect 1233 13967 1256 14019
rect 1256 13967 1285 14019
rect 1341 13967 1393 14019
rect 1233 13859 1256 13911
rect 1256 13859 1285 13911
rect 1341 13859 1393 13911
rect 1233 13751 1256 13803
rect 1256 13751 1285 13803
rect 1341 13751 1393 13803
rect 1233 13643 1256 13695
rect 1256 13643 1285 13695
rect 1341 13643 1393 13695
rect 1233 13535 1256 13587
rect 1256 13535 1285 13587
rect 1341 13535 1393 13587
rect 1233 13427 1256 13479
rect 1256 13427 1285 13479
rect 1341 13427 1393 13479
rect 1233 13319 1256 13371
rect 1256 13319 1285 13371
rect 1341 13319 1393 13371
rect 11569 17963 11621 18015
rect 11677 17963 11729 18015
rect 1505 17832 1557 17835
rect 1613 17832 1665 17835
rect 1721 17832 1773 17835
rect 1829 17832 1881 17835
rect 1937 17832 1989 17835
rect 2045 17832 2097 17835
rect 2153 17832 2205 17835
rect 2261 17832 2313 17835
rect 2369 17832 2421 17835
rect 2477 17832 2529 17835
rect 2585 17832 2637 17835
rect 2693 17832 2745 17835
rect 2801 17832 2853 17835
rect 2909 17832 2961 17835
rect 3017 17832 3069 17835
rect 3125 17832 3177 17835
rect 3233 17832 3285 17835
rect 5372 17832 5424 17835
rect 5480 17832 5532 17835
rect 5588 17832 5640 17835
rect 5696 17832 5748 17835
rect 5804 17832 5856 17835
rect 5912 17832 5964 17835
rect 6020 17832 6072 17835
rect 6128 17832 6180 17835
rect 6236 17832 6288 17835
rect 6344 17832 6396 17835
rect 7749 17832 7801 17835
rect 7857 17832 7909 17835
rect 7965 17832 8017 17835
rect 8073 17832 8125 17835
rect 8181 17832 8233 17835
rect 8289 17832 8341 17835
rect 8397 17832 8449 17835
rect 8505 17832 8557 17835
rect 8613 17832 8665 17835
rect 8721 17832 8773 17835
rect 8829 17832 8881 17835
rect 8937 17832 8989 17835
rect 9045 17832 9097 17835
rect 9153 17832 9205 17835
rect 9261 17832 9313 17835
rect 9369 17832 9421 17835
rect 9477 17832 9529 17835
rect 1505 17786 1557 17832
rect 1613 17786 1665 17832
rect 1721 17786 1773 17832
rect 1829 17786 1881 17832
rect 1937 17786 1989 17832
rect 2045 17786 2097 17832
rect 2153 17786 2205 17832
rect 2261 17786 2313 17832
rect 2369 17786 2421 17832
rect 2477 17786 2529 17832
rect 2585 17786 2637 17832
rect 2693 17786 2745 17832
rect 2801 17786 2853 17832
rect 2909 17786 2961 17832
rect 3017 17786 3069 17832
rect 3125 17786 3177 17832
rect 3233 17786 3285 17832
rect 5372 17786 5424 17832
rect 5480 17786 5532 17832
rect 5588 17786 5640 17832
rect 5696 17786 5748 17832
rect 5804 17786 5856 17832
rect 5912 17786 5964 17832
rect 6020 17786 6072 17832
rect 6128 17786 6180 17832
rect 6236 17786 6288 17832
rect 6344 17786 6396 17832
rect 7749 17786 7801 17832
rect 7857 17786 7909 17832
rect 7965 17786 8017 17832
rect 8073 17786 8125 17832
rect 8181 17786 8233 17832
rect 8289 17786 8341 17832
rect 8397 17786 8449 17832
rect 8505 17786 8557 17832
rect 8613 17786 8665 17832
rect 8721 17786 8773 17832
rect 8829 17786 8881 17832
rect 8937 17786 8989 17832
rect 9045 17786 9097 17832
rect 9153 17786 9205 17832
rect 9261 17786 9313 17832
rect 9369 17786 9421 17832
rect 9477 17786 9529 17832
rect 1505 17783 1557 17786
rect 1613 17783 1665 17786
rect 1721 17783 1773 17786
rect 1829 17783 1881 17786
rect 1937 17783 1989 17786
rect 2045 17783 2097 17786
rect 2153 17783 2205 17786
rect 2261 17783 2313 17786
rect 2369 17783 2421 17786
rect 2477 17783 2529 17786
rect 2585 17783 2637 17786
rect 2693 17783 2745 17786
rect 2801 17783 2853 17786
rect 2909 17783 2961 17786
rect 3017 17783 3069 17786
rect 3125 17783 3177 17786
rect 3233 17783 3285 17786
rect 5372 17783 5424 17786
rect 5480 17783 5532 17786
rect 5588 17783 5640 17786
rect 5696 17783 5748 17786
rect 5804 17783 5856 17786
rect 5912 17783 5964 17786
rect 6020 17783 6072 17786
rect 6128 17783 6180 17786
rect 6236 17783 6288 17786
rect 6344 17783 6396 17786
rect 7749 17783 7801 17786
rect 7857 17783 7909 17786
rect 7965 17783 8017 17786
rect 8073 17783 8125 17786
rect 8181 17783 8233 17786
rect 8289 17783 8341 17786
rect 8397 17783 8449 17786
rect 8505 17783 8557 17786
rect 8613 17783 8665 17786
rect 8721 17783 8773 17786
rect 8829 17783 8881 17786
rect 8937 17783 8989 17786
rect 9045 17783 9097 17786
rect 9153 17783 9205 17786
rect 9261 17783 9313 17786
rect 9369 17783 9421 17786
rect 9477 17783 9529 17786
rect 3433 17588 3485 17591
rect 3541 17588 3593 17591
rect 3649 17588 3701 17591
rect 3757 17588 3809 17591
rect 3865 17588 3917 17591
rect 3973 17588 4025 17591
rect 4081 17588 4133 17591
rect 4189 17588 4241 17591
rect 4297 17588 4349 17591
rect 4405 17588 4457 17591
rect 4513 17588 4565 17591
rect 4621 17588 4673 17591
rect 4729 17588 4781 17591
rect 4837 17588 4889 17591
rect 4945 17588 4997 17591
rect 5053 17588 5105 17591
rect 5161 17588 5213 17591
rect 6566 17588 6618 17591
rect 6674 17588 6726 17591
rect 6782 17588 6834 17591
rect 6890 17588 6942 17591
rect 6998 17588 7050 17591
rect 7106 17588 7158 17591
rect 7214 17588 7266 17591
rect 7322 17588 7374 17591
rect 7430 17588 7482 17591
rect 7538 17588 7590 17591
rect 9677 17588 9729 17591
rect 9785 17588 9837 17591
rect 9893 17588 9945 17591
rect 10001 17588 10053 17591
rect 10109 17588 10161 17591
rect 10217 17588 10269 17591
rect 10325 17588 10377 17591
rect 10433 17588 10485 17591
rect 10541 17588 10593 17591
rect 10649 17588 10701 17591
rect 10757 17588 10809 17591
rect 10865 17588 10917 17591
rect 10973 17588 11025 17591
rect 11081 17588 11133 17591
rect 11189 17588 11241 17591
rect 11297 17588 11349 17591
rect 11405 17588 11457 17591
rect 3433 17542 3485 17588
rect 3541 17542 3593 17588
rect 3649 17542 3701 17588
rect 3757 17542 3809 17588
rect 3865 17542 3917 17588
rect 3973 17542 4025 17588
rect 4081 17542 4133 17588
rect 4189 17542 4241 17588
rect 4297 17542 4349 17588
rect 4405 17542 4457 17588
rect 4513 17542 4565 17588
rect 4621 17542 4673 17588
rect 4729 17542 4781 17588
rect 4837 17542 4889 17588
rect 4945 17542 4997 17588
rect 5053 17542 5105 17588
rect 5161 17542 5213 17588
rect 6566 17542 6618 17588
rect 6674 17542 6726 17588
rect 6782 17542 6834 17588
rect 6890 17542 6942 17588
rect 6998 17542 7050 17588
rect 7106 17542 7158 17588
rect 7214 17542 7266 17588
rect 7322 17542 7374 17588
rect 7430 17542 7482 17588
rect 7538 17542 7590 17588
rect 9677 17542 9729 17588
rect 9785 17542 9837 17588
rect 9893 17542 9945 17588
rect 10001 17542 10053 17588
rect 10109 17542 10161 17588
rect 10217 17542 10269 17588
rect 10325 17542 10377 17588
rect 10433 17542 10485 17588
rect 10541 17542 10593 17588
rect 10649 17542 10701 17588
rect 10757 17542 10809 17588
rect 10865 17542 10917 17588
rect 10973 17542 11025 17588
rect 11081 17542 11133 17588
rect 11189 17542 11241 17588
rect 11297 17542 11349 17588
rect 11405 17542 11457 17588
rect 3433 17539 3485 17542
rect 3541 17539 3593 17542
rect 3649 17539 3701 17542
rect 3757 17539 3809 17542
rect 3865 17539 3917 17542
rect 3973 17539 4025 17542
rect 4081 17539 4133 17542
rect 4189 17539 4241 17542
rect 4297 17539 4349 17542
rect 4405 17539 4457 17542
rect 4513 17539 4565 17542
rect 4621 17539 4673 17542
rect 4729 17539 4781 17542
rect 4837 17539 4889 17542
rect 4945 17539 4997 17542
rect 5053 17539 5105 17542
rect 5161 17539 5213 17542
rect 6566 17539 6618 17542
rect 6674 17539 6726 17542
rect 6782 17539 6834 17542
rect 6890 17539 6942 17542
rect 6998 17539 7050 17542
rect 7106 17539 7158 17542
rect 7214 17539 7266 17542
rect 7322 17539 7374 17542
rect 7430 17539 7482 17542
rect 7538 17539 7590 17542
rect 9677 17539 9729 17542
rect 9785 17539 9837 17542
rect 9893 17539 9945 17542
rect 10001 17539 10053 17542
rect 10109 17539 10161 17542
rect 10217 17539 10269 17542
rect 10325 17539 10377 17542
rect 10433 17539 10485 17542
rect 10541 17539 10593 17542
rect 10649 17539 10701 17542
rect 10757 17539 10809 17542
rect 10865 17539 10917 17542
rect 10973 17539 11025 17542
rect 11081 17539 11133 17542
rect 11189 17539 11241 17542
rect 11297 17539 11349 17542
rect 11405 17539 11457 17542
rect 1505 17344 1557 17347
rect 1613 17344 1665 17347
rect 1721 17344 1773 17347
rect 1829 17344 1881 17347
rect 1937 17344 1989 17347
rect 2045 17344 2097 17347
rect 2153 17344 2205 17347
rect 2261 17344 2313 17347
rect 2369 17344 2421 17347
rect 2477 17344 2529 17347
rect 2585 17344 2637 17347
rect 2693 17344 2745 17347
rect 2801 17344 2853 17347
rect 2909 17344 2961 17347
rect 3017 17344 3069 17347
rect 3125 17344 3177 17347
rect 3233 17344 3285 17347
rect 5372 17344 5424 17347
rect 5480 17344 5532 17347
rect 5588 17344 5640 17347
rect 5696 17344 5748 17347
rect 5804 17344 5856 17347
rect 5912 17344 5964 17347
rect 6020 17344 6072 17347
rect 6128 17344 6180 17347
rect 6236 17344 6288 17347
rect 6344 17344 6396 17347
rect 7749 17344 7801 17347
rect 7857 17344 7909 17347
rect 7965 17344 8017 17347
rect 8073 17344 8125 17347
rect 8181 17344 8233 17347
rect 8289 17344 8341 17347
rect 8397 17344 8449 17347
rect 8505 17344 8557 17347
rect 8613 17344 8665 17347
rect 8721 17344 8773 17347
rect 8829 17344 8881 17347
rect 8937 17344 8989 17347
rect 9045 17344 9097 17347
rect 9153 17344 9205 17347
rect 9261 17344 9313 17347
rect 9369 17344 9421 17347
rect 9477 17344 9529 17347
rect 1505 17298 1557 17344
rect 1613 17298 1665 17344
rect 1721 17298 1773 17344
rect 1829 17298 1881 17344
rect 1937 17298 1989 17344
rect 2045 17298 2097 17344
rect 2153 17298 2205 17344
rect 2261 17298 2313 17344
rect 2369 17298 2421 17344
rect 2477 17298 2529 17344
rect 2585 17298 2637 17344
rect 2693 17298 2745 17344
rect 2801 17298 2853 17344
rect 2909 17298 2961 17344
rect 3017 17298 3069 17344
rect 3125 17298 3177 17344
rect 3233 17298 3285 17344
rect 5372 17298 5424 17344
rect 5480 17298 5532 17344
rect 5588 17298 5640 17344
rect 5696 17298 5748 17344
rect 5804 17298 5856 17344
rect 5912 17298 5964 17344
rect 6020 17298 6072 17344
rect 6128 17298 6180 17344
rect 6236 17298 6288 17344
rect 6344 17298 6396 17344
rect 7749 17298 7801 17344
rect 7857 17298 7909 17344
rect 7965 17298 8017 17344
rect 8073 17298 8125 17344
rect 8181 17298 8233 17344
rect 8289 17298 8341 17344
rect 8397 17298 8449 17344
rect 8505 17298 8557 17344
rect 8613 17298 8665 17344
rect 8721 17298 8773 17344
rect 8829 17298 8881 17344
rect 8937 17298 8989 17344
rect 9045 17298 9097 17344
rect 9153 17298 9205 17344
rect 9261 17298 9313 17344
rect 9369 17298 9421 17344
rect 9477 17298 9529 17344
rect 1505 17295 1557 17298
rect 1613 17295 1665 17298
rect 1721 17295 1773 17298
rect 1829 17295 1881 17298
rect 1937 17295 1989 17298
rect 2045 17295 2097 17298
rect 2153 17295 2205 17298
rect 2261 17295 2313 17298
rect 2369 17295 2421 17298
rect 2477 17295 2529 17298
rect 2585 17295 2637 17298
rect 2693 17295 2745 17298
rect 2801 17295 2853 17298
rect 2909 17295 2961 17298
rect 3017 17295 3069 17298
rect 3125 17295 3177 17298
rect 3233 17295 3285 17298
rect 5372 17295 5424 17298
rect 5480 17295 5532 17298
rect 5588 17295 5640 17298
rect 5696 17295 5748 17298
rect 5804 17295 5856 17298
rect 5912 17295 5964 17298
rect 6020 17295 6072 17298
rect 6128 17295 6180 17298
rect 6236 17295 6288 17298
rect 6344 17295 6396 17298
rect 7749 17295 7801 17298
rect 7857 17295 7909 17298
rect 7965 17295 8017 17298
rect 8073 17295 8125 17298
rect 8181 17295 8233 17298
rect 8289 17295 8341 17298
rect 8397 17295 8449 17298
rect 8505 17295 8557 17298
rect 8613 17295 8665 17298
rect 8721 17295 8773 17298
rect 8829 17295 8881 17298
rect 8937 17295 8989 17298
rect 9045 17295 9097 17298
rect 9153 17295 9205 17298
rect 9261 17295 9313 17298
rect 9369 17295 9421 17298
rect 9477 17295 9529 17298
rect 3433 17100 3485 17103
rect 3541 17100 3593 17103
rect 3649 17100 3701 17103
rect 3757 17100 3809 17103
rect 3865 17100 3917 17103
rect 3973 17100 4025 17103
rect 4081 17100 4133 17103
rect 4189 17100 4241 17103
rect 4297 17100 4349 17103
rect 4405 17100 4457 17103
rect 4513 17100 4565 17103
rect 4621 17100 4673 17103
rect 4729 17100 4781 17103
rect 4837 17100 4889 17103
rect 4945 17100 4997 17103
rect 5053 17100 5105 17103
rect 5161 17100 5213 17103
rect 6566 17100 6618 17103
rect 6674 17100 6726 17103
rect 6782 17100 6834 17103
rect 6890 17100 6942 17103
rect 6998 17100 7050 17103
rect 7106 17100 7158 17103
rect 7214 17100 7266 17103
rect 7322 17100 7374 17103
rect 7430 17100 7482 17103
rect 7538 17100 7590 17103
rect 9677 17100 9729 17103
rect 9785 17100 9837 17103
rect 9893 17100 9945 17103
rect 10001 17100 10053 17103
rect 10109 17100 10161 17103
rect 10217 17100 10269 17103
rect 10325 17100 10377 17103
rect 10433 17100 10485 17103
rect 10541 17100 10593 17103
rect 10649 17100 10701 17103
rect 10757 17100 10809 17103
rect 10865 17100 10917 17103
rect 10973 17100 11025 17103
rect 11081 17100 11133 17103
rect 11189 17100 11241 17103
rect 11297 17100 11349 17103
rect 11405 17100 11457 17103
rect 3433 17054 3485 17100
rect 3541 17054 3593 17100
rect 3649 17054 3701 17100
rect 3757 17054 3809 17100
rect 3865 17054 3917 17100
rect 3973 17054 4025 17100
rect 4081 17054 4133 17100
rect 4189 17054 4241 17100
rect 4297 17054 4349 17100
rect 4405 17054 4457 17100
rect 4513 17054 4565 17100
rect 4621 17054 4673 17100
rect 4729 17054 4781 17100
rect 4837 17054 4889 17100
rect 4945 17054 4997 17100
rect 5053 17054 5105 17100
rect 5161 17054 5213 17100
rect 6566 17054 6618 17100
rect 6674 17054 6726 17100
rect 6782 17054 6834 17100
rect 6890 17054 6942 17100
rect 6998 17054 7050 17100
rect 7106 17054 7158 17100
rect 7214 17054 7266 17100
rect 7322 17054 7374 17100
rect 7430 17054 7482 17100
rect 7538 17054 7590 17100
rect 9677 17054 9729 17100
rect 9785 17054 9837 17100
rect 9893 17054 9945 17100
rect 10001 17054 10053 17100
rect 10109 17054 10161 17100
rect 10217 17054 10269 17100
rect 10325 17054 10377 17100
rect 10433 17054 10485 17100
rect 10541 17054 10593 17100
rect 10649 17054 10701 17100
rect 10757 17054 10809 17100
rect 10865 17054 10917 17100
rect 10973 17054 11025 17100
rect 11081 17054 11133 17100
rect 11189 17054 11241 17100
rect 11297 17054 11349 17100
rect 11405 17054 11457 17100
rect 3433 17051 3485 17054
rect 3541 17051 3593 17054
rect 3649 17051 3701 17054
rect 3757 17051 3809 17054
rect 3865 17051 3917 17054
rect 3973 17051 4025 17054
rect 4081 17051 4133 17054
rect 4189 17051 4241 17054
rect 4297 17051 4349 17054
rect 4405 17051 4457 17054
rect 4513 17051 4565 17054
rect 4621 17051 4673 17054
rect 4729 17051 4781 17054
rect 4837 17051 4889 17054
rect 4945 17051 4997 17054
rect 5053 17051 5105 17054
rect 5161 17051 5213 17054
rect 6566 17051 6618 17054
rect 6674 17051 6726 17054
rect 6782 17051 6834 17054
rect 6890 17051 6942 17054
rect 6998 17051 7050 17054
rect 7106 17051 7158 17054
rect 7214 17051 7266 17054
rect 7322 17051 7374 17054
rect 7430 17051 7482 17054
rect 7538 17051 7590 17054
rect 9677 17051 9729 17054
rect 9785 17051 9837 17054
rect 9893 17051 9945 17054
rect 10001 17051 10053 17054
rect 10109 17051 10161 17054
rect 10217 17051 10269 17054
rect 10325 17051 10377 17054
rect 10433 17051 10485 17054
rect 10541 17051 10593 17054
rect 10649 17051 10701 17054
rect 10757 17051 10809 17054
rect 10865 17051 10917 17054
rect 10973 17051 11025 17054
rect 11081 17051 11133 17054
rect 11189 17051 11241 17054
rect 11297 17051 11349 17054
rect 11405 17051 11457 17054
rect 1505 16856 1557 16859
rect 1613 16856 1665 16859
rect 1721 16856 1773 16859
rect 1829 16856 1881 16859
rect 1937 16856 1989 16859
rect 2045 16856 2097 16859
rect 2153 16856 2205 16859
rect 2261 16856 2313 16859
rect 2369 16856 2421 16859
rect 2477 16856 2529 16859
rect 2585 16856 2637 16859
rect 2693 16856 2745 16859
rect 2801 16856 2853 16859
rect 2909 16856 2961 16859
rect 3017 16856 3069 16859
rect 3125 16856 3177 16859
rect 3233 16856 3285 16859
rect 5372 16856 5424 16859
rect 5480 16856 5532 16859
rect 5588 16856 5640 16859
rect 5696 16856 5748 16859
rect 5804 16856 5856 16859
rect 5912 16856 5964 16859
rect 6020 16856 6072 16859
rect 6128 16856 6180 16859
rect 6236 16856 6288 16859
rect 6344 16856 6396 16859
rect 7749 16856 7801 16859
rect 7857 16856 7909 16859
rect 7965 16856 8017 16859
rect 8073 16856 8125 16859
rect 8181 16856 8233 16859
rect 8289 16856 8341 16859
rect 8397 16856 8449 16859
rect 8505 16856 8557 16859
rect 8613 16856 8665 16859
rect 8721 16856 8773 16859
rect 8829 16856 8881 16859
rect 8937 16856 8989 16859
rect 9045 16856 9097 16859
rect 9153 16856 9205 16859
rect 9261 16856 9313 16859
rect 9369 16856 9421 16859
rect 9477 16856 9529 16859
rect 1505 16810 1557 16856
rect 1613 16810 1665 16856
rect 1721 16810 1773 16856
rect 1829 16810 1881 16856
rect 1937 16810 1989 16856
rect 2045 16810 2097 16856
rect 2153 16810 2205 16856
rect 2261 16810 2313 16856
rect 2369 16810 2421 16856
rect 2477 16810 2529 16856
rect 2585 16810 2637 16856
rect 2693 16810 2745 16856
rect 2801 16810 2853 16856
rect 2909 16810 2961 16856
rect 3017 16810 3069 16856
rect 3125 16810 3177 16856
rect 3233 16810 3285 16856
rect 5372 16810 5424 16856
rect 5480 16810 5532 16856
rect 5588 16810 5640 16856
rect 5696 16810 5748 16856
rect 5804 16810 5856 16856
rect 5912 16810 5964 16856
rect 6020 16810 6072 16856
rect 6128 16810 6180 16856
rect 6236 16810 6288 16856
rect 6344 16810 6396 16856
rect 7749 16810 7801 16856
rect 7857 16810 7909 16856
rect 7965 16810 8017 16856
rect 8073 16810 8125 16856
rect 8181 16810 8233 16856
rect 8289 16810 8341 16856
rect 8397 16810 8449 16856
rect 8505 16810 8557 16856
rect 8613 16810 8665 16856
rect 8721 16810 8773 16856
rect 8829 16810 8881 16856
rect 8937 16810 8989 16856
rect 9045 16810 9097 16856
rect 9153 16810 9205 16856
rect 9261 16810 9313 16856
rect 9369 16810 9421 16856
rect 9477 16810 9529 16856
rect 1505 16807 1557 16810
rect 1613 16807 1665 16810
rect 1721 16807 1773 16810
rect 1829 16807 1881 16810
rect 1937 16807 1989 16810
rect 2045 16807 2097 16810
rect 2153 16807 2205 16810
rect 2261 16807 2313 16810
rect 2369 16807 2421 16810
rect 2477 16807 2529 16810
rect 2585 16807 2637 16810
rect 2693 16807 2745 16810
rect 2801 16807 2853 16810
rect 2909 16807 2961 16810
rect 3017 16807 3069 16810
rect 3125 16807 3177 16810
rect 3233 16807 3285 16810
rect 5372 16807 5424 16810
rect 5480 16807 5532 16810
rect 5588 16807 5640 16810
rect 5696 16807 5748 16810
rect 5804 16807 5856 16810
rect 5912 16807 5964 16810
rect 6020 16807 6072 16810
rect 6128 16807 6180 16810
rect 6236 16807 6288 16810
rect 6344 16807 6396 16810
rect 7749 16807 7801 16810
rect 7857 16807 7909 16810
rect 7965 16807 8017 16810
rect 8073 16807 8125 16810
rect 8181 16807 8233 16810
rect 8289 16807 8341 16810
rect 8397 16807 8449 16810
rect 8505 16807 8557 16810
rect 8613 16807 8665 16810
rect 8721 16807 8773 16810
rect 8829 16807 8881 16810
rect 8937 16807 8989 16810
rect 9045 16807 9097 16810
rect 9153 16807 9205 16810
rect 9261 16807 9313 16810
rect 9369 16807 9421 16810
rect 9477 16807 9529 16810
rect 3433 16612 3485 16615
rect 3541 16612 3593 16615
rect 3649 16612 3701 16615
rect 3757 16612 3809 16615
rect 3865 16612 3917 16615
rect 3973 16612 4025 16615
rect 4081 16612 4133 16615
rect 4189 16612 4241 16615
rect 4297 16612 4349 16615
rect 4405 16612 4457 16615
rect 4513 16612 4565 16615
rect 4621 16612 4673 16615
rect 4729 16612 4781 16615
rect 4837 16612 4889 16615
rect 4945 16612 4997 16615
rect 5053 16612 5105 16615
rect 5161 16612 5213 16615
rect 6566 16612 6618 16615
rect 6674 16612 6726 16615
rect 6782 16612 6834 16615
rect 6890 16612 6942 16615
rect 6998 16612 7050 16615
rect 7106 16612 7158 16615
rect 7214 16612 7266 16615
rect 7322 16612 7374 16615
rect 7430 16612 7482 16615
rect 7538 16612 7590 16615
rect 9677 16612 9729 16615
rect 9785 16612 9837 16615
rect 9893 16612 9945 16615
rect 10001 16612 10053 16615
rect 10109 16612 10161 16615
rect 10217 16612 10269 16615
rect 10325 16612 10377 16615
rect 10433 16612 10485 16615
rect 10541 16612 10593 16615
rect 10649 16612 10701 16615
rect 10757 16612 10809 16615
rect 10865 16612 10917 16615
rect 10973 16612 11025 16615
rect 11081 16612 11133 16615
rect 11189 16612 11241 16615
rect 11297 16612 11349 16615
rect 11405 16612 11457 16615
rect 3433 16566 3485 16612
rect 3541 16566 3593 16612
rect 3649 16566 3701 16612
rect 3757 16566 3809 16612
rect 3865 16566 3917 16612
rect 3973 16566 4025 16612
rect 4081 16566 4133 16612
rect 4189 16566 4241 16612
rect 4297 16566 4349 16612
rect 4405 16566 4457 16612
rect 4513 16566 4565 16612
rect 4621 16566 4673 16612
rect 4729 16566 4781 16612
rect 4837 16566 4889 16612
rect 4945 16566 4997 16612
rect 5053 16566 5105 16612
rect 5161 16566 5213 16612
rect 6566 16566 6618 16612
rect 6674 16566 6726 16612
rect 6782 16566 6834 16612
rect 6890 16566 6942 16612
rect 6998 16566 7050 16612
rect 7106 16566 7158 16612
rect 7214 16566 7266 16612
rect 7322 16566 7374 16612
rect 7430 16566 7482 16612
rect 7538 16566 7590 16612
rect 9677 16566 9729 16612
rect 9785 16566 9837 16612
rect 9893 16566 9945 16612
rect 10001 16566 10053 16612
rect 10109 16566 10161 16612
rect 10217 16566 10269 16612
rect 10325 16566 10377 16612
rect 10433 16566 10485 16612
rect 10541 16566 10593 16612
rect 10649 16566 10701 16612
rect 10757 16566 10809 16612
rect 10865 16566 10917 16612
rect 10973 16566 11025 16612
rect 11081 16566 11133 16612
rect 11189 16566 11241 16612
rect 11297 16566 11349 16612
rect 11405 16566 11457 16612
rect 3433 16563 3485 16566
rect 3541 16563 3593 16566
rect 3649 16563 3701 16566
rect 3757 16563 3809 16566
rect 3865 16563 3917 16566
rect 3973 16563 4025 16566
rect 4081 16563 4133 16566
rect 4189 16563 4241 16566
rect 4297 16563 4349 16566
rect 4405 16563 4457 16566
rect 4513 16563 4565 16566
rect 4621 16563 4673 16566
rect 4729 16563 4781 16566
rect 4837 16563 4889 16566
rect 4945 16563 4997 16566
rect 5053 16563 5105 16566
rect 5161 16563 5213 16566
rect 6566 16563 6618 16566
rect 6674 16563 6726 16566
rect 6782 16563 6834 16566
rect 6890 16563 6942 16566
rect 6998 16563 7050 16566
rect 7106 16563 7158 16566
rect 7214 16563 7266 16566
rect 7322 16563 7374 16566
rect 7430 16563 7482 16566
rect 7538 16563 7590 16566
rect 9677 16563 9729 16566
rect 9785 16563 9837 16566
rect 9893 16563 9945 16566
rect 10001 16563 10053 16566
rect 10109 16563 10161 16566
rect 10217 16563 10269 16566
rect 10325 16563 10377 16566
rect 10433 16563 10485 16566
rect 10541 16563 10593 16566
rect 10649 16563 10701 16566
rect 10757 16563 10809 16566
rect 10865 16563 10917 16566
rect 10973 16563 11025 16566
rect 11081 16563 11133 16566
rect 11189 16563 11241 16566
rect 11297 16563 11349 16566
rect 11405 16563 11457 16566
rect 1505 16368 1557 16371
rect 1613 16368 1665 16371
rect 1721 16368 1773 16371
rect 1829 16368 1881 16371
rect 1937 16368 1989 16371
rect 2045 16368 2097 16371
rect 2153 16368 2205 16371
rect 2261 16368 2313 16371
rect 2369 16368 2421 16371
rect 2477 16368 2529 16371
rect 2585 16368 2637 16371
rect 2693 16368 2745 16371
rect 2801 16368 2853 16371
rect 2909 16368 2961 16371
rect 3017 16368 3069 16371
rect 3125 16368 3177 16371
rect 3233 16368 3285 16371
rect 5372 16368 5424 16371
rect 5480 16368 5532 16371
rect 5588 16368 5640 16371
rect 5696 16368 5748 16371
rect 5804 16368 5856 16371
rect 5912 16368 5964 16371
rect 6020 16368 6072 16371
rect 6128 16368 6180 16371
rect 6236 16368 6288 16371
rect 6344 16368 6396 16371
rect 7749 16368 7801 16371
rect 7857 16368 7909 16371
rect 7965 16368 8017 16371
rect 8073 16368 8125 16371
rect 8181 16368 8233 16371
rect 8289 16368 8341 16371
rect 8397 16368 8449 16371
rect 8505 16368 8557 16371
rect 8613 16368 8665 16371
rect 8721 16368 8773 16371
rect 8829 16368 8881 16371
rect 8937 16368 8989 16371
rect 9045 16368 9097 16371
rect 9153 16368 9205 16371
rect 9261 16368 9313 16371
rect 9369 16368 9421 16371
rect 9477 16368 9529 16371
rect 1505 16322 1557 16368
rect 1613 16322 1665 16368
rect 1721 16322 1773 16368
rect 1829 16322 1881 16368
rect 1937 16322 1989 16368
rect 2045 16322 2097 16368
rect 2153 16322 2205 16368
rect 2261 16322 2313 16368
rect 2369 16322 2421 16368
rect 2477 16322 2529 16368
rect 2585 16322 2637 16368
rect 2693 16322 2745 16368
rect 2801 16322 2853 16368
rect 2909 16322 2961 16368
rect 3017 16322 3069 16368
rect 3125 16322 3177 16368
rect 3233 16322 3285 16368
rect 5372 16322 5424 16368
rect 5480 16322 5532 16368
rect 5588 16322 5640 16368
rect 5696 16322 5748 16368
rect 5804 16322 5856 16368
rect 5912 16322 5964 16368
rect 6020 16322 6072 16368
rect 6128 16322 6180 16368
rect 6236 16322 6288 16368
rect 6344 16322 6396 16368
rect 7749 16322 7801 16368
rect 7857 16322 7909 16368
rect 7965 16322 8017 16368
rect 8073 16322 8125 16368
rect 8181 16322 8233 16368
rect 8289 16322 8341 16368
rect 8397 16322 8449 16368
rect 8505 16322 8557 16368
rect 8613 16322 8665 16368
rect 8721 16322 8773 16368
rect 8829 16322 8881 16368
rect 8937 16322 8989 16368
rect 9045 16322 9097 16368
rect 9153 16322 9205 16368
rect 9261 16322 9313 16368
rect 9369 16322 9421 16368
rect 9477 16322 9529 16368
rect 1505 16319 1557 16322
rect 1613 16319 1665 16322
rect 1721 16319 1773 16322
rect 1829 16319 1881 16322
rect 1937 16319 1989 16322
rect 2045 16319 2097 16322
rect 2153 16319 2205 16322
rect 2261 16319 2313 16322
rect 2369 16319 2421 16322
rect 2477 16319 2529 16322
rect 2585 16319 2637 16322
rect 2693 16319 2745 16322
rect 2801 16319 2853 16322
rect 2909 16319 2961 16322
rect 3017 16319 3069 16322
rect 3125 16319 3177 16322
rect 3233 16319 3285 16322
rect 5372 16319 5424 16322
rect 5480 16319 5532 16322
rect 5588 16319 5640 16322
rect 5696 16319 5748 16322
rect 5804 16319 5856 16322
rect 5912 16319 5964 16322
rect 6020 16319 6072 16322
rect 6128 16319 6180 16322
rect 6236 16319 6288 16322
rect 6344 16319 6396 16322
rect 7749 16319 7801 16322
rect 7857 16319 7909 16322
rect 7965 16319 8017 16322
rect 8073 16319 8125 16322
rect 8181 16319 8233 16322
rect 8289 16319 8341 16322
rect 8397 16319 8449 16322
rect 8505 16319 8557 16322
rect 8613 16319 8665 16322
rect 8721 16319 8773 16322
rect 8829 16319 8881 16322
rect 8937 16319 8989 16322
rect 9045 16319 9097 16322
rect 9153 16319 9205 16322
rect 9261 16319 9313 16322
rect 9369 16319 9421 16322
rect 9477 16319 9529 16322
rect 3433 16124 3485 16127
rect 3541 16124 3593 16127
rect 3649 16124 3701 16127
rect 3757 16124 3809 16127
rect 3865 16124 3917 16127
rect 3973 16124 4025 16127
rect 4081 16124 4133 16127
rect 4189 16124 4241 16127
rect 4297 16124 4349 16127
rect 4405 16124 4457 16127
rect 4513 16124 4565 16127
rect 4621 16124 4673 16127
rect 4729 16124 4781 16127
rect 4837 16124 4889 16127
rect 4945 16124 4997 16127
rect 5053 16124 5105 16127
rect 5161 16124 5213 16127
rect 6566 16124 6618 16127
rect 6674 16124 6726 16127
rect 6782 16124 6834 16127
rect 6890 16124 6942 16127
rect 6998 16124 7050 16127
rect 7106 16124 7158 16127
rect 7214 16124 7266 16127
rect 7322 16124 7374 16127
rect 7430 16124 7482 16127
rect 7538 16124 7590 16127
rect 9677 16124 9729 16127
rect 9785 16124 9837 16127
rect 9893 16124 9945 16127
rect 10001 16124 10053 16127
rect 10109 16124 10161 16127
rect 10217 16124 10269 16127
rect 10325 16124 10377 16127
rect 10433 16124 10485 16127
rect 10541 16124 10593 16127
rect 10649 16124 10701 16127
rect 10757 16124 10809 16127
rect 10865 16124 10917 16127
rect 10973 16124 11025 16127
rect 11081 16124 11133 16127
rect 11189 16124 11241 16127
rect 11297 16124 11349 16127
rect 11405 16124 11457 16127
rect 3433 16078 3485 16124
rect 3541 16078 3593 16124
rect 3649 16078 3701 16124
rect 3757 16078 3809 16124
rect 3865 16078 3917 16124
rect 3973 16078 4025 16124
rect 4081 16078 4133 16124
rect 4189 16078 4241 16124
rect 4297 16078 4349 16124
rect 4405 16078 4457 16124
rect 4513 16078 4565 16124
rect 4621 16078 4673 16124
rect 4729 16078 4781 16124
rect 4837 16078 4889 16124
rect 4945 16078 4997 16124
rect 5053 16078 5105 16124
rect 5161 16078 5213 16124
rect 6566 16078 6618 16124
rect 6674 16078 6726 16124
rect 6782 16078 6834 16124
rect 6890 16078 6942 16124
rect 6998 16078 7050 16124
rect 7106 16078 7158 16124
rect 7214 16078 7266 16124
rect 7322 16078 7374 16124
rect 7430 16078 7482 16124
rect 7538 16078 7590 16124
rect 9677 16078 9729 16124
rect 9785 16078 9837 16124
rect 9893 16078 9945 16124
rect 10001 16078 10053 16124
rect 10109 16078 10161 16124
rect 10217 16078 10269 16124
rect 10325 16078 10377 16124
rect 10433 16078 10485 16124
rect 10541 16078 10593 16124
rect 10649 16078 10701 16124
rect 10757 16078 10809 16124
rect 10865 16078 10917 16124
rect 10973 16078 11025 16124
rect 11081 16078 11133 16124
rect 11189 16078 11241 16124
rect 11297 16078 11349 16124
rect 11405 16078 11457 16124
rect 3433 16075 3485 16078
rect 3541 16075 3593 16078
rect 3649 16075 3701 16078
rect 3757 16075 3809 16078
rect 3865 16075 3917 16078
rect 3973 16075 4025 16078
rect 4081 16075 4133 16078
rect 4189 16075 4241 16078
rect 4297 16075 4349 16078
rect 4405 16075 4457 16078
rect 4513 16075 4565 16078
rect 4621 16075 4673 16078
rect 4729 16075 4781 16078
rect 4837 16075 4889 16078
rect 4945 16075 4997 16078
rect 5053 16075 5105 16078
rect 5161 16075 5213 16078
rect 6566 16075 6618 16078
rect 6674 16075 6726 16078
rect 6782 16075 6834 16078
rect 6890 16075 6942 16078
rect 6998 16075 7050 16078
rect 7106 16075 7158 16078
rect 7214 16075 7266 16078
rect 7322 16075 7374 16078
rect 7430 16075 7482 16078
rect 7538 16075 7590 16078
rect 9677 16075 9729 16078
rect 9785 16075 9837 16078
rect 9893 16075 9945 16078
rect 10001 16075 10053 16078
rect 10109 16075 10161 16078
rect 10217 16075 10269 16078
rect 10325 16075 10377 16078
rect 10433 16075 10485 16078
rect 10541 16075 10593 16078
rect 10649 16075 10701 16078
rect 10757 16075 10809 16078
rect 10865 16075 10917 16078
rect 10973 16075 11025 16078
rect 11081 16075 11133 16078
rect 11189 16075 11241 16078
rect 11297 16075 11349 16078
rect 11405 16075 11457 16078
rect 1505 15880 1557 15883
rect 1613 15880 1665 15883
rect 1721 15880 1773 15883
rect 1829 15880 1881 15883
rect 1937 15880 1989 15883
rect 2045 15880 2097 15883
rect 2153 15880 2205 15883
rect 2261 15880 2313 15883
rect 2369 15880 2421 15883
rect 2477 15880 2529 15883
rect 2585 15880 2637 15883
rect 2693 15880 2745 15883
rect 2801 15880 2853 15883
rect 2909 15880 2961 15883
rect 3017 15880 3069 15883
rect 3125 15880 3177 15883
rect 3233 15880 3285 15883
rect 5372 15880 5424 15883
rect 5480 15880 5532 15883
rect 5588 15880 5640 15883
rect 5696 15880 5748 15883
rect 5804 15880 5856 15883
rect 5912 15880 5964 15883
rect 6020 15880 6072 15883
rect 6128 15880 6180 15883
rect 6236 15880 6288 15883
rect 6344 15880 6396 15883
rect 7749 15880 7801 15883
rect 7857 15880 7909 15883
rect 7965 15880 8017 15883
rect 8073 15880 8125 15883
rect 8181 15880 8233 15883
rect 8289 15880 8341 15883
rect 8397 15880 8449 15883
rect 8505 15880 8557 15883
rect 8613 15880 8665 15883
rect 8721 15880 8773 15883
rect 8829 15880 8881 15883
rect 8937 15880 8989 15883
rect 9045 15880 9097 15883
rect 9153 15880 9205 15883
rect 9261 15880 9313 15883
rect 9369 15880 9421 15883
rect 9477 15880 9529 15883
rect 1505 15834 1557 15880
rect 1613 15834 1665 15880
rect 1721 15834 1773 15880
rect 1829 15834 1881 15880
rect 1937 15834 1989 15880
rect 2045 15834 2097 15880
rect 2153 15834 2205 15880
rect 2261 15834 2313 15880
rect 2369 15834 2421 15880
rect 2477 15834 2529 15880
rect 2585 15834 2637 15880
rect 2693 15834 2745 15880
rect 2801 15834 2853 15880
rect 2909 15834 2961 15880
rect 3017 15834 3069 15880
rect 3125 15834 3177 15880
rect 3233 15834 3285 15880
rect 5372 15834 5424 15880
rect 5480 15834 5532 15880
rect 5588 15834 5640 15880
rect 5696 15834 5748 15880
rect 5804 15834 5856 15880
rect 5912 15834 5964 15880
rect 6020 15834 6072 15880
rect 6128 15834 6180 15880
rect 6236 15834 6288 15880
rect 6344 15834 6396 15880
rect 7749 15834 7801 15880
rect 7857 15834 7909 15880
rect 7965 15834 8017 15880
rect 8073 15834 8125 15880
rect 8181 15834 8233 15880
rect 8289 15834 8341 15880
rect 8397 15834 8449 15880
rect 8505 15834 8557 15880
rect 8613 15834 8665 15880
rect 8721 15834 8773 15880
rect 8829 15834 8881 15880
rect 8937 15834 8989 15880
rect 9045 15834 9097 15880
rect 9153 15834 9205 15880
rect 9261 15834 9313 15880
rect 9369 15834 9421 15880
rect 9477 15834 9529 15880
rect 1505 15831 1557 15834
rect 1613 15831 1665 15834
rect 1721 15831 1773 15834
rect 1829 15831 1881 15834
rect 1937 15831 1989 15834
rect 2045 15831 2097 15834
rect 2153 15831 2205 15834
rect 2261 15831 2313 15834
rect 2369 15831 2421 15834
rect 2477 15831 2529 15834
rect 2585 15831 2637 15834
rect 2693 15831 2745 15834
rect 2801 15831 2853 15834
rect 2909 15831 2961 15834
rect 3017 15831 3069 15834
rect 3125 15831 3177 15834
rect 3233 15831 3285 15834
rect 5372 15831 5424 15834
rect 5480 15831 5532 15834
rect 5588 15831 5640 15834
rect 5696 15831 5748 15834
rect 5804 15831 5856 15834
rect 5912 15831 5964 15834
rect 6020 15831 6072 15834
rect 6128 15831 6180 15834
rect 6236 15831 6288 15834
rect 6344 15831 6396 15834
rect 7749 15831 7801 15834
rect 7857 15831 7909 15834
rect 7965 15831 8017 15834
rect 8073 15831 8125 15834
rect 8181 15831 8233 15834
rect 8289 15831 8341 15834
rect 8397 15831 8449 15834
rect 8505 15831 8557 15834
rect 8613 15831 8665 15834
rect 8721 15831 8773 15834
rect 8829 15831 8881 15834
rect 8937 15831 8989 15834
rect 9045 15831 9097 15834
rect 9153 15831 9205 15834
rect 9261 15831 9313 15834
rect 9369 15831 9421 15834
rect 9477 15831 9529 15834
rect 3433 15636 3485 15639
rect 3541 15636 3593 15639
rect 3649 15636 3701 15639
rect 3757 15636 3809 15639
rect 3865 15636 3917 15639
rect 3973 15636 4025 15639
rect 4081 15636 4133 15639
rect 4189 15636 4241 15639
rect 4297 15636 4349 15639
rect 4405 15636 4457 15639
rect 4513 15636 4565 15639
rect 4621 15636 4673 15639
rect 4729 15636 4781 15639
rect 4837 15636 4889 15639
rect 4945 15636 4997 15639
rect 5053 15636 5105 15639
rect 5161 15636 5213 15639
rect 6566 15636 6618 15639
rect 6674 15636 6726 15639
rect 6782 15636 6834 15639
rect 6890 15636 6942 15639
rect 6998 15636 7050 15639
rect 7106 15636 7158 15639
rect 7214 15636 7266 15639
rect 7322 15636 7374 15639
rect 7430 15636 7482 15639
rect 7538 15636 7590 15639
rect 9677 15636 9729 15639
rect 9785 15636 9837 15639
rect 9893 15636 9945 15639
rect 10001 15636 10053 15639
rect 10109 15636 10161 15639
rect 10217 15636 10269 15639
rect 10325 15636 10377 15639
rect 10433 15636 10485 15639
rect 10541 15636 10593 15639
rect 10649 15636 10701 15639
rect 10757 15636 10809 15639
rect 10865 15636 10917 15639
rect 10973 15636 11025 15639
rect 11081 15636 11133 15639
rect 11189 15636 11241 15639
rect 11297 15636 11349 15639
rect 11405 15636 11457 15639
rect 3433 15590 3485 15636
rect 3541 15590 3593 15636
rect 3649 15590 3701 15636
rect 3757 15590 3809 15636
rect 3865 15590 3917 15636
rect 3973 15590 4025 15636
rect 4081 15590 4133 15636
rect 4189 15590 4241 15636
rect 4297 15590 4349 15636
rect 4405 15590 4457 15636
rect 4513 15590 4565 15636
rect 4621 15590 4673 15636
rect 4729 15590 4781 15636
rect 4837 15590 4889 15636
rect 4945 15590 4997 15636
rect 5053 15590 5105 15636
rect 5161 15590 5213 15636
rect 6566 15590 6618 15636
rect 6674 15590 6726 15636
rect 6782 15590 6834 15636
rect 6890 15590 6942 15636
rect 6998 15590 7050 15636
rect 7106 15590 7158 15636
rect 7214 15590 7266 15636
rect 7322 15590 7374 15636
rect 7430 15590 7482 15636
rect 7538 15590 7590 15636
rect 9677 15590 9729 15636
rect 9785 15590 9837 15636
rect 9893 15590 9945 15636
rect 10001 15590 10053 15636
rect 10109 15590 10161 15636
rect 10217 15590 10269 15636
rect 10325 15590 10377 15636
rect 10433 15590 10485 15636
rect 10541 15590 10593 15636
rect 10649 15590 10701 15636
rect 10757 15590 10809 15636
rect 10865 15590 10917 15636
rect 10973 15590 11025 15636
rect 11081 15590 11133 15636
rect 11189 15590 11241 15636
rect 11297 15590 11349 15636
rect 11405 15590 11457 15636
rect 3433 15587 3485 15590
rect 3541 15587 3593 15590
rect 3649 15587 3701 15590
rect 3757 15587 3809 15590
rect 3865 15587 3917 15590
rect 3973 15587 4025 15590
rect 4081 15587 4133 15590
rect 4189 15587 4241 15590
rect 4297 15587 4349 15590
rect 4405 15587 4457 15590
rect 4513 15587 4565 15590
rect 4621 15587 4673 15590
rect 4729 15587 4781 15590
rect 4837 15587 4889 15590
rect 4945 15587 4997 15590
rect 5053 15587 5105 15590
rect 5161 15587 5213 15590
rect 6566 15587 6618 15590
rect 6674 15587 6726 15590
rect 6782 15587 6834 15590
rect 6890 15587 6942 15590
rect 6998 15587 7050 15590
rect 7106 15587 7158 15590
rect 7214 15587 7266 15590
rect 7322 15587 7374 15590
rect 7430 15587 7482 15590
rect 7538 15587 7590 15590
rect 9677 15587 9729 15590
rect 9785 15587 9837 15590
rect 9893 15587 9945 15590
rect 10001 15587 10053 15590
rect 10109 15587 10161 15590
rect 10217 15587 10269 15590
rect 10325 15587 10377 15590
rect 10433 15587 10485 15590
rect 10541 15587 10593 15590
rect 10649 15587 10701 15590
rect 10757 15587 10809 15590
rect 10865 15587 10917 15590
rect 10973 15587 11025 15590
rect 11081 15587 11133 15590
rect 11189 15587 11241 15590
rect 11297 15587 11349 15590
rect 11405 15587 11457 15590
rect 1505 15392 1557 15395
rect 1613 15392 1665 15395
rect 1721 15392 1773 15395
rect 1829 15392 1881 15395
rect 1937 15392 1989 15395
rect 2045 15392 2097 15395
rect 2153 15392 2205 15395
rect 2261 15392 2313 15395
rect 2369 15392 2421 15395
rect 2477 15392 2529 15395
rect 2585 15392 2637 15395
rect 2693 15392 2745 15395
rect 2801 15392 2853 15395
rect 2909 15392 2961 15395
rect 3017 15392 3069 15395
rect 3125 15392 3177 15395
rect 3233 15392 3285 15395
rect 5372 15392 5424 15395
rect 5480 15392 5532 15395
rect 5588 15392 5640 15395
rect 5696 15392 5748 15395
rect 5804 15392 5856 15395
rect 5912 15392 5964 15395
rect 6020 15392 6072 15395
rect 6128 15392 6180 15395
rect 6236 15392 6288 15395
rect 6344 15392 6396 15395
rect 7749 15392 7801 15395
rect 7857 15392 7909 15395
rect 7965 15392 8017 15395
rect 8073 15392 8125 15395
rect 8181 15392 8233 15395
rect 8289 15392 8341 15395
rect 8397 15392 8449 15395
rect 8505 15392 8557 15395
rect 8613 15392 8665 15395
rect 8721 15392 8773 15395
rect 8829 15392 8881 15395
rect 8937 15392 8989 15395
rect 9045 15392 9097 15395
rect 9153 15392 9205 15395
rect 9261 15392 9313 15395
rect 9369 15392 9421 15395
rect 9477 15392 9529 15395
rect 1505 15346 1557 15392
rect 1613 15346 1665 15392
rect 1721 15346 1773 15392
rect 1829 15346 1881 15392
rect 1937 15346 1989 15392
rect 2045 15346 2097 15392
rect 2153 15346 2205 15392
rect 2261 15346 2313 15392
rect 2369 15346 2421 15392
rect 2477 15346 2529 15392
rect 2585 15346 2637 15392
rect 2693 15346 2745 15392
rect 2801 15346 2853 15392
rect 2909 15346 2961 15392
rect 3017 15346 3069 15392
rect 3125 15346 3177 15392
rect 3233 15346 3285 15392
rect 5372 15346 5424 15392
rect 5480 15346 5532 15392
rect 5588 15346 5640 15392
rect 5696 15346 5748 15392
rect 5804 15346 5856 15392
rect 5912 15346 5964 15392
rect 6020 15346 6072 15392
rect 6128 15346 6180 15392
rect 6236 15346 6288 15392
rect 6344 15346 6396 15392
rect 7749 15346 7801 15392
rect 7857 15346 7909 15392
rect 7965 15346 8017 15392
rect 8073 15346 8125 15392
rect 8181 15346 8233 15392
rect 8289 15346 8341 15392
rect 8397 15346 8449 15392
rect 8505 15346 8557 15392
rect 8613 15346 8665 15392
rect 8721 15346 8773 15392
rect 8829 15346 8881 15392
rect 8937 15346 8989 15392
rect 9045 15346 9097 15392
rect 9153 15346 9205 15392
rect 9261 15346 9313 15392
rect 9369 15346 9421 15392
rect 9477 15346 9529 15392
rect 1505 15343 1557 15346
rect 1613 15343 1665 15346
rect 1721 15343 1773 15346
rect 1829 15343 1881 15346
rect 1937 15343 1989 15346
rect 2045 15343 2097 15346
rect 2153 15343 2205 15346
rect 2261 15343 2313 15346
rect 2369 15343 2421 15346
rect 2477 15343 2529 15346
rect 2585 15343 2637 15346
rect 2693 15343 2745 15346
rect 2801 15343 2853 15346
rect 2909 15343 2961 15346
rect 3017 15343 3069 15346
rect 3125 15343 3177 15346
rect 3233 15343 3285 15346
rect 5372 15343 5424 15346
rect 5480 15343 5532 15346
rect 5588 15343 5640 15346
rect 5696 15343 5748 15346
rect 5804 15343 5856 15346
rect 5912 15343 5964 15346
rect 6020 15343 6072 15346
rect 6128 15343 6180 15346
rect 6236 15343 6288 15346
rect 6344 15343 6396 15346
rect 7749 15343 7801 15346
rect 7857 15343 7909 15346
rect 7965 15343 8017 15346
rect 8073 15343 8125 15346
rect 8181 15343 8233 15346
rect 8289 15343 8341 15346
rect 8397 15343 8449 15346
rect 8505 15343 8557 15346
rect 8613 15343 8665 15346
rect 8721 15343 8773 15346
rect 8829 15343 8881 15346
rect 8937 15343 8989 15346
rect 9045 15343 9097 15346
rect 9153 15343 9205 15346
rect 9261 15343 9313 15346
rect 9369 15343 9421 15346
rect 9477 15343 9529 15346
rect 3433 15148 3485 15151
rect 3541 15148 3593 15151
rect 3649 15148 3701 15151
rect 3757 15148 3809 15151
rect 3865 15148 3917 15151
rect 3973 15148 4025 15151
rect 4081 15148 4133 15151
rect 4189 15148 4241 15151
rect 4297 15148 4349 15151
rect 4405 15148 4457 15151
rect 4513 15148 4565 15151
rect 4621 15148 4673 15151
rect 4729 15148 4781 15151
rect 4837 15148 4889 15151
rect 4945 15148 4997 15151
rect 5053 15148 5105 15151
rect 5161 15148 5213 15151
rect 6566 15148 6618 15151
rect 6674 15148 6726 15151
rect 6782 15148 6834 15151
rect 6890 15148 6942 15151
rect 6998 15148 7050 15151
rect 7106 15148 7158 15151
rect 7214 15148 7266 15151
rect 7322 15148 7374 15151
rect 7430 15148 7482 15151
rect 7538 15148 7590 15151
rect 9677 15148 9729 15151
rect 9785 15148 9837 15151
rect 9893 15148 9945 15151
rect 10001 15148 10053 15151
rect 10109 15148 10161 15151
rect 10217 15148 10269 15151
rect 10325 15148 10377 15151
rect 10433 15148 10485 15151
rect 10541 15148 10593 15151
rect 10649 15148 10701 15151
rect 10757 15148 10809 15151
rect 10865 15148 10917 15151
rect 10973 15148 11025 15151
rect 11081 15148 11133 15151
rect 11189 15148 11241 15151
rect 11297 15148 11349 15151
rect 11405 15148 11457 15151
rect 3433 15102 3485 15148
rect 3541 15102 3593 15148
rect 3649 15102 3701 15148
rect 3757 15102 3809 15148
rect 3865 15102 3917 15148
rect 3973 15102 4025 15148
rect 4081 15102 4133 15148
rect 4189 15102 4241 15148
rect 4297 15102 4349 15148
rect 4405 15102 4457 15148
rect 4513 15102 4565 15148
rect 4621 15102 4673 15148
rect 4729 15102 4781 15148
rect 4837 15102 4889 15148
rect 4945 15102 4997 15148
rect 5053 15102 5105 15148
rect 5161 15102 5213 15148
rect 6566 15102 6618 15148
rect 6674 15102 6726 15148
rect 6782 15102 6834 15148
rect 6890 15102 6942 15148
rect 6998 15102 7050 15148
rect 7106 15102 7158 15148
rect 7214 15102 7266 15148
rect 7322 15102 7374 15148
rect 7430 15102 7482 15148
rect 7538 15102 7590 15148
rect 9677 15102 9729 15148
rect 9785 15102 9837 15148
rect 9893 15102 9945 15148
rect 10001 15102 10053 15148
rect 10109 15102 10161 15148
rect 10217 15102 10269 15148
rect 10325 15102 10377 15148
rect 10433 15102 10485 15148
rect 10541 15102 10593 15148
rect 10649 15102 10701 15148
rect 10757 15102 10809 15148
rect 10865 15102 10917 15148
rect 10973 15102 11025 15148
rect 11081 15102 11133 15148
rect 11189 15102 11241 15148
rect 11297 15102 11349 15148
rect 11405 15102 11457 15148
rect 3433 15099 3485 15102
rect 3541 15099 3593 15102
rect 3649 15099 3701 15102
rect 3757 15099 3809 15102
rect 3865 15099 3917 15102
rect 3973 15099 4025 15102
rect 4081 15099 4133 15102
rect 4189 15099 4241 15102
rect 4297 15099 4349 15102
rect 4405 15099 4457 15102
rect 4513 15099 4565 15102
rect 4621 15099 4673 15102
rect 4729 15099 4781 15102
rect 4837 15099 4889 15102
rect 4945 15099 4997 15102
rect 5053 15099 5105 15102
rect 5161 15099 5213 15102
rect 6566 15099 6618 15102
rect 6674 15099 6726 15102
rect 6782 15099 6834 15102
rect 6890 15099 6942 15102
rect 6998 15099 7050 15102
rect 7106 15099 7158 15102
rect 7214 15099 7266 15102
rect 7322 15099 7374 15102
rect 7430 15099 7482 15102
rect 7538 15099 7590 15102
rect 9677 15099 9729 15102
rect 9785 15099 9837 15102
rect 9893 15099 9945 15102
rect 10001 15099 10053 15102
rect 10109 15099 10161 15102
rect 10217 15099 10269 15102
rect 10325 15099 10377 15102
rect 10433 15099 10485 15102
rect 10541 15099 10593 15102
rect 10649 15099 10701 15102
rect 10757 15099 10809 15102
rect 10865 15099 10917 15102
rect 10973 15099 11025 15102
rect 11081 15099 11133 15102
rect 11189 15099 11241 15102
rect 11297 15099 11349 15102
rect 11405 15099 11457 15102
rect 1505 14904 1557 14907
rect 1613 14904 1665 14907
rect 1721 14904 1773 14907
rect 1829 14904 1881 14907
rect 1937 14904 1989 14907
rect 2045 14904 2097 14907
rect 2153 14904 2205 14907
rect 2261 14904 2313 14907
rect 2369 14904 2421 14907
rect 2477 14904 2529 14907
rect 2585 14904 2637 14907
rect 2693 14904 2745 14907
rect 2801 14904 2853 14907
rect 2909 14904 2961 14907
rect 3017 14904 3069 14907
rect 3125 14904 3177 14907
rect 3233 14904 3285 14907
rect 5372 14904 5424 14907
rect 5480 14904 5532 14907
rect 5588 14904 5640 14907
rect 5696 14904 5748 14907
rect 5804 14904 5856 14907
rect 5912 14904 5964 14907
rect 6020 14904 6072 14907
rect 6128 14904 6180 14907
rect 6236 14904 6288 14907
rect 6344 14904 6396 14907
rect 7749 14904 7801 14907
rect 7857 14904 7909 14907
rect 7965 14904 8017 14907
rect 8073 14904 8125 14907
rect 8181 14904 8233 14907
rect 8289 14904 8341 14907
rect 8397 14904 8449 14907
rect 8505 14904 8557 14907
rect 8613 14904 8665 14907
rect 8721 14904 8773 14907
rect 8829 14904 8881 14907
rect 8937 14904 8989 14907
rect 9045 14904 9097 14907
rect 9153 14904 9205 14907
rect 9261 14904 9313 14907
rect 9369 14904 9421 14907
rect 9477 14904 9529 14907
rect 1505 14858 1557 14904
rect 1613 14858 1665 14904
rect 1721 14858 1773 14904
rect 1829 14858 1881 14904
rect 1937 14858 1989 14904
rect 2045 14858 2097 14904
rect 2153 14858 2205 14904
rect 2261 14858 2313 14904
rect 2369 14858 2421 14904
rect 2477 14858 2529 14904
rect 2585 14858 2637 14904
rect 2693 14858 2745 14904
rect 2801 14858 2853 14904
rect 2909 14858 2961 14904
rect 3017 14858 3069 14904
rect 3125 14858 3177 14904
rect 3233 14858 3285 14904
rect 5372 14858 5424 14904
rect 5480 14858 5532 14904
rect 5588 14858 5640 14904
rect 5696 14858 5748 14904
rect 5804 14858 5856 14904
rect 5912 14858 5964 14904
rect 6020 14858 6072 14904
rect 6128 14858 6180 14904
rect 6236 14858 6288 14904
rect 6344 14858 6396 14904
rect 7749 14858 7801 14904
rect 7857 14858 7909 14904
rect 7965 14858 8017 14904
rect 8073 14858 8125 14904
rect 8181 14858 8233 14904
rect 8289 14858 8341 14904
rect 8397 14858 8449 14904
rect 8505 14858 8557 14904
rect 8613 14858 8665 14904
rect 8721 14858 8773 14904
rect 8829 14858 8881 14904
rect 8937 14858 8989 14904
rect 9045 14858 9097 14904
rect 9153 14858 9205 14904
rect 9261 14858 9313 14904
rect 9369 14858 9421 14904
rect 9477 14858 9529 14904
rect 1505 14855 1557 14858
rect 1613 14855 1665 14858
rect 1721 14855 1773 14858
rect 1829 14855 1881 14858
rect 1937 14855 1989 14858
rect 2045 14855 2097 14858
rect 2153 14855 2205 14858
rect 2261 14855 2313 14858
rect 2369 14855 2421 14858
rect 2477 14855 2529 14858
rect 2585 14855 2637 14858
rect 2693 14855 2745 14858
rect 2801 14855 2853 14858
rect 2909 14855 2961 14858
rect 3017 14855 3069 14858
rect 3125 14855 3177 14858
rect 3233 14855 3285 14858
rect 5372 14855 5424 14858
rect 5480 14855 5532 14858
rect 5588 14855 5640 14858
rect 5696 14855 5748 14858
rect 5804 14855 5856 14858
rect 5912 14855 5964 14858
rect 6020 14855 6072 14858
rect 6128 14855 6180 14858
rect 6236 14855 6288 14858
rect 6344 14855 6396 14858
rect 7749 14855 7801 14858
rect 7857 14855 7909 14858
rect 7965 14855 8017 14858
rect 8073 14855 8125 14858
rect 8181 14855 8233 14858
rect 8289 14855 8341 14858
rect 8397 14855 8449 14858
rect 8505 14855 8557 14858
rect 8613 14855 8665 14858
rect 8721 14855 8773 14858
rect 8829 14855 8881 14858
rect 8937 14855 8989 14858
rect 9045 14855 9097 14858
rect 9153 14855 9205 14858
rect 9261 14855 9313 14858
rect 9369 14855 9421 14858
rect 9477 14855 9529 14858
rect 3433 14660 3485 14663
rect 3541 14660 3593 14663
rect 3649 14660 3701 14663
rect 3757 14660 3809 14663
rect 3865 14660 3917 14663
rect 3973 14660 4025 14663
rect 4081 14660 4133 14663
rect 4189 14660 4241 14663
rect 4297 14660 4349 14663
rect 4405 14660 4457 14663
rect 4513 14660 4565 14663
rect 4621 14660 4673 14663
rect 4729 14660 4781 14663
rect 4837 14660 4889 14663
rect 4945 14660 4997 14663
rect 5053 14660 5105 14663
rect 5161 14660 5213 14663
rect 6566 14660 6618 14663
rect 6674 14660 6726 14663
rect 6782 14660 6834 14663
rect 6890 14660 6942 14663
rect 6998 14660 7050 14663
rect 7106 14660 7158 14663
rect 7214 14660 7266 14663
rect 7322 14660 7374 14663
rect 7430 14660 7482 14663
rect 7538 14660 7590 14663
rect 9677 14660 9729 14663
rect 9785 14660 9837 14663
rect 9893 14660 9945 14663
rect 10001 14660 10053 14663
rect 10109 14660 10161 14663
rect 10217 14660 10269 14663
rect 10325 14660 10377 14663
rect 10433 14660 10485 14663
rect 10541 14660 10593 14663
rect 10649 14660 10701 14663
rect 10757 14660 10809 14663
rect 10865 14660 10917 14663
rect 10973 14660 11025 14663
rect 11081 14660 11133 14663
rect 11189 14660 11241 14663
rect 11297 14660 11349 14663
rect 11405 14660 11457 14663
rect 3433 14614 3485 14660
rect 3541 14614 3593 14660
rect 3649 14614 3701 14660
rect 3757 14614 3809 14660
rect 3865 14614 3917 14660
rect 3973 14614 4025 14660
rect 4081 14614 4133 14660
rect 4189 14614 4241 14660
rect 4297 14614 4349 14660
rect 4405 14614 4457 14660
rect 4513 14614 4565 14660
rect 4621 14614 4673 14660
rect 4729 14614 4781 14660
rect 4837 14614 4889 14660
rect 4945 14614 4997 14660
rect 5053 14614 5105 14660
rect 5161 14614 5213 14660
rect 6566 14614 6618 14660
rect 6674 14614 6726 14660
rect 6782 14614 6834 14660
rect 6890 14614 6942 14660
rect 6998 14614 7050 14660
rect 7106 14614 7158 14660
rect 7214 14614 7266 14660
rect 7322 14614 7374 14660
rect 7430 14614 7482 14660
rect 7538 14614 7590 14660
rect 9677 14614 9729 14660
rect 9785 14614 9837 14660
rect 9893 14614 9945 14660
rect 10001 14614 10053 14660
rect 10109 14614 10161 14660
rect 10217 14614 10269 14660
rect 10325 14614 10377 14660
rect 10433 14614 10485 14660
rect 10541 14614 10593 14660
rect 10649 14614 10701 14660
rect 10757 14614 10809 14660
rect 10865 14614 10917 14660
rect 10973 14614 11025 14660
rect 11081 14614 11133 14660
rect 11189 14614 11241 14660
rect 11297 14614 11349 14660
rect 11405 14614 11457 14660
rect 3433 14611 3485 14614
rect 3541 14611 3593 14614
rect 3649 14611 3701 14614
rect 3757 14611 3809 14614
rect 3865 14611 3917 14614
rect 3973 14611 4025 14614
rect 4081 14611 4133 14614
rect 4189 14611 4241 14614
rect 4297 14611 4349 14614
rect 4405 14611 4457 14614
rect 4513 14611 4565 14614
rect 4621 14611 4673 14614
rect 4729 14611 4781 14614
rect 4837 14611 4889 14614
rect 4945 14611 4997 14614
rect 5053 14611 5105 14614
rect 5161 14611 5213 14614
rect 6566 14611 6618 14614
rect 6674 14611 6726 14614
rect 6782 14611 6834 14614
rect 6890 14611 6942 14614
rect 6998 14611 7050 14614
rect 7106 14611 7158 14614
rect 7214 14611 7266 14614
rect 7322 14611 7374 14614
rect 7430 14611 7482 14614
rect 7538 14611 7590 14614
rect 9677 14611 9729 14614
rect 9785 14611 9837 14614
rect 9893 14611 9945 14614
rect 10001 14611 10053 14614
rect 10109 14611 10161 14614
rect 10217 14611 10269 14614
rect 10325 14611 10377 14614
rect 10433 14611 10485 14614
rect 10541 14611 10593 14614
rect 10649 14611 10701 14614
rect 10757 14611 10809 14614
rect 10865 14611 10917 14614
rect 10973 14611 11025 14614
rect 11081 14611 11133 14614
rect 11189 14611 11241 14614
rect 11297 14611 11349 14614
rect 11405 14611 11457 14614
rect 1505 14416 1557 14419
rect 1613 14416 1665 14419
rect 1721 14416 1773 14419
rect 1829 14416 1881 14419
rect 1937 14416 1989 14419
rect 2045 14416 2097 14419
rect 2153 14416 2205 14419
rect 2261 14416 2313 14419
rect 2369 14416 2421 14419
rect 2477 14416 2529 14419
rect 2585 14416 2637 14419
rect 2693 14416 2745 14419
rect 2801 14416 2853 14419
rect 2909 14416 2961 14419
rect 3017 14416 3069 14419
rect 3125 14416 3177 14419
rect 3233 14416 3285 14419
rect 5372 14416 5424 14419
rect 5480 14416 5532 14419
rect 5588 14416 5640 14419
rect 5696 14416 5748 14419
rect 5804 14416 5856 14419
rect 5912 14416 5964 14419
rect 6020 14416 6072 14419
rect 6128 14416 6180 14419
rect 6236 14416 6288 14419
rect 6344 14416 6396 14419
rect 7749 14416 7801 14419
rect 7857 14416 7909 14419
rect 7965 14416 8017 14419
rect 8073 14416 8125 14419
rect 8181 14416 8233 14419
rect 8289 14416 8341 14419
rect 8397 14416 8449 14419
rect 8505 14416 8557 14419
rect 8613 14416 8665 14419
rect 8721 14416 8773 14419
rect 8829 14416 8881 14419
rect 8937 14416 8989 14419
rect 9045 14416 9097 14419
rect 9153 14416 9205 14419
rect 9261 14416 9313 14419
rect 9369 14416 9421 14419
rect 9477 14416 9529 14419
rect 1505 14370 1557 14416
rect 1613 14370 1665 14416
rect 1721 14370 1773 14416
rect 1829 14370 1881 14416
rect 1937 14370 1989 14416
rect 2045 14370 2097 14416
rect 2153 14370 2205 14416
rect 2261 14370 2313 14416
rect 2369 14370 2421 14416
rect 2477 14370 2529 14416
rect 2585 14370 2637 14416
rect 2693 14370 2745 14416
rect 2801 14370 2853 14416
rect 2909 14370 2961 14416
rect 3017 14370 3069 14416
rect 3125 14370 3177 14416
rect 3233 14370 3285 14416
rect 5372 14370 5424 14416
rect 5480 14370 5532 14416
rect 5588 14370 5640 14416
rect 5696 14370 5748 14416
rect 5804 14370 5856 14416
rect 5912 14370 5964 14416
rect 6020 14370 6072 14416
rect 6128 14370 6180 14416
rect 6236 14370 6288 14416
rect 6344 14370 6396 14416
rect 7749 14370 7801 14416
rect 7857 14370 7909 14416
rect 7965 14370 8017 14416
rect 8073 14370 8125 14416
rect 8181 14370 8233 14416
rect 8289 14370 8341 14416
rect 8397 14370 8449 14416
rect 8505 14370 8557 14416
rect 8613 14370 8665 14416
rect 8721 14370 8773 14416
rect 8829 14370 8881 14416
rect 8937 14370 8989 14416
rect 9045 14370 9097 14416
rect 9153 14370 9205 14416
rect 9261 14370 9313 14416
rect 9369 14370 9421 14416
rect 9477 14370 9529 14416
rect 1505 14367 1557 14370
rect 1613 14367 1665 14370
rect 1721 14367 1773 14370
rect 1829 14367 1881 14370
rect 1937 14367 1989 14370
rect 2045 14367 2097 14370
rect 2153 14367 2205 14370
rect 2261 14367 2313 14370
rect 2369 14367 2421 14370
rect 2477 14367 2529 14370
rect 2585 14367 2637 14370
rect 2693 14367 2745 14370
rect 2801 14367 2853 14370
rect 2909 14367 2961 14370
rect 3017 14367 3069 14370
rect 3125 14367 3177 14370
rect 3233 14367 3285 14370
rect 5372 14367 5424 14370
rect 5480 14367 5532 14370
rect 5588 14367 5640 14370
rect 5696 14367 5748 14370
rect 5804 14367 5856 14370
rect 5912 14367 5964 14370
rect 6020 14367 6072 14370
rect 6128 14367 6180 14370
rect 6236 14367 6288 14370
rect 6344 14367 6396 14370
rect 7749 14367 7801 14370
rect 7857 14367 7909 14370
rect 7965 14367 8017 14370
rect 8073 14367 8125 14370
rect 8181 14367 8233 14370
rect 8289 14367 8341 14370
rect 8397 14367 8449 14370
rect 8505 14367 8557 14370
rect 8613 14367 8665 14370
rect 8721 14367 8773 14370
rect 8829 14367 8881 14370
rect 8937 14367 8989 14370
rect 9045 14367 9097 14370
rect 9153 14367 9205 14370
rect 9261 14367 9313 14370
rect 9369 14367 9421 14370
rect 9477 14367 9529 14370
rect 3433 14172 3485 14175
rect 3541 14172 3593 14175
rect 3649 14172 3701 14175
rect 3757 14172 3809 14175
rect 3865 14172 3917 14175
rect 3973 14172 4025 14175
rect 4081 14172 4133 14175
rect 4189 14172 4241 14175
rect 4297 14172 4349 14175
rect 4405 14172 4457 14175
rect 4513 14172 4565 14175
rect 4621 14172 4673 14175
rect 4729 14172 4781 14175
rect 4837 14172 4889 14175
rect 4945 14172 4997 14175
rect 5053 14172 5105 14175
rect 5161 14172 5213 14175
rect 6566 14172 6618 14175
rect 6674 14172 6726 14175
rect 6782 14172 6834 14175
rect 6890 14172 6942 14175
rect 6998 14172 7050 14175
rect 7106 14172 7158 14175
rect 7214 14172 7266 14175
rect 7322 14172 7374 14175
rect 7430 14172 7482 14175
rect 7538 14172 7590 14175
rect 9677 14172 9729 14175
rect 9785 14172 9837 14175
rect 9893 14172 9945 14175
rect 10001 14172 10053 14175
rect 10109 14172 10161 14175
rect 10217 14172 10269 14175
rect 10325 14172 10377 14175
rect 10433 14172 10485 14175
rect 10541 14172 10593 14175
rect 10649 14172 10701 14175
rect 10757 14172 10809 14175
rect 10865 14172 10917 14175
rect 10973 14172 11025 14175
rect 11081 14172 11133 14175
rect 11189 14172 11241 14175
rect 11297 14172 11349 14175
rect 11405 14172 11457 14175
rect 3433 14126 3485 14172
rect 3541 14126 3593 14172
rect 3649 14126 3701 14172
rect 3757 14126 3809 14172
rect 3865 14126 3917 14172
rect 3973 14126 4025 14172
rect 4081 14126 4133 14172
rect 4189 14126 4241 14172
rect 4297 14126 4349 14172
rect 4405 14126 4457 14172
rect 4513 14126 4565 14172
rect 4621 14126 4673 14172
rect 4729 14126 4781 14172
rect 4837 14126 4889 14172
rect 4945 14126 4997 14172
rect 5053 14126 5105 14172
rect 5161 14126 5213 14172
rect 6566 14126 6618 14172
rect 6674 14126 6726 14172
rect 6782 14126 6834 14172
rect 6890 14126 6942 14172
rect 6998 14126 7050 14172
rect 7106 14126 7158 14172
rect 7214 14126 7266 14172
rect 7322 14126 7374 14172
rect 7430 14126 7482 14172
rect 7538 14126 7590 14172
rect 9677 14126 9729 14172
rect 9785 14126 9837 14172
rect 9893 14126 9945 14172
rect 10001 14126 10053 14172
rect 10109 14126 10161 14172
rect 10217 14126 10269 14172
rect 10325 14126 10377 14172
rect 10433 14126 10485 14172
rect 10541 14126 10593 14172
rect 10649 14126 10701 14172
rect 10757 14126 10809 14172
rect 10865 14126 10917 14172
rect 10973 14126 11025 14172
rect 11081 14126 11133 14172
rect 11189 14126 11241 14172
rect 11297 14126 11349 14172
rect 11405 14126 11457 14172
rect 3433 14123 3485 14126
rect 3541 14123 3593 14126
rect 3649 14123 3701 14126
rect 3757 14123 3809 14126
rect 3865 14123 3917 14126
rect 3973 14123 4025 14126
rect 4081 14123 4133 14126
rect 4189 14123 4241 14126
rect 4297 14123 4349 14126
rect 4405 14123 4457 14126
rect 4513 14123 4565 14126
rect 4621 14123 4673 14126
rect 4729 14123 4781 14126
rect 4837 14123 4889 14126
rect 4945 14123 4997 14126
rect 5053 14123 5105 14126
rect 5161 14123 5213 14126
rect 6566 14123 6618 14126
rect 6674 14123 6726 14126
rect 6782 14123 6834 14126
rect 6890 14123 6942 14126
rect 6998 14123 7050 14126
rect 7106 14123 7158 14126
rect 7214 14123 7266 14126
rect 7322 14123 7374 14126
rect 7430 14123 7482 14126
rect 7538 14123 7590 14126
rect 9677 14123 9729 14126
rect 9785 14123 9837 14126
rect 9893 14123 9945 14126
rect 10001 14123 10053 14126
rect 10109 14123 10161 14126
rect 10217 14123 10269 14126
rect 10325 14123 10377 14126
rect 10433 14123 10485 14126
rect 10541 14123 10593 14126
rect 10649 14123 10701 14126
rect 10757 14123 10809 14126
rect 10865 14123 10917 14126
rect 10973 14123 11025 14126
rect 11081 14123 11133 14126
rect 11189 14123 11241 14126
rect 11297 14123 11349 14126
rect 11405 14123 11457 14126
rect 1505 13928 1557 13931
rect 1613 13928 1665 13931
rect 1721 13928 1773 13931
rect 1829 13928 1881 13931
rect 1937 13928 1989 13931
rect 2045 13928 2097 13931
rect 2153 13928 2205 13931
rect 2261 13928 2313 13931
rect 2369 13928 2421 13931
rect 2477 13928 2529 13931
rect 2585 13928 2637 13931
rect 2693 13928 2745 13931
rect 2801 13928 2853 13931
rect 2909 13928 2961 13931
rect 3017 13928 3069 13931
rect 3125 13928 3177 13931
rect 3233 13928 3285 13931
rect 5372 13928 5424 13931
rect 5480 13928 5532 13931
rect 5588 13928 5640 13931
rect 5696 13928 5748 13931
rect 5804 13928 5856 13931
rect 5912 13928 5964 13931
rect 6020 13928 6072 13931
rect 6128 13928 6180 13931
rect 6236 13928 6288 13931
rect 6344 13928 6396 13931
rect 7749 13928 7801 13931
rect 7857 13928 7909 13931
rect 7965 13928 8017 13931
rect 8073 13928 8125 13931
rect 8181 13928 8233 13931
rect 8289 13928 8341 13931
rect 8397 13928 8449 13931
rect 8505 13928 8557 13931
rect 8613 13928 8665 13931
rect 8721 13928 8773 13931
rect 8829 13928 8881 13931
rect 8937 13928 8989 13931
rect 9045 13928 9097 13931
rect 9153 13928 9205 13931
rect 9261 13928 9313 13931
rect 9369 13928 9421 13931
rect 9477 13928 9529 13931
rect 1505 13882 1557 13928
rect 1613 13882 1665 13928
rect 1721 13882 1773 13928
rect 1829 13882 1881 13928
rect 1937 13882 1989 13928
rect 2045 13882 2097 13928
rect 2153 13882 2205 13928
rect 2261 13882 2313 13928
rect 2369 13882 2421 13928
rect 2477 13882 2529 13928
rect 2585 13882 2637 13928
rect 2693 13882 2745 13928
rect 2801 13882 2853 13928
rect 2909 13882 2961 13928
rect 3017 13882 3069 13928
rect 3125 13882 3177 13928
rect 3233 13882 3285 13928
rect 5372 13882 5424 13928
rect 5480 13882 5532 13928
rect 5588 13882 5640 13928
rect 5696 13882 5748 13928
rect 5804 13882 5856 13928
rect 5912 13882 5964 13928
rect 6020 13882 6072 13928
rect 6128 13882 6180 13928
rect 6236 13882 6288 13928
rect 6344 13882 6396 13928
rect 7749 13882 7801 13928
rect 7857 13882 7909 13928
rect 7965 13882 8017 13928
rect 8073 13882 8125 13928
rect 8181 13882 8233 13928
rect 8289 13882 8341 13928
rect 8397 13882 8449 13928
rect 8505 13882 8557 13928
rect 8613 13882 8665 13928
rect 8721 13882 8773 13928
rect 8829 13882 8881 13928
rect 8937 13882 8989 13928
rect 9045 13882 9097 13928
rect 9153 13882 9205 13928
rect 9261 13882 9313 13928
rect 9369 13882 9421 13928
rect 9477 13882 9529 13928
rect 1505 13879 1557 13882
rect 1613 13879 1665 13882
rect 1721 13879 1773 13882
rect 1829 13879 1881 13882
rect 1937 13879 1989 13882
rect 2045 13879 2097 13882
rect 2153 13879 2205 13882
rect 2261 13879 2313 13882
rect 2369 13879 2421 13882
rect 2477 13879 2529 13882
rect 2585 13879 2637 13882
rect 2693 13879 2745 13882
rect 2801 13879 2853 13882
rect 2909 13879 2961 13882
rect 3017 13879 3069 13882
rect 3125 13879 3177 13882
rect 3233 13879 3285 13882
rect 5372 13879 5424 13882
rect 5480 13879 5532 13882
rect 5588 13879 5640 13882
rect 5696 13879 5748 13882
rect 5804 13879 5856 13882
rect 5912 13879 5964 13882
rect 6020 13879 6072 13882
rect 6128 13879 6180 13882
rect 6236 13879 6288 13882
rect 6344 13879 6396 13882
rect 7749 13879 7801 13882
rect 7857 13879 7909 13882
rect 7965 13879 8017 13882
rect 8073 13879 8125 13882
rect 8181 13879 8233 13882
rect 8289 13879 8341 13882
rect 8397 13879 8449 13882
rect 8505 13879 8557 13882
rect 8613 13879 8665 13882
rect 8721 13879 8773 13882
rect 8829 13879 8881 13882
rect 8937 13879 8989 13882
rect 9045 13879 9097 13882
rect 9153 13879 9205 13882
rect 9261 13879 9313 13882
rect 9369 13879 9421 13882
rect 9477 13879 9529 13882
rect 3433 13684 3485 13687
rect 3541 13684 3593 13687
rect 3649 13684 3701 13687
rect 3757 13684 3809 13687
rect 3865 13684 3917 13687
rect 3973 13684 4025 13687
rect 4081 13684 4133 13687
rect 4189 13684 4241 13687
rect 4297 13684 4349 13687
rect 4405 13684 4457 13687
rect 4513 13684 4565 13687
rect 4621 13684 4673 13687
rect 4729 13684 4781 13687
rect 4837 13684 4889 13687
rect 4945 13684 4997 13687
rect 5053 13684 5105 13687
rect 5161 13684 5213 13687
rect 6566 13684 6618 13687
rect 6674 13684 6726 13687
rect 6782 13684 6834 13687
rect 6890 13684 6942 13687
rect 6998 13684 7050 13687
rect 7106 13684 7158 13687
rect 7214 13684 7266 13687
rect 7322 13684 7374 13687
rect 7430 13684 7482 13687
rect 7538 13684 7590 13687
rect 9677 13684 9729 13687
rect 9785 13684 9837 13687
rect 9893 13684 9945 13687
rect 10001 13684 10053 13687
rect 10109 13684 10161 13687
rect 10217 13684 10269 13687
rect 10325 13684 10377 13687
rect 10433 13684 10485 13687
rect 10541 13684 10593 13687
rect 10649 13684 10701 13687
rect 10757 13684 10809 13687
rect 10865 13684 10917 13687
rect 10973 13684 11025 13687
rect 11081 13684 11133 13687
rect 11189 13684 11241 13687
rect 11297 13684 11349 13687
rect 11405 13684 11457 13687
rect 3433 13638 3485 13684
rect 3541 13638 3593 13684
rect 3649 13638 3701 13684
rect 3757 13638 3809 13684
rect 3865 13638 3917 13684
rect 3973 13638 4025 13684
rect 4081 13638 4133 13684
rect 4189 13638 4241 13684
rect 4297 13638 4349 13684
rect 4405 13638 4457 13684
rect 4513 13638 4565 13684
rect 4621 13638 4673 13684
rect 4729 13638 4781 13684
rect 4837 13638 4889 13684
rect 4945 13638 4997 13684
rect 5053 13638 5105 13684
rect 5161 13638 5213 13684
rect 6566 13638 6618 13684
rect 6674 13638 6726 13684
rect 6782 13638 6834 13684
rect 6890 13638 6942 13684
rect 6998 13638 7050 13684
rect 7106 13638 7158 13684
rect 7214 13638 7266 13684
rect 7322 13638 7374 13684
rect 7430 13638 7482 13684
rect 7538 13638 7590 13684
rect 9677 13638 9729 13684
rect 9785 13638 9837 13684
rect 9893 13638 9945 13684
rect 10001 13638 10053 13684
rect 10109 13638 10161 13684
rect 10217 13638 10269 13684
rect 10325 13638 10377 13684
rect 10433 13638 10485 13684
rect 10541 13638 10593 13684
rect 10649 13638 10701 13684
rect 10757 13638 10809 13684
rect 10865 13638 10917 13684
rect 10973 13638 11025 13684
rect 11081 13638 11133 13684
rect 11189 13638 11241 13684
rect 11297 13638 11349 13684
rect 11405 13638 11457 13684
rect 3433 13635 3485 13638
rect 3541 13635 3593 13638
rect 3649 13635 3701 13638
rect 3757 13635 3809 13638
rect 3865 13635 3917 13638
rect 3973 13635 4025 13638
rect 4081 13635 4133 13638
rect 4189 13635 4241 13638
rect 4297 13635 4349 13638
rect 4405 13635 4457 13638
rect 4513 13635 4565 13638
rect 4621 13635 4673 13638
rect 4729 13635 4781 13638
rect 4837 13635 4889 13638
rect 4945 13635 4997 13638
rect 5053 13635 5105 13638
rect 5161 13635 5213 13638
rect 6566 13635 6618 13638
rect 6674 13635 6726 13638
rect 6782 13635 6834 13638
rect 6890 13635 6942 13638
rect 6998 13635 7050 13638
rect 7106 13635 7158 13638
rect 7214 13635 7266 13638
rect 7322 13635 7374 13638
rect 7430 13635 7482 13638
rect 7538 13635 7590 13638
rect 9677 13635 9729 13638
rect 9785 13635 9837 13638
rect 9893 13635 9945 13638
rect 10001 13635 10053 13638
rect 10109 13635 10161 13638
rect 10217 13635 10269 13638
rect 10325 13635 10377 13638
rect 10433 13635 10485 13638
rect 10541 13635 10593 13638
rect 10649 13635 10701 13638
rect 10757 13635 10809 13638
rect 10865 13635 10917 13638
rect 10973 13635 11025 13638
rect 11081 13635 11133 13638
rect 11189 13635 11241 13638
rect 11297 13635 11349 13638
rect 11405 13635 11457 13638
rect 1505 13440 1557 13443
rect 1613 13440 1665 13443
rect 1721 13440 1773 13443
rect 1829 13440 1881 13443
rect 1937 13440 1989 13443
rect 2045 13440 2097 13443
rect 2153 13440 2205 13443
rect 2261 13440 2313 13443
rect 2369 13440 2421 13443
rect 2477 13440 2529 13443
rect 2585 13440 2637 13443
rect 2693 13440 2745 13443
rect 2801 13440 2853 13443
rect 2909 13440 2961 13443
rect 3017 13440 3069 13443
rect 3125 13440 3177 13443
rect 3233 13440 3285 13443
rect 5372 13440 5424 13443
rect 5480 13440 5532 13443
rect 5588 13440 5640 13443
rect 5696 13440 5748 13443
rect 5804 13440 5856 13443
rect 5912 13440 5964 13443
rect 6020 13440 6072 13443
rect 6128 13440 6180 13443
rect 6236 13440 6288 13443
rect 6344 13440 6396 13443
rect 7749 13440 7801 13443
rect 7857 13440 7909 13443
rect 7965 13440 8017 13443
rect 8073 13440 8125 13443
rect 8181 13440 8233 13443
rect 8289 13440 8341 13443
rect 8397 13440 8449 13443
rect 8505 13440 8557 13443
rect 8613 13440 8665 13443
rect 8721 13440 8773 13443
rect 8829 13440 8881 13443
rect 8937 13440 8989 13443
rect 9045 13440 9097 13443
rect 9153 13440 9205 13443
rect 9261 13440 9313 13443
rect 9369 13440 9421 13443
rect 9477 13440 9529 13443
rect 1505 13394 1557 13440
rect 1613 13394 1665 13440
rect 1721 13394 1773 13440
rect 1829 13394 1881 13440
rect 1937 13394 1989 13440
rect 2045 13394 2097 13440
rect 2153 13394 2205 13440
rect 2261 13394 2313 13440
rect 2369 13394 2421 13440
rect 2477 13394 2529 13440
rect 2585 13394 2637 13440
rect 2693 13394 2745 13440
rect 2801 13394 2853 13440
rect 2909 13394 2961 13440
rect 3017 13394 3069 13440
rect 3125 13394 3177 13440
rect 3233 13394 3285 13440
rect 5372 13394 5424 13440
rect 5480 13394 5532 13440
rect 5588 13394 5640 13440
rect 5696 13394 5748 13440
rect 5804 13394 5856 13440
rect 5912 13394 5964 13440
rect 6020 13394 6072 13440
rect 6128 13394 6180 13440
rect 6236 13394 6288 13440
rect 6344 13394 6396 13440
rect 7749 13394 7801 13440
rect 7857 13394 7909 13440
rect 7965 13394 8017 13440
rect 8073 13394 8125 13440
rect 8181 13394 8233 13440
rect 8289 13394 8341 13440
rect 8397 13394 8449 13440
rect 8505 13394 8557 13440
rect 8613 13394 8665 13440
rect 8721 13394 8773 13440
rect 8829 13394 8881 13440
rect 8937 13394 8989 13440
rect 9045 13394 9097 13440
rect 9153 13394 9205 13440
rect 9261 13394 9313 13440
rect 9369 13394 9421 13440
rect 9477 13394 9529 13440
rect 1505 13391 1557 13394
rect 1613 13391 1665 13394
rect 1721 13391 1773 13394
rect 1829 13391 1881 13394
rect 1937 13391 1989 13394
rect 2045 13391 2097 13394
rect 2153 13391 2205 13394
rect 2261 13391 2313 13394
rect 2369 13391 2421 13394
rect 2477 13391 2529 13394
rect 2585 13391 2637 13394
rect 2693 13391 2745 13394
rect 2801 13391 2853 13394
rect 2909 13391 2961 13394
rect 3017 13391 3069 13394
rect 3125 13391 3177 13394
rect 3233 13391 3285 13394
rect 5372 13391 5424 13394
rect 5480 13391 5532 13394
rect 5588 13391 5640 13394
rect 5696 13391 5748 13394
rect 5804 13391 5856 13394
rect 5912 13391 5964 13394
rect 6020 13391 6072 13394
rect 6128 13391 6180 13394
rect 6236 13391 6288 13394
rect 6344 13391 6396 13394
rect 7749 13391 7801 13394
rect 7857 13391 7909 13394
rect 7965 13391 8017 13394
rect 8073 13391 8125 13394
rect 8181 13391 8233 13394
rect 8289 13391 8341 13394
rect 8397 13391 8449 13394
rect 8505 13391 8557 13394
rect 8613 13391 8665 13394
rect 8721 13391 8773 13394
rect 8829 13391 8881 13394
rect 8937 13391 8989 13394
rect 9045 13391 9097 13394
rect 9153 13391 9205 13394
rect 9261 13391 9313 13394
rect 9369 13391 9421 13394
rect 9477 13391 9529 13394
rect 1233 13211 1285 13263
rect 1341 13211 1393 13263
rect 11569 17855 11621 17907
rect 11677 17855 11706 17907
rect 11706 17855 11729 17907
rect 11569 17747 11621 17799
rect 11677 17747 11706 17799
rect 11706 17747 11729 17799
rect 11569 17639 11621 17691
rect 11677 17639 11706 17691
rect 11706 17639 11729 17691
rect 11569 17531 11621 17583
rect 11677 17531 11706 17583
rect 11706 17531 11729 17583
rect 11569 17423 11621 17475
rect 11677 17423 11706 17475
rect 11706 17423 11729 17475
rect 11569 17315 11621 17367
rect 11677 17315 11706 17367
rect 11706 17315 11729 17367
rect 11569 17207 11621 17259
rect 11677 17207 11706 17259
rect 11706 17207 11729 17259
rect 11569 17099 11621 17151
rect 11677 17099 11706 17151
rect 11706 17099 11729 17151
rect 11569 16991 11621 17043
rect 11677 16991 11706 17043
rect 11706 16991 11729 17043
rect 11569 16883 11621 16935
rect 11677 16883 11706 16935
rect 11706 16883 11729 16935
rect 11569 16775 11621 16827
rect 11677 16775 11706 16827
rect 11706 16775 11729 16827
rect 11569 16667 11621 16719
rect 11677 16667 11706 16719
rect 11706 16667 11729 16719
rect 11569 16559 11621 16611
rect 11677 16559 11706 16611
rect 11706 16559 11729 16611
rect 11569 16451 11621 16503
rect 11677 16451 11706 16503
rect 11706 16451 11729 16503
rect 11569 16343 11621 16395
rect 11677 16343 11706 16395
rect 11706 16343 11729 16395
rect 11569 16235 11621 16287
rect 11677 16235 11706 16287
rect 11706 16235 11729 16287
rect 11569 16127 11621 16179
rect 11677 16127 11706 16179
rect 11706 16127 11729 16179
rect 11569 16019 11621 16071
rect 11677 16019 11706 16071
rect 11706 16019 11729 16071
rect 11569 15911 11621 15963
rect 11677 15911 11706 15963
rect 11706 15911 11729 15963
rect 11569 15803 11621 15855
rect 11677 15803 11706 15855
rect 11706 15803 11729 15855
rect 11569 15695 11621 15747
rect 11677 15695 11706 15747
rect 11706 15695 11729 15747
rect 11569 15587 11621 15639
rect 11677 15587 11706 15639
rect 11706 15587 11729 15639
rect 11569 15479 11621 15531
rect 11677 15479 11706 15531
rect 11706 15479 11729 15531
rect 11569 15371 11621 15423
rect 11677 15371 11706 15423
rect 11706 15371 11729 15423
rect 11569 15263 11621 15315
rect 11677 15263 11706 15315
rect 11706 15263 11729 15315
rect 11569 15155 11621 15207
rect 11677 15155 11706 15207
rect 11706 15155 11729 15207
rect 11569 15047 11621 15099
rect 11677 15047 11706 15099
rect 11706 15047 11729 15099
rect 11569 14939 11621 14991
rect 11677 14939 11706 14991
rect 11706 14939 11729 14991
rect 11569 14831 11621 14883
rect 11677 14831 11706 14883
rect 11706 14831 11729 14883
rect 11569 14723 11621 14775
rect 11677 14723 11706 14775
rect 11706 14723 11729 14775
rect 11569 14615 11621 14667
rect 11677 14615 11706 14667
rect 11706 14615 11729 14667
rect 11569 14507 11621 14559
rect 11677 14507 11706 14559
rect 11706 14507 11729 14559
rect 11569 14399 11621 14451
rect 11677 14399 11706 14451
rect 11706 14399 11729 14451
rect 11569 14291 11621 14343
rect 11677 14291 11706 14343
rect 11706 14291 11729 14343
rect 11569 14183 11621 14235
rect 11677 14183 11706 14235
rect 11706 14183 11729 14235
rect 11569 14075 11621 14127
rect 11677 14075 11706 14127
rect 11706 14075 11729 14127
rect 11569 13967 11621 14019
rect 11677 13967 11706 14019
rect 11706 13967 11729 14019
rect 11569 13859 11621 13911
rect 11677 13859 11706 13911
rect 11706 13859 11729 13911
rect 11569 13751 11621 13803
rect 11677 13751 11706 13803
rect 11706 13751 11729 13803
rect 11569 13643 11621 13695
rect 11677 13643 11706 13695
rect 11706 13643 11729 13695
rect 11569 13535 11621 13587
rect 11677 13535 11706 13587
rect 11706 13535 11729 13587
rect 11569 13427 11621 13479
rect 11677 13427 11706 13479
rect 11706 13427 11729 13479
rect 11569 13319 11621 13371
rect 11677 13319 11706 13371
rect 11706 13319 11729 13371
rect 11569 13211 11621 13263
rect 11677 13211 11729 13263
rect 3433 13196 3485 13199
rect 3541 13196 3593 13199
rect 3649 13196 3701 13199
rect 3757 13196 3809 13199
rect 3865 13196 3917 13199
rect 3973 13196 4025 13199
rect 4081 13196 4133 13199
rect 4189 13196 4241 13199
rect 4297 13196 4349 13199
rect 4405 13196 4457 13199
rect 4513 13196 4565 13199
rect 4621 13196 4673 13199
rect 4729 13196 4781 13199
rect 4837 13196 4889 13199
rect 4945 13196 4997 13199
rect 5053 13196 5105 13199
rect 5161 13196 5213 13199
rect 6566 13196 6618 13199
rect 6674 13196 6726 13199
rect 6782 13196 6834 13199
rect 6890 13196 6942 13199
rect 6998 13196 7050 13199
rect 7106 13196 7158 13199
rect 7214 13196 7266 13199
rect 7322 13196 7374 13199
rect 7430 13196 7482 13199
rect 7538 13196 7590 13199
rect 9677 13196 9729 13199
rect 9785 13196 9837 13199
rect 9893 13196 9945 13199
rect 10001 13196 10053 13199
rect 10109 13196 10161 13199
rect 10217 13196 10269 13199
rect 10325 13196 10377 13199
rect 10433 13196 10485 13199
rect 10541 13196 10593 13199
rect 10649 13196 10701 13199
rect 10757 13196 10809 13199
rect 10865 13196 10917 13199
rect 10973 13196 11025 13199
rect 11081 13196 11133 13199
rect 11189 13196 11241 13199
rect 11297 13196 11349 13199
rect 11405 13196 11457 13199
rect 3433 13150 3485 13196
rect 3541 13150 3593 13196
rect 3649 13150 3701 13196
rect 3757 13150 3809 13196
rect 3865 13150 3917 13196
rect 3973 13150 4025 13196
rect 4081 13150 4133 13196
rect 4189 13150 4241 13196
rect 4297 13150 4349 13196
rect 4405 13150 4457 13196
rect 4513 13150 4565 13196
rect 4621 13150 4673 13196
rect 4729 13150 4781 13196
rect 4837 13150 4889 13196
rect 4945 13150 4997 13196
rect 5053 13150 5105 13196
rect 5161 13150 5213 13196
rect 6566 13150 6618 13196
rect 6674 13150 6726 13196
rect 6782 13150 6834 13196
rect 6890 13150 6942 13196
rect 6998 13150 7050 13196
rect 7106 13150 7158 13196
rect 7214 13150 7266 13196
rect 7322 13150 7374 13196
rect 7430 13150 7482 13196
rect 7538 13150 7590 13196
rect 9677 13150 9729 13196
rect 9785 13150 9837 13196
rect 9893 13150 9945 13196
rect 10001 13150 10053 13196
rect 10109 13150 10161 13196
rect 10217 13150 10269 13196
rect 10325 13150 10377 13196
rect 10433 13150 10485 13196
rect 10541 13150 10593 13196
rect 10649 13150 10701 13196
rect 10757 13150 10809 13196
rect 10865 13150 10917 13196
rect 10973 13150 11025 13196
rect 11081 13150 11133 13196
rect 11189 13150 11241 13196
rect 11297 13150 11349 13196
rect 11405 13150 11457 13196
rect 3433 13147 3485 13150
rect 3541 13147 3593 13150
rect 3649 13147 3701 13150
rect 3757 13147 3809 13150
rect 3865 13147 3917 13150
rect 3973 13147 4025 13150
rect 4081 13147 4133 13150
rect 4189 13147 4241 13150
rect 4297 13147 4349 13150
rect 4405 13147 4457 13150
rect 4513 13147 4565 13150
rect 4621 13147 4673 13150
rect 4729 13147 4781 13150
rect 4837 13147 4889 13150
rect 4945 13147 4997 13150
rect 5053 13147 5105 13150
rect 5161 13147 5213 13150
rect 6566 13147 6618 13150
rect 6674 13147 6726 13150
rect 6782 13147 6834 13150
rect 6890 13147 6942 13150
rect 6998 13147 7050 13150
rect 7106 13147 7158 13150
rect 7214 13147 7266 13150
rect 7322 13147 7374 13150
rect 7430 13147 7482 13150
rect 7538 13147 7590 13150
rect 9677 13147 9729 13150
rect 9785 13147 9837 13150
rect 9893 13147 9945 13150
rect 10001 13147 10053 13150
rect 10109 13147 10161 13150
rect 10217 13147 10269 13150
rect 10325 13147 10377 13150
rect 10433 13147 10485 13150
rect 10541 13147 10593 13150
rect 10649 13147 10701 13150
rect 10757 13147 10809 13150
rect 10865 13147 10917 13150
rect 10973 13147 11025 13150
rect 11081 13147 11133 13150
rect 11189 13147 11241 13150
rect 11297 13147 11349 13150
rect 11405 13147 11457 13150
rect 12051 18429 12103 18481
rect 12159 18429 12211 18481
rect 12267 18429 12319 18481
rect 12051 18321 12103 18373
rect 12159 18321 12211 18373
rect 12267 18321 12319 18373
rect 12051 18213 12103 18265
rect 12159 18213 12211 18265
rect 12267 18213 12319 18265
rect 12051 18105 12103 18157
rect 12159 18105 12211 18157
rect 12267 18105 12319 18157
rect 12051 17997 12103 18049
rect 12159 17997 12211 18049
rect 12267 17997 12319 18049
rect 12051 17889 12103 17941
rect 12159 17889 12211 17941
rect 12267 17889 12319 17941
rect 12051 17781 12103 17833
rect 12159 17781 12211 17833
rect 12267 17781 12319 17833
rect 12051 17673 12103 17725
rect 12159 17673 12211 17725
rect 12267 17673 12319 17725
rect 12051 17565 12103 17617
rect 12159 17565 12211 17617
rect 12267 17565 12319 17617
rect 12051 17457 12103 17509
rect 12159 17457 12211 17509
rect 12267 17457 12319 17509
rect 12051 17349 12103 17401
rect 12159 17349 12211 17401
rect 12267 17349 12319 17401
rect 12051 17241 12103 17293
rect 12159 17241 12211 17293
rect 12267 17241 12319 17293
rect 12051 17133 12103 17185
rect 12159 17133 12211 17185
rect 12267 17133 12319 17185
rect 12051 17025 12103 17077
rect 12159 17025 12211 17077
rect 12267 17025 12319 17077
rect 12051 16917 12103 16969
rect 12159 16917 12211 16969
rect 12267 16917 12319 16969
rect 12051 16809 12103 16861
rect 12159 16809 12211 16861
rect 12267 16809 12319 16861
rect 12051 16701 12103 16753
rect 12159 16701 12211 16753
rect 12267 16701 12319 16753
rect 12051 16593 12103 16645
rect 12159 16593 12211 16645
rect 12267 16593 12319 16645
rect 12051 16485 12103 16537
rect 12159 16485 12211 16537
rect 12267 16485 12319 16537
rect 12051 16377 12103 16429
rect 12159 16377 12211 16429
rect 12267 16377 12319 16429
rect 12051 16269 12103 16321
rect 12159 16269 12211 16321
rect 12267 16269 12319 16321
rect 12051 16161 12103 16213
rect 12159 16161 12211 16213
rect 12267 16161 12319 16213
rect 12051 16053 12103 16105
rect 12159 16053 12211 16105
rect 12267 16053 12319 16105
rect 12051 15945 12103 15997
rect 12159 15945 12211 15997
rect 12267 15945 12319 15997
rect 12051 15837 12103 15889
rect 12159 15837 12211 15889
rect 12267 15837 12319 15889
rect 12051 15729 12103 15781
rect 12159 15729 12211 15781
rect 12267 15729 12319 15781
rect 12051 15621 12103 15673
rect 12159 15621 12211 15673
rect 12267 15621 12319 15673
rect 12051 15513 12103 15565
rect 12159 15513 12211 15565
rect 12267 15513 12319 15565
rect 12051 15405 12103 15457
rect 12159 15405 12211 15457
rect 12267 15405 12319 15457
rect 12051 15297 12103 15349
rect 12159 15297 12211 15349
rect 12267 15297 12319 15349
rect 12051 15189 12103 15241
rect 12159 15189 12211 15241
rect 12267 15189 12319 15241
rect 12051 15081 12103 15133
rect 12159 15081 12211 15133
rect 12267 15081 12319 15133
rect 12051 14973 12103 15025
rect 12159 14973 12211 15025
rect 12267 14973 12319 15025
rect 12051 14865 12103 14917
rect 12159 14865 12211 14917
rect 12267 14865 12319 14917
rect 12051 14757 12103 14809
rect 12159 14757 12211 14809
rect 12267 14757 12319 14809
rect 12051 14649 12103 14701
rect 12159 14649 12211 14701
rect 12267 14649 12319 14701
rect 12051 14541 12103 14593
rect 12159 14541 12211 14593
rect 12267 14541 12319 14593
rect 12051 14433 12103 14485
rect 12159 14433 12211 14485
rect 12267 14433 12319 14485
rect 12051 14325 12103 14377
rect 12159 14325 12211 14377
rect 12267 14325 12319 14377
rect 12051 14217 12103 14269
rect 12159 14217 12211 14269
rect 12267 14217 12319 14269
rect 12051 14109 12103 14161
rect 12159 14109 12211 14161
rect 12267 14109 12319 14161
rect 12051 14001 12103 14053
rect 12159 14001 12211 14053
rect 12267 14001 12319 14053
rect 12051 13893 12103 13945
rect 12159 13893 12211 13945
rect 12267 13893 12319 13945
rect 12051 13785 12103 13837
rect 12159 13785 12211 13837
rect 12267 13785 12319 13837
rect 12051 13677 12103 13729
rect 12159 13677 12211 13729
rect 12267 13677 12319 13729
rect 12051 13569 12103 13621
rect 12159 13569 12211 13621
rect 12267 13569 12319 13621
rect 12051 13461 12103 13513
rect 12159 13461 12211 13513
rect 12267 13461 12319 13513
rect 12051 13353 12103 13405
rect 12159 13353 12211 13405
rect 12267 13353 12319 13405
rect 12051 13245 12103 13297
rect 12159 13245 12211 13297
rect 12267 13245 12319 13297
rect 12051 13137 12103 13189
rect 12159 13137 12211 13189
rect 12267 13137 12319 13189
rect 12051 13029 12103 13081
rect 12159 13029 12211 13081
rect 12267 13029 12319 13081
rect 12051 12921 12103 12973
rect 12159 12921 12211 12973
rect 12267 12921 12319 12973
rect 12051 12813 12103 12865
rect 12159 12813 12211 12865
rect 12267 12813 12319 12865
rect 1505 12750 1557 12757
rect 1613 12750 1665 12757
rect 1721 12750 1773 12757
rect 1829 12750 1881 12757
rect 1937 12750 1989 12757
rect 2045 12750 2097 12757
rect 2153 12750 2205 12757
rect 2261 12750 2313 12757
rect 2369 12750 2421 12757
rect 2477 12750 2529 12757
rect 2585 12750 2637 12757
rect 2693 12750 2745 12757
rect 2801 12750 2853 12757
rect 2909 12750 2961 12757
rect 3017 12750 3069 12757
rect 3125 12750 3177 12757
rect 3233 12750 3285 12757
rect 5372 12750 5424 12757
rect 5480 12750 5532 12757
rect 5588 12750 5640 12757
rect 5696 12750 5748 12757
rect 5804 12750 5856 12757
rect 5912 12750 5964 12757
rect 6020 12750 6072 12757
rect 6128 12750 6180 12757
rect 6236 12750 6288 12757
rect 6344 12750 6396 12757
rect 7749 12750 7801 12757
rect 7857 12750 7909 12757
rect 7965 12750 8017 12757
rect 8073 12750 8125 12757
rect 8181 12750 8233 12757
rect 8289 12750 8341 12757
rect 8397 12750 8449 12757
rect 8505 12750 8557 12757
rect 8613 12750 8665 12757
rect 8721 12750 8773 12757
rect 8829 12750 8881 12757
rect 8937 12750 8989 12757
rect 9045 12750 9097 12757
rect 9153 12750 9205 12757
rect 9261 12750 9313 12757
rect 9369 12750 9421 12757
rect 9477 12750 9529 12757
rect 1505 12705 1557 12750
rect 1613 12705 1665 12750
rect 1721 12705 1773 12750
rect 1829 12705 1881 12750
rect 1937 12705 1989 12750
rect 2045 12705 2097 12750
rect 2153 12705 2205 12750
rect 2261 12705 2313 12750
rect 2369 12705 2421 12750
rect 2477 12705 2529 12750
rect 2585 12705 2637 12750
rect 2693 12705 2745 12750
rect 2801 12705 2853 12750
rect 2909 12705 2961 12750
rect 3017 12705 3069 12750
rect 3125 12705 3177 12750
rect 3233 12705 3285 12750
rect 5372 12705 5424 12750
rect 5480 12705 5532 12750
rect 5588 12705 5640 12750
rect 5696 12705 5748 12750
rect 5804 12705 5856 12750
rect 5912 12705 5964 12750
rect 6020 12705 6072 12750
rect 6128 12705 6180 12750
rect 6236 12705 6288 12750
rect 6344 12705 6396 12750
rect 7749 12705 7801 12750
rect 7857 12705 7909 12750
rect 7965 12705 8017 12750
rect 8073 12705 8125 12750
rect 8181 12705 8233 12750
rect 8289 12705 8341 12750
rect 8397 12705 8449 12750
rect 8505 12705 8557 12750
rect 8613 12705 8665 12750
rect 8721 12705 8773 12750
rect 8829 12705 8881 12750
rect 8937 12705 8989 12750
rect 9045 12705 9097 12750
rect 9153 12705 9205 12750
rect 9261 12705 9313 12750
rect 9369 12705 9421 12750
rect 9477 12705 9529 12750
rect 1505 12604 1557 12649
rect 1613 12604 1665 12649
rect 1721 12604 1773 12649
rect 1829 12604 1881 12649
rect 1937 12604 1989 12649
rect 2045 12604 2097 12649
rect 2153 12604 2205 12649
rect 2261 12604 2313 12649
rect 2369 12604 2421 12649
rect 2477 12604 2529 12649
rect 2585 12604 2637 12649
rect 2693 12604 2745 12649
rect 2801 12604 2853 12649
rect 2909 12604 2961 12649
rect 3017 12604 3069 12649
rect 3125 12604 3177 12649
rect 3233 12604 3285 12649
rect 5372 12604 5424 12649
rect 5480 12604 5532 12649
rect 5588 12604 5640 12649
rect 5696 12604 5748 12649
rect 5804 12604 5856 12649
rect 5912 12604 5964 12649
rect 6020 12604 6072 12649
rect 6128 12604 6180 12649
rect 6236 12604 6288 12649
rect 6344 12604 6396 12649
rect 7749 12604 7801 12649
rect 7857 12604 7909 12649
rect 7965 12604 8017 12649
rect 8073 12604 8125 12649
rect 8181 12604 8233 12649
rect 8289 12604 8341 12649
rect 8397 12604 8449 12649
rect 8505 12604 8557 12649
rect 8613 12604 8665 12649
rect 8721 12604 8773 12649
rect 8829 12604 8881 12649
rect 8937 12604 8989 12649
rect 9045 12604 9097 12649
rect 9153 12604 9205 12649
rect 9261 12604 9313 12649
rect 9369 12604 9421 12649
rect 9477 12604 9529 12649
rect 12051 12705 12103 12757
rect 12159 12705 12211 12757
rect 12267 12705 12319 12757
rect 1505 12597 1557 12604
rect 1613 12597 1665 12604
rect 1721 12597 1773 12604
rect 1829 12597 1881 12604
rect 1937 12597 1989 12604
rect 2045 12597 2097 12604
rect 2153 12597 2205 12604
rect 2261 12597 2313 12604
rect 2369 12597 2421 12604
rect 2477 12597 2529 12604
rect 2585 12597 2637 12604
rect 2693 12597 2745 12604
rect 2801 12597 2853 12604
rect 2909 12597 2961 12604
rect 3017 12597 3069 12604
rect 3125 12597 3177 12604
rect 3233 12597 3285 12604
rect 5372 12597 5424 12604
rect 5480 12597 5532 12604
rect 5588 12597 5640 12604
rect 5696 12597 5748 12604
rect 5804 12597 5856 12604
rect 5912 12597 5964 12604
rect 6020 12597 6072 12604
rect 6128 12597 6180 12604
rect 6236 12597 6288 12604
rect 6344 12597 6396 12604
rect 7749 12597 7801 12604
rect 7857 12597 7909 12604
rect 7965 12597 8017 12604
rect 8073 12597 8125 12604
rect 8181 12597 8233 12604
rect 8289 12597 8341 12604
rect 8397 12597 8449 12604
rect 8505 12597 8557 12604
rect 8613 12597 8665 12604
rect 8721 12597 8773 12604
rect 8829 12597 8881 12604
rect 8937 12597 8989 12604
rect 9045 12597 9097 12604
rect 9153 12597 9205 12604
rect 9261 12597 9313 12604
rect 9369 12597 9421 12604
rect 9477 12597 9529 12604
rect 12051 12597 12103 12649
rect 12159 12597 12211 12649
rect 12267 12597 12319 12649
rect 3433 12204 3485 12207
rect 3541 12204 3593 12207
rect 3649 12204 3701 12207
rect 3757 12204 3809 12207
rect 3865 12204 3917 12207
rect 3973 12204 4025 12207
rect 4081 12204 4133 12207
rect 4189 12204 4241 12207
rect 4297 12204 4349 12207
rect 4405 12204 4457 12207
rect 4513 12204 4565 12207
rect 4621 12204 4673 12207
rect 4729 12204 4781 12207
rect 4837 12204 4889 12207
rect 4945 12204 4997 12207
rect 5053 12204 5105 12207
rect 5161 12204 5213 12207
rect 6566 12204 6618 12207
rect 6674 12204 6726 12207
rect 6782 12204 6834 12207
rect 6890 12204 6942 12207
rect 6998 12204 7050 12207
rect 7106 12204 7158 12207
rect 7214 12204 7266 12207
rect 7322 12204 7374 12207
rect 7430 12204 7482 12207
rect 7538 12204 7590 12207
rect 9677 12204 9729 12207
rect 9785 12204 9837 12207
rect 9893 12204 9945 12207
rect 10001 12204 10053 12207
rect 10109 12204 10161 12207
rect 10217 12204 10269 12207
rect 10325 12204 10377 12207
rect 10433 12204 10485 12207
rect 10541 12204 10593 12207
rect 10649 12204 10701 12207
rect 10757 12204 10809 12207
rect 10865 12204 10917 12207
rect 10973 12204 11025 12207
rect 11081 12204 11133 12207
rect 11189 12204 11241 12207
rect 11297 12204 11349 12207
rect 11405 12204 11457 12207
rect 3433 12158 3485 12204
rect 3541 12158 3593 12204
rect 3649 12158 3701 12204
rect 3757 12158 3809 12204
rect 3865 12158 3917 12204
rect 3973 12158 4025 12204
rect 4081 12158 4133 12204
rect 4189 12158 4241 12204
rect 4297 12158 4349 12204
rect 4405 12158 4457 12204
rect 4513 12158 4565 12204
rect 4621 12158 4673 12204
rect 4729 12158 4781 12204
rect 4837 12158 4889 12204
rect 4945 12158 4997 12204
rect 5053 12158 5105 12204
rect 5161 12158 5213 12204
rect 6566 12158 6618 12204
rect 6674 12158 6726 12204
rect 6782 12158 6834 12204
rect 6890 12158 6942 12204
rect 6998 12158 7050 12204
rect 7106 12158 7158 12204
rect 7214 12158 7266 12204
rect 7322 12158 7374 12204
rect 7430 12158 7482 12204
rect 7538 12158 7590 12204
rect 9677 12158 9729 12204
rect 9785 12158 9837 12204
rect 9893 12158 9945 12204
rect 10001 12158 10053 12204
rect 10109 12158 10161 12204
rect 10217 12158 10269 12204
rect 10325 12158 10377 12204
rect 10433 12158 10485 12204
rect 10541 12158 10593 12204
rect 10649 12158 10701 12204
rect 10757 12158 10809 12204
rect 10865 12158 10917 12204
rect 10973 12158 11025 12204
rect 11081 12158 11133 12204
rect 11189 12158 11241 12204
rect 11297 12158 11349 12204
rect 11405 12158 11457 12204
rect 3433 12155 3485 12158
rect 3541 12155 3593 12158
rect 3649 12155 3701 12158
rect 3757 12155 3809 12158
rect 3865 12155 3917 12158
rect 3973 12155 4025 12158
rect 4081 12155 4133 12158
rect 4189 12155 4241 12158
rect 4297 12155 4349 12158
rect 4405 12155 4457 12158
rect 4513 12155 4565 12158
rect 4621 12155 4673 12158
rect 4729 12155 4781 12158
rect 4837 12155 4889 12158
rect 4945 12155 4997 12158
rect 5053 12155 5105 12158
rect 5161 12155 5213 12158
rect 6566 12155 6618 12158
rect 6674 12155 6726 12158
rect 6782 12155 6834 12158
rect 6890 12155 6942 12158
rect 6998 12155 7050 12158
rect 7106 12155 7158 12158
rect 7214 12155 7266 12158
rect 7322 12155 7374 12158
rect 7430 12155 7482 12158
rect 7538 12155 7590 12158
rect 9677 12155 9729 12158
rect 9785 12155 9837 12158
rect 9893 12155 9945 12158
rect 10001 12155 10053 12158
rect 10109 12155 10161 12158
rect 10217 12155 10269 12158
rect 10325 12155 10377 12158
rect 10433 12155 10485 12158
rect 10541 12155 10593 12158
rect 10649 12155 10701 12158
rect 10757 12155 10809 12158
rect 10865 12155 10917 12158
rect 10973 12155 11025 12158
rect 11081 12155 11133 12158
rect 11189 12155 11241 12158
rect 11297 12155 11349 12158
rect 11405 12155 11457 12158
rect 1233 12091 1285 12143
rect 1341 12091 1393 12143
rect 1233 11983 1256 12035
rect 1256 11983 1285 12035
rect 1341 11983 1393 12035
rect 1233 11875 1256 11927
rect 1256 11875 1285 11927
rect 1341 11875 1393 11927
rect 1233 11767 1256 11819
rect 1256 11767 1285 11819
rect 1341 11767 1393 11819
rect 1233 11659 1256 11711
rect 1256 11659 1285 11711
rect 1341 11659 1393 11711
rect 1233 11551 1256 11603
rect 1256 11551 1285 11603
rect 1341 11551 1393 11603
rect 1233 11443 1256 11495
rect 1256 11443 1285 11495
rect 1341 11443 1393 11495
rect 1233 11335 1256 11387
rect 1256 11335 1285 11387
rect 1341 11335 1393 11387
rect 1233 11227 1256 11279
rect 1256 11227 1285 11279
rect 1341 11227 1393 11279
rect 1233 11119 1256 11171
rect 1256 11119 1285 11171
rect 1341 11119 1393 11171
rect 1233 11011 1256 11063
rect 1256 11011 1285 11063
rect 1341 11011 1393 11063
rect 1233 10903 1256 10955
rect 1256 10903 1285 10955
rect 1341 10903 1393 10955
rect 1233 10795 1256 10847
rect 1256 10795 1285 10847
rect 1341 10795 1393 10847
rect 1233 10687 1256 10739
rect 1256 10687 1285 10739
rect 1341 10687 1393 10739
rect 1233 10579 1256 10631
rect 1256 10579 1285 10631
rect 1341 10579 1393 10631
rect 1233 10471 1256 10523
rect 1256 10471 1285 10523
rect 1341 10471 1393 10523
rect 1233 10363 1256 10415
rect 1256 10363 1285 10415
rect 1341 10363 1393 10415
rect 1233 10255 1256 10307
rect 1256 10255 1285 10307
rect 1341 10255 1393 10307
rect 1233 10147 1256 10199
rect 1256 10147 1285 10199
rect 1341 10147 1393 10199
rect 1233 10039 1256 10091
rect 1256 10039 1285 10091
rect 1341 10039 1393 10091
rect 1233 9931 1256 9983
rect 1256 9931 1285 9983
rect 1341 9931 1393 9983
rect 1233 9823 1256 9875
rect 1256 9823 1285 9875
rect 1341 9823 1393 9875
rect 1233 9715 1256 9767
rect 1256 9715 1285 9767
rect 1341 9715 1393 9767
rect 1233 9607 1256 9659
rect 1256 9607 1285 9659
rect 1341 9607 1393 9659
rect 1233 9499 1256 9551
rect 1256 9499 1285 9551
rect 1341 9499 1393 9551
rect 1233 9391 1256 9443
rect 1256 9391 1285 9443
rect 1341 9391 1393 9443
rect 1233 9283 1256 9335
rect 1256 9283 1285 9335
rect 1341 9283 1393 9335
rect 1233 9175 1256 9227
rect 1256 9175 1285 9227
rect 1341 9175 1393 9227
rect 1233 9067 1256 9119
rect 1256 9067 1285 9119
rect 1341 9067 1393 9119
rect 1233 8959 1256 9011
rect 1256 8959 1285 9011
rect 1341 8959 1393 9011
rect 1233 8851 1256 8903
rect 1256 8851 1285 8903
rect 1341 8851 1393 8903
rect 1233 8743 1256 8795
rect 1256 8743 1285 8795
rect 1341 8743 1393 8795
rect 1233 8635 1256 8687
rect 1256 8635 1285 8687
rect 1341 8635 1393 8687
rect 1233 8527 1256 8579
rect 1256 8527 1285 8579
rect 1341 8527 1393 8579
rect 1233 8419 1256 8471
rect 1256 8419 1285 8471
rect 1341 8419 1393 8471
rect 1233 8311 1256 8363
rect 1256 8311 1285 8363
rect 1341 8311 1393 8363
rect 1233 8203 1256 8255
rect 1256 8203 1285 8255
rect 1341 8203 1393 8255
rect 1233 8095 1256 8147
rect 1256 8095 1285 8147
rect 1341 8095 1393 8147
rect 1233 7987 1256 8039
rect 1256 7987 1285 8039
rect 1341 7987 1393 8039
rect 1233 7879 1256 7931
rect 1256 7879 1285 7931
rect 1341 7879 1393 7931
rect 1233 7771 1256 7823
rect 1256 7771 1285 7823
rect 1341 7771 1393 7823
rect 1233 7663 1256 7715
rect 1256 7663 1285 7715
rect 1341 7663 1393 7715
rect 1233 7555 1256 7607
rect 1256 7555 1285 7607
rect 1341 7555 1393 7607
rect 1233 7447 1256 7499
rect 1256 7447 1285 7499
rect 1341 7447 1393 7499
rect 11569 12091 11621 12143
rect 11677 12091 11729 12143
rect 1505 11960 1557 11963
rect 1613 11960 1665 11963
rect 1721 11960 1773 11963
rect 1829 11960 1881 11963
rect 1937 11960 1989 11963
rect 2045 11960 2097 11963
rect 2153 11960 2205 11963
rect 2261 11960 2313 11963
rect 2369 11960 2421 11963
rect 2477 11960 2529 11963
rect 2585 11960 2637 11963
rect 2693 11960 2745 11963
rect 2801 11960 2853 11963
rect 2909 11960 2961 11963
rect 3017 11960 3069 11963
rect 3125 11960 3177 11963
rect 3233 11960 3285 11963
rect 5372 11960 5424 11963
rect 5480 11960 5532 11963
rect 5588 11960 5640 11963
rect 5696 11960 5748 11963
rect 5804 11960 5856 11963
rect 5912 11960 5964 11963
rect 6020 11960 6072 11963
rect 6128 11960 6180 11963
rect 6236 11960 6288 11963
rect 6344 11960 6396 11963
rect 7749 11960 7801 11963
rect 7857 11960 7909 11963
rect 7965 11960 8017 11963
rect 8073 11960 8125 11963
rect 8181 11960 8233 11963
rect 8289 11960 8341 11963
rect 8397 11960 8449 11963
rect 8505 11960 8557 11963
rect 8613 11960 8665 11963
rect 8721 11960 8773 11963
rect 8829 11960 8881 11963
rect 8937 11960 8989 11963
rect 9045 11960 9097 11963
rect 9153 11960 9205 11963
rect 9261 11960 9313 11963
rect 9369 11960 9421 11963
rect 9477 11960 9529 11963
rect 1505 11914 1557 11960
rect 1613 11914 1665 11960
rect 1721 11914 1773 11960
rect 1829 11914 1881 11960
rect 1937 11914 1989 11960
rect 2045 11914 2097 11960
rect 2153 11914 2205 11960
rect 2261 11914 2313 11960
rect 2369 11914 2421 11960
rect 2477 11914 2529 11960
rect 2585 11914 2637 11960
rect 2693 11914 2745 11960
rect 2801 11914 2853 11960
rect 2909 11914 2961 11960
rect 3017 11914 3069 11960
rect 3125 11914 3177 11960
rect 3233 11914 3285 11960
rect 5372 11914 5424 11960
rect 5480 11914 5532 11960
rect 5588 11914 5640 11960
rect 5696 11914 5748 11960
rect 5804 11914 5856 11960
rect 5912 11914 5964 11960
rect 6020 11914 6072 11960
rect 6128 11914 6180 11960
rect 6236 11914 6288 11960
rect 6344 11914 6396 11960
rect 7749 11914 7801 11960
rect 7857 11914 7909 11960
rect 7965 11914 8017 11960
rect 8073 11914 8125 11960
rect 8181 11914 8233 11960
rect 8289 11914 8341 11960
rect 8397 11914 8449 11960
rect 8505 11914 8557 11960
rect 8613 11914 8665 11960
rect 8721 11914 8773 11960
rect 8829 11914 8881 11960
rect 8937 11914 8989 11960
rect 9045 11914 9097 11960
rect 9153 11914 9205 11960
rect 9261 11914 9313 11960
rect 9369 11914 9421 11960
rect 9477 11914 9529 11960
rect 1505 11911 1557 11914
rect 1613 11911 1665 11914
rect 1721 11911 1773 11914
rect 1829 11911 1881 11914
rect 1937 11911 1989 11914
rect 2045 11911 2097 11914
rect 2153 11911 2205 11914
rect 2261 11911 2313 11914
rect 2369 11911 2421 11914
rect 2477 11911 2529 11914
rect 2585 11911 2637 11914
rect 2693 11911 2745 11914
rect 2801 11911 2853 11914
rect 2909 11911 2961 11914
rect 3017 11911 3069 11914
rect 3125 11911 3177 11914
rect 3233 11911 3285 11914
rect 5372 11911 5424 11914
rect 5480 11911 5532 11914
rect 5588 11911 5640 11914
rect 5696 11911 5748 11914
rect 5804 11911 5856 11914
rect 5912 11911 5964 11914
rect 6020 11911 6072 11914
rect 6128 11911 6180 11914
rect 6236 11911 6288 11914
rect 6344 11911 6396 11914
rect 7749 11911 7801 11914
rect 7857 11911 7909 11914
rect 7965 11911 8017 11914
rect 8073 11911 8125 11914
rect 8181 11911 8233 11914
rect 8289 11911 8341 11914
rect 8397 11911 8449 11914
rect 8505 11911 8557 11914
rect 8613 11911 8665 11914
rect 8721 11911 8773 11914
rect 8829 11911 8881 11914
rect 8937 11911 8989 11914
rect 9045 11911 9097 11914
rect 9153 11911 9205 11914
rect 9261 11911 9313 11914
rect 9369 11911 9421 11914
rect 9477 11911 9529 11914
rect 3433 11716 3485 11719
rect 3541 11716 3593 11719
rect 3649 11716 3701 11719
rect 3757 11716 3809 11719
rect 3865 11716 3917 11719
rect 3973 11716 4025 11719
rect 4081 11716 4133 11719
rect 4189 11716 4241 11719
rect 4297 11716 4349 11719
rect 4405 11716 4457 11719
rect 4513 11716 4565 11719
rect 4621 11716 4673 11719
rect 4729 11716 4781 11719
rect 4837 11716 4889 11719
rect 4945 11716 4997 11719
rect 5053 11716 5105 11719
rect 5161 11716 5213 11719
rect 6566 11716 6618 11719
rect 6674 11716 6726 11719
rect 6782 11716 6834 11719
rect 6890 11716 6942 11719
rect 6998 11716 7050 11719
rect 7106 11716 7158 11719
rect 7214 11716 7266 11719
rect 7322 11716 7374 11719
rect 7430 11716 7482 11719
rect 7538 11716 7590 11719
rect 9677 11716 9729 11719
rect 9785 11716 9837 11719
rect 9893 11716 9945 11719
rect 10001 11716 10053 11719
rect 10109 11716 10161 11719
rect 10217 11716 10269 11719
rect 10325 11716 10377 11719
rect 10433 11716 10485 11719
rect 10541 11716 10593 11719
rect 10649 11716 10701 11719
rect 10757 11716 10809 11719
rect 10865 11716 10917 11719
rect 10973 11716 11025 11719
rect 11081 11716 11133 11719
rect 11189 11716 11241 11719
rect 11297 11716 11349 11719
rect 11405 11716 11457 11719
rect 3433 11670 3485 11716
rect 3541 11670 3593 11716
rect 3649 11670 3701 11716
rect 3757 11670 3809 11716
rect 3865 11670 3917 11716
rect 3973 11670 4025 11716
rect 4081 11670 4133 11716
rect 4189 11670 4241 11716
rect 4297 11670 4349 11716
rect 4405 11670 4457 11716
rect 4513 11670 4565 11716
rect 4621 11670 4673 11716
rect 4729 11670 4781 11716
rect 4837 11670 4889 11716
rect 4945 11670 4997 11716
rect 5053 11670 5105 11716
rect 5161 11670 5213 11716
rect 6566 11670 6618 11716
rect 6674 11670 6726 11716
rect 6782 11670 6834 11716
rect 6890 11670 6942 11716
rect 6998 11670 7050 11716
rect 7106 11670 7158 11716
rect 7214 11670 7266 11716
rect 7322 11670 7374 11716
rect 7430 11670 7482 11716
rect 7538 11670 7590 11716
rect 9677 11670 9729 11716
rect 9785 11670 9837 11716
rect 9893 11670 9945 11716
rect 10001 11670 10053 11716
rect 10109 11670 10161 11716
rect 10217 11670 10269 11716
rect 10325 11670 10377 11716
rect 10433 11670 10485 11716
rect 10541 11670 10593 11716
rect 10649 11670 10701 11716
rect 10757 11670 10809 11716
rect 10865 11670 10917 11716
rect 10973 11670 11025 11716
rect 11081 11670 11133 11716
rect 11189 11670 11241 11716
rect 11297 11670 11349 11716
rect 11405 11670 11457 11716
rect 3433 11667 3485 11670
rect 3541 11667 3593 11670
rect 3649 11667 3701 11670
rect 3757 11667 3809 11670
rect 3865 11667 3917 11670
rect 3973 11667 4025 11670
rect 4081 11667 4133 11670
rect 4189 11667 4241 11670
rect 4297 11667 4349 11670
rect 4405 11667 4457 11670
rect 4513 11667 4565 11670
rect 4621 11667 4673 11670
rect 4729 11667 4781 11670
rect 4837 11667 4889 11670
rect 4945 11667 4997 11670
rect 5053 11667 5105 11670
rect 5161 11667 5213 11670
rect 6566 11667 6618 11670
rect 6674 11667 6726 11670
rect 6782 11667 6834 11670
rect 6890 11667 6942 11670
rect 6998 11667 7050 11670
rect 7106 11667 7158 11670
rect 7214 11667 7266 11670
rect 7322 11667 7374 11670
rect 7430 11667 7482 11670
rect 7538 11667 7590 11670
rect 9677 11667 9729 11670
rect 9785 11667 9837 11670
rect 9893 11667 9945 11670
rect 10001 11667 10053 11670
rect 10109 11667 10161 11670
rect 10217 11667 10269 11670
rect 10325 11667 10377 11670
rect 10433 11667 10485 11670
rect 10541 11667 10593 11670
rect 10649 11667 10701 11670
rect 10757 11667 10809 11670
rect 10865 11667 10917 11670
rect 10973 11667 11025 11670
rect 11081 11667 11133 11670
rect 11189 11667 11241 11670
rect 11297 11667 11349 11670
rect 11405 11667 11457 11670
rect 1505 11472 1557 11475
rect 1613 11472 1665 11475
rect 1721 11472 1773 11475
rect 1829 11472 1881 11475
rect 1937 11472 1989 11475
rect 2045 11472 2097 11475
rect 2153 11472 2205 11475
rect 2261 11472 2313 11475
rect 2369 11472 2421 11475
rect 2477 11472 2529 11475
rect 2585 11472 2637 11475
rect 2693 11472 2745 11475
rect 2801 11472 2853 11475
rect 2909 11472 2961 11475
rect 3017 11472 3069 11475
rect 3125 11472 3177 11475
rect 3233 11472 3285 11475
rect 5372 11472 5424 11475
rect 5480 11472 5532 11475
rect 5588 11472 5640 11475
rect 5696 11472 5748 11475
rect 5804 11472 5856 11475
rect 5912 11472 5964 11475
rect 6020 11472 6072 11475
rect 6128 11472 6180 11475
rect 6236 11472 6288 11475
rect 6344 11472 6396 11475
rect 7749 11472 7801 11475
rect 7857 11472 7909 11475
rect 7965 11472 8017 11475
rect 8073 11472 8125 11475
rect 8181 11472 8233 11475
rect 8289 11472 8341 11475
rect 8397 11472 8449 11475
rect 8505 11472 8557 11475
rect 8613 11472 8665 11475
rect 8721 11472 8773 11475
rect 8829 11472 8881 11475
rect 8937 11472 8989 11475
rect 9045 11472 9097 11475
rect 9153 11472 9205 11475
rect 9261 11472 9313 11475
rect 9369 11472 9421 11475
rect 9477 11472 9529 11475
rect 1505 11426 1557 11472
rect 1613 11426 1665 11472
rect 1721 11426 1773 11472
rect 1829 11426 1881 11472
rect 1937 11426 1989 11472
rect 2045 11426 2097 11472
rect 2153 11426 2205 11472
rect 2261 11426 2313 11472
rect 2369 11426 2421 11472
rect 2477 11426 2529 11472
rect 2585 11426 2637 11472
rect 2693 11426 2745 11472
rect 2801 11426 2853 11472
rect 2909 11426 2961 11472
rect 3017 11426 3069 11472
rect 3125 11426 3177 11472
rect 3233 11426 3285 11472
rect 5372 11426 5424 11472
rect 5480 11426 5532 11472
rect 5588 11426 5640 11472
rect 5696 11426 5748 11472
rect 5804 11426 5856 11472
rect 5912 11426 5964 11472
rect 6020 11426 6072 11472
rect 6128 11426 6180 11472
rect 6236 11426 6288 11472
rect 6344 11426 6396 11472
rect 7749 11426 7801 11472
rect 7857 11426 7909 11472
rect 7965 11426 8017 11472
rect 8073 11426 8125 11472
rect 8181 11426 8233 11472
rect 8289 11426 8341 11472
rect 8397 11426 8449 11472
rect 8505 11426 8557 11472
rect 8613 11426 8665 11472
rect 8721 11426 8773 11472
rect 8829 11426 8881 11472
rect 8937 11426 8989 11472
rect 9045 11426 9097 11472
rect 9153 11426 9205 11472
rect 9261 11426 9313 11472
rect 9369 11426 9421 11472
rect 9477 11426 9529 11472
rect 1505 11423 1557 11426
rect 1613 11423 1665 11426
rect 1721 11423 1773 11426
rect 1829 11423 1881 11426
rect 1937 11423 1989 11426
rect 2045 11423 2097 11426
rect 2153 11423 2205 11426
rect 2261 11423 2313 11426
rect 2369 11423 2421 11426
rect 2477 11423 2529 11426
rect 2585 11423 2637 11426
rect 2693 11423 2745 11426
rect 2801 11423 2853 11426
rect 2909 11423 2961 11426
rect 3017 11423 3069 11426
rect 3125 11423 3177 11426
rect 3233 11423 3285 11426
rect 5372 11423 5424 11426
rect 5480 11423 5532 11426
rect 5588 11423 5640 11426
rect 5696 11423 5748 11426
rect 5804 11423 5856 11426
rect 5912 11423 5964 11426
rect 6020 11423 6072 11426
rect 6128 11423 6180 11426
rect 6236 11423 6288 11426
rect 6344 11423 6396 11426
rect 7749 11423 7801 11426
rect 7857 11423 7909 11426
rect 7965 11423 8017 11426
rect 8073 11423 8125 11426
rect 8181 11423 8233 11426
rect 8289 11423 8341 11426
rect 8397 11423 8449 11426
rect 8505 11423 8557 11426
rect 8613 11423 8665 11426
rect 8721 11423 8773 11426
rect 8829 11423 8881 11426
rect 8937 11423 8989 11426
rect 9045 11423 9097 11426
rect 9153 11423 9205 11426
rect 9261 11423 9313 11426
rect 9369 11423 9421 11426
rect 9477 11423 9529 11426
rect 3433 11228 3485 11231
rect 3541 11228 3593 11231
rect 3649 11228 3701 11231
rect 3757 11228 3809 11231
rect 3865 11228 3917 11231
rect 3973 11228 4025 11231
rect 4081 11228 4133 11231
rect 4189 11228 4241 11231
rect 4297 11228 4349 11231
rect 4405 11228 4457 11231
rect 4513 11228 4565 11231
rect 4621 11228 4673 11231
rect 4729 11228 4781 11231
rect 4837 11228 4889 11231
rect 4945 11228 4997 11231
rect 5053 11228 5105 11231
rect 5161 11228 5213 11231
rect 6566 11228 6618 11231
rect 6674 11228 6726 11231
rect 6782 11228 6834 11231
rect 6890 11228 6942 11231
rect 6998 11228 7050 11231
rect 7106 11228 7158 11231
rect 7214 11228 7266 11231
rect 7322 11228 7374 11231
rect 7430 11228 7482 11231
rect 7538 11228 7590 11231
rect 9677 11228 9729 11231
rect 9785 11228 9837 11231
rect 9893 11228 9945 11231
rect 10001 11228 10053 11231
rect 10109 11228 10161 11231
rect 10217 11228 10269 11231
rect 10325 11228 10377 11231
rect 10433 11228 10485 11231
rect 10541 11228 10593 11231
rect 10649 11228 10701 11231
rect 10757 11228 10809 11231
rect 10865 11228 10917 11231
rect 10973 11228 11025 11231
rect 11081 11228 11133 11231
rect 11189 11228 11241 11231
rect 11297 11228 11349 11231
rect 11405 11228 11457 11231
rect 3433 11182 3485 11228
rect 3541 11182 3593 11228
rect 3649 11182 3701 11228
rect 3757 11182 3809 11228
rect 3865 11182 3917 11228
rect 3973 11182 4025 11228
rect 4081 11182 4133 11228
rect 4189 11182 4241 11228
rect 4297 11182 4349 11228
rect 4405 11182 4457 11228
rect 4513 11182 4565 11228
rect 4621 11182 4673 11228
rect 4729 11182 4781 11228
rect 4837 11182 4889 11228
rect 4945 11182 4997 11228
rect 5053 11182 5105 11228
rect 5161 11182 5213 11228
rect 6566 11182 6618 11228
rect 6674 11182 6726 11228
rect 6782 11182 6834 11228
rect 6890 11182 6942 11228
rect 6998 11182 7050 11228
rect 7106 11182 7158 11228
rect 7214 11182 7266 11228
rect 7322 11182 7374 11228
rect 7430 11182 7482 11228
rect 7538 11182 7590 11228
rect 9677 11182 9729 11228
rect 9785 11182 9837 11228
rect 9893 11182 9945 11228
rect 10001 11182 10053 11228
rect 10109 11182 10161 11228
rect 10217 11182 10269 11228
rect 10325 11182 10377 11228
rect 10433 11182 10485 11228
rect 10541 11182 10593 11228
rect 10649 11182 10701 11228
rect 10757 11182 10809 11228
rect 10865 11182 10917 11228
rect 10973 11182 11025 11228
rect 11081 11182 11133 11228
rect 11189 11182 11241 11228
rect 11297 11182 11349 11228
rect 11405 11182 11457 11228
rect 3433 11179 3485 11182
rect 3541 11179 3593 11182
rect 3649 11179 3701 11182
rect 3757 11179 3809 11182
rect 3865 11179 3917 11182
rect 3973 11179 4025 11182
rect 4081 11179 4133 11182
rect 4189 11179 4241 11182
rect 4297 11179 4349 11182
rect 4405 11179 4457 11182
rect 4513 11179 4565 11182
rect 4621 11179 4673 11182
rect 4729 11179 4781 11182
rect 4837 11179 4889 11182
rect 4945 11179 4997 11182
rect 5053 11179 5105 11182
rect 5161 11179 5213 11182
rect 6566 11179 6618 11182
rect 6674 11179 6726 11182
rect 6782 11179 6834 11182
rect 6890 11179 6942 11182
rect 6998 11179 7050 11182
rect 7106 11179 7158 11182
rect 7214 11179 7266 11182
rect 7322 11179 7374 11182
rect 7430 11179 7482 11182
rect 7538 11179 7590 11182
rect 9677 11179 9729 11182
rect 9785 11179 9837 11182
rect 9893 11179 9945 11182
rect 10001 11179 10053 11182
rect 10109 11179 10161 11182
rect 10217 11179 10269 11182
rect 10325 11179 10377 11182
rect 10433 11179 10485 11182
rect 10541 11179 10593 11182
rect 10649 11179 10701 11182
rect 10757 11179 10809 11182
rect 10865 11179 10917 11182
rect 10973 11179 11025 11182
rect 11081 11179 11133 11182
rect 11189 11179 11241 11182
rect 11297 11179 11349 11182
rect 11405 11179 11457 11182
rect 1505 10984 1557 10987
rect 1613 10984 1665 10987
rect 1721 10984 1773 10987
rect 1829 10984 1881 10987
rect 1937 10984 1989 10987
rect 2045 10984 2097 10987
rect 2153 10984 2205 10987
rect 2261 10984 2313 10987
rect 2369 10984 2421 10987
rect 2477 10984 2529 10987
rect 2585 10984 2637 10987
rect 2693 10984 2745 10987
rect 2801 10984 2853 10987
rect 2909 10984 2961 10987
rect 3017 10984 3069 10987
rect 3125 10984 3177 10987
rect 3233 10984 3285 10987
rect 5372 10984 5424 10987
rect 5480 10984 5532 10987
rect 5588 10984 5640 10987
rect 5696 10984 5748 10987
rect 5804 10984 5856 10987
rect 5912 10984 5964 10987
rect 6020 10984 6072 10987
rect 6128 10984 6180 10987
rect 6236 10984 6288 10987
rect 6344 10984 6396 10987
rect 7749 10984 7801 10987
rect 7857 10984 7909 10987
rect 7965 10984 8017 10987
rect 8073 10984 8125 10987
rect 8181 10984 8233 10987
rect 8289 10984 8341 10987
rect 8397 10984 8449 10987
rect 8505 10984 8557 10987
rect 8613 10984 8665 10987
rect 8721 10984 8773 10987
rect 8829 10984 8881 10987
rect 8937 10984 8989 10987
rect 9045 10984 9097 10987
rect 9153 10984 9205 10987
rect 9261 10984 9313 10987
rect 9369 10984 9421 10987
rect 9477 10984 9529 10987
rect 1505 10938 1557 10984
rect 1613 10938 1665 10984
rect 1721 10938 1773 10984
rect 1829 10938 1881 10984
rect 1937 10938 1989 10984
rect 2045 10938 2097 10984
rect 2153 10938 2205 10984
rect 2261 10938 2313 10984
rect 2369 10938 2421 10984
rect 2477 10938 2529 10984
rect 2585 10938 2637 10984
rect 2693 10938 2745 10984
rect 2801 10938 2853 10984
rect 2909 10938 2961 10984
rect 3017 10938 3069 10984
rect 3125 10938 3177 10984
rect 3233 10938 3285 10984
rect 5372 10938 5424 10984
rect 5480 10938 5532 10984
rect 5588 10938 5640 10984
rect 5696 10938 5748 10984
rect 5804 10938 5856 10984
rect 5912 10938 5964 10984
rect 6020 10938 6072 10984
rect 6128 10938 6180 10984
rect 6236 10938 6288 10984
rect 6344 10938 6396 10984
rect 7749 10938 7801 10984
rect 7857 10938 7909 10984
rect 7965 10938 8017 10984
rect 8073 10938 8125 10984
rect 8181 10938 8233 10984
rect 8289 10938 8341 10984
rect 8397 10938 8449 10984
rect 8505 10938 8557 10984
rect 8613 10938 8665 10984
rect 8721 10938 8773 10984
rect 8829 10938 8881 10984
rect 8937 10938 8989 10984
rect 9045 10938 9097 10984
rect 9153 10938 9205 10984
rect 9261 10938 9313 10984
rect 9369 10938 9421 10984
rect 9477 10938 9529 10984
rect 1505 10935 1557 10938
rect 1613 10935 1665 10938
rect 1721 10935 1773 10938
rect 1829 10935 1881 10938
rect 1937 10935 1989 10938
rect 2045 10935 2097 10938
rect 2153 10935 2205 10938
rect 2261 10935 2313 10938
rect 2369 10935 2421 10938
rect 2477 10935 2529 10938
rect 2585 10935 2637 10938
rect 2693 10935 2745 10938
rect 2801 10935 2853 10938
rect 2909 10935 2961 10938
rect 3017 10935 3069 10938
rect 3125 10935 3177 10938
rect 3233 10935 3285 10938
rect 5372 10935 5424 10938
rect 5480 10935 5532 10938
rect 5588 10935 5640 10938
rect 5696 10935 5748 10938
rect 5804 10935 5856 10938
rect 5912 10935 5964 10938
rect 6020 10935 6072 10938
rect 6128 10935 6180 10938
rect 6236 10935 6288 10938
rect 6344 10935 6396 10938
rect 7749 10935 7801 10938
rect 7857 10935 7909 10938
rect 7965 10935 8017 10938
rect 8073 10935 8125 10938
rect 8181 10935 8233 10938
rect 8289 10935 8341 10938
rect 8397 10935 8449 10938
rect 8505 10935 8557 10938
rect 8613 10935 8665 10938
rect 8721 10935 8773 10938
rect 8829 10935 8881 10938
rect 8937 10935 8989 10938
rect 9045 10935 9097 10938
rect 9153 10935 9205 10938
rect 9261 10935 9313 10938
rect 9369 10935 9421 10938
rect 9477 10935 9529 10938
rect 3433 10740 3485 10743
rect 3541 10740 3593 10743
rect 3649 10740 3701 10743
rect 3757 10740 3809 10743
rect 3865 10740 3917 10743
rect 3973 10740 4025 10743
rect 4081 10740 4133 10743
rect 4189 10740 4241 10743
rect 4297 10740 4349 10743
rect 4405 10740 4457 10743
rect 4513 10740 4565 10743
rect 4621 10740 4673 10743
rect 4729 10740 4781 10743
rect 4837 10740 4889 10743
rect 4945 10740 4997 10743
rect 5053 10740 5105 10743
rect 5161 10740 5213 10743
rect 6566 10740 6618 10743
rect 6674 10740 6726 10743
rect 6782 10740 6834 10743
rect 6890 10740 6942 10743
rect 6998 10740 7050 10743
rect 7106 10740 7158 10743
rect 7214 10740 7266 10743
rect 7322 10740 7374 10743
rect 7430 10740 7482 10743
rect 7538 10740 7590 10743
rect 9677 10740 9729 10743
rect 9785 10740 9837 10743
rect 9893 10740 9945 10743
rect 10001 10740 10053 10743
rect 10109 10740 10161 10743
rect 10217 10740 10269 10743
rect 10325 10740 10377 10743
rect 10433 10740 10485 10743
rect 10541 10740 10593 10743
rect 10649 10740 10701 10743
rect 10757 10740 10809 10743
rect 10865 10740 10917 10743
rect 10973 10740 11025 10743
rect 11081 10740 11133 10743
rect 11189 10740 11241 10743
rect 11297 10740 11349 10743
rect 11405 10740 11457 10743
rect 3433 10694 3485 10740
rect 3541 10694 3593 10740
rect 3649 10694 3701 10740
rect 3757 10694 3809 10740
rect 3865 10694 3917 10740
rect 3973 10694 4025 10740
rect 4081 10694 4133 10740
rect 4189 10694 4241 10740
rect 4297 10694 4349 10740
rect 4405 10694 4457 10740
rect 4513 10694 4565 10740
rect 4621 10694 4673 10740
rect 4729 10694 4781 10740
rect 4837 10694 4889 10740
rect 4945 10694 4997 10740
rect 5053 10694 5105 10740
rect 5161 10694 5213 10740
rect 6566 10694 6618 10740
rect 6674 10694 6726 10740
rect 6782 10694 6834 10740
rect 6890 10694 6942 10740
rect 6998 10694 7050 10740
rect 7106 10694 7158 10740
rect 7214 10694 7266 10740
rect 7322 10694 7374 10740
rect 7430 10694 7482 10740
rect 7538 10694 7590 10740
rect 9677 10694 9729 10740
rect 9785 10694 9837 10740
rect 9893 10694 9945 10740
rect 10001 10694 10053 10740
rect 10109 10694 10161 10740
rect 10217 10694 10269 10740
rect 10325 10694 10377 10740
rect 10433 10694 10485 10740
rect 10541 10694 10593 10740
rect 10649 10694 10701 10740
rect 10757 10694 10809 10740
rect 10865 10694 10917 10740
rect 10973 10694 11025 10740
rect 11081 10694 11133 10740
rect 11189 10694 11241 10740
rect 11297 10694 11349 10740
rect 11405 10694 11457 10740
rect 3433 10691 3485 10694
rect 3541 10691 3593 10694
rect 3649 10691 3701 10694
rect 3757 10691 3809 10694
rect 3865 10691 3917 10694
rect 3973 10691 4025 10694
rect 4081 10691 4133 10694
rect 4189 10691 4241 10694
rect 4297 10691 4349 10694
rect 4405 10691 4457 10694
rect 4513 10691 4565 10694
rect 4621 10691 4673 10694
rect 4729 10691 4781 10694
rect 4837 10691 4889 10694
rect 4945 10691 4997 10694
rect 5053 10691 5105 10694
rect 5161 10691 5213 10694
rect 6566 10691 6618 10694
rect 6674 10691 6726 10694
rect 6782 10691 6834 10694
rect 6890 10691 6942 10694
rect 6998 10691 7050 10694
rect 7106 10691 7158 10694
rect 7214 10691 7266 10694
rect 7322 10691 7374 10694
rect 7430 10691 7482 10694
rect 7538 10691 7590 10694
rect 9677 10691 9729 10694
rect 9785 10691 9837 10694
rect 9893 10691 9945 10694
rect 10001 10691 10053 10694
rect 10109 10691 10161 10694
rect 10217 10691 10269 10694
rect 10325 10691 10377 10694
rect 10433 10691 10485 10694
rect 10541 10691 10593 10694
rect 10649 10691 10701 10694
rect 10757 10691 10809 10694
rect 10865 10691 10917 10694
rect 10973 10691 11025 10694
rect 11081 10691 11133 10694
rect 11189 10691 11241 10694
rect 11297 10691 11349 10694
rect 11405 10691 11457 10694
rect 1505 10496 1557 10499
rect 1613 10496 1665 10499
rect 1721 10496 1773 10499
rect 1829 10496 1881 10499
rect 1937 10496 1989 10499
rect 2045 10496 2097 10499
rect 2153 10496 2205 10499
rect 2261 10496 2313 10499
rect 2369 10496 2421 10499
rect 2477 10496 2529 10499
rect 2585 10496 2637 10499
rect 2693 10496 2745 10499
rect 2801 10496 2853 10499
rect 2909 10496 2961 10499
rect 3017 10496 3069 10499
rect 3125 10496 3177 10499
rect 3233 10496 3285 10499
rect 5372 10496 5424 10499
rect 5480 10496 5532 10499
rect 5588 10496 5640 10499
rect 5696 10496 5748 10499
rect 5804 10496 5856 10499
rect 5912 10496 5964 10499
rect 6020 10496 6072 10499
rect 6128 10496 6180 10499
rect 6236 10496 6288 10499
rect 6344 10496 6396 10499
rect 7749 10496 7801 10499
rect 7857 10496 7909 10499
rect 7965 10496 8017 10499
rect 8073 10496 8125 10499
rect 8181 10496 8233 10499
rect 8289 10496 8341 10499
rect 8397 10496 8449 10499
rect 8505 10496 8557 10499
rect 8613 10496 8665 10499
rect 8721 10496 8773 10499
rect 8829 10496 8881 10499
rect 8937 10496 8989 10499
rect 9045 10496 9097 10499
rect 9153 10496 9205 10499
rect 9261 10496 9313 10499
rect 9369 10496 9421 10499
rect 9477 10496 9529 10499
rect 1505 10450 1557 10496
rect 1613 10450 1665 10496
rect 1721 10450 1773 10496
rect 1829 10450 1881 10496
rect 1937 10450 1989 10496
rect 2045 10450 2097 10496
rect 2153 10450 2205 10496
rect 2261 10450 2313 10496
rect 2369 10450 2421 10496
rect 2477 10450 2529 10496
rect 2585 10450 2637 10496
rect 2693 10450 2745 10496
rect 2801 10450 2853 10496
rect 2909 10450 2961 10496
rect 3017 10450 3069 10496
rect 3125 10450 3177 10496
rect 3233 10450 3285 10496
rect 5372 10450 5424 10496
rect 5480 10450 5532 10496
rect 5588 10450 5640 10496
rect 5696 10450 5748 10496
rect 5804 10450 5856 10496
rect 5912 10450 5964 10496
rect 6020 10450 6072 10496
rect 6128 10450 6180 10496
rect 6236 10450 6288 10496
rect 6344 10450 6396 10496
rect 7749 10450 7801 10496
rect 7857 10450 7909 10496
rect 7965 10450 8017 10496
rect 8073 10450 8125 10496
rect 8181 10450 8233 10496
rect 8289 10450 8341 10496
rect 8397 10450 8449 10496
rect 8505 10450 8557 10496
rect 8613 10450 8665 10496
rect 8721 10450 8773 10496
rect 8829 10450 8881 10496
rect 8937 10450 8989 10496
rect 9045 10450 9097 10496
rect 9153 10450 9205 10496
rect 9261 10450 9313 10496
rect 9369 10450 9421 10496
rect 9477 10450 9529 10496
rect 1505 10447 1557 10450
rect 1613 10447 1665 10450
rect 1721 10447 1773 10450
rect 1829 10447 1881 10450
rect 1937 10447 1989 10450
rect 2045 10447 2097 10450
rect 2153 10447 2205 10450
rect 2261 10447 2313 10450
rect 2369 10447 2421 10450
rect 2477 10447 2529 10450
rect 2585 10447 2637 10450
rect 2693 10447 2745 10450
rect 2801 10447 2853 10450
rect 2909 10447 2961 10450
rect 3017 10447 3069 10450
rect 3125 10447 3177 10450
rect 3233 10447 3285 10450
rect 5372 10447 5424 10450
rect 5480 10447 5532 10450
rect 5588 10447 5640 10450
rect 5696 10447 5748 10450
rect 5804 10447 5856 10450
rect 5912 10447 5964 10450
rect 6020 10447 6072 10450
rect 6128 10447 6180 10450
rect 6236 10447 6288 10450
rect 6344 10447 6396 10450
rect 7749 10447 7801 10450
rect 7857 10447 7909 10450
rect 7965 10447 8017 10450
rect 8073 10447 8125 10450
rect 8181 10447 8233 10450
rect 8289 10447 8341 10450
rect 8397 10447 8449 10450
rect 8505 10447 8557 10450
rect 8613 10447 8665 10450
rect 8721 10447 8773 10450
rect 8829 10447 8881 10450
rect 8937 10447 8989 10450
rect 9045 10447 9097 10450
rect 9153 10447 9205 10450
rect 9261 10447 9313 10450
rect 9369 10447 9421 10450
rect 9477 10447 9529 10450
rect 3433 10252 3485 10255
rect 3541 10252 3593 10255
rect 3649 10252 3701 10255
rect 3757 10252 3809 10255
rect 3865 10252 3917 10255
rect 3973 10252 4025 10255
rect 4081 10252 4133 10255
rect 4189 10252 4241 10255
rect 4297 10252 4349 10255
rect 4405 10252 4457 10255
rect 4513 10252 4565 10255
rect 4621 10252 4673 10255
rect 4729 10252 4781 10255
rect 4837 10252 4889 10255
rect 4945 10252 4997 10255
rect 5053 10252 5105 10255
rect 5161 10252 5213 10255
rect 6566 10252 6618 10255
rect 6674 10252 6726 10255
rect 6782 10252 6834 10255
rect 6890 10252 6942 10255
rect 6998 10252 7050 10255
rect 7106 10252 7158 10255
rect 7214 10252 7266 10255
rect 7322 10252 7374 10255
rect 7430 10252 7482 10255
rect 7538 10252 7590 10255
rect 9677 10252 9729 10255
rect 9785 10252 9837 10255
rect 9893 10252 9945 10255
rect 10001 10252 10053 10255
rect 10109 10252 10161 10255
rect 10217 10252 10269 10255
rect 10325 10252 10377 10255
rect 10433 10252 10485 10255
rect 10541 10252 10593 10255
rect 10649 10252 10701 10255
rect 10757 10252 10809 10255
rect 10865 10252 10917 10255
rect 10973 10252 11025 10255
rect 11081 10252 11133 10255
rect 11189 10252 11241 10255
rect 11297 10252 11349 10255
rect 11405 10252 11457 10255
rect 3433 10206 3485 10252
rect 3541 10206 3593 10252
rect 3649 10206 3701 10252
rect 3757 10206 3809 10252
rect 3865 10206 3917 10252
rect 3973 10206 4025 10252
rect 4081 10206 4133 10252
rect 4189 10206 4241 10252
rect 4297 10206 4349 10252
rect 4405 10206 4457 10252
rect 4513 10206 4565 10252
rect 4621 10206 4673 10252
rect 4729 10206 4781 10252
rect 4837 10206 4889 10252
rect 4945 10206 4997 10252
rect 5053 10206 5105 10252
rect 5161 10206 5213 10252
rect 6566 10206 6618 10252
rect 6674 10206 6726 10252
rect 6782 10206 6834 10252
rect 6890 10206 6942 10252
rect 6998 10206 7050 10252
rect 7106 10206 7158 10252
rect 7214 10206 7266 10252
rect 7322 10206 7374 10252
rect 7430 10206 7482 10252
rect 7538 10206 7590 10252
rect 9677 10206 9729 10252
rect 9785 10206 9837 10252
rect 9893 10206 9945 10252
rect 10001 10206 10053 10252
rect 10109 10206 10161 10252
rect 10217 10206 10269 10252
rect 10325 10206 10377 10252
rect 10433 10206 10485 10252
rect 10541 10206 10593 10252
rect 10649 10206 10701 10252
rect 10757 10206 10809 10252
rect 10865 10206 10917 10252
rect 10973 10206 11025 10252
rect 11081 10206 11133 10252
rect 11189 10206 11241 10252
rect 11297 10206 11349 10252
rect 11405 10206 11457 10252
rect 3433 10203 3485 10206
rect 3541 10203 3593 10206
rect 3649 10203 3701 10206
rect 3757 10203 3809 10206
rect 3865 10203 3917 10206
rect 3973 10203 4025 10206
rect 4081 10203 4133 10206
rect 4189 10203 4241 10206
rect 4297 10203 4349 10206
rect 4405 10203 4457 10206
rect 4513 10203 4565 10206
rect 4621 10203 4673 10206
rect 4729 10203 4781 10206
rect 4837 10203 4889 10206
rect 4945 10203 4997 10206
rect 5053 10203 5105 10206
rect 5161 10203 5213 10206
rect 6566 10203 6618 10206
rect 6674 10203 6726 10206
rect 6782 10203 6834 10206
rect 6890 10203 6942 10206
rect 6998 10203 7050 10206
rect 7106 10203 7158 10206
rect 7214 10203 7266 10206
rect 7322 10203 7374 10206
rect 7430 10203 7482 10206
rect 7538 10203 7590 10206
rect 9677 10203 9729 10206
rect 9785 10203 9837 10206
rect 9893 10203 9945 10206
rect 10001 10203 10053 10206
rect 10109 10203 10161 10206
rect 10217 10203 10269 10206
rect 10325 10203 10377 10206
rect 10433 10203 10485 10206
rect 10541 10203 10593 10206
rect 10649 10203 10701 10206
rect 10757 10203 10809 10206
rect 10865 10203 10917 10206
rect 10973 10203 11025 10206
rect 11081 10203 11133 10206
rect 11189 10203 11241 10206
rect 11297 10203 11349 10206
rect 11405 10203 11457 10206
rect 1505 10008 1557 10011
rect 1613 10008 1665 10011
rect 1721 10008 1773 10011
rect 1829 10008 1881 10011
rect 1937 10008 1989 10011
rect 2045 10008 2097 10011
rect 2153 10008 2205 10011
rect 2261 10008 2313 10011
rect 2369 10008 2421 10011
rect 2477 10008 2529 10011
rect 2585 10008 2637 10011
rect 2693 10008 2745 10011
rect 2801 10008 2853 10011
rect 2909 10008 2961 10011
rect 3017 10008 3069 10011
rect 3125 10008 3177 10011
rect 3233 10008 3285 10011
rect 5372 10008 5424 10011
rect 5480 10008 5532 10011
rect 5588 10008 5640 10011
rect 5696 10008 5748 10011
rect 5804 10008 5856 10011
rect 5912 10008 5964 10011
rect 6020 10008 6072 10011
rect 6128 10008 6180 10011
rect 6236 10008 6288 10011
rect 6344 10008 6396 10011
rect 7749 10008 7801 10011
rect 7857 10008 7909 10011
rect 7965 10008 8017 10011
rect 8073 10008 8125 10011
rect 8181 10008 8233 10011
rect 8289 10008 8341 10011
rect 8397 10008 8449 10011
rect 8505 10008 8557 10011
rect 8613 10008 8665 10011
rect 8721 10008 8773 10011
rect 8829 10008 8881 10011
rect 8937 10008 8989 10011
rect 9045 10008 9097 10011
rect 9153 10008 9205 10011
rect 9261 10008 9313 10011
rect 9369 10008 9421 10011
rect 9477 10008 9529 10011
rect 1505 9962 1557 10008
rect 1613 9962 1665 10008
rect 1721 9962 1773 10008
rect 1829 9962 1881 10008
rect 1937 9962 1989 10008
rect 2045 9962 2097 10008
rect 2153 9962 2205 10008
rect 2261 9962 2313 10008
rect 2369 9962 2421 10008
rect 2477 9962 2529 10008
rect 2585 9962 2637 10008
rect 2693 9962 2745 10008
rect 2801 9962 2853 10008
rect 2909 9962 2961 10008
rect 3017 9962 3069 10008
rect 3125 9962 3177 10008
rect 3233 9962 3285 10008
rect 5372 9962 5424 10008
rect 5480 9962 5532 10008
rect 5588 9962 5640 10008
rect 5696 9962 5748 10008
rect 5804 9962 5856 10008
rect 5912 9962 5964 10008
rect 6020 9962 6072 10008
rect 6128 9962 6180 10008
rect 6236 9962 6288 10008
rect 6344 9962 6396 10008
rect 7749 9962 7801 10008
rect 7857 9962 7909 10008
rect 7965 9962 8017 10008
rect 8073 9962 8125 10008
rect 8181 9962 8233 10008
rect 8289 9962 8341 10008
rect 8397 9962 8449 10008
rect 8505 9962 8557 10008
rect 8613 9962 8665 10008
rect 8721 9962 8773 10008
rect 8829 9962 8881 10008
rect 8937 9962 8989 10008
rect 9045 9962 9097 10008
rect 9153 9962 9205 10008
rect 9261 9962 9313 10008
rect 9369 9962 9421 10008
rect 9477 9962 9529 10008
rect 1505 9959 1557 9962
rect 1613 9959 1665 9962
rect 1721 9959 1773 9962
rect 1829 9959 1881 9962
rect 1937 9959 1989 9962
rect 2045 9959 2097 9962
rect 2153 9959 2205 9962
rect 2261 9959 2313 9962
rect 2369 9959 2421 9962
rect 2477 9959 2529 9962
rect 2585 9959 2637 9962
rect 2693 9959 2745 9962
rect 2801 9959 2853 9962
rect 2909 9959 2961 9962
rect 3017 9959 3069 9962
rect 3125 9959 3177 9962
rect 3233 9959 3285 9962
rect 5372 9959 5424 9962
rect 5480 9959 5532 9962
rect 5588 9959 5640 9962
rect 5696 9959 5748 9962
rect 5804 9959 5856 9962
rect 5912 9959 5964 9962
rect 6020 9959 6072 9962
rect 6128 9959 6180 9962
rect 6236 9959 6288 9962
rect 6344 9959 6396 9962
rect 7749 9959 7801 9962
rect 7857 9959 7909 9962
rect 7965 9959 8017 9962
rect 8073 9959 8125 9962
rect 8181 9959 8233 9962
rect 8289 9959 8341 9962
rect 8397 9959 8449 9962
rect 8505 9959 8557 9962
rect 8613 9959 8665 9962
rect 8721 9959 8773 9962
rect 8829 9959 8881 9962
rect 8937 9959 8989 9962
rect 9045 9959 9097 9962
rect 9153 9959 9205 9962
rect 9261 9959 9313 9962
rect 9369 9959 9421 9962
rect 9477 9959 9529 9962
rect 3433 9764 3485 9767
rect 3541 9764 3593 9767
rect 3649 9764 3701 9767
rect 3757 9764 3809 9767
rect 3865 9764 3917 9767
rect 3973 9764 4025 9767
rect 4081 9764 4133 9767
rect 4189 9764 4241 9767
rect 4297 9764 4349 9767
rect 4405 9764 4457 9767
rect 4513 9764 4565 9767
rect 4621 9764 4673 9767
rect 4729 9764 4781 9767
rect 4837 9764 4889 9767
rect 4945 9764 4997 9767
rect 5053 9764 5105 9767
rect 5161 9764 5213 9767
rect 6566 9764 6618 9767
rect 6674 9764 6726 9767
rect 6782 9764 6834 9767
rect 6890 9764 6942 9767
rect 6998 9764 7050 9767
rect 7106 9764 7158 9767
rect 7214 9764 7266 9767
rect 7322 9764 7374 9767
rect 7430 9764 7482 9767
rect 7538 9764 7590 9767
rect 9677 9764 9729 9767
rect 9785 9764 9837 9767
rect 9893 9764 9945 9767
rect 10001 9764 10053 9767
rect 10109 9764 10161 9767
rect 10217 9764 10269 9767
rect 10325 9764 10377 9767
rect 10433 9764 10485 9767
rect 10541 9764 10593 9767
rect 10649 9764 10701 9767
rect 10757 9764 10809 9767
rect 10865 9764 10917 9767
rect 10973 9764 11025 9767
rect 11081 9764 11133 9767
rect 11189 9764 11241 9767
rect 11297 9764 11349 9767
rect 11405 9764 11457 9767
rect 3433 9718 3485 9764
rect 3541 9718 3593 9764
rect 3649 9718 3701 9764
rect 3757 9718 3809 9764
rect 3865 9718 3917 9764
rect 3973 9718 4025 9764
rect 4081 9718 4133 9764
rect 4189 9718 4241 9764
rect 4297 9718 4349 9764
rect 4405 9718 4457 9764
rect 4513 9718 4565 9764
rect 4621 9718 4673 9764
rect 4729 9718 4781 9764
rect 4837 9718 4889 9764
rect 4945 9718 4997 9764
rect 5053 9718 5105 9764
rect 5161 9718 5213 9764
rect 6566 9718 6618 9764
rect 6674 9718 6726 9764
rect 6782 9718 6834 9764
rect 6890 9718 6942 9764
rect 6998 9718 7050 9764
rect 7106 9718 7158 9764
rect 7214 9718 7266 9764
rect 7322 9718 7374 9764
rect 7430 9718 7482 9764
rect 7538 9718 7590 9764
rect 9677 9718 9729 9764
rect 9785 9718 9837 9764
rect 9893 9718 9945 9764
rect 10001 9718 10053 9764
rect 10109 9718 10161 9764
rect 10217 9718 10269 9764
rect 10325 9718 10377 9764
rect 10433 9718 10485 9764
rect 10541 9718 10593 9764
rect 10649 9718 10701 9764
rect 10757 9718 10809 9764
rect 10865 9718 10917 9764
rect 10973 9718 11025 9764
rect 11081 9718 11133 9764
rect 11189 9718 11241 9764
rect 11297 9718 11349 9764
rect 11405 9718 11457 9764
rect 3433 9715 3485 9718
rect 3541 9715 3593 9718
rect 3649 9715 3701 9718
rect 3757 9715 3809 9718
rect 3865 9715 3917 9718
rect 3973 9715 4025 9718
rect 4081 9715 4133 9718
rect 4189 9715 4241 9718
rect 4297 9715 4349 9718
rect 4405 9715 4457 9718
rect 4513 9715 4565 9718
rect 4621 9715 4673 9718
rect 4729 9715 4781 9718
rect 4837 9715 4889 9718
rect 4945 9715 4997 9718
rect 5053 9715 5105 9718
rect 5161 9715 5213 9718
rect 6566 9715 6618 9718
rect 6674 9715 6726 9718
rect 6782 9715 6834 9718
rect 6890 9715 6942 9718
rect 6998 9715 7050 9718
rect 7106 9715 7158 9718
rect 7214 9715 7266 9718
rect 7322 9715 7374 9718
rect 7430 9715 7482 9718
rect 7538 9715 7590 9718
rect 9677 9715 9729 9718
rect 9785 9715 9837 9718
rect 9893 9715 9945 9718
rect 10001 9715 10053 9718
rect 10109 9715 10161 9718
rect 10217 9715 10269 9718
rect 10325 9715 10377 9718
rect 10433 9715 10485 9718
rect 10541 9715 10593 9718
rect 10649 9715 10701 9718
rect 10757 9715 10809 9718
rect 10865 9715 10917 9718
rect 10973 9715 11025 9718
rect 11081 9715 11133 9718
rect 11189 9715 11241 9718
rect 11297 9715 11349 9718
rect 11405 9715 11457 9718
rect 1505 9520 1557 9523
rect 1613 9520 1665 9523
rect 1721 9520 1773 9523
rect 1829 9520 1881 9523
rect 1937 9520 1989 9523
rect 2045 9520 2097 9523
rect 2153 9520 2205 9523
rect 2261 9520 2313 9523
rect 2369 9520 2421 9523
rect 2477 9520 2529 9523
rect 2585 9520 2637 9523
rect 2693 9520 2745 9523
rect 2801 9520 2853 9523
rect 2909 9520 2961 9523
rect 3017 9520 3069 9523
rect 3125 9520 3177 9523
rect 3233 9520 3285 9523
rect 5372 9520 5424 9523
rect 5480 9520 5532 9523
rect 5588 9520 5640 9523
rect 5696 9520 5748 9523
rect 5804 9520 5856 9523
rect 5912 9520 5964 9523
rect 6020 9520 6072 9523
rect 6128 9520 6180 9523
rect 6236 9520 6288 9523
rect 6344 9520 6396 9523
rect 7749 9520 7801 9523
rect 7857 9520 7909 9523
rect 7965 9520 8017 9523
rect 8073 9520 8125 9523
rect 8181 9520 8233 9523
rect 8289 9520 8341 9523
rect 8397 9520 8449 9523
rect 8505 9520 8557 9523
rect 8613 9520 8665 9523
rect 8721 9520 8773 9523
rect 8829 9520 8881 9523
rect 8937 9520 8989 9523
rect 9045 9520 9097 9523
rect 9153 9520 9205 9523
rect 9261 9520 9313 9523
rect 9369 9520 9421 9523
rect 9477 9520 9529 9523
rect 1505 9474 1557 9520
rect 1613 9474 1665 9520
rect 1721 9474 1773 9520
rect 1829 9474 1881 9520
rect 1937 9474 1989 9520
rect 2045 9474 2097 9520
rect 2153 9474 2205 9520
rect 2261 9474 2313 9520
rect 2369 9474 2421 9520
rect 2477 9474 2529 9520
rect 2585 9474 2637 9520
rect 2693 9474 2745 9520
rect 2801 9474 2853 9520
rect 2909 9474 2961 9520
rect 3017 9474 3069 9520
rect 3125 9474 3177 9520
rect 3233 9474 3285 9520
rect 5372 9474 5424 9520
rect 5480 9474 5532 9520
rect 5588 9474 5640 9520
rect 5696 9474 5748 9520
rect 5804 9474 5856 9520
rect 5912 9474 5964 9520
rect 6020 9474 6072 9520
rect 6128 9474 6180 9520
rect 6236 9474 6288 9520
rect 6344 9474 6396 9520
rect 7749 9474 7801 9520
rect 7857 9474 7909 9520
rect 7965 9474 8017 9520
rect 8073 9474 8125 9520
rect 8181 9474 8233 9520
rect 8289 9474 8341 9520
rect 8397 9474 8449 9520
rect 8505 9474 8557 9520
rect 8613 9474 8665 9520
rect 8721 9474 8773 9520
rect 8829 9474 8881 9520
rect 8937 9474 8989 9520
rect 9045 9474 9097 9520
rect 9153 9474 9205 9520
rect 9261 9474 9313 9520
rect 9369 9474 9421 9520
rect 9477 9474 9529 9520
rect 1505 9471 1557 9474
rect 1613 9471 1665 9474
rect 1721 9471 1773 9474
rect 1829 9471 1881 9474
rect 1937 9471 1989 9474
rect 2045 9471 2097 9474
rect 2153 9471 2205 9474
rect 2261 9471 2313 9474
rect 2369 9471 2421 9474
rect 2477 9471 2529 9474
rect 2585 9471 2637 9474
rect 2693 9471 2745 9474
rect 2801 9471 2853 9474
rect 2909 9471 2961 9474
rect 3017 9471 3069 9474
rect 3125 9471 3177 9474
rect 3233 9471 3285 9474
rect 5372 9471 5424 9474
rect 5480 9471 5532 9474
rect 5588 9471 5640 9474
rect 5696 9471 5748 9474
rect 5804 9471 5856 9474
rect 5912 9471 5964 9474
rect 6020 9471 6072 9474
rect 6128 9471 6180 9474
rect 6236 9471 6288 9474
rect 6344 9471 6396 9474
rect 7749 9471 7801 9474
rect 7857 9471 7909 9474
rect 7965 9471 8017 9474
rect 8073 9471 8125 9474
rect 8181 9471 8233 9474
rect 8289 9471 8341 9474
rect 8397 9471 8449 9474
rect 8505 9471 8557 9474
rect 8613 9471 8665 9474
rect 8721 9471 8773 9474
rect 8829 9471 8881 9474
rect 8937 9471 8989 9474
rect 9045 9471 9097 9474
rect 9153 9471 9205 9474
rect 9261 9471 9313 9474
rect 9369 9471 9421 9474
rect 9477 9471 9529 9474
rect 3433 9276 3485 9279
rect 3541 9276 3593 9279
rect 3649 9276 3701 9279
rect 3757 9276 3809 9279
rect 3865 9276 3917 9279
rect 3973 9276 4025 9279
rect 4081 9276 4133 9279
rect 4189 9276 4241 9279
rect 4297 9276 4349 9279
rect 4405 9276 4457 9279
rect 4513 9276 4565 9279
rect 4621 9276 4673 9279
rect 4729 9276 4781 9279
rect 4837 9276 4889 9279
rect 4945 9276 4997 9279
rect 5053 9276 5105 9279
rect 5161 9276 5213 9279
rect 6566 9276 6618 9279
rect 6674 9276 6726 9279
rect 6782 9276 6834 9279
rect 6890 9276 6942 9279
rect 6998 9276 7050 9279
rect 7106 9276 7158 9279
rect 7214 9276 7266 9279
rect 7322 9276 7374 9279
rect 7430 9276 7482 9279
rect 7538 9276 7590 9279
rect 9677 9276 9729 9279
rect 9785 9276 9837 9279
rect 9893 9276 9945 9279
rect 10001 9276 10053 9279
rect 10109 9276 10161 9279
rect 10217 9276 10269 9279
rect 10325 9276 10377 9279
rect 10433 9276 10485 9279
rect 10541 9276 10593 9279
rect 10649 9276 10701 9279
rect 10757 9276 10809 9279
rect 10865 9276 10917 9279
rect 10973 9276 11025 9279
rect 11081 9276 11133 9279
rect 11189 9276 11241 9279
rect 11297 9276 11349 9279
rect 11405 9276 11457 9279
rect 3433 9230 3485 9276
rect 3541 9230 3593 9276
rect 3649 9230 3701 9276
rect 3757 9230 3809 9276
rect 3865 9230 3917 9276
rect 3973 9230 4025 9276
rect 4081 9230 4133 9276
rect 4189 9230 4241 9276
rect 4297 9230 4349 9276
rect 4405 9230 4457 9276
rect 4513 9230 4565 9276
rect 4621 9230 4673 9276
rect 4729 9230 4781 9276
rect 4837 9230 4889 9276
rect 4945 9230 4997 9276
rect 5053 9230 5105 9276
rect 5161 9230 5213 9276
rect 6566 9230 6618 9276
rect 6674 9230 6726 9276
rect 6782 9230 6834 9276
rect 6890 9230 6942 9276
rect 6998 9230 7050 9276
rect 7106 9230 7158 9276
rect 7214 9230 7266 9276
rect 7322 9230 7374 9276
rect 7430 9230 7482 9276
rect 7538 9230 7590 9276
rect 9677 9230 9729 9276
rect 9785 9230 9837 9276
rect 9893 9230 9945 9276
rect 10001 9230 10053 9276
rect 10109 9230 10161 9276
rect 10217 9230 10269 9276
rect 10325 9230 10377 9276
rect 10433 9230 10485 9276
rect 10541 9230 10593 9276
rect 10649 9230 10701 9276
rect 10757 9230 10809 9276
rect 10865 9230 10917 9276
rect 10973 9230 11025 9276
rect 11081 9230 11133 9276
rect 11189 9230 11241 9276
rect 11297 9230 11349 9276
rect 11405 9230 11457 9276
rect 3433 9227 3485 9230
rect 3541 9227 3593 9230
rect 3649 9227 3701 9230
rect 3757 9227 3809 9230
rect 3865 9227 3917 9230
rect 3973 9227 4025 9230
rect 4081 9227 4133 9230
rect 4189 9227 4241 9230
rect 4297 9227 4349 9230
rect 4405 9227 4457 9230
rect 4513 9227 4565 9230
rect 4621 9227 4673 9230
rect 4729 9227 4781 9230
rect 4837 9227 4889 9230
rect 4945 9227 4997 9230
rect 5053 9227 5105 9230
rect 5161 9227 5213 9230
rect 6566 9227 6618 9230
rect 6674 9227 6726 9230
rect 6782 9227 6834 9230
rect 6890 9227 6942 9230
rect 6998 9227 7050 9230
rect 7106 9227 7158 9230
rect 7214 9227 7266 9230
rect 7322 9227 7374 9230
rect 7430 9227 7482 9230
rect 7538 9227 7590 9230
rect 9677 9227 9729 9230
rect 9785 9227 9837 9230
rect 9893 9227 9945 9230
rect 10001 9227 10053 9230
rect 10109 9227 10161 9230
rect 10217 9227 10269 9230
rect 10325 9227 10377 9230
rect 10433 9227 10485 9230
rect 10541 9227 10593 9230
rect 10649 9227 10701 9230
rect 10757 9227 10809 9230
rect 10865 9227 10917 9230
rect 10973 9227 11025 9230
rect 11081 9227 11133 9230
rect 11189 9227 11241 9230
rect 11297 9227 11349 9230
rect 11405 9227 11457 9230
rect 1505 9032 1557 9035
rect 1613 9032 1665 9035
rect 1721 9032 1773 9035
rect 1829 9032 1881 9035
rect 1937 9032 1989 9035
rect 2045 9032 2097 9035
rect 2153 9032 2205 9035
rect 2261 9032 2313 9035
rect 2369 9032 2421 9035
rect 2477 9032 2529 9035
rect 2585 9032 2637 9035
rect 2693 9032 2745 9035
rect 2801 9032 2853 9035
rect 2909 9032 2961 9035
rect 3017 9032 3069 9035
rect 3125 9032 3177 9035
rect 3233 9032 3285 9035
rect 5372 9032 5424 9035
rect 5480 9032 5532 9035
rect 5588 9032 5640 9035
rect 5696 9032 5748 9035
rect 5804 9032 5856 9035
rect 5912 9032 5964 9035
rect 6020 9032 6072 9035
rect 6128 9032 6180 9035
rect 6236 9032 6288 9035
rect 6344 9032 6396 9035
rect 7749 9032 7801 9035
rect 7857 9032 7909 9035
rect 7965 9032 8017 9035
rect 8073 9032 8125 9035
rect 8181 9032 8233 9035
rect 8289 9032 8341 9035
rect 8397 9032 8449 9035
rect 8505 9032 8557 9035
rect 8613 9032 8665 9035
rect 8721 9032 8773 9035
rect 8829 9032 8881 9035
rect 8937 9032 8989 9035
rect 9045 9032 9097 9035
rect 9153 9032 9205 9035
rect 9261 9032 9313 9035
rect 9369 9032 9421 9035
rect 9477 9032 9529 9035
rect 1505 8986 1557 9032
rect 1613 8986 1665 9032
rect 1721 8986 1773 9032
rect 1829 8986 1881 9032
rect 1937 8986 1989 9032
rect 2045 8986 2097 9032
rect 2153 8986 2205 9032
rect 2261 8986 2313 9032
rect 2369 8986 2421 9032
rect 2477 8986 2529 9032
rect 2585 8986 2637 9032
rect 2693 8986 2745 9032
rect 2801 8986 2853 9032
rect 2909 8986 2961 9032
rect 3017 8986 3069 9032
rect 3125 8986 3177 9032
rect 3233 8986 3285 9032
rect 5372 8986 5424 9032
rect 5480 8986 5532 9032
rect 5588 8986 5640 9032
rect 5696 8986 5748 9032
rect 5804 8986 5856 9032
rect 5912 8986 5964 9032
rect 6020 8986 6072 9032
rect 6128 8986 6180 9032
rect 6236 8986 6288 9032
rect 6344 8986 6396 9032
rect 7749 8986 7801 9032
rect 7857 8986 7909 9032
rect 7965 8986 8017 9032
rect 8073 8986 8125 9032
rect 8181 8986 8233 9032
rect 8289 8986 8341 9032
rect 8397 8986 8449 9032
rect 8505 8986 8557 9032
rect 8613 8986 8665 9032
rect 8721 8986 8773 9032
rect 8829 8986 8881 9032
rect 8937 8986 8989 9032
rect 9045 8986 9097 9032
rect 9153 8986 9205 9032
rect 9261 8986 9313 9032
rect 9369 8986 9421 9032
rect 9477 8986 9529 9032
rect 1505 8983 1557 8986
rect 1613 8983 1665 8986
rect 1721 8983 1773 8986
rect 1829 8983 1881 8986
rect 1937 8983 1989 8986
rect 2045 8983 2097 8986
rect 2153 8983 2205 8986
rect 2261 8983 2313 8986
rect 2369 8983 2421 8986
rect 2477 8983 2529 8986
rect 2585 8983 2637 8986
rect 2693 8983 2745 8986
rect 2801 8983 2853 8986
rect 2909 8983 2961 8986
rect 3017 8983 3069 8986
rect 3125 8983 3177 8986
rect 3233 8983 3285 8986
rect 5372 8983 5424 8986
rect 5480 8983 5532 8986
rect 5588 8983 5640 8986
rect 5696 8983 5748 8986
rect 5804 8983 5856 8986
rect 5912 8983 5964 8986
rect 6020 8983 6072 8986
rect 6128 8983 6180 8986
rect 6236 8983 6288 8986
rect 6344 8983 6396 8986
rect 7749 8983 7801 8986
rect 7857 8983 7909 8986
rect 7965 8983 8017 8986
rect 8073 8983 8125 8986
rect 8181 8983 8233 8986
rect 8289 8983 8341 8986
rect 8397 8983 8449 8986
rect 8505 8983 8557 8986
rect 8613 8983 8665 8986
rect 8721 8983 8773 8986
rect 8829 8983 8881 8986
rect 8937 8983 8989 8986
rect 9045 8983 9097 8986
rect 9153 8983 9205 8986
rect 9261 8983 9313 8986
rect 9369 8983 9421 8986
rect 9477 8983 9529 8986
rect 3433 8788 3485 8791
rect 3541 8788 3593 8791
rect 3649 8788 3701 8791
rect 3757 8788 3809 8791
rect 3865 8788 3917 8791
rect 3973 8788 4025 8791
rect 4081 8788 4133 8791
rect 4189 8788 4241 8791
rect 4297 8788 4349 8791
rect 4405 8788 4457 8791
rect 4513 8788 4565 8791
rect 4621 8788 4673 8791
rect 4729 8788 4781 8791
rect 4837 8788 4889 8791
rect 4945 8788 4997 8791
rect 5053 8788 5105 8791
rect 5161 8788 5213 8791
rect 6566 8788 6618 8791
rect 6674 8788 6726 8791
rect 6782 8788 6834 8791
rect 6890 8788 6942 8791
rect 6998 8788 7050 8791
rect 7106 8788 7158 8791
rect 7214 8788 7266 8791
rect 7322 8788 7374 8791
rect 7430 8788 7482 8791
rect 7538 8788 7590 8791
rect 9677 8788 9729 8791
rect 9785 8788 9837 8791
rect 9893 8788 9945 8791
rect 10001 8788 10053 8791
rect 10109 8788 10161 8791
rect 10217 8788 10269 8791
rect 10325 8788 10377 8791
rect 10433 8788 10485 8791
rect 10541 8788 10593 8791
rect 10649 8788 10701 8791
rect 10757 8788 10809 8791
rect 10865 8788 10917 8791
rect 10973 8788 11025 8791
rect 11081 8788 11133 8791
rect 11189 8788 11241 8791
rect 11297 8788 11349 8791
rect 11405 8788 11457 8791
rect 3433 8742 3485 8788
rect 3541 8742 3593 8788
rect 3649 8742 3701 8788
rect 3757 8742 3809 8788
rect 3865 8742 3917 8788
rect 3973 8742 4025 8788
rect 4081 8742 4133 8788
rect 4189 8742 4241 8788
rect 4297 8742 4349 8788
rect 4405 8742 4457 8788
rect 4513 8742 4565 8788
rect 4621 8742 4673 8788
rect 4729 8742 4781 8788
rect 4837 8742 4889 8788
rect 4945 8742 4997 8788
rect 5053 8742 5105 8788
rect 5161 8742 5213 8788
rect 6566 8742 6618 8788
rect 6674 8742 6726 8788
rect 6782 8742 6834 8788
rect 6890 8742 6942 8788
rect 6998 8742 7050 8788
rect 7106 8742 7158 8788
rect 7214 8742 7266 8788
rect 7322 8742 7374 8788
rect 7430 8742 7482 8788
rect 7538 8742 7590 8788
rect 9677 8742 9729 8788
rect 9785 8742 9837 8788
rect 9893 8742 9945 8788
rect 10001 8742 10053 8788
rect 10109 8742 10161 8788
rect 10217 8742 10269 8788
rect 10325 8742 10377 8788
rect 10433 8742 10485 8788
rect 10541 8742 10593 8788
rect 10649 8742 10701 8788
rect 10757 8742 10809 8788
rect 10865 8742 10917 8788
rect 10973 8742 11025 8788
rect 11081 8742 11133 8788
rect 11189 8742 11241 8788
rect 11297 8742 11349 8788
rect 11405 8742 11457 8788
rect 3433 8739 3485 8742
rect 3541 8739 3593 8742
rect 3649 8739 3701 8742
rect 3757 8739 3809 8742
rect 3865 8739 3917 8742
rect 3973 8739 4025 8742
rect 4081 8739 4133 8742
rect 4189 8739 4241 8742
rect 4297 8739 4349 8742
rect 4405 8739 4457 8742
rect 4513 8739 4565 8742
rect 4621 8739 4673 8742
rect 4729 8739 4781 8742
rect 4837 8739 4889 8742
rect 4945 8739 4997 8742
rect 5053 8739 5105 8742
rect 5161 8739 5213 8742
rect 6566 8739 6618 8742
rect 6674 8739 6726 8742
rect 6782 8739 6834 8742
rect 6890 8739 6942 8742
rect 6998 8739 7050 8742
rect 7106 8739 7158 8742
rect 7214 8739 7266 8742
rect 7322 8739 7374 8742
rect 7430 8739 7482 8742
rect 7538 8739 7590 8742
rect 9677 8739 9729 8742
rect 9785 8739 9837 8742
rect 9893 8739 9945 8742
rect 10001 8739 10053 8742
rect 10109 8739 10161 8742
rect 10217 8739 10269 8742
rect 10325 8739 10377 8742
rect 10433 8739 10485 8742
rect 10541 8739 10593 8742
rect 10649 8739 10701 8742
rect 10757 8739 10809 8742
rect 10865 8739 10917 8742
rect 10973 8739 11025 8742
rect 11081 8739 11133 8742
rect 11189 8739 11241 8742
rect 11297 8739 11349 8742
rect 11405 8739 11457 8742
rect 1505 8544 1557 8547
rect 1613 8544 1665 8547
rect 1721 8544 1773 8547
rect 1829 8544 1881 8547
rect 1937 8544 1989 8547
rect 2045 8544 2097 8547
rect 2153 8544 2205 8547
rect 2261 8544 2313 8547
rect 2369 8544 2421 8547
rect 2477 8544 2529 8547
rect 2585 8544 2637 8547
rect 2693 8544 2745 8547
rect 2801 8544 2853 8547
rect 2909 8544 2961 8547
rect 3017 8544 3069 8547
rect 3125 8544 3177 8547
rect 3233 8544 3285 8547
rect 5372 8544 5424 8547
rect 5480 8544 5532 8547
rect 5588 8544 5640 8547
rect 5696 8544 5748 8547
rect 5804 8544 5856 8547
rect 5912 8544 5964 8547
rect 6020 8544 6072 8547
rect 6128 8544 6180 8547
rect 6236 8544 6288 8547
rect 6344 8544 6396 8547
rect 7749 8544 7801 8547
rect 7857 8544 7909 8547
rect 7965 8544 8017 8547
rect 8073 8544 8125 8547
rect 8181 8544 8233 8547
rect 8289 8544 8341 8547
rect 8397 8544 8449 8547
rect 8505 8544 8557 8547
rect 8613 8544 8665 8547
rect 8721 8544 8773 8547
rect 8829 8544 8881 8547
rect 8937 8544 8989 8547
rect 9045 8544 9097 8547
rect 9153 8544 9205 8547
rect 9261 8544 9313 8547
rect 9369 8544 9421 8547
rect 9477 8544 9529 8547
rect 1505 8498 1557 8544
rect 1613 8498 1665 8544
rect 1721 8498 1773 8544
rect 1829 8498 1881 8544
rect 1937 8498 1989 8544
rect 2045 8498 2097 8544
rect 2153 8498 2205 8544
rect 2261 8498 2313 8544
rect 2369 8498 2421 8544
rect 2477 8498 2529 8544
rect 2585 8498 2637 8544
rect 2693 8498 2745 8544
rect 2801 8498 2853 8544
rect 2909 8498 2961 8544
rect 3017 8498 3069 8544
rect 3125 8498 3177 8544
rect 3233 8498 3285 8544
rect 5372 8498 5424 8544
rect 5480 8498 5532 8544
rect 5588 8498 5640 8544
rect 5696 8498 5748 8544
rect 5804 8498 5856 8544
rect 5912 8498 5964 8544
rect 6020 8498 6072 8544
rect 6128 8498 6180 8544
rect 6236 8498 6288 8544
rect 6344 8498 6396 8544
rect 7749 8498 7801 8544
rect 7857 8498 7909 8544
rect 7965 8498 8017 8544
rect 8073 8498 8125 8544
rect 8181 8498 8233 8544
rect 8289 8498 8341 8544
rect 8397 8498 8449 8544
rect 8505 8498 8557 8544
rect 8613 8498 8665 8544
rect 8721 8498 8773 8544
rect 8829 8498 8881 8544
rect 8937 8498 8989 8544
rect 9045 8498 9097 8544
rect 9153 8498 9205 8544
rect 9261 8498 9313 8544
rect 9369 8498 9421 8544
rect 9477 8498 9529 8544
rect 1505 8495 1557 8498
rect 1613 8495 1665 8498
rect 1721 8495 1773 8498
rect 1829 8495 1881 8498
rect 1937 8495 1989 8498
rect 2045 8495 2097 8498
rect 2153 8495 2205 8498
rect 2261 8495 2313 8498
rect 2369 8495 2421 8498
rect 2477 8495 2529 8498
rect 2585 8495 2637 8498
rect 2693 8495 2745 8498
rect 2801 8495 2853 8498
rect 2909 8495 2961 8498
rect 3017 8495 3069 8498
rect 3125 8495 3177 8498
rect 3233 8495 3285 8498
rect 5372 8495 5424 8498
rect 5480 8495 5532 8498
rect 5588 8495 5640 8498
rect 5696 8495 5748 8498
rect 5804 8495 5856 8498
rect 5912 8495 5964 8498
rect 6020 8495 6072 8498
rect 6128 8495 6180 8498
rect 6236 8495 6288 8498
rect 6344 8495 6396 8498
rect 7749 8495 7801 8498
rect 7857 8495 7909 8498
rect 7965 8495 8017 8498
rect 8073 8495 8125 8498
rect 8181 8495 8233 8498
rect 8289 8495 8341 8498
rect 8397 8495 8449 8498
rect 8505 8495 8557 8498
rect 8613 8495 8665 8498
rect 8721 8495 8773 8498
rect 8829 8495 8881 8498
rect 8937 8495 8989 8498
rect 9045 8495 9097 8498
rect 9153 8495 9205 8498
rect 9261 8495 9313 8498
rect 9369 8495 9421 8498
rect 9477 8495 9529 8498
rect 3433 8300 3485 8303
rect 3541 8300 3593 8303
rect 3649 8300 3701 8303
rect 3757 8300 3809 8303
rect 3865 8300 3917 8303
rect 3973 8300 4025 8303
rect 4081 8300 4133 8303
rect 4189 8300 4241 8303
rect 4297 8300 4349 8303
rect 4405 8300 4457 8303
rect 4513 8300 4565 8303
rect 4621 8300 4673 8303
rect 4729 8300 4781 8303
rect 4837 8300 4889 8303
rect 4945 8300 4997 8303
rect 5053 8300 5105 8303
rect 5161 8300 5213 8303
rect 6566 8300 6618 8303
rect 6674 8300 6726 8303
rect 6782 8300 6834 8303
rect 6890 8300 6942 8303
rect 6998 8300 7050 8303
rect 7106 8300 7158 8303
rect 7214 8300 7266 8303
rect 7322 8300 7374 8303
rect 7430 8300 7482 8303
rect 7538 8300 7590 8303
rect 9677 8300 9729 8303
rect 9785 8300 9837 8303
rect 9893 8300 9945 8303
rect 10001 8300 10053 8303
rect 10109 8300 10161 8303
rect 10217 8300 10269 8303
rect 10325 8300 10377 8303
rect 10433 8300 10485 8303
rect 10541 8300 10593 8303
rect 10649 8300 10701 8303
rect 10757 8300 10809 8303
rect 10865 8300 10917 8303
rect 10973 8300 11025 8303
rect 11081 8300 11133 8303
rect 11189 8300 11241 8303
rect 11297 8300 11349 8303
rect 11405 8300 11457 8303
rect 3433 8254 3485 8300
rect 3541 8254 3593 8300
rect 3649 8254 3701 8300
rect 3757 8254 3809 8300
rect 3865 8254 3917 8300
rect 3973 8254 4025 8300
rect 4081 8254 4133 8300
rect 4189 8254 4241 8300
rect 4297 8254 4349 8300
rect 4405 8254 4457 8300
rect 4513 8254 4565 8300
rect 4621 8254 4673 8300
rect 4729 8254 4781 8300
rect 4837 8254 4889 8300
rect 4945 8254 4997 8300
rect 5053 8254 5105 8300
rect 5161 8254 5213 8300
rect 6566 8254 6618 8300
rect 6674 8254 6726 8300
rect 6782 8254 6834 8300
rect 6890 8254 6942 8300
rect 6998 8254 7050 8300
rect 7106 8254 7158 8300
rect 7214 8254 7266 8300
rect 7322 8254 7374 8300
rect 7430 8254 7482 8300
rect 7538 8254 7590 8300
rect 9677 8254 9729 8300
rect 9785 8254 9837 8300
rect 9893 8254 9945 8300
rect 10001 8254 10053 8300
rect 10109 8254 10161 8300
rect 10217 8254 10269 8300
rect 10325 8254 10377 8300
rect 10433 8254 10485 8300
rect 10541 8254 10593 8300
rect 10649 8254 10701 8300
rect 10757 8254 10809 8300
rect 10865 8254 10917 8300
rect 10973 8254 11025 8300
rect 11081 8254 11133 8300
rect 11189 8254 11241 8300
rect 11297 8254 11349 8300
rect 11405 8254 11457 8300
rect 3433 8251 3485 8254
rect 3541 8251 3593 8254
rect 3649 8251 3701 8254
rect 3757 8251 3809 8254
rect 3865 8251 3917 8254
rect 3973 8251 4025 8254
rect 4081 8251 4133 8254
rect 4189 8251 4241 8254
rect 4297 8251 4349 8254
rect 4405 8251 4457 8254
rect 4513 8251 4565 8254
rect 4621 8251 4673 8254
rect 4729 8251 4781 8254
rect 4837 8251 4889 8254
rect 4945 8251 4997 8254
rect 5053 8251 5105 8254
rect 5161 8251 5213 8254
rect 6566 8251 6618 8254
rect 6674 8251 6726 8254
rect 6782 8251 6834 8254
rect 6890 8251 6942 8254
rect 6998 8251 7050 8254
rect 7106 8251 7158 8254
rect 7214 8251 7266 8254
rect 7322 8251 7374 8254
rect 7430 8251 7482 8254
rect 7538 8251 7590 8254
rect 9677 8251 9729 8254
rect 9785 8251 9837 8254
rect 9893 8251 9945 8254
rect 10001 8251 10053 8254
rect 10109 8251 10161 8254
rect 10217 8251 10269 8254
rect 10325 8251 10377 8254
rect 10433 8251 10485 8254
rect 10541 8251 10593 8254
rect 10649 8251 10701 8254
rect 10757 8251 10809 8254
rect 10865 8251 10917 8254
rect 10973 8251 11025 8254
rect 11081 8251 11133 8254
rect 11189 8251 11241 8254
rect 11297 8251 11349 8254
rect 11405 8251 11457 8254
rect 1505 8056 1557 8059
rect 1613 8056 1665 8059
rect 1721 8056 1773 8059
rect 1829 8056 1881 8059
rect 1937 8056 1989 8059
rect 2045 8056 2097 8059
rect 2153 8056 2205 8059
rect 2261 8056 2313 8059
rect 2369 8056 2421 8059
rect 2477 8056 2529 8059
rect 2585 8056 2637 8059
rect 2693 8056 2745 8059
rect 2801 8056 2853 8059
rect 2909 8056 2961 8059
rect 3017 8056 3069 8059
rect 3125 8056 3177 8059
rect 3233 8056 3285 8059
rect 5372 8056 5424 8059
rect 5480 8056 5532 8059
rect 5588 8056 5640 8059
rect 5696 8056 5748 8059
rect 5804 8056 5856 8059
rect 5912 8056 5964 8059
rect 6020 8056 6072 8059
rect 6128 8056 6180 8059
rect 6236 8056 6288 8059
rect 6344 8056 6396 8059
rect 7749 8056 7801 8059
rect 7857 8056 7909 8059
rect 7965 8056 8017 8059
rect 8073 8056 8125 8059
rect 8181 8056 8233 8059
rect 8289 8056 8341 8059
rect 8397 8056 8449 8059
rect 8505 8056 8557 8059
rect 8613 8056 8665 8059
rect 8721 8056 8773 8059
rect 8829 8056 8881 8059
rect 8937 8056 8989 8059
rect 9045 8056 9097 8059
rect 9153 8056 9205 8059
rect 9261 8056 9313 8059
rect 9369 8056 9421 8059
rect 9477 8056 9529 8059
rect 1505 8010 1557 8056
rect 1613 8010 1665 8056
rect 1721 8010 1773 8056
rect 1829 8010 1881 8056
rect 1937 8010 1989 8056
rect 2045 8010 2097 8056
rect 2153 8010 2205 8056
rect 2261 8010 2313 8056
rect 2369 8010 2421 8056
rect 2477 8010 2529 8056
rect 2585 8010 2637 8056
rect 2693 8010 2745 8056
rect 2801 8010 2853 8056
rect 2909 8010 2961 8056
rect 3017 8010 3069 8056
rect 3125 8010 3177 8056
rect 3233 8010 3285 8056
rect 5372 8010 5424 8056
rect 5480 8010 5532 8056
rect 5588 8010 5640 8056
rect 5696 8010 5748 8056
rect 5804 8010 5856 8056
rect 5912 8010 5964 8056
rect 6020 8010 6072 8056
rect 6128 8010 6180 8056
rect 6236 8010 6288 8056
rect 6344 8010 6396 8056
rect 7749 8010 7801 8056
rect 7857 8010 7909 8056
rect 7965 8010 8017 8056
rect 8073 8010 8125 8056
rect 8181 8010 8233 8056
rect 8289 8010 8341 8056
rect 8397 8010 8449 8056
rect 8505 8010 8557 8056
rect 8613 8010 8665 8056
rect 8721 8010 8773 8056
rect 8829 8010 8881 8056
rect 8937 8010 8989 8056
rect 9045 8010 9097 8056
rect 9153 8010 9205 8056
rect 9261 8010 9313 8056
rect 9369 8010 9421 8056
rect 9477 8010 9529 8056
rect 1505 8007 1557 8010
rect 1613 8007 1665 8010
rect 1721 8007 1773 8010
rect 1829 8007 1881 8010
rect 1937 8007 1989 8010
rect 2045 8007 2097 8010
rect 2153 8007 2205 8010
rect 2261 8007 2313 8010
rect 2369 8007 2421 8010
rect 2477 8007 2529 8010
rect 2585 8007 2637 8010
rect 2693 8007 2745 8010
rect 2801 8007 2853 8010
rect 2909 8007 2961 8010
rect 3017 8007 3069 8010
rect 3125 8007 3177 8010
rect 3233 8007 3285 8010
rect 5372 8007 5424 8010
rect 5480 8007 5532 8010
rect 5588 8007 5640 8010
rect 5696 8007 5748 8010
rect 5804 8007 5856 8010
rect 5912 8007 5964 8010
rect 6020 8007 6072 8010
rect 6128 8007 6180 8010
rect 6236 8007 6288 8010
rect 6344 8007 6396 8010
rect 7749 8007 7801 8010
rect 7857 8007 7909 8010
rect 7965 8007 8017 8010
rect 8073 8007 8125 8010
rect 8181 8007 8233 8010
rect 8289 8007 8341 8010
rect 8397 8007 8449 8010
rect 8505 8007 8557 8010
rect 8613 8007 8665 8010
rect 8721 8007 8773 8010
rect 8829 8007 8881 8010
rect 8937 8007 8989 8010
rect 9045 8007 9097 8010
rect 9153 8007 9205 8010
rect 9261 8007 9313 8010
rect 9369 8007 9421 8010
rect 9477 8007 9529 8010
rect 3433 7812 3485 7815
rect 3541 7812 3593 7815
rect 3649 7812 3701 7815
rect 3757 7812 3809 7815
rect 3865 7812 3917 7815
rect 3973 7812 4025 7815
rect 4081 7812 4133 7815
rect 4189 7812 4241 7815
rect 4297 7812 4349 7815
rect 4405 7812 4457 7815
rect 4513 7812 4565 7815
rect 4621 7812 4673 7815
rect 4729 7812 4781 7815
rect 4837 7812 4889 7815
rect 4945 7812 4997 7815
rect 5053 7812 5105 7815
rect 5161 7812 5213 7815
rect 6566 7812 6618 7815
rect 6674 7812 6726 7815
rect 6782 7812 6834 7815
rect 6890 7812 6942 7815
rect 6998 7812 7050 7815
rect 7106 7812 7158 7815
rect 7214 7812 7266 7815
rect 7322 7812 7374 7815
rect 7430 7812 7482 7815
rect 7538 7812 7590 7815
rect 9677 7812 9729 7815
rect 9785 7812 9837 7815
rect 9893 7812 9945 7815
rect 10001 7812 10053 7815
rect 10109 7812 10161 7815
rect 10217 7812 10269 7815
rect 10325 7812 10377 7815
rect 10433 7812 10485 7815
rect 10541 7812 10593 7815
rect 10649 7812 10701 7815
rect 10757 7812 10809 7815
rect 10865 7812 10917 7815
rect 10973 7812 11025 7815
rect 11081 7812 11133 7815
rect 11189 7812 11241 7815
rect 11297 7812 11349 7815
rect 11405 7812 11457 7815
rect 3433 7766 3485 7812
rect 3541 7766 3593 7812
rect 3649 7766 3701 7812
rect 3757 7766 3809 7812
rect 3865 7766 3917 7812
rect 3973 7766 4025 7812
rect 4081 7766 4133 7812
rect 4189 7766 4241 7812
rect 4297 7766 4349 7812
rect 4405 7766 4457 7812
rect 4513 7766 4565 7812
rect 4621 7766 4673 7812
rect 4729 7766 4781 7812
rect 4837 7766 4889 7812
rect 4945 7766 4997 7812
rect 5053 7766 5105 7812
rect 5161 7766 5213 7812
rect 6566 7766 6618 7812
rect 6674 7766 6726 7812
rect 6782 7766 6834 7812
rect 6890 7766 6942 7812
rect 6998 7766 7050 7812
rect 7106 7766 7158 7812
rect 7214 7766 7266 7812
rect 7322 7766 7374 7812
rect 7430 7766 7482 7812
rect 7538 7766 7590 7812
rect 9677 7766 9729 7812
rect 9785 7766 9837 7812
rect 9893 7766 9945 7812
rect 10001 7766 10053 7812
rect 10109 7766 10161 7812
rect 10217 7766 10269 7812
rect 10325 7766 10377 7812
rect 10433 7766 10485 7812
rect 10541 7766 10593 7812
rect 10649 7766 10701 7812
rect 10757 7766 10809 7812
rect 10865 7766 10917 7812
rect 10973 7766 11025 7812
rect 11081 7766 11133 7812
rect 11189 7766 11241 7812
rect 11297 7766 11349 7812
rect 11405 7766 11457 7812
rect 3433 7763 3485 7766
rect 3541 7763 3593 7766
rect 3649 7763 3701 7766
rect 3757 7763 3809 7766
rect 3865 7763 3917 7766
rect 3973 7763 4025 7766
rect 4081 7763 4133 7766
rect 4189 7763 4241 7766
rect 4297 7763 4349 7766
rect 4405 7763 4457 7766
rect 4513 7763 4565 7766
rect 4621 7763 4673 7766
rect 4729 7763 4781 7766
rect 4837 7763 4889 7766
rect 4945 7763 4997 7766
rect 5053 7763 5105 7766
rect 5161 7763 5213 7766
rect 6566 7763 6618 7766
rect 6674 7763 6726 7766
rect 6782 7763 6834 7766
rect 6890 7763 6942 7766
rect 6998 7763 7050 7766
rect 7106 7763 7158 7766
rect 7214 7763 7266 7766
rect 7322 7763 7374 7766
rect 7430 7763 7482 7766
rect 7538 7763 7590 7766
rect 9677 7763 9729 7766
rect 9785 7763 9837 7766
rect 9893 7763 9945 7766
rect 10001 7763 10053 7766
rect 10109 7763 10161 7766
rect 10217 7763 10269 7766
rect 10325 7763 10377 7766
rect 10433 7763 10485 7766
rect 10541 7763 10593 7766
rect 10649 7763 10701 7766
rect 10757 7763 10809 7766
rect 10865 7763 10917 7766
rect 10973 7763 11025 7766
rect 11081 7763 11133 7766
rect 11189 7763 11241 7766
rect 11297 7763 11349 7766
rect 11405 7763 11457 7766
rect 1505 7568 1557 7571
rect 1613 7568 1665 7571
rect 1721 7568 1773 7571
rect 1829 7568 1881 7571
rect 1937 7568 1989 7571
rect 2045 7568 2097 7571
rect 2153 7568 2205 7571
rect 2261 7568 2313 7571
rect 2369 7568 2421 7571
rect 2477 7568 2529 7571
rect 2585 7568 2637 7571
rect 2693 7568 2745 7571
rect 2801 7568 2853 7571
rect 2909 7568 2961 7571
rect 3017 7568 3069 7571
rect 3125 7568 3177 7571
rect 3233 7568 3285 7571
rect 5372 7568 5424 7571
rect 5480 7568 5532 7571
rect 5588 7568 5640 7571
rect 5696 7568 5748 7571
rect 5804 7568 5856 7571
rect 5912 7568 5964 7571
rect 6020 7568 6072 7571
rect 6128 7568 6180 7571
rect 6236 7568 6288 7571
rect 6344 7568 6396 7571
rect 7749 7568 7801 7571
rect 7857 7568 7909 7571
rect 7965 7568 8017 7571
rect 8073 7568 8125 7571
rect 8181 7568 8233 7571
rect 8289 7568 8341 7571
rect 8397 7568 8449 7571
rect 8505 7568 8557 7571
rect 8613 7568 8665 7571
rect 8721 7568 8773 7571
rect 8829 7568 8881 7571
rect 8937 7568 8989 7571
rect 9045 7568 9097 7571
rect 9153 7568 9205 7571
rect 9261 7568 9313 7571
rect 9369 7568 9421 7571
rect 9477 7568 9529 7571
rect 1505 7522 1557 7568
rect 1613 7522 1665 7568
rect 1721 7522 1773 7568
rect 1829 7522 1881 7568
rect 1937 7522 1989 7568
rect 2045 7522 2097 7568
rect 2153 7522 2205 7568
rect 2261 7522 2313 7568
rect 2369 7522 2421 7568
rect 2477 7522 2529 7568
rect 2585 7522 2637 7568
rect 2693 7522 2745 7568
rect 2801 7522 2853 7568
rect 2909 7522 2961 7568
rect 3017 7522 3069 7568
rect 3125 7522 3177 7568
rect 3233 7522 3285 7568
rect 5372 7522 5424 7568
rect 5480 7522 5532 7568
rect 5588 7522 5640 7568
rect 5696 7522 5748 7568
rect 5804 7522 5856 7568
rect 5912 7522 5964 7568
rect 6020 7522 6072 7568
rect 6128 7522 6180 7568
rect 6236 7522 6288 7568
rect 6344 7522 6396 7568
rect 7749 7522 7801 7568
rect 7857 7522 7909 7568
rect 7965 7522 8017 7568
rect 8073 7522 8125 7568
rect 8181 7522 8233 7568
rect 8289 7522 8341 7568
rect 8397 7522 8449 7568
rect 8505 7522 8557 7568
rect 8613 7522 8665 7568
rect 8721 7522 8773 7568
rect 8829 7522 8881 7568
rect 8937 7522 8989 7568
rect 9045 7522 9097 7568
rect 9153 7522 9205 7568
rect 9261 7522 9313 7568
rect 9369 7522 9421 7568
rect 9477 7522 9529 7568
rect 1505 7519 1557 7522
rect 1613 7519 1665 7522
rect 1721 7519 1773 7522
rect 1829 7519 1881 7522
rect 1937 7519 1989 7522
rect 2045 7519 2097 7522
rect 2153 7519 2205 7522
rect 2261 7519 2313 7522
rect 2369 7519 2421 7522
rect 2477 7519 2529 7522
rect 2585 7519 2637 7522
rect 2693 7519 2745 7522
rect 2801 7519 2853 7522
rect 2909 7519 2961 7522
rect 3017 7519 3069 7522
rect 3125 7519 3177 7522
rect 3233 7519 3285 7522
rect 5372 7519 5424 7522
rect 5480 7519 5532 7522
rect 5588 7519 5640 7522
rect 5696 7519 5748 7522
rect 5804 7519 5856 7522
rect 5912 7519 5964 7522
rect 6020 7519 6072 7522
rect 6128 7519 6180 7522
rect 6236 7519 6288 7522
rect 6344 7519 6396 7522
rect 7749 7519 7801 7522
rect 7857 7519 7909 7522
rect 7965 7519 8017 7522
rect 8073 7519 8125 7522
rect 8181 7519 8233 7522
rect 8289 7519 8341 7522
rect 8397 7519 8449 7522
rect 8505 7519 8557 7522
rect 8613 7519 8665 7522
rect 8721 7519 8773 7522
rect 8829 7519 8881 7522
rect 8937 7519 8989 7522
rect 9045 7519 9097 7522
rect 9153 7519 9205 7522
rect 9261 7519 9313 7522
rect 9369 7519 9421 7522
rect 9477 7519 9529 7522
rect 1233 7339 1285 7391
rect 1341 7339 1393 7391
rect 11569 11983 11621 12035
rect 11677 11983 11706 12035
rect 11706 11983 11729 12035
rect 11569 11875 11621 11927
rect 11677 11875 11706 11927
rect 11706 11875 11729 11927
rect 11569 11767 11621 11819
rect 11677 11767 11706 11819
rect 11706 11767 11729 11819
rect 11569 11659 11621 11711
rect 11677 11659 11706 11711
rect 11706 11659 11729 11711
rect 11569 11551 11621 11603
rect 11677 11551 11706 11603
rect 11706 11551 11729 11603
rect 11569 11443 11621 11495
rect 11677 11443 11706 11495
rect 11706 11443 11729 11495
rect 11569 11335 11621 11387
rect 11677 11335 11706 11387
rect 11706 11335 11729 11387
rect 11569 11227 11621 11279
rect 11677 11227 11706 11279
rect 11706 11227 11729 11279
rect 11569 11119 11621 11171
rect 11677 11119 11706 11171
rect 11706 11119 11729 11171
rect 11569 11011 11621 11063
rect 11677 11011 11706 11063
rect 11706 11011 11729 11063
rect 11569 10903 11621 10955
rect 11677 10903 11706 10955
rect 11706 10903 11729 10955
rect 11569 10795 11621 10847
rect 11677 10795 11706 10847
rect 11706 10795 11729 10847
rect 11569 10687 11621 10739
rect 11677 10687 11706 10739
rect 11706 10687 11729 10739
rect 11569 10579 11621 10631
rect 11677 10579 11706 10631
rect 11706 10579 11729 10631
rect 11569 10471 11621 10523
rect 11677 10471 11706 10523
rect 11706 10471 11729 10523
rect 11569 10363 11621 10415
rect 11677 10363 11706 10415
rect 11706 10363 11729 10415
rect 11569 10255 11621 10307
rect 11677 10255 11706 10307
rect 11706 10255 11729 10307
rect 11569 10147 11621 10199
rect 11677 10147 11706 10199
rect 11706 10147 11729 10199
rect 11569 10039 11621 10091
rect 11677 10039 11706 10091
rect 11706 10039 11729 10091
rect 11569 9931 11621 9983
rect 11677 9931 11706 9983
rect 11706 9931 11729 9983
rect 11569 9823 11621 9875
rect 11677 9823 11706 9875
rect 11706 9823 11729 9875
rect 11569 9715 11621 9767
rect 11677 9715 11706 9767
rect 11706 9715 11729 9767
rect 11569 9607 11621 9659
rect 11677 9607 11706 9659
rect 11706 9607 11729 9659
rect 11569 9499 11621 9551
rect 11677 9499 11706 9551
rect 11706 9499 11729 9551
rect 11569 9391 11621 9443
rect 11677 9391 11706 9443
rect 11706 9391 11729 9443
rect 11569 9283 11621 9335
rect 11677 9283 11706 9335
rect 11706 9283 11729 9335
rect 11569 9175 11621 9227
rect 11677 9175 11706 9227
rect 11706 9175 11729 9227
rect 11569 9067 11621 9119
rect 11677 9067 11706 9119
rect 11706 9067 11729 9119
rect 11569 8959 11621 9011
rect 11677 8959 11706 9011
rect 11706 8959 11729 9011
rect 11569 8851 11621 8903
rect 11677 8851 11706 8903
rect 11706 8851 11729 8903
rect 11569 8743 11621 8795
rect 11677 8743 11706 8795
rect 11706 8743 11729 8795
rect 11569 8635 11621 8687
rect 11677 8635 11706 8687
rect 11706 8635 11729 8687
rect 11569 8527 11621 8579
rect 11677 8527 11706 8579
rect 11706 8527 11729 8579
rect 11569 8419 11621 8471
rect 11677 8419 11706 8471
rect 11706 8419 11729 8471
rect 11569 8311 11621 8363
rect 11677 8311 11706 8363
rect 11706 8311 11729 8363
rect 11569 8203 11621 8255
rect 11677 8203 11706 8255
rect 11706 8203 11729 8255
rect 11569 8095 11621 8147
rect 11677 8095 11706 8147
rect 11706 8095 11729 8147
rect 11569 7987 11621 8039
rect 11677 7987 11706 8039
rect 11706 7987 11729 8039
rect 11569 7879 11621 7931
rect 11677 7879 11706 7931
rect 11706 7879 11729 7931
rect 11569 7771 11621 7823
rect 11677 7771 11706 7823
rect 11706 7771 11729 7823
rect 11569 7663 11621 7715
rect 11677 7663 11706 7715
rect 11706 7663 11729 7715
rect 11569 7555 11621 7607
rect 11677 7555 11706 7607
rect 11706 7555 11729 7607
rect 11569 7447 11621 7499
rect 11677 7447 11706 7499
rect 11706 7447 11729 7499
rect 11569 7339 11621 7391
rect 11677 7339 11729 7391
rect 3433 7324 3485 7327
rect 3541 7324 3593 7327
rect 3649 7324 3701 7327
rect 3757 7324 3809 7327
rect 3865 7324 3917 7327
rect 3973 7324 4025 7327
rect 4081 7324 4133 7327
rect 4189 7324 4241 7327
rect 4297 7324 4349 7327
rect 4405 7324 4457 7327
rect 4513 7324 4565 7327
rect 4621 7324 4673 7327
rect 4729 7324 4781 7327
rect 4837 7324 4889 7327
rect 4945 7324 4997 7327
rect 5053 7324 5105 7327
rect 5161 7324 5213 7327
rect 6566 7324 6618 7327
rect 6674 7324 6726 7327
rect 6782 7324 6834 7327
rect 6890 7324 6942 7327
rect 6998 7324 7050 7327
rect 7106 7324 7158 7327
rect 7214 7324 7266 7327
rect 7322 7324 7374 7327
rect 7430 7324 7482 7327
rect 7538 7324 7590 7327
rect 9677 7324 9729 7327
rect 9785 7324 9837 7327
rect 9893 7324 9945 7327
rect 10001 7324 10053 7327
rect 10109 7324 10161 7327
rect 10217 7324 10269 7327
rect 10325 7324 10377 7327
rect 10433 7324 10485 7327
rect 10541 7324 10593 7327
rect 10649 7324 10701 7327
rect 10757 7324 10809 7327
rect 10865 7324 10917 7327
rect 10973 7324 11025 7327
rect 11081 7324 11133 7327
rect 11189 7324 11241 7327
rect 11297 7324 11349 7327
rect 11405 7324 11457 7327
rect 3433 7278 3485 7324
rect 3541 7278 3593 7324
rect 3649 7278 3701 7324
rect 3757 7278 3809 7324
rect 3865 7278 3917 7324
rect 3973 7278 4025 7324
rect 4081 7278 4133 7324
rect 4189 7278 4241 7324
rect 4297 7278 4349 7324
rect 4405 7278 4457 7324
rect 4513 7278 4565 7324
rect 4621 7278 4673 7324
rect 4729 7278 4781 7324
rect 4837 7278 4889 7324
rect 4945 7278 4997 7324
rect 5053 7278 5105 7324
rect 5161 7278 5213 7324
rect 6566 7278 6618 7324
rect 6674 7278 6726 7324
rect 6782 7278 6834 7324
rect 6890 7278 6942 7324
rect 6998 7278 7050 7324
rect 7106 7278 7158 7324
rect 7214 7278 7266 7324
rect 7322 7278 7374 7324
rect 7430 7278 7482 7324
rect 7538 7278 7590 7324
rect 9677 7278 9729 7324
rect 9785 7278 9837 7324
rect 9893 7278 9945 7324
rect 10001 7278 10053 7324
rect 10109 7278 10161 7324
rect 10217 7278 10269 7324
rect 10325 7278 10377 7324
rect 10433 7278 10485 7324
rect 10541 7278 10593 7324
rect 10649 7278 10701 7324
rect 10757 7278 10809 7324
rect 10865 7278 10917 7324
rect 10973 7278 11025 7324
rect 11081 7278 11133 7324
rect 11189 7278 11241 7324
rect 11297 7278 11349 7324
rect 11405 7278 11457 7324
rect 3433 7275 3485 7278
rect 3541 7275 3593 7278
rect 3649 7275 3701 7278
rect 3757 7275 3809 7278
rect 3865 7275 3917 7278
rect 3973 7275 4025 7278
rect 4081 7275 4133 7278
rect 4189 7275 4241 7278
rect 4297 7275 4349 7278
rect 4405 7275 4457 7278
rect 4513 7275 4565 7278
rect 4621 7275 4673 7278
rect 4729 7275 4781 7278
rect 4837 7275 4889 7278
rect 4945 7275 4997 7278
rect 5053 7275 5105 7278
rect 5161 7275 5213 7278
rect 6566 7275 6618 7278
rect 6674 7275 6726 7278
rect 6782 7275 6834 7278
rect 6890 7275 6942 7278
rect 6998 7275 7050 7278
rect 7106 7275 7158 7278
rect 7214 7275 7266 7278
rect 7322 7275 7374 7278
rect 7430 7275 7482 7278
rect 7538 7275 7590 7278
rect 9677 7275 9729 7278
rect 9785 7275 9837 7278
rect 9893 7275 9945 7278
rect 10001 7275 10053 7278
rect 10109 7275 10161 7278
rect 10217 7275 10269 7278
rect 10325 7275 10377 7278
rect 10433 7275 10485 7278
rect 10541 7275 10593 7278
rect 10649 7275 10701 7278
rect 10757 7275 10809 7278
rect 10865 7275 10917 7278
rect 10973 7275 11025 7278
rect 11081 7275 11133 7278
rect 11189 7275 11241 7278
rect 11297 7275 11349 7278
rect 11405 7275 11457 7278
rect 12051 12489 12103 12541
rect 12159 12489 12211 12541
rect 12267 12489 12319 12541
rect 12051 12381 12103 12433
rect 12159 12381 12211 12433
rect 12267 12381 12319 12433
rect 12051 12273 12103 12325
rect 12159 12273 12211 12325
rect 12267 12273 12319 12325
rect 12051 12165 12103 12217
rect 12159 12165 12211 12217
rect 12267 12165 12319 12217
rect 12051 12057 12103 12109
rect 12159 12057 12211 12109
rect 12267 12057 12319 12109
rect 12051 11949 12103 12001
rect 12159 11949 12211 12001
rect 12267 11949 12319 12001
rect 12051 11841 12103 11893
rect 12159 11841 12211 11893
rect 12267 11841 12319 11893
rect 12051 11733 12103 11785
rect 12159 11733 12211 11785
rect 12267 11733 12319 11785
rect 12051 11625 12103 11677
rect 12159 11625 12211 11677
rect 12267 11625 12319 11677
rect 12051 11517 12103 11569
rect 12159 11517 12211 11569
rect 12267 11517 12319 11569
rect 12051 11409 12103 11461
rect 12159 11409 12211 11461
rect 12267 11409 12319 11461
rect 12051 11301 12103 11353
rect 12159 11301 12211 11353
rect 12267 11301 12319 11353
rect 12051 11193 12103 11245
rect 12159 11193 12211 11245
rect 12267 11193 12319 11245
rect 12051 11085 12103 11137
rect 12159 11085 12211 11137
rect 12267 11085 12319 11137
rect 12051 10977 12103 11029
rect 12159 10977 12211 11029
rect 12267 10977 12319 11029
rect 12051 10869 12103 10921
rect 12159 10869 12211 10921
rect 12267 10869 12319 10921
rect 12051 10761 12103 10813
rect 12159 10761 12211 10813
rect 12267 10761 12319 10813
rect 12051 10653 12103 10705
rect 12159 10653 12211 10705
rect 12267 10653 12319 10705
rect 12051 10545 12103 10597
rect 12159 10545 12211 10597
rect 12267 10545 12319 10597
rect 12051 10437 12103 10489
rect 12159 10437 12211 10489
rect 12267 10437 12319 10489
rect 12051 10329 12103 10381
rect 12159 10329 12211 10381
rect 12267 10329 12319 10381
rect 12051 10221 12103 10273
rect 12159 10221 12211 10273
rect 12267 10221 12319 10273
rect 12051 10113 12103 10165
rect 12159 10113 12211 10165
rect 12267 10113 12319 10165
rect 12051 10005 12103 10057
rect 12159 10005 12211 10057
rect 12267 10005 12319 10057
rect 12051 9897 12103 9949
rect 12159 9897 12211 9949
rect 12267 9897 12319 9949
rect 12051 9789 12103 9841
rect 12159 9789 12211 9841
rect 12267 9789 12319 9841
rect 12051 9681 12103 9733
rect 12159 9681 12211 9733
rect 12267 9681 12319 9733
rect 12051 9573 12103 9625
rect 12159 9573 12211 9625
rect 12267 9573 12319 9625
rect 12051 9465 12103 9517
rect 12159 9465 12211 9517
rect 12267 9465 12319 9517
rect 12051 9357 12103 9409
rect 12159 9357 12211 9409
rect 12267 9357 12319 9409
rect 12051 9249 12103 9301
rect 12159 9249 12211 9301
rect 12267 9249 12319 9301
rect 12051 9141 12103 9193
rect 12159 9141 12211 9193
rect 12267 9141 12319 9193
rect 12051 9033 12103 9085
rect 12159 9033 12211 9085
rect 12267 9033 12319 9085
rect 12051 8925 12103 8977
rect 12159 8925 12211 8977
rect 12267 8925 12319 8977
rect 12051 8817 12103 8869
rect 12159 8817 12211 8869
rect 12267 8817 12319 8869
rect 12051 8709 12103 8761
rect 12159 8709 12211 8761
rect 12267 8709 12319 8761
rect 12051 8601 12103 8653
rect 12159 8601 12211 8653
rect 12267 8601 12319 8653
rect 12051 8493 12103 8545
rect 12159 8493 12211 8545
rect 12267 8493 12319 8545
rect 12051 8385 12103 8437
rect 12159 8385 12211 8437
rect 12267 8385 12319 8437
rect 12051 8277 12103 8329
rect 12159 8277 12211 8329
rect 12267 8277 12319 8329
rect 12051 8169 12103 8221
rect 12159 8169 12211 8221
rect 12267 8169 12319 8221
rect 12051 8061 12103 8113
rect 12159 8061 12211 8113
rect 12267 8061 12319 8113
rect 12051 7953 12103 8005
rect 12159 7953 12211 8005
rect 12267 7953 12319 8005
rect 12051 7845 12103 7897
rect 12159 7845 12211 7897
rect 12267 7845 12319 7897
rect 12051 7737 12103 7789
rect 12159 7737 12211 7789
rect 12267 7737 12319 7789
rect 12051 7629 12103 7681
rect 12159 7629 12211 7681
rect 12267 7629 12319 7681
rect 12051 7521 12103 7573
rect 12159 7521 12211 7573
rect 12267 7521 12319 7573
rect 12051 7413 12103 7465
rect 12159 7413 12211 7465
rect 12267 7413 12319 7465
rect 12051 7305 12103 7357
rect 12159 7305 12211 7357
rect 12267 7305 12319 7357
rect 12051 7197 12103 7249
rect 12159 7197 12211 7249
rect 12267 7197 12319 7249
rect 12051 7089 12103 7141
rect 12159 7089 12211 7141
rect 12267 7089 12319 7141
rect 12051 6981 12103 7033
rect 12159 6981 12211 7033
rect 12267 6981 12319 7033
rect 1505 6878 1557 6885
rect 1613 6878 1665 6885
rect 1721 6878 1773 6885
rect 1829 6878 1881 6885
rect 1937 6878 1989 6885
rect 2045 6878 2097 6885
rect 2153 6878 2205 6885
rect 2261 6878 2313 6885
rect 2369 6878 2421 6885
rect 2477 6878 2529 6885
rect 2585 6878 2637 6885
rect 2693 6878 2745 6885
rect 2801 6878 2853 6885
rect 2909 6878 2961 6885
rect 3017 6878 3069 6885
rect 3125 6878 3177 6885
rect 3233 6878 3285 6885
rect 5372 6878 5424 6885
rect 5480 6878 5532 6885
rect 5588 6878 5640 6885
rect 5696 6878 5748 6885
rect 5804 6878 5856 6885
rect 5912 6878 5964 6885
rect 6020 6878 6072 6885
rect 6128 6878 6180 6885
rect 6236 6878 6288 6885
rect 6344 6878 6396 6885
rect 7749 6878 7801 6885
rect 7857 6878 7909 6885
rect 7965 6878 8017 6885
rect 8073 6878 8125 6885
rect 8181 6878 8233 6885
rect 8289 6878 8341 6885
rect 8397 6878 8449 6885
rect 8505 6878 8557 6885
rect 8613 6878 8665 6885
rect 8721 6878 8773 6885
rect 8829 6878 8881 6885
rect 8937 6878 8989 6885
rect 9045 6878 9097 6885
rect 9153 6878 9205 6885
rect 9261 6878 9313 6885
rect 9369 6878 9421 6885
rect 9477 6878 9529 6885
rect 1505 6833 1557 6878
rect 1613 6833 1665 6878
rect 1721 6833 1773 6878
rect 1829 6833 1881 6878
rect 1937 6833 1989 6878
rect 2045 6833 2097 6878
rect 2153 6833 2205 6878
rect 2261 6833 2313 6878
rect 2369 6833 2421 6878
rect 2477 6833 2529 6878
rect 2585 6833 2637 6878
rect 2693 6833 2745 6878
rect 2801 6833 2853 6878
rect 2909 6833 2961 6878
rect 3017 6833 3069 6878
rect 3125 6833 3177 6878
rect 3233 6833 3285 6878
rect 5372 6833 5424 6878
rect 5480 6833 5532 6878
rect 5588 6833 5640 6878
rect 5696 6833 5748 6878
rect 5804 6833 5856 6878
rect 5912 6833 5964 6878
rect 6020 6833 6072 6878
rect 6128 6833 6180 6878
rect 6236 6833 6288 6878
rect 6344 6833 6396 6878
rect 7749 6833 7801 6878
rect 7857 6833 7909 6878
rect 7965 6833 8017 6878
rect 8073 6833 8125 6878
rect 8181 6833 8233 6878
rect 8289 6833 8341 6878
rect 8397 6833 8449 6878
rect 8505 6833 8557 6878
rect 8613 6833 8665 6878
rect 8721 6833 8773 6878
rect 8829 6833 8881 6878
rect 8937 6833 8989 6878
rect 9045 6833 9097 6878
rect 9153 6833 9205 6878
rect 9261 6833 9313 6878
rect 9369 6833 9421 6878
rect 9477 6833 9529 6878
rect 1505 6732 1557 6777
rect 1613 6732 1665 6777
rect 1721 6732 1773 6777
rect 1829 6732 1881 6777
rect 1937 6732 1989 6777
rect 2045 6732 2097 6777
rect 2153 6732 2205 6777
rect 2261 6732 2313 6777
rect 2369 6732 2421 6777
rect 2477 6732 2529 6777
rect 2585 6732 2637 6777
rect 2693 6732 2745 6777
rect 2801 6732 2853 6777
rect 2909 6732 2961 6777
rect 3017 6732 3069 6777
rect 3125 6732 3177 6777
rect 3233 6732 3285 6777
rect 5372 6732 5424 6777
rect 5480 6732 5532 6777
rect 5588 6732 5640 6777
rect 5696 6732 5748 6777
rect 5804 6732 5856 6777
rect 5912 6732 5964 6777
rect 6020 6732 6072 6777
rect 6128 6732 6180 6777
rect 6236 6732 6288 6777
rect 6344 6732 6396 6777
rect 7749 6732 7801 6777
rect 7857 6732 7909 6777
rect 7965 6732 8017 6777
rect 8073 6732 8125 6777
rect 8181 6732 8233 6777
rect 8289 6732 8341 6777
rect 8397 6732 8449 6777
rect 8505 6732 8557 6777
rect 8613 6732 8665 6777
rect 8721 6732 8773 6777
rect 8829 6732 8881 6777
rect 8937 6732 8989 6777
rect 9045 6732 9097 6777
rect 9153 6732 9205 6777
rect 9261 6732 9313 6777
rect 9369 6732 9421 6777
rect 9477 6732 9529 6777
rect 12051 6873 12103 6925
rect 12159 6873 12211 6925
rect 12267 6873 12319 6925
rect 12051 6765 12103 6817
rect 12159 6765 12211 6817
rect 12267 6765 12319 6817
rect 1505 6725 1557 6732
rect 1613 6725 1665 6732
rect 1721 6725 1773 6732
rect 1829 6725 1881 6732
rect 1937 6725 1989 6732
rect 2045 6725 2097 6732
rect 2153 6725 2205 6732
rect 2261 6725 2313 6732
rect 2369 6725 2421 6732
rect 2477 6725 2529 6732
rect 2585 6725 2637 6732
rect 2693 6725 2745 6732
rect 2801 6725 2853 6732
rect 2909 6725 2961 6732
rect 3017 6725 3069 6732
rect 3125 6725 3177 6732
rect 3233 6725 3285 6732
rect 5372 6725 5424 6732
rect 5480 6725 5532 6732
rect 5588 6725 5640 6732
rect 5696 6725 5748 6732
rect 5804 6725 5856 6732
rect 5912 6725 5964 6732
rect 6020 6725 6072 6732
rect 6128 6725 6180 6732
rect 6236 6725 6288 6732
rect 6344 6725 6396 6732
rect 7749 6725 7801 6732
rect 7857 6725 7909 6732
rect 7965 6725 8017 6732
rect 8073 6725 8125 6732
rect 8181 6725 8233 6732
rect 8289 6725 8341 6732
rect 8397 6725 8449 6732
rect 8505 6725 8557 6732
rect 8613 6725 8665 6732
rect 8721 6725 8773 6732
rect 8829 6725 8881 6732
rect 8937 6725 8989 6732
rect 9045 6725 9097 6732
rect 9153 6725 9205 6732
rect 9261 6725 9313 6732
rect 9369 6725 9421 6732
rect 9477 6725 9529 6732
rect 3433 6332 3485 6335
rect 3541 6332 3593 6335
rect 3649 6332 3701 6335
rect 3757 6332 3809 6335
rect 3865 6332 3917 6335
rect 3973 6332 4025 6335
rect 4081 6332 4133 6335
rect 4189 6332 4241 6335
rect 4297 6332 4349 6335
rect 4405 6332 4457 6335
rect 4513 6332 4565 6335
rect 4621 6332 4673 6335
rect 4729 6332 4781 6335
rect 4837 6332 4889 6335
rect 4945 6332 4997 6335
rect 5053 6332 5105 6335
rect 5161 6332 5213 6335
rect 6566 6332 6618 6335
rect 6674 6332 6726 6335
rect 6782 6332 6834 6335
rect 6890 6332 6942 6335
rect 6998 6332 7050 6335
rect 7106 6332 7158 6335
rect 7214 6332 7266 6335
rect 7322 6332 7374 6335
rect 7430 6332 7482 6335
rect 7538 6332 7590 6335
rect 9677 6332 9729 6335
rect 9785 6332 9837 6335
rect 9893 6332 9945 6335
rect 10001 6332 10053 6335
rect 10109 6332 10161 6335
rect 10217 6332 10269 6335
rect 10325 6332 10377 6335
rect 10433 6332 10485 6335
rect 10541 6332 10593 6335
rect 10649 6332 10701 6335
rect 10757 6332 10809 6335
rect 10865 6332 10917 6335
rect 10973 6332 11025 6335
rect 11081 6332 11133 6335
rect 11189 6332 11241 6335
rect 11297 6332 11349 6335
rect 11405 6332 11457 6335
rect 3433 6286 3485 6332
rect 3541 6286 3593 6332
rect 3649 6286 3701 6332
rect 3757 6286 3809 6332
rect 3865 6286 3917 6332
rect 3973 6286 4025 6332
rect 4081 6286 4133 6332
rect 4189 6286 4241 6332
rect 4297 6286 4349 6332
rect 4405 6286 4457 6332
rect 4513 6286 4565 6332
rect 4621 6286 4673 6332
rect 4729 6286 4781 6332
rect 4837 6286 4889 6332
rect 4945 6286 4997 6332
rect 5053 6286 5105 6332
rect 5161 6286 5213 6332
rect 6566 6286 6618 6332
rect 6674 6286 6726 6332
rect 6782 6286 6834 6332
rect 6890 6286 6942 6332
rect 6998 6286 7050 6332
rect 7106 6286 7158 6332
rect 7214 6286 7266 6332
rect 7322 6286 7374 6332
rect 7430 6286 7482 6332
rect 7538 6286 7590 6332
rect 9677 6286 9729 6332
rect 9785 6286 9837 6332
rect 9893 6286 9945 6332
rect 10001 6286 10053 6332
rect 10109 6286 10161 6332
rect 10217 6286 10269 6332
rect 10325 6286 10377 6332
rect 10433 6286 10485 6332
rect 10541 6286 10593 6332
rect 10649 6286 10701 6332
rect 10757 6286 10809 6332
rect 10865 6286 10917 6332
rect 10973 6286 11025 6332
rect 11081 6286 11133 6332
rect 11189 6286 11241 6332
rect 11297 6286 11349 6332
rect 11405 6286 11457 6332
rect 3433 6283 3485 6286
rect 3541 6283 3593 6286
rect 3649 6283 3701 6286
rect 3757 6283 3809 6286
rect 3865 6283 3917 6286
rect 3973 6283 4025 6286
rect 4081 6283 4133 6286
rect 4189 6283 4241 6286
rect 4297 6283 4349 6286
rect 4405 6283 4457 6286
rect 4513 6283 4565 6286
rect 4621 6283 4673 6286
rect 4729 6283 4781 6286
rect 4837 6283 4889 6286
rect 4945 6283 4997 6286
rect 5053 6283 5105 6286
rect 5161 6283 5213 6286
rect 6566 6283 6618 6286
rect 6674 6283 6726 6286
rect 6782 6283 6834 6286
rect 6890 6283 6942 6286
rect 6998 6283 7050 6286
rect 7106 6283 7158 6286
rect 7214 6283 7266 6286
rect 7322 6283 7374 6286
rect 7430 6283 7482 6286
rect 7538 6283 7590 6286
rect 9677 6283 9729 6286
rect 9785 6283 9837 6286
rect 9893 6283 9945 6286
rect 10001 6283 10053 6286
rect 10109 6283 10161 6286
rect 10217 6283 10269 6286
rect 10325 6283 10377 6286
rect 10433 6283 10485 6286
rect 10541 6283 10593 6286
rect 10649 6283 10701 6286
rect 10757 6283 10809 6286
rect 10865 6283 10917 6286
rect 10973 6283 11025 6286
rect 11081 6283 11133 6286
rect 11189 6283 11241 6286
rect 11297 6283 11349 6286
rect 11405 6283 11457 6286
rect 1233 6219 1285 6271
rect 1341 6219 1393 6271
rect 1233 6111 1256 6163
rect 1256 6111 1285 6163
rect 1341 6111 1393 6163
rect 1233 6003 1256 6055
rect 1256 6003 1285 6055
rect 1341 6003 1393 6055
rect 1233 5895 1256 5947
rect 1256 5895 1285 5947
rect 1341 5895 1393 5947
rect 1233 5787 1256 5839
rect 1256 5787 1285 5839
rect 1341 5787 1393 5839
rect 1233 5679 1256 5731
rect 1256 5679 1285 5731
rect 1341 5679 1393 5731
rect 1233 5571 1256 5623
rect 1256 5571 1285 5623
rect 1341 5571 1393 5623
rect 1233 5463 1256 5515
rect 1256 5463 1285 5515
rect 1341 5463 1393 5515
rect 1233 5355 1256 5407
rect 1256 5355 1285 5407
rect 1341 5355 1393 5407
rect 1233 5247 1256 5299
rect 1256 5247 1285 5299
rect 1341 5247 1393 5299
rect 1233 5139 1256 5191
rect 1256 5139 1285 5191
rect 1341 5139 1393 5191
rect 1233 5031 1256 5083
rect 1256 5031 1285 5083
rect 1341 5031 1393 5083
rect 1233 4923 1256 4975
rect 1256 4923 1285 4975
rect 1341 4923 1393 4975
rect 1233 4815 1256 4867
rect 1256 4815 1285 4867
rect 1341 4815 1393 4867
rect 1233 4707 1256 4759
rect 1256 4707 1285 4759
rect 1341 4707 1393 4759
rect 1233 4599 1256 4651
rect 1256 4599 1285 4651
rect 1341 4599 1393 4651
rect 1233 4491 1256 4543
rect 1256 4491 1285 4543
rect 1341 4491 1393 4543
rect 1233 4383 1256 4435
rect 1256 4383 1285 4435
rect 1341 4383 1393 4435
rect 1233 4275 1256 4327
rect 1256 4275 1285 4327
rect 1341 4275 1393 4327
rect 1233 4167 1256 4219
rect 1256 4167 1285 4219
rect 1341 4167 1393 4219
rect 1233 4059 1256 4111
rect 1256 4059 1285 4111
rect 1341 4059 1393 4111
rect 1233 3951 1256 4003
rect 1256 3951 1285 4003
rect 1341 3951 1393 4003
rect 1233 3843 1256 3895
rect 1256 3843 1285 3895
rect 1341 3843 1393 3895
rect 1233 3735 1256 3787
rect 1256 3735 1285 3787
rect 1341 3735 1393 3787
rect 1233 3627 1256 3679
rect 1256 3627 1285 3679
rect 1341 3627 1393 3679
rect 1233 3519 1256 3571
rect 1256 3519 1285 3571
rect 1341 3519 1393 3571
rect 1233 3411 1256 3463
rect 1256 3411 1285 3463
rect 1341 3411 1393 3463
rect 1233 3303 1256 3355
rect 1256 3303 1285 3355
rect 1341 3303 1393 3355
rect 1233 3195 1256 3247
rect 1256 3195 1285 3247
rect 1341 3195 1393 3247
rect 1233 3087 1256 3139
rect 1256 3087 1285 3139
rect 1341 3087 1393 3139
rect 1233 2979 1256 3031
rect 1256 2979 1285 3031
rect 1341 2979 1393 3031
rect 1233 2871 1256 2923
rect 1256 2871 1285 2923
rect 1341 2871 1393 2923
rect 1233 2763 1256 2815
rect 1256 2763 1285 2815
rect 1341 2763 1393 2815
rect 1233 2655 1256 2707
rect 1256 2655 1285 2707
rect 1341 2655 1393 2707
rect 1233 2547 1256 2599
rect 1256 2547 1285 2599
rect 1341 2547 1393 2599
rect 1233 2439 1256 2491
rect 1256 2439 1285 2491
rect 1341 2439 1393 2491
rect 1233 2331 1256 2383
rect 1256 2331 1285 2383
rect 1341 2331 1393 2383
rect 1233 2223 1256 2275
rect 1256 2223 1285 2275
rect 1341 2223 1393 2275
rect 1233 2115 1256 2167
rect 1256 2115 1285 2167
rect 1341 2115 1393 2167
rect 1233 2007 1256 2059
rect 1256 2007 1285 2059
rect 1341 2007 1393 2059
rect 1233 1899 1256 1951
rect 1256 1899 1285 1951
rect 1341 1899 1393 1951
rect 1233 1791 1256 1843
rect 1256 1791 1285 1843
rect 1341 1791 1393 1843
rect 1233 1683 1256 1735
rect 1256 1683 1285 1735
rect 1341 1683 1393 1735
rect 1233 1575 1256 1627
rect 1256 1575 1285 1627
rect 1341 1575 1393 1627
rect 11569 6219 11621 6271
rect 11677 6219 11729 6271
rect 1505 6088 1557 6091
rect 1613 6088 1665 6091
rect 1721 6088 1773 6091
rect 1829 6088 1881 6091
rect 1937 6088 1989 6091
rect 2045 6088 2097 6091
rect 2153 6088 2205 6091
rect 2261 6088 2313 6091
rect 2369 6088 2421 6091
rect 2477 6088 2529 6091
rect 2585 6088 2637 6091
rect 2693 6088 2745 6091
rect 2801 6088 2853 6091
rect 2909 6088 2961 6091
rect 3017 6088 3069 6091
rect 3125 6088 3177 6091
rect 3233 6088 3285 6091
rect 5372 6088 5424 6091
rect 5480 6088 5532 6091
rect 5588 6088 5640 6091
rect 5696 6088 5748 6091
rect 5804 6088 5856 6091
rect 5912 6088 5964 6091
rect 6020 6088 6072 6091
rect 6128 6088 6180 6091
rect 6236 6088 6288 6091
rect 6344 6088 6396 6091
rect 7749 6088 7801 6091
rect 7857 6088 7909 6091
rect 7965 6088 8017 6091
rect 8073 6088 8125 6091
rect 8181 6088 8233 6091
rect 8289 6088 8341 6091
rect 8397 6088 8449 6091
rect 8505 6088 8557 6091
rect 8613 6088 8665 6091
rect 8721 6088 8773 6091
rect 8829 6088 8881 6091
rect 8937 6088 8989 6091
rect 9045 6088 9097 6091
rect 9153 6088 9205 6091
rect 9261 6088 9313 6091
rect 9369 6088 9421 6091
rect 9477 6088 9529 6091
rect 1505 6042 1557 6088
rect 1613 6042 1665 6088
rect 1721 6042 1773 6088
rect 1829 6042 1881 6088
rect 1937 6042 1989 6088
rect 2045 6042 2097 6088
rect 2153 6042 2205 6088
rect 2261 6042 2313 6088
rect 2369 6042 2421 6088
rect 2477 6042 2529 6088
rect 2585 6042 2637 6088
rect 2693 6042 2745 6088
rect 2801 6042 2853 6088
rect 2909 6042 2961 6088
rect 3017 6042 3069 6088
rect 3125 6042 3177 6088
rect 3233 6042 3285 6088
rect 5372 6042 5424 6088
rect 5480 6042 5532 6088
rect 5588 6042 5640 6088
rect 5696 6042 5748 6088
rect 5804 6042 5856 6088
rect 5912 6042 5964 6088
rect 6020 6042 6072 6088
rect 6128 6042 6180 6088
rect 6236 6042 6288 6088
rect 6344 6042 6396 6088
rect 7749 6042 7801 6088
rect 7857 6042 7909 6088
rect 7965 6042 8017 6088
rect 8073 6042 8125 6088
rect 8181 6042 8233 6088
rect 8289 6042 8341 6088
rect 8397 6042 8449 6088
rect 8505 6042 8557 6088
rect 8613 6042 8665 6088
rect 8721 6042 8773 6088
rect 8829 6042 8881 6088
rect 8937 6042 8989 6088
rect 9045 6042 9097 6088
rect 9153 6042 9205 6088
rect 9261 6042 9313 6088
rect 9369 6042 9421 6088
rect 9477 6042 9529 6088
rect 1505 6039 1557 6042
rect 1613 6039 1665 6042
rect 1721 6039 1773 6042
rect 1829 6039 1881 6042
rect 1937 6039 1989 6042
rect 2045 6039 2097 6042
rect 2153 6039 2205 6042
rect 2261 6039 2313 6042
rect 2369 6039 2421 6042
rect 2477 6039 2529 6042
rect 2585 6039 2637 6042
rect 2693 6039 2745 6042
rect 2801 6039 2853 6042
rect 2909 6039 2961 6042
rect 3017 6039 3069 6042
rect 3125 6039 3177 6042
rect 3233 6039 3285 6042
rect 5372 6039 5424 6042
rect 5480 6039 5532 6042
rect 5588 6039 5640 6042
rect 5696 6039 5748 6042
rect 5804 6039 5856 6042
rect 5912 6039 5964 6042
rect 6020 6039 6072 6042
rect 6128 6039 6180 6042
rect 6236 6039 6288 6042
rect 6344 6039 6396 6042
rect 7749 6039 7801 6042
rect 7857 6039 7909 6042
rect 7965 6039 8017 6042
rect 8073 6039 8125 6042
rect 8181 6039 8233 6042
rect 8289 6039 8341 6042
rect 8397 6039 8449 6042
rect 8505 6039 8557 6042
rect 8613 6039 8665 6042
rect 8721 6039 8773 6042
rect 8829 6039 8881 6042
rect 8937 6039 8989 6042
rect 9045 6039 9097 6042
rect 9153 6039 9205 6042
rect 9261 6039 9313 6042
rect 9369 6039 9421 6042
rect 9477 6039 9529 6042
rect 3433 5844 3485 5847
rect 3541 5844 3593 5847
rect 3649 5844 3701 5847
rect 3757 5844 3809 5847
rect 3865 5844 3917 5847
rect 3973 5844 4025 5847
rect 4081 5844 4133 5847
rect 4189 5844 4241 5847
rect 4297 5844 4349 5847
rect 4405 5844 4457 5847
rect 4513 5844 4565 5847
rect 4621 5844 4673 5847
rect 4729 5844 4781 5847
rect 4837 5844 4889 5847
rect 4945 5844 4997 5847
rect 5053 5844 5105 5847
rect 5161 5844 5213 5847
rect 6566 5844 6618 5847
rect 6674 5844 6726 5847
rect 6782 5844 6834 5847
rect 6890 5844 6942 5847
rect 6998 5844 7050 5847
rect 7106 5844 7158 5847
rect 7214 5844 7266 5847
rect 7322 5844 7374 5847
rect 7430 5844 7482 5847
rect 7538 5844 7590 5847
rect 9677 5844 9729 5847
rect 9785 5844 9837 5847
rect 9893 5844 9945 5847
rect 10001 5844 10053 5847
rect 10109 5844 10161 5847
rect 10217 5844 10269 5847
rect 10325 5844 10377 5847
rect 10433 5844 10485 5847
rect 10541 5844 10593 5847
rect 10649 5844 10701 5847
rect 10757 5844 10809 5847
rect 10865 5844 10917 5847
rect 10973 5844 11025 5847
rect 11081 5844 11133 5847
rect 11189 5844 11241 5847
rect 11297 5844 11349 5847
rect 11405 5844 11457 5847
rect 3433 5798 3485 5844
rect 3541 5798 3593 5844
rect 3649 5798 3701 5844
rect 3757 5798 3809 5844
rect 3865 5798 3917 5844
rect 3973 5798 4025 5844
rect 4081 5798 4133 5844
rect 4189 5798 4241 5844
rect 4297 5798 4349 5844
rect 4405 5798 4457 5844
rect 4513 5798 4565 5844
rect 4621 5798 4673 5844
rect 4729 5798 4781 5844
rect 4837 5798 4889 5844
rect 4945 5798 4997 5844
rect 5053 5798 5105 5844
rect 5161 5798 5213 5844
rect 6566 5798 6618 5844
rect 6674 5798 6726 5844
rect 6782 5798 6834 5844
rect 6890 5798 6942 5844
rect 6998 5798 7050 5844
rect 7106 5798 7158 5844
rect 7214 5798 7266 5844
rect 7322 5798 7374 5844
rect 7430 5798 7482 5844
rect 7538 5798 7590 5844
rect 9677 5798 9729 5844
rect 9785 5798 9837 5844
rect 9893 5798 9945 5844
rect 10001 5798 10053 5844
rect 10109 5798 10161 5844
rect 10217 5798 10269 5844
rect 10325 5798 10377 5844
rect 10433 5798 10485 5844
rect 10541 5798 10593 5844
rect 10649 5798 10701 5844
rect 10757 5798 10809 5844
rect 10865 5798 10917 5844
rect 10973 5798 11025 5844
rect 11081 5798 11133 5844
rect 11189 5798 11241 5844
rect 11297 5798 11349 5844
rect 11405 5798 11457 5844
rect 3433 5795 3485 5798
rect 3541 5795 3593 5798
rect 3649 5795 3701 5798
rect 3757 5795 3809 5798
rect 3865 5795 3917 5798
rect 3973 5795 4025 5798
rect 4081 5795 4133 5798
rect 4189 5795 4241 5798
rect 4297 5795 4349 5798
rect 4405 5795 4457 5798
rect 4513 5795 4565 5798
rect 4621 5795 4673 5798
rect 4729 5795 4781 5798
rect 4837 5795 4889 5798
rect 4945 5795 4997 5798
rect 5053 5795 5105 5798
rect 5161 5795 5213 5798
rect 6566 5795 6618 5798
rect 6674 5795 6726 5798
rect 6782 5795 6834 5798
rect 6890 5795 6942 5798
rect 6998 5795 7050 5798
rect 7106 5795 7158 5798
rect 7214 5795 7266 5798
rect 7322 5795 7374 5798
rect 7430 5795 7482 5798
rect 7538 5795 7590 5798
rect 9677 5795 9729 5798
rect 9785 5795 9837 5798
rect 9893 5795 9945 5798
rect 10001 5795 10053 5798
rect 10109 5795 10161 5798
rect 10217 5795 10269 5798
rect 10325 5795 10377 5798
rect 10433 5795 10485 5798
rect 10541 5795 10593 5798
rect 10649 5795 10701 5798
rect 10757 5795 10809 5798
rect 10865 5795 10917 5798
rect 10973 5795 11025 5798
rect 11081 5795 11133 5798
rect 11189 5795 11241 5798
rect 11297 5795 11349 5798
rect 11405 5795 11457 5798
rect 1505 5600 1557 5603
rect 1613 5600 1665 5603
rect 1721 5600 1773 5603
rect 1829 5600 1881 5603
rect 1937 5600 1989 5603
rect 2045 5600 2097 5603
rect 2153 5600 2205 5603
rect 2261 5600 2313 5603
rect 2369 5600 2421 5603
rect 2477 5600 2529 5603
rect 2585 5600 2637 5603
rect 2693 5600 2745 5603
rect 2801 5600 2853 5603
rect 2909 5600 2961 5603
rect 3017 5600 3069 5603
rect 3125 5600 3177 5603
rect 3233 5600 3285 5603
rect 5372 5600 5424 5603
rect 5480 5600 5532 5603
rect 5588 5600 5640 5603
rect 5696 5600 5748 5603
rect 5804 5600 5856 5603
rect 5912 5600 5964 5603
rect 6020 5600 6072 5603
rect 6128 5600 6180 5603
rect 6236 5600 6288 5603
rect 6344 5600 6396 5603
rect 7749 5600 7801 5603
rect 7857 5600 7909 5603
rect 7965 5600 8017 5603
rect 8073 5600 8125 5603
rect 8181 5600 8233 5603
rect 8289 5600 8341 5603
rect 8397 5600 8449 5603
rect 8505 5600 8557 5603
rect 8613 5600 8665 5603
rect 8721 5600 8773 5603
rect 8829 5600 8881 5603
rect 8937 5600 8989 5603
rect 9045 5600 9097 5603
rect 9153 5600 9205 5603
rect 9261 5600 9313 5603
rect 9369 5600 9421 5603
rect 9477 5600 9529 5603
rect 1505 5554 1557 5600
rect 1613 5554 1665 5600
rect 1721 5554 1773 5600
rect 1829 5554 1881 5600
rect 1937 5554 1989 5600
rect 2045 5554 2097 5600
rect 2153 5554 2205 5600
rect 2261 5554 2313 5600
rect 2369 5554 2421 5600
rect 2477 5554 2529 5600
rect 2585 5554 2637 5600
rect 2693 5554 2745 5600
rect 2801 5554 2853 5600
rect 2909 5554 2961 5600
rect 3017 5554 3069 5600
rect 3125 5554 3177 5600
rect 3233 5554 3285 5600
rect 5372 5554 5424 5600
rect 5480 5554 5532 5600
rect 5588 5554 5640 5600
rect 5696 5554 5748 5600
rect 5804 5554 5856 5600
rect 5912 5554 5964 5600
rect 6020 5554 6072 5600
rect 6128 5554 6180 5600
rect 6236 5554 6288 5600
rect 6344 5554 6396 5600
rect 7749 5554 7801 5600
rect 7857 5554 7909 5600
rect 7965 5554 8017 5600
rect 8073 5554 8125 5600
rect 8181 5554 8233 5600
rect 8289 5554 8341 5600
rect 8397 5554 8449 5600
rect 8505 5554 8557 5600
rect 8613 5554 8665 5600
rect 8721 5554 8773 5600
rect 8829 5554 8881 5600
rect 8937 5554 8989 5600
rect 9045 5554 9097 5600
rect 9153 5554 9205 5600
rect 9261 5554 9313 5600
rect 9369 5554 9421 5600
rect 9477 5554 9529 5600
rect 1505 5551 1557 5554
rect 1613 5551 1665 5554
rect 1721 5551 1773 5554
rect 1829 5551 1881 5554
rect 1937 5551 1989 5554
rect 2045 5551 2097 5554
rect 2153 5551 2205 5554
rect 2261 5551 2313 5554
rect 2369 5551 2421 5554
rect 2477 5551 2529 5554
rect 2585 5551 2637 5554
rect 2693 5551 2745 5554
rect 2801 5551 2853 5554
rect 2909 5551 2961 5554
rect 3017 5551 3069 5554
rect 3125 5551 3177 5554
rect 3233 5551 3285 5554
rect 5372 5551 5424 5554
rect 5480 5551 5532 5554
rect 5588 5551 5640 5554
rect 5696 5551 5748 5554
rect 5804 5551 5856 5554
rect 5912 5551 5964 5554
rect 6020 5551 6072 5554
rect 6128 5551 6180 5554
rect 6236 5551 6288 5554
rect 6344 5551 6396 5554
rect 7749 5551 7801 5554
rect 7857 5551 7909 5554
rect 7965 5551 8017 5554
rect 8073 5551 8125 5554
rect 8181 5551 8233 5554
rect 8289 5551 8341 5554
rect 8397 5551 8449 5554
rect 8505 5551 8557 5554
rect 8613 5551 8665 5554
rect 8721 5551 8773 5554
rect 8829 5551 8881 5554
rect 8937 5551 8989 5554
rect 9045 5551 9097 5554
rect 9153 5551 9205 5554
rect 9261 5551 9313 5554
rect 9369 5551 9421 5554
rect 9477 5551 9529 5554
rect 3433 5356 3485 5359
rect 3541 5356 3593 5359
rect 3649 5356 3701 5359
rect 3757 5356 3809 5359
rect 3865 5356 3917 5359
rect 3973 5356 4025 5359
rect 4081 5356 4133 5359
rect 4189 5356 4241 5359
rect 4297 5356 4349 5359
rect 4405 5356 4457 5359
rect 4513 5356 4565 5359
rect 4621 5356 4673 5359
rect 4729 5356 4781 5359
rect 4837 5356 4889 5359
rect 4945 5356 4997 5359
rect 5053 5356 5105 5359
rect 5161 5356 5213 5359
rect 6566 5356 6618 5359
rect 6674 5356 6726 5359
rect 6782 5356 6834 5359
rect 6890 5356 6942 5359
rect 6998 5356 7050 5359
rect 7106 5356 7158 5359
rect 7214 5356 7266 5359
rect 7322 5356 7374 5359
rect 7430 5356 7482 5359
rect 7538 5356 7590 5359
rect 9677 5356 9729 5359
rect 9785 5356 9837 5359
rect 9893 5356 9945 5359
rect 10001 5356 10053 5359
rect 10109 5356 10161 5359
rect 10217 5356 10269 5359
rect 10325 5356 10377 5359
rect 10433 5356 10485 5359
rect 10541 5356 10593 5359
rect 10649 5356 10701 5359
rect 10757 5356 10809 5359
rect 10865 5356 10917 5359
rect 10973 5356 11025 5359
rect 11081 5356 11133 5359
rect 11189 5356 11241 5359
rect 11297 5356 11349 5359
rect 11405 5356 11457 5359
rect 3433 5310 3485 5356
rect 3541 5310 3593 5356
rect 3649 5310 3701 5356
rect 3757 5310 3809 5356
rect 3865 5310 3917 5356
rect 3973 5310 4025 5356
rect 4081 5310 4133 5356
rect 4189 5310 4241 5356
rect 4297 5310 4349 5356
rect 4405 5310 4457 5356
rect 4513 5310 4565 5356
rect 4621 5310 4673 5356
rect 4729 5310 4781 5356
rect 4837 5310 4889 5356
rect 4945 5310 4997 5356
rect 5053 5310 5105 5356
rect 5161 5310 5213 5356
rect 6566 5310 6618 5356
rect 6674 5310 6726 5356
rect 6782 5310 6834 5356
rect 6890 5310 6942 5356
rect 6998 5310 7050 5356
rect 7106 5310 7158 5356
rect 7214 5310 7266 5356
rect 7322 5310 7374 5356
rect 7430 5310 7482 5356
rect 7538 5310 7590 5356
rect 9677 5310 9729 5356
rect 9785 5310 9837 5356
rect 9893 5310 9945 5356
rect 10001 5310 10053 5356
rect 10109 5310 10161 5356
rect 10217 5310 10269 5356
rect 10325 5310 10377 5356
rect 10433 5310 10485 5356
rect 10541 5310 10593 5356
rect 10649 5310 10701 5356
rect 10757 5310 10809 5356
rect 10865 5310 10917 5356
rect 10973 5310 11025 5356
rect 11081 5310 11133 5356
rect 11189 5310 11241 5356
rect 11297 5310 11349 5356
rect 11405 5310 11457 5356
rect 3433 5307 3485 5310
rect 3541 5307 3593 5310
rect 3649 5307 3701 5310
rect 3757 5307 3809 5310
rect 3865 5307 3917 5310
rect 3973 5307 4025 5310
rect 4081 5307 4133 5310
rect 4189 5307 4241 5310
rect 4297 5307 4349 5310
rect 4405 5307 4457 5310
rect 4513 5307 4565 5310
rect 4621 5307 4673 5310
rect 4729 5307 4781 5310
rect 4837 5307 4889 5310
rect 4945 5307 4997 5310
rect 5053 5307 5105 5310
rect 5161 5307 5213 5310
rect 6566 5307 6618 5310
rect 6674 5307 6726 5310
rect 6782 5307 6834 5310
rect 6890 5307 6942 5310
rect 6998 5307 7050 5310
rect 7106 5307 7158 5310
rect 7214 5307 7266 5310
rect 7322 5307 7374 5310
rect 7430 5307 7482 5310
rect 7538 5307 7590 5310
rect 9677 5307 9729 5310
rect 9785 5307 9837 5310
rect 9893 5307 9945 5310
rect 10001 5307 10053 5310
rect 10109 5307 10161 5310
rect 10217 5307 10269 5310
rect 10325 5307 10377 5310
rect 10433 5307 10485 5310
rect 10541 5307 10593 5310
rect 10649 5307 10701 5310
rect 10757 5307 10809 5310
rect 10865 5307 10917 5310
rect 10973 5307 11025 5310
rect 11081 5307 11133 5310
rect 11189 5307 11241 5310
rect 11297 5307 11349 5310
rect 11405 5307 11457 5310
rect 1505 5112 1557 5115
rect 1613 5112 1665 5115
rect 1721 5112 1773 5115
rect 1829 5112 1881 5115
rect 1937 5112 1989 5115
rect 2045 5112 2097 5115
rect 2153 5112 2205 5115
rect 2261 5112 2313 5115
rect 2369 5112 2421 5115
rect 2477 5112 2529 5115
rect 2585 5112 2637 5115
rect 2693 5112 2745 5115
rect 2801 5112 2853 5115
rect 2909 5112 2961 5115
rect 3017 5112 3069 5115
rect 3125 5112 3177 5115
rect 3233 5112 3285 5115
rect 5372 5112 5424 5115
rect 5480 5112 5532 5115
rect 5588 5112 5640 5115
rect 5696 5112 5748 5115
rect 5804 5112 5856 5115
rect 5912 5112 5964 5115
rect 6020 5112 6072 5115
rect 6128 5112 6180 5115
rect 6236 5112 6288 5115
rect 6344 5112 6396 5115
rect 7749 5112 7801 5115
rect 7857 5112 7909 5115
rect 7965 5112 8017 5115
rect 8073 5112 8125 5115
rect 8181 5112 8233 5115
rect 8289 5112 8341 5115
rect 8397 5112 8449 5115
rect 8505 5112 8557 5115
rect 8613 5112 8665 5115
rect 8721 5112 8773 5115
rect 8829 5112 8881 5115
rect 8937 5112 8989 5115
rect 9045 5112 9097 5115
rect 9153 5112 9205 5115
rect 9261 5112 9313 5115
rect 9369 5112 9421 5115
rect 9477 5112 9529 5115
rect 1505 5066 1557 5112
rect 1613 5066 1665 5112
rect 1721 5066 1773 5112
rect 1829 5066 1881 5112
rect 1937 5066 1989 5112
rect 2045 5066 2097 5112
rect 2153 5066 2205 5112
rect 2261 5066 2313 5112
rect 2369 5066 2421 5112
rect 2477 5066 2529 5112
rect 2585 5066 2637 5112
rect 2693 5066 2745 5112
rect 2801 5066 2853 5112
rect 2909 5066 2961 5112
rect 3017 5066 3069 5112
rect 3125 5066 3177 5112
rect 3233 5066 3285 5112
rect 5372 5066 5424 5112
rect 5480 5066 5532 5112
rect 5588 5066 5640 5112
rect 5696 5066 5748 5112
rect 5804 5066 5856 5112
rect 5912 5066 5964 5112
rect 6020 5066 6072 5112
rect 6128 5066 6180 5112
rect 6236 5066 6288 5112
rect 6344 5066 6396 5112
rect 7749 5066 7801 5112
rect 7857 5066 7909 5112
rect 7965 5066 8017 5112
rect 8073 5066 8125 5112
rect 8181 5066 8233 5112
rect 8289 5066 8341 5112
rect 8397 5066 8449 5112
rect 8505 5066 8557 5112
rect 8613 5066 8665 5112
rect 8721 5066 8773 5112
rect 8829 5066 8881 5112
rect 8937 5066 8989 5112
rect 9045 5066 9097 5112
rect 9153 5066 9205 5112
rect 9261 5066 9313 5112
rect 9369 5066 9421 5112
rect 9477 5066 9529 5112
rect 1505 5063 1557 5066
rect 1613 5063 1665 5066
rect 1721 5063 1773 5066
rect 1829 5063 1881 5066
rect 1937 5063 1989 5066
rect 2045 5063 2097 5066
rect 2153 5063 2205 5066
rect 2261 5063 2313 5066
rect 2369 5063 2421 5066
rect 2477 5063 2529 5066
rect 2585 5063 2637 5066
rect 2693 5063 2745 5066
rect 2801 5063 2853 5066
rect 2909 5063 2961 5066
rect 3017 5063 3069 5066
rect 3125 5063 3177 5066
rect 3233 5063 3285 5066
rect 5372 5063 5424 5066
rect 5480 5063 5532 5066
rect 5588 5063 5640 5066
rect 5696 5063 5748 5066
rect 5804 5063 5856 5066
rect 5912 5063 5964 5066
rect 6020 5063 6072 5066
rect 6128 5063 6180 5066
rect 6236 5063 6288 5066
rect 6344 5063 6396 5066
rect 7749 5063 7801 5066
rect 7857 5063 7909 5066
rect 7965 5063 8017 5066
rect 8073 5063 8125 5066
rect 8181 5063 8233 5066
rect 8289 5063 8341 5066
rect 8397 5063 8449 5066
rect 8505 5063 8557 5066
rect 8613 5063 8665 5066
rect 8721 5063 8773 5066
rect 8829 5063 8881 5066
rect 8937 5063 8989 5066
rect 9045 5063 9097 5066
rect 9153 5063 9205 5066
rect 9261 5063 9313 5066
rect 9369 5063 9421 5066
rect 9477 5063 9529 5066
rect 3433 4868 3485 4871
rect 3541 4868 3593 4871
rect 3649 4868 3701 4871
rect 3757 4868 3809 4871
rect 3865 4868 3917 4871
rect 3973 4868 4025 4871
rect 4081 4868 4133 4871
rect 4189 4868 4241 4871
rect 4297 4868 4349 4871
rect 4405 4868 4457 4871
rect 4513 4868 4565 4871
rect 4621 4868 4673 4871
rect 4729 4868 4781 4871
rect 4837 4868 4889 4871
rect 4945 4868 4997 4871
rect 5053 4868 5105 4871
rect 5161 4868 5213 4871
rect 6566 4868 6618 4871
rect 6674 4868 6726 4871
rect 6782 4868 6834 4871
rect 6890 4868 6942 4871
rect 6998 4868 7050 4871
rect 7106 4868 7158 4871
rect 7214 4868 7266 4871
rect 7322 4868 7374 4871
rect 7430 4868 7482 4871
rect 7538 4868 7590 4871
rect 9677 4868 9729 4871
rect 9785 4868 9837 4871
rect 9893 4868 9945 4871
rect 10001 4868 10053 4871
rect 10109 4868 10161 4871
rect 10217 4868 10269 4871
rect 10325 4868 10377 4871
rect 10433 4868 10485 4871
rect 10541 4868 10593 4871
rect 10649 4868 10701 4871
rect 10757 4868 10809 4871
rect 10865 4868 10917 4871
rect 10973 4868 11025 4871
rect 11081 4868 11133 4871
rect 11189 4868 11241 4871
rect 11297 4868 11349 4871
rect 11405 4868 11457 4871
rect 3433 4822 3485 4868
rect 3541 4822 3593 4868
rect 3649 4822 3701 4868
rect 3757 4822 3809 4868
rect 3865 4822 3917 4868
rect 3973 4822 4025 4868
rect 4081 4822 4133 4868
rect 4189 4822 4241 4868
rect 4297 4822 4349 4868
rect 4405 4822 4457 4868
rect 4513 4822 4565 4868
rect 4621 4822 4673 4868
rect 4729 4822 4781 4868
rect 4837 4822 4889 4868
rect 4945 4822 4997 4868
rect 5053 4822 5105 4868
rect 5161 4822 5213 4868
rect 6566 4822 6618 4868
rect 6674 4822 6726 4868
rect 6782 4822 6834 4868
rect 6890 4822 6942 4868
rect 6998 4822 7050 4868
rect 7106 4822 7158 4868
rect 7214 4822 7266 4868
rect 7322 4822 7374 4868
rect 7430 4822 7482 4868
rect 7538 4822 7590 4868
rect 9677 4822 9729 4868
rect 9785 4822 9837 4868
rect 9893 4822 9945 4868
rect 10001 4822 10053 4868
rect 10109 4822 10161 4868
rect 10217 4822 10269 4868
rect 10325 4822 10377 4868
rect 10433 4822 10485 4868
rect 10541 4822 10593 4868
rect 10649 4822 10701 4868
rect 10757 4822 10809 4868
rect 10865 4822 10917 4868
rect 10973 4822 11025 4868
rect 11081 4822 11133 4868
rect 11189 4822 11241 4868
rect 11297 4822 11349 4868
rect 11405 4822 11457 4868
rect 3433 4819 3485 4822
rect 3541 4819 3593 4822
rect 3649 4819 3701 4822
rect 3757 4819 3809 4822
rect 3865 4819 3917 4822
rect 3973 4819 4025 4822
rect 4081 4819 4133 4822
rect 4189 4819 4241 4822
rect 4297 4819 4349 4822
rect 4405 4819 4457 4822
rect 4513 4819 4565 4822
rect 4621 4819 4673 4822
rect 4729 4819 4781 4822
rect 4837 4819 4889 4822
rect 4945 4819 4997 4822
rect 5053 4819 5105 4822
rect 5161 4819 5213 4822
rect 6566 4819 6618 4822
rect 6674 4819 6726 4822
rect 6782 4819 6834 4822
rect 6890 4819 6942 4822
rect 6998 4819 7050 4822
rect 7106 4819 7158 4822
rect 7214 4819 7266 4822
rect 7322 4819 7374 4822
rect 7430 4819 7482 4822
rect 7538 4819 7590 4822
rect 9677 4819 9729 4822
rect 9785 4819 9837 4822
rect 9893 4819 9945 4822
rect 10001 4819 10053 4822
rect 10109 4819 10161 4822
rect 10217 4819 10269 4822
rect 10325 4819 10377 4822
rect 10433 4819 10485 4822
rect 10541 4819 10593 4822
rect 10649 4819 10701 4822
rect 10757 4819 10809 4822
rect 10865 4819 10917 4822
rect 10973 4819 11025 4822
rect 11081 4819 11133 4822
rect 11189 4819 11241 4822
rect 11297 4819 11349 4822
rect 11405 4819 11457 4822
rect 1505 4624 1557 4627
rect 1613 4624 1665 4627
rect 1721 4624 1773 4627
rect 1829 4624 1881 4627
rect 1937 4624 1989 4627
rect 2045 4624 2097 4627
rect 2153 4624 2205 4627
rect 2261 4624 2313 4627
rect 2369 4624 2421 4627
rect 2477 4624 2529 4627
rect 2585 4624 2637 4627
rect 2693 4624 2745 4627
rect 2801 4624 2853 4627
rect 2909 4624 2961 4627
rect 3017 4624 3069 4627
rect 3125 4624 3177 4627
rect 3233 4624 3285 4627
rect 5372 4624 5424 4627
rect 5480 4624 5532 4627
rect 5588 4624 5640 4627
rect 5696 4624 5748 4627
rect 5804 4624 5856 4627
rect 5912 4624 5964 4627
rect 6020 4624 6072 4627
rect 6128 4624 6180 4627
rect 6236 4624 6288 4627
rect 6344 4624 6396 4627
rect 7749 4624 7801 4627
rect 7857 4624 7909 4627
rect 7965 4624 8017 4627
rect 8073 4624 8125 4627
rect 8181 4624 8233 4627
rect 8289 4624 8341 4627
rect 8397 4624 8449 4627
rect 8505 4624 8557 4627
rect 8613 4624 8665 4627
rect 8721 4624 8773 4627
rect 8829 4624 8881 4627
rect 8937 4624 8989 4627
rect 9045 4624 9097 4627
rect 9153 4624 9205 4627
rect 9261 4624 9313 4627
rect 9369 4624 9421 4627
rect 9477 4624 9529 4627
rect 1505 4578 1557 4624
rect 1613 4578 1665 4624
rect 1721 4578 1773 4624
rect 1829 4578 1881 4624
rect 1937 4578 1989 4624
rect 2045 4578 2097 4624
rect 2153 4578 2205 4624
rect 2261 4578 2313 4624
rect 2369 4578 2421 4624
rect 2477 4578 2529 4624
rect 2585 4578 2637 4624
rect 2693 4578 2745 4624
rect 2801 4578 2853 4624
rect 2909 4578 2961 4624
rect 3017 4578 3069 4624
rect 3125 4578 3177 4624
rect 3233 4578 3285 4624
rect 5372 4578 5424 4624
rect 5480 4578 5532 4624
rect 5588 4578 5640 4624
rect 5696 4578 5748 4624
rect 5804 4578 5856 4624
rect 5912 4578 5964 4624
rect 6020 4578 6072 4624
rect 6128 4578 6180 4624
rect 6236 4578 6288 4624
rect 6344 4578 6396 4624
rect 7749 4578 7801 4624
rect 7857 4578 7909 4624
rect 7965 4578 8017 4624
rect 8073 4578 8125 4624
rect 8181 4578 8233 4624
rect 8289 4578 8341 4624
rect 8397 4578 8449 4624
rect 8505 4578 8557 4624
rect 8613 4578 8665 4624
rect 8721 4578 8773 4624
rect 8829 4578 8881 4624
rect 8937 4578 8989 4624
rect 9045 4578 9097 4624
rect 9153 4578 9205 4624
rect 9261 4578 9313 4624
rect 9369 4578 9421 4624
rect 9477 4578 9529 4624
rect 1505 4575 1557 4578
rect 1613 4575 1665 4578
rect 1721 4575 1773 4578
rect 1829 4575 1881 4578
rect 1937 4575 1989 4578
rect 2045 4575 2097 4578
rect 2153 4575 2205 4578
rect 2261 4575 2313 4578
rect 2369 4575 2421 4578
rect 2477 4575 2529 4578
rect 2585 4575 2637 4578
rect 2693 4575 2745 4578
rect 2801 4575 2853 4578
rect 2909 4575 2961 4578
rect 3017 4575 3069 4578
rect 3125 4575 3177 4578
rect 3233 4575 3285 4578
rect 5372 4575 5424 4578
rect 5480 4575 5532 4578
rect 5588 4575 5640 4578
rect 5696 4575 5748 4578
rect 5804 4575 5856 4578
rect 5912 4575 5964 4578
rect 6020 4575 6072 4578
rect 6128 4575 6180 4578
rect 6236 4575 6288 4578
rect 6344 4575 6396 4578
rect 7749 4575 7801 4578
rect 7857 4575 7909 4578
rect 7965 4575 8017 4578
rect 8073 4575 8125 4578
rect 8181 4575 8233 4578
rect 8289 4575 8341 4578
rect 8397 4575 8449 4578
rect 8505 4575 8557 4578
rect 8613 4575 8665 4578
rect 8721 4575 8773 4578
rect 8829 4575 8881 4578
rect 8937 4575 8989 4578
rect 9045 4575 9097 4578
rect 9153 4575 9205 4578
rect 9261 4575 9313 4578
rect 9369 4575 9421 4578
rect 9477 4575 9529 4578
rect 3433 4380 3485 4383
rect 3541 4380 3593 4383
rect 3649 4380 3701 4383
rect 3757 4380 3809 4383
rect 3865 4380 3917 4383
rect 3973 4380 4025 4383
rect 4081 4380 4133 4383
rect 4189 4380 4241 4383
rect 4297 4380 4349 4383
rect 4405 4380 4457 4383
rect 4513 4380 4565 4383
rect 4621 4380 4673 4383
rect 4729 4380 4781 4383
rect 4837 4380 4889 4383
rect 4945 4380 4997 4383
rect 5053 4380 5105 4383
rect 5161 4380 5213 4383
rect 6566 4380 6618 4383
rect 6674 4380 6726 4383
rect 6782 4380 6834 4383
rect 6890 4380 6942 4383
rect 6998 4380 7050 4383
rect 7106 4380 7158 4383
rect 7214 4380 7266 4383
rect 7322 4380 7374 4383
rect 7430 4380 7482 4383
rect 7538 4380 7590 4383
rect 9677 4380 9729 4383
rect 9785 4380 9837 4383
rect 9893 4380 9945 4383
rect 10001 4380 10053 4383
rect 10109 4380 10161 4383
rect 10217 4380 10269 4383
rect 10325 4380 10377 4383
rect 10433 4380 10485 4383
rect 10541 4380 10593 4383
rect 10649 4380 10701 4383
rect 10757 4380 10809 4383
rect 10865 4380 10917 4383
rect 10973 4380 11025 4383
rect 11081 4380 11133 4383
rect 11189 4380 11241 4383
rect 11297 4380 11349 4383
rect 11405 4380 11457 4383
rect 3433 4334 3485 4380
rect 3541 4334 3593 4380
rect 3649 4334 3701 4380
rect 3757 4334 3809 4380
rect 3865 4334 3917 4380
rect 3973 4334 4025 4380
rect 4081 4334 4133 4380
rect 4189 4334 4241 4380
rect 4297 4334 4349 4380
rect 4405 4334 4457 4380
rect 4513 4334 4565 4380
rect 4621 4334 4673 4380
rect 4729 4334 4781 4380
rect 4837 4334 4889 4380
rect 4945 4334 4997 4380
rect 5053 4334 5105 4380
rect 5161 4334 5213 4380
rect 6566 4334 6618 4380
rect 6674 4334 6726 4380
rect 6782 4334 6834 4380
rect 6890 4334 6942 4380
rect 6998 4334 7050 4380
rect 7106 4334 7158 4380
rect 7214 4334 7266 4380
rect 7322 4334 7374 4380
rect 7430 4334 7482 4380
rect 7538 4334 7590 4380
rect 9677 4334 9729 4380
rect 9785 4334 9837 4380
rect 9893 4334 9945 4380
rect 10001 4334 10053 4380
rect 10109 4334 10161 4380
rect 10217 4334 10269 4380
rect 10325 4334 10377 4380
rect 10433 4334 10485 4380
rect 10541 4334 10593 4380
rect 10649 4334 10701 4380
rect 10757 4334 10809 4380
rect 10865 4334 10917 4380
rect 10973 4334 11025 4380
rect 11081 4334 11133 4380
rect 11189 4334 11241 4380
rect 11297 4334 11349 4380
rect 11405 4334 11457 4380
rect 3433 4331 3485 4334
rect 3541 4331 3593 4334
rect 3649 4331 3701 4334
rect 3757 4331 3809 4334
rect 3865 4331 3917 4334
rect 3973 4331 4025 4334
rect 4081 4331 4133 4334
rect 4189 4331 4241 4334
rect 4297 4331 4349 4334
rect 4405 4331 4457 4334
rect 4513 4331 4565 4334
rect 4621 4331 4673 4334
rect 4729 4331 4781 4334
rect 4837 4331 4889 4334
rect 4945 4331 4997 4334
rect 5053 4331 5105 4334
rect 5161 4331 5213 4334
rect 6566 4331 6618 4334
rect 6674 4331 6726 4334
rect 6782 4331 6834 4334
rect 6890 4331 6942 4334
rect 6998 4331 7050 4334
rect 7106 4331 7158 4334
rect 7214 4331 7266 4334
rect 7322 4331 7374 4334
rect 7430 4331 7482 4334
rect 7538 4331 7590 4334
rect 9677 4331 9729 4334
rect 9785 4331 9837 4334
rect 9893 4331 9945 4334
rect 10001 4331 10053 4334
rect 10109 4331 10161 4334
rect 10217 4331 10269 4334
rect 10325 4331 10377 4334
rect 10433 4331 10485 4334
rect 10541 4331 10593 4334
rect 10649 4331 10701 4334
rect 10757 4331 10809 4334
rect 10865 4331 10917 4334
rect 10973 4331 11025 4334
rect 11081 4331 11133 4334
rect 11189 4331 11241 4334
rect 11297 4331 11349 4334
rect 11405 4331 11457 4334
rect 1505 4136 1557 4139
rect 1613 4136 1665 4139
rect 1721 4136 1773 4139
rect 1829 4136 1881 4139
rect 1937 4136 1989 4139
rect 2045 4136 2097 4139
rect 2153 4136 2205 4139
rect 2261 4136 2313 4139
rect 2369 4136 2421 4139
rect 2477 4136 2529 4139
rect 2585 4136 2637 4139
rect 2693 4136 2745 4139
rect 2801 4136 2853 4139
rect 2909 4136 2961 4139
rect 3017 4136 3069 4139
rect 3125 4136 3177 4139
rect 3233 4136 3285 4139
rect 5372 4136 5424 4139
rect 5480 4136 5532 4139
rect 5588 4136 5640 4139
rect 5696 4136 5748 4139
rect 5804 4136 5856 4139
rect 5912 4136 5964 4139
rect 6020 4136 6072 4139
rect 6128 4136 6180 4139
rect 6236 4136 6288 4139
rect 6344 4136 6396 4139
rect 7749 4136 7801 4139
rect 7857 4136 7909 4139
rect 7965 4136 8017 4139
rect 8073 4136 8125 4139
rect 8181 4136 8233 4139
rect 8289 4136 8341 4139
rect 8397 4136 8449 4139
rect 8505 4136 8557 4139
rect 8613 4136 8665 4139
rect 8721 4136 8773 4139
rect 8829 4136 8881 4139
rect 8937 4136 8989 4139
rect 9045 4136 9097 4139
rect 9153 4136 9205 4139
rect 9261 4136 9313 4139
rect 9369 4136 9421 4139
rect 9477 4136 9529 4139
rect 1505 4090 1557 4136
rect 1613 4090 1665 4136
rect 1721 4090 1773 4136
rect 1829 4090 1881 4136
rect 1937 4090 1989 4136
rect 2045 4090 2097 4136
rect 2153 4090 2205 4136
rect 2261 4090 2313 4136
rect 2369 4090 2421 4136
rect 2477 4090 2529 4136
rect 2585 4090 2637 4136
rect 2693 4090 2745 4136
rect 2801 4090 2853 4136
rect 2909 4090 2961 4136
rect 3017 4090 3069 4136
rect 3125 4090 3177 4136
rect 3233 4090 3285 4136
rect 5372 4090 5424 4136
rect 5480 4090 5532 4136
rect 5588 4090 5640 4136
rect 5696 4090 5748 4136
rect 5804 4090 5856 4136
rect 5912 4090 5964 4136
rect 6020 4090 6072 4136
rect 6128 4090 6180 4136
rect 6236 4090 6288 4136
rect 6344 4090 6396 4136
rect 7749 4090 7801 4136
rect 7857 4090 7909 4136
rect 7965 4090 8017 4136
rect 8073 4090 8125 4136
rect 8181 4090 8233 4136
rect 8289 4090 8341 4136
rect 8397 4090 8449 4136
rect 8505 4090 8557 4136
rect 8613 4090 8665 4136
rect 8721 4090 8773 4136
rect 8829 4090 8881 4136
rect 8937 4090 8989 4136
rect 9045 4090 9097 4136
rect 9153 4090 9205 4136
rect 9261 4090 9313 4136
rect 9369 4090 9421 4136
rect 9477 4090 9529 4136
rect 1505 4087 1557 4090
rect 1613 4087 1665 4090
rect 1721 4087 1773 4090
rect 1829 4087 1881 4090
rect 1937 4087 1989 4090
rect 2045 4087 2097 4090
rect 2153 4087 2205 4090
rect 2261 4087 2313 4090
rect 2369 4087 2421 4090
rect 2477 4087 2529 4090
rect 2585 4087 2637 4090
rect 2693 4087 2745 4090
rect 2801 4087 2853 4090
rect 2909 4087 2961 4090
rect 3017 4087 3069 4090
rect 3125 4087 3177 4090
rect 3233 4087 3285 4090
rect 5372 4087 5424 4090
rect 5480 4087 5532 4090
rect 5588 4087 5640 4090
rect 5696 4087 5748 4090
rect 5804 4087 5856 4090
rect 5912 4087 5964 4090
rect 6020 4087 6072 4090
rect 6128 4087 6180 4090
rect 6236 4087 6288 4090
rect 6344 4087 6396 4090
rect 7749 4087 7801 4090
rect 7857 4087 7909 4090
rect 7965 4087 8017 4090
rect 8073 4087 8125 4090
rect 8181 4087 8233 4090
rect 8289 4087 8341 4090
rect 8397 4087 8449 4090
rect 8505 4087 8557 4090
rect 8613 4087 8665 4090
rect 8721 4087 8773 4090
rect 8829 4087 8881 4090
rect 8937 4087 8989 4090
rect 9045 4087 9097 4090
rect 9153 4087 9205 4090
rect 9261 4087 9313 4090
rect 9369 4087 9421 4090
rect 9477 4087 9529 4090
rect 3433 3892 3485 3895
rect 3541 3892 3593 3895
rect 3649 3892 3701 3895
rect 3757 3892 3809 3895
rect 3865 3892 3917 3895
rect 3973 3892 4025 3895
rect 4081 3892 4133 3895
rect 4189 3892 4241 3895
rect 4297 3892 4349 3895
rect 4405 3892 4457 3895
rect 4513 3892 4565 3895
rect 4621 3892 4673 3895
rect 4729 3892 4781 3895
rect 4837 3892 4889 3895
rect 4945 3892 4997 3895
rect 5053 3892 5105 3895
rect 5161 3892 5213 3895
rect 6566 3892 6618 3895
rect 6674 3892 6726 3895
rect 6782 3892 6834 3895
rect 6890 3892 6942 3895
rect 6998 3892 7050 3895
rect 7106 3892 7158 3895
rect 7214 3892 7266 3895
rect 7322 3892 7374 3895
rect 7430 3892 7482 3895
rect 7538 3892 7590 3895
rect 9677 3892 9729 3895
rect 9785 3892 9837 3895
rect 9893 3892 9945 3895
rect 10001 3892 10053 3895
rect 10109 3892 10161 3895
rect 10217 3892 10269 3895
rect 10325 3892 10377 3895
rect 10433 3892 10485 3895
rect 10541 3892 10593 3895
rect 10649 3892 10701 3895
rect 10757 3892 10809 3895
rect 10865 3892 10917 3895
rect 10973 3892 11025 3895
rect 11081 3892 11133 3895
rect 11189 3892 11241 3895
rect 11297 3892 11349 3895
rect 11405 3892 11457 3895
rect 3433 3846 3485 3892
rect 3541 3846 3593 3892
rect 3649 3846 3701 3892
rect 3757 3846 3809 3892
rect 3865 3846 3917 3892
rect 3973 3846 4025 3892
rect 4081 3846 4133 3892
rect 4189 3846 4241 3892
rect 4297 3846 4349 3892
rect 4405 3846 4457 3892
rect 4513 3846 4565 3892
rect 4621 3846 4673 3892
rect 4729 3846 4781 3892
rect 4837 3846 4889 3892
rect 4945 3846 4997 3892
rect 5053 3846 5105 3892
rect 5161 3846 5213 3892
rect 6566 3846 6618 3892
rect 6674 3846 6726 3892
rect 6782 3846 6834 3892
rect 6890 3846 6942 3892
rect 6998 3846 7050 3892
rect 7106 3846 7158 3892
rect 7214 3846 7266 3892
rect 7322 3846 7374 3892
rect 7430 3846 7482 3892
rect 7538 3846 7590 3892
rect 9677 3846 9729 3892
rect 9785 3846 9837 3892
rect 9893 3846 9945 3892
rect 10001 3846 10053 3892
rect 10109 3846 10161 3892
rect 10217 3846 10269 3892
rect 10325 3846 10377 3892
rect 10433 3846 10485 3892
rect 10541 3846 10593 3892
rect 10649 3846 10701 3892
rect 10757 3846 10809 3892
rect 10865 3846 10917 3892
rect 10973 3846 11025 3892
rect 11081 3846 11133 3892
rect 11189 3846 11241 3892
rect 11297 3846 11349 3892
rect 11405 3846 11457 3892
rect 3433 3843 3485 3846
rect 3541 3843 3593 3846
rect 3649 3843 3701 3846
rect 3757 3843 3809 3846
rect 3865 3843 3917 3846
rect 3973 3843 4025 3846
rect 4081 3843 4133 3846
rect 4189 3843 4241 3846
rect 4297 3843 4349 3846
rect 4405 3843 4457 3846
rect 4513 3843 4565 3846
rect 4621 3843 4673 3846
rect 4729 3843 4781 3846
rect 4837 3843 4889 3846
rect 4945 3843 4997 3846
rect 5053 3843 5105 3846
rect 5161 3843 5213 3846
rect 6566 3843 6618 3846
rect 6674 3843 6726 3846
rect 6782 3843 6834 3846
rect 6890 3843 6942 3846
rect 6998 3843 7050 3846
rect 7106 3843 7158 3846
rect 7214 3843 7266 3846
rect 7322 3843 7374 3846
rect 7430 3843 7482 3846
rect 7538 3843 7590 3846
rect 9677 3843 9729 3846
rect 9785 3843 9837 3846
rect 9893 3843 9945 3846
rect 10001 3843 10053 3846
rect 10109 3843 10161 3846
rect 10217 3843 10269 3846
rect 10325 3843 10377 3846
rect 10433 3843 10485 3846
rect 10541 3843 10593 3846
rect 10649 3843 10701 3846
rect 10757 3843 10809 3846
rect 10865 3843 10917 3846
rect 10973 3843 11025 3846
rect 11081 3843 11133 3846
rect 11189 3843 11241 3846
rect 11297 3843 11349 3846
rect 11405 3843 11457 3846
rect 1505 3648 1557 3651
rect 1613 3648 1665 3651
rect 1721 3648 1773 3651
rect 1829 3648 1881 3651
rect 1937 3648 1989 3651
rect 2045 3648 2097 3651
rect 2153 3648 2205 3651
rect 2261 3648 2313 3651
rect 2369 3648 2421 3651
rect 2477 3648 2529 3651
rect 2585 3648 2637 3651
rect 2693 3648 2745 3651
rect 2801 3648 2853 3651
rect 2909 3648 2961 3651
rect 3017 3648 3069 3651
rect 3125 3648 3177 3651
rect 3233 3648 3285 3651
rect 5372 3648 5424 3651
rect 5480 3648 5532 3651
rect 5588 3648 5640 3651
rect 5696 3648 5748 3651
rect 5804 3648 5856 3651
rect 5912 3648 5964 3651
rect 6020 3648 6072 3651
rect 6128 3648 6180 3651
rect 6236 3648 6288 3651
rect 6344 3648 6396 3651
rect 7749 3648 7801 3651
rect 7857 3648 7909 3651
rect 7965 3648 8017 3651
rect 8073 3648 8125 3651
rect 8181 3648 8233 3651
rect 8289 3648 8341 3651
rect 8397 3648 8449 3651
rect 8505 3648 8557 3651
rect 8613 3648 8665 3651
rect 8721 3648 8773 3651
rect 8829 3648 8881 3651
rect 8937 3648 8989 3651
rect 9045 3648 9097 3651
rect 9153 3648 9205 3651
rect 9261 3648 9313 3651
rect 9369 3648 9421 3651
rect 9477 3648 9529 3651
rect 1505 3602 1557 3648
rect 1613 3602 1665 3648
rect 1721 3602 1773 3648
rect 1829 3602 1881 3648
rect 1937 3602 1989 3648
rect 2045 3602 2097 3648
rect 2153 3602 2205 3648
rect 2261 3602 2313 3648
rect 2369 3602 2421 3648
rect 2477 3602 2529 3648
rect 2585 3602 2637 3648
rect 2693 3602 2745 3648
rect 2801 3602 2853 3648
rect 2909 3602 2961 3648
rect 3017 3602 3069 3648
rect 3125 3602 3177 3648
rect 3233 3602 3285 3648
rect 5372 3602 5424 3648
rect 5480 3602 5532 3648
rect 5588 3602 5640 3648
rect 5696 3602 5748 3648
rect 5804 3602 5856 3648
rect 5912 3602 5964 3648
rect 6020 3602 6072 3648
rect 6128 3602 6180 3648
rect 6236 3602 6288 3648
rect 6344 3602 6396 3648
rect 7749 3602 7801 3648
rect 7857 3602 7909 3648
rect 7965 3602 8017 3648
rect 8073 3602 8125 3648
rect 8181 3602 8233 3648
rect 8289 3602 8341 3648
rect 8397 3602 8449 3648
rect 8505 3602 8557 3648
rect 8613 3602 8665 3648
rect 8721 3602 8773 3648
rect 8829 3602 8881 3648
rect 8937 3602 8989 3648
rect 9045 3602 9097 3648
rect 9153 3602 9205 3648
rect 9261 3602 9313 3648
rect 9369 3602 9421 3648
rect 9477 3602 9529 3648
rect 1505 3599 1557 3602
rect 1613 3599 1665 3602
rect 1721 3599 1773 3602
rect 1829 3599 1881 3602
rect 1937 3599 1989 3602
rect 2045 3599 2097 3602
rect 2153 3599 2205 3602
rect 2261 3599 2313 3602
rect 2369 3599 2421 3602
rect 2477 3599 2529 3602
rect 2585 3599 2637 3602
rect 2693 3599 2745 3602
rect 2801 3599 2853 3602
rect 2909 3599 2961 3602
rect 3017 3599 3069 3602
rect 3125 3599 3177 3602
rect 3233 3599 3285 3602
rect 5372 3599 5424 3602
rect 5480 3599 5532 3602
rect 5588 3599 5640 3602
rect 5696 3599 5748 3602
rect 5804 3599 5856 3602
rect 5912 3599 5964 3602
rect 6020 3599 6072 3602
rect 6128 3599 6180 3602
rect 6236 3599 6288 3602
rect 6344 3599 6396 3602
rect 7749 3599 7801 3602
rect 7857 3599 7909 3602
rect 7965 3599 8017 3602
rect 8073 3599 8125 3602
rect 8181 3599 8233 3602
rect 8289 3599 8341 3602
rect 8397 3599 8449 3602
rect 8505 3599 8557 3602
rect 8613 3599 8665 3602
rect 8721 3599 8773 3602
rect 8829 3599 8881 3602
rect 8937 3599 8989 3602
rect 9045 3599 9097 3602
rect 9153 3599 9205 3602
rect 9261 3599 9313 3602
rect 9369 3599 9421 3602
rect 9477 3599 9529 3602
rect 3433 3404 3485 3407
rect 3541 3404 3593 3407
rect 3649 3404 3701 3407
rect 3757 3404 3809 3407
rect 3865 3404 3917 3407
rect 3973 3404 4025 3407
rect 4081 3404 4133 3407
rect 4189 3404 4241 3407
rect 4297 3404 4349 3407
rect 4405 3404 4457 3407
rect 4513 3404 4565 3407
rect 4621 3404 4673 3407
rect 4729 3404 4781 3407
rect 4837 3404 4889 3407
rect 4945 3404 4997 3407
rect 5053 3404 5105 3407
rect 5161 3404 5213 3407
rect 6566 3404 6618 3407
rect 6674 3404 6726 3407
rect 6782 3404 6834 3407
rect 6890 3404 6942 3407
rect 6998 3404 7050 3407
rect 7106 3404 7158 3407
rect 7214 3404 7266 3407
rect 7322 3404 7374 3407
rect 7430 3404 7482 3407
rect 7538 3404 7590 3407
rect 9677 3404 9729 3407
rect 9785 3404 9837 3407
rect 9893 3404 9945 3407
rect 10001 3404 10053 3407
rect 10109 3404 10161 3407
rect 10217 3404 10269 3407
rect 10325 3404 10377 3407
rect 10433 3404 10485 3407
rect 10541 3404 10593 3407
rect 10649 3404 10701 3407
rect 10757 3404 10809 3407
rect 10865 3404 10917 3407
rect 10973 3404 11025 3407
rect 11081 3404 11133 3407
rect 11189 3404 11241 3407
rect 11297 3404 11349 3407
rect 11405 3404 11457 3407
rect 3433 3358 3485 3404
rect 3541 3358 3593 3404
rect 3649 3358 3701 3404
rect 3757 3358 3809 3404
rect 3865 3358 3917 3404
rect 3973 3358 4025 3404
rect 4081 3358 4133 3404
rect 4189 3358 4241 3404
rect 4297 3358 4349 3404
rect 4405 3358 4457 3404
rect 4513 3358 4565 3404
rect 4621 3358 4673 3404
rect 4729 3358 4781 3404
rect 4837 3358 4889 3404
rect 4945 3358 4997 3404
rect 5053 3358 5105 3404
rect 5161 3358 5213 3404
rect 6566 3358 6618 3404
rect 6674 3358 6726 3404
rect 6782 3358 6834 3404
rect 6890 3358 6942 3404
rect 6998 3358 7050 3404
rect 7106 3358 7158 3404
rect 7214 3358 7266 3404
rect 7322 3358 7374 3404
rect 7430 3358 7482 3404
rect 7538 3358 7590 3404
rect 9677 3358 9729 3404
rect 9785 3358 9837 3404
rect 9893 3358 9945 3404
rect 10001 3358 10053 3404
rect 10109 3358 10161 3404
rect 10217 3358 10269 3404
rect 10325 3358 10377 3404
rect 10433 3358 10485 3404
rect 10541 3358 10593 3404
rect 10649 3358 10701 3404
rect 10757 3358 10809 3404
rect 10865 3358 10917 3404
rect 10973 3358 11025 3404
rect 11081 3358 11133 3404
rect 11189 3358 11241 3404
rect 11297 3358 11349 3404
rect 11405 3358 11457 3404
rect 3433 3355 3485 3358
rect 3541 3355 3593 3358
rect 3649 3355 3701 3358
rect 3757 3355 3809 3358
rect 3865 3355 3917 3358
rect 3973 3355 4025 3358
rect 4081 3355 4133 3358
rect 4189 3355 4241 3358
rect 4297 3355 4349 3358
rect 4405 3355 4457 3358
rect 4513 3355 4565 3358
rect 4621 3355 4673 3358
rect 4729 3355 4781 3358
rect 4837 3355 4889 3358
rect 4945 3355 4997 3358
rect 5053 3355 5105 3358
rect 5161 3355 5213 3358
rect 6566 3355 6618 3358
rect 6674 3355 6726 3358
rect 6782 3355 6834 3358
rect 6890 3355 6942 3358
rect 6998 3355 7050 3358
rect 7106 3355 7158 3358
rect 7214 3355 7266 3358
rect 7322 3355 7374 3358
rect 7430 3355 7482 3358
rect 7538 3355 7590 3358
rect 9677 3355 9729 3358
rect 9785 3355 9837 3358
rect 9893 3355 9945 3358
rect 10001 3355 10053 3358
rect 10109 3355 10161 3358
rect 10217 3355 10269 3358
rect 10325 3355 10377 3358
rect 10433 3355 10485 3358
rect 10541 3355 10593 3358
rect 10649 3355 10701 3358
rect 10757 3355 10809 3358
rect 10865 3355 10917 3358
rect 10973 3355 11025 3358
rect 11081 3355 11133 3358
rect 11189 3355 11241 3358
rect 11297 3355 11349 3358
rect 11405 3355 11457 3358
rect 1505 3160 1557 3163
rect 1613 3160 1665 3163
rect 1721 3160 1773 3163
rect 1829 3160 1881 3163
rect 1937 3160 1989 3163
rect 2045 3160 2097 3163
rect 2153 3160 2205 3163
rect 2261 3160 2313 3163
rect 2369 3160 2421 3163
rect 2477 3160 2529 3163
rect 2585 3160 2637 3163
rect 2693 3160 2745 3163
rect 2801 3160 2853 3163
rect 2909 3160 2961 3163
rect 3017 3160 3069 3163
rect 3125 3160 3177 3163
rect 3233 3160 3285 3163
rect 5372 3160 5424 3163
rect 5480 3160 5532 3163
rect 5588 3160 5640 3163
rect 5696 3160 5748 3163
rect 5804 3160 5856 3163
rect 5912 3160 5964 3163
rect 6020 3160 6072 3163
rect 6128 3160 6180 3163
rect 6236 3160 6288 3163
rect 6344 3160 6396 3163
rect 7749 3160 7801 3163
rect 7857 3160 7909 3163
rect 7965 3160 8017 3163
rect 8073 3160 8125 3163
rect 8181 3160 8233 3163
rect 8289 3160 8341 3163
rect 8397 3160 8449 3163
rect 8505 3160 8557 3163
rect 8613 3160 8665 3163
rect 8721 3160 8773 3163
rect 8829 3160 8881 3163
rect 8937 3160 8989 3163
rect 9045 3160 9097 3163
rect 9153 3160 9205 3163
rect 9261 3160 9313 3163
rect 9369 3160 9421 3163
rect 9477 3160 9529 3163
rect 1505 3114 1557 3160
rect 1613 3114 1665 3160
rect 1721 3114 1773 3160
rect 1829 3114 1881 3160
rect 1937 3114 1989 3160
rect 2045 3114 2097 3160
rect 2153 3114 2205 3160
rect 2261 3114 2313 3160
rect 2369 3114 2421 3160
rect 2477 3114 2529 3160
rect 2585 3114 2637 3160
rect 2693 3114 2745 3160
rect 2801 3114 2853 3160
rect 2909 3114 2961 3160
rect 3017 3114 3069 3160
rect 3125 3114 3177 3160
rect 3233 3114 3285 3160
rect 5372 3114 5424 3160
rect 5480 3114 5532 3160
rect 5588 3114 5640 3160
rect 5696 3114 5748 3160
rect 5804 3114 5856 3160
rect 5912 3114 5964 3160
rect 6020 3114 6072 3160
rect 6128 3114 6180 3160
rect 6236 3114 6288 3160
rect 6344 3114 6396 3160
rect 7749 3114 7801 3160
rect 7857 3114 7909 3160
rect 7965 3114 8017 3160
rect 8073 3114 8125 3160
rect 8181 3114 8233 3160
rect 8289 3114 8341 3160
rect 8397 3114 8449 3160
rect 8505 3114 8557 3160
rect 8613 3114 8665 3160
rect 8721 3114 8773 3160
rect 8829 3114 8881 3160
rect 8937 3114 8989 3160
rect 9045 3114 9097 3160
rect 9153 3114 9205 3160
rect 9261 3114 9313 3160
rect 9369 3114 9421 3160
rect 9477 3114 9529 3160
rect 1505 3111 1557 3114
rect 1613 3111 1665 3114
rect 1721 3111 1773 3114
rect 1829 3111 1881 3114
rect 1937 3111 1989 3114
rect 2045 3111 2097 3114
rect 2153 3111 2205 3114
rect 2261 3111 2313 3114
rect 2369 3111 2421 3114
rect 2477 3111 2529 3114
rect 2585 3111 2637 3114
rect 2693 3111 2745 3114
rect 2801 3111 2853 3114
rect 2909 3111 2961 3114
rect 3017 3111 3069 3114
rect 3125 3111 3177 3114
rect 3233 3111 3285 3114
rect 5372 3111 5424 3114
rect 5480 3111 5532 3114
rect 5588 3111 5640 3114
rect 5696 3111 5748 3114
rect 5804 3111 5856 3114
rect 5912 3111 5964 3114
rect 6020 3111 6072 3114
rect 6128 3111 6180 3114
rect 6236 3111 6288 3114
rect 6344 3111 6396 3114
rect 7749 3111 7801 3114
rect 7857 3111 7909 3114
rect 7965 3111 8017 3114
rect 8073 3111 8125 3114
rect 8181 3111 8233 3114
rect 8289 3111 8341 3114
rect 8397 3111 8449 3114
rect 8505 3111 8557 3114
rect 8613 3111 8665 3114
rect 8721 3111 8773 3114
rect 8829 3111 8881 3114
rect 8937 3111 8989 3114
rect 9045 3111 9097 3114
rect 9153 3111 9205 3114
rect 9261 3111 9313 3114
rect 9369 3111 9421 3114
rect 9477 3111 9529 3114
rect 3433 2916 3485 2919
rect 3541 2916 3593 2919
rect 3649 2916 3701 2919
rect 3757 2916 3809 2919
rect 3865 2916 3917 2919
rect 3973 2916 4025 2919
rect 4081 2916 4133 2919
rect 4189 2916 4241 2919
rect 4297 2916 4349 2919
rect 4405 2916 4457 2919
rect 4513 2916 4565 2919
rect 4621 2916 4673 2919
rect 4729 2916 4781 2919
rect 4837 2916 4889 2919
rect 4945 2916 4997 2919
rect 5053 2916 5105 2919
rect 5161 2916 5213 2919
rect 6566 2916 6618 2919
rect 6674 2916 6726 2919
rect 6782 2916 6834 2919
rect 6890 2916 6942 2919
rect 6998 2916 7050 2919
rect 7106 2916 7158 2919
rect 7214 2916 7266 2919
rect 7322 2916 7374 2919
rect 7430 2916 7482 2919
rect 7538 2916 7590 2919
rect 9677 2916 9729 2919
rect 9785 2916 9837 2919
rect 9893 2916 9945 2919
rect 10001 2916 10053 2919
rect 10109 2916 10161 2919
rect 10217 2916 10269 2919
rect 10325 2916 10377 2919
rect 10433 2916 10485 2919
rect 10541 2916 10593 2919
rect 10649 2916 10701 2919
rect 10757 2916 10809 2919
rect 10865 2916 10917 2919
rect 10973 2916 11025 2919
rect 11081 2916 11133 2919
rect 11189 2916 11241 2919
rect 11297 2916 11349 2919
rect 11405 2916 11457 2919
rect 3433 2870 3485 2916
rect 3541 2870 3593 2916
rect 3649 2870 3701 2916
rect 3757 2870 3809 2916
rect 3865 2870 3917 2916
rect 3973 2870 4025 2916
rect 4081 2870 4133 2916
rect 4189 2870 4241 2916
rect 4297 2870 4349 2916
rect 4405 2870 4457 2916
rect 4513 2870 4565 2916
rect 4621 2870 4673 2916
rect 4729 2870 4781 2916
rect 4837 2870 4889 2916
rect 4945 2870 4997 2916
rect 5053 2870 5105 2916
rect 5161 2870 5213 2916
rect 6566 2870 6618 2916
rect 6674 2870 6726 2916
rect 6782 2870 6834 2916
rect 6890 2870 6942 2916
rect 6998 2870 7050 2916
rect 7106 2870 7158 2916
rect 7214 2870 7266 2916
rect 7322 2870 7374 2916
rect 7430 2870 7482 2916
rect 7538 2870 7590 2916
rect 9677 2870 9729 2916
rect 9785 2870 9837 2916
rect 9893 2870 9945 2916
rect 10001 2870 10053 2916
rect 10109 2870 10161 2916
rect 10217 2870 10269 2916
rect 10325 2870 10377 2916
rect 10433 2870 10485 2916
rect 10541 2870 10593 2916
rect 10649 2870 10701 2916
rect 10757 2870 10809 2916
rect 10865 2870 10917 2916
rect 10973 2870 11025 2916
rect 11081 2870 11133 2916
rect 11189 2870 11241 2916
rect 11297 2870 11349 2916
rect 11405 2870 11457 2916
rect 3433 2867 3485 2870
rect 3541 2867 3593 2870
rect 3649 2867 3701 2870
rect 3757 2867 3809 2870
rect 3865 2867 3917 2870
rect 3973 2867 4025 2870
rect 4081 2867 4133 2870
rect 4189 2867 4241 2870
rect 4297 2867 4349 2870
rect 4405 2867 4457 2870
rect 4513 2867 4565 2870
rect 4621 2867 4673 2870
rect 4729 2867 4781 2870
rect 4837 2867 4889 2870
rect 4945 2867 4997 2870
rect 5053 2867 5105 2870
rect 5161 2867 5213 2870
rect 6566 2867 6618 2870
rect 6674 2867 6726 2870
rect 6782 2867 6834 2870
rect 6890 2867 6942 2870
rect 6998 2867 7050 2870
rect 7106 2867 7158 2870
rect 7214 2867 7266 2870
rect 7322 2867 7374 2870
rect 7430 2867 7482 2870
rect 7538 2867 7590 2870
rect 9677 2867 9729 2870
rect 9785 2867 9837 2870
rect 9893 2867 9945 2870
rect 10001 2867 10053 2870
rect 10109 2867 10161 2870
rect 10217 2867 10269 2870
rect 10325 2867 10377 2870
rect 10433 2867 10485 2870
rect 10541 2867 10593 2870
rect 10649 2867 10701 2870
rect 10757 2867 10809 2870
rect 10865 2867 10917 2870
rect 10973 2867 11025 2870
rect 11081 2867 11133 2870
rect 11189 2867 11241 2870
rect 11297 2867 11349 2870
rect 11405 2867 11457 2870
rect 1505 2672 1557 2675
rect 1613 2672 1665 2675
rect 1721 2672 1773 2675
rect 1829 2672 1881 2675
rect 1937 2672 1989 2675
rect 2045 2672 2097 2675
rect 2153 2672 2205 2675
rect 2261 2672 2313 2675
rect 2369 2672 2421 2675
rect 2477 2672 2529 2675
rect 2585 2672 2637 2675
rect 2693 2672 2745 2675
rect 2801 2672 2853 2675
rect 2909 2672 2961 2675
rect 3017 2672 3069 2675
rect 3125 2672 3177 2675
rect 3233 2672 3285 2675
rect 5372 2672 5424 2675
rect 5480 2672 5532 2675
rect 5588 2672 5640 2675
rect 5696 2672 5748 2675
rect 5804 2672 5856 2675
rect 5912 2672 5964 2675
rect 6020 2672 6072 2675
rect 6128 2672 6180 2675
rect 6236 2672 6288 2675
rect 6344 2672 6396 2675
rect 7749 2672 7801 2675
rect 7857 2672 7909 2675
rect 7965 2672 8017 2675
rect 8073 2672 8125 2675
rect 8181 2672 8233 2675
rect 8289 2672 8341 2675
rect 8397 2672 8449 2675
rect 8505 2672 8557 2675
rect 8613 2672 8665 2675
rect 8721 2672 8773 2675
rect 8829 2672 8881 2675
rect 8937 2672 8989 2675
rect 9045 2672 9097 2675
rect 9153 2672 9205 2675
rect 9261 2672 9313 2675
rect 9369 2672 9421 2675
rect 9477 2672 9529 2675
rect 1505 2626 1557 2672
rect 1613 2626 1665 2672
rect 1721 2626 1773 2672
rect 1829 2626 1881 2672
rect 1937 2626 1989 2672
rect 2045 2626 2097 2672
rect 2153 2626 2205 2672
rect 2261 2626 2313 2672
rect 2369 2626 2421 2672
rect 2477 2626 2529 2672
rect 2585 2626 2637 2672
rect 2693 2626 2745 2672
rect 2801 2626 2853 2672
rect 2909 2626 2961 2672
rect 3017 2626 3069 2672
rect 3125 2626 3177 2672
rect 3233 2626 3285 2672
rect 5372 2626 5424 2672
rect 5480 2626 5532 2672
rect 5588 2626 5640 2672
rect 5696 2626 5748 2672
rect 5804 2626 5856 2672
rect 5912 2626 5964 2672
rect 6020 2626 6072 2672
rect 6128 2626 6180 2672
rect 6236 2626 6288 2672
rect 6344 2626 6396 2672
rect 7749 2626 7801 2672
rect 7857 2626 7909 2672
rect 7965 2626 8017 2672
rect 8073 2626 8125 2672
rect 8181 2626 8233 2672
rect 8289 2626 8341 2672
rect 8397 2626 8449 2672
rect 8505 2626 8557 2672
rect 8613 2626 8665 2672
rect 8721 2626 8773 2672
rect 8829 2626 8881 2672
rect 8937 2626 8989 2672
rect 9045 2626 9097 2672
rect 9153 2626 9205 2672
rect 9261 2626 9313 2672
rect 9369 2626 9421 2672
rect 9477 2626 9529 2672
rect 1505 2623 1557 2626
rect 1613 2623 1665 2626
rect 1721 2623 1773 2626
rect 1829 2623 1881 2626
rect 1937 2623 1989 2626
rect 2045 2623 2097 2626
rect 2153 2623 2205 2626
rect 2261 2623 2313 2626
rect 2369 2623 2421 2626
rect 2477 2623 2529 2626
rect 2585 2623 2637 2626
rect 2693 2623 2745 2626
rect 2801 2623 2853 2626
rect 2909 2623 2961 2626
rect 3017 2623 3069 2626
rect 3125 2623 3177 2626
rect 3233 2623 3285 2626
rect 5372 2623 5424 2626
rect 5480 2623 5532 2626
rect 5588 2623 5640 2626
rect 5696 2623 5748 2626
rect 5804 2623 5856 2626
rect 5912 2623 5964 2626
rect 6020 2623 6072 2626
rect 6128 2623 6180 2626
rect 6236 2623 6288 2626
rect 6344 2623 6396 2626
rect 7749 2623 7801 2626
rect 7857 2623 7909 2626
rect 7965 2623 8017 2626
rect 8073 2623 8125 2626
rect 8181 2623 8233 2626
rect 8289 2623 8341 2626
rect 8397 2623 8449 2626
rect 8505 2623 8557 2626
rect 8613 2623 8665 2626
rect 8721 2623 8773 2626
rect 8829 2623 8881 2626
rect 8937 2623 8989 2626
rect 9045 2623 9097 2626
rect 9153 2623 9205 2626
rect 9261 2623 9313 2626
rect 9369 2623 9421 2626
rect 9477 2623 9529 2626
rect 3433 2428 3485 2431
rect 3541 2428 3593 2431
rect 3649 2428 3701 2431
rect 3757 2428 3809 2431
rect 3865 2428 3917 2431
rect 3973 2428 4025 2431
rect 4081 2428 4133 2431
rect 4189 2428 4241 2431
rect 4297 2428 4349 2431
rect 4405 2428 4457 2431
rect 4513 2428 4565 2431
rect 4621 2428 4673 2431
rect 4729 2428 4781 2431
rect 4837 2428 4889 2431
rect 4945 2428 4997 2431
rect 5053 2428 5105 2431
rect 5161 2428 5213 2431
rect 6566 2428 6618 2431
rect 6674 2428 6726 2431
rect 6782 2428 6834 2431
rect 6890 2428 6942 2431
rect 6998 2428 7050 2431
rect 7106 2428 7158 2431
rect 7214 2428 7266 2431
rect 7322 2428 7374 2431
rect 7430 2428 7482 2431
rect 7538 2428 7590 2431
rect 9677 2428 9729 2431
rect 9785 2428 9837 2431
rect 9893 2428 9945 2431
rect 10001 2428 10053 2431
rect 10109 2428 10161 2431
rect 10217 2428 10269 2431
rect 10325 2428 10377 2431
rect 10433 2428 10485 2431
rect 10541 2428 10593 2431
rect 10649 2428 10701 2431
rect 10757 2428 10809 2431
rect 10865 2428 10917 2431
rect 10973 2428 11025 2431
rect 11081 2428 11133 2431
rect 11189 2428 11241 2431
rect 11297 2428 11349 2431
rect 11405 2428 11457 2431
rect 3433 2382 3485 2428
rect 3541 2382 3593 2428
rect 3649 2382 3701 2428
rect 3757 2382 3809 2428
rect 3865 2382 3917 2428
rect 3973 2382 4025 2428
rect 4081 2382 4133 2428
rect 4189 2382 4241 2428
rect 4297 2382 4349 2428
rect 4405 2382 4457 2428
rect 4513 2382 4565 2428
rect 4621 2382 4673 2428
rect 4729 2382 4781 2428
rect 4837 2382 4889 2428
rect 4945 2382 4997 2428
rect 5053 2382 5105 2428
rect 5161 2382 5213 2428
rect 6566 2382 6618 2428
rect 6674 2382 6726 2428
rect 6782 2382 6834 2428
rect 6890 2382 6942 2428
rect 6998 2382 7050 2428
rect 7106 2382 7158 2428
rect 7214 2382 7266 2428
rect 7322 2382 7374 2428
rect 7430 2382 7482 2428
rect 7538 2382 7590 2428
rect 9677 2382 9729 2428
rect 9785 2382 9837 2428
rect 9893 2382 9945 2428
rect 10001 2382 10053 2428
rect 10109 2382 10161 2428
rect 10217 2382 10269 2428
rect 10325 2382 10377 2428
rect 10433 2382 10485 2428
rect 10541 2382 10593 2428
rect 10649 2382 10701 2428
rect 10757 2382 10809 2428
rect 10865 2382 10917 2428
rect 10973 2382 11025 2428
rect 11081 2382 11133 2428
rect 11189 2382 11241 2428
rect 11297 2382 11349 2428
rect 11405 2382 11457 2428
rect 3433 2379 3485 2382
rect 3541 2379 3593 2382
rect 3649 2379 3701 2382
rect 3757 2379 3809 2382
rect 3865 2379 3917 2382
rect 3973 2379 4025 2382
rect 4081 2379 4133 2382
rect 4189 2379 4241 2382
rect 4297 2379 4349 2382
rect 4405 2379 4457 2382
rect 4513 2379 4565 2382
rect 4621 2379 4673 2382
rect 4729 2379 4781 2382
rect 4837 2379 4889 2382
rect 4945 2379 4997 2382
rect 5053 2379 5105 2382
rect 5161 2379 5213 2382
rect 6566 2379 6618 2382
rect 6674 2379 6726 2382
rect 6782 2379 6834 2382
rect 6890 2379 6942 2382
rect 6998 2379 7050 2382
rect 7106 2379 7158 2382
rect 7214 2379 7266 2382
rect 7322 2379 7374 2382
rect 7430 2379 7482 2382
rect 7538 2379 7590 2382
rect 9677 2379 9729 2382
rect 9785 2379 9837 2382
rect 9893 2379 9945 2382
rect 10001 2379 10053 2382
rect 10109 2379 10161 2382
rect 10217 2379 10269 2382
rect 10325 2379 10377 2382
rect 10433 2379 10485 2382
rect 10541 2379 10593 2382
rect 10649 2379 10701 2382
rect 10757 2379 10809 2382
rect 10865 2379 10917 2382
rect 10973 2379 11025 2382
rect 11081 2379 11133 2382
rect 11189 2379 11241 2382
rect 11297 2379 11349 2382
rect 11405 2379 11457 2382
rect 1505 2184 1557 2187
rect 1613 2184 1665 2187
rect 1721 2184 1773 2187
rect 1829 2184 1881 2187
rect 1937 2184 1989 2187
rect 2045 2184 2097 2187
rect 2153 2184 2205 2187
rect 2261 2184 2313 2187
rect 2369 2184 2421 2187
rect 2477 2184 2529 2187
rect 2585 2184 2637 2187
rect 2693 2184 2745 2187
rect 2801 2184 2853 2187
rect 2909 2184 2961 2187
rect 3017 2184 3069 2187
rect 3125 2184 3177 2187
rect 3233 2184 3285 2187
rect 5372 2184 5424 2187
rect 5480 2184 5532 2187
rect 5588 2184 5640 2187
rect 5696 2184 5748 2187
rect 5804 2184 5856 2187
rect 5912 2184 5964 2187
rect 6020 2184 6072 2187
rect 6128 2184 6180 2187
rect 6236 2184 6288 2187
rect 6344 2184 6396 2187
rect 7749 2184 7801 2187
rect 7857 2184 7909 2187
rect 7965 2184 8017 2187
rect 8073 2184 8125 2187
rect 8181 2184 8233 2187
rect 8289 2184 8341 2187
rect 8397 2184 8449 2187
rect 8505 2184 8557 2187
rect 8613 2184 8665 2187
rect 8721 2184 8773 2187
rect 8829 2184 8881 2187
rect 8937 2184 8989 2187
rect 9045 2184 9097 2187
rect 9153 2184 9205 2187
rect 9261 2184 9313 2187
rect 9369 2184 9421 2187
rect 9477 2184 9529 2187
rect 1505 2138 1557 2184
rect 1613 2138 1665 2184
rect 1721 2138 1773 2184
rect 1829 2138 1881 2184
rect 1937 2138 1989 2184
rect 2045 2138 2097 2184
rect 2153 2138 2205 2184
rect 2261 2138 2313 2184
rect 2369 2138 2421 2184
rect 2477 2138 2529 2184
rect 2585 2138 2637 2184
rect 2693 2138 2745 2184
rect 2801 2138 2853 2184
rect 2909 2138 2961 2184
rect 3017 2138 3069 2184
rect 3125 2138 3177 2184
rect 3233 2138 3285 2184
rect 5372 2138 5424 2184
rect 5480 2138 5532 2184
rect 5588 2138 5640 2184
rect 5696 2138 5748 2184
rect 5804 2138 5856 2184
rect 5912 2138 5964 2184
rect 6020 2138 6072 2184
rect 6128 2138 6180 2184
rect 6236 2138 6288 2184
rect 6344 2138 6396 2184
rect 7749 2138 7801 2184
rect 7857 2138 7909 2184
rect 7965 2138 8017 2184
rect 8073 2138 8125 2184
rect 8181 2138 8233 2184
rect 8289 2138 8341 2184
rect 8397 2138 8449 2184
rect 8505 2138 8557 2184
rect 8613 2138 8665 2184
rect 8721 2138 8773 2184
rect 8829 2138 8881 2184
rect 8937 2138 8989 2184
rect 9045 2138 9097 2184
rect 9153 2138 9205 2184
rect 9261 2138 9313 2184
rect 9369 2138 9421 2184
rect 9477 2138 9529 2184
rect 1505 2135 1557 2138
rect 1613 2135 1665 2138
rect 1721 2135 1773 2138
rect 1829 2135 1881 2138
rect 1937 2135 1989 2138
rect 2045 2135 2097 2138
rect 2153 2135 2205 2138
rect 2261 2135 2313 2138
rect 2369 2135 2421 2138
rect 2477 2135 2529 2138
rect 2585 2135 2637 2138
rect 2693 2135 2745 2138
rect 2801 2135 2853 2138
rect 2909 2135 2961 2138
rect 3017 2135 3069 2138
rect 3125 2135 3177 2138
rect 3233 2135 3285 2138
rect 5372 2135 5424 2138
rect 5480 2135 5532 2138
rect 5588 2135 5640 2138
rect 5696 2135 5748 2138
rect 5804 2135 5856 2138
rect 5912 2135 5964 2138
rect 6020 2135 6072 2138
rect 6128 2135 6180 2138
rect 6236 2135 6288 2138
rect 6344 2135 6396 2138
rect 7749 2135 7801 2138
rect 7857 2135 7909 2138
rect 7965 2135 8017 2138
rect 8073 2135 8125 2138
rect 8181 2135 8233 2138
rect 8289 2135 8341 2138
rect 8397 2135 8449 2138
rect 8505 2135 8557 2138
rect 8613 2135 8665 2138
rect 8721 2135 8773 2138
rect 8829 2135 8881 2138
rect 8937 2135 8989 2138
rect 9045 2135 9097 2138
rect 9153 2135 9205 2138
rect 9261 2135 9313 2138
rect 9369 2135 9421 2138
rect 9477 2135 9529 2138
rect 3433 1940 3485 1943
rect 3541 1940 3593 1943
rect 3649 1940 3701 1943
rect 3757 1940 3809 1943
rect 3865 1940 3917 1943
rect 3973 1940 4025 1943
rect 4081 1940 4133 1943
rect 4189 1940 4241 1943
rect 4297 1940 4349 1943
rect 4405 1940 4457 1943
rect 4513 1940 4565 1943
rect 4621 1940 4673 1943
rect 4729 1940 4781 1943
rect 4837 1940 4889 1943
rect 4945 1940 4997 1943
rect 5053 1940 5105 1943
rect 5161 1940 5213 1943
rect 6566 1940 6618 1943
rect 6674 1940 6726 1943
rect 6782 1940 6834 1943
rect 6890 1940 6942 1943
rect 6998 1940 7050 1943
rect 7106 1940 7158 1943
rect 7214 1940 7266 1943
rect 7322 1940 7374 1943
rect 7430 1940 7482 1943
rect 7538 1940 7590 1943
rect 9677 1940 9729 1943
rect 9785 1940 9837 1943
rect 9893 1940 9945 1943
rect 10001 1940 10053 1943
rect 10109 1940 10161 1943
rect 10217 1940 10269 1943
rect 10325 1940 10377 1943
rect 10433 1940 10485 1943
rect 10541 1940 10593 1943
rect 10649 1940 10701 1943
rect 10757 1940 10809 1943
rect 10865 1940 10917 1943
rect 10973 1940 11025 1943
rect 11081 1940 11133 1943
rect 11189 1940 11241 1943
rect 11297 1940 11349 1943
rect 11405 1940 11457 1943
rect 3433 1894 3485 1940
rect 3541 1894 3593 1940
rect 3649 1894 3701 1940
rect 3757 1894 3809 1940
rect 3865 1894 3917 1940
rect 3973 1894 4025 1940
rect 4081 1894 4133 1940
rect 4189 1894 4241 1940
rect 4297 1894 4349 1940
rect 4405 1894 4457 1940
rect 4513 1894 4565 1940
rect 4621 1894 4673 1940
rect 4729 1894 4781 1940
rect 4837 1894 4889 1940
rect 4945 1894 4997 1940
rect 5053 1894 5105 1940
rect 5161 1894 5213 1940
rect 6566 1894 6618 1940
rect 6674 1894 6726 1940
rect 6782 1894 6834 1940
rect 6890 1894 6942 1940
rect 6998 1894 7050 1940
rect 7106 1894 7158 1940
rect 7214 1894 7266 1940
rect 7322 1894 7374 1940
rect 7430 1894 7482 1940
rect 7538 1894 7590 1940
rect 9677 1894 9729 1940
rect 9785 1894 9837 1940
rect 9893 1894 9945 1940
rect 10001 1894 10053 1940
rect 10109 1894 10161 1940
rect 10217 1894 10269 1940
rect 10325 1894 10377 1940
rect 10433 1894 10485 1940
rect 10541 1894 10593 1940
rect 10649 1894 10701 1940
rect 10757 1894 10809 1940
rect 10865 1894 10917 1940
rect 10973 1894 11025 1940
rect 11081 1894 11133 1940
rect 11189 1894 11241 1940
rect 11297 1894 11349 1940
rect 11405 1894 11457 1940
rect 3433 1891 3485 1894
rect 3541 1891 3593 1894
rect 3649 1891 3701 1894
rect 3757 1891 3809 1894
rect 3865 1891 3917 1894
rect 3973 1891 4025 1894
rect 4081 1891 4133 1894
rect 4189 1891 4241 1894
rect 4297 1891 4349 1894
rect 4405 1891 4457 1894
rect 4513 1891 4565 1894
rect 4621 1891 4673 1894
rect 4729 1891 4781 1894
rect 4837 1891 4889 1894
rect 4945 1891 4997 1894
rect 5053 1891 5105 1894
rect 5161 1891 5213 1894
rect 6566 1891 6618 1894
rect 6674 1891 6726 1894
rect 6782 1891 6834 1894
rect 6890 1891 6942 1894
rect 6998 1891 7050 1894
rect 7106 1891 7158 1894
rect 7214 1891 7266 1894
rect 7322 1891 7374 1894
rect 7430 1891 7482 1894
rect 7538 1891 7590 1894
rect 9677 1891 9729 1894
rect 9785 1891 9837 1894
rect 9893 1891 9945 1894
rect 10001 1891 10053 1894
rect 10109 1891 10161 1894
rect 10217 1891 10269 1894
rect 10325 1891 10377 1894
rect 10433 1891 10485 1894
rect 10541 1891 10593 1894
rect 10649 1891 10701 1894
rect 10757 1891 10809 1894
rect 10865 1891 10917 1894
rect 10973 1891 11025 1894
rect 11081 1891 11133 1894
rect 11189 1891 11241 1894
rect 11297 1891 11349 1894
rect 11405 1891 11457 1894
rect 1505 1696 1557 1699
rect 1613 1696 1665 1699
rect 1721 1696 1773 1699
rect 1829 1696 1881 1699
rect 1937 1696 1989 1699
rect 2045 1696 2097 1699
rect 2153 1696 2205 1699
rect 2261 1696 2313 1699
rect 2369 1696 2421 1699
rect 2477 1696 2529 1699
rect 2585 1696 2637 1699
rect 2693 1696 2745 1699
rect 2801 1696 2853 1699
rect 2909 1696 2961 1699
rect 3017 1696 3069 1699
rect 3125 1696 3177 1699
rect 3233 1696 3285 1699
rect 5372 1696 5424 1699
rect 5480 1696 5532 1699
rect 5588 1696 5640 1699
rect 5696 1696 5748 1699
rect 5804 1696 5856 1699
rect 5912 1696 5964 1699
rect 6020 1696 6072 1699
rect 6128 1696 6180 1699
rect 6236 1696 6288 1699
rect 6344 1696 6396 1699
rect 7749 1696 7801 1699
rect 7857 1696 7909 1699
rect 7965 1696 8017 1699
rect 8073 1696 8125 1699
rect 8181 1696 8233 1699
rect 8289 1696 8341 1699
rect 8397 1696 8449 1699
rect 8505 1696 8557 1699
rect 8613 1696 8665 1699
rect 8721 1696 8773 1699
rect 8829 1696 8881 1699
rect 8937 1696 8989 1699
rect 9045 1696 9097 1699
rect 9153 1696 9205 1699
rect 9261 1696 9313 1699
rect 9369 1696 9421 1699
rect 9477 1696 9529 1699
rect 1505 1650 1557 1696
rect 1613 1650 1665 1696
rect 1721 1650 1773 1696
rect 1829 1650 1881 1696
rect 1937 1650 1989 1696
rect 2045 1650 2097 1696
rect 2153 1650 2205 1696
rect 2261 1650 2313 1696
rect 2369 1650 2421 1696
rect 2477 1650 2529 1696
rect 2585 1650 2637 1696
rect 2693 1650 2745 1696
rect 2801 1650 2853 1696
rect 2909 1650 2961 1696
rect 3017 1650 3069 1696
rect 3125 1650 3177 1696
rect 3233 1650 3285 1696
rect 5372 1650 5424 1696
rect 5480 1650 5532 1696
rect 5588 1650 5640 1696
rect 5696 1650 5748 1696
rect 5804 1650 5856 1696
rect 5912 1650 5964 1696
rect 6020 1650 6072 1696
rect 6128 1650 6180 1696
rect 6236 1650 6288 1696
rect 6344 1650 6396 1696
rect 7749 1650 7801 1696
rect 7857 1650 7909 1696
rect 7965 1650 8017 1696
rect 8073 1650 8125 1696
rect 8181 1650 8233 1696
rect 8289 1650 8341 1696
rect 8397 1650 8449 1696
rect 8505 1650 8557 1696
rect 8613 1650 8665 1696
rect 8721 1650 8773 1696
rect 8829 1650 8881 1696
rect 8937 1650 8989 1696
rect 9045 1650 9097 1696
rect 9153 1650 9205 1696
rect 9261 1650 9313 1696
rect 9369 1650 9421 1696
rect 9477 1650 9529 1696
rect 1505 1647 1557 1650
rect 1613 1647 1665 1650
rect 1721 1647 1773 1650
rect 1829 1647 1881 1650
rect 1937 1647 1989 1650
rect 2045 1647 2097 1650
rect 2153 1647 2205 1650
rect 2261 1647 2313 1650
rect 2369 1647 2421 1650
rect 2477 1647 2529 1650
rect 2585 1647 2637 1650
rect 2693 1647 2745 1650
rect 2801 1647 2853 1650
rect 2909 1647 2961 1650
rect 3017 1647 3069 1650
rect 3125 1647 3177 1650
rect 3233 1647 3285 1650
rect 5372 1647 5424 1650
rect 5480 1647 5532 1650
rect 5588 1647 5640 1650
rect 5696 1647 5748 1650
rect 5804 1647 5856 1650
rect 5912 1647 5964 1650
rect 6020 1647 6072 1650
rect 6128 1647 6180 1650
rect 6236 1647 6288 1650
rect 6344 1647 6396 1650
rect 7749 1647 7801 1650
rect 7857 1647 7909 1650
rect 7965 1647 8017 1650
rect 8073 1647 8125 1650
rect 8181 1647 8233 1650
rect 8289 1647 8341 1650
rect 8397 1647 8449 1650
rect 8505 1647 8557 1650
rect 8613 1647 8665 1650
rect 8721 1647 8773 1650
rect 8829 1647 8881 1650
rect 8937 1647 8989 1650
rect 9045 1647 9097 1650
rect 9153 1647 9205 1650
rect 9261 1647 9313 1650
rect 9369 1647 9421 1650
rect 9477 1647 9529 1650
rect 1233 1467 1285 1519
rect 1341 1467 1393 1519
rect 11569 6111 11621 6163
rect 11677 6111 11706 6163
rect 11706 6111 11729 6163
rect 11569 6003 11621 6055
rect 11677 6003 11706 6055
rect 11706 6003 11729 6055
rect 11569 5895 11621 5947
rect 11677 5895 11706 5947
rect 11706 5895 11729 5947
rect 11569 5787 11621 5839
rect 11677 5787 11706 5839
rect 11706 5787 11729 5839
rect 11569 5679 11621 5731
rect 11677 5679 11706 5731
rect 11706 5679 11729 5731
rect 11569 5571 11621 5623
rect 11677 5571 11706 5623
rect 11706 5571 11729 5623
rect 11569 5463 11621 5515
rect 11677 5463 11706 5515
rect 11706 5463 11729 5515
rect 11569 5355 11621 5407
rect 11677 5355 11706 5407
rect 11706 5355 11729 5407
rect 11569 5247 11621 5299
rect 11677 5247 11706 5299
rect 11706 5247 11729 5299
rect 11569 5139 11621 5191
rect 11677 5139 11706 5191
rect 11706 5139 11729 5191
rect 11569 5031 11621 5083
rect 11677 5031 11706 5083
rect 11706 5031 11729 5083
rect 11569 4923 11621 4975
rect 11677 4923 11706 4975
rect 11706 4923 11729 4975
rect 11569 4815 11621 4867
rect 11677 4815 11706 4867
rect 11706 4815 11729 4867
rect 11569 4707 11621 4759
rect 11677 4707 11706 4759
rect 11706 4707 11729 4759
rect 11569 4599 11621 4651
rect 11677 4599 11706 4651
rect 11706 4599 11729 4651
rect 11569 4491 11621 4543
rect 11677 4491 11706 4543
rect 11706 4491 11729 4543
rect 11569 4383 11621 4435
rect 11677 4383 11706 4435
rect 11706 4383 11729 4435
rect 11569 4275 11621 4327
rect 11677 4275 11706 4327
rect 11706 4275 11729 4327
rect 11569 4167 11621 4219
rect 11677 4167 11706 4219
rect 11706 4167 11729 4219
rect 11569 4059 11621 4111
rect 11677 4059 11706 4111
rect 11706 4059 11729 4111
rect 11569 3951 11621 4003
rect 11677 3951 11706 4003
rect 11706 3951 11729 4003
rect 11569 3843 11621 3895
rect 11677 3843 11706 3895
rect 11706 3843 11729 3895
rect 11569 3735 11621 3787
rect 11677 3735 11706 3787
rect 11706 3735 11729 3787
rect 11569 3627 11621 3679
rect 11677 3627 11706 3679
rect 11706 3627 11729 3679
rect 11569 3519 11621 3571
rect 11677 3519 11706 3571
rect 11706 3519 11729 3571
rect 11569 3411 11621 3463
rect 11677 3411 11706 3463
rect 11706 3411 11729 3463
rect 11569 3303 11621 3355
rect 11677 3303 11706 3355
rect 11706 3303 11729 3355
rect 11569 3195 11621 3247
rect 11677 3195 11706 3247
rect 11706 3195 11729 3247
rect 11569 3087 11621 3139
rect 11677 3087 11706 3139
rect 11706 3087 11729 3139
rect 11569 2979 11621 3031
rect 11677 2979 11706 3031
rect 11706 2979 11729 3031
rect 11569 2871 11621 2923
rect 11677 2871 11706 2923
rect 11706 2871 11729 2923
rect 11569 2763 11621 2815
rect 11677 2763 11706 2815
rect 11706 2763 11729 2815
rect 11569 2655 11621 2707
rect 11677 2655 11706 2707
rect 11706 2655 11729 2707
rect 11569 2547 11621 2599
rect 11677 2547 11706 2599
rect 11706 2547 11729 2599
rect 11569 2439 11621 2491
rect 11677 2439 11706 2491
rect 11706 2439 11729 2491
rect 11569 2331 11621 2383
rect 11677 2331 11706 2383
rect 11706 2331 11729 2383
rect 11569 2223 11621 2275
rect 11677 2223 11706 2275
rect 11706 2223 11729 2275
rect 11569 2115 11621 2167
rect 11677 2115 11706 2167
rect 11706 2115 11729 2167
rect 11569 2007 11621 2059
rect 11677 2007 11706 2059
rect 11706 2007 11729 2059
rect 11569 1899 11621 1951
rect 11677 1899 11706 1951
rect 11706 1899 11729 1951
rect 11569 1791 11621 1843
rect 11677 1791 11706 1843
rect 11706 1791 11729 1843
rect 11569 1683 11621 1735
rect 11677 1683 11706 1735
rect 11706 1683 11729 1735
rect 11569 1575 11621 1627
rect 11677 1575 11706 1627
rect 11706 1575 11729 1627
rect 11569 1467 11621 1519
rect 11677 1467 11729 1519
rect 3433 1452 3485 1455
rect 3541 1452 3593 1455
rect 3649 1452 3701 1455
rect 3757 1452 3809 1455
rect 3865 1452 3917 1455
rect 3973 1452 4025 1455
rect 4081 1452 4133 1455
rect 4189 1452 4241 1455
rect 4297 1452 4349 1455
rect 4405 1452 4457 1455
rect 4513 1452 4565 1455
rect 4621 1452 4673 1455
rect 4729 1452 4781 1455
rect 4837 1452 4889 1455
rect 4945 1452 4997 1455
rect 5053 1452 5105 1455
rect 5161 1452 5213 1455
rect 6566 1452 6618 1455
rect 6674 1452 6726 1455
rect 6782 1452 6834 1455
rect 6890 1452 6942 1455
rect 6998 1452 7050 1455
rect 7106 1452 7158 1455
rect 7214 1452 7266 1455
rect 7322 1452 7374 1455
rect 7430 1452 7482 1455
rect 7538 1452 7590 1455
rect 9677 1452 9729 1455
rect 9785 1452 9837 1455
rect 9893 1452 9945 1455
rect 10001 1452 10053 1455
rect 10109 1452 10161 1455
rect 10217 1452 10269 1455
rect 10325 1452 10377 1455
rect 10433 1452 10485 1455
rect 10541 1452 10593 1455
rect 10649 1452 10701 1455
rect 10757 1452 10809 1455
rect 10865 1452 10917 1455
rect 10973 1452 11025 1455
rect 11081 1452 11133 1455
rect 11189 1452 11241 1455
rect 11297 1452 11349 1455
rect 11405 1452 11457 1455
rect 3433 1406 3485 1452
rect 3541 1406 3593 1452
rect 3649 1406 3701 1452
rect 3757 1406 3809 1452
rect 3865 1406 3917 1452
rect 3973 1406 4025 1452
rect 4081 1406 4133 1452
rect 4189 1406 4241 1452
rect 4297 1406 4349 1452
rect 4405 1406 4457 1452
rect 4513 1406 4565 1452
rect 4621 1406 4673 1452
rect 4729 1406 4781 1452
rect 4837 1406 4889 1452
rect 4945 1406 4997 1452
rect 5053 1406 5105 1452
rect 5161 1406 5213 1452
rect 6566 1406 6618 1452
rect 6674 1406 6726 1452
rect 6782 1406 6834 1452
rect 6890 1406 6942 1452
rect 6998 1406 7050 1452
rect 7106 1406 7158 1452
rect 7214 1406 7266 1452
rect 7322 1406 7374 1452
rect 7430 1406 7482 1452
rect 7538 1406 7590 1452
rect 9677 1406 9729 1452
rect 9785 1406 9837 1452
rect 9893 1406 9945 1452
rect 10001 1406 10053 1452
rect 10109 1406 10161 1452
rect 10217 1406 10269 1452
rect 10325 1406 10377 1452
rect 10433 1406 10485 1452
rect 10541 1406 10593 1452
rect 10649 1406 10701 1452
rect 10757 1406 10809 1452
rect 10865 1406 10917 1452
rect 10973 1406 11025 1452
rect 11081 1406 11133 1452
rect 11189 1406 11241 1452
rect 11297 1406 11349 1452
rect 11405 1406 11457 1452
rect 3433 1403 3485 1406
rect 3541 1403 3593 1406
rect 3649 1403 3701 1406
rect 3757 1403 3809 1406
rect 3865 1403 3917 1406
rect 3973 1403 4025 1406
rect 4081 1403 4133 1406
rect 4189 1403 4241 1406
rect 4297 1403 4349 1406
rect 4405 1403 4457 1406
rect 4513 1403 4565 1406
rect 4621 1403 4673 1406
rect 4729 1403 4781 1406
rect 4837 1403 4889 1406
rect 4945 1403 4997 1406
rect 5053 1403 5105 1406
rect 5161 1403 5213 1406
rect 6566 1403 6618 1406
rect 6674 1403 6726 1406
rect 6782 1403 6834 1406
rect 6890 1403 6942 1406
rect 6998 1403 7050 1406
rect 7106 1403 7158 1406
rect 7214 1403 7266 1406
rect 7322 1403 7374 1406
rect 7430 1403 7482 1406
rect 7538 1403 7590 1406
rect 9677 1403 9729 1406
rect 9785 1403 9837 1406
rect 9893 1403 9945 1406
rect 10001 1403 10053 1406
rect 10109 1403 10161 1406
rect 10217 1403 10269 1406
rect 10325 1403 10377 1406
rect 10433 1403 10485 1406
rect 10541 1403 10593 1406
rect 10649 1403 10701 1406
rect 10757 1403 10809 1406
rect 10865 1403 10917 1406
rect 10973 1403 11025 1406
rect 11081 1403 11133 1406
rect 11189 1403 11241 1406
rect 11297 1403 11349 1406
rect 11405 1403 11457 1406
rect 12051 6657 12103 6709
rect 12159 6657 12211 6709
rect 12267 6657 12319 6709
rect 12051 6549 12103 6601
rect 12159 6549 12211 6601
rect 12267 6549 12319 6601
rect 12051 6441 12103 6493
rect 12159 6441 12211 6493
rect 12267 6441 12319 6493
rect 12051 6333 12103 6385
rect 12159 6333 12211 6385
rect 12267 6333 12319 6385
rect 12051 6225 12103 6277
rect 12159 6225 12211 6277
rect 12267 6225 12319 6277
rect 12051 6117 12103 6169
rect 12159 6117 12211 6169
rect 12267 6117 12319 6169
rect 12051 6009 12103 6061
rect 12159 6009 12211 6061
rect 12267 6009 12319 6061
rect 12051 5901 12103 5953
rect 12159 5901 12211 5953
rect 12267 5901 12319 5953
rect 12051 5793 12103 5845
rect 12159 5793 12211 5845
rect 12267 5793 12319 5845
rect 12051 5685 12103 5737
rect 12159 5685 12211 5737
rect 12267 5685 12319 5737
rect 12051 5577 12103 5629
rect 12159 5577 12211 5629
rect 12267 5577 12319 5629
rect 12051 5469 12103 5521
rect 12159 5469 12211 5521
rect 12267 5469 12319 5521
rect 12051 5361 12103 5413
rect 12159 5361 12211 5413
rect 12267 5361 12319 5413
rect 12051 5253 12103 5305
rect 12159 5253 12211 5305
rect 12267 5253 12319 5305
rect 12051 5145 12103 5197
rect 12159 5145 12211 5197
rect 12267 5145 12319 5197
rect 12051 5037 12103 5089
rect 12159 5037 12211 5089
rect 12267 5037 12319 5089
rect 12051 4929 12103 4981
rect 12159 4929 12211 4981
rect 12267 4929 12319 4981
rect 12051 4821 12103 4873
rect 12159 4821 12211 4873
rect 12267 4821 12319 4873
rect 12051 4713 12103 4765
rect 12159 4713 12211 4765
rect 12267 4713 12319 4765
rect 12051 4605 12103 4657
rect 12159 4605 12211 4657
rect 12267 4605 12319 4657
rect 12051 4497 12103 4549
rect 12159 4497 12211 4549
rect 12267 4497 12319 4549
rect 12051 4389 12103 4441
rect 12159 4389 12211 4441
rect 12267 4389 12319 4441
rect 12051 4281 12103 4333
rect 12159 4281 12211 4333
rect 12267 4281 12319 4333
rect 12051 4173 12103 4225
rect 12159 4173 12211 4225
rect 12267 4173 12319 4225
rect 12051 4065 12103 4117
rect 12159 4065 12211 4117
rect 12267 4065 12319 4117
rect 12051 3957 12103 4009
rect 12159 3957 12211 4009
rect 12267 3957 12319 4009
rect 12051 3849 12103 3901
rect 12159 3849 12211 3901
rect 12267 3849 12319 3901
rect 12051 3741 12103 3793
rect 12159 3741 12211 3793
rect 12267 3741 12319 3793
rect 12051 3633 12103 3685
rect 12159 3633 12211 3685
rect 12267 3633 12319 3685
rect 12051 3525 12103 3577
rect 12159 3525 12211 3577
rect 12267 3525 12319 3577
rect 12051 3417 12103 3469
rect 12159 3417 12211 3469
rect 12267 3417 12319 3469
rect 12051 3309 12103 3361
rect 12159 3309 12211 3361
rect 12267 3309 12319 3361
rect 12051 3201 12103 3253
rect 12159 3201 12211 3253
rect 12267 3201 12319 3253
rect 12051 3093 12103 3145
rect 12159 3093 12211 3145
rect 12267 3093 12319 3145
rect 12051 2985 12103 3037
rect 12159 2985 12211 3037
rect 12267 2985 12319 3037
rect 12051 2877 12103 2929
rect 12159 2877 12211 2929
rect 12267 2877 12319 2929
rect 12051 2769 12103 2821
rect 12159 2769 12211 2821
rect 12267 2769 12319 2821
rect 12051 2661 12103 2713
rect 12159 2661 12211 2713
rect 12267 2661 12319 2713
rect 12051 2553 12103 2605
rect 12159 2553 12211 2605
rect 12267 2553 12319 2605
rect 12051 2445 12103 2497
rect 12159 2445 12211 2497
rect 12267 2445 12319 2497
rect 12051 2337 12103 2389
rect 12159 2337 12211 2389
rect 12267 2337 12319 2389
rect 12051 2229 12103 2281
rect 12159 2229 12211 2281
rect 12267 2229 12319 2281
rect 12051 2121 12103 2173
rect 12159 2121 12211 2173
rect 12267 2121 12319 2173
rect 12051 2013 12103 2065
rect 12159 2013 12211 2065
rect 12267 2013 12319 2065
rect 12051 1905 12103 1957
rect 12159 1905 12211 1957
rect 12267 1905 12319 1957
rect 12051 1797 12103 1849
rect 12159 1797 12211 1849
rect 12267 1797 12319 1849
rect 12051 1689 12103 1741
rect 12159 1689 12211 1741
rect 12267 1689 12319 1741
rect 12051 1581 12103 1633
rect 12159 1581 12211 1633
rect 12267 1581 12319 1633
rect 12051 1473 12103 1525
rect 12159 1473 12211 1525
rect 12267 1473 12319 1525
rect 12051 1365 12103 1417
rect 12159 1365 12211 1417
rect 12267 1365 12319 1417
rect 12051 1257 12103 1309
rect 12159 1257 12211 1309
rect 12267 1257 12319 1309
rect 12051 1149 12103 1201
rect 12159 1149 12211 1201
rect 12267 1149 12319 1201
rect 12051 1041 12103 1093
rect 12159 1041 12211 1093
rect 12267 1041 12319 1093
rect 1505 909 1557 961
rect 1613 909 1665 961
rect 1721 909 1773 961
rect 1829 909 1881 961
rect 1937 909 1989 961
rect 2045 909 2097 961
rect 2153 909 2205 961
rect 2261 909 2313 961
rect 2369 909 2421 961
rect 2477 909 2529 961
rect 2585 909 2637 961
rect 2693 909 2745 961
rect 2801 909 2853 961
rect 2909 909 2961 961
rect 3017 909 3069 961
rect 3125 909 3177 961
rect 3233 909 3285 961
rect 5372 909 5424 961
rect 5480 909 5532 961
rect 5588 909 5640 961
rect 5696 909 5748 961
rect 5804 909 5856 961
rect 5912 909 5964 961
rect 6020 909 6072 961
rect 6128 909 6180 961
rect 6236 909 6288 961
rect 6344 909 6396 961
rect 7749 909 7801 961
rect 7857 909 7909 961
rect 7965 909 8017 961
rect 8073 909 8125 961
rect 8181 909 8233 961
rect 8289 909 8341 961
rect 8397 909 8449 961
rect 8505 909 8557 961
rect 8613 909 8665 961
rect 8721 909 8773 961
rect 8829 909 8881 961
rect 8937 909 8989 961
rect 9045 909 9097 961
rect 9153 909 9205 961
rect 9261 909 9313 961
rect 9369 909 9421 961
rect 9477 909 9529 961
rect 1505 801 1557 853
rect 1613 801 1665 853
rect 1721 801 1773 853
rect 1829 801 1881 853
rect 1937 801 1989 853
rect 2045 801 2097 853
rect 2153 801 2205 853
rect 2261 801 2313 853
rect 2369 801 2421 853
rect 2477 801 2529 853
rect 2585 801 2637 853
rect 2693 801 2745 853
rect 2801 801 2853 853
rect 2909 801 2961 853
rect 3017 801 3069 853
rect 3125 801 3177 853
rect 3233 801 3285 853
rect 5372 801 5424 853
rect 5480 801 5532 853
rect 5588 801 5640 853
rect 5696 801 5748 853
rect 5804 801 5856 853
rect 5912 801 5964 853
rect 6020 801 6072 853
rect 6128 801 6180 853
rect 6236 801 6288 853
rect 6344 801 6396 853
rect 7749 801 7801 853
rect 7857 801 7909 853
rect 7965 801 8017 853
rect 8073 801 8125 853
rect 8181 801 8233 853
rect 8289 801 8341 853
rect 8397 801 8449 853
rect 8505 801 8557 853
rect 8613 801 8665 853
rect 8721 801 8773 853
rect 8829 801 8881 853
rect 8937 801 8989 853
rect 9045 801 9097 853
rect 9153 801 9205 853
rect 9261 801 9313 853
rect 9369 801 9421 853
rect 9477 801 9529 853
rect 1505 693 1557 745
rect 1613 693 1665 745
rect 1721 693 1773 745
rect 1829 693 1881 745
rect 1937 693 1989 745
rect 2045 693 2097 745
rect 2153 693 2205 745
rect 2261 693 2313 745
rect 2369 693 2421 745
rect 2477 693 2529 745
rect 2585 693 2637 745
rect 2693 693 2745 745
rect 2801 693 2853 745
rect 2909 693 2961 745
rect 3017 693 3069 745
rect 3125 693 3177 745
rect 3233 693 3285 745
rect 5372 693 5424 745
rect 5480 693 5532 745
rect 5588 693 5640 745
rect 5696 693 5748 745
rect 5804 693 5856 745
rect 5912 693 5964 745
rect 6020 693 6072 745
rect 6128 693 6180 745
rect 6236 693 6288 745
rect 6344 693 6396 745
rect 7749 693 7801 745
rect 7857 693 7909 745
rect 7965 693 8017 745
rect 8073 693 8125 745
rect 8181 693 8233 745
rect 8289 693 8341 745
rect 8397 693 8449 745
rect 8505 693 8557 745
rect 8613 693 8665 745
rect 8721 693 8773 745
rect 8829 693 8881 745
rect 8937 693 8989 745
rect 9045 693 9097 745
rect 9153 693 9205 745
rect 9261 693 9313 745
rect 9369 693 9421 745
rect 9477 693 9529 745
rect 12051 933 12103 985
rect 12159 933 12211 985
rect 12267 933 12319 985
rect 12051 825 12103 877
rect 12159 825 12211 877
rect 12267 825 12319 877
rect 12051 717 12103 769
rect 12159 717 12211 769
rect 12267 717 12319 769
rect 82 309 134 361
rect 190 309 242 361
rect 298 309 350 361
rect 406 309 458 361
rect 514 309 566 361
rect 622 309 674 361
rect 730 309 782 361
rect 838 309 890 361
rect 946 309 998 361
rect 1054 309 1106 361
rect 3433 309 3485 361
rect 3541 309 3593 361
rect 3649 309 3701 361
rect 3757 309 3809 361
rect 3865 309 3917 361
rect 3973 309 4025 361
rect 4081 309 4133 361
rect 4189 309 4241 361
rect 4297 309 4349 361
rect 4405 309 4457 361
rect 4513 309 4565 361
rect 4621 309 4673 361
rect 4729 309 4781 361
rect 4837 309 4889 361
rect 4945 309 4997 361
rect 5053 309 5105 361
rect 5161 309 5213 361
rect 6566 309 6618 361
rect 6674 309 6726 361
rect 6782 309 6834 361
rect 6890 309 6942 361
rect 6998 309 7050 361
rect 7106 309 7158 361
rect 7214 309 7266 361
rect 7322 309 7374 361
rect 7430 309 7482 361
rect 7538 309 7590 361
rect 9677 309 9729 361
rect 9785 309 9837 361
rect 9893 309 9945 361
rect 10001 309 10053 361
rect 10109 309 10161 361
rect 10217 309 10269 361
rect 10325 309 10377 361
rect 10433 309 10485 361
rect 10541 309 10593 361
rect 10649 309 10701 361
rect 10757 309 10809 361
rect 10865 309 10917 361
rect 10973 309 11025 361
rect 11081 309 11133 361
rect 11189 309 11241 361
rect 11297 309 11349 361
rect 11405 309 11457 361
rect 82 201 134 253
rect 190 201 242 253
rect 298 201 350 253
rect 406 201 458 253
rect 514 201 566 253
rect 622 201 674 253
rect 730 201 782 253
rect 838 201 890 253
rect 946 201 998 253
rect 1054 201 1106 253
rect 3433 201 3485 253
rect 3541 201 3593 253
rect 3649 201 3701 253
rect 3757 201 3809 253
rect 3865 201 3917 253
rect 3973 201 4025 253
rect 4081 201 4133 253
rect 4189 201 4241 253
rect 4297 201 4349 253
rect 4405 201 4457 253
rect 4513 201 4565 253
rect 4621 201 4673 253
rect 4729 201 4781 253
rect 4837 201 4889 253
rect 4945 201 4997 253
rect 5053 201 5105 253
rect 5161 201 5213 253
rect 6566 201 6618 253
rect 6674 201 6726 253
rect 6782 201 6834 253
rect 6890 201 6942 253
rect 6998 201 7050 253
rect 7106 201 7158 253
rect 7214 201 7266 253
rect 7322 201 7374 253
rect 7430 201 7482 253
rect 7538 201 7590 253
rect 9677 201 9729 253
rect 9785 201 9837 253
rect 9893 201 9945 253
rect 10001 201 10053 253
rect 10109 201 10161 253
rect 10217 201 10269 253
rect 10325 201 10377 253
rect 10433 201 10485 253
rect 10541 201 10593 253
rect 10649 201 10701 253
rect 10757 201 10809 253
rect 10865 201 10917 253
rect 10973 201 11025 253
rect 11081 201 11133 253
rect 11189 201 11241 253
rect 11297 201 11349 253
rect 11405 201 11457 253
rect 82 93 134 145
rect 190 93 242 145
rect 298 93 350 145
rect 406 93 458 145
rect 514 93 566 145
rect 622 93 674 145
rect 730 93 782 145
rect 838 93 890 145
rect 946 93 998 145
rect 1054 93 1106 145
rect 3433 93 3485 145
rect 3541 93 3593 145
rect 3649 93 3701 145
rect 3757 93 3809 145
rect 3865 93 3917 145
rect 3973 93 4025 145
rect 4081 93 4133 145
rect 4189 93 4241 145
rect 4297 93 4349 145
rect 4405 93 4457 145
rect 4513 93 4565 145
rect 4621 93 4673 145
rect 4729 93 4781 145
rect 4837 93 4889 145
rect 4945 93 4997 145
rect 5053 93 5105 145
rect 5161 93 5213 145
rect 6566 93 6618 145
rect 6674 93 6726 145
rect 6782 93 6834 145
rect 6890 93 6942 145
rect 6998 93 7050 145
rect 7106 93 7158 145
rect 7214 93 7266 145
rect 7322 93 7374 145
rect 7430 93 7482 145
rect 7538 93 7590 145
rect 9677 93 9729 145
rect 9785 93 9837 145
rect 9893 93 9945 145
rect 10001 93 10053 145
rect 10109 93 10161 145
rect 10217 93 10269 145
rect 10325 93 10377 145
rect 10433 93 10485 145
rect 10541 93 10593 145
rect 10649 93 10701 145
rect 10757 93 10809 145
rect 10865 93 10917 145
rect 10973 93 11025 145
rect 11081 93 11133 145
rect 11189 93 11241 145
rect 11297 93 11349 145
rect 11405 93 11457 145
<< metal2 >>
rect 43 25261 1145 25617
rect 43 25209 82 25261
rect 134 25209 190 25261
rect 242 25209 298 25261
rect 350 25209 406 25261
rect 458 25209 514 25261
rect 566 25209 622 25261
rect 674 25209 730 25261
rect 782 25209 838 25261
rect 890 25209 946 25261
rect 998 25209 1054 25261
rect 1106 25209 1145 25261
rect 43 25153 1145 25209
rect 43 25101 82 25153
rect 134 25101 190 25153
rect 242 25101 298 25153
rect 350 25101 406 25153
rect 458 25101 514 25153
rect 566 25101 622 25153
rect 674 25101 730 25153
rect 782 25101 838 25153
rect 890 25101 946 25153
rect 998 25101 1054 25153
rect 1106 25101 1145 25153
rect 43 25045 1145 25101
rect 43 24993 82 25045
rect 134 24993 190 25045
rect 242 24993 298 25045
rect 350 24993 406 25045
rect 458 24993 514 25045
rect 566 24993 622 25045
rect 674 24993 730 25045
rect 782 24993 838 25045
rect 890 24993 946 25045
rect 998 24993 1054 25045
rect 1106 24993 1145 25045
rect 43 24853 1145 24993
rect 43 24801 93 24853
rect 145 24801 201 24853
rect 253 24801 309 24853
rect 361 24801 1145 24853
rect 43 24745 1145 24801
rect 43 24693 93 24745
rect 145 24693 201 24745
rect 253 24693 309 24745
rect 361 24693 1145 24745
rect 43 24637 1145 24693
rect 43 24585 93 24637
rect 145 24585 201 24637
rect 253 24585 309 24637
rect 361 24585 1145 24637
rect 43 24529 1145 24585
rect 43 24477 93 24529
rect 145 24477 201 24529
rect 253 24477 309 24529
rect 361 24477 1145 24529
rect 43 24421 1145 24477
rect 43 24369 93 24421
rect 145 24369 201 24421
rect 253 24369 309 24421
rect 361 24369 1145 24421
rect 43 24313 1145 24369
rect 43 24261 93 24313
rect 145 24261 201 24313
rect 253 24261 309 24313
rect 361 24261 1145 24313
rect 43 24205 1145 24261
rect 43 24153 93 24205
rect 145 24153 201 24205
rect 253 24153 309 24205
rect 361 24153 1145 24205
rect 43 24097 1145 24153
rect 43 24045 93 24097
rect 145 24045 201 24097
rect 253 24045 309 24097
rect 361 24045 1145 24097
rect 43 23989 1145 24045
rect 43 23937 93 23989
rect 145 23937 201 23989
rect 253 23937 309 23989
rect 361 23937 1145 23989
rect 43 23881 1145 23937
rect 43 23829 93 23881
rect 145 23829 201 23881
rect 253 23829 309 23881
rect 361 23829 1145 23881
rect 43 23773 1145 23829
rect 43 23721 93 23773
rect 145 23721 201 23773
rect 253 23721 309 23773
rect 361 23721 1145 23773
rect 43 23665 1145 23721
rect 43 23613 93 23665
rect 145 23613 201 23665
rect 253 23613 309 23665
rect 361 23613 1145 23665
rect 43 23557 1145 23613
rect 43 23505 93 23557
rect 145 23505 201 23557
rect 253 23505 309 23557
rect 361 23505 1145 23557
rect 43 23449 1145 23505
rect 43 23397 93 23449
rect 145 23397 201 23449
rect 253 23397 309 23449
rect 361 23397 1145 23449
rect 43 23341 1145 23397
rect 43 23289 93 23341
rect 145 23289 201 23341
rect 253 23289 309 23341
rect 361 23289 1145 23341
rect 43 23233 1145 23289
rect 43 23181 93 23233
rect 145 23181 201 23233
rect 253 23181 309 23233
rect 361 23181 1145 23233
rect 43 23125 1145 23181
rect 43 23073 93 23125
rect 145 23073 201 23125
rect 253 23073 309 23125
rect 361 23073 1145 23125
rect 43 23017 1145 23073
rect 43 22965 93 23017
rect 145 22965 201 23017
rect 253 22965 309 23017
rect 361 22965 1145 23017
rect 43 22909 1145 22965
rect 43 22857 93 22909
rect 145 22857 201 22909
rect 253 22857 309 22909
rect 361 22857 1145 22909
rect 43 22801 1145 22857
rect 43 22749 93 22801
rect 145 22749 201 22801
rect 253 22749 309 22801
rect 361 22749 1145 22801
rect 43 22693 1145 22749
rect 43 22641 93 22693
rect 145 22641 201 22693
rect 253 22641 309 22693
rect 361 22641 1145 22693
rect 43 22585 1145 22641
rect 43 22533 93 22585
rect 145 22533 201 22585
rect 253 22533 309 22585
rect 361 22533 1145 22585
rect 43 22477 1145 22533
rect 43 22425 93 22477
rect 145 22425 201 22477
rect 253 22425 309 22477
rect 361 22425 1145 22477
rect 43 22369 1145 22425
rect 43 22317 93 22369
rect 145 22317 201 22369
rect 253 22317 309 22369
rect 361 22317 1145 22369
rect 43 22261 1145 22317
rect 43 22209 93 22261
rect 145 22209 201 22261
rect 253 22209 309 22261
rect 361 22209 1145 22261
rect 43 22153 1145 22209
rect 43 22101 93 22153
rect 145 22101 201 22153
rect 253 22101 309 22153
rect 361 22101 1145 22153
rect 43 22045 1145 22101
rect 43 21993 93 22045
rect 145 21993 201 22045
rect 253 21993 309 22045
rect 361 21993 1145 22045
rect 43 21937 1145 21993
rect 43 21885 93 21937
rect 145 21885 201 21937
rect 253 21885 309 21937
rect 361 21885 1145 21937
rect 43 21829 1145 21885
rect 43 21777 93 21829
rect 145 21777 201 21829
rect 253 21777 309 21829
rect 361 21777 1145 21829
rect 43 21721 1145 21777
rect 43 21669 93 21721
rect 145 21669 201 21721
rect 253 21669 309 21721
rect 361 21669 1145 21721
rect 43 21613 1145 21669
rect 43 21561 93 21613
rect 145 21561 201 21613
rect 253 21561 309 21613
rect 361 21561 1145 21613
rect 43 21505 1145 21561
rect 43 21453 93 21505
rect 145 21453 201 21505
rect 253 21453 309 21505
rect 361 21453 1145 21505
rect 43 21397 1145 21453
rect 43 21345 93 21397
rect 145 21345 201 21397
rect 253 21345 309 21397
rect 361 21345 1145 21397
rect 43 21289 1145 21345
rect 43 21237 93 21289
rect 145 21237 201 21289
rect 253 21237 309 21289
rect 361 21237 1145 21289
rect 43 21181 1145 21237
rect 43 21129 93 21181
rect 145 21129 201 21181
rect 253 21129 309 21181
rect 361 21129 1145 21181
rect 43 21073 1145 21129
rect 43 21021 93 21073
rect 145 21021 201 21073
rect 253 21021 309 21073
rect 361 21021 1145 21073
rect 43 20965 1145 21021
rect 43 20913 93 20965
rect 145 20913 201 20965
rect 253 20913 309 20965
rect 361 20913 1145 20965
rect 43 20857 1145 20913
rect 43 20805 93 20857
rect 145 20805 201 20857
rect 253 20805 309 20857
rect 361 20805 1145 20857
rect 43 20749 1145 20805
rect 43 20697 93 20749
rect 145 20697 201 20749
rect 253 20697 309 20749
rect 361 20697 1145 20749
rect 43 20641 1145 20697
rect 43 20589 93 20641
rect 145 20589 201 20641
rect 253 20589 309 20641
rect 361 20589 1145 20641
rect 43 20533 1145 20589
rect 43 20481 93 20533
rect 145 20481 201 20533
rect 253 20481 309 20533
rect 361 20481 1145 20533
rect 43 20425 1145 20481
rect 43 20373 93 20425
rect 145 20373 201 20425
rect 253 20373 309 20425
rect 361 20373 1145 20425
rect 43 20317 1145 20373
rect 43 20265 93 20317
rect 145 20265 201 20317
rect 253 20265 309 20317
rect 361 20265 1145 20317
rect 43 20209 1145 20265
rect 43 20157 93 20209
rect 145 20157 201 20209
rect 253 20157 309 20209
rect 361 20157 1145 20209
rect 43 20101 1145 20157
rect 43 20049 93 20101
rect 145 20049 201 20101
rect 253 20049 309 20101
rect 361 20049 1145 20101
rect 43 19993 1145 20049
rect 43 19941 93 19993
rect 145 19941 201 19993
rect 253 19941 309 19993
rect 361 19941 1145 19993
rect 43 19885 1145 19941
rect 43 19833 93 19885
rect 145 19833 201 19885
rect 253 19833 309 19885
rect 361 19833 1145 19885
rect 43 19777 1145 19833
rect 43 19725 93 19777
rect 145 19725 201 19777
rect 253 19725 309 19777
rect 361 19725 1145 19777
rect 43 19669 1145 19725
rect 43 19617 93 19669
rect 145 19617 201 19669
rect 253 19617 309 19669
rect 361 19617 1145 19669
rect 43 19561 1145 19617
rect 43 19509 93 19561
rect 145 19509 201 19561
rect 253 19509 309 19561
rect 361 19509 1145 19561
rect 43 19453 1145 19509
rect 43 19401 93 19453
rect 145 19401 201 19453
rect 253 19401 309 19453
rect 361 19401 1145 19453
rect 43 19345 1145 19401
rect 43 19293 93 19345
rect 145 19293 201 19345
rect 253 19293 309 19345
rect 361 19293 1145 19345
rect 43 19237 1145 19293
rect 43 19185 93 19237
rect 145 19185 201 19237
rect 253 19185 309 19237
rect 361 19185 1145 19237
rect 43 19129 1145 19185
rect 43 19077 93 19129
rect 145 19077 201 19129
rect 253 19077 309 19129
rect 361 19077 1145 19129
rect 43 19021 1145 19077
rect 43 18969 93 19021
rect 145 18969 201 19021
rect 253 18969 309 19021
rect 361 18969 1145 19021
rect 43 18913 1145 18969
rect 43 18861 93 18913
rect 145 18861 201 18913
rect 253 18861 309 18913
rect 361 18861 1145 18913
rect 43 18805 1145 18861
rect 43 18753 93 18805
rect 145 18753 201 18805
rect 253 18753 309 18805
rect 361 18753 1145 18805
rect 43 18697 1145 18753
rect 43 18645 93 18697
rect 145 18645 201 18697
rect 253 18645 309 18697
rect 361 18645 1145 18697
rect 43 18589 1145 18645
rect 43 18537 93 18589
rect 145 18537 201 18589
rect 253 18537 309 18589
rect 361 18537 1145 18589
rect 43 18481 1145 18537
rect 43 18429 93 18481
rect 145 18429 201 18481
rect 253 18429 309 18481
rect 361 18429 1145 18481
rect 43 18373 1145 18429
rect 43 18321 93 18373
rect 145 18321 201 18373
rect 253 18321 309 18373
rect 361 18321 1145 18373
rect 43 18265 1145 18321
rect 43 18213 93 18265
rect 145 18213 201 18265
rect 253 18213 309 18265
rect 361 18213 1145 18265
rect 43 18157 1145 18213
rect 43 18105 93 18157
rect 145 18105 201 18157
rect 253 18105 309 18157
rect 361 18105 1145 18157
rect 43 18049 1145 18105
rect 43 17997 93 18049
rect 145 17997 201 18049
rect 253 17997 309 18049
rect 361 17997 1145 18049
rect 43 17941 1145 17997
rect 43 17889 93 17941
rect 145 17889 201 17941
rect 253 17889 309 17941
rect 361 17889 1145 17941
rect 43 17833 1145 17889
rect 43 17781 93 17833
rect 145 17781 201 17833
rect 253 17781 309 17833
rect 361 17781 1145 17833
rect 43 17725 1145 17781
rect 43 17673 93 17725
rect 145 17673 201 17725
rect 253 17673 309 17725
rect 361 17673 1145 17725
rect 43 17617 1145 17673
rect 43 17565 93 17617
rect 145 17565 201 17617
rect 253 17565 309 17617
rect 361 17565 1145 17617
rect 43 17509 1145 17565
rect 43 17457 93 17509
rect 145 17457 201 17509
rect 253 17457 309 17509
rect 361 17457 1145 17509
rect 43 17401 1145 17457
rect 43 17349 93 17401
rect 145 17349 201 17401
rect 253 17349 309 17401
rect 361 17349 1145 17401
rect 43 17293 1145 17349
rect 43 17241 93 17293
rect 145 17241 201 17293
rect 253 17241 309 17293
rect 361 17241 1145 17293
rect 43 17185 1145 17241
rect 43 17133 93 17185
rect 145 17133 201 17185
rect 253 17133 309 17185
rect 361 17133 1145 17185
rect 43 17077 1145 17133
rect 43 17025 93 17077
rect 145 17025 201 17077
rect 253 17025 309 17077
rect 361 17025 1145 17077
rect 43 16969 1145 17025
rect 43 16917 93 16969
rect 145 16917 201 16969
rect 253 16917 309 16969
rect 361 16917 1145 16969
rect 43 16861 1145 16917
rect 43 16809 93 16861
rect 145 16809 201 16861
rect 253 16809 309 16861
rect 361 16809 1145 16861
rect 43 16753 1145 16809
rect 43 16701 93 16753
rect 145 16701 201 16753
rect 253 16701 309 16753
rect 361 16701 1145 16753
rect 43 16645 1145 16701
rect 43 16593 93 16645
rect 145 16593 201 16645
rect 253 16593 309 16645
rect 361 16593 1145 16645
rect 43 16537 1145 16593
rect 43 16485 93 16537
rect 145 16485 201 16537
rect 253 16485 309 16537
rect 361 16485 1145 16537
rect 43 16429 1145 16485
rect 43 16377 93 16429
rect 145 16377 201 16429
rect 253 16377 309 16429
rect 361 16377 1145 16429
rect 43 16321 1145 16377
rect 43 16269 93 16321
rect 145 16269 201 16321
rect 253 16269 309 16321
rect 361 16269 1145 16321
rect 43 16213 1145 16269
rect 43 16161 93 16213
rect 145 16161 201 16213
rect 253 16161 309 16213
rect 361 16161 1145 16213
rect 43 16105 1145 16161
rect 43 16053 93 16105
rect 145 16053 201 16105
rect 253 16053 309 16105
rect 361 16053 1145 16105
rect 43 15997 1145 16053
rect 43 15945 93 15997
rect 145 15945 201 15997
rect 253 15945 309 15997
rect 361 15945 1145 15997
rect 43 15889 1145 15945
rect 43 15837 93 15889
rect 145 15837 201 15889
rect 253 15837 309 15889
rect 361 15837 1145 15889
rect 43 15781 1145 15837
rect 43 15729 93 15781
rect 145 15729 201 15781
rect 253 15729 309 15781
rect 361 15729 1145 15781
rect 43 15673 1145 15729
rect 43 15621 93 15673
rect 145 15621 201 15673
rect 253 15621 309 15673
rect 361 15621 1145 15673
rect 43 15565 1145 15621
rect 43 15513 93 15565
rect 145 15513 201 15565
rect 253 15513 309 15565
rect 361 15513 1145 15565
rect 43 15457 1145 15513
rect 43 15405 93 15457
rect 145 15405 201 15457
rect 253 15405 309 15457
rect 361 15405 1145 15457
rect 43 15349 1145 15405
rect 43 15297 93 15349
rect 145 15297 201 15349
rect 253 15297 309 15349
rect 361 15297 1145 15349
rect 43 15241 1145 15297
rect 43 15189 93 15241
rect 145 15189 201 15241
rect 253 15189 309 15241
rect 361 15189 1145 15241
rect 43 15133 1145 15189
rect 43 15081 93 15133
rect 145 15081 201 15133
rect 253 15081 309 15133
rect 361 15081 1145 15133
rect 43 15025 1145 15081
rect 43 14973 93 15025
rect 145 14973 201 15025
rect 253 14973 309 15025
rect 361 14973 1145 15025
rect 43 14917 1145 14973
rect 43 14865 93 14917
rect 145 14865 201 14917
rect 253 14865 309 14917
rect 361 14865 1145 14917
rect 43 14809 1145 14865
rect 43 14757 93 14809
rect 145 14757 201 14809
rect 253 14757 309 14809
rect 361 14757 1145 14809
rect 43 14701 1145 14757
rect 43 14649 93 14701
rect 145 14649 201 14701
rect 253 14649 309 14701
rect 361 14649 1145 14701
rect 43 14593 1145 14649
rect 43 14541 93 14593
rect 145 14541 201 14593
rect 253 14541 309 14593
rect 361 14541 1145 14593
rect 43 14485 1145 14541
rect 43 14433 93 14485
rect 145 14433 201 14485
rect 253 14433 309 14485
rect 361 14433 1145 14485
rect 43 14377 1145 14433
rect 43 14325 93 14377
rect 145 14325 201 14377
rect 253 14325 309 14377
rect 361 14325 1145 14377
rect 43 14269 1145 14325
rect 43 14217 93 14269
rect 145 14217 201 14269
rect 253 14217 309 14269
rect 361 14217 1145 14269
rect 43 14161 1145 14217
rect 43 14109 93 14161
rect 145 14109 201 14161
rect 253 14109 309 14161
rect 361 14109 1145 14161
rect 43 14053 1145 14109
rect 43 14001 93 14053
rect 145 14001 201 14053
rect 253 14001 309 14053
rect 361 14001 1145 14053
rect 43 13945 1145 14001
rect 43 13893 93 13945
rect 145 13893 201 13945
rect 253 13893 309 13945
rect 361 13893 1145 13945
rect 43 13837 1145 13893
rect 43 13785 93 13837
rect 145 13785 201 13837
rect 253 13785 309 13837
rect 361 13785 1145 13837
rect 43 13729 1145 13785
rect 43 13677 93 13729
rect 145 13677 201 13729
rect 253 13677 309 13729
rect 361 13677 1145 13729
rect 43 13621 1145 13677
rect 43 13569 93 13621
rect 145 13569 201 13621
rect 253 13569 309 13621
rect 361 13569 1145 13621
rect 43 13513 1145 13569
rect 43 13461 93 13513
rect 145 13461 201 13513
rect 253 13461 309 13513
rect 361 13461 1145 13513
rect 43 13405 1145 13461
rect 43 13353 93 13405
rect 145 13353 201 13405
rect 253 13353 309 13405
rect 361 13353 1145 13405
rect 43 13297 1145 13353
rect 43 13245 93 13297
rect 145 13245 201 13297
rect 253 13245 309 13297
rect 361 13245 1145 13297
rect 43 13189 1145 13245
rect 43 13137 93 13189
rect 145 13137 201 13189
rect 253 13137 309 13189
rect 361 13137 1145 13189
rect 43 13081 1145 13137
rect 43 13029 93 13081
rect 145 13029 201 13081
rect 253 13029 309 13081
rect 361 13029 1145 13081
rect 43 12973 1145 13029
rect 43 12921 93 12973
rect 145 12921 201 12973
rect 253 12921 309 12973
rect 361 12921 1145 12973
rect 43 12865 1145 12921
rect 43 12813 93 12865
rect 145 12813 201 12865
rect 253 12813 309 12865
rect 361 12813 1145 12865
rect 43 12757 1145 12813
rect 43 12705 93 12757
rect 145 12705 201 12757
rect 253 12705 309 12757
rect 361 12705 1145 12757
rect 43 12649 1145 12705
rect 43 12597 93 12649
rect 145 12597 201 12649
rect 253 12597 309 12649
rect 361 12597 1145 12649
rect 43 12541 1145 12597
rect 43 12489 93 12541
rect 145 12489 201 12541
rect 253 12489 309 12541
rect 361 12489 1145 12541
rect 43 12433 1145 12489
rect 43 12381 93 12433
rect 145 12381 201 12433
rect 253 12381 309 12433
rect 361 12381 1145 12433
rect 43 12325 1145 12381
rect 43 12273 93 12325
rect 145 12273 201 12325
rect 253 12273 309 12325
rect 361 12273 1145 12325
rect 43 12217 1145 12273
rect 43 12165 93 12217
rect 145 12165 201 12217
rect 253 12165 309 12217
rect 361 12165 1145 12217
rect 43 12109 1145 12165
rect 43 12057 93 12109
rect 145 12057 201 12109
rect 253 12057 309 12109
rect 361 12057 1145 12109
rect 43 12001 1145 12057
rect 43 11949 93 12001
rect 145 11949 201 12001
rect 253 11949 309 12001
rect 361 11949 1145 12001
rect 43 11893 1145 11949
rect 43 11841 93 11893
rect 145 11841 201 11893
rect 253 11841 309 11893
rect 361 11841 1145 11893
rect 43 11785 1145 11841
rect 43 11733 93 11785
rect 145 11733 201 11785
rect 253 11733 309 11785
rect 361 11733 1145 11785
rect 43 11677 1145 11733
rect 43 11625 93 11677
rect 145 11625 201 11677
rect 253 11625 309 11677
rect 361 11625 1145 11677
rect 43 11569 1145 11625
rect 43 11517 93 11569
rect 145 11517 201 11569
rect 253 11517 309 11569
rect 361 11517 1145 11569
rect 43 11461 1145 11517
rect 43 11409 93 11461
rect 145 11409 201 11461
rect 253 11409 309 11461
rect 361 11409 1145 11461
rect 43 11353 1145 11409
rect 43 11301 93 11353
rect 145 11301 201 11353
rect 253 11301 309 11353
rect 361 11301 1145 11353
rect 43 11245 1145 11301
rect 43 11193 93 11245
rect 145 11193 201 11245
rect 253 11193 309 11245
rect 361 11193 1145 11245
rect 43 11137 1145 11193
rect 43 11085 93 11137
rect 145 11085 201 11137
rect 253 11085 309 11137
rect 361 11085 1145 11137
rect 43 11029 1145 11085
rect 43 10977 93 11029
rect 145 10977 201 11029
rect 253 10977 309 11029
rect 361 10977 1145 11029
rect 43 10921 1145 10977
rect 43 10869 93 10921
rect 145 10869 201 10921
rect 253 10869 309 10921
rect 361 10869 1145 10921
rect 43 10813 1145 10869
rect 43 10761 93 10813
rect 145 10761 201 10813
rect 253 10761 309 10813
rect 361 10761 1145 10813
rect 43 10705 1145 10761
rect 43 10653 93 10705
rect 145 10653 201 10705
rect 253 10653 309 10705
rect 361 10653 1145 10705
rect 43 10597 1145 10653
rect 43 10545 93 10597
rect 145 10545 201 10597
rect 253 10545 309 10597
rect 361 10545 1145 10597
rect 43 10489 1145 10545
rect 43 10437 93 10489
rect 145 10437 201 10489
rect 253 10437 309 10489
rect 361 10437 1145 10489
rect 43 10381 1145 10437
rect 43 10329 93 10381
rect 145 10329 201 10381
rect 253 10329 309 10381
rect 361 10329 1145 10381
rect 43 10273 1145 10329
rect 43 10221 93 10273
rect 145 10221 201 10273
rect 253 10221 309 10273
rect 361 10221 1145 10273
rect 43 10165 1145 10221
rect 43 10113 93 10165
rect 145 10113 201 10165
rect 253 10113 309 10165
rect 361 10113 1145 10165
rect 43 10057 1145 10113
rect 43 10005 93 10057
rect 145 10005 201 10057
rect 253 10005 309 10057
rect 361 10005 1145 10057
rect 43 9949 1145 10005
rect 43 9897 93 9949
rect 145 9897 201 9949
rect 253 9897 309 9949
rect 361 9897 1145 9949
rect 43 9841 1145 9897
rect 43 9789 93 9841
rect 145 9789 201 9841
rect 253 9789 309 9841
rect 361 9789 1145 9841
rect 43 9733 1145 9789
rect 43 9681 93 9733
rect 145 9681 201 9733
rect 253 9681 309 9733
rect 361 9681 1145 9733
rect 43 9625 1145 9681
rect 43 9573 93 9625
rect 145 9573 201 9625
rect 253 9573 309 9625
rect 361 9573 1145 9625
rect 43 9517 1145 9573
rect 43 9465 93 9517
rect 145 9465 201 9517
rect 253 9465 309 9517
rect 361 9465 1145 9517
rect 43 9409 1145 9465
rect 43 9357 93 9409
rect 145 9357 201 9409
rect 253 9357 309 9409
rect 361 9357 1145 9409
rect 43 9301 1145 9357
rect 43 9249 93 9301
rect 145 9249 201 9301
rect 253 9249 309 9301
rect 361 9249 1145 9301
rect 43 9193 1145 9249
rect 43 9141 93 9193
rect 145 9141 201 9193
rect 253 9141 309 9193
rect 361 9141 1145 9193
rect 43 9085 1145 9141
rect 43 9033 93 9085
rect 145 9033 201 9085
rect 253 9033 309 9085
rect 361 9033 1145 9085
rect 43 8977 1145 9033
rect 43 8925 93 8977
rect 145 8925 201 8977
rect 253 8925 309 8977
rect 361 8925 1145 8977
rect 43 8869 1145 8925
rect 43 8817 93 8869
rect 145 8817 201 8869
rect 253 8817 309 8869
rect 361 8817 1145 8869
rect 43 8761 1145 8817
rect 43 8709 93 8761
rect 145 8709 201 8761
rect 253 8709 309 8761
rect 361 8709 1145 8761
rect 43 8653 1145 8709
rect 43 8601 93 8653
rect 145 8601 201 8653
rect 253 8601 309 8653
rect 361 8601 1145 8653
rect 43 8545 1145 8601
rect 43 8493 93 8545
rect 145 8493 201 8545
rect 253 8493 309 8545
rect 361 8493 1145 8545
rect 43 8437 1145 8493
rect 43 8385 93 8437
rect 145 8385 201 8437
rect 253 8385 309 8437
rect 361 8385 1145 8437
rect 43 8329 1145 8385
rect 43 8277 93 8329
rect 145 8277 201 8329
rect 253 8277 309 8329
rect 361 8277 1145 8329
rect 43 8221 1145 8277
rect 43 8169 93 8221
rect 145 8169 201 8221
rect 253 8169 309 8221
rect 361 8169 1145 8221
rect 43 8113 1145 8169
rect 43 8061 93 8113
rect 145 8061 201 8113
rect 253 8061 309 8113
rect 361 8061 1145 8113
rect 43 8005 1145 8061
rect 43 7953 93 8005
rect 145 7953 201 8005
rect 253 7953 309 8005
rect 361 7953 1145 8005
rect 43 7897 1145 7953
rect 43 7845 93 7897
rect 145 7845 201 7897
rect 253 7845 309 7897
rect 361 7845 1145 7897
rect 43 7789 1145 7845
rect 43 7737 93 7789
rect 145 7737 201 7789
rect 253 7737 309 7789
rect 361 7737 1145 7789
rect 43 7681 1145 7737
rect 43 7629 93 7681
rect 145 7629 201 7681
rect 253 7629 309 7681
rect 361 7629 1145 7681
rect 43 7573 1145 7629
rect 43 7521 93 7573
rect 145 7521 201 7573
rect 253 7521 309 7573
rect 361 7521 1145 7573
rect 43 7465 1145 7521
rect 43 7413 93 7465
rect 145 7413 201 7465
rect 253 7413 309 7465
rect 361 7413 1145 7465
rect 43 7357 1145 7413
rect 43 7305 93 7357
rect 145 7305 201 7357
rect 253 7305 309 7357
rect 361 7305 1145 7357
rect 43 7249 1145 7305
rect 43 7197 93 7249
rect 145 7197 201 7249
rect 253 7197 309 7249
rect 361 7197 1145 7249
rect 43 7141 1145 7197
rect 43 7089 93 7141
rect 145 7089 201 7141
rect 253 7089 309 7141
rect 361 7089 1145 7141
rect 43 7033 1145 7089
rect 43 6981 93 7033
rect 145 6981 201 7033
rect 253 6981 309 7033
rect 361 6981 1145 7033
rect 43 6925 1145 6981
rect 43 6873 93 6925
rect 145 6873 201 6925
rect 253 6873 309 6925
rect 361 6873 1145 6925
rect 43 6817 1145 6873
rect 43 6765 93 6817
rect 145 6765 201 6817
rect 253 6765 309 6817
rect 361 6765 1145 6817
rect 43 6709 1145 6765
rect 43 6657 93 6709
rect 145 6657 201 6709
rect 253 6657 309 6709
rect 361 6657 1145 6709
rect 43 6601 1145 6657
rect 43 6549 93 6601
rect 145 6549 201 6601
rect 253 6549 309 6601
rect 361 6549 1145 6601
rect 43 6493 1145 6549
rect 43 6441 93 6493
rect 145 6441 201 6493
rect 253 6441 309 6493
rect 361 6441 1145 6493
rect 43 6385 1145 6441
rect 43 6333 93 6385
rect 145 6333 201 6385
rect 253 6333 309 6385
rect 361 6333 1145 6385
rect 43 6277 1145 6333
rect 43 6225 93 6277
rect 145 6225 201 6277
rect 253 6225 309 6277
rect 361 6225 1145 6277
rect 43 6169 1145 6225
rect 43 6117 93 6169
rect 145 6117 201 6169
rect 253 6117 309 6169
rect 361 6117 1145 6169
rect 43 6061 1145 6117
rect 43 6009 93 6061
rect 145 6009 201 6061
rect 253 6009 309 6061
rect 361 6009 1145 6061
rect 43 5953 1145 6009
rect 43 5901 93 5953
rect 145 5901 201 5953
rect 253 5901 309 5953
rect 361 5901 1145 5953
rect 43 5845 1145 5901
rect 43 5793 93 5845
rect 145 5793 201 5845
rect 253 5793 309 5845
rect 361 5793 1145 5845
rect 43 5737 1145 5793
rect 43 5685 93 5737
rect 145 5685 201 5737
rect 253 5685 309 5737
rect 361 5685 1145 5737
rect 43 5629 1145 5685
rect 43 5577 93 5629
rect 145 5577 201 5629
rect 253 5577 309 5629
rect 361 5577 1145 5629
rect 43 5521 1145 5577
rect 43 5469 93 5521
rect 145 5469 201 5521
rect 253 5469 309 5521
rect 361 5469 1145 5521
rect 43 5413 1145 5469
rect 43 5361 93 5413
rect 145 5361 201 5413
rect 253 5361 309 5413
rect 361 5361 1145 5413
rect 43 5305 1145 5361
rect 43 5253 93 5305
rect 145 5253 201 5305
rect 253 5253 309 5305
rect 361 5253 1145 5305
rect 43 5197 1145 5253
rect 43 5145 93 5197
rect 145 5145 201 5197
rect 253 5145 309 5197
rect 361 5145 1145 5197
rect 43 5089 1145 5145
rect 43 5037 93 5089
rect 145 5037 201 5089
rect 253 5037 309 5089
rect 361 5037 1145 5089
rect 43 4981 1145 5037
rect 43 4929 93 4981
rect 145 4929 201 4981
rect 253 4929 309 4981
rect 361 4929 1145 4981
rect 43 4873 1145 4929
rect 43 4821 93 4873
rect 145 4821 201 4873
rect 253 4821 309 4873
rect 361 4821 1145 4873
rect 43 4765 1145 4821
rect 43 4713 93 4765
rect 145 4713 201 4765
rect 253 4713 309 4765
rect 361 4713 1145 4765
rect 43 4657 1145 4713
rect 43 4605 93 4657
rect 145 4605 201 4657
rect 253 4605 309 4657
rect 361 4605 1145 4657
rect 43 4549 1145 4605
rect 43 4497 93 4549
rect 145 4497 201 4549
rect 253 4497 309 4549
rect 361 4497 1145 4549
rect 43 4441 1145 4497
rect 43 4389 93 4441
rect 145 4389 201 4441
rect 253 4389 309 4441
rect 361 4389 1145 4441
rect 43 4333 1145 4389
rect 43 4281 93 4333
rect 145 4281 201 4333
rect 253 4281 309 4333
rect 361 4281 1145 4333
rect 43 4225 1145 4281
rect 43 4173 93 4225
rect 145 4173 201 4225
rect 253 4173 309 4225
rect 361 4173 1145 4225
rect 43 4117 1145 4173
rect 43 4065 93 4117
rect 145 4065 201 4117
rect 253 4065 309 4117
rect 361 4065 1145 4117
rect 43 4009 1145 4065
rect 43 3957 93 4009
rect 145 3957 201 4009
rect 253 3957 309 4009
rect 361 3957 1145 4009
rect 43 3901 1145 3957
rect 43 3849 93 3901
rect 145 3849 201 3901
rect 253 3849 309 3901
rect 361 3849 1145 3901
rect 43 3793 1145 3849
rect 43 3741 93 3793
rect 145 3741 201 3793
rect 253 3741 309 3793
rect 361 3741 1145 3793
rect 43 3685 1145 3741
rect 43 3633 93 3685
rect 145 3633 201 3685
rect 253 3633 309 3685
rect 361 3633 1145 3685
rect 43 3577 1145 3633
rect 43 3525 93 3577
rect 145 3525 201 3577
rect 253 3525 309 3577
rect 361 3525 1145 3577
rect 43 3469 1145 3525
rect 43 3417 93 3469
rect 145 3417 201 3469
rect 253 3417 309 3469
rect 361 3417 1145 3469
rect 43 3361 1145 3417
rect 43 3309 93 3361
rect 145 3309 201 3361
rect 253 3309 309 3361
rect 361 3309 1145 3361
rect 43 3253 1145 3309
rect 43 3201 93 3253
rect 145 3201 201 3253
rect 253 3201 309 3253
rect 361 3201 1145 3253
rect 43 3145 1145 3201
rect 43 3093 93 3145
rect 145 3093 201 3145
rect 253 3093 309 3145
rect 361 3093 1145 3145
rect 43 3037 1145 3093
rect 43 2985 93 3037
rect 145 2985 201 3037
rect 253 2985 309 3037
rect 361 2985 1145 3037
rect 43 2929 1145 2985
rect 43 2877 93 2929
rect 145 2877 201 2929
rect 253 2877 309 2929
rect 361 2877 1145 2929
rect 43 2821 1145 2877
rect 43 2769 93 2821
rect 145 2769 201 2821
rect 253 2769 309 2821
rect 361 2769 1145 2821
rect 43 2713 1145 2769
rect 43 2661 93 2713
rect 145 2661 201 2713
rect 253 2661 309 2713
rect 361 2661 1145 2713
rect 43 2605 1145 2661
rect 43 2553 93 2605
rect 145 2553 201 2605
rect 253 2553 309 2605
rect 361 2553 1145 2605
rect 43 2497 1145 2553
rect 43 2445 93 2497
rect 145 2445 201 2497
rect 253 2445 309 2497
rect 361 2445 1145 2497
rect 43 2389 1145 2445
rect 43 2337 93 2389
rect 145 2337 201 2389
rect 253 2337 309 2389
rect 361 2337 1145 2389
rect 43 2281 1145 2337
rect 43 2229 93 2281
rect 145 2229 201 2281
rect 253 2229 309 2281
rect 361 2229 1145 2281
rect 43 2173 1145 2229
rect 43 2121 93 2173
rect 145 2121 201 2173
rect 253 2121 309 2173
rect 361 2121 1145 2173
rect 43 2065 1145 2121
rect 43 2013 93 2065
rect 145 2013 201 2065
rect 253 2013 309 2065
rect 361 2013 1145 2065
rect 43 1957 1145 2013
rect 43 1905 93 1957
rect 145 1905 201 1957
rect 253 1905 309 1957
rect 361 1905 1145 1957
rect 43 1849 1145 1905
rect 43 1797 93 1849
rect 145 1797 201 1849
rect 253 1797 309 1849
rect 361 1797 1145 1849
rect 43 1741 1145 1797
rect 43 1689 93 1741
rect 145 1689 201 1741
rect 253 1689 309 1741
rect 361 1689 1145 1741
rect 43 1633 1145 1689
rect 43 1581 93 1633
rect 145 1581 201 1633
rect 253 1581 309 1633
rect 361 1581 1145 1633
rect 43 1525 1145 1581
rect 43 1473 93 1525
rect 145 1473 201 1525
rect 253 1473 309 1525
rect 361 1473 1145 1525
rect 43 1417 1145 1473
rect 1213 23887 1413 25617
rect 1213 23835 1233 23887
rect 1285 23835 1341 23887
rect 1393 23835 1413 23887
rect 1213 23779 1413 23835
rect 1213 23727 1233 23779
rect 1285 23727 1341 23779
rect 1393 23727 1413 23779
rect 1213 23671 1413 23727
rect 1213 23619 1233 23671
rect 1285 23619 1341 23671
rect 1393 23619 1413 23671
rect 1213 23563 1413 23619
rect 1213 23511 1233 23563
rect 1285 23511 1341 23563
rect 1393 23511 1413 23563
rect 1213 23455 1413 23511
rect 1213 23403 1233 23455
rect 1285 23403 1341 23455
rect 1393 23403 1413 23455
rect 1213 23347 1413 23403
rect 1213 23295 1233 23347
rect 1285 23295 1341 23347
rect 1393 23295 1413 23347
rect 1213 23239 1413 23295
rect 1213 23187 1233 23239
rect 1285 23187 1341 23239
rect 1393 23187 1413 23239
rect 1213 23131 1413 23187
rect 1213 23079 1233 23131
rect 1285 23079 1341 23131
rect 1393 23079 1413 23131
rect 1213 23023 1413 23079
rect 1213 22971 1233 23023
rect 1285 22971 1341 23023
rect 1393 22971 1413 23023
rect 1213 22915 1413 22971
rect 1213 22863 1233 22915
rect 1285 22863 1341 22915
rect 1393 22863 1413 22915
rect 1213 22807 1413 22863
rect 1213 22755 1233 22807
rect 1285 22755 1341 22807
rect 1393 22755 1413 22807
rect 1213 22699 1413 22755
rect 1213 22647 1233 22699
rect 1285 22647 1341 22699
rect 1393 22647 1413 22699
rect 1213 22591 1413 22647
rect 1213 22539 1233 22591
rect 1285 22539 1341 22591
rect 1393 22539 1413 22591
rect 1213 22483 1413 22539
rect 1213 22431 1233 22483
rect 1285 22431 1341 22483
rect 1393 22431 1413 22483
rect 1213 22375 1413 22431
rect 1213 22323 1233 22375
rect 1285 22323 1341 22375
rect 1393 22323 1413 22375
rect 1213 22267 1413 22323
rect 1213 22215 1233 22267
rect 1285 22215 1341 22267
rect 1393 22215 1413 22267
rect 1213 22159 1413 22215
rect 1213 22107 1233 22159
rect 1285 22107 1341 22159
rect 1393 22107 1413 22159
rect 1213 22051 1413 22107
rect 1213 21999 1233 22051
rect 1285 21999 1341 22051
rect 1393 21999 1413 22051
rect 1213 21943 1413 21999
rect 1213 21891 1233 21943
rect 1285 21891 1341 21943
rect 1393 21891 1413 21943
rect 1213 21835 1413 21891
rect 1213 21783 1233 21835
rect 1285 21783 1341 21835
rect 1393 21783 1413 21835
rect 1213 21727 1413 21783
rect 1213 21675 1233 21727
rect 1285 21675 1341 21727
rect 1393 21675 1413 21727
rect 1213 21619 1413 21675
rect 1213 21567 1233 21619
rect 1285 21567 1341 21619
rect 1393 21567 1413 21619
rect 1213 21511 1413 21567
rect 1213 21459 1233 21511
rect 1285 21459 1341 21511
rect 1393 21459 1413 21511
rect 1213 21403 1413 21459
rect 1213 21351 1233 21403
rect 1285 21351 1341 21403
rect 1393 21351 1413 21403
rect 1213 21295 1413 21351
rect 1213 21243 1233 21295
rect 1285 21243 1341 21295
rect 1393 21243 1413 21295
rect 1213 21187 1413 21243
rect 1213 21135 1233 21187
rect 1285 21135 1341 21187
rect 1393 21135 1413 21187
rect 1213 21079 1413 21135
rect 1213 21027 1233 21079
rect 1285 21027 1341 21079
rect 1393 21027 1413 21079
rect 1213 20971 1413 21027
rect 1213 20919 1233 20971
rect 1285 20919 1341 20971
rect 1393 20919 1413 20971
rect 1213 20863 1413 20919
rect 1213 20811 1233 20863
rect 1285 20811 1341 20863
rect 1393 20811 1413 20863
rect 1213 20755 1413 20811
rect 1213 20703 1233 20755
rect 1285 20703 1341 20755
rect 1393 20703 1413 20755
rect 1213 20647 1413 20703
rect 1213 20595 1233 20647
rect 1285 20595 1341 20647
rect 1393 20595 1413 20647
rect 1213 20539 1413 20595
rect 1213 20487 1233 20539
rect 1285 20487 1341 20539
rect 1393 20487 1413 20539
rect 1213 20431 1413 20487
rect 1213 20379 1233 20431
rect 1285 20379 1341 20431
rect 1393 20379 1413 20431
rect 1213 20323 1413 20379
rect 1213 20271 1233 20323
rect 1285 20271 1341 20323
rect 1393 20271 1413 20323
rect 1213 20215 1413 20271
rect 1213 20163 1233 20215
rect 1285 20163 1341 20215
rect 1393 20163 1413 20215
rect 1213 20107 1413 20163
rect 1213 20055 1233 20107
rect 1285 20055 1341 20107
rect 1393 20055 1413 20107
rect 1213 19999 1413 20055
rect 1213 19947 1233 19999
rect 1285 19947 1341 19999
rect 1393 19947 1413 19999
rect 1213 19891 1413 19947
rect 1213 19839 1233 19891
rect 1285 19839 1341 19891
rect 1393 19839 1413 19891
rect 1213 19783 1413 19839
rect 1213 19731 1233 19783
rect 1285 19731 1341 19783
rect 1393 19731 1413 19783
rect 1213 19675 1413 19731
rect 1213 19623 1233 19675
rect 1285 19623 1341 19675
rect 1393 19623 1413 19675
rect 1213 19567 1413 19623
rect 1213 19515 1233 19567
rect 1285 19515 1341 19567
rect 1393 19515 1413 19567
rect 1213 19459 1413 19515
rect 1213 19407 1233 19459
rect 1285 19407 1341 19459
rect 1393 19407 1413 19459
rect 1213 19351 1413 19407
rect 1213 19299 1233 19351
rect 1285 19299 1341 19351
rect 1393 19299 1413 19351
rect 1213 19243 1413 19299
rect 1213 19191 1233 19243
rect 1285 19191 1341 19243
rect 1393 19191 1413 19243
rect 1213 19135 1413 19191
rect 1213 19083 1233 19135
rect 1285 19083 1341 19135
rect 1393 19083 1413 19135
rect 1213 18015 1413 19083
rect 1213 17963 1233 18015
rect 1285 17963 1341 18015
rect 1393 17963 1413 18015
rect 1213 17907 1413 17963
rect 1213 17855 1233 17907
rect 1285 17855 1341 17907
rect 1393 17855 1413 17907
rect 1213 17799 1413 17855
rect 1213 17747 1233 17799
rect 1285 17747 1341 17799
rect 1393 17747 1413 17799
rect 1213 17691 1413 17747
rect 1213 17639 1233 17691
rect 1285 17639 1341 17691
rect 1393 17639 1413 17691
rect 1213 17583 1413 17639
rect 1213 17531 1233 17583
rect 1285 17531 1341 17583
rect 1393 17531 1413 17583
rect 1213 17475 1413 17531
rect 1213 17423 1233 17475
rect 1285 17423 1341 17475
rect 1393 17423 1413 17475
rect 1213 17367 1413 17423
rect 1213 17315 1233 17367
rect 1285 17315 1341 17367
rect 1393 17315 1413 17367
rect 1213 17259 1413 17315
rect 1213 17207 1233 17259
rect 1285 17207 1341 17259
rect 1393 17207 1413 17259
rect 1213 17151 1413 17207
rect 1213 17099 1233 17151
rect 1285 17099 1341 17151
rect 1393 17099 1413 17151
rect 1213 17043 1413 17099
rect 1213 16991 1233 17043
rect 1285 16991 1341 17043
rect 1393 16991 1413 17043
rect 1213 16935 1413 16991
rect 1213 16883 1233 16935
rect 1285 16883 1341 16935
rect 1393 16883 1413 16935
rect 1213 16827 1413 16883
rect 1213 16775 1233 16827
rect 1285 16775 1341 16827
rect 1393 16775 1413 16827
rect 1213 16719 1413 16775
rect 1213 16667 1233 16719
rect 1285 16667 1341 16719
rect 1393 16667 1413 16719
rect 1213 16611 1413 16667
rect 1213 16559 1233 16611
rect 1285 16559 1341 16611
rect 1393 16559 1413 16611
rect 1213 16503 1413 16559
rect 1213 16451 1233 16503
rect 1285 16451 1341 16503
rect 1393 16451 1413 16503
rect 1213 16395 1413 16451
rect 1213 16343 1233 16395
rect 1285 16343 1341 16395
rect 1393 16343 1413 16395
rect 1213 16287 1413 16343
rect 1213 16235 1233 16287
rect 1285 16235 1341 16287
rect 1393 16235 1413 16287
rect 1213 16179 1413 16235
rect 1213 16127 1233 16179
rect 1285 16127 1341 16179
rect 1393 16127 1413 16179
rect 1213 16071 1413 16127
rect 1213 16019 1233 16071
rect 1285 16019 1341 16071
rect 1393 16019 1413 16071
rect 1213 15963 1413 16019
rect 1213 15911 1233 15963
rect 1285 15911 1341 15963
rect 1393 15911 1413 15963
rect 1213 15855 1413 15911
rect 1213 15803 1233 15855
rect 1285 15803 1341 15855
rect 1393 15803 1413 15855
rect 1213 15747 1413 15803
rect 1213 15695 1233 15747
rect 1285 15695 1341 15747
rect 1393 15695 1413 15747
rect 1213 15639 1413 15695
rect 1213 15587 1233 15639
rect 1285 15587 1341 15639
rect 1393 15587 1413 15639
rect 1213 15531 1413 15587
rect 1213 15479 1233 15531
rect 1285 15479 1341 15531
rect 1393 15479 1413 15531
rect 1213 15423 1413 15479
rect 1213 15371 1233 15423
rect 1285 15371 1341 15423
rect 1393 15371 1413 15423
rect 1213 15315 1413 15371
rect 1213 15263 1233 15315
rect 1285 15263 1341 15315
rect 1393 15263 1413 15315
rect 1213 15207 1413 15263
rect 1213 15155 1233 15207
rect 1285 15155 1341 15207
rect 1393 15155 1413 15207
rect 1213 15099 1413 15155
rect 1213 15047 1233 15099
rect 1285 15047 1341 15099
rect 1393 15047 1413 15099
rect 1213 14991 1413 15047
rect 1213 14939 1233 14991
rect 1285 14939 1341 14991
rect 1393 14939 1413 14991
rect 1213 14883 1413 14939
rect 1213 14831 1233 14883
rect 1285 14831 1341 14883
rect 1393 14831 1413 14883
rect 1213 14775 1413 14831
rect 1213 14723 1233 14775
rect 1285 14723 1341 14775
rect 1393 14723 1413 14775
rect 1213 14667 1413 14723
rect 1213 14615 1233 14667
rect 1285 14615 1341 14667
rect 1393 14615 1413 14667
rect 1213 14559 1413 14615
rect 1213 14507 1233 14559
rect 1285 14507 1341 14559
rect 1393 14507 1413 14559
rect 1213 14451 1413 14507
rect 1213 14399 1233 14451
rect 1285 14399 1341 14451
rect 1393 14399 1413 14451
rect 1213 14343 1413 14399
rect 1213 14291 1233 14343
rect 1285 14291 1341 14343
rect 1393 14291 1413 14343
rect 1213 14235 1413 14291
rect 1213 14183 1233 14235
rect 1285 14183 1341 14235
rect 1393 14183 1413 14235
rect 1213 14127 1413 14183
rect 1213 14075 1233 14127
rect 1285 14075 1341 14127
rect 1393 14075 1413 14127
rect 1213 14019 1413 14075
rect 1213 13967 1233 14019
rect 1285 13967 1341 14019
rect 1393 13967 1413 14019
rect 1213 13911 1413 13967
rect 1213 13859 1233 13911
rect 1285 13859 1341 13911
rect 1393 13859 1413 13911
rect 1213 13803 1413 13859
rect 1213 13751 1233 13803
rect 1285 13751 1341 13803
rect 1393 13751 1413 13803
rect 1213 13695 1413 13751
rect 1213 13643 1233 13695
rect 1285 13643 1341 13695
rect 1393 13643 1413 13695
rect 1213 13587 1413 13643
rect 1213 13535 1233 13587
rect 1285 13535 1341 13587
rect 1393 13535 1413 13587
rect 1213 13479 1413 13535
rect 1213 13427 1233 13479
rect 1285 13427 1341 13479
rect 1393 13427 1413 13479
rect 1213 13371 1413 13427
rect 1213 13319 1233 13371
rect 1285 13319 1341 13371
rect 1393 13319 1413 13371
rect 1213 13263 1413 13319
rect 1213 13211 1233 13263
rect 1285 13211 1341 13263
rect 1393 13211 1413 13263
rect 1213 12143 1413 13211
rect 1213 12091 1233 12143
rect 1285 12091 1341 12143
rect 1393 12091 1413 12143
rect 1213 12035 1413 12091
rect 1213 11983 1233 12035
rect 1285 11983 1341 12035
rect 1393 11983 1413 12035
rect 1213 11927 1413 11983
rect 1213 11875 1233 11927
rect 1285 11875 1341 11927
rect 1393 11875 1413 11927
rect 1213 11819 1413 11875
rect 1213 11767 1233 11819
rect 1285 11767 1341 11819
rect 1393 11767 1413 11819
rect 1213 11711 1413 11767
rect 1213 11659 1233 11711
rect 1285 11659 1341 11711
rect 1393 11659 1413 11711
rect 1213 11603 1413 11659
rect 1213 11551 1233 11603
rect 1285 11551 1341 11603
rect 1393 11551 1413 11603
rect 1213 11495 1413 11551
rect 1213 11443 1233 11495
rect 1285 11443 1341 11495
rect 1393 11443 1413 11495
rect 1213 11387 1413 11443
rect 1213 11335 1233 11387
rect 1285 11335 1341 11387
rect 1393 11335 1413 11387
rect 1213 11279 1413 11335
rect 1213 11227 1233 11279
rect 1285 11227 1341 11279
rect 1393 11227 1413 11279
rect 1213 11171 1413 11227
rect 1213 11119 1233 11171
rect 1285 11119 1341 11171
rect 1393 11119 1413 11171
rect 1213 11063 1413 11119
rect 1213 11011 1233 11063
rect 1285 11011 1341 11063
rect 1393 11011 1413 11063
rect 1213 10955 1413 11011
rect 1213 10903 1233 10955
rect 1285 10903 1341 10955
rect 1393 10903 1413 10955
rect 1213 10847 1413 10903
rect 1213 10795 1233 10847
rect 1285 10795 1341 10847
rect 1393 10795 1413 10847
rect 1213 10739 1413 10795
rect 1213 10687 1233 10739
rect 1285 10687 1341 10739
rect 1393 10687 1413 10739
rect 1213 10631 1413 10687
rect 1213 10579 1233 10631
rect 1285 10579 1341 10631
rect 1393 10579 1413 10631
rect 1213 10523 1413 10579
rect 1213 10471 1233 10523
rect 1285 10471 1341 10523
rect 1393 10471 1413 10523
rect 1213 10415 1413 10471
rect 1213 10363 1233 10415
rect 1285 10363 1341 10415
rect 1393 10363 1413 10415
rect 1213 10307 1413 10363
rect 1213 10255 1233 10307
rect 1285 10255 1341 10307
rect 1393 10255 1413 10307
rect 1213 10199 1413 10255
rect 1213 10147 1233 10199
rect 1285 10147 1341 10199
rect 1393 10147 1413 10199
rect 1213 10091 1413 10147
rect 1213 10039 1233 10091
rect 1285 10039 1341 10091
rect 1393 10039 1413 10091
rect 1213 9983 1413 10039
rect 1213 9931 1233 9983
rect 1285 9931 1341 9983
rect 1393 9931 1413 9983
rect 1213 9875 1413 9931
rect 1213 9823 1233 9875
rect 1285 9823 1341 9875
rect 1393 9823 1413 9875
rect 1213 9767 1413 9823
rect 1213 9715 1233 9767
rect 1285 9715 1341 9767
rect 1393 9715 1413 9767
rect 1213 9659 1413 9715
rect 1213 9607 1233 9659
rect 1285 9607 1341 9659
rect 1393 9607 1413 9659
rect 1213 9551 1413 9607
rect 1213 9499 1233 9551
rect 1285 9499 1341 9551
rect 1393 9499 1413 9551
rect 1213 9443 1413 9499
rect 1213 9391 1233 9443
rect 1285 9391 1341 9443
rect 1393 9391 1413 9443
rect 1213 9335 1413 9391
rect 1213 9283 1233 9335
rect 1285 9283 1341 9335
rect 1393 9283 1413 9335
rect 1213 9227 1413 9283
rect 1213 9175 1233 9227
rect 1285 9175 1341 9227
rect 1393 9175 1413 9227
rect 1213 9119 1413 9175
rect 1213 9067 1233 9119
rect 1285 9067 1341 9119
rect 1393 9067 1413 9119
rect 1213 9011 1413 9067
rect 1213 8959 1233 9011
rect 1285 8959 1341 9011
rect 1393 8959 1413 9011
rect 1213 8903 1413 8959
rect 1213 8851 1233 8903
rect 1285 8851 1341 8903
rect 1393 8851 1413 8903
rect 1213 8795 1413 8851
rect 1213 8743 1233 8795
rect 1285 8743 1341 8795
rect 1393 8743 1413 8795
rect 1213 8687 1413 8743
rect 1213 8635 1233 8687
rect 1285 8635 1341 8687
rect 1393 8635 1413 8687
rect 1213 8579 1413 8635
rect 1213 8527 1233 8579
rect 1285 8527 1341 8579
rect 1393 8527 1413 8579
rect 1213 8471 1413 8527
rect 1213 8419 1233 8471
rect 1285 8419 1341 8471
rect 1393 8419 1413 8471
rect 1213 8363 1413 8419
rect 1213 8311 1233 8363
rect 1285 8311 1341 8363
rect 1393 8311 1413 8363
rect 1213 8255 1413 8311
rect 1213 8203 1233 8255
rect 1285 8203 1341 8255
rect 1393 8203 1413 8255
rect 1213 8147 1413 8203
rect 1213 8095 1233 8147
rect 1285 8095 1341 8147
rect 1393 8095 1413 8147
rect 1213 8039 1413 8095
rect 1213 7987 1233 8039
rect 1285 7987 1341 8039
rect 1393 7987 1413 8039
rect 1213 7931 1413 7987
rect 1213 7879 1233 7931
rect 1285 7879 1341 7931
rect 1393 7879 1413 7931
rect 1213 7823 1413 7879
rect 1213 7771 1233 7823
rect 1285 7771 1341 7823
rect 1393 7771 1413 7823
rect 1213 7715 1413 7771
rect 1213 7663 1233 7715
rect 1285 7663 1341 7715
rect 1393 7663 1413 7715
rect 1213 7607 1413 7663
rect 1213 7555 1233 7607
rect 1285 7555 1341 7607
rect 1393 7555 1413 7607
rect 1213 7499 1413 7555
rect 1213 7447 1233 7499
rect 1285 7447 1341 7499
rect 1393 7447 1413 7499
rect 1213 7391 1413 7447
rect 1213 7339 1233 7391
rect 1285 7339 1341 7391
rect 1393 7339 1413 7391
rect 1213 6271 1413 7339
rect 1213 6219 1233 6271
rect 1285 6219 1341 6271
rect 1393 6219 1413 6271
rect 1213 6163 1413 6219
rect 1213 6111 1233 6163
rect 1285 6111 1341 6163
rect 1393 6111 1413 6163
rect 1213 6055 1413 6111
rect 1213 6003 1233 6055
rect 1285 6003 1341 6055
rect 1393 6003 1413 6055
rect 1213 5947 1413 6003
rect 1213 5895 1233 5947
rect 1285 5895 1341 5947
rect 1393 5895 1413 5947
rect 1213 5839 1413 5895
rect 1213 5787 1233 5839
rect 1285 5787 1341 5839
rect 1393 5787 1413 5839
rect 1213 5731 1413 5787
rect 1213 5679 1233 5731
rect 1285 5679 1341 5731
rect 1393 5679 1413 5731
rect 1213 5623 1413 5679
rect 1213 5571 1233 5623
rect 1285 5571 1341 5623
rect 1393 5571 1413 5623
rect 1213 5515 1413 5571
rect 1213 5463 1233 5515
rect 1285 5463 1341 5515
rect 1393 5463 1413 5515
rect 1213 5407 1413 5463
rect 1213 5355 1233 5407
rect 1285 5355 1341 5407
rect 1393 5355 1413 5407
rect 1213 5299 1413 5355
rect 1213 5247 1233 5299
rect 1285 5247 1341 5299
rect 1393 5247 1413 5299
rect 1213 5191 1413 5247
rect 1213 5139 1233 5191
rect 1285 5139 1341 5191
rect 1393 5139 1413 5191
rect 1213 5083 1413 5139
rect 1213 5031 1233 5083
rect 1285 5031 1341 5083
rect 1393 5031 1413 5083
rect 1213 4975 1413 5031
rect 1213 4923 1233 4975
rect 1285 4923 1341 4975
rect 1393 4923 1413 4975
rect 1213 4867 1413 4923
rect 1213 4815 1233 4867
rect 1285 4815 1341 4867
rect 1393 4815 1413 4867
rect 1213 4759 1413 4815
rect 1213 4707 1233 4759
rect 1285 4707 1341 4759
rect 1393 4707 1413 4759
rect 1213 4651 1413 4707
rect 1213 4599 1233 4651
rect 1285 4599 1341 4651
rect 1393 4599 1413 4651
rect 1213 4543 1413 4599
rect 1213 4491 1233 4543
rect 1285 4491 1341 4543
rect 1393 4491 1413 4543
rect 1213 4435 1413 4491
rect 1213 4383 1233 4435
rect 1285 4383 1341 4435
rect 1393 4383 1413 4435
rect 1213 4327 1413 4383
rect 1213 4275 1233 4327
rect 1285 4275 1341 4327
rect 1393 4275 1413 4327
rect 1213 4219 1413 4275
rect 1213 4167 1233 4219
rect 1285 4167 1341 4219
rect 1393 4167 1413 4219
rect 1213 4111 1413 4167
rect 1213 4059 1233 4111
rect 1285 4059 1341 4111
rect 1393 4059 1413 4111
rect 1213 4003 1413 4059
rect 1213 3951 1233 4003
rect 1285 3951 1341 4003
rect 1393 3951 1413 4003
rect 1213 3895 1413 3951
rect 1213 3843 1233 3895
rect 1285 3843 1341 3895
rect 1393 3843 1413 3895
rect 1213 3787 1413 3843
rect 1213 3735 1233 3787
rect 1285 3735 1341 3787
rect 1393 3735 1413 3787
rect 1213 3679 1413 3735
rect 1213 3627 1233 3679
rect 1285 3627 1341 3679
rect 1393 3627 1413 3679
rect 1213 3571 1413 3627
rect 1213 3519 1233 3571
rect 1285 3519 1341 3571
rect 1393 3519 1413 3571
rect 1213 3463 1413 3519
rect 1213 3411 1233 3463
rect 1285 3411 1341 3463
rect 1393 3411 1413 3463
rect 1213 3355 1413 3411
rect 1213 3303 1233 3355
rect 1285 3303 1341 3355
rect 1393 3303 1413 3355
rect 1213 3247 1413 3303
rect 1213 3195 1233 3247
rect 1285 3195 1341 3247
rect 1393 3195 1413 3247
rect 1213 3139 1413 3195
rect 1213 3087 1233 3139
rect 1285 3087 1341 3139
rect 1393 3087 1413 3139
rect 1213 3031 1413 3087
rect 1213 2979 1233 3031
rect 1285 2979 1341 3031
rect 1393 2979 1413 3031
rect 1213 2923 1413 2979
rect 1213 2871 1233 2923
rect 1285 2871 1341 2923
rect 1393 2871 1413 2923
rect 1213 2815 1413 2871
rect 1213 2763 1233 2815
rect 1285 2763 1341 2815
rect 1393 2763 1413 2815
rect 1213 2707 1413 2763
rect 1213 2655 1233 2707
rect 1285 2655 1341 2707
rect 1393 2655 1413 2707
rect 1213 2599 1413 2655
rect 1213 2547 1233 2599
rect 1285 2547 1341 2599
rect 1393 2547 1413 2599
rect 1213 2491 1413 2547
rect 1213 2439 1233 2491
rect 1285 2439 1341 2491
rect 1393 2439 1413 2491
rect 1213 2383 1413 2439
rect 1213 2331 1233 2383
rect 1285 2331 1341 2383
rect 1393 2331 1413 2383
rect 1213 2275 1413 2331
rect 1213 2223 1233 2275
rect 1285 2223 1341 2275
rect 1393 2223 1413 2275
rect 1213 2167 1413 2223
rect 1213 2115 1233 2167
rect 1285 2115 1341 2167
rect 1393 2115 1413 2167
rect 1213 2059 1413 2115
rect 1213 2007 1233 2059
rect 1285 2007 1341 2059
rect 1393 2007 1413 2059
rect 1213 1951 1413 2007
rect 1213 1899 1233 1951
rect 1285 1899 1341 1951
rect 1393 1899 1413 1951
rect 1213 1843 1413 1899
rect 1213 1791 1233 1843
rect 1285 1791 1341 1843
rect 1393 1791 1413 1843
rect 1213 1735 1413 1791
rect 1213 1683 1233 1735
rect 1285 1683 1341 1735
rect 1393 1683 1413 1735
rect 1213 1627 1413 1683
rect 1213 1575 1233 1627
rect 1285 1575 1341 1627
rect 1393 1575 1413 1627
rect 1213 1519 1413 1575
rect 1213 1467 1233 1519
rect 1285 1467 1341 1519
rect 1393 1467 1413 1519
rect 1213 1455 1413 1467
rect 1481 24661 3309 25617
rect 1481 24609 1505 24661
rect 1557 24609 1613 24661
rect 1665 24609 1721 24661
rect 1773 24609 1829 24661
rect 1881 24609 1937 24661
rect 1989 24609 2045 24661
rect 2097 24609 2153 24661
rect 2205 24609 2261 24661
rect 2313 24609 2369 24661
rect 2421 24609 2477 24661
rect 2529 24609 2585 24661
rect 2637 24609 2693 24661
rect 2745 24609 2801 24661
rect 2853 24609 2909 24661
rect 2961 24609 3017 24661
rect 3069 24609 3125 24661
rect 3177 24609 3233 24661
rect 3285 24609 3309 24661
rect 1481 24553 3309 24609
rect 1481 24501 1505 24553
rect 1557 24501 1613 24553
rect 1665 24501 1721 24553
rect 1773 24501 1829 24553
rect 1881 24501 1937 24553
rect 1989 24501 2045 24553
rect 2097 24501 2153 24553
rect 2205 24501 2261 24553
rect 2313 24501 2369 24553
rect 2421 24501 2477 24553
rect 2529 24501 2585 24553
rect 2637 24501 2693 24553
rect 2745 24501 2801 24553
rect 2853 24501 2909 24553
rect 2961 24501 3017 24553
rect 3069 24501 3125 24553
rect 3177 24501 3233 24553
rect 3285 24501 3309 24553
rect 1481 24445 3309 24501
rect 1481 24393 1505 24445
rect 1557 24393 1613 24445
rect 1665 24393 1721 24445
rect 1773 24393 1829 24445
rect 1881 24393 1937 24445
rect 1989 24393 2045 24445
rect 2097 24393 2153 24445
rect 2205 24393 2261 24445
rect 2313 24393 2369 24445
rect 2421 24393 2477 24445
rect 2529 24393 2585 24445
rect 2637 24393 2693 24445
rect 2745 24393 2801 24445
rect 2853 24393 2909 24445
rect 2961 24393 3017 24445
rect 3069 24393 3125 24445
rect 3177 24393 3233 24445
rect 3285 24393 3309 24445
rect 1481 23707 3309 24393
rect 1481 23655 1505 23707
rect 1557 23655 1613 23707
rect 1665 23655 1721 23707
rect 1773 23655 1829 23707
rect 1881 23655 1937 23707
rect 1989 23655 2045 23707
rect 2097 23655 2153 23707
rect 2205 23655 2261 23707
rect 2313 23655 2369 23707
rect 2421 23655 2477 23707
rect 2529 23655 2585 23707
rect 2637 23655 2693 23707
rect 2745 23655 2801 23707
rect 2853 23655 2909 23707
rect 2961 23655 3017 23707
rect 3069 23655 3125 23707
rect 3177 23655 3233 23707
rect 3285 23655 3309 23707
rect 1481 23219 3309 23655
rect 1481 23167 1505 23219
rect 1557 23167 1613 23219
rect 1665 23167 1721 23219
rect 1773 23167 1829 23219
rect 1881 23167 1937 23219
rect 1989 23167 2045 23219
rect 2097 23167 2153 23219
rect 2205 23167 2261 23219
rect 2313 23167 2369 23219
rect 2421 23167 2477 23219
rect 2529 23167 2585 23219
rect 2637 23167 2693 23219
rect 2745 23167 2801 23219
rect 2853 23167 2909 23219
rect 2961 23167 3017 23219
rect 3069 23167 3125 23219
rect 3177 23167 3233 23219
rect 3285 23167 3309 23219
rect 1481 22731 3309 23167
rect 1481 22679 1505 22731
rect 1557 22679 1613 22731
rect 1665 22679 1721 22731
rect 1773 22679 1829 22731
rect 1881 22679 1937 22731
rect 1989 22679 2045 22731
rect 2097 22679 2153 22731
rect 2205 22679 2261 22731
rect 2313 22679 2369 22731
rect 2421 22679 2477 22731
rect 2529 22679 2585 22731
rect 2637 22679 2693 22731
rect 2745 22679 2801 22731
rect 2853 22679 2909 22731
rect 2961 22679 3017 22731
rect 3069 22679 3125 22731
rect 3177 22679 3233 22731
rect 3285 22679 3309 22731
rect 1481 22243 3309 22679
rect 1481 22191 1505 22243
rect 1557 22191 1613 22243
rect 1665 22191 1721 22243
rect 1773 22191 1829 22243
rect 1881 22191 1937 22243
rect 1989 22191 2045 22243
rect 2097 22191 2153 22243
rect 2205 22191 2261 22243
rect 2313 22191 2369 22243
rect 2421 22191 2477 22243
rect 2529 22191 2585 22243
rect 2637 22191 2693 22243
rect 2745 22191 2801 22243
rect 2853 22191 2909 22243
rect 2961 22191 3017 22243
rect 3069 22191 3125 22243
rect 3177 22191 3233 22243
rect 3285 22191 3309 22243
rect 1481 21755 3309 22191
rect 1481 21703 1505 21755
rect 1557 21703 1613 21755
rect 1665 21703 1721 21755
rect 1773 21703 1829 21755
rect 1881 21703 1937 21755
rect 1989 21703 2045 21755
rect 2097 21703 2153 21755
rect 2205 21703 2261 21755
rect 2313 21703 2369 21755
rect 2421 21703 2477 21755
rect 2529 21703 2585 21755
rect 2637 21703 2693 21755
rect 2745 21703 2801 21755
rect 2853 21703 2909 21755
rect 2961 21703 3017 21755
rect 3069 21703 3125 21755
rect 3177 21703 3233 21755
rect 3285 21703 3309 21755
rect 1481 21267 3309 21703
rect 1481 21215 1505 21267
rect 1557 21215 1613 21267
rect 1665 21215 1721 21267
rect 1773 21215 1829 21267
rect 1881 21215 1937 21267
rect 1989 21215 2045 21267
rect 2097 21215 2153 21267
rect 2205 21215 2261 21267
rect 2313 21215 2369 21267
rect 2421 21215 2477 21267
rect 2529 21215 2585 21267
rect 2637 21215 2693 21267
rect 2745 21215 2801 21267
rect 2853 21215 2909 21267
rect 2961 21215 3017 21267
rect 3069 21215 3125 21267
rect 3177 21215 3233 21267
rect 3285 21215 3309 21267
rect 1481 20779 3309 21215
rect 1481 20727 1505 20779
rect 1557 20727 1613 20779
rect 1665 20727 1721 20779
rect 1773 20727 1829 20779
rect 1881 20727 1937 20779
rect 1989 20727 2045 20779
rect 2097 20727 2153 20779
rect 2205 20727 2261 20779
rect 2313 20727 2369 20779
rect 2421 20727 2477 20779
rect 2529 20727 2585 20779
rect 2637 20727 2693 20779
rect 2745 20727 2801 20779
rect 2853 20727 2909 20779
rect 2961 20727 3017 20779
rect 3069 20727 3125 20779
rect 3177 20727 3233 20779
rect 3285 20727 3309 20779
rect 1481 20291 3309 20727
rect 1481 20239 1505 20291
rect 1557 20239 1613 20291
rect 1665 20239 1721 20291
rect 1773 20239 1829 20291
rect 1881 20239 1937 20291
rect 1989 20239 2045 20291
rect 2097 20239 2153 20291
rect 2205 20239 2261 20291
rect 2313 20239 2369 20291
rect 2421 20239 2477 20291
rect 2529 20239 2585 20291
rect 2637 20239 2693 20291
rect 2745 20239 2801 20291
rect 2853 20239 2909 20291
rect 2961 20239 3017 20291
rect 3069 20239 3125 20291
rect 3177 20239 3233 20291
rect 3285 20239 3309 20291
rect 1481 19803 3309 20239
rect 1481 19751 1505 19803
rect 1557 19751 1613 19803
rect 1665 19751 1721 19803
rect 1773 19751 1829 19803
rect 1881 19751 1937 19803
rect 1989 19751 2045 19803
rect 2097 19751 2153 19803
rect 2205 19751 2261 19803
rect 2313 19751 2369 19803
rect 2421 19751 2477 19803
rect 2529 19751 2585 19803
rect 2637 19751 2693 19803
rect 2745 19751 2801 19803
rect 2853 19751 2909 19803
rect 2961 19751 3017 19803
rect 3069 19751 3125 19803
rect 3177 19751 3233 19803
rect 3285 19751 3309 19803
rect 1481 19315 3309 19751
rect 1481 19263 1505 19315
rect 1557 19263 1613 19315
rect 1665 19263 1721 19315
rect 1773 19263 1829 19315
rect 1881 19263 1937 19315
rect 1989 19263 2045 19315
rect 2097 19263 2153 19315
rect 2205 19263 2261 19315
rect 2313 19263 2369 19315
rect 2421 19263 2477 19315
rect 2529 19263 2585 19315
rect 2637 19263 2693 19315
rect 2745 19263 2801 19315
rect 2853 19263 2909 19315
rect 2961 19263 3017 19315
rect 3069 19263 3125 19315
rect 3177 19263 3233 19315
rect 3285 19263 3309 19315
rect 1481 18629 3309 19263
rect 1481 18577 1505 18629
rect 1557 18577 1613 18629
rect 1665 18577 1721 18629
rect 1773 18577 1829 18629
rect 1881 18577 1937 18629
rect 1989 18577 2045 18629
rect 2097 18577 2153 18629
rect 2205 18577 2261 18629
rect 2313 18577 2369 18629
rect 2421 18577 2477 18629
rect 2529 18577 2585 18629
rect 2637 18577 2693 18629
rect 2745 18577 2801 18629
rect 2853 18577 2909 18629
rect 2961 18577 3017 18629
rect 3069 18577 3125 18629
rect 3177 18577 3233 18629
rect 3285 18577 3309 18629
rect 1481 18521 3309 18577
rect 1481 18469 1505 18521
rect 1557 18469 1613 18521
rect 1665 18469 1721 18521
rect 1773 18469 1829 18521
rect 1881 18469 1937 18521
rect 1989 18469 2045 18521
rect 2097 18469 2153 18521
rect 2205 18469 2261 18521
rect 2313 18469 2369 18521
rect 2421 18469 2477 18521
rect 2529 18469 2585 18521
rect 2637 18469 2693 18521
rect 2745 18469 2801 18521
rect 2853 18469 2909 18521
rect 2961 18469 3017 18521
rect 3069 18469 3125 18521
rect 3177 18469 3233 18521
rect 3285 18469 3309 18521
rect 1481 17835 3309 18469
rect 1481 17783 1505 17835
rect 1557 17783 1613 17835
rect 1665 17783 1721 17835
rect 1773 17783 1829 17835
rect 1881 17783 1937 17835
rect 1989 17783 2045 17835
rect 2097 17783 2153 17835
rect 2205 17783 2261 17835
rect 2313 17783 2369 17835
rect 2421 17783 2477 17835
rect 2529 17783 2585 17835
rect 2637 17783 2693 17835
rect 2745 17783 2801 17835
rect 2853 17783 2909 17835
rect 2961 17783 3017 17835
rect 3069 17783 3125 17835
rect 3177 17783 3233 17835
rect 3285 17783 3309 17835
rect 1481 17347 3309 17783
rect 1481 17295 1505 17347
rect 1557 17295 1613 17347
rect 1665 17295 1721 17347
rect 1773 17295 1829 17347
rect 1881 17295 1937 17347
rect 1989 17295 2045 17347
rect 2097 17295 2153 17347
rect 2205 17295 2261 17347
rect 2313 17295 2369 17347
rect 2421 17295 2477 17347
rect 2529 17295 2585 17347
rect 2637 17295 2693 17347
rect 2745 17295 2801 17347
rect 2853 17295 2909 17347
rect 2961 17295 3017 17347
rect 3069 17295 3125 17347
rect 3177 17295 3233 17347
rect 3285 17295 3309 17347
rect 1481 16859 3309 17295
rect 1481 16807 1505 16859
rect 1557 16807 1613 16859
rect 1665 16807 1721 16859
rect 1773 16807 1829 16859
rect 1881 16807 1937 16859
rect 1989 16807 2045 16859
rect 2097 16807 2153 16859
rect 2205 16807 2261 16859
rect 2313 16807 2369 16859
rect 2421 16807 2477 16859
rect 2529 16807 2585 16859
rect 2637 16807 2693 16859
rect 2745 16807 2801 16859
rect 2853 16807 2909 16859
rect 2961 16807 3017 16859
rect 3069 16807 3125 16859
rect 3177 16807 3233 16859
rect 3285 16807 3309 16859
rect 1481 16371 3309 16807
rect 1481 16319 1505 16371
rect 1557 16319 1613 16371
rect 1665 16319 1721 16371
rect 1773 16319 1829 16371
rect 1881 16319 1937 16371
rect 1989 16319 2045 16371
rect 2097 16319 2153 16371
rect 2205 16319 2261 16371
rect 2313 16319 2369 16371
rect 2421 16319 2477 16371
rect 2529 16319 2585 16371
rect 2637 16319 2693 16371
rect 2745 16319 2801 16371
rect 2853 16319 2909 16371
rect 2961 16319 3017 16371
rect 3069 16319 3125 16371
rect 3177 16319 3233 16371
rect 3285 16319 3309 16371
rect 1481 15883 3309 16319
rect 1481 15831 1505 15883
rect 1557 15831 1613 15883
rect 1665 15831 1721 15883
rect 1773 15831 1829 15883
rect 1881 15831 1937 15883
rect 1989 15831 2045 15883
rect 2097 15831 2153 15883
rect 2205 15831 2261 15883
rect 2313 15831 2369 15883
rect 2421 15831 2477 15883
rect 2529 15831 2585 15883
rect 2637 15831 2693 15883
rect 2745 15831 2801 15883
rect 2853 15831 2909 15883
rect 2961 15831 3017 15883
rect 3069 15831 3125 15883
rect 3177 15831 3233 15883
rect 3285 15831 3309 15883
rect 1481 15395 3309 15831
rect 1481 15343 1505 15395
rect 1557 15343 1613 15395
rect 1665 15343 1721 15395
rect 1773 15343 1829 15395
rect 1881 15343 1937 15395
rect 1989 15343 2045 15395
rect 2097 15343 2153 15395
rect 2205 15343 2261 15395
rect 2313 15343 2369 15395
rect 2421 15343 2477 15395
rect 2529 15343 2585 15395
rect 2637 15343 2693 15395
rect 2745 15343 2801 15395
rect 2853 15343 2909 15395
rect 2961 15343 3017 15395
rect 3069 15343 3125 15395
rect 3177 15343 3233 15395
rect 3285 15343 3309 15395
rect 1481 14907 3309 15343
rect 1481 14855 1505 14907
rect 1557 14855 1613 14907
rect 1665 14855 1721 14907
rect 1773 14855 1829 14907
rect 1881 14855 1937 14907
rect 1989 14855 2045 14907
rect 2097 14855 2153 14907
rect 2205 14855 2261 14907
rect 2313 14855 2369 14907
rect 2421 14855 2477 14907
rect 2529 14855 2585 14907
rect 2637 14855 2693 14907
rect 2745 14855 2801 14907
rect 2853 14855 2909 14907
rect 2961 14855 3017 14907
rect 3069 14855 3125 14907
rect 3177 14855 3233 14907
rect 3285 14855 3309 14907
rect 1481 14419 3309 14855
rect 1481 14367 1505 14419
rect 1557 14367 1613 14419
rect 1665 14367 1721 14419
rect 1773 14367 1829 14419
rect 1881 14367 1937 14419
rect 1989 14367 2045 14419
rect 2097 14367 2153 14419
rect 2205 14367 2261 14419
rect 2313 14367 2369 14419
rect 2421 14367 2477 14419
rect 2529 14367 2585 14419
rect 2637 14367 2693 14419
rect 2745 14367 2801 14419
rect 2853 14367 2909 14419
rect 2961 14367 3017 14419
rect 3069 14367 3125 14419
rect 3177 14367 3233 14419
rect 3285 14367 3309 14419
rect 1481 13931 3309 14367
rect 1481 13879 1505 13931
rect 1557 13879 1613 13931
rect 1665 13879 1721 13931
rect 1773 13879 1829 13931
rect 1881 13879 1937 13931
rect 1989 13879 2045 13931
rect 2097 13879 2153 13931
rect 2205 13879 2261 13931
rect 2313 13879 2369 13931
rect 2421 13879 2477 13931
rect 2529 13879 2585 13931
rect 2637 13879 2693 13931
rect 2745 13879 2801 13931
rect 2853 13879 2909 13931
rect 2961 13879 3017 13931
rect 3069 13879 3125 13931
rect 3177 13879 3233 13931
rect 3285 13879 3309 13931
rect 1481 13443 3309 13879
rect 1481 13391 1505 13443
rect 1557 13391 1613 13443
rect 1665 13391 1721 13443
rect 1773 13391 1829 13443
rect 1881 13391 1937 13443
rect 1989 13391 2045 13443
rect 2097 13391 2153 13443
rect 2205 13391 2261 13443
rect 2313 13391 2369 13443
rect 2421 13391 2477 13443
rect 2529 13391 2585 13443
rect 2637 13391 2693 13443
rect 2745 13391 2801 13443
rect 2853 13391 2909 13443
rect 2961 13391 3017 13443
rect 3069 13391 3125 13443
rect 3177 13391 3233 13443
rect 3285 13391 3309 13443
rect 1481 12757 3309 13391
rect 1481 12705 1505 12757
rect 1557 12705 1613 12757
rect 1665 12705 1721 12757
rect 1773 12705 1829 12757
rect 1881 12705 1937 12757
rect 1989 12705 2045 12757
rect 2097 12705 2153 12757
rect 2205 12705 2261 12757
rect 2313 12705 2369 12757
rect 2421 12705 2477 12757
rect 2529 12705 2585 12757
rect 2637 12705 2693 12757
rect 2745 12705 2801 12757
rect 2853 12705 2909 12757
rect 2961 12705 3017 12757
rect 3069 12705 3125 12757
rect 3177 12705 3233 12757
rect 3285 12705 3309 12757
rect 1481 12649 3309 12705
rect 1481 12597 1505 12649
rect 1557 12597 1613 12649
rect 1665 12597 1721 12649
rect 1773 12597 1829 12649
rect 1881 12597 1937 12649
rect 1989 12597 2045 12649
rect 2097 12597 2153 12649
rect 2205 12597 2261 12649
rect 2313 12597 2369 12649
rect 2421 12597 2477 12649
rect 2529 12597 2585 12649
rect 2637 12597 2693 12649
rect 2745 12597 2801 12649
rect 2853 12597 2909 12649
rect 2961 12597 3017 12649
rect 3069 12597 3125 12649
rect 3177 12597 3233 12649
rect 3285 12597 3309 12649
rect 1481 11963 3309 12597
rect 1481 11911 1505 11963
rect 1557 11911 1613 11963
rect 1665 11911 1721 11963
rect 1773 11911 1829 11963
rect 1881 11911 1937 11963
rect 1989 11911 2045 11963
rect 2097 11911 2153 11963
rect 2205 11911 2261 11963
rect 2313 11911 2369 11963
rect 2421 11911 2477 11963
rect 2529 11911 2585 11963
rect 2637 11911 2693 11963
rect 2745 11911 2801 11963
rect 2853 11911 2909 11963
rect 2961 11911 3017 11963
rect 3069 11911 3125 11963
rect 3177 11911 3233 11963
rect 3285 11911 3309 11963
rect 1481 11475 3309 11911
rect 1481 11423 1505 11475
rect 1557 11423 1613 11475
rect 1665 11423 1721 11475
rect 1773 11423 1829 11475
rect 1881 11423 1937 11475
rect 1989 11423 2045 11475
rect 2097 11423 2153 11475
rect 2205 11423 2261 11475
rect 2313 11423 2369 11475
rect 2421 11423 2477 11475
rect 2529 11423 2585 11475
rect 2637 11423 2693 11475
rect 2745 11423 2801 11475
rect 2853 11423 2909 11475
rect 2961 11423 3017 11475
rect 3069 11423 3125 11475
rect 3177 11423 3233 11475
rect 3285 11423 3309 11475
rect 1481 10987 3309 11423
rect 1481 10935 1505 10987
rect 1557 10935 1613 10987
rect 1665 10935 1721 10987
rect 1773 10935 1829 10987
rect 1881 10935 1937 10987
rect 1989 10935 2045 10987
rect 2097 10935 2153 10987
rect 2205 10935 2261 10987
rect 2313 10935 2369 10987
rect 2421 10935 2477 10987
rect 2529 10935 2585 10987
rect 2637 10935 2693 10987
rect 2745 10935 2801 10987
rect 2853 10935 2909 10987
rect 2961 10935 3017 10987
rect 3069 10935 3125 10987
rect 3177 10935 3233 10987
rect 3285 10935 3309 10987
rect 1481 10499 3309 10935
rect 1481 10447 1505 10499
rect 1557 10447 1613 10499
rect 1665 10447 1721 10499
rect 1773 10447 1829 10499
rect 1881 10447 1937 10499
rect 1989 10447 2045 10499
rect 2097 10447 2153 10499
rect 2205 10447 2261 10499
rect 2313 10447 2369 10499
rect 2421 10447 2477 10499
rect 2529 10447 2585 10499
rect 2637 10447 2693 10499
rect 2745 10447 2801 10499
rect 2853 10447 2909 10499
rect 2961 10447 3017 10499
rect 3069 10447 3125 10499
rect 3177 10447 3233 10499
rect 3285 10447 3309 10499
rect 1481 10011 3309 10447
rect 1481 9959 1505 10011
rect 1557 9959 1613 10011
rect 1665 9959 1721 10011
rect 1773 9959 1829 10011
rect 1881 9959 1937 10011
rect 1989 9959 2045 10011
rect 2097 9959 2153 10011
rect 2205 9959 2261 10011
rect 2313 9959 2369 10011
rect 2421 9959 2477 10011
rect 2529 9959 2585 10011
rect 2637 9959 2693 10011
rect 2745 9959 2801 10011
rect 2853 9959 2909 10011
rect 2961 9959 3017 10011
rect 3069 9959 3125 10011
rect 3177 9959 3233 10011
rect 3285 9959 3309 10011
rect 1481 9523 3309 9959
rect 1481 9471 1505 9523
rect 1557 9471 1613 9523
rect 1665 9471 1721 9523
rect 1773 9471 1829 9523
rect 1881 9471 1937 9523
rect 1989 9471 2045 9523
rect 2097 9471 2153 9523
rect 2205 9471 2261 9523
rect 2313 9471 2369 9523
rect 2421 9471 2477 9523
rect 2529 9471 2585 9523
rect 2637 9471 2693 9523
rect 2745 9471 2801 9523
rect 2853 9471 2909 9523
rect 2961 9471 3017 9523
rect 3069 9471 3125 9523
rect 3177 9471 3233 9523
rect 3285 9471 3309 9523
rect 1481 9035 3309 9471
rect 1481 8983 1505 9035
rect 1557 8983 1613 9035
rect 1665 8983 1721 9035
rect 1773 8983 1829 9035
rect 1881 8983 1937 9035
rect 1989 8983 2045 9035
rect 2097 8983 2153 9035
rect 2205 8983 2261 9035
rect 2313 8983 2369 9035
rect 2421 8983 2477 9035
rect 2529 8983 2585 9035
rect 2637 8983 2693 9035
rect 2745 8983 2801 9035
rect 2853 8983 2909 9035
rect 2961 8983 3017 9035
rect 3069 8983 3125 9035
rect 3177 8983 3233 9035
rect 3285 8983 3309 9035
rect 1481 8547 3309 8983
rect 1481 8495 1505 8547
rect 1557 8495 1613 8547
rect 1665 8495 1721 8547
rect 1773 8495 1829 8547
rect 1881 8495 1937 8547
rect 1989 8495 2045 8547
rect 2097 8495 2153 8547
rect 2205 8495 2261 8547
rect 2313 8495 2369 8547
rect 2421 8495 2477 8547
rect 2529 8495 2585 8547
rect 2637 8495 2693 8547
rect 2745 8495 2801 8547
rect 2853 8495 2909 8547
rect 2961 8495 3017 8547
rect 3069 8495 3125 8547
rect 3177 8495 3233 8547
rect 3285 8495 3309 8547
rect 1481 8059 3309 8495
rect 1481 8007 1505 8059
rect 1557 8007 1613 8059
rect 1665 8007 1721 8059
rect 1773 8007 1829 8059
rect 1881 8007 1937 8059
rect 1989 8007 2045 8059
rect 2097 8007 2153 8059
rect 2205 8007 2261 8059
rect 2313 8007 2369 8059
rect 2421 8007 2477 8059
rect 2529 8007 2585 8059
rect 2637 8007 2693 8059
rect 2745 8007 2801 8059
rect 2853 8007 2909 8059
rect 2961 8007 3017 8059
rect 3069 8007 3125 8059
rect 3177 8007 3233 8059
rect 3285 8007 3309 8059
rect 1481 7571 3309 8007
rect 1481 7519 1505 7571
rect 1557 7519 1613 7571
rect 1665 7519 1721 7571
rect 1773 7519 1829 7571
rect 1881 7519 1937 7571
rect 1989 7519 2045 7571
rect 2097 7519 2153 7571
rect 2205 7519 2261 7571
rect 2313 7519 2369 7571
rect 2421 7519 2477 7571
rect 2529 7519 2585 7571
rect 2637 7519 2693 7571
rect 2745 7519 2801 7571
rect 2853 7519 2909 7571
rect 2961 7519 3017 7571
rect 3069 7519 3125 7571
rect 3177 7519 3233 7571
rect 3285 7519 3309 7571
rect 1481 6885 3309 7519
rect 1481 6833 1505 6885
rect 1557 6833 1613 6885
rect 1665 6833 1721 6885
rect 1773 6833 1829 6885
rect 1881 6833 1937 6885
rect 1989 6833 2045 6885
rect 2097 6833 2153 6885
rect 2205 6833 2261 6885
rect 2313 6833 2369 6885
rect 2421 6833 2477 6885
rect 2529 6833 2585 6885
rect 2637 6833 2693 6885
rect 2745 6833 2801 6885
rect 2853 6833 2909 6885
rect 2961 6833 3017 6885
rect 3069 6833 3125 6885
rect 3177 6833 3233 6885
rect 3285 6833 3309 6885
rect 1481 6777 3309 6833
rect 1481 6725 1505 6777
rect 1557 6725 1613 6777
rect 1665 6725 1721 6777
rect 1773 6725 1829 6777
rect 1881 6725 1937 6777
rect 1989 6725 2045 6777
rect 2097 6725 2153 6777
rect 2205 6725 2261 6777
rect 2313 6725 2369 6777
rect 2421 6725 2477 6777
rect 2529 6725 2585 6777
rect 2637 6725 2693 6777
rect 2745 6725 2801 6777
rect 2853 6725 2909 6777
rect 2961 6725 3017 6777
rect 3069 6725 3125 6777
rect 3177 6725 3233 6777
rect 3285 6725 3309 6777
rect 1481 6091 3309 6725
rect 1481 6039 1505 6091
rect 1557 6039 1613 6091
rect 1665 6039 1721 6091
rect 1773 6039 1829 6091
rect 1881 6039 1937 6091
rect 1989 6039 2045 6091
rect 2097 6039 2153 6091
rect 2205 6039 2261 6091
rect 2313 6039 2369 6091
rect 2421 6039 2477 6091
rect 2529 6039 2585 6091
rect 2637 6039 2693 6091
rect 2745 6039 2801 6091
rect 2853 6039 2909 6091
rect 2961 6039 3017 6091
rect 3069 6039 3125 6091
rect 3177 6039 3233 6091
rect 3285 6039 3309 6091
rect 1481 5603 3309 6039
rect 1481 5551 1505 5603
rect 1557 5551 1613 5603
rect 1665 5551 1721 5603
rect 1773 5551 1829 5603
rect 1881 5551 1937 5603
rect 1989 5551 2045 5603
rect 2097 5551 2153 5603
rect 2205 5551 2261 5603
rect 2313 5551 2369 5603
rect 2421 5551 2477 5603
rect 2529 5551 2585 5603
rect 2637 5551 2693 5603
rect 2745 5551 2801 5603
rect 2853 5551 2909 5603
rect 2961 5551 3017 5603
rect 3069 5551 3125 5603
rect 3177 5551 3233 5603
rect 3285 5551 3309 5603
rect 1481 5115 3309 5551
rect 1481 5063 1505 5115
rect 1557 5063 1613 5115
rect 1665 5063 1721 5115
rect 1773 5063 1829 5115
rect 1881 5063 1937 5115
rect 1989 5063 2045 5115
rect 2097 5063 2153 5115
rect 2205 5063 2261 5115
rect 2313 5063 2369 5115
rect 2421 5063 2477 5115
rect 2529 5063 2585 5115
rect 2637 5063 2693 5115
rect 2745 5063 2801 5115
rect 2853 5063 2909 5115
rect 2961 5063 3017 5115
rect 3069 5063 3125 5115
rect 3177 5063 3233 5115
rect 3285 5063 3309 5115
rect 1481 4627 3309 5063
rect 1481 4575 1505 4627
rect 1557 4575 1613 4627
rect 1665 4575 1721 4627
rect 1773 4575 1829 4627
rect 1881 4575 1937 4627
rect 1989 4575 2045 4627
rect 2097 4575 2153 4627
rect 2205 4575 2261 4627
rect 2313 4575 2369 4627
rect 2421 4575 2477 4627
rect 2529 4575 2585 4627
rect 2637 4575 2693 4627
rect 2745 4575 2801 4627
rect 2853 4575 2909 4627
rect 2961 4575 3017 4627
rect 3069 4575 3125 4627
rect 3177 4575 3233 4627
rect 3285 4575 3309 4627
rect 1481 4139 3309 4575
rect 1481 4087 1505 4139
rect 1557 4087 1613 4139
rect 1665 4087 1721 4139
rect 1773 4087 1829 4139
rect 1881 4087 1937 4139
rect 1989 4087 2045 4139
rect 2097 4087 2153 4139
rect 2205 4087 2261 4139
rect 2313 4087 2369 4139
rect 2421 4087 2477 4139
rect 2529 4087 2585 4139
rect 2637 4087 2693 4139
rect 2745 4087 2801 4139
rect 2853 4087 2909 4139
rect 2961 4087 3017 4139
rect 3069 4087 3125 4139
rect 3177 4087 3233 4139
rect 3285 4087 3309 4139
rect 1481 3651 3309 4087
rect 1481 3599 1505 3651
rect 1557 3599 1613 3651
rect 1665 3599 1721 3651
rect 1773 3599 1829 3651
rect 1881 3599 1937 3651
rect 1989 3599 2045 3651
rect 2097 3599 2153 3651
rect 2205 3599 2261 3651
rect 2313 3599 2369 3651
rect 2421 3599 2477 3651
rect 2529 3599 2585 3651
rect 2637 3599 2693 3651
rect 2745 3599 2801 3651
rect 2853 3599 2909 3651
rect 2961 3599 3017 3651
rect 3069 3599 3125 3651
rect 3177 3599 3233 3651
rect 3285 3599 3309 3651
rect 1481 3163 3309 3599
rect 1481 3111 1505 3163
rect 1557 3111 1613 3163
rect 1665 3111 1721 3163
rect 1773 3111 1829 3163
rect 1881 3111 1937 3163
rect 1989 3111 2045 3163
rect 2097 3111 2153 3163
rect 2205 3111 2261 3163
rect 2313 3111 2369 3163
rect 2421 3111 2477 3163
rect 2529 3111 2585 3163
rect 2637 3111 2693 3163
rect 2745 3111 2801 3163
rect 2853 3111 2909 3163
rect 2961 3111 3017 3163
rect 3069 3111 3125 3163
rect 3177 3111 3233 3163
rect 3285 3111 3309 3163
rect 1481 2675 3309 3111
rect 1481 2623 1505 2675
rect 1557 2623 1613 2675
rect 1665 2623 1721 2675
rect 1773 2623 1829 2675
rect 1881 2623 1937 2675
rect 1989 2623 2045 2675
rect 2097 2623 2153 2675
rect 2205 2623 2261 2675
rect 2313 2623 2369 2675
rect 2421 2623 2477 2675
rect 2529 2623 2585 2675
rect 2637 2623 2693 2675
rect 2745 2623 2801 2675
rect 2853 2623 2909 2675
rect 2961 2623 3017 2675
rect 3069 2623 3125 2675
rect 3177 2623 3233 2675
rect 3285 2623 3309 2675
rect 1481 2187 3309 2623
rect 1481 2135 1505 2187
rect 1557 2135 1613 2187
rect 1665 2135 1721 2187
rect 1773 2135 1829 2187
rect 1881 2135 1937 2187
rect 1989 2135 2045 2187
rect 2097 2135 2153 2187
rect 2205 2135 2261 2187
rect 2313 2135 2369 2187
rect 2421 2135 2477 2187
rect 2529 2135 2585 2187
rect 2637 2135 2693 2187
rect 2745 2135 2801 2187
rect 2853 2135 2909 2187
rect 2961 2135 3017 2187
rect 3069 2135 3125 2187
rect 3177 2135 3233 2187
rect 3285 2135 3309 2187
rect 1481 1699 3309 2135
rect 1481 1647 1505 1699
rect 1557 1647 1613 1699
rect 1665 1647 1721 1699
rect 1773 1647 1829 1699
rect 1881 1647 1937 1699
rect 1989 1647 2045 1699
rect 2097 1647 2153 1699
rect 2205 1647 2261 1699
rect 2313 1647 2369 1699
rect 2421 1647 2477 1699
rect 2529 1647 2585 1699
rect 2637 1647 2693 1699
rect 2745 1647 2801 1699
rect 2853 1647 2909 1699
rect 2961 1647 3017 1699
rect 3069 1647 3125 1699
rect 3177 1647 3233 1699
rect 3285 1647 3309 1699
rect 43 1365 93 1417
rect 145 1365 201 1417
rect 253 1365 309 1417
rect 361 1365 1145 1417
rect 43 1309 1145 1365
rect 43 1257 93 1309
rect 145 1257 201 1309
rect 253 1257 309 1309
rect 361 1257 1145 1309
rect 43 1201 1145 1257
rect 43 1149 93 1201
rect 145 1149 201 1201
rect 253 1149 309 1201
rect 361 1149 1145 1201
rect 43 1093 1145 1149
rect 43 1041 93 1093
rect 145 1041 201 1093
rect 253 1041 309 1093
rect 361 1041 1145 1093
rect 43 985 1145 1041
rect 43 933 93 985
rect 145 933 201 985
rect 253 933 309 985
rect 361 933 1145 985
rect 43 877 1145 933
rect 43 825 93 877
rect 145 825 201 877
rect 253 825 309 877
rect 361 825 1145 877
rect 43 769 1145 825
rect 43 717 93 769
rect 145 717 201 769
rect 253 717 309 769
rect 361 717 1145 769
rect 43 661 1145 717
rect 43 609 93 661
rect 145 609 201 661
rect 253 609 309 661
rect 361 609 1145 661
rect 43 553 1145 609
rect 43 501 93 553
rect 145 501 201 553
rect 253 501 309 553
rect 361 501 1145 553
rect 43 361 1145 501
rect 43 309 82 361
rect 134 309 190 361
rect 242 309 298 361
rect 350 309 406 361
rect 458 309 514 361
rect 566 309 622 361
rect 674 309 730 361
rect 782 309 838 361
rect 890 309 946 361
rect 998 309 1054 361
rect 1106 309 1145 361
rect 43 253 1145 309
rect 43 201 82 253
rect 134 201 190 253
rect 242 201 298 253
rect 350 201 406 253
rect 458 201 514 253
rect 566 201 622 253
rect 674 201 730 253
rect 782 201 838 253
rect 890 201 946 253
rect 998 201 1054 253
rect 1106 201 1145 253
rect 43 145 1145 201
rect 43 93 82 145
rect 134 93 190 145
rect 242 93 298 145
rect 350 93 406 145
rect 458 93 514 145
rect 566 93 622 145
rect 674 93 730 145
rect 782 93 838 145
rect 890 93 946 145
rect 998 93 1054 145
rect 1106 93 1145 145
rect 43 43 1145 93
rect 1481 961 3309 1647
rect 1481 909 1505 961
rect 1557 909 1613 961
rect 1665 909 1721 961
rect 1773 909 1829 961
rect 1881 909 1937 961
rect 1989 909 2045 961
rect 2097 909 2153 961
rect 2205 909 2261 961
rect 2313 909 2369 961
rect 2421 909 2477 961
rect 2529 909 2585 961
rect 2637 909 2693 961
rect 2745 909 2801 961
rect 2853 909 2909 961
rect 2961 909 3017 961
rect 3069 909 3125 961
rect 3177 909 3233 961
rect 3285 909 3309 961
rect 1481 853 3309 909
rect 1481 801 1505 853
rect 1557 801 1613 853
rect 1665 801 1721 853
rect 1773 801 1829 853
rect 1881 801 1937 853
rect 1989 801 2045 853
rect 2097 801 2153 853
rect 2205 801 2261 853
rect 2313 801 2369 853
rect 2421 801 2477 853
rect 2529 801 2585 853
rect 2637 801 2693 853
rect 2745 801 2801 853
rect 2853 801 2909 853
rect 2961 801 3017 853
rect 3069 801 3125 853
rect 3177 801 3233 853
rect 3285 801 3309 853
rect 1481 745 3309 801
rect 1481 693 1505 745
rect 1557 693 1613 745
rect 1665 693 1721 745
rect 1773 693 1829 745
rect 1881 693 1937 745
rect 1989 693 2045 745
rect 2097 693 2153 745
rect 2205 693 2261 745
rect 2313 693 2369 745
rect 2421 693 2477 745
rect 2529 693 2585 745
rect 2637 693 2693 745
rect 2745 693 2801 745
rect 2853 693 2909 745
rect 2961 693 3017 745
rect 3069 693 3125 745
rect 3177 693 3233 745
rect 3285 693 3309 745
rect 1481 43 3309 693
rect 3409 25261 5237 25617
rect 3409 25209 3433 25261
rect 3485 25209 3541 25261
rect 3593 25209 3649 25261
rect 3701 25209 3757 25261
rect 3809 25209 3865 25261
rect 3917 25209 3973 25261
rect 4025 25209 4081 25261
rect 4133 25209 4189 25261
rect 4241 25209 4297 25261
rect 4349 25209 4405 25261
rect 4457 25209 4513 25261
rect 4565 25209 4621 25261
rect 4673 25209 4729 25261
rect 4781 25209 4837 25261
rect 4889 25209 4945 25261
rect 4997 25209 5053 25261
rect 5105 25209 5161 25261
rect 5213 25209 5237 25261
rect 3409 25153 5237 25209
rect 3409 25101 3433 25153
rect 3485 25101 3541 25153
rect 3593 25101 3649 25153
rect 3701 25101 3757 25153
rect 3809 25101 3865 25153
rect 3917 25101 3973 25153
rect 4025 25101 4081 25153
rect 4133 25101 4189 25153
rect 4241 25101 4297 25153
rect 4349 25101 4405 25153
rect 4457 25101 4513 25153
rect 4565 25101 4621 25153
rect 4673 25101 4729 25153
rect 4781 25101 4837 25153
rect 4889 25101 4945 25153
rect 4997 25101 5053 25153
rect 5105 25101 5161 25153
rect 5213 25101 5237 25153
rect 3409 25045 5237 25101
rect 3409 24993 3433 25045
rect 3485 24993 3541 25045
rect 3593 24993 3649 25045
rect 3701 24993 3757 25045
rect 3809 24993 3865 25045
rect 3917 24993 3973 25045
rect 4025 24993 4081 25045
rect 4133 24993 4189 25045
rect 4241 24993 4297 25045
rect 4349 24993 4405 25045
rect 4457 24993 4513 25045
rect 4565 24993 4621 25045
rect 4673 24993 4729 25045
rect 4781 24993 4837 25045
rect 4889 24993 4945 25045
rect 4997 24993 5053 25045
rect 5105 24993 5161 25045
rect 5213 24993 5237 25045
rect 3409 23951 5237 24993
rect 3409 23899 3433 23951
rect 3485 23899 3541 23951
rect 3593 23899 3649 23951
rect 3701 23899 3757 23951
rect 3809 23899 3865 23951
rect 3917 23899 3973 23951
rect 4025 23899 4081 23951
rect 4133 23899 4189 23951
rect 4241 23899 4297 23951
rect 4349 23899 4405 23951
rect 4457 23899 4513 23951
rect 4565 23899 4621 23951
rect 4673 23899 4729 23951
rect 4781 23899 4837 23951
rect 4889 23899 4945 23951
rect 4997 23899 5053 23951
rect 5105 23899 5161 23951
rect 5213 23899 5237 23951
rect 3409 23463 5237 23899
rect 3409 23411 3433 23463
rect 3485 23411 3541 23463
rect 3593 23411 3649 23463
rect 3701 23411 3757 23463
rect 3809 23411 3865 23463
rect 3917 23411 3973 23463
rect 4025 23411 4081 23463
rect 4133 23411 4189 23463
rect 4241 23411 4297 23463
rect 4349 23411 4405 23463
rect 4457 23411 4513 23463
rect 4565 23411 4621 23463
rect 4673 23411 4729 23463
rect 4781 23411 4837 23463
rect 4889 23411 4945 23463
rect 4997 23411 5053 23463
rect 5105 23411 5161 23463
rect 5213 23411 5237 23463
rect 3409 22975 5237 23411
rect 3409 22923 3433 22975
rect 3485 22923 3541 22975
rect 3593 22923 3649 22975
rect 3701 22923 3757 22975
rect 3809 22923 3865 22975
rect 3917 22923 3973 22975
rect 4025 22923 4081 22975
rect 4133 22923 4189 22975
rect 4241 22923 4297 22975
rect 4349 22923 4405 22975
rect 4457 22923 4513 22975
rect 4565 22923 4621 22975
rect 4673 22923 4729 22975
rect 4781 22923 4837 22975
rect 4889 22923 4945 22975
rect 4997 22923 5053 22975
rect 5105 22923 5161 22975
rect 5213 22923 5237 22975
rect 3409 22487 5237 22923
rect 3409 22435 3433 22487
rect 3485 22435 3541 22487
rect 3593 22435 3649 22487
rect 3701 22435 3757 22487
rect 3809 22435 3865 22487
rect 3917 22435 3973 22487
rect 4025 22435 4081 22487
rect 4133 22435 4189 22487
rect 4241 22435 4297 22487
rect 4349 22435 4405 22487
rect 4457 22435 4513 22487
rect 4565 22435 4621 22487
rect 4673 22435 4729 22487
rect 4781 22435 4837 22487
rect 4889 22435 4945 22487
rect 4997 22435 5053 22487
rect 5105 22435 5161 22487
rect 5213 22435 5237 22487
rect 3409 21999 5237 22435
rect 3409 21947 3433 21999
rect 3485 21947 3541 21999
rect 3593 21947 3649 21999
rect 3701 21947 3757 21999
rect 3809 21947 3865 21999
rect 3917 21947 3973 21999
rect 4025 21947 4081 21999
rect 4133 21947 4189 21999
rect 4241 21947 4297 21999
rect 4349 21947 4405 21999
rect 4457 21947 4513 21999
rect 4565 21947 4621 21999
rect 4673 21947 4729 21999
rect 4781 21947 4837 21999
rect 4889 21947 4945 21999
rect 4997 21947 5053 21999
rect 5105 21947 5161 21999
rect 5213 21947 5237 21999
rect 3409 21511 5237 21947
rect 3409 21459 3433 21511
rect 3485 21459 3541 21511
rect 3593 21459 3649 21511
rect 3701 21459 3757 21511
rect 3809 21459 3865 21511
rect 3917 21459 3973 21511
rect 4025 21459 4081 21511
rect 4133 21459 4189 21511
rect 4241 21459 4297 21511
rect 4349 21459 4405 21511
rect 4457 21459 4513 21511
rect 4565 21459 4621 21511
rect 4673 21459 4729 21511
rect 4781 21459 4837 21511
rect 4889 21459 4945 21511
rect 4997 21459 5053 21511
rect 5105 21459 5161 21511
rect 5213 21459 5237 21511
rect 3409 21023 5237 21459
rect 3409 20971 3433 21023
rect 3485 20971 3541 21023
rect 3593 20971 3649 21023
rect 3701 20971 3757 21023
rect 3809 20971 3865 21023
rect 3917 20971 3973 21023
rect 4025 20971 4081 21023
rect 4133 20971 4189 21023
rect 4241 20971 4297 21023
rect 4349 20971 4405 21023
rect 4457 20971 4513 21023
rect 4565 20971 4621 21023
rect 4673 20971 4729 21023
rect 4781 20971 4837 21023
rect 4889 20971 4945 21023
rect 4997 20971 5053 21023
rect 5105 20971 5161 21023
rect 5213 20971 5237 21023
rect 3409 20535 5237 20971
rect 3409 20483 3433 20535
rect 3485 20483 3541 20535
rect 3593 20483 3649 20535
rect 3701 20483 3757 20535
rect 3809 20483 3865 20535
rect 3917 20483 3973 20535
rect 4025 20483 4081 20535
rect 4133 20483 4189 20535
rect 4241 20483 4297 20535
rect 4349 20483 4405 20535
rect 4457 20483 4513 20535
rect 4565 20483 4621 20535
rect 4673 20483 4729 20535
rect 4781 20483 4837 20535
rect 4889 20483 4945 20535
rect 4997 20483 5053 20535
rect 5105 20483 5161 20535
rect 5213 20483 5237 20535
rect 3409 20047 5237 20483
rect 3409 19995 3433 20047
rect 3485 19995 3541 20047
rect 3593 19995 3649 20047
rect 3701 19995 3757 20047
rect 3809 19995 3865 20047
rect 3917 19995 3973 20047
rect 4025 19995 4081 20047
rect 4133 19995 4189 20047
rect 4241 19995 4297 20047
rect 4349 19995 4405 20047
rect 4457 19995 4513 20047
rect 4565 19995 4621 20047
rect 4673 19995 4729 20047
rect 4781 19995 4837 20047
rect 4889 19995 4945 20047
rect 4997 19995 5053 20047
rect 5105 19995 5161 20047
rect 5213 19995 5237 20047
rect 3409 19559 5237 19995
rect 3409 19507 3433 19559
rect 3485 19507 3541 19559
rect 3593 19507 3649 19559
rect 3701 19507 3757 19559
rect 3809 19507 3865 19559
rect 3917 19507 3973 19559
rect 4025 19507 4081 19559
rect 4133 19507 4189 19559
rect 4241 19507 4297 19559
rect 4349 19507 4405 19559
rect 4457 19507 4513 19559
rect 4565 19507 4621 19559
rect 4673 19507 4729 19559
rect 4781 19507 4837 19559
rect 4889 19507 4945 19559
rect 4997 19507 5053 19559
rect 5105 19507 5161 19559
rect 5213 19507 5237 19559
rect 3409 19071 5237 19507
rect 3409 19019 3433 19071
rect 3485 19019 3541 19071
rect 3593 19019 3649 19071
rect 3701 19019 3757 19071
rect 3809 19019 3865 19071
rect 3917 19019 3973 19071
rect 4025 19019 4081 19071
rect 4133 19019 4189 19071
rect 4241 19019 4297 19071
rect 4349 19019 4405 19071
rect 4457 19019 4513 19071
rect 4565 19019 4621 19071
rect 4673 19019 4729 19071
rect 4781 19019 4837 19071
rect 4889 19019 4945 19071
rect 4997 19019 5053 19071
rect 5105 19019 5161 19071
rect 5213 19019 5237 19071
rect 3409 18079 5237 19019
rect 3409 18027 3433 18079
rect 3485 18027 3541 18079
rect 3593 18027 3649 18079
rect 3701 18027 3757 18079
rect 3809 18027 3865 18079
rect 3917 18027 3973 18079
rect 4025 18027 4081 18079
rect 4133 18027 4189 18079
rect 4241 18027 4297 18079
rect 4349 18027 4405 18079
rect 4457 18027 4513 18079
rect 4565 18027 4621 18079
rect 4673 18027 4729 18079
rect 4781 18027 4837 18079
rect 4889 18027 4945 18079
rect 4997 18027 5053 18079
rect 5105 18027 5161 18079
rect 5213 18027 5237 18079
rect 3409 17591 5237 18027
rect 3409 17539 3433 17591
rect 3485 17539 3541 17591
rect 3593 17539 3649 17591
rect 3701 17539 3757 17591
rect 3809 17539 3865 17591
rect 3917 17539 3973 17591
rect 4025 17539 4081 17591
rect 4133 17539 4189 17591
rect 4241 17539 4297 17591
rect 4349 17539 4405 17591
rect 4457 17539 4513 17591
rect 4565 17539 4621 17591
rect 4673 17539 4729 17591
rect 4781 17539 4837 17591
rect 4889 17539 4945 17591
rect 4997 17539 5053 17591
rect 5105 17539 5161 17591
rect 5213 17539 5237 17591
rect 3409 17103 5237 17539
rect 3409 17051 3433 17103
rect 3485 17051 3541 17103
rect 3593 17051 3649 17103
rect 3701 17051 3757 17103
rect 3809 17051 3865 17103
rect 3917 17051 3973 17103
rect 4025 17051 4081 17103
rect 4133 17051 4189 17103
rect 4241 17051 4297 17103
rect 4349 17051 4405 17103
rect 4457 17051 4513 17103
rect 4565 17051 4621 17103
rect 4673 17051 4729 17103
rect 4781 17051 4837 17103
rect 4889 17051 4945 17103
rect 4997 17051 5053 17103
rect 5105 17051 5161 17103
rect 5213 17051 5237 17103
rect 3409 16615 5237 17051
rect 3409 16563 3433 16615
rect 3485 16563 3541 16615
rect 3593 16563 3649 16615
rect 3701 16563 3757 16615
rect 3809 16563 3865 16615
rect 3917 16563 3973 16615
rect 4025 16563 4081 16615
rect 4133 16563 4189 16615
rect 4241 16563 4297 16615
rect 4349 16563 4405 16615
rect 4457 16563 4513 16615
rect 4565 16563 4621 16615
rect 4673 16563 4729 16615
rect 4781 16563 4837 16615
rect 4889 16563 4945 16615
rect 4997 16563 5053 16615
rect 5105 16563 5161 16615
rect 5213 16563 5237 16615
rect 3409 16127 5237 16563
rect 3409 16075 3433 16127
rect 3485 16075 3541 16127
rect 3593 16075 3649 16127
rect 3701 16075 3757 16127
rect 3809 16075 3865 16127
rect 3917 16075 3973 16127
rect 4025 16075 4081 16127
rect 4133 16075 4189 16127
rect 4241 16075 4297 16127
rect 4349 16075 4405 16127
rect 4457 16075 4513 16127
rect 4565 16075 4621 16127
rect 4673 16075 4729 16127
rect 4781 16075 4837 16127
rect 4889 16075 4945 16127
rect 4997 16075 5053 16127
rect 5105 16075 5161 16127
rect 5213 16075 5237 16127
rect 3409 15639 5237 16075
rect 3409 15587 3433 15639
rect 3485 15587 3541 15639
rect 3593 15587 3649 15639
rect 3701 15587 3757 15639
rect 3809 15587 3865 15639
rect 3917 15587 3973 15639
rect 4025 15587 4081 15639
rect 4133 15587 4189 15639
rect 4241 15587 4297 15639
rect 4349 15587 4405 15639
rect 4457 15587 4513 15639
rect 4565 15587 4621 15639
rect 4673 15587 4729 15639
rect 4781 15587 4837 15639
rect 4889 15587 4945 15639
rect 4997 15587 5053 15639
rect 5105 15587 5161 15639
rect 5213 15587 5237 15639
rect 3409 15151 5237 15587
rect 3409 15099 3433 15151
rect 3485 15099 3541 15151
rect 3593 15099 3649 15151
rect 3701 15099 3757 15151
rect 3809 15099 3865 15151
rect 3917 15099 3973 15151
rect 4025 15099 4081 15151
rect 4133 15099 4189 15151
rect 4241 15099 4297 15151
rect 4349 15099 4405 15151
rect 4457 15099 4513 15151
rect 4565 15099 4621 15151
rect 4673 15099 4729 15151
rect 4781 15099 4837 15151
rect 4889 15099 4945 15151
rect 4997 15099 5053 15151
rect 5105 15099 5161 15151
rect 5213 15099 5237 15151
rect 3409 14663 5237 15099
rect 3409 14611 3433 14663
rect 3485 14611 3541 14663
rect 3593 14611 3649 14663
rect 3701 14611 3757 14663
rect 3809 14611 3865 14663
rect 3917 14611 3973 14663
rect 4025 14611 4081 14663
rect 4133 14611 4189 14663
rect 4241 14611 4297 14663
rect 4349 14611 4405 14663
rect 4457 14611 4513 14663
rect 4565 14611 4621 14663
rect 4673 14611 4729 14663
rect 4781 14611 4837 14663
rect 4889 14611 4945 14663
rect 4997 14611 5053 14663
rect 5105 14611 5161 14663
rect 5213 14611 5237 14663
rect 3409 14175 5237 14611
rect 3409 14123 3433 14175
rect 3485 14123 3541 14175
rect 3593 14123 3649 14175
rect 3701 14123 3757 14175
rect 3809 14123 3865 14175
rect 3917 14123 3973 14175
rect 4025 14123 4081 14175
rect 4133 14123 4189 14175
rect 4241 14123 4297 14175
rect 4349 14123 4405 14175
rect 4457 14123 4513 14175
rect 4565 14123 4621 14175
rect 4673 14123 4729 14175
rect 4781 14123 4837 14175
rect 4889 14123 4945 14175
rect 4997 14123 5053 14175
rect 5105 14123 5161 14175
rect 5213 14123 5237 14175
rect 3409 13687 5237 14123
rect 3409 13635 3433 13687
rect 3485 13635 3541 13687
rect 3593 13635 3649 13687
rect 3701 13635 3757 13687
rect 3809 13635 3865 13687
rect 3917 13635 3973 13687
rect 4025 13635 4081 13687
rect 4133 13635 4189 13687
rect 4241 13635 4297 13687
rect 4349 13635 4405 13687
rect 4457 13635 4513 13687
rect 4565 13635 4621 13687
rect 4673 13635 4729 13687
rect 4781 13635 4837 13687
rect 4889 13635 4945 13687
rect 4997 13635 5053 13687
rect 5105 13635 5161 13687
rect 5213 13635 5237 13687
rect 3409 13199 5237 13635
rect 3409 13147 3433 13199
rect 3485 13147 3541 13199
rect 3593 13147 3649 13199
rect 3701 13147 3757 13199
rect 3809 13147 3865 13199
rect 3917 13147 3973 13199
rect 4025 13147 4081 13199
rect 4133 13147 4189 13199
rect 4241 13147 4297 13199
rect 4349 13147 4405 13199
rect 4457 13147 4513 13199
rect 4565 13147 4621 13199
rect 4673 13147 4729 13199
rect 4781 13147 4837 13199
rect 4889 13147 4945 13199
rect 4997 13147 5053 13199
rect 5105 13147 5161 13199
rect 5213 13147 5237 13199
rect 3409 12207 5237 13147
rect 3409 12155 3433 12207
rect 3485 12155 3541 12207
rect 3593 12155 3649 12207
rect 3701 12155 3757 12207
rect 3809 12155 3865 12207
rect 3917 12155 3973 12207
rect 4025 12155 4081 12207
rect 4133 12155 4189 12207
rect 4241 12155 4297 12207
rect 4349 12155 4405 12207
rect 4457 12155 4513 12207
rect 4565 12155 4621 12207
rect 4673 12155 4729 12207
rect 4781 12155 4837 12207
rect 4889 12155 4945 12207
rect 4997 12155 5053 12207
rect 5105 12155 5161 12207
rect 5213 12155 5237 12207
rect 3409 11719 5237 12155
rect 3409 11667 3433 11719
rect 3485 11667 3541 11719
rect 3593 11667 3649 11719
rect 3701 11667 3757 11719
rect 3809 11667 3865 11719
rect 3917 11667 3973 11719
rect 4025 11667 4081 11719
rect 4133 11667 4189 11719
rect 4241 11667 4297 11719
rect 4349 11667 4405 11719
rect 4457 11667 4513 11719
rect 4565 11667 4621 11719
rect 4673 11667 4729 11719
rect 4781 11667 4837 11719
rect 4889 11667 4945 11719
rect 4997 11667 5053 11719
rect 5105 11667 5161 11719
rect 5213 11667 5237 11719
rect 3409 11231 5237 11667
rect 3409 11179 3433 11231
rect 3485 11179 3541 11231
rect 3593 11179 3649 11231
rect 3701 11179 3757 11231
rect 3809 11179 3865 11231
rect 3917 11179 3973 11231
rect 4025 11179 4081 11231
rect 4133 11179 4189 11231
rect 4241 11179 4297 11231
rect 4349 11179 4405 11231
rect 4457 11179 4513 11231
rect 4565 11179 4621 11231
rect 4673 11179 4729 11231
rect 4781 11179 4837 11231
rect 4889 11179 4945 11231
rect 4997 11179 5053 11231
rect 5105 11179 5161 11231
rect 5213 11179 5237 11231
rect 3409 10743 5237 11179
rect 3409 10691 3433 10743
rect 3485 10691 3541 10743
rect 3593 10691 3649 10743
rect 3701 10691 3757 10743
rect 3809 10691 3865 10743
rect 3917 10691 3973 10743
rect 4025 10691 4081 10743
rect 4133 10691 4189 10743
rect 4241 10691 4297 10743
rect 4349 10691 4405 10743
rect 4457 10691 4513 10743
rect 4565 10691 4621 10743
rect 4673 10691 4729 10743
rect 4781 10691 4837 10743
rect 4889 10691 4945 10743
rect 4997 10691 5053 10743
rect 5105 10691 5161 10743
rect 5213 10691 5237 10743
rect 3409 10255 5237 10691
rect 3409 10203 3433 10255
rect 3485 10203 3541 10255
rect 3593 10203 3649 10255
rect 3701 10203 3757 10255
rect 3809 10203 3865 10255
rect 3917 10203 3973 10255
rect 4025 10203 4081 10255
rect 4133 10203 4189 10255
rect 4241 10203 4297 10255
rect 4349 10203 4405 10255
rect 4457 10203 4513 10255
rect 4565 10203 4621 10255
rect 4673 10203 4729 10255
rect 4781 10203 4837 10255
rect 4889 10203 4945 10255
rect 4997 10203 5053 10255
rect 5105 10203 5161 10255
rect 5213 10203 5237 10255
rect 3409 9767 5237 10203
rect 3409 9715 3433 9767
rect 3485 9715 3541 9767
rect 3593 9715 3649 9767
rect 3701 9715 3757 9767
rect 3809 9715 3865 9767
rect 3917 9715 3973 9767
rect 4025 9715 4081 9767
rect 4133 9715 4189 9767
rect 4241 9715 4297 9767
rect 4349 9715 4405 9767
rect 4457 9715 4513 9767
rect 4565 9715 4621 9767
rect 4673 9715 4729 9767
rect 4781 9715 4837 9767
rect 4889 9715 4945 9767
rect 4997 9715 5053 9767
rect 5105 9715 5161 9767
rect 5213 9715 5237 9767
rect 3409 9279 5237 9715
rect 3409 9227 3433 9279
rect 3485 9227 3541 9279
rect 3593 9227 3649 9279
rect 3701 9227 3757 9279
rect 3809 9227 3865 9279
rect 3917 9227 3973 9279
rect 4025 9227 4081 9279
rect 4133 9227 4189 9279
rect 4241 9227 4297 9279
rect 4349 9227 4405 9279
rect 4457 9227 4513 9279
rect 4565 9227 4621 9279
rect 4673 9227 4729 9279
rect 4781 9227 4837 9279
rect 4889 9227 4945 9279
rect 4997 9227 5053 9279
rect 5105 9227 5161 9279
rect 5213 9227 5237 9279
rect 3409 8791 5237 9227
rect 3409 8739 3433 8791
rect 3485 8739 3541 8791
rect 3593 8739 3649 8791
rect 3701 8739 3757 8791
rect 3809 8739 3865 8791
rect 3917 8739 3973 8791
rect 4025 8739 4081 8791
rect 4133 8739 4189 8791
rect 4241 8739 4297 8791
rect 4349 8739 4405 8791
rect 4457 8739 4513 8791
rect 4565 8739 4621 8791
rect 4673 8739 4729 8791
rect 4781 8739 4837 8791
rect 4889 8739 4945 8791
rect 4997 8739 5053 8791
rect 5105 8739 5161 8791
rect 5213 8739 5237 8791
rect 3409 8303 5237 8739
rect 3409 8251 3433 8303
rect 3485 8251 3541 8303
rect 3593 8251 3649 8303
rect 3701 8251 3757 8303
rect 3809 8251 3865 8303
rect 3917 8251 3973 8303
rect 4025 8251 4081 8303
rect 4133 8251 4189 8303
rect 4241 8251 4297 8303
rect 4349 8251 4405 8303
rect 4457 8251 4513 8303
rect 4565 8251 4621 8303
rect 4673 8251 4729 8303
rect 4781 8251 4837 8303
rect 4889 8251 4945 8303
rect 4997 8251 5053 8303
rect 5105 8251 5161 8303
rect 5213 8251 5237 8303
rect 3409 7815 5237 8251
rect 3409 7763 3433 7815
rect 3485 7763 3541 7815
rect 3593 7763 3649 7815
rect 3701 7763 3757 7815
rect 3809 7763 3865 7815
rect 3917 7763 3973 7815
rect 4025 7763 4081 7815
rect 4133 7763 4189 7815
rect 4241 7763 4297 7815
rect 4349 7763 4405 7815
rect 4457 7763 4513 7815
rect 4565 7763 4621 7815
rect 4673 7763 4729 7815
rect 4781 7763 4837 7815
rect 4889 7763 4945 7815
rect 4997 7763 5053 7815
rect 5105 7763 5161 7815
rect 5213 7763 5237 7815
rect 3409 7327 5237 7763
rect 3409 7275 3433 7327
rect 3485 7275 3541 7327
rect 3593 7275 3649 7327
rect 3701 7275 3757 7327
rect 3809 7275 3865 7327
rect 3917 7275 3973 7327
rect 4025 7275 4081 7327
rect 4133 7275 4189 7327
rect 4241 7275 4297 7327
rect 4349 7275 4405 7327
rect 4457 7275 4513 7327
rect 4565 7275 4621 7327
rect 4673 7275 4729 7327
rect 4781 7275 4837 7327
rect 4889 7275 4945 7327
rect 4997 7275 5053 7327
rect 5105 7275 5161 7327
rect 5213 7275 5237 7327
rect 3409 6335 5237 7275
rect 3409 6283 3433 6335
rect 3485 6283 3541 6335
rect 3593 6283 3649 6335
rect 3701 6283 3757 6335
rect 3809 6283 3865 6335
rect 3917 6283 3973 6335
rect 4025 6283 4081 6335
rect 4133 6283 4189 6335
rect 4241 6283 4297 6335
rect 4349 6283 4405 6335
rect 4457 6283 4513 6335
rect 4565 6283 4621 6335
rect 4673 6283 4729 6335
rect 4781 6283 4837 6335
rect 4889 6283 4945 6335
rect 4997 6283 5053 6335
rect 5105 6283 5161 6335
rect 5213 6283 5237 6335
rect 3409 5847 5237 6283
rect 3409 5795 3433 5847
rect 3485 5795 3541 5847
rect 3593 5795 3649 5847
rect 3701 5795 3757 5847
rect 3809 5795 3865 5847
rect 3917 5795 3973 5847
rect 4025 5795 4081 5847
rect 4133 5795 4189 5847
rect 4241 5795 4297 5847
rect 4349 5795 4405 5847
rect 4457 5795 4513 5847
rect 4565 5795 4621 5847
rect 4673 5795 4729 5847
rect 4781 5795 4837 5847
rect 4889 5795 4945 5847
rect 4997 5795 5053 5847
rect 5105 5795 5161 5847
rect 5213 5795 5237 5847
rect 3409 5359 5237 5795
rect 3409 5307 3433 5359
rect 3485 5307 3541 5359
rect 3593 5307 3649 5359
rect 3701 5307 3757 5359
rect 3809 5307 3865 5359
rect 3917 5307 3973 5359
rect 4025 5307 4081 5359
rect 4133 5307 4189 5359
rect 4241 5307 4297 5359
rect 4349 5307 4405 5359
rect 4457 5307 4513 5359
rect 4565 5307 4621 5359
rect 4673 5307 4729 5359
rect 4781 5307 4837 5359
rect 4889 5307 4945 5359
rect 4997 5307 5053 5359
rect 5105 5307 5161 5359
rect 5213 5307 5237 5359
rect 3409 4871 5237 5307
rect 3409 4819 3433 4871
rect 3485 4819 3541 4871
rect 3593 4819 3649 4871
rect 3701 4819 3757 4871
rect 3809 4819 3865 4871
rect 3917 4819 3973 4871
rect 4025 4819 4081 4871
rect 4133 4819 4189 4871
rect 4241 4819 4297 4871
rect 4349 4819 4405 4871
rect 4457 4819 4513 4871
rect 4565 4819 4621 4871
rect 4673 4819 4729 4871
rect 4781 4819 4837 4871
rect 4889 4819 4945 4871
rect 4997 4819 5053 4871
rect 5105 4819 5161 4871
rect 5213 4819 5237 4871
rect 3409 4383 5237 4819
rect 3409 4331 3433 4383
rect 3485 4331 3541 4383
rect 3593 4331 3649 4383
rect 3701 4331 3757 4383
rect 3809 4331 3865 4383
rect 3917 4331 3973 4383
rect 4025 4331 4081 4383
rect 4133 4331 4189 4383
rect 4241 4331 4297 4383
rect 4349 4331 4405 4383
rect 4457 4331 4513 4383
rect 4565 4331 4621 4383
rect 4673 4331 4729 4383
rect 4781 4331 4837 4383
rect 4889 4331 4945 4383
rect 4997 4331 5053 4383
rect 5105 4331 5161 4383
rect 5213 4331 5237 4383
rect 3409 3895 5237 4331
rect 3409 3843 3433 3895
rect 3485 3843 3541 3895
rect 3593 3843 3649 3895
rect 3701 3843 3757 3895
rect 3809 3843 3865 3895
rect 3917 3843 3973 3895
rect 4025 3843 4081 3895
rect 4133 3843 4189 3895
rect 4241 3843 4297 3895
rect 4349 3843 4405 3895
rect 4457 3843 4513 3895
rect 4565 3843 4621 3895
rect 4673 3843 4729 3895
rect 4781 3843 4837 3895
rect 4889 3843 4945 3895
rect 4997 3843 5053 3895
rect 5105 3843 5161 3895
rect 5213 3843 5237 3895
rect 3409 3407 5237 3843
rect 3409 3355 3433 3407
rect 3485 3355 3541 3407
rect 3593 3355 3649 3407
rect 3701 3355 3757 3407
rect 3809 3355 3865 3407
rect 3917 3355 3973 3407
rect 4025 3355 4081 3407
rect 4133 3355 4189 3407
rect 4241 3355 4297 3407
rect 4349 3355 4405 3407
rect 4457 3355 4513 3407
rect 4565 3355 4621 3407
rect 4673 3355 4729 3407
rect 4781 3355 4837 3407
rect 4889 3355 4945 3407
rect 4997 3355 5053 3407
rect 5105 3355 5161 3407
rect 5213 3355 5237 3407
rect 3409 2919 5237 3355
rect 3409 2867 3433 2919
rect 3485 2867 3541 2919
rect 3593 2867 3649 2919
rect 3701 2867 3757 2919
rect 3809 2867 3865 2919
rect 3917 2867 3973 2919
rect 4025 2867 4081 2919
rect 4133 2867 4189 2919
rect 4241 2867 4297 2919
rect 4349 2867 4405 2919
rect 4457 2867 4513 2919
rect 4565 2867 4621 2919
rect 4673 2867 4729 2919
rect 4781 2867 4837 2919
rect 4889 2867 4945 2919
rect 4997 2867 5053 2919
rect 5105 2867 5161 2919
rect 5213 2867 5237 2919
rect 3409 2431 5237 2867
rect 3409 2379 3433 2431
rect 3485 2379 3541 2431
rect 3593 2379 3649 2431
rect 3701 2379 3757 2431
rect 3809 2379 3865 2431
rect 3917 2379 3973 2431
rect 4025 2379 4081 2431
rect 4133 2379 4189 2431
rect 4241 2379 4297 2431
rect 4349 2379 4405 2431
rect 4457 2379 4513 2431
rect 4565 2379 4621 2431
rect 4673 2379 4729 2431
rect 4781 2379 4837 2431
rect 4889 2379 4945 2431
rect 4997 2379 5053 2431
rect 5105 2379 5161 2431
rect 5213 2379 5237 2431
rect 3409 1943 5237 2379
rect 3409 1891 3433 1943
rect 3485 1891 3541 1943
rect 3593 1891 3649 1943
rect 3701 1891 3757 1943
rect 3809 1891 3865 1943
rect 3917 1891 3973 1943
rect 4025 1891 4081 1943
rect 4133 1891 4189 1943
rect 4241 1891 4297 1943
rect 4349 1891 4405 1943
rect 4457 1891 4513 1943
rect 4565 1891 4621 1943
rect 4673 1891 4729 1943
rect 4781 1891 4837 1943
rect 4889 1891 4945 1943
rect 4997 1891 5053 1943
rect 5105 1891 5161 1943
rect 5213 1891 5237 1943
rect 3409 1455 5237 1891
rect 3409 1403 3433 1455
rect 3485 1403 3541 1455
rect 3593 1403 3649 1455
rect 3701 1403 3757 1455
rect 3809 1403 3865 1455
rect 3917 1403 3973 1455
rect 4025 1403 4081 1455
rect 4133 1403 4189 1455
rect 4241 1403 4297 1455
rect 4349 1403 4405 1455
rect 4457 1403 4513 1455
rect 4565 1403 4621 1455
rect 4673 1403 4729 1455
rect 4781 1403 4837 1455
rect 4889 1403 4945 1455
rect 4997 1403 5053 1455
rect 5105 1403 5161 1455
rect 5213 1403 5237 1455
rect 3409 361 5237 1403
rect 3409 309 3433 361
rect 3485 309 3541 361
rect 3593 309 3649 361
rect 3701 309 3757 361
rect 3809 309 3865 361
rect 3917 309 3973 361
rect 4025 309 4081 361
rect 4133 309 4189 361
rect 4241 309 4297 361
rect 4349 309 4405 361
rect 4457 309 4513 361
rect 4565 309 4621 361
rect 4673 309 4729 361
rect 4781 309 4837 361
rect 4889 309 4945 361
rect 4997 309 5053 361
rect 5105 309 5161 361
rect 5213 309 5237 361
rect 3409 253 5237 309
rect 3409 201 3433 253
rect 3485 201 3541 253
rect 3593 201 3649 253
rect 3701 201 3757 253
rect 3809 201 3865 253
rect 3917 201 3973 253
rect 4025 201 4081 253
rect 4133 201 4189 253
rect 4241 201 4297 253
rect 4349 201 4405 253
rect 4457 201 4513 253
rect 4565 201 4621 253
rect 4673 201 4729 253
rect 4781 201 4837 253
rect 4889 201 4945 253
rect 4997 201 5053 253
rect 5105 201 5161 253
rect 5213 201 5237 253
rect 3409 145 5237 201
rect 3409 93 3433 145
rect 3485 93 3541 145
rect 3593 93 3649 145
rect 3701 93 3757 145
rect 3809 93 3865 145
rect 3917 93 3973 145
rect 4025 93 4081 145
rect 4133 93 4189 145
rect 4241 93 4297 145
rect 4349 93 4405 145
rect 4457 93 4513 145
rect 4565 93 4621 145
rect 4673 93 4729 145
rect 4781 93 4837 145
rect 4889 93 4945 145
rect 4997 93 5053 145
rect 5105 93 5161 145
rect 5213 93 5237 145
rect 3409 43 5237 93
rect 5337 24661 6431 25617
rect 5337 24609 5372 24661
rect 5424 24609 5480 24661
rect 5532 24609 5588 24661
rect 5640 24609 5696 24661
rect 5748 24609 5804 24661
rect 5856 24609 5912 24661
rect 5964 24609 6020 24661
rect 6072 24609 6128 24661
rect 6180 24609 6236 24661
rect 6288 24609 6344 24661
rect 6396 24609 6431 24661
rect 5337 24553 6431 24609
rect 5337 24501 5372 24553
rect 5424 24501 5480 24553
rect 5532 24501 5588 24553
rect 5640 24501 5696 24553
rect 5748 24501 5804 24553
rect 5856 24501 5912 24553
rect 5964 24501 6020 24553
rect 6072 24501 6128 24553
rect 6180 24501 6236 24553
rect 6288 24501 6344 24553
rect 6396 24501 6431 24553
rect 5337 24445 6431 24501
rect 5337 24393 5372 24445
rect 5424 24393 5480 24445
rect 5532 24393 5588 24445
rect 5640 24393 5696 24445
rect 5748 24393 5804 24445
rect 5856 24393 5912 24445
rect 5964 24393 6020 24445
rect 6072 24393 6128 24445
rect 6180 24393 6236 24445
rect 6288 24393 6344 24445
rect 6396 24393 6431 24445
rect 5337 23707 6431 24393
rect 5337 23655 5372 23707
rect 5424 23655 5480 23707
rect 5532 23655 5588 23707
rect 5640 23655 5696 23707
rect 5748 23655 5804 23707
rect 5856 23655 5912 23707
rect 5964 23655 6020 23707
rect 6072 23655 6128 23707
rect 6180 23655 6236 23707
rect 6288 23655 6344 23707
rect 6396 23655 6431 23707
rect 5337 23219 6431 23655
rect 5337 23167 5372 23219
rect 5424 23167 5480 23219
rect 5532 23167 5588 23219
rect 5640 23167 5696 23219
rect 5748 23167 5804 23219
rect 5856 23167 5912 23219
rect 5964 23167 6020 23219
rect 6072 23167 6128 23219
rect 6180 23167 6236 23219
rect 6288 23167 6344 23219
rect 6396 23167 6431 23219
rect 5337 22731 6431 23167
rect 5337 22679 5372 22731
rect 5424 22679 5480 22731
rect 5532 22679 5588 22731
rect 5640 22679 5696 22731
rect 5748 22679 5804 22731
rect 5856 22679 5912 22731
rect 5964 22679 6020 22731
rect 6072 22679 6128 22731
rect 6180 22679 6236 22731
rect 6288 22679 6344 22731
rect 6396 22679 6431 22731
rect 5337 22243 6431 22679
rect 5337 22191 5372 22243
rect 5424 22191 5480 22243
rect 5532 22191 5588 22243
rect 5640 22191 5696 22243
rect 5748 22191 5804 22243
rect 5856 22191 5912 22243
rect 5964 22191 6020 22243
rect 6072 22191 6128 22243
rect 6180 22191 6236 22243
rect 6288 22191 6344 22243
rect 6396 22191 6431 22243
rect 5337 21755 6431 22191
rect 5337 21703 5372 21755
rect 5424 21703 5480 21755
rect 5532 21703 5588 21755
rect 5640 21703 5696 21755
rect 5748 21703 5804 21755
rect 5856 21703 5912 21755
rect 5964 21703 6020 21755
rect 6072 21703 6128 21755
rect 6180 21703 6236 21755
rect 6288 21703 6344 21755
rect 6396 21703 6431 21755
rect 5337 21267 6431 21703
rect 5337 21215 5372 21267
rect 5424 21215 5480 21267
rect 5532 21215 5588 21267
rect 5640 21215 5696 21267
rect 5748 21215 5804 21267
rect 5856 21215 5912 21267
rect 5964 21215 6020 21267
rect 6072 21215 6128 21267
rect 6180 21215 6236 21267
rect 6288 21215 6344 21267
rect 6396 21215 6431 21267
rect 5337 20779 6431 21215
rect 5337 20727 5372 20779
rect 5424 20727 5480 20779
rect 5532 20727 5588 20779
rect 5640 20727 5696 20779
rect 5748 20727 5804 20779
rect 5856 20727 5912 20779
rect 5964 20727 6020 20779
rect 6072 20727 6128 20779
rect 6180 20727 6236 20779
rect 6288 20727 6344 20779
rect 6396 20727 6431 20779
rect 5337 20291 6431 20727
rect 5337 20239 5372 20291
rect 5424 20239 5480 20291
rect 5532 20239 5588 20291
rect 5640 20239 5696 20291
rect 5748 20239 5804 20291
rect 5856 20239 5912 20291
rect 5964 20239 6020 20291
rect 6072 20239 6128 20291
rect 6180 20239 6236 20291
rect 6288 20239 6344 20291
rect 6396 20239 6431 20291
rect 5337 19803 6431 20239
rect 5337 19751 5372 19803
rect 5424 19751 5480 19803
rect 5532 19751 5588 19803
rect 5640 19751 5696 19803
rect 5748 19751 5804 19803
rect 5856 19751 5912 19803
rect 5964 19751 6020 19803
rect 6072 19751 6128 19803
rect 6180 19751 6236 19803
rect 6288 19751 6344 19803
rect 6396 19751 6431 19803
rect 5337 19315 6431 19751
rect 5337 19263 5372 19315
rect 5424 19263 5480 19315
rect 5532 19263 5588 19315
rect 5640 19263 5696 19315
rect 5748 19263 5804 19315
rect 5856 19263 5912 19315
rect 5964 19263 6020 19315
rect 6072 19263 6128 19315
rect 6180 19263 6236 19315
rect 6288 19263 6344 19315
rect 6396 19263 6431 19315
rect 5337 18629 6431 19263
rect 5337 18577 5372 18629
rect 5424 18577 5480 18629
rect 5532 18577 5588 18629
rect 5640 18577 5696 18629
rect 5748 18577 5804 18629
rect 5856 18577 5912 18629
rect 5964 18577 6020 18629
rect 6072 18577 6128 18629
rect 6180 18577 6236 18629
rect 6288 18577 6344 18629
rect 6396 18577 6431 18629
rect 5337 18521 6431 18577
rect 5337 18469 5372 18521
rect 5424 18469 5480 18521
rect 5532 18469 5588 18521
rect 5640 18469 5696 18521
rect 5748 18469 5804 18521
rect 5856 18469 5912 18521
rect 5964 18469 6020 18521
rect 6072 18469 6128 18521
rect 6180 18469 6236 18521
rect 6288 18469 6344 18521
rect 6396 18469 6431 18521
rect 5337 17835 6431 18469
rect 5337 17783 5372 17835
rect 5424 17783 5480 17835
rect 5532 17783 5588 17835
rect 5640 17783 5696 17835
rect 5748 17783 5804 17835
rect 5856 17783 5912 17835
rect 5964 17783 6020 17835
rect 6072 17783 6128 17835
rect 6180 17783 6236 17835
rect 6288 17783 6344 17835
rect 6396 17783 6431 17835
rect 5337 17347 6431 17783
rect 5337 17295 5372 17347
rect 5424 17295 5480 17347
rect 5532 17295 5588 17347
rect 5640 17295 5696 17347
rect 5748 17295 5804 17347
rect 5856 17295 5912 17347
rect 5964 17295 6020 17347
rect 6072 17295 6128 17347
rect 6180 17295 6236 17347
rect 6288 17295 6344 17347
rect 6396 17295 6431 17347
rect 5337 16859 6431 17295
rect 5337 16807 5372 16859
rect 5424 16807 5480 16859
rect 5532 16807 5588 16859
rect 5640 16807 5696 16859
rect 5748 16807 5804 16859
rect 5856 16807 5912 16859
rect 5964 16807 6020 16859
rect 6072 16807 6128 16859
rect 6180 16807 6236 16859
rect 6288 16807 6344 16859
rect 6396 16807 6431 16859
rect 5337 16371 6431 16807
rect 5337 16319 5372 16371
rect 5424 16319 5480 16371
rect 5532 16319 5588 16371
rect 5640 16319 5696 16371
rect 5748 16319 5804 16371
rect 5856 16319 5912 16371
rect 5964 16319 6020 16371
rect 6072 16319 6128 16371
rect 6180 16319 6236 16371
rect 6288 16319 6344 16371
rect 6396 16319 6431 16371
rect 5337 15883 6431 16319
rect 5337 15831 5372 15883
rect 5424 15831 5480 15883
rect 5532 15831 5588 15883
rect 5640 15831 5696 15883
rect 5748 15831 5804 15883
rect 5856 15831 5912 15883
rect 5964 15831 6020 15883
rect 6072 15831 6128 15883
rect 6180 15831 6236 15883
rect 6288 15831 6344 15883
rect 6396 15831 6431 15883
rect 5337 15395 6431 15831
rect 5337 15343 5372 15395
rect 5424 15343 5480 15395
rect 5532 15343 5588 15395
rect 5640 15343 5696 15395
rect 5748 15343 5804 15395
rect 5856 15343 5912 15395
rect 5964 15343 6020 15395
rect 6072 15343 6128 15395
rect 6180 15343 6236 15395
rect 6288 15343 6344 15395
rect 6396 15343 6431 15395
rect 5337 14907 6431 15343
rect 5337 14855 5372 14907
rect 5424 14855 5480 14907
rect 5532 14855 5588 14907
rect 5640 14855 5696 14907
rect 5748 14855 5804 14907
rect 5856 14855 5912 14907
rect 5964 14855 6020 14907
rect 6072 14855 6128 14907
rect 6180 14855 6236 14907
rect 6288 14855 6344 14907
rect 6396 14855 6431 14907
rect 5337 14419 6431 14855
rect 5337 14367 5372 14419
rect 5424 14367 5480 14419
rect 5532 14367 5588 14419
rect 5640 14367 5696 14419
rect 5748 14367 5804 14419
rect 5856 14367 5912 14419
rect 5964 14367 6020 14419
rect 6072 14367 6128 14419
rect 6180 14367 6236 14419
rect 6288 14367 6344 14419
rect 6396 14367 6431 14419
rect 5337 13931 6431 14367
rect 5337 13879 5372 13931
rect 5424 13879 5480 13931
rect 5532 13879 5588 13931
rect 5640 13879 5696 13931
rect 5748 13879 5804 13931
rect 5856 13879 5912 13931
rect 5964 13879 6020 13931
rect 6072 13879 6128 13931
rect 6180 13879 6236 13931
rect 6288 13879 6344 13931
rect 6396 13879 6431 13931
rect 5337 13443 6431 13879
rect 5337 13391 5372 13443
rect 5424 13391 5480 13443
rect 5532 13391 5588 13443
rect 5640 13391 5696 13443
rect 5748 13391 5804 13443
rect 5856 13391 5912 13443
rect 5964 13391 6020 13443
rect 6072 13391 6128 13443
rect 6180 13391 6236 13443
rect 6288 13391 6344 13443
rect 6396 13391 6431 13443
rect 5337 12757 6431 13391
rect 5337 12705 5372 12757
rect 5424 12705 5480 12757
rect 5532 12705 5588 12757
rect 5640 12705 5696 12757
rect 5748 12705 5804 12757
rect 5856 12705 5912 12757
rect 5964 12705 6020 12757
rect 6072 12705 6128 12757
rect 6180 12705 6236 12757
rect 6288 12705 6344 12757
rect 6396 12705 6431 12757
rect 5337 12649 6431 12705
rect 5337 12597 5372 12649
rect 5424 12597 5480 12649
rect 5532 12597 5588 12649
rect 5640 12597 5696 12649
rect 5748 12597 5804 12649
rect 5856 12597 5912 12649
rect 5964 12597 6020 12649
rect 6072 12597 6128 12649
rect 6180 12597 6236 12649
rect 6288 12597 6344 12649
rect 6396 12597 6431 12649
rect 5337 11963 6431 12597
rect 5337 11911 5372 11963
rect 5424 11911 5480 11963
rect 5532 11911 5588 11963
rect 5640 11911 5696 11963
rect 5748 11911 5804 11963
rect 5856 11911 5912 11963
rect 5964 11911 6020 11963
rect 6072 11911 6128 11963
rect 6180 11911 6236 11963
rect 6288 11911 6344 11963
rect 6396 11911 6431 11963
rect 5337 11475 6431 11911
rect 5337 11423 5372 11475
rect 5424 11423 5480 11475
rect 5532 11423 5588 11475
rect 5640 11423 5696 11475
rect 5748 11423 5804 11475
rect 5856 11423 5912 11475
rect 5964 11423 6020 11475
rect 6072 11423 6128 11475
rect 6180 11423 6236 11475
rect 6288 11423 6344 11475
rect 6396 11423 6431 11475
rect 5337 10987 6431 11423
rect 5337 10935 5372 10987
rect 5424 10935 5480 10987
rect 5532 10935 5588 10987
rect 5640 10935 5696 10987
rect 5748 10935 5804 10987
rect 5856 10935 5912 10987
rect 5964 10935 6020 10987
rect 6072 10935 6128 10987
rect 6180 10935 6236 10987
rect 6288 10935 6344 10987
rect 6396 10935 6431 10987
rect 5337 10499 6431 10935
rect 5337 10447 5372 10499
rect 5424 10447 5480 10499
rect 5532 10447 5588 10499
rect 5640 10447 5696 10499
rect 5748 10447 5804 10499
rect 5856 10447 5912 10499
rect 5964 10447 6020 10499
rect 6072 10447 6128 10499
rect 6180 10447 6236 10499
rect 6288 10447 6344 10499
rect 6396 10447 6431 10499
rect 5337 10011 6431 10447
rect 5337 9959 5372 10011
rect 5424 9959 5480 10011
rect 5532 9959 5588 10011
rect 5640 9959 5696 10011
rect 5748 9959 5804 10011
rect 5856 9959 5912 10011
rect 5964 9959 6020 10011
rect 6072 9959 6128 10011
rect 6180 9959 6236 10011
rect 6288 9959 6344 10011
rect 6396 9959 6431 10011
rect 5337 9523 6431 9959
rect 5337 9471 5372 9523
rect 5424 9471 5480 9523
rect 5532 9471 5588 9523
rect 5640 9471 5696 9523
rect 5748 9471 5804 9523
rect 5856 9471 5912 9523
rect 5964 9471 6020 9523
rect 6072 9471 6128 9523
rect 6180 9471 6236 9523
rect 6288 9471 6344 9523
rect 6396 9471 6431 9523
rect 5337 9035 6431 9471
rect 5337 8983 5372 9035
rect 5424 8983 5480 9035
rect 5532 8983 5588 9035
rect 5640 8983 5696 9035
rect 5748 8983 5804 9035
rect 5856 8983 5912 9035
rect 5964 8983 6020 9035
rect 6072 8983 6128 9035
rect 6180 8983 6236 9035
rect 6288 8983 6344 9035
rect 6396 8983 6431 9035
rect 5337 8547 6431 8983
rect 5337 8495 5372 8547
rect 5424 8495 5480 8547
rect 5532 8495 5588 8547
rect 5640 8495 5696 8547
rect 5748 8495 5804 8547
rect 5856 8495 5912 8547
rect 5964 8495 6020 8547
rect 6072 8495 6128 8547
rect 6180 8495 6236 8547
rect 6288 8495 6344 8547
rect 6396 8495 6431 8547
rect 5337 8059 6431 8495
rect 5337 8007 5372 8059
rect 5424 8007 5480 8059
rect 5532 8007 5588 8059
rect 5640 8007 5696 8059
rect 5748 8007 5804 8059
rect 5856 8007 5912 8059
rect 5964 8007 6020 8059
rect 6072 8007 6128 8059
rect 6180 8007 6236 8059
rect 6288 8007 6344 8059
rect 6396 8007 6431 8059
rect 5337 7571 6431 8007
rect 5337 7519 5372 7571
rect 5424 7519 5480 7571
rect 5532 7519 5588 7571
rect 5640 7519 5696 7571
rect 5748 7519 5804 7571
rect 5856 7519 5912 7571
rect 5964 7519 6020 7571
rect 6072 7519 6128 7571
rect 6180 7519 6236 7571
rect 6288 7519 6344 7571
rect 6396 7519 6431 7571
rect 5337 6885 6431 7519
rect 5337 6833 5372 6885
rect 5424 6833 5480 6885
rect 5532 6833 5588 6885
rect 5640 6833 5696 6885
rect 5748 6833 5804 6885
rect 5856 6833 5912 6885
rect 5964 6833 6020 6885
rect 6072 6833 6128 6885
rect 6180 6833 6236 6885
rect 6288 6833 6344 6885
rect 6396 6833 6431 6885
rect 5337 6777 6431 6833
rect 5337 6725 5372 6777
rect 5424 6725 5480 6777
rect 5532 6725 5588 6777
rect 5640 6725 5696 6777
rect 5748 6725 5804 6777
rect 5856 6725 5912 6777
rect 5964 6725 6020 6777
rect 6072 6725 6128 6777
rect 6180 6725 6236 6777
rect 6288 6725 6344 6777
rect 6396 6725 6431 6777
rect 5337 6091 6431 6725
rect 5337 6039 5372 6091
rect 5424 6039 5480 6091
rect 5532 6039 5588 6091
rect 5640 6039 5696 6091
rect 5748 6039 5804 6091
rect 5856 6039 5912 6091
rect 5964 6039 6020 6091
rect 6072 6039 6128 6091
rect 6180 6039 6236 6091
rect 6288 6039 6344 6091
rect 6396 6039 6431 6091
rect 5337 5603 6431 6039
rect 5337 5551 5372 5603
rect 5424 5551 5480 5603
rect 5532 5551 5588 5603
rect 5640 5551 5696 5603
rect 5748 5551 5804 5603
rect 5856 5551 5912 5603
rect 5964 5551 6020 5603
rect 6072 5551 6128 5603
rect 6180 5551 6236 5603
rect 6288 5551 6344 5603
rect 6396 5551 6431 5603
rect 5337 5115 6431 5551
rect 5337 5063 5372 5115
rect 5424 5063 5480 5115
rect 5532 5063 5588 5115
rect 5640 5063 5696 5115
rect 5748 5063 5804 5115
rect 5856 5063 5912 5115
rect 5964 5063 6020 5115
rect 6072 5063 6128 5115
rect 6180 5063 6236 5115
rect 6288 5063 6344 5115
rect 6396 5063 6431 5115
rect 5337 4627 6431 5063
rect 5337 4575 5372 4627
rect 5424 4575 5480 4627
rect 5532 4575 5588 4627
rect 5640 4575 5696 4627
rect 5748 4575 5804 4627
rect 5856 4575 5912 4627
rect 5964 4575 6020 4627
rect 6072 4575 6128 4627
rect 6180 4575 6236 4627
rect 6288 4575 6344 4627
rect 6396 4575 6431 4627
rect 5337 4139 6431 4575
rect 5337 4087 5372 4139
rect 5424 4087 5480 4139
rect 5532 4087 5588 4139
rect 5640 4087 5696 4139
rect 5748 4087 5804 4139
rect 5856 4087 5912 4139
rect 5964 4087 6020 4139
rect 6072 4087 6128 4139
rect 6180 4087 6236 4139
rect 6288 4087 6344 4139
rect 6396 4087 6431 4139
rect 5337 3651 6431 4087
rect 5337 3599 5372 3651
rect 5424 3599 5480 3651
rect 5532 3599 5588 3651
rect 5640 3599 5696 3651
rect 5748 3599 5804 3651
rect 5856 3599 5912 3651
rect 5964 3599 6020 3651
rect 6072 3599 6128 3651
rect 6180 3599 6236 3651
rect 6288 3599 6344 3651
rect 6396 3599 6431 3651
rect 5337 3163 6431 3599
rect 5337 3111 5372 3163
rect 5424 3111 5480 3163
rect 5532 3111 5588 3163
rect 5640 3111 5696 3163
rect 5748 3111 5804 3163
rect 5856 3111 5912 3163
rect 5964 3111 6020 3163
rect 6072 3111 6128 3163
rect 6180 3111 6236 3163
rect 6288 3111 6344 3163
rect 6396 3111 6431 3163
rect 5337 2675 6431 3111
rect 5337 2623 5372 2675
rect 5424 2623 5480 2675
rect 5532 2623 5588 2675
rect 5640 2623 5696 2675
rect 5748 2623 5804 2675
rect 5856 2623 5912 2675
rect 5964 2623 6020 2675
rect 6072 2623 6128 2675
rect 6180 2623 6236 2675
rect 6288 2623 6344 2675
rect 6396 2623 6431 2675
rect 5337 2187 6431 2623
rect 5337 2135 5372 2187
rect 5424 2135 5480 2187
rect 5532 2135 5588 2187
rect 5640 2135 5696 2187
rect 5748 2135 5804 2187
rect 5856 2135 5912 2187
rect 5964 2135 6020 2187
rect 6072 2135 6128 2187
rect 6180 2135 6236 2187
rect 6288 2135 6344 2187
rect 6396 2135 6431 2187
rect 5337 1699 6431 2135
rect 5337 1647 5372 1699
rect 5424 1647 5480 1699
rect 5532 1647 5588 1699
rect 5640 1647 5696 1699
rect 5748 1647 5804 1699
rect 5856 1647 5912 1699
rect 5964 1647 6020 1699
rect 6072 1647 6128 1699
rect 6180 1647 6236 1699
rect 6288 1647 6344 1699
rect 6396 1647 6431 1699
rect 5337 961 6431 1647
rect 5337 909 5372 961
rect 5424 909 5480 961
rect 5532 909 5588 961
rect 5640 909 5696 961
rect 5748 909 5804 961
rect 5856 909 5912 961
rect 5964 909 6020 961
rect 6072 909 6128 961
rect 6180 909 6236 961
rect 6288 909 6344 961
rect 6396 909 6431 961
rect 5337 853 6431 909
rect 5337 801 5372 853
rect 5424 801 5480 853
rect 5532 801 5588 853
rect 5640 801 5696 853
rect 5748 801 5804 853
rect 5856 801 5912 853
rect 5964 801 6020 853
rect 6072 801 6128 853
rect 6180 801 6236 853
rect 6288 801 6344 853
rect 6396 801 6431 853
rect 5337 745 6431 801
rect 5337 693 5372 745
rect 5424 693 5480 745
rect 5532 693 5588 745
rect 5640 693 5696 745
rect 5748 693 5804 745
rect 5856 693 5912 745
rect 5964 693 6020 745
rect 6072 693 6128 745
rect 6180 693 6236 745
rect 6288 693 6344 745
rect 6396 693 6431 745
rect 5337 43 6431 693
rect 6531 25261 7625 25617
rect 6531 25209 6566 25261
rect 6618 25209 6674 25261
rect 6726 25209 6782 25261
rect 6834 25209 6890 25261
rect 6942 25209 6998 25261
rect 7050 25209 7106 25261
rect 7158 25209 7214 25261
rect 7266 25209 7322 25261
rect 7374 25209 7430 25261
rect 7482 25209 7538 25261
rect 7590 25209 7625 25261
rect 6531 25153 7625 25209
rect 6531 25101 6566 25153
rect 6618 25101 6674 25153
rect 6726 25101 6782 25153
rect 6834 25101 6890 25153
rect 6942 25101 6998 25153
rect 7050 25101 7106 25153
rect 7158 25101 7214 25153
rect 7266 25101 7322 25153
rect 7374 25101 7430 25153
rect 7482 25101 7538 25153
rect 7590 25101 7625 25153
rect 6531 25045 7625 25101
rect 6531 24993 6566 25045
rect 6618 24993 6674 25045
rect 6726 24993 6782 25045
rect 6834 24993 6890 25045
rect 6942 24993 6998 25045
rect 7050 24993 7106 25045
rect 7158 24993 7214 25045
rect 7266 24993 7322 25045
rect 7374 24993 7430 25045
rect 7482 24993 7538 25045
rect 7590 24993 7625 25045
rect 6531 23951 7625 24993
rect 6531 23899 6566 23951
rect 6618 23899 6674 23951
rect 6726 23899 6782 23951
rect 6834 23899 6890 23951
rect 6942 23899 6998 23951
rect 7050 23899 7106 23951
rect 7158 23899 7214 23951
rect 7266 23899 7322 23951
rect 7374 23899 7430 23951
rect 7482 23899 7538 23951
rect 7590 23899 7625 23951
rect 6531 23463 7625 23899
rect 6531 23411 6566 23463
rect 6618 23411 6674 23463
rect 6726 23411 6782 23463
rect 6834 23411 6890 23463
rect 6942 23411 6998 23463
rect 7050 23411 7106 23463
rect 7158 23411 7214 23463
rect 7266 23411 7322 23463
rect 7374 23411 7430 23463
rect 7482 23411 7538 23463
rect 7590 23411 7625 23463
rect 6531 22975 7625 23411
rect 6531 22923 6566 22975
rect 6618 22923 6674 22975
rect 6726 22923 6782 22975
rect 6834 22923 6890 22975
rect 6942 22923 6998 22975
rect 7050 22923 7106 22975
rect 7158 22923 7214 22975
rect 7266 22923 7322 22975
rect 7374 22923 7430 22975
rect 7482 22923 7538 22975
rect 7590 22923 7625 22975
rect 6531 22487 7625 22923
rect 6531 22435 6566 22487
rect 6618 22435 6674 22487
rect 6726 22435 6782 22487
rect 6834 22435 6890 22487
rect 6942 22435 6998 22487
rect 7050 22435 7106 22487
rect 7158 22435 7214 22487
rect 7266 22435 7322 22487
rect 7374 22435 7430 22487
rect 7482 22435 7538 22487
rect 7590 22435 7625 22487
rect 6531 21999 7625 22435
rect 6531 21947 6566 21999
rect 6618 21947 6674 21999
rect 6726 21947 6782 21999
rect 6834 21947 6890 21999
rect 6942 21947 6998 21999
rect 7050 21947 7106 21999
rect 7158 21947 7214 21999
rect 7266 21947 7322 21999
rect 7374 21947 7430 21999
rect 7482 21947 7538 21999
rect 7590 21947 7625 21999
rect 6531 21511 7625 21947
rect 6531 21459 6566 21511
rect 6618 21459 6674 21511
rect 6726 21459 6782 21511
rect 6834 21459 6890 21511
rect 6942 21459 6998 21511
rect 7050 21459 7106 21511
rect 7158 21459 7214 21511
rect 7266 21459 7322 21511
rect 7374 21459 7430 21511
rect 7482 21459 7538 21511
rect 7590 21459 7625 21511
rect 6531 21023 7625 21459
rect 6531 20971 6566 21023
rect 6618 20971 6674 21023
rect 6726 20971 6782 21023
rect 6834 20971 6890 21023
rect 6942 20971 6998 21023
rect 7050 20971 7106 21023
rect 7158 20971 7214 21023
rect 7266 20971 7322 21023
rect 7374 20971 7430 21023
rect 7482 20971 7538 21023
rect 7590 20971 7625 21023
rect 6531 20535 7625 20971
rect 6531 20483 6566 20535
rect 6618 20483 6674 20535
rect 6726 20483 6782 20535
rect 6834 20483 6890 20535
rect 6942 20483 6998 20535
rect 7050 20483 7106 20535
rect 7158 20483 7214 20535
rect 7266 20483 7322 20535
rect 7374 20483 7430 20535
rect 7482 20483 7538 20535
rect 7590 20483 7625 20535
rect 6531 20047 7625 20483
rect 6531 19995 6566 20047
rect 6618 19995 6674 20047
rect 6726 19995 6782 20047
rect 6834 19995 6890 20047
rect 6942 19995 6998 20047
rect 7050 19995 7106 20047
rect 7158 19995 7214 20047
rect 7266 19995 7322 20047
rect 7374 19995 7430 20047
rect 7482 19995 7538 20047
rect 7590 19995 7625 20047
rect 6531 19559 7625 19995
rect 6531 19507 6566 19559
rect 6618 19507 6674 19559
rect 6726 19507 6782 19559
rect 6834 19507 6890 19559
rect 6942 19507 6998 19559
rect 7050 19507 7106 19559
rect 7158 19507 7214 19559
rect 7266 19507 7322 19559
rect 7374 19507 7430 19559
rect 7482 19507 7538 19559
rect 7590 19507 7625 19559
rect 6531 19071 7625 19507
rect 6531 19019 6566 19071
rect 6618 19019 6674 19071
rect 6726 19019 6782 19071
rect 6834 19019 6890 19071
rect 6942 19019 6998 19071
rect 7050 19019 7106 19071
rect 7158 19019 7214 19071
rect 7266 19019 7322 19071
rect 7374 19019 7430 19071
rect 7482 19019 7538 19071
rect 7590 19019 7625 19071
rect 6531 18079 7625 19019
rect 6531 18027 6566 18079
rect 6618 18027 6674 18079
rect 6726 18027 6782 18079
rect 6834 18027 6890 18079
rect 6942 18027 6998 18079
rect 7050 18027 7106 18079
rect 7158 18027 7214 18079
rect 7266 18027 7322 18079
rect 7374 18027 7430 18079
rect 7482 18027 7538 18079
rect 7590 18027 7625 18079
rect 6531 17591 7625 18027
rect 6531 17539 6566 17591
rect 6618 17539 6674 17591
rect 6726 17539 6782 17591
rect 6834 17539 6890 17591
rect 6942 17539 6998 17591
rect 7050 17539 7106 17591
rect 7158 17539 7214 17591
rect 7266 17539 7322 17591
rect 7374 17539 7430 17591
rect 7482 17539 7538 17591
rect 7590 17539 7625 17591
rect 6531 17103 7625 17539
rect 6531 17051 6566 17103
rect 6618 17051 6674 17103
rect 6726 17051 6782 17103
rect 6834 17051 6890 17103
rect 6942 17051 6998 17103
rect 7050 17051 7106 17103
rect 7158 17051 7214 17103
rect 7266 17051 7322 17103
rect 7374 17051 7430 17103
rect 7482 17051 7538 17103
rect 7590 17051 7625 17103
rect 6531 16615 7625 17051
rect 6531 16563 6566 16615
rect 6618 16563 6674 16615
rect 6726 16563 6782 16615
rect 6834 16563 6890 16615
rect 6942 16563 6998 16615
rect 7050 16563 7106 16615
rect 7158 16563 7214 16615
rect 7266 16563 7322 16615
rect 7374 16563 7430 16615
rect 7482 16563 7538 16615
rect 7590 16563 7625 16615
rect 6531 16127 7625 16563
rect 6531 16075 6566 16127
rect 6618 16075 6674 16127
rect 6726 16075 6782 16127
rect 6834 16075 6890 16127
rect 6942 16075 6998 16127
rect 7050 16075 7106 16127
rect 7158 16075 7214 16127
rect 7266 16075 7322 16127
rect 7374 16075 7430 16127
rect 7482 16075 7538 16127
rect 7590 16075 7625 16127
rect 6531 15639 7625 16075
rect 6531 15587 6566 15639
rect 6618 15587 6674 15639
rect 6726 15587 6782 15639
rect 6834 15587 6890 15639
rect 6942 15587 6998 15639
rect 7050 15587 7106 15639
rect 7158 15587 7214 15639
rect 7266 15587 7322 15639
rect 7374 15587 7430 15639
rect 7482 15587 7538 15639
rect 7590 15587 7625 15639
rect 6531 15151 7625 15587
rect 6531 15099 6566 15151
rect 6618 15099 6674 15151
rect 6726 15099 6782 15151
rect 6834 15099 6890 15151
rect 6942 15099 6998 15151
rect 7050 15099 7106 15151
rect 7158 15099 7214 15151
rect 7266 15099 7322 15151
rect 7374 15099 7430 15151
rect 7482 15099 7538 15151
rect 7590 15099 7625 15151
rect 6531 14663 7625 15099
rect 6531 14611 6566 14663
rect 6618 14611 6674 14663
rect 6726 14611 6782 14663
rect 6834 14611 6890 14663
rect 6942 14611 6998 14663
rect 7050 14611 7106 14663
rect 7158 14611 7214 14663
rect 7266 14611 7322 14663
rect 7374 14611 7430 14663
rect 7482 14611 7538 14663
rect 7590 14611 7625 14663
rect 6531 14175 7625 14611
rect 6531 14123 6566 14175
rect 6618 14123 6674 14175
rect 6726 14123 6782 14175
rect 6834 14123 6890 14175
rect 6942 14123 6998 14175
rect 7050 14123 7106 14175
rect 7158 14123 7214 14175
rect 7266 14123 7322 14175
rect 7374 14123 7430 14175
rect 7482 14123 7538 14175
rect 7590 14123 7625 14175
rect 6531 13687 7625 14123
rect 6531 13635 6566 13687
rect 6618 13635 6674 13687
rect 6726 13635 6782 13687
rect 6834 13635 6890 13687
rect 6942 13635 6998 13687
rect 7050 13635 7106 13687
rect 7158 13635 7214 13687
rect 7266 13635 7322 13687
rect 7374 13635 7430 13687
rect 7482 13635 7538 13687
rect 7590 13635 7625 13687
rect 6531 13199 7625 13635
rect 6531 13147 6566 13199
rect 6618 13147 6674 13199
rect 6726 13147 6782 13199
rect 6834 13147 6890 13199
rect 6942 13147 6998 13199
rect 7050 13147 7106 13199
rect 7158 13147 7214 13199
rect 7266 13147 7322 13199
rect 7374 13147 7430 13199
rect 7482 13147 7538 13199
rect 7590 13147 7625 13199
rect 6531 12207 7625 13147
rect 6531 12155 6566 12207
rect 6618 12155 6674 12207
rect 6726 12155 6782 12207
rect 6834 12155 6890 12207
rect 6942 12155 6998 12207
rect 7050 12155 7106 12207
rect 7158 12155 7214 12207
rect 7266 12155 7322 12207
rect 7374 12155 7430 12207
rect 7482 12155 7538 12207
rect 7590 12155 7625 12207
rect 6531 11719 7625 12155
rect 6531 11667 6566 11719
rect 6618 11667 6674 11719
rect 6726 11667 6782 11719
rect 6834 11667 6890 11719
rect 6942 11667 6998 11719
rect 7050 11667 7106 11719
rect 7158 11667 7214 11719
rect 7266 11667 7322 11719
rect 7374 11667 7430 11719
rect 7482 11667 7538 11719
rect 7590 11667 7625 11719
rect 6531 11231 7625 11667
rect 6531 11179 6566 11231
rect 6618 11179 6674 11231
rect 6726 11179 6782 11231
rect 6834 11179 6890 11231
rect 6942 11179 6998 11231
rect 7050 11179 7106 11231
rect 7158 11179 7214 11231
rect 7266 11179 7322 11231
rect 7374 11179 7430 11231
rect 7482 11179 7538 11231
rect 7590 11179 7625 11231
rect 6531 10743 7625 11179
rect 6531 10691 6566 10743
rect 6618 10691 6674 10743
rect 6726 10691 6782 10743
rect 6834 10691 6890 10743
rect 6942 10691 6998 10743
rect 7050 10691 7106 10743
rect 7158 10691 7214 10743
rect 7266 10691 7322 10743
rect 7374 10691 7430 10743
rect 7482 10691 7538 10743
rect 7590 10691 7625 10743
rect 6531 10255 7625 10691
rect 6531 10203 6566 10255
rect 6618 10203 6674 10255
rect 6726 10203 6782 10255
rect 6834 10203 6890 10255
rect 6942 10203 6998 10255
rect 7050 10203 7106 10255
rect 7158 10203 7214 10255
rect 7266 10203 7322 10255
rect 7374 10203 7430 10255
rect 7482 10203 7538 10255
rect 7590 10203 7625 10255
rect 6531 9767 7625 10203
rect 6531 9715 6566 9767
rect 6618 9715 6674 9767
rect 6726 9715 6782 9767
rect 6834 9715 6890 9767
rect 6942 9715 6998 9767
rect 7050 9715 7106 9767
rect 7158 9715 7214 9767
rect 7266 9715 7322 9767
rect 7374 9715 7430 9767
rect 7482 9715 7538 9767
rect 7590 9715 7625 9767
rect 6531 9279 7625 9715
rect 6531 9227 6566 9279
rect 6618 9227 6674 9279
rect 6726 9227 6782 9279
rect 6834 9227 6890 9279
rect 6942 9227 6998 9279
rect 7050 9227 7106 9279
rect 7158 9227 7214 9279
rect 7266 9227 7322 9279
rect 7374 9227 7430 9279
rect 7482 9227 7538 9279
rect 7590 9227 7625 9279
rect 6531 8791 7625 9227
rect 6531 8739 6566 8791
rect 6618 8739 6674 8791
rect 6726 8739 6782 8791
rect 6834 8739 6890 8791
rect 6942 8739 6998 8791
rect 7050 8739 7106 8791
rect 7158 8739 7214 8791
rect 7266 8739 7322 8791
rect 7374 8739 7430 8791
rect 7482 8739 7538 8791
rect 7590 8739 7625 8791
rect 6531 8303 7625 8739
rect 6531 8251 6566 8303
rect 6618 8251 6674 8303
rect 6726 8251 6782 8303
rect 6834 8251 6890 8303
rect 6942 8251 6998 8303
rect 7050 8251 7106 8303
rect 7158 8251 7214 8303
rect 7266 8251 7322 8303
rect 7374 8251 7430 8303
rect 7482 8251 7538 8303
rect 7590 8251 7625 8303
rect 6531 7815 7625 8251
rect 6531 7763 6566 7815
rect 6618 7763 6674 7815
rect 6726 7763 6782 7815
rect 6834 7763 6890 7815
rect 6942 7763 6998 7815
rect 7050 7763 7106 7815
rect 7158 7763 7214 7815
rect 7266 7763 7322 7815
rect 7374 7763 7430 7815
rect 7482 7763 7538 7815
rect 7590 7763 7625 7815
rect 6531 7327 7625 7763
rect 6531 7275 6566 7327
rect 6618 7275 6674 7327
rect 6726 7275 6782 7327
rect 6834 7275 6890 7327
rect 6942 7275 6998 7327
rect 7050 7275 7106 7327
rect 7158 7275 7214 7327
rect 7266 7275 7322 7327
rect 7374 7275 7430 7327
rect 7482 7275 7538 7327
rect 7590 7275 7625 7327
rect 6531 6335 7625 7275
rect 6531 6283 6566 6335
rect 6618 6283 6674 6335
rect 6726 6283 6782 6335
rect 6834 6283 6890 6335
rect 6942 6283 6998 6335
rect 7050 6283 7106 6335
rect 7158 6283 7214 6335
rect 7266 6283 7322 6335
rect 7374 6283 7430 6335
rect 7482 6283 7538 6335
rect 7590 6283 7625 6335
rect 6531 5847 7625 6283
rect 6531 5795 6566 5847
rect 6618 5795 6674 5847
rect 6726 5795 6782 5847
rect 6834 5795 6890 5847
rect 6942 5795 6998 5847
rect 7050 5795 7106 5847
rect 7158 5795 7214 5847
rect 7266 5795 7322 5847
rect 7374 5795 7430 5847
rect 7482 5795 7538 5847
rect 7590 5795 7625 5847
rect 6531 5359 7625 5795
rect 6531 5307 6566 5359
rect 6618 5307 6674 5359
rect 6726 5307 6782 5359
rect 6834 5307 6890 5359
rect 6942 5307 6998 5359
rect 7050 5307 7106 5359
rect 7158 5307 7214 5359
rect 7266 5307 7322 5359
rect 7374 5307 7430 5359
rect 7482 5307 7538 5359
rect 7590 5307 7625 5359
rect 6531 4871 7625 5307
rect 6531 4819 6566 4871
rect 6618 4819 6674 4871
rect 6726 4819 6782 4871
rect 6834 4819 6890 4871
rect 6942 4819 6998 4871
rect 7050 4819 7106 4871
rect 7158 4819 7214 4871
rect 7266 4819 7322 4871
rect 7374 4819 7430 4871
rect 7482 4819 7538 4871
rect 7590 4819 7625 4871
rect 6531 4383 7625 4819
rect 6531 4331 6566 4383
rect 6618 4331 6674 4383
rect 6726 4331 6782 4383
rect 6834 4331 6890 4383
rect 6942 4331 6998 4383
rect 7050 4331 7106 4383
rect 7158 4331 7214 4383
rect 7266 4331 7322 4383
rect 7374 4331 7430 4383
rect 7482 4331 7538 4383
rect 7590 4331 7625 4383
rect 6531 3895 7625 4331
rect 6531 3843 6566 3895
rect 6618 3843 6674 3895
rect 6726 3843 6782 3895
rect 6834 3843 6890 3895
rect 6942 3843 6998 3895
rect 7050 3843 7106 3895
rect 7158 3843 7214 3895
rect 7266 3843 7322 3895
rect 7374 3843 7430 3895
rect 7482 3843 7538 3895
rect 7590 3843 7625 3895
rect 6531 3407 7625 3843
rect 6531 3355 6566 3407
rect 6618 3355 6674 3407
rect 6726 3355 6782 3407
rect 6834 3355 6890 3407
rect 6942 3355 6998 3407
rect 7050 3355 7106 3407
rect 7158 3355 7214 3407
rect 7266 3355 7322 3407
rect 7374 3355 7430 3407
rect 7482 3355 7538 3407
rect 7590 3355 7625 3407
rect 6531 2919 7625 3355
rect 6531 2867 6566 2919
rect 6618 2867 6674 2919
rect 6726 2867 6782 2919
rect 6834 2867 6890 2919
rect 6942 2867 6998 2919
rect 7050 2867 7106 2919
rect 7158 2867 7214 2919
rect 7266 2867 7322 2919
rect 7374 2867 7430 2919
rect 7482 2867 7538 2919
rect 7590 2867 7625 2919
rect 6531 2431 7625 2867
rect 6531 2379 6566 2431
rect 6618 2379 6674 2431
rect 6726 2379 6782 2431
rect 6834 2379 6890 2431
rect 6942 2379 6998 2431
rect 7050 2379 7106 2431
rect 7158 2379 7214 2431
rect 7266 2379 7322 2431
rect 7374 2379 7430 2431
rect 7482 2379 7538 2431
rect 7590 2379 7625 2431
rect 6531 1943 7625 2379
rect 6531 1891 6566 1943
rect 6618 1891 6674 1943
rect 6726 1891 6782 1943
rect 6834 1891 6890 1943
rect 6942 1891 6998 1943
rect 7050 1891 7106 1943
rect 7158 1891 7214 1943
rect 7266 1891 7322 1943
rect 7374 1891 7430 1943
rect 7482 1891 7538 1943
rect 7590 1891 7625 1943
rect 6531 1455 7625 1891
rect 6531 1403 6566 1455
rect 6618 1403 6674 1455
rect 6726 1403 6782 1455
rect 6834 1403 6890 1455
rect 6942 1403 6998 1455
rect 7050 1403 7106 1455
rect 7158 1403 7214 1455
rect 7266 1403 7322 1455
rect 7374 1403 7430 1455
rect 7482 1403 7538 1455
rect 7590 1403 7625 1455
rect 6531 361 7625 1403
rect 6531 309 6566 361
rect 6618 309 6674 361
rect 6726 309 6782 361
rect 6834 309 6890 361
rect 6942 309 6998 361
rect 7050 309 7106 361
rect 7158 309 7214 361
rect 7266 309 7322 361
rect 7374 309 7430 361
rect 7482 309 7538 361
rect 7590 309 7625 361
rect 6531 253 7625 309
rect 6531 201 6566 253
rect 6618 201 6674 253
rect 6726 201 6782 253
rect 6834 201 6890 253
rect 6942 201 6998 253
rect 7050 201 7106 253
rect 7158 201 7214 253
rect 7266 201 7322 253
rect 7374 201 7430 253
rect 7482 201 7538 253
rect 7590 201 7625 253
rect 6531 145 7625 201
rect 6531 93 6566 145
rect 6618 93 6674 145
rect 6726 93 6782 145
rect 6834 93 6890 145
rect 6942 93 6998 145
rect 7050 93 7106 145
rect 7158 93 7214 145
rect 7266 93 7322 145
rect 7374 93 7430 145
rect 7482 93 7538 145
rect 7590 93 7625 145
rect 6531 43 7625 93
rect 7725 24661 9553 25617
rect 7725 24609 7749 24661
rect 7801 24609 7857 24661
rect 7909 24609 7965 24661
rect 8017 24609 8073 24661
rect 8125 24609 8181 24661
rect 8233 24609 8289 24661
rect 8341 24609 8397 24661
rect 8449 24609 8505 24661
rect 8557 24609 8613 24661
rect 8665 24609 8721 24661
rect 8773 24609 8829 24661
rect 8881 24609 8937 24661
rect 8989 24609 9045 24661
rect 9097 24609 9153 24661
rect 9205 24609 9261 24661
rect 9313 24609 9369 24661
rect 9421 24609 9477 24661
rect 9529 24609 9553 24661
rect 7725 24553 9553 24609
rect 7725 24501 7749 24553
rect 7801 24501 7857 24553
rect 7909 24501 7965 24553
rect 8017 24501 8073 24553
rect 8125 24501 8181 24553
rect 8233 24501 8289 24553
rect 8341 24501 8397 24553
rect 8449 24501 8505 24553
rect 8557 24501 8613 24553
rect 8665 24501 8721 24553
rect 8773 24501 8829 24553
rect 8881 24501 8937 24553
rect 8989 24501 9045 24553
rect 9097 24501 9153 24553
rect 9205 24501 9261 24553
rect 9313 24501 9369 24553
rect 9421 24501 9477 24553
rect 9529 24501 9553 24553
rect 7725 24445 9553 24501
rect 7725 24393 7749 24445
rect 7801 24393 7857 24445
rect 7909 24393 7965 24445
rect 8017 24393 8073 24445
rect 8125 24393 8181 24445
rect 8233 24393 8289 24445
rect 8341 24393 8397 24445
rect 8449 24393 8505 24445
rect 8557 24393 8613 24445
rect 8665 24393 8721 24445
rect 8773 24393 8829 24445
rect 8881 24393 8937 24445
rect 8989 24393 9045 24445
rect 9097 24393 9153 24445
rect 9205 24393 9261 24445
rect 9313 24393 9369 24445
rect 9421 24393 9477 24445
rect 9529 24393 9553 24445
rect 7725 23707 9553 24393
rect 7725 23655 7749 23707
rect 7801 23655 7857 23707
rect 7909 23655 7965 23707
rect 8017 23655 8073 23707
rect 8125 23655 8181 23707
rect 8233 23655 8289 23707
rect 8341 23655 8397 23707
rect 8449 23655 8505 23707
rect 8557 23655 8613 23707
rect 8665 23655 8721 23707
rect 8773 23655 8829 23707
rect 8881 23655 8937 23707
rect 8989 23655 9045 23707
rect 9097 23655 9153 23707
rect 9205 23655 9261 23707
rect 9313 23655 9369 23707
rect 9421 23655 9477 23707
rect 9529 23655 9553 23707
rect 7725 23219 9553 23655
rect 7725 23167 7749 23219
rect 7801 23167 7857 23219
rect 7909 23167 7965 23219
rect 8017 23167 8073 23219
rect 8125 23167 8181 23219
rect 8233 23167 8289 23219
rect 8341 23167 8397 23219
rect 8449 23167 8505 23219
rect 8557 23167 8613 23219
rect 8665 23167 8721 23219
rect 8773 23167 8829 23219
rect 8881 23167 8937 23219
rect 8989 23167 9045 23219
rect 9097 23167 9153 23219
rect 9205 23167 9261 23219
rect 9313 23167 9369 23219
rect 9421 23167 9477 23219
rect 9529 23167 9553 23219
rect 7725 22731 9553 23167
rect 7725 22679 7749 22731
rect 7801 22679 7857 22731
rect 7909 22679 7965 22731
rect 8017 22679 8073 22731
rect 8125 22679 8181 22731
rect 8233 22679 8289 22731
rect 8341 22679 8397 22731
rect 8449 22679 8505 22731
rect 8557 22679 8613 22731
rect 8665 22679 8721 22731
rect 8773 22679 8829 22731
rect 8881 22679 8937 22731
rect 8989 22679 9045 22731
rect 9097 22679 9153 22731
rect 9205 22679 9261 22731
rect 9313 22679 9369 22731
rect 9421 22679 9477 22731
rect 9529 22679 9553 22731
rect 7725 22243 9553 22679
rect 7725 22191 7749 22243
rect 7801 22191 7857 22243
rect 7909 22191 7965 22243
rect 8017 22191 8073 22243
rect 8125 22191 8181 22243
rect 8233 22191 8289 22243
rect 8341 22191 8397 22243
rect 8449 22191 8505 22243
rect 8557 22191 8613 22243
rect 8665 22191 8721 22243
rect 8773 22191 8829 22243
rect 8881 22191 8937 22243
rect 8989 22191 9045 22243
rect 9097 22191 9153 22243
rect 9205 22191 9261 22243
rect 9313 22191 9369 22243
rect 9421 22191 9477 22243
rect 9529 22191 9553 22243
rect 7725 21755 9553 22191
rect 7725 21703 7749 21755
rect 7801 21703 7857 21755
rect 7909 21703 7965 21755
rect 8017 21703 8073 21755
rect 8125 21703 8181 21755
rect 8233 21703 8289 21755
rect 8341 21703 8397 21755
rect 8449 21703 8505 21755
rect 8557 21703 8613 21755
rect 8665 21703 8721 21755
rect 8773 21703 8829 21755
rect 8881 21703 8937 21755
rect 8989 21703 9045 21755
rect 9097 21703 9153 21755
rect 9205 21703 9261 21755
rect 9313 21703 9369 21755
rect 9421 21703 9477 21755
rect 9529 21703 9553 21755
rect 7725 21267 9553 21703
rect 7725 21215 7749 21267
rect 7801 21215 7857 21267
rect 7909 21215 7965 21267
rect 8017 21215 8073 21267
rect 8125 21215 8181 21267
rect 8233 21215 8289 21267
rect 8341 21215 8397 21267
rect 8449 21215 8505 21267
rect 8557 21215 8613 21267
rect 8665 21215 8721 21267
rect 8773 21215 8829 21267
rect 8881 21215 8937 21267
rect 8989 21215 9045 21267
rect 9097 21215 9153 21267
rect 9205 21215 9261 21267
rect 9313 21215 9369 21267
rect 9421 21215 9477 21267
rect 9529 21215 9553 21267
rect 7725 20779 9553 21215
rect 7725 20727 7749 20779
rect 7801 20727 7857 20779
rect 7909 20727 7965 20779
rect 8017 20727 8073 20779
rect 8125 20727 8181 20779
rect 8233 20727 8289 20779
rect 8341 20727 8397 20779
rect 8449 20727 8505 20779
rect 8557 20727 8613 20779
rect 8665 20727 8721 20779
rect 8773 20727 8829 20779
rect 8881 20727 8937 20779
rect 8989 20727 9045 20779
rect 9097 20727 9153 20779
rect 9205 20727 9261 20779
rect 9313 20727 9369 20779
rect 9421 20727 9477 20779
rect 9529 20727 9553 20779
rect 7725 20291 9553 20727
rect 7725 20239 7749 20291
rect 7801 20239 7857 20291
rect 7909 20239 7965 20291
rect 8017 20239 8073 20291
rect 8125 20239 8181 20291
rect 8233 20239 8289 20291
rect 8341 20239 8397 20291
rect 8449 20239 8505 20291
rect 8557 20239 8613 20291
rect 8665 20239 8721 20291
rect 8773 20239 8829 20291
rect 8881 20239 8937 20291
rect 8989 20239 9045 20291
rect 9097 20239 9153 20291
rect 9205 20239 9261 20291
rect 9313 20239 9369 20291
rect 9421 20239 9477 20291
rect 9529 20239 9553 20291
rect 7725 19803 9553 20239
rect 7725 19751 7749 19803
rect 7801 19751 7857 19803
rect 7909 19751 7965 19803
rect 8017 19751 8073 19803
rect 8125 19751 8181 19803
rect 8233 19751 8289 19803
rect 8341 19751 8397 19803
rect 8449 19751 8505 19803
rect 8557 19751 8613 19803
rect 8665 19751 8721 19803
rect 8773 19751 8829 19803
rect 8881 19751 8937 19803
rect 8989 19751 9045 19803
rect 9097 19751 9153 19803
rect 9205 19751 9261 19803
rect 9313 19751 9369 19803
rect 9421 19751 9477 19803
rect 9529 19751 9553 19803
rect 7725 19315 9553 19751
rect 7725 19263 7749 19315
rect 7801 19263 7857 19315
rect 7909 19263 7965 19315
rect 8017 19263 8073 19315
rect 8125 19263 8181 19315
rect 8233 19263 8289 19315
rect 8341 19263 8397 19315
rect 8449 19263 8505 19315
rect 8557 19263 8613 19315
rect 8665 19263 8721 19315
rect 8773 19263 8829 19315
rect 8881 19263 8937 19315
rect 8989 19263 9045 19315
rect 9097 19263 9153 19315
rect 9205 19263 9261 19315
rect 9313 19263 9369 19315
rect 9421 19263 9477 19315
rect 9529 19263 9553 19315
rect 7725 18629 9553 19263
rect 7725 18577 7749 18629
rect 7801 18577 7857 18629
rect 7909 18577 7965 18629
rect 8017 18577 8073 18629
rect 8125 18577 8181 18629
rect 8233 18577 8289 18629
rect 8341 18577 8397 18629
rect 8449 18577 8505 18629
rect 8557 18577 8613 18629
rect 8665 18577 8721 18629
rect 8773 18577 8829 18629
rect 8881 18577 8937 18629
rect 8989 18577 9045 18629
rect 9097 18577 9153 18629
rect 9205 18577 9261 18629
rect 9313 18577 9369 18629
rect 9421 18577 9477 18629
rect 9529 18577 9553 18629
rect 7725 18521 9553 18577
rect 7725 18469 7749 18521
rect 7801 18469 7857 18521
rect 7909 18469 7965 18521
rect 8017 18469 8073 18521
rect 8125 18469 8181 18521
rect 8233 18469 8289 18521
rect 8341 18469 8397 18521
rect 8449 18469 8505 18521
rect 8557 18469 8613 18521
rect 8665 18469 8721 18521
rect 8773 18469 8829 18521
rect 8881 18469 8937 18521
rect 8989 18469 9045 18521
rect 9097 18469 9153 18521
rect 9205 18469 9261 18521
rect 9313 18469 9369 18521
rect 9421 18469 9477 18521
rect 9529 18469 9553 18521
rect 7725 17835 9553 18469
rect 7725 17783 7749 17835
rect 7801 17783 7857 17835
rect 7909 17783 7965 17835
rect 8017 17783 8073 17835
rect 8125 17783 8181 17835
rect 8233 17783 8289 17835
rect 8341 17783 8397 17835
rect 8449 17783 8505 17835
rect 8557 17783 8613 17835
rect 8665 17783 8721 17835
rect 8773 17783 8829 17835
rect 8881 17783 8937 17835
rect 8989 17783 9045 17835
rect 9097 17783 9153 17835
rect 9205 17783 9261 17835
rect 9313 17783 9369 17835
rect 9421 17783 9477 17835
rect 9529 17783 9553 17835
rect 7725 17347 9553 17783
rect 7725 17295 7749 17347
rect 7801 17295 7857 17347
rect 7909 17295 7965 17347
rect 8017 17295 8073 17347
rect 8125 17295 8181 17347
rect 8233 17295 8289 17347
rect 8341 17295 8397 17347
rect 8449 17295 8505 17347
rect 8557 17295 8613 17347
rect 8665 17295 8721 17347
rect 8773 17295 8829 17347
rect 8881 17295 8937 17347
rect 8989 17295 9045 17347
rect 9097 17295 9153 17347
rect 9205 17295 9261 17347
rect 9313 17295 9369 17347
rect 9421 17295 9477 17347
rect 9529 17295 9553 17347
rect 7725 16859 9553 17295
rect 7725 16807 7749 16859
rect 7801 16807 7857 16859
rect 7909 16807 7965 16859
rect 8017 16807 8073 16859
rect 8125 16807 8181 16859
rect 8233 16807 8289 16859
rect 8341 16807 8397 16859
rect 8449 16807 8505 16859
rect 8557 16807 8613 16859
rect 8665 16807 8721 16859
rect 8773 16807 8829 16859
rect 8881 16807 8937 16859
rect 8989 16807 9045 16859
rect 9097 16807 9153 16859
rect 9205 16807 9261 16859
rect 9313 16807 9369 16859
rect 9421 16807 9477 16859
rect 9529 16807 9553 16859
rect 7725 16371 9553 16807
rect 7725 16319 7749 16371
rect 7801 16319 7857 16371
rect 7909 16319 7965 16371
rect 8017 16319 8073 16371
rect 8125 16319 8181 16371
rect 8233 16319 8289 16371
rect 8341 16319 8397 16371
rect 8449 16319 8505 16371
rect 8557 16319 8613 16371
rect 8665 16319 8721 16371
rect 8773 16319 8829 16371
rect 8881 16319 8937 16371
rect 8989 16319 9045 16371
rect 9097 16319 9153 16371
rect 9205 16319 9261 16371
rect 9313 16319 9369 16371
rect 9421 16319 9477 16371
rect 9529 16319 9553 16371
rect 7725 15883 9553 16319
rect 7725 15831 7749 15883
rect 7801 15831 7857 15883
rect 7909 15831 7965 15883
rect 8017 15831 8073 15883
rect 8125 15831 8181 15883
rect 8233 15831 8289 15883
rect 8341 15831 8397 15883
rect 8449 15831 8505 15883
rect 8557 15831 8613 15883
rect 8665 15831 8721 15883
rect 8773 15831 8829 15883
rect 8881 15831 8937 15883
rect 8989 15831 9045 15883
rect 9097 15831 9153 15883
rect 9205 15831 9261 15883
rect 9313 15831 9369 15883
rect 9421 15831 9477 15883
rect 9529 15831 9553 15883
rect 7725 15395 9553 15831
rect 7725 15343 7749 15395
rect 7801 15343 7857 15395
rect 7909 15343 7965 15395
rect 8017 15343 8073 15395
rect 8125 15343 8181 15395
rect 8233 15343 8289 15395
rect 8341 15343 8397 15395
rect 8449 15343 8505 15395
rect 8557 15343 8613 15395
rect 8665 15343 8721 15395
rect 8773 15343 8829 15395
rect 8881 15343 8937 15395
rect 8989 15343 9045 15395
rect 9097 15343 9153 15395
rect 9205 15343 9261 15395
rect 9313 15343 9369 15395
rect 9421 15343 9477 15395
rect 9529 15343 9553 15395
rect 7725 14907 9553 15343
rect 7725 14855 7749 14907
rect 7801 14855 7857 14907
rect 7909 14855 7965 14907
rect 8017 14855 8073 14907
rect 8125 14855 8181 14907
rect 8233 14855 8289 14907
rect 8341 14855 8397 14907
rect 8449 14855 8505 14907
rect 8557 14855 8613 14907
rect 8665 14855 8721 14907
rect 8773 14855 8829 14907
rect 8881 14855 8937 14907
rect 8989 14855 9045 14907
rect 9097 14855 9153 14907
rect 9205 14855 9261 14907
rect 9313 14855 9369 14907
rect 9421 14855 9477 14907
rect 9529 14855 9553 14907
rect 7725 14419 9553 14855
rect 7725 14367 7749 14419
rect 7801 14367 7857 14419
rect 7909 14367 7965 14419
rect 8017 14367 8073 14419
rect 8125 14367 8181 14419
rect 8233 14367 8289 14419
rect 8341 14367 8397 14419
rect 8449 14367 8505 14419
rect 8557 14367 8613 14419
rect 8665 14367 8721 14419
rect 8773 14367 8829 14419
rect 8881 14367 8937 14419
rect 8989 14367 9045 14419
rect 9097 14367 9153 14419
rect 9205 14367 9261 14419
rect 9313 14367 9369 14419
rect 9421 14367 9477 14419
rect 9529 14367 9553 14419
rect 7725 13931 9553 14367
rect 7725 13879 7749 13931
rect 7801 13879 7857 13931
rect 7909 13879 7965 13931
rect 8017 13879 8073 13931
rect 8125 13879 8181 13931
rect 8233 13879 8289 13931
rect 8341 13879 8397 13931
rect 8449 13879 8505 13931
rect 8557 13879 8613 13931
rect 8665 13879 8721 13931
rect 8773 13879 8829 13931
rect 8881 13879 8937 13931
rect 8989 13879 9045 13931
rect 9097 13879 9153 13931
rect 9205 13879 9261 13931
rect 9313 13879 9369 13931
rect 9421 13879 9477 13931
rect 9529 13879 9553 13931
rect 7725 13443 9553 13879
rect 7725 13391 7749 13443
rect 7801 13391 7857 13443
rect 7909 13391 7965 13443
rect 8017 13391 8073 13443
rect 8125 13391 8181 13443
rect 8233 13391 8289 13443
rect 8341 13391 8397 13443
rect 8449 13391 8505 13443
rect 8557 13391 8613 13443
rect 8665 13391 8721 13443
rect 8773 13391 8829 13443
rect 8881 13391 8937 13443
rect 8989 13391 9045 13443
rect 9097 13391 9153 13443
rect 9205 13391 9261 13443
rect 9313 13391 9369 13443
rect 9421 13391 9477 13443
rect 9529 13391 9553 13443
rect 7725 12757 9553 13391
rect 7725 12705 7749 12757
rect 7801 12705 7857 12757
rect 7909 12705 7965 12757
rect 8017 12705 8073 12757
rect 8125 12705 8181 12757
rect 8233 12705 8289 12757
rect 8341 12705 8397 12757
rect 8449 12705 8505 12757
rect 8557 12705 8613 12757
rect 8665 12705 8721 12757
rect 8773 12705 8829 12757
rect 8881 12705 8937 12757
rect 8989 12705 9045 12757
rect 9097 12705 9153 12757
rect 9205 12705 9261 12757
rect 9313 12705 9369 12757
rect 9421 12705 9477 12757
rect 9529 12705 9553 12757
rect 7725 12649 9553 12705
rect 7725 12597 7749 12649
rect 7801 12597 7857 12649
rect 7909 12597 7965 12649
rect 8017 12597 8073 12649
rect 8125 12597 8181 12649
rect 8233 12597 8289 12649
rect 8341 12597 8397 12649
rect 8449 12597 8505 12649
rect 8557 12597 8613 12649
rect 8665 12597 8721 12649
rect 8773 12597 8829 12649
rect 8881 12597 8937 12649
rect 8989 12597 9045 12649
rect 9097 12597 9153 12649
rect 9205 12597 9261 12649
rect 9313 12597 9369 12649
rect 9421 12597 9477 12649
rect 9529 12597 9553 12649
rect 7725 11963 9553 12597
rect 7725 11911 7749 11963
rect 7801 11911 7857 11963
rect 7909 11911 7965 11963
rect 8017 11911 8073 11963
rect 8125 11911 8181 11963
rect 8233 11911 8289 11963
rect 8341 11911 8397 11963
rect 8449 11911 8505 11963
rect 8557 11911 8613 11963
rect 8665 11911 8721 11963
rect 8773 11911 8829 11963
rect 8881 11911 8937 11963
rect 8989 11911 9045 11963
rect 9097 11911 9153 11963
rect 9205 11911 9261 11963
rect 9313 11911 9369 11963
rect 9421 11911 9477 11963
rect 9529 11911 9553 11963
rect 7725 11475 9553 11911
rect 7725 11423 7749 11475
rect 7801 11423 7857 11475
rect 7909 11423 7965 11475
rect 8017 11423 8073 11475
rect 8125 11423 8181 11475
rect 8233 11423 8289 11475
rect 8341 11423 8397 11475
rect 8449 11423 8505 11475
rect 8557 11423 8613 11475
rect 8665 11423 8721 11475
rect 8773 11423 8829 11475
rect 8881 11423 8937 11475
rect 8989 11423 9045 11475
rect 9097 11423 9153 11475
rect 9205 11423 9261 11475
rect 9313 11423 9369 11475
rect 9421 11423 9477 11475
rect 9529 11423 9553 11475
rect 7725 10987 9553 11423
rect 7725 10935 7749 10987
rect 7801 10935 7857 10987
rect 7909 10935 7965 10987
rect 8017 10935 8073 10987
rect 8125 10935 8181 10987
rect 8233 10935 8289 10987
rect 8341 10935 8397 10987
rect 8449 10935 8505 10987
rect 8557 10935 8613 10987
rect 8665 10935 8721 10987
rect 8773 10935 8829 10987
rect 8881 10935 8937 10987
rect 8989 10935 9045 10987
rect 9097 10935 9153 10987
rect 9205 10935 9261 10987
rect 9313 10935 9369 10987
rect 9421 10935 9477 10987
rect 9529 10935 9553 10987
rect 7725 10499 9553 10935
rect 7725 10447 7749 10499
rect 7801 10447 7857 10499
rect 7909 10447 7965 10499
rect 8017 10447 8073 10499
rect 8125 10447 8181 10499
rect 8233 10447 8289 10499
rect 8341 10447 8397 10499
rect 8449 10447 8505 10499
rect 8557 10447 8613 10499
rect 8665 10447 8721 10499
rect 8773 10447 8829 10499
rect 8881 10447 8937 10499
rect 8989 10447 9045 10499
rect 9097 10447 9153 10499
rect 9205 10447 9261 10499
rect 9313 10447 9369 10499
rect 9421 10447 9477 10499
rect 9529 10447 9553 10499
rect 7725 10011 9553 10447
rect 7725 9959 7749 10011
rect 7801 9959 7857 10011
rect 7909 9959 7965 10011
rect 8017 9959 8073 10011
rect 8125 9959 8181 10011
rect 8233 9959 8289 10011
rect 8341 9959 8397 10011
rect 8449 9959 8505 10011
rect 8557 9959 8613 10011
rect 8665 9959 8721 10011
rect 8773 9959 8829 10011
rect 8881 9959 8937 10011
rect 8989 9959 9045 10011
rect 9097 9959 9153 10011
rect 9205 9959 9261 10011
rect 9313 9959 9369 10011
rect 9421 9959 9477 10011
rect 9529 9959 9553 10011
rect 7725 9523 9553 9959
rect 7725 9471 7749 9523
rect 7801 9471 7857 9523
rect 7909 9471 7965 9523
rect 8017 9471 8073 9523
rect 8125 9471 8181 9523
rect 8233 9471 8289 9523
rect 8341 9471 8397 9523
rect 8449 9471 8505 9523
rect 8557 9471 8613 9523
rect 8665 9471 8721 9523
rect 8773 9471 8829 9523
rect 8881 9471 8937 9523
rect 8989 9471 9045 9523
rect 9097 9471 9153 9523
rect 9205 9471 9261 9523
rect 9313 9471 9369 9523
rect 9421 9471 9477 9523
rect 9529 9471 9553 9523
rect 7725 9035 9553 9471
rect 7725 8983 7749 9035
rect 7801 8983 7857 9035
rect 7909 8983 7965 9035
rect 8017 8983 8073 9035
rect 8125 8983 8181 9035
rect 8233 8983 8289 9035
rect 8341 8983 8397 9035
rect 8449 8983 8505 9035
rect 8557 8983 8613 9035
rect 8665 8983 8721 9035
rect 8773 8983 8829 9035
rect 8881 8983 8937 9035
rect 8989 8983 9045 9035
rect 9097 8983 9153 9035
rect 9205 8983 9261 9035
rect 9313 8983 9369 9035
rect 9421 8983 9477 9035
rect 9529 8983 9553 9035
rect 7725 8547 9553 8983
rect 7725 8495 7749 8547
rect 7801 8495 7857 8547
rect 7909 8495 7965 8547
rect 8017 8495 8073 8547
rect 8125 8495 8181 8547
rect 8233 8495 8289 8547
rect 8341 8495 8397 8547
rect 8449 8495 8505 8547
rect 8557 8495 8613 8547
rect 8665 8495 8721 8547
rect 8773 8495 8829 8547
rect 8881 8495 8937 8547
rect 8989 8495 9045 8547
rect 9097 8495 9153 8547
rect 9205 8495 9261 8547
rect 9313 8495 9369 8547
rect 9421 8495 9477 8547
rect 9529 8495 9553 8547
rect 7725 8059 9553 8495
rect 7725 8007 7749 8059
rect 7801 8007 7857 8059
rect 7909 8007 7965 8059
rect 8017 8007 8073 8059
rect 8125 8007 8181 8059
rect 8233 8007 8289 8059
rect 8341 8007 8397 8059
rect 8449 8007 8505 8059
rect 8557 8007 8613 8059
rect 8665 8007 8721 8059
rect 8773 8007 8829 8059
rect 8881 8007 8937 8059
rect 8989 8007 9045 8059
rect 9097 8007 9153 8059
rect 9205 8007 9261 8059
rect 9313 8007 9369 8059
rect 9421 8007 9477 8059
rect 9529 8007 9553 8059
rect 7725 7571 9553 8007
rect 7725 7519 7749 7571
rect 7801 7519 7857 7571
rect 7909 7519 7965 7571
rect 8017 7519 8073 7571
rect 8125 7519 8181 7571
rect 8233 7519 8289 7571
rect 8341 7519 8397 7571
rect 8449 7519 8505 7571
rect 8557 7519 8613 7571
rect 8665 7519 8721 7571
rect 8773 7519 8829 7571
rect 8881 7519 8937 7571
rect 8989 7519 9045 7571
rect 9097 7519 9153 7571
rect 9205 7519 9261 7571
rect 9313 7519 9369 7571
rect 9421 7519 9477 7571
rect 9529 7519 9553 7571
rect 7725 6885 9553 7519
rect 7725 6833 7749 6885
rect 7801 6833 7857 6885
rect 7909 6833 7965 6885
rect 8017 6833 8073 6885
rect 8125 6833 8181 6885
rect 8233 6833 8289 6885
rect 8341 6833 8397 6885
rect 8449 6833 8505 6885
rect 8557 6833 8613 6885
rect 8665 6833 8721 6885
rect 8773 6833 8829 6885
rect 8881 6833 8937 6885
rect 8989 6833 9045 6885
rect 9097 6833 9153 6885
rect 9205 6833 9261 6885
rect 9313 6833 9369 6885
rect 9421 6833 9477 6885
rect 9529 6833 9553 6885
rect 7725 6777 9553 6833
rect 7725 6725 7749 6777
rect 7801 6725 7857 6777
rect 7909 6725 7965 6777
rect 8017 6725 8073 6777
rect 8125 6725 8181 6777
rect 8233 6725 8289 6777
rect 8341 6725 8397 6777
rect 8449 6725 8505 6777
rect 8557 6725 8613 6777
rect 8665 6725 8721 6777
rect 8773 6725 8829 6777
rect 8881 6725 8937 6777
rect 8989 6725 9045 6777
rect 9097 6725 9153 6777
rect 9205 6725 9261 6777
rect 9313 6725 9369 6777
rect 9421 6725 9477 6777
rect 9529 6725 9553 6777
rect 7725 6091 9553 6725
rect 7725 6039 7749 6091
rect 7801 6039 7857 6091
rect 7909 6039 7965 6091
rect 8017 6039 8073 6091
rect 8125 6039 8181 6091
rect 8233 6039 8289 6091
rect 8341 6039 8397 6091
rect 8449 6039 8505 6091
rect 8557 6039 8613 6091
rect 8665 6039 8721 6091
rect 8773 6039 8829 6091
rect 8881 6039 8937 6091
rect 8989 6039 9045 6091
rect 9097 6039 9153 6091
rect 9205 6039 9261 6091
rect 9313 6039 9369 6091
rect 9421 6039 9477 6091
rect 9529 6039 9553 6091
rect 7725 5603 9553 6039
rect 7725 5551 7749 5603
rect 7801 5551 7857 5603
rect 7909 5551 7965 5603
rect 8017 5551 8073 5603
rect 8125 5551 8181 5603
rect 8233 5551 8289 5603
rect 8341 5551 8397 5603
rect 8449 5551 8505 5603
rect 8557 5551 8613 5603
rect 8665 5551 8721 5603
rect 8773 5551 8829 5603
rect 8881 5551 8937 5603
rect 8989 5551 9045 5603
rect 9097 5551 9153 5603
rect 9205 5551 9261 5603
rect 9313 5551 9369 5603
rect 9421 5551 9477 5603
rect 9529 5551 9553 5603
rect 7725 5115 9553 5551
rect 7725 5063 7749 5115
rect 7801 5063 7857 5115
rect 7909 5063 7965 5115
rect 8017 5063 8073 5115
rect 8125 5063 8181 5115
rect 8233 5063 8289 5115
rect 8341 5063 8397 5115
rect 8449 5063 8505 5115
rect 8557 5063 8613 5115
rect 8665 5063 8721 5115
rect 8773 5063 8829 5115
rect 8881 5063 8937 5115
rect 8989 5063 9045 5115
rect 9097 5063 9153 5115
rect 9205 5063 9261 5115
rect 9313 5063 9369 5115
rect 9421 5063 9477 5115
rect 9529 5063 9553 5115
rect 7725 4627 9553 5063
rect 7725 4575 7749 4627
rect 7801 4575 7857 4627
rect 7909 4575 7965 4627
rect 8017 4575 8073 4627
rect 8125 4575 8181 4627
rect 8233 4575 8289 4627
rect 8341 4575 8397 4627
rect 8449 4575 8505 4627
rect 8557 4575 8613 4627
rect 8665 4575 8721 4627
rect 8773 4575 8829 4627
rect 8881 4575 8937 4627
rect 8989 4575 9045 4627
rect 9097 4575 9153 4627
rect 9205 4575 9261 4627
rect 9313 4575 9369 4627
rect 9421 4575 9477 4627
rect 9529 4575 9553 4627
rect 7725 4139 9553 4575
rect 7725 4087 7749 4139
rect 7801 4087 7857 4139
rect 7909 4087 7965 4139
rect 8017 4087 8073 4139
rect 8125 4087 8181 4139
rect 8233 4087 8289 4139
rect 8341 4087 8397 4139
rect 8449 4087 8505 4139
rect 8557 4087 8613 4139
rect 8665 4087 8721 4139
rect 8773 4087 8829 4139
rect 8881 4087 8937 4139
rect 8989 4087 9045 4139
rect 9097 4087 9153 4139
rect 9205 4087 9261 4139
rect 9313 4087 9369 4139
rect 9421 4087 9477 4139
rect 9529 4087 9553 4139
rect 7725 3651 9553 4087
rect 7725 3599 7749 3651
rect 7801 3599 7857 3651
rect 7909 3599 7965 3651
rect 8017 3599 8073 3651
rect 8125 3599 8181 3651
rect 8233 3599 8289 3651
rect 8341 3599 8397 3651
rect 8449 3599 8505 3651
rect 8557 3599 8613 3651
rect 8665 3599 8721 3651
rect 8773 3599 8829 3651
rect 8881 3599 8937 3651
rect 8989 3599 9045 3651
rect 9097 3599 9153 3651
rect 9205 3599 9261 3651
rect 9313 3599 9369 3651
rect 9421 3599 9477 3651
rect 9529 3599 9553 3651
rect 7725 3163 9553 3599
rect 7725 3111 7749 3163
rect 7801 3111 7857 3163
rect 7909 3111 7965 3163
rect 8017 3111 8073 3163
rect 8125 3111 8181 3163
rect 8233 3111 8289 3163
rect 8341 3111 8397 3163
rect 8449 3111 8505 3163
rect 8557 3111 8613 3163
rect 8665 3111 8721 3163
rect 8773 3111 8829 3163
rect 8881 3111 8937 3163
rect 8989 3111 9045 3163
rect 9097 3111 9153 3163
rect 9205 3111 9261 3163
rect 9313 3111 9369 3163
rect 9421 3111 9477 3163
rect 9529 3111 9553 3163
rect 7725 2675 9553 3111
rect 7725 2623 7749 2675
rect 7801 2623 7857 2675
rect 7909 2623 7965 2675
rect 8017 2623 8073 2675
rect 8125 2623 8181 2675
rect 8233 2623 8289 2675
rect 8341 2623 8397 2675
rect 8449 2623 8505 2675
rect 8557 2623 8613 2675
rect 8665 2623 8721 2675
rect 8773 2623 8829 2675
rect 8881 2623 8937 2675
rect 8989 2623 9045 2675
rect 9097 2623 9153 2675
rect 9205 2623 9261 2675
rect 9313 2623 9369 2675
rect 9421 2623 9477 2675
rect 9529 2623 9553 2675
rect 7725 2187 9553 2623
rect 7725 2135 7749 2187
rect 7801 2135 7857 2187
rect 7909 2135 7965 2187
rect 8017 2135 8073 2187
rect 8125 2135 8181 2187
rect 8233 2135 8289 2187
rect 8341 2135 8397 2187
rect 8449 2135 8505 2187
rect 8557 2135 8613 2187
rect 8665 2135 8721 2187
rect 8773 2135 8829 2187
rect 8881 2135 8937 2187
rect 8989 2135 9045 2187
rect 9097 2135 9153 2187
rect 9205 2135 9261 2187
rect 9313 2135 9369 2187
rect 9421 2135 9477 2187
rect 9529 2135 9553 2187
rect 7725 1699 9553 2135
rect 7725 1647 7749 1699
rect 7801 1647 7857 1699
rect 7909 1647 7965 1699
rect 8017 1647 8073 1699
rect 8125 1647 8181 1699
rect 8233 1647 8289 1699
rect 8341 1647 8397 1699
rect 8449 1647 8505 1699
rect 8557 1647 8613 1699
rect 8665 1647 8721 1699
rect 8773 1647 8829 1699
rect 8881 1647 8937 1699
rect 8989 1647 9045 1699
rect 9097 1647 9153 1699
rect 9205 1647 9261 1699
rect 9313 1647 9369 1699
rect 9421 1647 9477 1699
rect 9529 1647 9553 1699
rect 7725 961 9553 1647
rect 7725 909 7749 961
rect 7801 909 7857 961
rect 7909 909 7965 961
rect 8017 909 8073 961
rect 8125 909 8181 961
rect 8233 909 8289 961
rect 8341 909 8397 961
rect 8449 909 8505 961
rect 8557 909 8613 961
rect 8665 909 8721 961
rect 8773 909 8829 961
rect 8881 909 8937 961
rect 8989 909 9045 961
rect 9097 909 9153 961
rect 9205 909 9261 961
rect 9313 909 9369 961
rect 9421 909 9477 961
rect 9529 909 9553 961
rect 7725 853 9553 909
rect 7725 801 7749 853
rect 7801 801 7857 853
rect 7909 801 7965 853
rect 8017 801 8073 853
rect 8125 801 8181 853
rect 8233 801 8289 853
rect 8341 801 8397 853
rect 8449 801 8505 853
rect 8557 801 8613 853
rect 8665 801 8721 853
rect 8773 801 8829 853
rect 8881 801 8937 853
rect 8989 801 9045 853
rect 9097 801 9153 853
rect 9205 801 9261 853
rect 9313 801 9369 853
rect 9421 801 9477 853
rect 9529 801 9553 853
rect 7725 745 9553 801
rect 7725 693 7749 745
rect 7801 693 7857 745
rect 7909 693 7965 745
rect 8017 693 8073 745
rect 8125 693 8181 745
rect 8233 693 8289 745
rect 8341 693 8397 745
rect 8449 693 8505 745
rect 8557 693 8613 745
rect 8665 693 8721 745
rect 8773 693 8829 745
rect 8881 693 8937 745
rect 8989 693 9045 745
rect 9097 693 9153 745
rect 9205 693 9261 745
rect 9313 693 9369 745
rect 9421 693 9477 745
rect 9529 693 9553 745
rect 7725 43 9553 693
rect 9653 25261 11481 25617
rect 9653 25209 9677 25261
rect 9729 25209 9785 25261
rect 9837 25209 9893 25261
rect 9945 25209 10001 25261
rect 10053 25209 10109 25261
rect 10161 25209 10217 25261
rect 10269 25209 10325 25261
rect 10377 25209 10433 25261
rect 10485 25209 10541 25261
rect 10593 25209 10649 25261
rect 10701 25209 10757 25261
rect 10809 25209 10865 25261
rect 10917 25209 10973 25261
rect 11025 25209 11081 25261
rect 11133 25209 11189 25261
rect 11241 25209 11297 25261
rect 11349 25209 11405 25261
rect 11457 25209 11481 25261
rect 9653 25153 11481 25209
rect 9653 25101 9677 25153
rect 9729 25101 9785 25153
rect 9837 25101 9893 25153
rect 9945 25101 10001 25153
rect 10053 25101 10109 25153
rect 10161 25101 10217 25153
rect 10269 25101 10325 25153
rect 10377 25101 10433 25153
rect 10485 25101 10541 25153
rect 10593 25101 10649 25153
rect 10701 25101 10757 25153
rect 10809 25101 10865 25153
rect 10917 25101 10973 25153
rect 11025 25101 11081 25153
rect 11133 25101 11189 25153
rect 11241 25101 11297 25153
rect 11349 25101 11405 25153
rect 11457 25101 11481 25153
rect 9653 25045 11481 25101
rect 9653 24993 9677 25045
rect 9729 24993 9785 25045
rect 9837 24993 9893 25045
rect 9945 24993 10001 25045
rect 10053 24993 10109 25045
rect 10161 24993 10217 25045
rect 10269 24993 10325 25045
rect 10377 24993 10433 25045
rect 10485 24993 10541 25045
rect 10593 24993 10649 25045
rect 10701 24993 10757 25045
rect 10809 24993 10865 25045
rect 10917 24993 10973 25045
rect 11025 24993 11081 25045
rect 11133 24993 11189 25045
rect 11241 24993 11297 25045
rect 11349 24993 11405 25045
rect 11457 24993 11481 25045
rect 9653 23951 11481 24993
rect 9653 23899 9677 23951
rect 9729 23899 9785 23951
rect 9837 23899 9893 23951
rect 9945 23899 10001 23951
rect 10053 23899 10109 23951
rect 10161 23899 10217 23951
rect 10269 23899 10325 23951
rect 10377 23899 10433 23951
rect 10485 23899 10541 23951
rect 10593 23899 10649 23951
rect 10701 23899 10757 23951
rect 10809 23899 10865 23951
rect 10917 23899 10973 23951
rect 11025 23899 11081 23951
rect 11133 23899 11189 23951
rect 11241 23899 11297 23951
rect 11349 23899 11405 23951
rect 11457 23899 11481 23951
rect 9653 23463 11481 23899
rect 9653 23411 9677 23463
rect 9729 23411 9785 23463
rect 9837 23411 9893 23463
rect 9945 23411 10001 23463
rect 10053 23411 10109 23463
rect 10161 23411 10217 23463
rect 10269 23411 10325 23463
rect 10377 23411 10433 23463
rect 10485 23411 10541 23463
rect 10593 23411 10649 23463
rect 10701 23411 10757 23463
rect 10809 23411 10865 23463
rect 10917 23411 10973 23463
rect 11025 23411 11081 23463
rect 11133 23411 11189 23463
rect 11241 23411 11297 23463
rect 11349 23411 11405 23463
rect 11457 23411 11481 23463
rect 9653 22975 11481 23411
rect 9653 22923 9677 22975
rect 9729 22923 9785 22975
rect 9837 22923 9893 22975
rect 9945 22923 10001 22975
rect 10053 22923 10109 22975
rect 10161 22923 10217 22975
rect 10269 22923 10325 22975
rect 10377 22923 10433 22975
rect 10485 22923 10541 22975
rect 10593 22923 10649 22975
rect 10701 22923 10757 22975
rect 10809 22923 10865 22975
rect 10917 22923 10973 22975
rect 11025 22923 11081 22975
rect 11133 22923 11189 22975
rect 11241 22923 11297 22975
rect 11349 22923 11405 22975
rect 11457 22923 11481 22975
rect 9653 22487 11481 22923
rect 9653 22435 9677 22487
rect 9729 22435 9785 22487
rect 9837 22435 9893 22487
rect 9945 22435 10001 22487
rect 10053 22435 10109 22487
rect 10161 22435 10217 22487
rect 10269 22435 10325 22487
rect 10377 22435 10433 22487
rect 10485 22435 10541 22487
rect 10593 22435 10649 22487
rect 10701 22435 10757 22487
rect 10809 22435 10865 22487
rect 10917 22435 10973 22487
rect 11025 22435 11081 22487
rect 11133 22435 11189 22487
rect 11241 22435 11297 22487
rect 11349 22435 11405 22487
rect 11457 22435 11481 22487
rect 9653 21999 11481 22435
rect 9653 21947 9677 21999
rect 9729 21947 9785 21999
rect 9837 21947 9893 21999
rect 9945 21947 10001 21999
rect 10053 21947 10109 21999
rect 10161 21947 10217 21999
rect 10269 21947 10325 21999
rect 10377 21947 10433 21999
rect 10485 21947 10541 21999
rect 10593 21947 10649 21999
rect 10701 21947 10757 21999
rect 10809 21947 10865 21999
rect 10917 21947 10973 21999
rect 11025 21947 11081 21999
rect 11133 21947 11189 21999
rect 11241 21947 11297 21999
rect 11349 21947 11405 21999
rect 11457 21947 11481 21999
rect 9653 21511 11481 21947
rect 9653 21459 9677 21511
rect 9729 21459 9785 21511
rect 9837 21459 9893 21511
rect 9945 21459 10001 21511
rect 10053 21459 10109 21511
rect 10161 21459 10217 21511
rect 10269 21459 10325 21511
rect 10377 21459 10433 21511
rect 10485 21459 10541 21511
rect 10593 21459 10649 21511
rect 10701 21459 10757 21511
rect 10809 21459 10865 21511
rect 10917 21459 10973 21511
rect 11025 21459 11081 21511
rect 11133 21459 11189 21511
rect 11241 21459 11297 21511
rect 11349 21459 11405 21511
rect 11457 21459 11481 21511
rect 9653 21023 11481 21459
rect 9653 20971 9677 21023
rect 9729 20971 9785 21023
rect 9837 20971 9893 21023
rect 9945 20971 10001 21023
rect 10053 20971 10109 21023
rect 10161 20971 10217 21023
rect 10269 20971 10325 21023
rect 10377 20971 10433 21023
rect 10485 20971 10541 21023
rect 10593 20971 10649 21023
rect 10701 20971 10757 21023
rect 10809 20971 10865 21023
rect 10917 20971 10973 21023
rect 11025 20971 11081 21023
rect 11133 20971 11189 21023
rect 11241 20971 11297 21023
rect 11349 20971 11405 21023
rect 11457 20971 11481 21023
rect 9653 20535 11481 20971
rect 9653 20483 9677 20535
rect 9729 20483 9785 20535
rect 9837 20483 9893 20535
rect 9945 20483 10001 20535
rect 10053 20483 10109 20535
rect 10161 20483 10217 20535
rect 10269 20483 10325 20535
rect 10377 20483 10433 20535
rect 10485 20483 10541 20535
rect 10593 20483 10649 20535
rect 10701 20483 10757 20535
rect 10809 20483 10865 20535
rect 10917 20483 10973 20535
rect 11025 20483 11081 20535
rect 11133 20483 11189 20535
rect 11241 20483 11297 20535
rect 11349 20483 11405 20535
rect 11457 20483 11481 20535
rect 9653 20047 11481 20483
rect 9653 19995 9677 20047
rect 9729 19995 9785 20047
rect 9837 19995 9893 20047
rect 9945 19995 10001 20047
rect 10053 19995 10109 20047
rect 10161 19995 10217 20047
rect 10269 19995 10325 20047
rect 10377 19995 10433 20047
rect 10485 19995 10541 20047
rect 10593 19995 10649 20047
rect 10701 19995 10757 20047
rect 10809 19995 10865 20047
rect 10917 19995 10973 20047
rect 11025 19995 11081 20047
rect 11133 19995 11189 20047
rect 11241 19995 11297 20047
rect 11349 19995 11405 20047
rect 11457 19995 11481 20047
rect 9653 19559 11481 19995
rect 9653 19507 9677 19559
rect 9729 19507 9785 19559
rect 9837 19507 9893 19559
rect 9945 19507 10001 19559
rect 10053 19507 10109 19559
rect 10161 19507 10217 19559
rect 10269 19507 10325 19559
rect 10377 19507 10433 19559
rect 10485 19507 10541 19559
rect 10593 19507 10649 19559
rect 10701 19507 10757 19559
rect 10809 19507 10865 19559
rect 10917 19507 10973 19559
rect 11025 19507 11081 19559
rect 11133 19507 11189 19559
rect 11241 19507 11297 19559
rect 11349 19507 11405 19559
rect 11457 19507 11481 19559
rect 9653 19071 11481 19507
rect 9653 19019 9677 19071
rect 9729 19019 9785 19071
rect 9837 19019 9893 19071
rect 9945 19019 10001 19071
rect 10053 19019 10109 19071
rect 10161 19019 10217 19071
rect 10269 19019 10325 19071
rect 10377 19019 10433 19071
rect 10485 19019 10541 19071
rect 10593 19019 10649 19071
rect 10701 19019 10757 19071
rect 10809 19019 10865 19071
rect 10917 19019 10973 19071
rect 11025 19019 11081 19071
rect 11133 19019 11189 19071
rect 11241 19019 11297 19071
rect 11349 19019 11405 19071
rect 11457 19019 11481 19071
rect 9653 18079 11481 19019
rect 9653 18027 9677 18079
rect 9729 18027 9785 18079
rect 9837 18027 9893 18079
rect 9945 18027 10001 18079
rect 10053 18027 10109 18079
rect 10161 18027 10217 18079
rect 10269 18027 10325 18079
rect 10377 18027 10433 18079
rect 10485 18027 10541 18079
rect 10593 18027 10649 18079
rect 10701 18027 10757 18079
rect 10809 18027 10865 18079
rect 10917 18027 10973 18079
rect 11025 18027 11081 18079
rect 11133 18027 11189 18079
rect 11241 18027 11297 18079
rect 11349 18027 11405 18079
rect 11457 18027 11481 18079
rect 9653 17591 11481 18027
rect 9653 17539 9677 17591
rect 9729 17539 9785 17591
rect 9837 17539 9893 17591
rect 9945 17539 10001 17591
rect 10053 17539 10109 17591
rect 10161 17539 10217 17591
rect 10269 17539 10325 17591
rect 10377 17539 10433 17591
rect 10485 17539 10541 17591
rect 10593 17539 10649 17591
rect 10701 17539 10757 17591
rect 10809 17539 10865 17591
rect 10917 17539 10973 17591
rect 11025 17539 11081 17591
rect 11133 17539 11189 17591
rect 11241 17539 11297 17591
rect 11349 17539 11405 17591
rect 11457 17539 11481 17591
rect 9653 17103 11481 17539
rect 9653 17051 9677 17103
rect 9729 17051 9785 17103
rect 9837 17051 9893 17103
rect 9945 17051 10001 17103
rect 10053 17051 10109 17103
rect 10161 17051 10217 17103
rect 10269 17051 10325 17103
rect 10377 17051 10433 17103
rect 10485 17051 10541 17103
rect 10593 17051 10649 17103
rect 10701 17051 10757 17103
rect 10809 17051 10865 17103
rect 10917 17051 10973 17103
rect 11025 17051 11081 17103
rect 11133 17051 11189 17103
rect 11241 17051 11297 17103
rect 11349 17051 11405 17103
rect 11457 17051 11481 17103
rect 9653 16615 11481 17051
rect 9653 16563 9677 16615
rect 9729 16563 9785 16615
rect 9837 16563 9893 16615
rect 9945 16563 10001 16615
rect 10053 16563 10109 16615
rect 10161 16563 10217 16615
rect 10269 16563 10325 16615
rect 10377 16563 10433 16615
rect 10485 16563 10541 16615
rect 10593 16563 10649 16615
rect 10701 16563 10757 16615
rect 10809 16563 10865 16615
rect 10917 16563 10973 16615
rect 11025 16563 11081 16615
rect 11133 16563 11189 16615
rect 11241 16563 11297 16615
rect 11349 16563 11405 16615
rect 11457 16563 11481 16615
rect 9653 16127 11481 16563
rect 9653 16075 9677 16127
rect 9729 16075 9785 16127
rect 9837 16075 9893 16127
rect 9945 16075 10001 16127
rect 10053 16075 10109 16127
rect 10161 16075 10217 16127
rect 10269 16075 10325 16127
rect 10377 16075 10433 16127
rect 10485 16075 10541 16127
rect 10593 16075 10649 16127
rect 10701 16075 10757 16127
rect 10809 16075 10865 16127
rect 10917 16075 10973 16127
rect 11025 16075 11081 16127
rect 11133 16075 11189 16127
rect 11241 16075 11297 16127
rect 11349 16075 11405 16127
rect 11457 16075 11481 16127
rect 9653 15639 11481 16075
rect 9653 15587 9677 15639
rect 9729 15587 9785 15639
rect 9837 15587 9893 15639
rect 9945 15587 10001 15639
rect 10053 15587 10109 15639
rect 10161 15587 10217 15639
rect 10269 15587 10325 15639
rect 10377 15587 10433 15639
rect 10485 15587 10541 15639
rect 10593 15587 10649 15639
rect 10701 15587 10757 15639
rect 10809 15587 10865 15639
rect 10917 15587 10973 15639
rect 11025 15587 11081 15639
rect 11133 15587 11189 15639
rect 11241 15587 11297 15639
rect 11349 15587 11405 15639
rect 11457 15587 11481 15639
rect 9653 15151 11481 15587
rect 9653 15099 9677 15151
rect 9729 15099 9785 15151
rect 9837 15099 9893 15151
rect 9945 15099 10001 15151
rect 10053 15099 10109 15151
rect 10161 15099 10217 15151
rect 10269 15099 10325 15151
rect 10377 15099 10433 15151
rect 10485 15099 10541 15151
rect 10593 15099 10649 15151
rect 10701 15099 10757 15151
rect 10809 15099 10865 15151
rect 10917 15099 10973 15151
rect 11025 15099 11081 15151
rect 11133 15099 11189 15151
rect 11241 15099 11297 15151
rect 11349 15099 11405 15151
rect 11457 15099 11481 15151
rect 9653 14663 11481 15099
rect 9653 14611 9677 14663
rect 9729 14611 9785 14663
rect 9837 14611 9893 14663
rect 9945 14611 10001 14663
rect 10053 14611 10109 14663
rect 10161 14611 10217 14663
rect 10269 14611 10325 14663
rect 10377 14611 10433 14663
rect 10485 14611 10541 14663
rect 10593 14611 10649 14663
rect 10701 14611 10757 14663
rect 10809 14611 10865 14663
rect 10917 14611 10973 14663
rect 11025 14611 11081 14663
rect 11133 14611 11189 14663
rect 11241 14611 11297 14663
rect 11349 14611 11405 14663
rect 11457 14611 11481 14663
rect 9653 14175 11481 14611
rect 9653 14123 9677 14175
rect 9729 14123 9785 14175
rect 9837 14123 9893 14175
rect 9945 14123 10001 14175
rect 10053 14123 10109 14175
rect 10161 14123 10217 14175
rect 10269 14123 10325 14175
rect 10377 14123 10433 14175
rect 10485 14123 10541 14175
rect 10593 14123 10649 14175
rect 10701 14123 10757 14175
rect 10809 14123 10865 14175
rect 10917 14123 10973 14175
rect 11025 14123 11081 14175
rect 11133 14123 11189 14175
rect 11241 14123 11297 14175
rect 11349 14123 11405 14175
rect 11457 14123 11481 14175
rect 9653 13687 11481 14123
rect 9653 13635 9677 13687
rect 9729 13635 9785 13687
rect 9837 13635 9893 13687
rect 9945 13635 10001 13687
rect 10053 13635 10109 13687
rect 10161 13635 10217 13687
rect 10269 13635 10325 13687
rect 10377 13635 10433 13687
rect 10485 13635 10541 13687
rect 10593 13635 10649 13687
rect 10701 13635 10757 13687
rect 10809 13635 10865 13687
rect 10917 13635 10973 13687
rect 11025 13635 11081 13687
rect 11133 13635 11189 13687
rect 11241 13635 11297 13687
rect 11349 13635 11405 13687
rect 11457 13635 11481 13687
rect 9653 13199 11481 13635
rect 9653 13147 9677 13199
rect 9729 13147 9785 13199
rect 9837 13147 9893 13199
rect 9945 13147 10001 13199
rect 10053 13147 10109 13199
rect 10161 13147 10217 13199
rect 10269 13147 10325 13199
rect 10377 13147 10433 13199
rect 10485 13147 10541 13199
rect 10593 13147 10649 13199
rect 10701 13147 10757 13199
rect 10809 13147 10865 13199
rect 10917 13147 10973 13199
rect 11025 13147 11081 13199
rect 11133 13147 11189 13199
rect 11241 13147 11297 13199
rect 11349 13147 11405 13199
rect 11457 13147 11481 13199
rect 9653 12207 11481 13147
rect 9653 12155 9677 12207
rect 9729 12155 9785 12207
rect 9837 12155 9893 12207
rect 9945 12155 10001 12207
rect 10053 12155 10109 12207
rect 10161 12155 10217 12207
rect 10269 12155 10325 12207
rect 10377 12155 10433 12207
rect 10485 12155 10541 12207
rect 10593 12155 10649 12207
rect 10701 12155 10757 12207
rect 10809 12155 10865 12207
rect 10917 12155 10973 12207
rect 11025 12155 11081 12207
rect 11133 12155 11189 12207
rect 11241 12155 11297 12207
rect 11349 12155 11405 12207
rect 11457 12155 11481 12207
rect 9653 11719 11481 12155
rect 9653 11667 9677 11719
rect 9729 11667 9785 11719
rect 9837 11667 9893 11719
rect 9945 11667 10001 11719
rect 10053 11667 10109 11719
rect 10161 11667 10217 11719
rect 10269 11667 10325 11719
rect 10377 11667 10433 11719
rect 10485 11667 10541 11719
rect 10593 11667 10649 11719
rect 10701 11667 10757 11719
rect 10809 11667 10865 11719
rect 10917 11667 10973 11719
rect 11025 11667 11081 11719
rect 11133 11667 11189 11719
rect 11241 11667 11297 11719
rect 11349 11667 11405 11719
rect 11457 11667 11481 11719
rect 9653 11231 11481 11667
rect 9653 11179 9677 11231
rect 9729 11179 9785 11231
rect 9837 11179 9893 11231
rect 9945 11179 10001 11231
rect 10053 11179 10109 11231
rect 10161 11179 10217 11231
rect 10269 11179 10325 11231
rect 10377 11179 10433 11231
rect 10485 11179 10541 11231
rect 10593 11179 10649 11231
rect 10701 11179 10757 11231
rect 10809 11179 10865 11231
rect 10917 11179 10973 11231
rect 11025 11179 11081 11231
rect 11133 11179 11189 11231
rect 11241 11179 11297 11231
rect 11349 11179 11405 11231
rect 11457 11179 11481 11231
rect 9653 10743 11481 11179
rect 9653 10691 9677 10743
rect 9729 10691 9785 10743
rect 9837 10691 9893 10743
rect 9945 10691 10001 10743
rect 10053 10691 10109 10743
rect 10161 10691 10217 10743
rect 10269 10691 10325 10743
rect 10377 10691 10433 10743
rect 10485 10691 10541 10743
rect 10593 10691 10649 10743
rect 10701 10691 10757 10743
rect 10809 10691 10865 10743
rect 10917 10691 10973 10743
rect 11025 10691 11081 10743
rect 11133 10691 11189 10743
rect 11241 10691 11297 10743
rect 11349 10691 11405 10743
rect 11457 10691 11481 10743
rect 9653 10255 11481 10691
rect 9653 10203 9677 10255
rect 9729 10203 9785 10255
rect 9837 10203 9893 10255
rect 9945 10203 10001 10255
rect 10053 10203 10109 10255
rect 10161 10203 10217 10255
rect 10269 10203 10325 10255
rect 10377 10203 10433 10255
rect 10485 10203 10541 10255
rect 10593 10203 10649 10255
rect 10701 10203 10757 10255
rect 10809 10203 10865 10255
rect 10917 10203 10973 10255
rect 11025 10203 11081 10255
rect 11133 10203 11189 10255
rect 11241 10203 11297 10255
rect 11349 10203 11405 10255
rect 11457 10203 11481 10255
rect 9653 9767 11481 10203
rect 9653 9715 9677 9767
rect 9729 9715 9785 9767
rect 9837 9715 9893 9767
rect 9945 9715 10001 9767
rect 10053 9715 10109 9767
rect 10161 9715 10217 9767
rect 10269 9715 10325 9767
rect 10377 9715 10433 9767
rect 10485 9715 10541 9767
rect 10593 9715 10649 9767
rect 10701 9715 10757 9767
rect 10809 9715 10865 9767
rect 10917 9715 10973 9767
rect 11025 9715 11081 9767
rect 11133 9715 11189 9767
rect 11241 9715 11297 9767
rect 11349 9715 11405 9767
rect 11457 9715 11481 9767
rect 9653 9279 11481 9715
rect 9653 9227 9677 9279
rect 9729 9227 9785 9279
rect 9837 9227 9893 9279
rect 9945 9227 10001 9279
rect 10053 9227 10109 9279
rect 10161 9227 10217 9279
rect 10269 9227 10325 9279
rect 10377 9227 10433 9279
rect 10485 9227 10541 9279
rect 10593 9227 10649 9279
rect 10701 9227 10757 9279
rect 10809 9227 10865 9279
rect 10917 9227 10973 9279
rect 11025 9227 11081 9279
rect 11133 9227 11189 9279
rect 11241 9227 11297 9279
rect 11349 9227 11405 9279
rect 11457 9227 11481 9279
rect 9653 8791 11481 9227
rect 9653 8739 9677 8791
rect 9729 8739 9785 8791
rect 9837 8739 9893 8791
rect 9945 8739 10001 8791
rect 10053 8739 10109 8791
rect 10161 8739 10217 8791
rect 10269 8739 10325 8791
rect 10377 8739 10433 8791
rect 10485 8739 10541 8791
rect 10593 8739 10649 8791
rect 10701 8739 10757 8791
rect 10809 8739 10865 8791
rect 10917 8739 10973 8791
rect 11025 8739 11081 8791
rect 11133 8739 11189 8791
rect 11241 8739 11297 8791
rect 11349 8739 11405 8791
rect 11457 8739 11481 8791
rect 9653 8303 11481 8739
rect 9653 8251 9677 8303
rect 9729 8251 9785 8303
rect 9837 8251 9893 8303
rect 9945 8251 10001 8303
rect 10053 8251 10109 8303
rect 10161 8251 10217 8303
rect 10269 8251 10325 8303
rect 10377 8251 10433 8303
rect 10485 8251 10541 8303
rect 10593 8251 10649 8303
rect 10701 8251 10757 8303
rect 10809 8251 10865 8303
rect 10917 8251 10973 8303
rect 11025 8251 11081 8303
rect 11133 8251 11189 8303
rect 11241 8251 11297 8303
rect 11349 8251 11405 8303
rect 11457 8251 11481 8303
rect 9653 7815 11481 8251
rect 9653 7763 9677 7815
rect 9729 7763 9785 7815
rect 9837 7763 9893 7815
rect 9945 7763 10001 7815
rect 10053 7763 10109 7815
rect 10161 7763 10217 7815
rect 10269 7763 10325 7815
rect 10377 7763 10433 7815
rect 10485 7763 10541 7815
rect 10593 7763 10649 7815
rect 10701 7763 10757 7815
rect 10809 7763 10865 7815
rect 10917 7763 10973 7815
rect 11025 7763 11081 7815
rect 11133 7763 11189 7815
rect 11241 7763 11297 7815
rect 11349 7763 11405 7815
rect 11457 7763 11481 7815
rect 9653 7327 11481 7763
rect 9653 7275 9677 7327
rect 9729 7275 9785 7327
rect 9837 7275 9893 7327
rect 9945 7275 10001 7327
rect 10053 7275 10109 7327
rect 10161 7275 10217 7327
rect 10269 7275 10325 7327
rect 10377 7275 10433 7327
rect 10485 7275 10541 7327
rect 10593 7275 10649 7327
rect 10701 7275 10757 7327
rect 10809 7275 10865 7327
rect 10917 7275 10973 7327
rect 11025 7275 11081 7327
rect 11133 7275 11189 7327
rect 11241 7275 11297 7327
rect 11349 7275 11405 7327
rect 11457 7275 11481 7327
rect 9653 6335 11481 7275
rect 9653 6283 9677 6335
rect 9729 6283 9785 6335
rect 9837 6283 9893 6335
rect 9945 6283 10001 6335
rect 10053 6283 10109 6335
rect 10161 6283 10217 6335
rect 10269 6283 10325 6335
rect 10377 6283 10433 6335
rect 10485 6283 10541 6335
rect 10593 6283 10649 6335
rect 10701 6283 10757 6335
rect 10809 6283 10865 6335
rect 10917 6283 10973 6335
rect 11025 6283 11081 6335
rect 11133 6283 11189 6335
rect 11241 6283 11297 6335
rect 11349 6283 11405 6335
rect 11457 6283 11481 6335
rect 9653 5847 11481 6283
rect 9653 5795 9677 5847
rect 9729 5795 9785 5847
rect 9837 5795 9893 5847
rect 9945 5795 10001 5847
rect 10053 5795 10109 5847
rect 10161 5795 10217 5847
rect 10269 5795 10325 5847
rect 10377 5795 10433 5847
rect 10485 5795 10541 5847
rect 10593 5795 10649 5847
rect 10701 5795 10757 5847
rect 10809 5795 10865 5847
rect 10917 5795 10973 5847
rect 11025 5795 11081 5847
rect 11133 5795 11189 5847
rect 11241 5795 11297 5847
rect 11349 5795 11405 5847
rect 11457 5795 11481 5847
rect 9653 5359 11481 5795
rect 9653 5307 9677 5359
rect 9729 5307 9785 5359
rect 9837 5307 9893 5359
rect 9945 5307 10001 5359
rect 10053 5307 10109 5359
rect 10161 5307 10217 5359
rect 10269 5307 10325 5359
rect 10377 5307 10433 5359
rect 10485 5307 10541 5359
rect 10593 5307 10649 5359
rect 10701 5307 10757 5359
rect 10809 5307 10865 5359
rect 10917 5307 10973 5359
rect 11025 5307 11081 5359
rect 11133 5307 11189 5359
rect 11241 5307 11297 5359
rect 11349 5307 11405 5359
rect 11457 5307 11481 5359
rect 9653 4871 11481 5307
rect 9653 4819 9677 4871
rect 9729 4819 9785 4871
rect 9837 4819 9893 4871
rect 9945 4819 10001 4871
rect 10053 4819 10109 4871
rect 10161 4819 10217 4871
rect 10269 4819 10325 4871
rect 10377 4819 10433 4871
rect 10485 4819 10541 4871
rect 10593 4819 10649 4871
rect 10701 4819 10757 4871
rect 10809 4819 10865 4871
rect 10917 4819 10973 4871
rect 11025 4819 11081 4871
rect 11133 4819 11189 4871
rect 11241 4819 11297 4871
rect 11349 4819 11405 4871
rect 11457 4819 11481 4871
rect 9653 4383 11481 4819
rect 9653 4331 9677 4383
rect 9729 4331 9785 4383
rect 9837 4331 9893 4383
rect 9945 4331 10001 4383
rect 10053 4331 10109 4383
rect 10161 4331 10217 4383
rect 10269 4331 10325 4383
rect 10377 4331 10433 4383
rect 10485 4331 10541 4383
rect 10593 4331 10649 4383
rect 10701 4331 10757 4383
rect 10809 4331 10865 4383
rect 10917 4331 10973 4383
rect 11025 4331 11081 4383
rect 11133 4331 11189 4383
rect 11241 4331 11297 4383
rect 11349 4331 11405 4383
rect 11457 4331 11481 4383
rect 9653 3895 11481 4331
rect 9653 3843 9677 3895
rect 9729 3843 9785 3895
rect 9837 3843 9893 3895
rect 9945 3843 10001 3895
rect 10053 3843 10109 3895
rect 10161 3843 10217 3895
rect 10269 3843 10325 3895
rect 10377 3843 10433 3895
rect 10485 3843 10541 3895
rect 10593 3843 10649 3895
rect 10701 3843 10757 3895
rect 10809 3843 10865 3895
rect 10917 3843 10973 3895
rect 11025 3843 11081 3895
rect 11133 3843 11189 3895
rect 11241 3843 11297 3895
rect 11349 3843 11405 3895
rect 11457 3843 11481 3895
rect 9653 3407 11481 3843
rect 9653 3355 9677 3407
rect 9729 3355 9785 3407
rect 9837 3355 9893 3407
rect 9945 3355 10001 3407
rect 10053 3355 10109 3407
rect 10161 3355 10217 3407
rect 10269 3355 10325 3407
rect 10377 3355 10433 3407
rect 10485 3355 10541 3407
rect 10593 3355 10649 3407
rect 10701 3355 10757 3407
rect 10809 3355 10865 3407
rect 10917 3355 10973 3407
rect 11025 3355 11081 3407
rect 11133 3355 11189 3407
rect 11241 3355 11297 3407
rect 11349 3355 11405 3407
rect 11457 3355 11481 3407
rect 9653 2919 11481 3355
rect 9653 2867 9677 2919
rect 9729 2867 9785 2919
rect 9837 2867 9893 2919
rect 9945 2867 10001 2919
rect 10053 2867 10109 2919
rect 10161 2867 10217 2919
rect 10269 2867 10325 2919
rect 10377 2867 10433 2919
rect 10485 2867 10541 2919
rect 10593 2867 10649 2919
rect 10701 2867 10757 2919
rect 10809 2867 10865 2919
rect 10917 2867 10973 2919
rect 11025 2867 11081 2919
rect 11133 2867 11189 2919
rect 11241 2867 11297 2919
rect 11349 2867 11405 2919
rect 11457 2867 11481 2919
rect 9653 2431 11481 2867
rect 9653 2379 9677 2431
rect 9729 2379 9785 2431
rect 9837 2379 9893 2431
rect 9945 2379 10001 2431
rect 10053 2379 10109 2431
rect 10161 2379 10217 2431
rect 10269 2379 10325 2431
rect 10377 2379 10433 2431
rect 10485 2379 10541 2431
rect 10593 2379 10649 2431
rect 10701 2379 10757 2431
rect 10809 2379 10865 2431
rect 10917 2379 10973 2431
rect 11025 2379 11081 2431
rect 11133 2379 11189 2431
rect 11241 2379 11297 2431
rect 11349 2379 11405 2431
rect 11457 2379 11481 2431
rect 9653 1943 11481 2379
rect 9653 1891 9677 1943
rect 9729 1891 9785 1943
rect 9837 1891 9893 1943
rect 9945 1891 10001 1943
rect 10053 1891 10109 1943
rect 10161 1891 10217 1943
rect 10269 1891 10325 1943
rect 10377 1891 10433 1943
rect 10485 1891 10541 1943
rect 10593 1891 10649 1943
rect 10701 1891 10757 1943
rect 10809 1891 10865 1943
rect 10917 1891 10973 1943
rect 11025 1891 11081 1943
rect 11133 1891 11189 1943
rect 11241 1891 11297 1943
rect 11349 1891 11405 1943
rect 11457 1891 11481 1943
rect 9653 1455 11481 1891
rect 11549 23887 11749 25617
rect 11549 23835 11569 23887
rect 11621 23835 11677 23887
rect 11729 23835 11749 23887
rect 11549 23779 11749 23835
rect 11549 23727 11569 23779
rect 11621 23727 11677 23779
rect 11729 23727 11749 23779
rect 11549 23671 11749 23727
rect 11549 23619 11569 23671
rect 11621 23619 11677 23671
rect 11729 23619 11749 23671
rect 11549 23563 11749 23619
rect 11549 23511 11569 23563
rect 11621 23511 11677 23563
rect 11729 23511 11749 23563
rect 11549 23455 11749 23511
rect 11549 23403 11569 23455
rect 11621 23403 11677 23455
rect 11729 23403 11749 23455
rect 11549 23347 11749 23403
rect 11549 23295 11569 23347
rect 11621 23295 11677 23347
rect 11729 23295 11749 23347
rect 11549 23239 11749 23295
rect 11549 23187 11569 23239
rect 11621 23187 11677 23239
rect 11729 23187 11749 23239
rect 11549 23131 11749 23187
rect 11549 23079 11569 23131
rect 11621 23079 11677 23131
rect 11729 23079 11749 23131
rect 11549 23023 11749 23079
rect 11549 22971 11569 23023
rect 11621 22971 11677 23023
rect 11729 22971 11749 23023
rect 11549 22915 11749 22971
rect 11549 22863 11569 22915
rect 11621 22863 11677 22915
rect 11729 22863 11749 22915
rect 11549 22807 11749 22863
rect 11549 22755 11569 22807
rect 11621 22755 11677 22807
rect 11729 22755 11749 22807
rect 11549 22699 11749 22755
rect 11549 22647 11569 22699
rect 11621 22647 11677 22699
rect 11729 22647 11749 22699
rect 11549 22591 11749 22647
rect 11549 22539 11569 22591
rect 11621 22539 11677 22591
rect 11729 22539 11749 22591
rect 11549 22483 11749 22539
rect 11549 22431 11569 22483
rect 11621 22431 11677 22483
rect 11729 22431 11749 22483
rect 11549 22375 11749 22431
rect 11549 22323 11569 22375
rect 11621 22323 11677 22375
rect 11729 22323 11749 22375
rect 11549 22267 11749 22323
rect 11549 22215 11569 22267
rect 11621 22215 11677 22267
rect 11729 22215 11749 22267
rect 11549 22159 11749 22215
rect 11549 22107 11569 22159
rect 11621 22107 11677 22159
rect 11729 22107 11749 22159
rect 11549 22051 11749 22107
rect 11549 21999 11569 22051
rect 11621 21999 11677 22051
rect 11729 21999 11749 22051
rect 11549 21943 11749 21999
rect 11549 21891 11569 21943
rect 11621 21891 11677 21943
rect 11729 21891 11749 21943
rect 11549 21835 11749 21891
rect 11549 21783 11569 21835
rect 11621 21783 11677 21835
rect 11729 21783 11749 21835
rect 11549 21727 11749 21783
rect 11549 21675 11569 21727
rect 11621 21675 11677 21727
rect 11729 21675 11749 21727
rect 11549 21619 11749 21675
rect 11549 21567 11569 21619
rect 11621 21567 11677 21619
rect 11729 21567 11749 21619
rect 11549 21511 11749 21567
rect 11549 21459 11569 21511
rect 11621 21459 11677 21511
rect 11729 21459 11749 21511
rect 11549 21403 11749 21459
rect 11549 21351 11569 21403
rect 11621 21351 11677 21403
rect 11729 21351 11749 21403
rect 11549 21295 11749 21351
rect 11549 21243 11569 21295
rect 11621 21243 11677 21295
rect 11729 21243 11749 21295
rect 11549 21187 11749 21243
rect 11549 21135 11569 21187
rect 11621 21135 11677 21187
rect 11729 21135 11749 21187
rect 11549 21079 11749 21135
rect 11549 21027 11569 21079
rect 11621 21027 11677 21079
rect 11729 21027 11749 21079
rect 11549 20971 11749 21027
rect 11549 20919 11569 20971
rect 11621 20919 11677 20971
rect 11729 20919 11749 20971
rect 11549 20863 11749 20919
rect 11549 20811 11569 20863
rect 11621 20811 11677 20863
rect 11729 20811 11749 20863
rect 11549 20755 11749 20811
rect 11549 20703 11569 20755
rect 11621 20703 11677 20755
rect 11729 20703 11749 20755
rect 11549 20647 11749 20703
rect 11549 20595 11569 20647
rect 11621 20595 11677 20647
rect 11729 20595 11749 20647
rect 11549 20539 11749 20595
rect 11549 20487 11569 20539
rect 11621 20487 11677 20539
rect 11729 20487 11749 20539
rect 11549 20431 11749 20487
rect 11549 20379 11569 20431
rect 11621 20379 11677 20431
rect 11729 20379 11749 20431
rect 11549 20323 11749 20379
rect 11549 20271 11569 20323
rect 11621 20271 11677 20323
rect 11729 20271 11749 20323
rect 11549 20215 11749 20271
rect 11549 20163 11569 20215
rect 11621 20163 11677 20215
rect 11729 20163 11749 20215
rect 11549 20107 11749 20163
rect 11549 20055 11569 20107
rect 11621 20055 11677 20107
rect 11729 20055 11749 20107
rect 11549 19999 11749 20055
rect 11549 19947 11569 19999
rect 11621 19947 11677 19999
rect 11729 19947 11749 19999
rect 11549 19891 11749 19947
rect 11549 19839 11569 19891
rect 11621 19839 11677 19891
rect 11729 19839 11749 19891
rect 11549 19783 11749 19839
rect 11549 19731 11569 19783
rect 11621 19731 11677 19783
rect 11729 19731 11749 19783
rect 11549 19675 11749 19731
rect 11549 19623 11569 19675
rect 11621 19623 11677 19675
rect 11729 19623 11749 19675
rect 11549 19567 11749 19623
rect 11549 19515 11569 19567
rect 11621 19515 11677 19567
rect 11729 19515 11749 19567
rect 11549 19459 11749 19515
rect 11549 19407 11569 19459
rect 11621 19407 11677 19459
rect 11729 19407 11749 19459
rect 11549 19351 11749 19407
rect 11549 19299 11569 19351
rect 11621 19299 11677 19351
rect 11729 19299 11749 19351
rect 11549 19243 11749 19299
rect 11549 19191 11569 19243
rect 11621 19191 11677 19243
rect 11729 19191 11749 19243
rect 11549 19135 11749 19191
rect 11549 19083 11569 19135
rect 11621 19083 11677 19135
rect 11729 19083 11749 19135
rect 11549 18015 11749 19083
rect 11549 17963 11569 18015
rect 11621 17963 11677 18015
rect 11729 17963 11749 18015
rect 11549 17907 11749 17963
rect 11549 17855 11569 17907
rect 11621 17855 11677 17907
rect 11729 17855 11749 17907
rect 11549 17799 11749 17855
rect 11549 17747 11569 17799
rect 11621 17747 11677 17799
rect 11729 17747 11749 17799
rect 11549 17691 11749 17747
rect 11549 17639 11569 17691
rect 11621 17639 11677 17691
rect 11729 17639 11749 17691
rect 11549 17583 11749 17639
rect 11549 17531 11569 17583
rect 11621 17531 11677 17583
rect 11729 17531 11749 17583
rect 11549 17475 11749 17531
rect 11549 17423 11569 17475
rect 11621 17423 11677 17475
rect 11729 17423 11749 17475
rect 11549 17367 11749 17423
rect 11549 17315 11569 17367
rect 11621 17315 11677 17367
rect 11729 17315 11749 17367
rect 11549 17259 11749 17315
rect 11549 17207 11569 17259
rect 11621 17207 11677 17259
rect 11729 17207 11749 17259
rect 11549 17151 11749 17207
rect 11549 17099 11569 17151
rect 11621 17099 11677 17151
rect 11729 17099 11749 17151
rect 11549 17043 11749 17099
rect 11549 16991 11569 17043
rect 11621 16991 11677 17043
rect 11729 16991 11749 17043
rect 11549 16935 11749 16991
rect 11549 16883 11569 16935
rect 11621 16883 11677 16935
rect 11729 16883 11749 16935
rect 11549 16827 11749 16883
rect 11549 16775 11569 16827
rect 11621 16775 11677 16827
rect 11729 16775 11749 16827
rect 11549 16719 11749 16775
rect 11549 16667 11569 16719
rect 11621 16667 11677 16719
rect 11729 16667 11749 16719
rect 11549 16611 11749 16667
rect 11549 16559 11569 16611
rect 11621 16559 11677 16611
rect 11729 16559 11749 16611
rect 11549 16503 11749 16559
rect 11549 16451 11569 16503
rect 11621 16451 11677 16503
rect 11729 16451 11749 16503
rect 11549 16395 11749 16451
rect 11549 16343 11569 16395
rect 11621 16343 11677 16395
rect 11729 16343 11749 16395
rect 11549 16287 11749 16343
rect 11549 16235 11569 16287
rect 11621 16235 11677 16287
rect 11729 16235 11749 16287
rect 11549 16179 11749 16235
rect 11549 16127 11569 16179
rect 11621 16127 11677 16179
rect 11729 16127 11749 16179
rect 11549 16071 11749 16127
rect 11549 16019 11569 16071
rect 11621 16019 11677 16071
rect 11729 16019 11749 16071
rect 11549 15963 11749 16019
rect 11549 15911 11569 15963
rect 11621 15911 11677 15963
rect 11729 15911 11749 15963
rect 11549 15855 11749 15911
rect 11549 15803 11569 15855
rect 11621 15803 11677 15855
rect 11729 15803 11749 15855
rect 11549 15747 11749 15803
rect 11549 15695 11569 15747
rect 11621 15695 11677 15747
rect 11729 15695 11749 15747
rect 11549 15639 11749 15695
rect 11549 15587 11569 15639
rect 11621 15587 11677 15639
rect 11729 15587 11749 15639
rect 11549 15531 11749 15587
rect 11549 15479 11569 15531
rect 11621 15479 11677 15531
rect 11729 15479 11749 15531
rect 11549 15423 11749 15479
rect 11549 15371 11569 15423
rect 11621 15371 11677 15423
rect 11729 15371 11749 15423
rect 11549 15315 11749 15371
rect 11549 15263 11569 15315
rect 11621 15263 11677 15315
rect 11729 15263 11749 15315
rect 11549 15207 11749 15263
rect 11549 15155 11569 15207
rect 11621 15155 11677 15207
rect 11729 15155 11749 15207
rect 11549 15099 11749 15155
rect 11549 15047 11569 15099
rect 11621 15047 11677 15099
rect 11729 15047 11749 15099
rect 11549 14991 11749 15047
rect 11549 14939 11569 14991
rect 11621 14939 11677 14991
rect 11729 14939 11749 14991
rect 11549 14883 11749 14939
rect 11549 14831 11569 14883
rect 11621 14831 11677 14883
rect 11729 14831 11749 14883
rect 11549 14775 11749 14831
rect 11549 14723 11569 14775
rect 11621 14723 11677 14775
rect 11729 14723 11749 14775
rect 11549 14667 11749 14723
rect 11549 14615 11569 14667
rect 11621 14615 11677 14667
rect 11729 14615 11749 14667
rect 11549 14559 11749 14615
rect 11549 14507 11569 14559
rect 11621 14507 11677 14559
rect 11729 14507 11749 14559
rect 11549 14451 11749 14507
rect 11549 14399 11569 14451
rect 11621 14399 11677 14451
rect 11729 14399 11749 14451
rect 11549 14343 11749 14399
rect 11549 14291 11569 14343
rect 11621 14291 11677 14343
rect 11729 14291 11749 14343
rect 11549 14235 11749 14291
rect 11549 14183 11569 14235
rect 11621 14183 11677 14235
rect 11729 14183 11749 14235
rect 11549 14127 11749 14183
rect 11549 14075 11569 14127
rect 11621 14075 11677 14127
rect 11729 14075 11749 14127
rect 11549 14019 11749 14075
rect 11549 13967 11569 14019
rect 11621 13967 11677 14019
rect 11729 13967 11749 14019
rect 11549 13911 11749 13967
rect 11549 13859 11569 13911
rect 11621 13859 11677 13911
rect 11729 13859 11749 13911
rect 11549 13803 11749 13859
rect 11549 13751 11569 13803
rect 11621 13751 11677 13803
rect 11729 13751 11749 13803
rect 11549 13695 11749 13751
rect 11549 13643 11569 13695
rect 11621 13643 11677 13695
rect 11729 13643 11749 13695
rect 11549 13587 11749 13643
rect 11549 13535 11569 13587
rect 11621 13535 11677 13587
rect 11729 13535 11749 13587
rect 11549 13479 11749 13535
rect 11549 13427 11569 13479
rect 11621 13427 11677 13479
rect 11729 13427 11749 13479
rect 11549 13371 11749 13427
rect 11549 13319 11569 13371
rect 11621 13319 11677 13371
rect 11729 13319 11749 13371
rect 11549 13263 11749 13319
rect 11549 13211 11569 13263
rect 11621 13211 11677 13263
rect 11729 13211 11749 13263
rect 11549 12143 11749 13211
rect 11549 12091 11569 12143
rect 11621 12091 11677 12143
rect 11729 12091 11749 12143
rect 11549 12035 11749 12091
rect 11549 11983 11569 12035
rect 11621 11983 11677 12035
rect 11729 11983 11749 12035
rect 11549 11927 11749 11983
rect 11549 11875 11569 11927
rect 11621 11875 11677 11927
rect 11729 11875 11749 11927
rect 11549 11819 11749 11875
rect 11549 11767 11569 11819
rect 11621 11767 11677 11819
rect 11729 11767 11749 11819
rect 11549 11711 11749 11767
rect 11549 11659 11569 11711
rect 11621 11659 11677 11711
rect 11729 11659 11749 11711
rect 11549 11603 11749 11659
rect 11549 11551 11569 11603
rect 11621 11551 11677 11603
rect 11729 11551 11749 11603
rect 11549 11495 11749 11551
rect 11549 11443 11569 11495
rect 11621 11443 11677 11495
rect 11729 11443 11749 11495
rect 11549 11387 11749 11443
rect 11549 11335 11569 11387
rect 11621 11335 11677 11387
rect 11729 11335 11749 11387
rect 11549 11279 11749 11335
rect 11549 11227 11569 11279
rect 11621 11227 11677 11279
rect 11729 11227 11749 11279
rect 11549 11171 11749 11227
rect 11549 11119 11569 11171
rect 11621 11119 11677 11171
rect 11729 11119 11749 11171
rect 11549 11063 11749 11119
rect 11549 11011 11569 11063
rect 11621 11011 11677 11063
rect 11729 11011 11749 11063
rect 11549 10955 11749 11011
rect 11549 10903 11569 10955
rect 11621 10903 11677 10955
rect 11729 10903 11749 10955
rect 11549 10847 11749 10903
rect 11549 10795 11569 10847
rect 11621 10795 11677 10847
rect 11729 10795 11749 10847
rect 11549 10739 11749 10795
rect 11549 10687 11569 10739
rect 11621 10687 11677 10739
rect 11729 10687 11749 10739
rect 11549 10631 11749 10687
rect 11549 10579 11569 10631
rect 11621 10579 11677 10631
rect 11729 10579 11749 10631
rect 11549 10523 11749 10579
rect 11549 10471 11569 10523
rect 11621 10471 11677 10523
rect 11729 10471 11749 10523
rect 11549 10415 11749 10471
rect 11549 10363 11569 10415
rect 11621 10363 11677 10415
rect 11729 10363 11749 10415
rect 11549 10307 11749 10363
rect 11549 10255 11569 10307
rect 11621 10255 11677 10307
rect 11729 10255 11749 10307
rect 11549 10199 11749 10255
rect 11549 10147 11569 10199
rect 11621 10147 11677 10199
rect 11729 10147 11749 10199
rect 11549 10091 11749 10147
rect 11549 10039 11569 10091
rect 11621 10039 11677 10091
rect 11729 10039 11749 10091
rect 11549 9983 11749 10039
rect 11549 9931 11569 9983
rect 11621 9931 11677 9983
rect 11729 9931 11749 9983
rect 11549 9875 11749 9931
rect 11549 9823 11569 9875
rect 11621 9823 11677 9875
rect 11729 9823 11749 9875
rect 11549 9767 11749 9823
rect 11549 9715 11569 9767
rect 11621 9715 11677 9767
rect 11729 9715 11749 9767
rect 11549 9659 11749 9715
rect 11549 9607 11569 9659
rect 11621 9607 11677 9659
rect 11729 9607 11749 9659
rect 11549 9551 11749 9607
rect 11549 9499 11569 9551
rect 11621 9499 11677 9551
rect 11729 9499 11749 9551
rect 11549 9443 11749 9499
rect 11549 9391 11569 9443
rect 11621 9391 11677 9443
rect 11729 9391 11749 9443
rect 11549 9335 11749 9391
rect 11549 9283 11569 9335
rect 11621 9283 11677 9335
rect 11729 9283 11749 9335
rect 11549 9227 11749 9283
rect 11549 9175 11569 9227
rect 11621 9175 11677 9227
rect 11729 9175 11749 9227
rect 11549 9119 11749 9175
rect 11549 9067 11569 9119
rect 11621 9067 11677 9119
rect 11729 9067 11749 9119
rect 11549 9011 11749 9067
rect 11549 8959 11569 9011
rect 11621 8959 11677 9011
rect 11729 8959 11749 9011
rect 11549 8903 11749 8959
rect 11549 8851 11569 8903
rect 11621 8851 11677 8903
rect 11729 8851 11749 8903
rect 11549 8795 11749 8851
rect 11549 8743 11569 8795
rect 11621 8743 11677 8795
rect 11729 8743 11749 8795
rect 11549 8687 11749 8743
rect 11549 8635 11569 8687
rect 11621 8635 11677 8687
rect 11729 8635 11749 8687
rect 11549 8579 11749 8635
rect 11549 8527 11569 8579
rect 11621 8527 11677 8579
rect 11729 8527 11749 8579
rect 11549 8471 11749 8527
rect 11549 8419 11569 8471
rect 11621 8419 11677 8471
rect 11729 8419 11749 8471
rect 11549 8363 11749 8419
rect 11549 8311 11569 8363
rect 11621 8311 11677 8363
rect 11729 8311 11749 8363
rect 11549 8255 11749 8311
rect 11549 8203 11569 8255
rect 11621 8203 11677 8255
rect 11729 8203 11749 8255
rect 11549 8147 11749 8203
rect 11549 8095 11569 8147
rect 11621 8095 11677 8147
rect 11729 8095 11749 8147
rect 11549 8039 11749 8095
rect 11549 7987 11569 8039
rect 11621 7987 11677 8039
rect 11729 7987 11749 8039
rect 11549 7931 11749 7987
rect 11549 7879 11569 7931
rect 11621 7879 11677 7931
rect 11729 7879 11749 7931
rect 11549 7823 11749 7879
rect 11549 7771 11569 7823
rect 11621 7771 11677 7823
rect 11729 7771 11749 7823
rect 11549 7715 11749 7771
rect 11549 7663 11569 7715
rect 11621 7663 11677 7715
rect 11729 7663 11749 7715
rect 11549 7607 11749 7663
rect 11549 7555 11569 7607
rect 11621 7555 11677 7607
rect 11729 7555 11749 7607
rect 11549 7499 11749 7555
rect 11549 7447 11569 7499
rect 11621 7447 11677 7499
rect 11729 7447 11749 7499
rect 11549 7391 11749 7447
rect 11549 7339 11569 7391
rect 11621 7339 11677 7391
rect 11729 7339 11749 7391
rect 11549 6271 11749 7339
rect 11549 6219 11569 6271
rect 11621 6219 11677 6271
rect 11729 6219 11749 6271
rect 11549 6163 11749 6219
rect 11549 6111 11569 6163
rect 11621 6111 11677 6163
rect 11729 6111 11749 6163
rect 11549 6055 11749 6111
rect 11549 6003 11569 6055
rect 11621 6003 11677 6055
rect 11729 6003 11749 6055
rect 11549 5947 11749 6003
rect 11549 5895 11569 5947
rect 11621 5895 11677 5947
rect 11729 5895 11749 5947
rect 11549 5839 11749 5895
rect 11549 5787 11569 5839
rect 11621 5787 11677 5839
rect 11729 5787 11749 5839
rect 11549 5731 11749 5787
rect 11549 5679 11569 5731
rect 11621 5679 11677 5731
rect 11729 5679 11749 5731
rect 11549 5623 11749 5679
rect 11549 5571 11569 5623
rect 11621 5571 11677 5623
rect 11729 5571 11749 5623
rect 11549 5515 11749 5571
rect 11549 5463 11569 5515
rect 11621 5463 11677 5515
rect 11729 5463 11749 5515
rect 11549 5407 11749 5463
rect 11549 5355 11569 5407
rect 11621 5355 11677 5407
rect 11729 5355 11749 5407
rect 11549 5299 11749 5355
rect 11549 5247 11569 5299
rect 11621 5247 11677 5299
rect 11729 5247 11749 5299
rect 11549 5191 11749 5247
rect 11549 5139 11569 5191
rect 11621 5139 11677 5191
rect 11729 5139 11749 5191
rect 11549 5083 11749 5139
rect 11549 5031 11569 5083
rect 11621 5031 11677 5083
rect 11729 5031 11749 5083
rect 11549 4975 11749 5031
rect 11549 4923 11569 4975
rect 11621 4923 11677 4975
rect 11729 4923 11749 4975
rect 11549 4867 11749 4923
rect 11549 4815 11569 4867
rect 11621 4815 11677 4867
rect 11729 4815 11749 4867
rect 11549 4759 11749 4815
rect 11549 4707 11569 4759
rect 11621 4707 11677 4759
rect 11729 4707 11749 4759
rect 11549 4651 11749 4707
rect 11549 4599 11569 4651
rect 11621 4599 11677 4651
rect 11729 4599 11749 4651
rect 11549 4543 11749 4599
rect 11549 4491 11569 4543
rect 11621 4491 11677 4543
rect 11729 4491 11749 4543
rect 11549 4435 11749 4491
rect 11549 4383 11569 4435
rect 11621 4383 11677 4435
rect 11729 4383 11749 4435
rect 11549 4327 11749 4383
rect 11549 4275 11569 4327
rect 11621 4275 11677 4327
rect 11729 4275 11749 4327
rect 11549 4219 11749 4275
rect 11549 4167 11569 4219
rect 11621 4167 11677 4219
rect 11729 4167 11749 4219
rect 11549 4111 11749 4167
rect 11549 4059 11569 4111
rect 11621 4059 11677 4111
rect 11729 4059 11749 4111
rect 11549 4003 11749 4059
rect 11549 3951 11569 4003
rect 11621 3951 11677 4003
rect 11729 3951 11749 4003
rect 11549 3895 11749 3951
rect 11549 3843 11569 3895
rect 11621 3843 11677 3895
rect 11729 3843 11749 3895
rect 11549 3787 11749 3843
rect 11549 3735 11569 3787
rect 11621 3735 11677 3787
rect 11729 3735 11749 3787
rect 11549 3679 11749 3735
rect 11549 3627 11569 3679
rect 11621 3627 11677 3679
rect 11729 3627 11749 3679
rect 11549 3571 11749 3627
rect 11549 3519 11569 3571
rect 11621 3519 11677 3571
rect 11729 3519 11749 3571
rect 11549 3463 11749 3519
rect 11549 3411 11569 3463
rect 11621 3411 11677 3463
rect 11729 3411 11749 3463
rect 11549 3355 11749 3411
rect 11549 3303 11569 3355
rect 11621 3303 11677 3355
rect 11729 3303 11749 3355
rect 11549 3247 11749 3303
rect 11549 3195 11569 3247
rect 11621 3195 11677 3247
rect 11729 3195 11749 3247
rect 11549 3139 11749 3195
rect 11549 3087 11569 3139
rect 11621 3087 11677 3139
rect 11729 3087 11749 3139
rect 11549 3031 11749 3087
rect 11549 2979 11569 3031
rect 11621 2979 11677 3031
rect 11729 2979 11749 3031
rect 11549 2923 11749 2979
rect 11549 2871 11569 2923
rect 11621 2871 11677 2923
rect 11729 2871 11749 2923
rect 11549 2815 11749 2871
rect 11549 2763 11569 2815
rect 11621 2763 11677 2815
rect 11729 2763 11749 2815
rect 11549 2707 11749 2763
rect 11549 2655 11569 2707
rect 11621 2655 11677 2707
rect 11729 2655 11749 2707
rect 11549 2599 11749 2655
rect 11549 2547 11569 2599
rect 11621 2547 11677 2599
rect 11729 2547 11749 2599
rect 11549 2491 11749 2547
rect 11549 2439 11569 2491
rect 11621 2439 11677 2491
rect 11729 2439 11749 2491
rect 11549 2383 11749 2439
rect 11549 2331 11569 2383
rect 11621 2331 11677 2383
rect 11729 2331 11749 2383
rect 11549 2275 11749 2331
rect 11549 2223 11569 2275
rect 11621 2223 11677 2275
rect 11729 2223 11749 2275
rect 11549 2167 11749 2223
rect 11549 2115 11569 2167
rect 11621 2115 11677 2167
rect 11729 2115 11749 2167
rect 11549 2059 11749 2115
rect 11549 2007 11569 2059
rect 11621 2007 11677 2059
rect 11729 2007 11749 2059
rect 11549 1951 11749 2007
rect 11549 1899 11569 1951
rect 11621 1899 11677 1951
rect 11729 1899 11749 1951
rect 11549 1843 11749 1899
rect 11549 1791 11569 1843
rect 11621 1791 11677 1843
rect 11729 1791 11749 1843
rect 11549 1735 11749 1791
rect 11549 1683 11569 1735
rect 11621 1683 11677 1735
rect 11729 1683 11749 1735
rect 11549 1627 11749 1683
rect 11549 1575 11569 1627
rect 11621 1575 11677 1627
rect 11729 1575 11749 1627
rect 11549 1519 11749 1575
rect 11549 1467 11569 1519
rect 11621 1467 11677 1519
rect 11729 1467 11749 1519
rect 11549 1455 11749 1467
rect 11817 24637 12919 25617
rect 11817 24585 12051 24637
rect 12103 24585 12159 24637
rect 12211 24585 12267 24637
rect 12319 24585 12919 24637
rect 11817 24529 12919 24585
rect 11817 24477 12051 24529
rect 12103 24477 12159 24529
rect 12211 24477 12267 24529
rect 12319 24477 12919 24529
rect 11817 24421 12919 24477
rect 11817 24369 12051 24421
rect 12103 24369 12159 24421
rect 12211 24369 12267 24421
rect 12319 24369 12919 24421
rect 11817 24313 12919 24369
rect 11817 24261 12051 24313
rect 12103 24261 12159 24313
rect 12211 24261 12267 24313
rect 12319 24261 12919 24313
rect 11817 24205 12919 24261
rect 11817 24153 12051 24205
rect 12103 24153 12159 24205
rect 12211 24153 12267 24205
rect 12319 24153 12919 24205
rect 11817 24097 12919 24153
rect 11817 24045 12051 24097
rect 12103 24045 12159 24097
rect 12211 24045 12267 24097
rect 12319 24045 12919 24097
rect 11817 23989 12919 24045
rect 11817 23937 12051 23989
rect 12103 23937 12159 23989
rect 12211 23937 12267 23989
rect 12319 23937 12919 23989
rect 11817 23881 12919 23937
rect 11817 23829 12051 23881
rect 12103 23829 12159 23881
rect 12211 23829 12267 23881
rect 12319 23829 12919 23881
rect 11817 23773 12919 23829
rect 11817 23721 12051 23773
rect 12103 23721 12159 23773
rect 12211 23721 12267 23773
rect 12319 23721 12919 23773
rect 11817 23665 12919 23721
rect 11817 23613 12051 23665
rect 12103 23613 12159 23665
rect 12211 23613 12267 23665
rect 12319 23613 12919 23665
rect 11817 23557 12919 23613
rect 11817 23505 12051 23557
rect 12103 23505 12159 23557
rect 12211 23505 12267 23557
rect 12319 23505 12919 23557
rect 11817 23449 12919 23505
rect 11817 23397 12051 23449
rect 12103 23397 12159 23449
rect 12211 23397 12267 23449
rect 12319 23397 12919 23449
rect 11817 23341 12919 23397
rect 11817 23289 12051 23341
rect 12103 23289 12159 23341
rect 12211 23289 12267 23341
rect 12319 23289 12919 23341
rect 11817 23233 12919 23289
rect 11817 23181 12051 23233
rect 12103 23181 12159 23233
rect 12211 23181 12267 23233
rect 12319 23181 12919 23233
rect 11817 23125 12919 23181
rect 11817 23073 12051 23125
rect 12103 23073 12159 23125
rect 12211 23073 12267 23125
rect 12319 23073 12919 23125
rect 11817 23017 12919 23073
rect 11817 22965 12051 23017
rect 12103 22965 12159 23017
rect 12211 22965 12267 23017
rect 12319 22965 12919 23017
rect 11817 22909 12919 22965
rect 11817 22857 12051 22909
rect 12103 22857 12159 22909
rect 12211 22857 12267 22909
rect 12319 22857 12919 22909
rect 11817 22801 12919 22857
rect 11817 22749 12051 22801
rect 12103 22749 12159 22801
rect 12211 22749 12267 22801
rect 12319 22749 12919 22801
rect 11817 22693 12919 22749
rect 11817 22641 12051 22693
rect 12103 22641 12159 22693
rect 12211 22641 12267 22693
rect 12319 22641 12919 22693
rect 11817 22585 12919 22641
rect 11817 22533 12051 22585
rect 12103 22533 12159 22585
rect 12211 22533 12267 22585
rect 12319 22533 12919 22585
rect 11817 22477 12919 22533
rect 11817 22425 12051 22477
rect 12103 22425 12159 22477
rect 12211 22425 12267 22477
rect 12319 22425 12919 22477
rect 11817 22369 12919 22425
rect 11817 22317 12051 22369
rect 12103 22317 12159 22369
rect 12211 22317 12267 22369
rect 12319 22317 12919 22369
rect 11817 22261 12919 22317
rect 11817 22209 12051 22261
rect 12103 22209 12159 22261
rect 12211 22209 12267 22261
rect 12319 22209 12919 22261
rect 11817 22153 12919 22209
rect 11817 22101 12051 22153
rect 12103 22101 12159 22153
rect 12211 22101 12267 22153
rect 12319 22101 12919 22153
rect 11817 22045 12919 22101
rect 11817 21993 12051 22045
rect 12103 21993 12159 22045
rect 12211 21993 12267 22045
rect 12319 21993 12919 22045
rect 11817 21937 12919 21993
rect 11817 21885 12051 21937
rect 12103 21885 12159 21937
rect 12211 21885 12267 21937
rect 12319 21885 12919 21937
rect 11817 21829 12919 21885
rect 11817 21777 12051 21829
rect 12103 21777 12159 21829
rect 12211 21777 12267 21829
rect 12319 21777 12919 21829
rect 11817 21721 12919 21777
rect 11817 21669 12051 21721
rect 12103 21669 12159 21721
rect 12211 21669 12267 21721
rect 12319 21669 12919 21721
rect 11817 21613 12919 21669
rect 11817 21561 12051 21613
rect 12103 21561 12159 21613
rect 12211 21561 12267 21613
rect 12319 21561 12919 21613
rect 11817 21505 12919 21561
rect 11817 21453 12051 21505
rect 12103 21453 12159 21505
rect 12211 21453 12267 21505
rect 12319 21453 12919 21505
rect 11817 21397 12919 21453
rect 11817 21345 12051 21397
rect 12103 21345 12159 21397
rect 12211 21345 12267 21397
rect 12319 21345 12919 21397
rect 11817 21289 12919 21345
rect 11817 21237 12051 21289
rect 12103 21237 12159 21289
rect 12211 21237 12267 21289
rect 12319 21237 12919 21289
rect 11817 21181 12919 21237
rect 11817 21129 12051 21181
rect 12103 21129 12159 21181
rect 12211 21129 12267 21181
rect 12319 21129 12919 21181
rect 11817 21073 12919 21129
rect 11817 21021 12051 21073
rect 12103 21021 12159 21073
rect 12211 21021 12267 21073
rect 12319 21021 12919 21073
rect 11817 20965 12919 21021
rect 11817 20913 12051 20965
rect 12103 20913 12159 20965
rect 12211 20913 12267 20965
rect 12319 20913 12919 20965
rect 11817 20857 12919 20913
rect 11817 20805 12051 20857
rect 12103 20805 12159 20857
rect 12211 20805 12267 20857
rect 12319 20805 12919 20857
rect 11817 20749 12919 20805
rect 11817 20697 12051 20749
rect 12103 20697 12159 20749
rect 12211 20697 12267 20749
rect 12319 20697 12919 20749
rect 11817 20641 12919 20697
rect 11817 20589 12051 20641
rect 12103 20589 12159 20641
rect 12211 20589 12267 20641
rect 12319 20589 12919 20641
rect 11817 20533 12919 20589
rect 11817 20481 12051 20533
rect 12103 20481 12159 20533
rect 12211 20481 12267 20533
rect 12319 20481 12919 20533
rect 11817 20425 12919 20481
rect 11817 20373 12051 20425
rect 12103 20373 12159 20425
rect 12211 20373 12267 20425
rect 12319 20373 12919 20425
rect 11817 20317 12919 20373
rect 11817 20265 12051 20317
rect 12103 20265 12159 20317
rect 12211 20265 12267 20317
rect 12319 20265 12919 20317
rect 11817 20209 12919 20265
rect 11817 20157 12051 20209
rect 12103 20157 12159 20209
rect 12211 20157 12267 20209
rect 12319 20157 12919 20209
rect 11817 20101 12919 20157
rect 11817 20049 12051 20101
rect 12103 20049 12159 20101
rect 12211 20049 12267 20101
rect 12319 20049 12919 20101
rect 11817 19993 12919 20049
rect 11817 19941 12051 19993
rect 12103 19941 12159 19993
rect 12211 19941 12267 19993
rect 12319 19941 12919 19993
rect 11817 19885 12919 19941
rect 11817 19833 12051 19885
rect 12103 19833 12159 19885
rect 12211 19833 12267 19885
rect 12319 19833 12919 19885
rect 11817 19777 12919 19833
rect 11817 19725 12051 19777
rect 12103 19725 12159 19777
rect 12211 19725 12267 19777
rect 12319 19725 12919 19777
rect 11817 19669 12919 19725
rect 11817 19617 12051 19669
rect 12103 19617 12159 19669
rect 12211 19617 12267 19669
rect 12319 19617 12919 19669
rect 11817 19561 12919 19617
rect 11817 19509 12051 19561
rect 12103 19509 12159 19561
rect 12211 19509 12267 19561
rect 12319 19509 12919 19561
rect 11817 19453 12919 19509
rect 11817 19401 12051 19453
rect 12103 19401 12159 19453
rect 12211 19401 12267 19453
rect 12319 19401 12919 19453
rect 11817 19345 12919 19401
rect 11817 19293 12051 19345
rect 12103 19293 12159 19345
rect 12211 19293 12267 19345
rect 12319 19293 12919 19345
rect 11817 19237 12919 19293
rect 11817 19185 12051 19237
rect 12103 19185 12159 19237
rect 12211 19185 12267 19237
rect 12319 19185 12919 19237
rect 11817 19129 12919 19185
rect 11817 19077 12051 19129
rect 12103 19077 12159 19129
rect 12211 19077 12267 19129
rect 12319 19077 12919 19129
rect 11817 19021 12919 19077
rect 11817 18969 12051 19021
rect 12103 18969 12159 19021
rect 12211 18969 12267 19021
rect 12319 18969 12919 19021
rect 11817 18913 12919 18969
rect 11817 18861 12051 18913
rect 12103 18861 12159 18913
rect 12211 18861 12267 18913
rect 12319 18861 12919 18913
rect 11817 18805 12919 18861
rect 11817 18753 12051 18805
rect 12103 18753 12159 18805
rect 12211 18753 12267 18805
rect 12319 18753 12919 18805
rect 11817 18697 12919 18753
rect 11817 18645 12051 18697
rect 12103 18645 12159 18697
rect 12211 18645 12267 18697
rect 12319 18645 12919 18697
rect 11817 18589 12919 18645
rect 11817 18537 12051 18589
rect 12103 18537 12159 18589
rect 12211 18537 12267 18589
rect 12319 18537 12919 18589
rect 11817 18481 12919 18537
rect 11817 18429 12051 18481
rect 12103 18429 12159 18481
rect 12211 18429 12267 18481
rect 12319 18429 12919 18481
rect 11817 18373 12919 18429
rect 11817 18321 12051 18373
rect 12103 18321 12159 18373
rect 12211 18321 12267 18373
rect 12319 18321 12919 18373
rect 11817 18265 12919 18321
rect 11817 18213 12051 18265
rect 12103 18213 12159 18265
rect 12211 18213 12267 18265
rect 12319 18213 12919 18265
rect 11817 18157 12919 18213
rect 11817 18105 12051 18157
rect 12103 18105 12159 18157
rect 12211 18105 12267 18157
rect 12319 18105 12919 18157
rect 11817 18049 12919 18105
rect 11817 17997 12051 18049
rect 12103 17997 12159 18049
rect 12211 17997 12267 18049
rect 12319 17997 12919 18049
rect 11817 17941 12919 17997
rect 11817 17889 12051 17941
rect 12103 17889 12159 17941
rect 12211 17889 12267 17941
rect 12319 17889 12919 17941
rect 11817 17833 12919 17889
rect 11817 17781 12051 17833
rect 12103 17781 12159 17833
rect 12211 17781 12267 17833
rect 12319 17781 12919 17833
rect 11817 17725 12919 17781
rect 11817 17673 12051 17725
rect 12103 17673 12159 17725
rect 12211 17673 12267 17725
rect 12319 17673 12919 17725
rect 11817 17617 12919 17673
rect 11817 17565 12051 17617
rect 12103 17565 12159 17617
rect 12211 17565 12267 17617
rect 12319 17565 12919 17617
rect 11817 17509 12919 17565
rect 11817 17457 12051 17509
rect 12103 17457 12159 17509
rect 12211 17457 12267 17509
rect 12319 17457 12919 17509
rect 11817 17401 12919 17457
rect 11817 17349 12051 17401
rect 12103 17349 12159 17401
rect 12211 17349 12267 17401
rect 12319 17349 12919 17401
rect 11817 17293 12919 17349
rect 11817 17241 12051 17293
rect 12103 17241 12159 17293
rect 12211 17241 12267 17293
rect 12319 17241 12919 17293
rect 11817 17185 12919 17241
rect 11817 17133 12051 17185
rect 12103 17133 12159 17185
rect 12211 17133 12267 17185
rect 12319 17133 12919 17185
rect 11817 17077 12919 17133
rect 11817 17025 12051 17077
rect 12103 17025 12159 17077
rect 12211 17025 12267 17077
rect 12319 17025 12919 17077
rect 11817 16969 12919 17025
rect 11817 16917 12051 16969
rect 12103 16917 12159 16969
rect 12211 16917 12267 16969
rect 12319 16917 12919 16969
rect 11817 16861 12919 16917
rect 11817 16809 12051 16861
rect 12103 16809 12159 16861
rect 12211 16809 12267 16861
rect 12319 16809 12919 16861
rect 11817 16753 12919 16809
rect 11817 16701 12051 16753
rect 12103 16701 12159 16753
rect 12211 16701 12267 16753
rect 12319 16701 12919 16753
rect 11817 16645 12919 16701
rect 11817 16593 12051 16645
rect 12103 16593 12159 16645
rect 12211 16593 12267 16645
rect 12319 16593 12919 16645
rect 11817 16537 12919 16593
rect 11817 16485 12051 16537
rect 12103 16485 12159 16537
rect 12211 16485 12267 16537
rect 12319 16485 12919 16537
rect 11817 16429 12919 16485
rect 11817 16377 12051 16429
rect 12103 16377 12159 16429
rect 12211 16377 12267 16429
rect 12319 16377 12919 16429
rect 11817 16321 12919 16377
rect 11817 16269 12051 16321
rect 12103 16269 12159 16321
rect 12211 16269 12267 16321
rect 12319 16269 12919 16321
rect 11817 16213 12919 16269
rect 11817 16161 12051 16213
rect 12103 16161 12159 16213
rect 12211 16161 12267 16213
rect 12319 16161 12919 16213
rect 11817 16105 12919 16161
rect 11817 16053 12051 16105
rect 12103 16053 12159 16105
rect 12211 16053 12267 16105
rect 12319 16053 12919 16105
rect 11817 15997 12919 16053
rect 11817 15945 12051 15997
rect 12103 15945 12159 15997
rect 12211 15945 12267 15997
rect 12319 15945 12919 15997
rect 11817 15889 12919 15945
rect 11817 15837 12051 15889
rect 12103 15837 12159 15889
rect 12211 15837 12267 15889
rect 12319 15837 12919 15889
rect 11817 15781 12919 15837
rect 11817 15729 12051 15781
rect 12103 15729 12159 15781
rect 12211 15729 12267 15781
rect 12319 15729 12919 15781
rect 11817 15673 12919 15729
rect 11817 15621 12051 15673
rect 12103 15621 12159 15673
rect 12211 15621 12267 15673
rect 12319 15621 12919 15673
rect 11817 15565 12919 15621
rect 11817 15513 12051 15565
rect 12103 15513 12159 15565
rect 12211 15513 12267 15565
rect 12319 15513 12919 15565
rect 11817 15457 12919 15513
rect 11817 15405 12051 15457
rect 12103 15405 12159 15457
rect 12211 15405 12267 15457
rect 12319 15405 12919 15457
rect 11817 15349 12919 15405
rect 11817 15297 12051 15349
rect 12103 15297 12159 15349
rect 12211 15297 12267 15349
rect 12319 15297 12919 15349
rect 11817 15241 12919 15297
rect 11817 15189 12051 15241
rect 12103 15189 12159 15241
rect 12211 15189 12267 15241
rect 12319 15189 12919 15241
rect 11817 15133 12919 15189
rect 11817 15081 12051 15133
rect 12103 15081 12159 15133
rect 12211 15081 12267 15133
rect 12319 15081 12919 15133
rect 11817 15025 12919 15081
rect 11817 14973 12051 15025
rect 12103 14973 12159 15025
rect 12211 14973 12267 15025
rect 12319 14973 12919 15025
rect 11817 14917 12919 14973
rect 11817 14865 12051 14917
rect 12103 14865 12159 14917
rect 12211 14865 12267 14917
rect 12319 14865 12919 14917
rect 11817 14809 12919 14865
rect 11817 14757 12051 14809
rect 12103 14757 12159 14809
rect 12211 14757 12267 14809
rect 12319 14757 12919 14809
rect 11817 14701 12919 14757
rect 11817 14649 12051 14701
rect 12103 14649 12159 14701
rect 12211 14649 12267 14701
rect 12319 14649 12919 14701
rect 11817 14593 12919 14649
rect 11817 14541 12051 14593
rect 12103 14541 12159 14593
rect 12211 14541 12267 14593
rect 12319 14541 12919 14593
rect 11817 14485 12919 14541
rect 11817 14433 12051 14485
rect 12103 14433 12159 14485
rect 12211 14433 12267 14485
rect 12319 14433 12919 14485
rect 11817 14377 12919 14433
rect 11817 14325 12051 14377
rect 12103 14325 12159 14377
rect 12211 14325 12267 14377
rect 12319 14325 12919 14377
rect 11817 14269 12919 14325
rect 11817 14217 12051 14269
rect 12103 14217 12159 14269
rect 12211 14217 12267 14269
rect 12319 14217 12919 14269
rect 11817 14161 12919 14217
rect 11817 14109 12051 14161
rect 12103 14109 12159 14161
rect 12211 14109 12267 14161
rect 12319 14109 12919 14161
rect 11817 14053 12919 14109
rect 11817 14001 12051 14053
rect 12103 14001 12159 14053
rect 12211 14001 12267 14053
rect 12319 14001 12919 14053
rect 11817 13945 12919 14001
rect 11817 13893 12051 13945
rect 12103 13893 12159 13945
rect 12211 13893 12267 13945
rect 12319 13893 12919 13945
rect 11817 13837 12919 13893
rect 11817 13785 12051 13837
rect 12103 13785 12159 13837
rect 12211 13785 12267 13837
rect 12319 13785 12919 13837
rect 11817 13729 12919 13785
rect 11817 13677 12051 13729
rect 12103 13677 12159 13729
rect 12211 13677 12267 13729
rect 12319 13677 12919 13729
rect 11817 13621 12919 13677
rect 11817 13569 12051 13621
rect 12103 13569 12159 13621
rect 12211 13569 12267 13621
rect 12319 13569 12919 13621
rect 11817 13513 12919 13569
rect 11817 13461 12051 13513
rect 12103 13461 12159 13513
rect 12211 13461 12267 13513
rect 12319 13461 12919 13513
rect 11817 13405 12919 13461
rect 11817 13353 12051 13405
rect 12103 13353 12159 13405
rect 12211 13353 12267 13405
rect 12319 13353 12919 13405
rect 11817 13297 12919 13353
rect 11817 13245 12051 13297
rect 12103 13245 12159 13297
rect 12211 13245 12267 13297
rect 12319 13245 12919 13297
rect 11817 13189 12919 13245
rect 11817 13137 12051 13189
rect 12103 13137 12159 13189
rect 12211 13137 12267 13189
rect 12319 13137 12919 13189
rect 11817 13081 12919 13137
rect 11817 13029 12051 13081
rect 12103 13029 12159 13081
rect 12211 13029 12267 13081
rect 12319 13029 12919 13081
rect 11817 12973 12919 13029
rect 11817 12921 12051 12973
rect 12103 12921 12159 12973
rect 12211 12921 12267 12973
rect 12319 12921 12919 12973
rect 11817 12865 12919 12921
rect 11817 12813 12051 12865
rect 12103 12813 12159 12865
rect 12211 12813 12267 12865
rect 12319 12813 12919 12865
rect 11817 12757 12919 12813
rect 11817 12705 12051 12757
rect 12103 12705 12159 12757
rect 12211 12705 12267 12757
rect 12319 12705 12919 12757
rect 11817 12649 12919 12705
rect 11817 12597 12051 12649
rect 12103 12597 12159 12649
rect 12211 12597 12267 12649
rect 12319 12597 12919 12649
rect 11817 12541 12919 12597
rect 11817 12489 12051 12541
rect 12103 12489 12159 12541
rect 12211 12489 12267 12541
rect 12319 12489 12919 12541
rect 11817 12433 12919 12489
rect 11817 12381 12051 12433
rect 12103 12381 12159 12433
rect 12211 12381 12267 12433
rect 12319 12381 12919 12433
rect 11817 12325 12919 12381
rect 11817 12273 12051 12325
rect 12103 12273 12159 12325
rect 12211 12273 12267 12325
rect 12319 12273 12919 12325
rect 11817 12217 12919 12273
rect 11817 12165 12051 12217
rect 12103 12165 12159 12217
rect 12211 12165 12267 12217
rect 12319 12165 12919 12217
rect 11817 12109 12919 12165
rect 11817 12057 12051 12109
rect 12103 12057 12159 12109
rect 12211 12057 12267 12109
rect 12319 12057 12919 12109
rect 11817 12001 12919 12057
rect 11817 11949 12051 12001
rect 12103 11949 12159 12001
rect 12211 11949 12267 12001
rect 12319 11949 12919 12001
rect 11817 11893 12919 11949
rect 11817 11841 12051 11893
rect 12103 11841 12159 11893
rect 12211 11841 12267 11893
rect 12319 11841 12919 11893
rect 11817 11785 12919 11841
rect 11817 11733 12051 11785
rect 12103 11733 12159 11785
rect 12211 11733 12267 11785
rect 12319 11733 12919 11785
rect 11817 11677 12919 11733
rect 11817 11625 12051 11677
rect 12103 11625 12159 11677
rect 12211 11625 12267 11677
rect 12319 11625 12919 11677
rect 11817 11569 12919 11625
rect 11817 11517 12051 11569
rect 12103 11517 12159 11569
rect 12211 11517 12267 11569
rect 12319 11517 12919 11569
rect 11817 11461 12919 11517
rect 11817 11409 12051 11461
rect 12103 11409 12159 11461
rect 12211 11409 12267 11461
rect 12319 11409 12919 11461
rect 11817 11353 12919 11409
rect 11817 11301 12051 11353
rect 12103 11301 12159 11353
rect 12211 11301 12267 11353
rect 12319 11301 12919 11353
rect 11817 11245 12919 11301
rect 11817 11193 12051 11245
rect 12103 11193 12159 11245
rect 12211 11193 12267 11245
rect 12319 11193 12919 11245
rect 11817 11137 12919 11193
rect 11817 11085 12051 11137
rect 12103 11085 12159 11137
rect 12211 11085 12267 11137
rect 12319 11085 12919 11137
rect 11817 11029 12919 11085
rect 11817 10977 12051 11029
rect 12103 10977 12159 11029
rect 12211 10977 12267 11029
rect 12319 10977 12919 11029
rect 11817 10921 12919 10977
rect 11817 10869 12051 10921
rect 12103 10869 12159 10921
rect 12211 10869 12267 10921
rect 12319 10869 12919 10921
rect 11817 10813 12919 10869
rect 11817 10761 12051 10813
rect 12103 10761 12159 10813
rect 12211 10761 12267 10813
rect 12319 10761 12919 10813
rect 11817 10705 12919 10761
rect 11817 10653 12051 10705
rect 12103 10653 12159 10705
rect 12211 10653 12267 10705
rect 12319 10653 12919 10705
rect 11817 10597 12919 10653
rect 11817 10545 12051 10597
rect 12103 10545 12159 10597
rect 12211 10545 12267 10597
rect 12319 10545 12919 10597
rect 11817 10489 12919 10545
rect 11817 10437 12051 10489
rect 12103 10437 12159 10489
rect 12211 10437 12267 10489
rect 12319 10437 12919 10489
rect 11817 10381 12919 10437
rect 11817 10329 12051 10381
rect 12103 10329 12159 10381
rect 12211 10329 12267 10381
rect 12319 10329 12919 10381
rect 11817 10273 12919 10329
rect 11817 10221 12051 10273
rect 12103 10221 12159 10273
rect 12211 10221 12267 10273
rect 12319 10221 12919 10273
rect 11817 10165 12919 10221
rect 11817 10113 12051 10165
rect 12103 10113 12159 10165
rect 12211 10113 12267 10165
rect 12319 10113 12919 10165
rect 11817 10057 12919 10113
rect 11817 10005 12051 10057
rect 12103 10005 12159 10057
rect 12211 10005 12267 10057
rect 12319 10005 12919 10057
rect 11817 9949 12919 10005
rect 11817 9897 12051 9949
rect 12103 9897 12159 9949
rect 12211 9897 12267 9949
rect 12319 9897 12919 9949
rect 11817 9841 12919 9897
rect 11817 9789 12051 9841
rect 12103 9789 12159 9841
rect 12211 9789 12267 9841
rect 12319 9789 12919 9841
rect 11817 9733 12919 9789
rect 11817 9681 12051 9733
rect 12103 9681 12159 9733
rect 12211 9681 12267 9733
rect 12319 9681 12919 9733
rect 11817 9625 12919 9681
rect 11817 9573 12051 9625
rect 12103 9573 12159 9625
rect 12211 9573 12267 9625
rect 12319 9573 12919 9625
rect 11817 9517 12919 9573
rect 11817 9465 12051 9517
rect 12103 9465 12159 9517
rect 12211 9465 12267 9517
rect 12319 9465 12919 9517
rect 11817 9409 12919 9465
rect 11817 9357 12051 9409
rect 12103 9357 12159 9409
rect 12211 9357 12267 9409
rect 12319 9357 12919 9409
rect 11817 9301 12919 9357
rect 11817 9249 12051 9301
rect 12103 9249 12159 9301
rect 12211 9249 12267 9301
rect 12319 9249 12919 9301
rect 11817 9193 12919 9249
rect 11817 9141 12051 9193
rect 12103 9141 12159 9193
rect 12211 9141 12267 9193
rect 12319 9141 12919 9193
rect 11817 9085 12919 9141
rect 11817 9033 12051 9085
rect 12103 9033 12159 9085
rect 12211 9033 12267 9085
rect 12319 9033 12919 9085
rect 11817 8977 12919 9033
rect 11817 8925 12051 8977
rect 12103 8925 12159 8977
rect 12211 8925 12267 8977
rect 12319 8925 12919 8977
rect 11817 8869 12919 8925
rect 11817 8817 12051 8869
rect 12103 8817 12159 8869
rect 12211 8817 12267 8869
rect 12319 8817 12919 8869
rect 11817 8761 12919 8817
rect 11817 8709 12051 8761
rect 12103 8709 12159 8761
rect 12211 8709 12267 8761
rect 12319 8709 12919 8761
rect 11817 8653 12919 8709
rect 11817 8601 12051 8653
rect 12103 8601 12159 8653
rect 12211 8601 12267 8653
rect 12319 8601 12919 8653
rect 11817 8545 12919 8601
rect 11817 8493 12051 8545
rect 12103 8493 12159 8545
rect 12211 8493 12267 8545
rect 12319 8493 12919 8545
rect 11817 8437 12919 8493
rect 11817 8385 12051 8437
rect 12103 8385 12159 8437
rect 12211 8385 12267 8437
rect 12319 8385 12919 8437
rect 11817 8329 12919 8385
rect 11817 8277 12051 8329
rect 12103 8277 12159 8329
rect 12211 8277 12267 8329
rect 12319 8277 12919 8329
rect 11817 8221 12919 8277
rect 11817 8169 12051 8221
rect 12103 8169 12159 8221
rect 12211 8169 12267 8221
rect 12319 8169 12919 8221
rect 11817 8113 12919 8169
rect 11817 8061 12051 8113
rect 12103 8061 12159 8113
rect 12211 8061 12267 8113
rect 12319 8061 12919 8113
rect 11817 8005 12919 8061
rect 11817 7953 12051 8005
rect 12103 7953 12159 8005
rect 12211 7953 12267 8005
rect 12319 7953 12919 8005
rect 11817 7897 12919 7953
rect 11817 7845 12051 7897
rect 12103 7845 12159 7897
rect 12211 7845 12267 7897
rect 12319 7845 12919 7897
rect 11817 7789 12919 7845
rect 11817 7737 12051 7789
rect 12103 7737 12159 7789
rect 12211 7737 12267 7789
rect 12319 7737 12919 7789
rect 11817 7681 12919 7737
rect 11817 7629 12051 7681
rect 12103 7629 12159 7681
rect 12211 7629 12267 7681
rect 12319 7629 12919 7681
rect 11817 7573 12919 7629
rect 11817 7521 12051 7573
rect 12103 7521 12159 7573
rect 12211 7521 12267 7573
rect 12319 7521 12919 7573
rect 11817 7465 12919 7521
rect 11817 7413 12051 7465
rect 12103 7413 12159 7465
rect 12211 7413 12267 7465
rect 12319 7413 12919 7465
rect 11817 7357 12919 7413
rect 11817 7305 12051 7357
rect 12103 7305 12159 7357
rect 12211 7305 12267 7357
rect 12319 7305 12919 7357
rect 11817 7249 12919 7305
rect 11817 7197 12051 7249
rect 12103 7197 12159 7249
rect 12211 7197 12267 7249
rect 12319 7197 12919 7249
rect 11817 7141 12919 7197
rect 11817 7089 12051 7141
rect 12103 7089 12159 7141
rect 12211 7089 12267 7141
rect 12319 7089 12919 7141
rect 11817 7033 12919 7089
rect 11817 6981 12051 7033
rect 12103 6981 12159 7033
rect 12211 6981 12267 7033
rect 12319 6981 12919 7033
rect 11817 6925 12919 6981
rect 11817 6873 12051 6925
rect 12103 6873 12159 6925
rect 12211 6873 12267 6925
rect 12319 6873 12919 6925
rect 11817 6817 12919 6873
rect 11817 6765 12051 6817
rect 12103 6765 12159 6817
rect 12211 6765 12267 6817
rect 12319 6765 12919 6817
rect 11817 6709 12919 6765
rect 11817 6657 12051 6709
rect 12103 6657 12159 6709
rect 12211 6657 12267 6709
rect 12319 6657 12919 6709
rect 11817 6601 12919 6657
rect 11817 6549 12051 6601
rect 12103 6549 12159 6601
rect 12211 6549 12267 6601
rect 12319 6549 12919 6601
rect 11817 6493 12919 6549
rect 11817 6441 12051 6493
rect 12103 6441 12159 6493
rect 12211 6441 12267 6493
rect 12319 6441 12919 6493
rect 11817 6385 12919 6441
rect 11817 6333 12051 6385
rect 12103 6333 12159 6385
rect 12211 6333 12267 6385
rect 12319 6333 12919 6385
rect 11817 6277 12919 6333
rect 11817 6225 12051 6277
rect 12103 6225 12159 6277
rect 12211 6225 12267 6277
rect 12319 6225 12919 6277
rect 11817 6169 12919 6225
rect 11817 6117 12051 6169
rect 12103 6117 12159 6169
rect 12211 6117 12267 6169
rect 12319 6117 12919 6169
rect 11817 6061 12919 6117
rect 11817 6009 12051 6061
rect 12103 6009 12159 6061
rect 12211 6009 12267 6061
rect 12319 6009 12919 6061
rect 11817 5953 12919 6009
rect 11817 5901 12051 5953
rect 12103 5901 12159 5953
rect 12211 5901 12267 5953
rect 12319 5901 12919 5953
rect 11817 5845 12919 5901
rect 11817 5793 12051 5845
rect 12103 5793 12159 5845
rect 12211 5793 12267 5845
rect 12319 5793 12919 5845
rect 11817 5737 12919 5793
rect 11817 5685 12051 5737
rect 12103 5685 12159 5737
rect 12211 5685 12267 5737
rect 12319 5685 12919 5737
rect 11817 5629 12919 5685
rect 11817 5577 12051 5629
rect 12103 5577 12159 5629
rect 12211 5577 12267 5629
rect 12319 5577 12919 5629
rect 11817 5521 12919 5577
rect 11817 5469 12051 5521
rect 12103 5469 12159 5521
rect 12211 5469 12267 5521
rect 12319 5469 12919 5521
rect 11817 5413 12919 5469
rect 11817 5361 12051 5413
rect 12103 5361 12159 5413
rect 12211 5361 12267 5413
rect 12319 5361 12919 5413
rect 11817 5305 12919 5361
rect 11817 5253 12051 5305
rect 12103 5253 12159 5305
rect 12211 5253 12267 5305
rect 12319 5253 12919 5305
rect 11817 5197 12919 5253
rect 11817 5145 12051 5197
rect 12103 5145 12159 5197
rect 12211 5145 12267 5197
rect 12319 5145 12919 5197
rect 11817 5089 12919 5145
rect 11817 5037 12051 5089
rect 12103 5037 12159 5089
rect 12211 5037 12267 5089
rect 12319 5037 12919 5089
rect 11817 4981 12919 5037
rect 11817 4929 12051 4981
rect 12103 4929 12159 4981
rect 12211 4929 12267 4981
rect 12319 4929 12919 4981
rect 11817 4873 12919 4929
rect 11817 4821 12051 4873
rect 12103 4821 12159 4873
rect 12211 4821 12267 4873
rect 12319 4821 12919 4873
rect 11817 4765 12919 4821
rect 11817 4713 12051 4765
rect 12103 4713 12159 4765
rect 12211 4713 12267 4765
rect 12319 4713 12919 4765
rect 11817 4657 12919 4713
rect 11817 4605 12051 4657
rect 12103 4605 12159 4657
rect 12211 4605 12267 4657
rect 12319 4605 12919 4657
rect 11817 4549 12919 4605
rect 11817 4497 12051 4549
rect 12103 4497 12159 4549
rect 12211 4497 12267 4549
rect 12319 4497 12919 4549
rect 11817 4441 12919 4497
rect 11817 4389 12051 4441
rect 12103 4389 12159 4441
rect 12211 4389 12267 4441
rect 12319 4389 12919 4441
rect 11817 4333 12919 4389
rect 11817 4281 12051 4333
rect 12103 4281 12159 4333
rect 12211 4281 12267 4333
rect 12319 4281 12919 4333
rect 11817 4225 12919 4281
rect 11817 4173 12051 4225
rect 12103 4173 12159 4225
rect 12211 4173 12267 4225
rect 12319 4173 12919 4225
rect 11817 4117 12919 4173
rect 11817 4065 12051 4117
rect 12103 4065 12159 4117
rect 12211 4065 12267 4117
rect 12319 4065 12919 4117
rect 11817 4009 12919 4065
rect 11817 3957 12051 4009
rect 12103 3957 12159 4009
rect 12211 3957 12267 4009
rect 12319 3957 12919 4009
rect 11817 3901 12919 3957
rect 11817 3849 12051 3901
rect 12103 3849 12159 3901
rect 12211 3849 12267 3901
rect 12319 3849 12919 3901
rect 11817 3793 12919 3849
rect 11817 3741 12051 3793
rect 12103 3741 12159 3793
rect 12211 3741 12267 3793
rect 12319 3741 12919 3793
rect 11817 3685 12919 3741
rect 11817 3633 12051 3685
rect 12103 3633 12159 3685
rect 12211 3633 12267 3685
rect 12319 3633 12919 3685
rect 11817 3577 12919 3633
rect 11817 3525 12051 3577
rect 12103 3525 12159 3577
rect 12211 3525 12267 3577
rect 12319 3525 12919 3577
rect 11817 3469 12919 3525
rect 11817 3417 12051 3469
rect 12103 3417 12159 3469
rect 12211 3417 12267 3469
rect 12319 3417 12919 3469
rect 11817 3361 12919 3417
rect 11817 3309 12051 3361
rect 12103 3309 12159 3361
rect 12211 3309 12267 3361
rect 12319 3309 12919 3361
rect 11817 3253 12919 3309
rect 11817 3201 12051 3253
rect 12103 3201 12159 3253
rect 12211 3201 12267 3253
rect 12319 3201 12919 3253
rect 11817 3145 12919 3201
rect 11817 3093 12051 3145
rect 12103 3093 12159 3145
rect 12211 3093 12267 3145
rect 12319 3093 12919 3145
rect 11817 3037 12919 3093
rect 11817 2985 12051 3037
rect 12103 2985 12159 3037
rect 12211 2985 12267 3037
rect 12319 2985 12919 3037
rect 11817 2929 12919 2985
rect 11817 2877 12051 2929
rect 12103 2877 12159 2929
rect 12211 2877 12267 2929
rect 12319 2877 12919 2929
rect 11817 2821 12919 2877
rect 11817 2769 12051 2821
rect 12103 2769 12159 2821
rect 12211 2769 12267 2821
rect 12319 2769 12919 2821
rect 11817 2713 12919 2769
rect 11817 2661 12051 2713
rect 12103 2661 12159 2713
rect 12211 2661 12267 2713
rect 12319 2661 12919 2713
rect 11817 2605 12919 2661
rect 11817 2553 12051 2605
rect 12103 2553 12159 2605
rect 12211 2553 12267 2605
rect 12319 2553 12919 2605
rect 11817 2497 12919 2553
rect 11817 2445 12051 2497
rect 12103 2445 12159 2497
rect 12211 2445 12267 2497
rect 12319 2445 12919 2497
rect 11817 2389 12919 2445
rect 11817 2337 12051 2389
rect 12103 2337 12159 2389
rect 12211 2337 12267 2389
rect 12319 2337 12919 2389
rect 11817 2281 12919 2337
rect 11817 2229 12051 2281
rect 12103 2229 12159 2281
rect 12211 2229 12267 2281
rect 12319 2229 12919 2281
rect 11817 2173 12919 2229
rect 11817 2121 12051 2173
rect 12103 2121 12159 2173
rect 12211 2121 12267 2173
rect 12319 2121 12919 2173
rect 11817 2065 12919 2121
rect 11817 2013 12051 2065
rect 12103 2013 12159 2065
rect 12211 2013 12267 2065
rect 12319 2013 12919 2065
rect 11817 1957 12919 2013
rect 11817 1905 12051 1957
rect 12103 1905 12159 1957
rect 12211 1905 12267 1957
rect 12319 1905 12919 1957
rect 11817 1849 12919 1905
rect 11817 1797 12051 1849
rect 12103 1797 12159 1849
rect 12211 1797 12267 1849
rect 12319 1797 12919 1849
rect 11817 1741 12919 1797
rect 11817 1689 12051 1741
rect 12103 1689 12159 1741
rect 12211 1689 12267 1741
rect 12319 1689 12919 1741
rect 11817 1633 12919 1689
rect 11817 1581 12051 1633
rect 12103 1581 12159 1633
rect 12211 1581 12267 1633
rect 12319 1581 12919 1633
rect 11817 1525 12919 1581
rect 11817 1473 12051 1525
rect 12103 1473 12159 1525
rect 12211 1473 12267 1525
rect 12319 1473 12919 1525
rect 9653 1403 9677 1455
rect 9729 1403 9785 1455
rect 9837 1403 9893 1455
rect 9945 1403 10001 1455
rect 10053 1403 10109 1455
rect 10161 1403 10217 1455
rect 10269 1403 10325 1455
rect 10377 1403 10433 1455
rect 10485 1403 10541 1455
rect 10593 1403 10649 1455
rect 10701 1403 10757 1455
rect 10809 1403 10865 1455
rect 10917 1403 10973 1455
rect 11025 1403 11081 1455
rect 11133 1403 11189 1455
rect 11241 1403 11297 1455
rect 11349 1403 11405 1455
rect 11457 1403 11481 1455
rect 9653 361 11481 1403
rect 9653 309 9677 361
rect 9729 309 9785 361
rect 9837 309 9893 361
rect 9945 309 10001 361
rect 10053 309 10109 361
rect 10161 309 10217 361
rect 10269 309 10325 361
rect 10377 309 10433 361
rect 10485 309 10541 361
rect 10593 309 10649 361
rect 10701 309 10757 361
rect 10809 309 10865 361
rect 10917 309 10973 361
rect 11025 309 11081 361
rect 11133 309 11189 361
rect 11241 309 11297 361
rect 11349 309 11405 361
rect 11457 309 11481 361
rect 9653 253 11481 309
rect 9653 201 9677 253
rect 9729 201 9785 253
rect 9837 201 9893 253
rect 9945 201 10001 253
rect 10053 201 10109 253
rect 10161 201 10217 253
rect 10269 201 10325 253
rect 10377 201 10433 253
rect 10485 201 10541 253
rect 10593 201 10649 253
rect 10701 201 10757 253
rect 10809 201 10865 253
rect 10917 201 10973 253
rect 11025 201 11081 253
rect 11133 201 11189 253
rect 11241 201 11297 253
rect 11349 201 11405 253
rect 11457 201 11481 253
rect 9653 145 11481 201
rect 9653 93 9677 145
rect 9729 93 9785 145
rect 9837 93 9893 145
rect 9945 93 10001 145
rect 10053 93 10109 145
rect 10161 93 10217 145
rect 10269 93 10325 145
rect 10377 93 10433 145
rect 10485 93 10541 145
rect 10593 93 10649 145
rect 10701 93 10757 145
rect 10809 93 10865 145
rect 10917 93 10973 145
rect 11025 93 11081 145
rect 11133 93 11189 145
rect 11241 93 11297 145
rect 11349 93 11405 145
rect 11457 93 11481 145
rect 9653 43 11481 93
rect 11817 1417 12919 1473
rect 11817 1365 12051 1417
rect 12103 1365 12159 1417
rect 12211 1365 12267 1417
rect 12319 1365 12919 1417
rect 11817 1309 12919 1365
rect 11817 1257 12051 1309
rect 12103 1257 12159 1309
rect 12211 1257 12267 1309
rect 12319 1257 12919 1309
rect 11817 1201 12919 1257
rect 11817 1149 12051 1201
rect 12103 1149 12159 1201
rect 12211 1149 12267 1201
rect 12319 1149 12919 1201
rect 11817 1093 12919 1149
rect 11817 1041 12051 1093
rect 12103 1041 12159 1093
rect 12211 1041 12267 1093
rect 12319 1041 12919 1093
rect 11817 985 12919 1041
rect 11817 933 12051 985
rect 12103 933 12159 985
rect 12211 933 12267 985
rect 12319 933 12919 985
rect 11817 877 12919 933
rect 11817 825 12051 877
rect 12103 825 12159 877
rect 12211 825 12267 877
rect 12319 825 12919 877
rect 11817 769 12919 825
rect 11817 717 12051 769
rect 12103 717 12159 769
rect 12211 717 12267 769
rect 12319 717 12919 769
rect 11817 43 12919 717
use M1_NWELL_CDNS_40661956134135  M1_NWELL_CDNS_40661956134135_0
timestamp 1698431365
transform 1 0 227 0 1 12677
box 0 0 1 1
use M1_NWELL_CDNS_40661956134135  M1_NWELL_CDNS_40661956134135_1
timestamp 1698431365
transform 1 0 12735 0 1 12677
box 0 0 1 1
use M1_NWELL_CDNS_40661956134139  M1_NWELL_CDNS_40661956134139_0
timestamp 1698431365
transform 1 0 6481 0 1 227
box 0 0 1 1
use M1_NWELL_CDNS_40661956134139  M1_NWELL_CDNS_40661956134139_1
timestamp 1698431365
transform 1 0 6481 0 1 25127
box 0 0 1 1
use M1_POLY2_CDNS_40661956134136  M1_POLY2_CDNS_40661956134136_0
timestamp 1698431365
transform -1 0 11633 0 1 9741
box 0 0 1 1
use M1_POLY2_CDNS_40661956134136  M1_POLY2_CDNS_40661956134136_1
timestamp 1698431365
transform -1 0 11633 0 1 3869
box 0 0 1 1
use M1_POLY2_CDNS_40661956134136  M1_POLY2_CDNS_40661956134136_2
timestamp 1698431365
transform 1 0 1329 0 1 3869
box 0 0 1 1
use M1_POLY2_CDNS_40661956134136  M1_POLY2_CDNS_40661956134136_3
timestamp 1698431365
transform 1 0 1329 0 1 9741
box 0 0 1 1
use M1_POLY2_CDNS_40661956134136  M1_POLY2_CDNS_40661956134136_4
timestamp 1698431365
transform 1 0 1329 0 1 15613
box 0 0 1 1
use M1_POLY2_CDNS_40661956134136  M1_POLY2_CDNS_40661956134136_5
timestamp 1698431365
transform 1 0 1329 0 1 21485
box 0 0 1 1
use M1_POLY2_CDNS_40661956134136  M1_POLY2_CDNS_40661956134136_6
timestamp 1698431365
transform -1 0 11633 0 1 15613
box 0 0 1 1
use M1_POLY2_CDNS_40661956134136  M1_POLY2_CDNS_40661956134136_7
timestamp 1698431365
transform -1 0 11633 0 1 21485
box 0 0 1 1
use M1_PSUB_CDNS_40661956134134  M1_PSUB_CDNS_40661956134134_0
timestamp 1698431365
transform 1 0 6481 0 1 6805
box 0 0 1 1
use M1_PSUB_CDNS_40661956134134  M1_PSUB_CDNS_40661956134134_1
timestamp 1698431365
transform 1 0 6481 0 1 18549
box 0 0 1 1
use M1_PSUB_CDNS_40661956134134  M1_PSUB_CDNS_40661956134134_2
timestamp 1698431365
transform 1 0 6481 0 1 12677
box 0 0 1 1
use M1_PSUB_CDNS_40661956134137  M1_PSUB_CDNS_40661956134137_0
timestamp 1698431365
transform 1 0 12185 0 1 12677
box 0 0 1 1
use M1_PSUB_CDNS_40661956134137  M1_PSUB_CDNS_40661956134137_1
timestamp 1698431365
transform 1 0 777 0 1 12677
box 0 0 1 1
use M1_PSUB_CDNS_40661956134138  M1_PSUB_CDNS_40661956134138_0
timestamp 1698431365
transform 1 0 6481 0 1 24527
box 0 0 1 1
use M1_PSUB_CDNS_40661956134138  M1_PSUB_CDNS_40661956134138_1
timestamp 1698431365
transform 1 0 6481 0 1 827
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_0
timestamp 1698431365
transform 1 0 10567 0 1 4845
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_1
timestamp 1698431365
transform 1 0 10567 0 1 4357
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_2
timestamp 1698431365
transform 1 0 10567 0 1 3869
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_3
timestamp 1698431365
transform 1 0 10567 0 1 3381
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_4
timestamp 1698431365
transform 1 0 10567 0 1 2893
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_5
timestamp 1698431365
transform 1 0 10567 0 1 2405
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_6
timestamp 1698431365
transform 1 0 10567 0 1 1917
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_7
timestamp 1698431365
transform 1 0 8639 0 1 6065
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_8
timestamp 1698431365
transform 1 0 8639 0 1 5577
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_9
timestamp 1698431365
transform 1 0 8639 0 1 5089
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_10
timestamp 1698431365
transform 1 0 8639 0 1 4601
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_11
timestamp 1698431365
transform 1 0 8639 0 1 4113
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_12
timestamp 1698431365
transform 1 0 8639 0 1 3625
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_13
timestamp 1698431365
transform 1 0 8639 0 1 3137
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_14
timestamp 1698431365
transform 1 0 8639 0 1 2649
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_15
timestamp 1698431365
transform 1 0 8639 0 1 2161
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_16
timestamp 1698431365
transform 1 0 8639 0 1 1673
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_17
timestamp 1698431365
transform 1 0 8639 0 1 11937
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_18
timestamp 1698431365
transform 1 0 8639 0 1 11449
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_19
timestamp 1698431365
transform 1 0 8639 0 1 10961
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_20
timestamp 1698431365
transform 1 0 8639 0 1 10473
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_21
timestamp 1698431365
transform 1 0 8639 0 1 9985
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_22
timestamp 1698431365
transform 1 0 8639 0 1 9497
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_23
timestamp 1698431365
transform 1 0 8639 0 1 9009
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_24
timestamp 1698431365
transform 1 0 8639 0 1 8521
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_25
timestamp 1698431365
transform 1 0 8639 0 1 8033
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_26
timestamp 1698431365
transform 1 0 10567 0 1 1429
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_27
timestamp 1698431365
transform 1 0 10567 0 1 7301
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_28
timestamp 1698431365
transform 1 0 10567 0 1 8277
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_29
timestamp 1698431365
transform 1 0 10567 0 1 8765
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_30
timestamp 1698431365
transform 1 0 10567 0 1 9253
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_31
timestamp 1698431365
transform 1 0 10567 0 1 9741
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_32
timestamp 1698431365
transform 1 0 10567 0 1 10229
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_33
timestamp 1698431365
transform 1 0 10567 0 1 10717
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_34
timestamp 1698431365
transform 1 0 10567 0 1 11205
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_35
timestamp 1698431365
transform 1 0 10567 0 1 11693
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_36
timestamp 1698431365
transform 1 0 10567 0 1 12181
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_37
timestamp 1698431365
transform 1 0 8639 0 1 7545
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_38
timestamp 1698431365
transform 1 0 10567 0 1 6309
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_39
timestamp 1698431365
transform 1 0 10567 0 1 5821
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_40
timestamp 1698431365
transform 1 0 10567 0 1 7789
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_41
timestamp 1698431365
transform 1 0 10567 0 1 5333
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_42
timestamp 1698431365
transform 1 0 4323 0 1 5333
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_43
timestamp 1698431365
transform 1 0 4323 0 1 4845
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_44
timestamp 1698431365
transform 1 0 4323 0 1 4357
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_45
timestamp 1698431365
transform 1 0 4323 0 1 3869
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_46
timestamp 1698431365
transform 1 0 4323 0 1 3381
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_47
timestamp 1698431365
transform 1 0 4323 0 1 2893
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_48
timestamp 1698431365
transform 1 0 4323 0 1 2405
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_49
timestamp 1698431365
transform 1 0 4323 0 1 1917
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_50
timestamp 1698431365
transform 1 0 4323 0 1 1429
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_51
timestamp 1698431365
transform 1 0 4323 0 1 5821
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_52
timestamp 1698431365
transform 1 0 2395 0 1 6065
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_53
timestamp 1698431365
transform 1 0 2395 0 1 9985
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_54
timestamp 1698431365
transform 1 0 2395 0 1 11937
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_55
timestamp 1698431365
transform 1 0 4323 0 1 11693
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_56
timestamp 1698431365
transform 1 0 2395 0 1 11449
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_57
timestamp 1698431365
transform 1 0 4323 0 1 11205
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_58
timestamp 1698431365
transform 1 0 2395 0 1 10961
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_59
timestamp 1698431365
transform 1 0 4323 0 1 10717
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_60
timestamp 1698431365
transform 1 0 2395 0 1 10473
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_61
timestamp 1698431365
transform 1 0 4323 0 1 10229
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_62
timestamp 1698431365
transform 1 0 4323 0 1 9741
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_63
timestamp 1698431365
transform 1 0 2395 0 1 9497
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_64
timestamp 1698431365
transform 1 0 4323 0 1 9253
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_65
timestamp 1698431365
transform 1 0 2395 0 1 9009
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_66
timestamp 1698431365
transform 1 0 4323 0 1 8765
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_67
timestamp 1698431365
transform 1 0 2395 0 1 8521
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_68
timestamp 1698431365
transform 1 0 4323 0 1 8277
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_69
timestamp 1698431365
transform 1 0 2395 0 1 8033
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_70
timestamp 1698431365
transform 1 0 4323 0 1 7789
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_71
timestamp 1698431365
transform 1 0 4323 0 1 7301
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_72
timestamp 1698431365
transform 1 0 4323 0 1 12181
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_73
timestamp 1698431365
transform 1 0 2395 0 1 7545
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_74
timestamp 1698431365
transform 1 0 2395 0 1 5577
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_75
timestamp 1698431365
transform 1 0 2395 0 1 5089
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_76
timestamp 1698431365
transform 1 0 2395 0 1 4601
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_77
timestamp 1698431365
transform 1 0 2395 0 1 4113
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_78
timestamp 1698431365
transform 1 0 2395 0 1 3625
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_79
timestamp 1698431365
transform 1 0 2395 0 1 3137
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_80
timestamp 1698431365
transform 1 0 2395 0 1 2649
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_81
timestamp 1698431365
transform 1 0 2395 0 1 2161
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_82
timestamp 1698431365
transform 1 0 2395 0 1 1673
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_83
timestamp 1698431365
transform 1 0 4323 0 1 6309
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_84
timestamp 1698431365
transform 1 0 4323 0 1 21973
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_85
timestamp 1698431365
transform 1 0 2395 0 1 19289
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_86
timestamp 1698431365
transform 1 0 4323 0 1 21485
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_87
timestamp 1698431365
transform 1 0 2395 0 1 21241
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_88
timestamp 1698431365
transform 1 0 4323 0 1 20997
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_89
timestamp 1698431365
transform 1 0 2395 0 1 20753
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_90
timestamp 1698431365
transform 1 0 4323 0 1 20509
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_91
timestamp 1698431365
transform 1 0 2395 0 1 20265
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_92
timestamp 1698431365
transform 1 0 4323 0 1 20021
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_93
timestamp 1698431365
transform 1 0 2395 0 1 19777
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_94
timestamp 1698431365
transform 1 0 4323 0 1 19533
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_95
timestamp 1698431365
transform 1 0 2395 0 1 21729
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_96
timestamp 1698431365
transform 1 0 4323 0 1 18053
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_97
timestamp 1698431365
transform 1 0 2395 0 1 17809
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_98
timestamp 1698431365
transform 1 0 4323 0 1 17565
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_99
timestamp 1698431365
transform 1 0 2395 0 1 17321
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_100
timestamp 1698431365
transform 1 0 4323 0 1 17077
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_101
timestamp 1698431365
transform 1 0 2395 0 1 16833
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_102
timestamp 1698431365
transform 1 0 4323 0 1 16589
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_103
timestamp 1698431365
transform 1 0 2395 0 1 16345
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_104
timestamp 1698431365
transform 1 0 2395 0 1 15857
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_105
timestamp 1698431365
transform 1 0 4323 0 1 15613
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_106
timestamp 1698431365
transform 1 0 2395 0 1 15369
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_107
timestamp 1698431365
transform 1 0 4323 0 1 15125
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_108
timestamp 1698431365
transform 1 0 2395 0 1 14881
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_109
timestamp 1698431365
transform 1 0 4323 0 1 14637
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_110
timestamp 1698431365
transform 1 0 2395 0 1 14393
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_111
timestamp 1698431365
transform 1 0 4323 0 1 14149
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_112
timestamp 1698431365
transform 1 0 2395 0 1 13905
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_113
timestamp 1698431365
transform 1 0 4323 0 1 16101
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_114
timestamp 1698431365
transform 1 0 4323 0 1 13661
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_115
timestamp 1698431365
transform 1 0 4323 0 1 19045
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_116
timestamp 1698431365
transform 1 0 4323 0 1 13173
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_117
timestamp 1698431365
transform 1 0 2395 0 1 13417
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_118
timestamp 1698431365
transform 1 0 4323 0 1 23925
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_119
timestamp 1698431365
transform 1 0 2395 0 1 23681
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_120
timestamp 1698431365
transform 1 0 4323 0 1 23437
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_121
timestamp 1698431365
transform 1 0 2395 0 1 23193
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_122
timestamp 1698431365
transform 1 0 4323 0 1 22949
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_123
timestamp 1698431365
transform 1 0 2395 0 1 22705
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_124
timestamp 1698431365
transform 1 0 4323 0 1 22461
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_125
timestamp 1698431365
transform 1 0 2395 0 1 22217
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_126
timestamp 1698431365
transform 1 0 10567 0 1 14637
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_127
timestamp 1698431365
transform 1 0 10567 0 1 14149
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_128
timestamp 1698431365
transform 1 0 10567 0 1 13173
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_129
timestamp 1698431365
transform 1 0 8639 0 1 13417
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_130
timestamp 1698431365
transform 1 0 8639 0 1 23681
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_131
timestamp 1698431365
transform 1 0 8639 0 1 23193
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_132
timestamp 1698431365
transform 1 0 8639 0 1 22705
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_133
timestamp 1698431365
transform 1 0 8639 0 1 22217
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_134
timestamp 1698431365
transform 1 0 8639 0 1 21729
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_135
timestamp 1698431365
transform 1 0 8639 0 1 21241
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_136
timestamp 1698431365
transform 1 0 8639 0 1 20753
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_137
timestamp 1698431365
transform 1 0 8639 0 1 20265
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_138
timestamp 1698431365
transform 1 0 8639 0 1 19777
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_139
timestamp 1698431365
transform 1 0 10567 0 1 19533
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_140
timestamp 1698431365
transform 1 0 10567 0 1 19045
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_141
timestamp 1698431365
transform 1 0 10567 0 1 20021
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_142
timestamp 1698431365
transform 1 0 10567 0 1 20509
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_143
timestamp 1698431365
transform 1 0 10567 0 1 20997
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_144
timestamp 1698431365
transform 1 0 10567 0 1 21485
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_145
timestamp 1698431365
transform 1 0 10567 0 1 21973
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_146
timestamp 1698431365
transform 1 0 10567 0 1 22461
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_147
timestamp 1698431365
transform 1 0 10567 0 1 22949
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_148
timestamp 1698431365
transform 1 0 10567 0 1 23437
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_149
timestamp 1698431365
transform 1 0 10567 0 1 23925
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_150
timestamp 1698431365
transform 1 0 8639 0 1 19289
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_151
timestamp 1698431365
transform 1 0 10567 0 1 13661
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_152
timestamp 1698431365
transform 1 0 10567 0 1 18053
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_153
timestamp 1698431365
transform 1 0 8639 0 1 17809
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_154
timestamp 1698431365
transform 1 0 8639 0 1 17321
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_155
timestamp 1698431365
transform 1 0 8639 0 1 16833
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_156
timestamp 1698431365
transform 1 0 8639 0 1 16345
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_157
timestamp 1698431365
transform 1 0 8639 0 1 15857
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_158
timestamp 1698431365
transform 1 0 8639 0 1 15369
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_159
timestamp 1698431365
transform 1 0 8639 0 1 14881
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_160
timestamp 1698431365
transform 1 0 8639 0 1 14393
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_161
timestamp 1698431365
transform 1 0 8639 0 1 13905
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_162
timestamp 1698431365
transform 1 0 10567 0 1 17565
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_163
timestamp 1698431365
transform 1 0 10567 0 1 17077
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_164
timestamp 1698431365
transform 1 0 10567 0 1 16589
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_165
timestamp 1698431365
transform 1 0 10567 0 1 16101
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_166
timestamp 1698431365
transform 1 0 10567 0 1 15613
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_167
timestamp 1698431365
transform 1 0 10567 0 1 15125
box 0 0 1 1
use M2_M1_CDNS_40661956134141  M2_M1_CDNS_40661956134141_0
timestamp 1698431365
transform 1 0 11649 0 1 3869
box 0 0 1 1
use M2_M1_CDNS_40661956134141  M2_M1_CDNS_40661956134141_1
timestamp 1698431365
transform 1 0 11649 0 1 9741
box 0 0 1 1
use M2_M1_CDNS_40661956134141  M2_M1_CDNS_40661956134141_2
timestamp 1698431365
transform 1 0 1313 0 1 9741
box 0 0 1 1
use M2_M1_CDNS_40661956134141  M2_M1_CDNS_40661956134141_3
timestamp 1698431365
transform 1 0 1313 0 1 3869
box 0 0 1 1
use M2_M1_CDNS_40661956134141  M2_M1_CDNS_40661956134141_4
timestamp 1698431365
transform 1 0 1313 0 1 21485
box 0 0 1 1
use M2_M1_CDNS_40661956134141  M2_M1_CDNS_40661956134141_5
timestamp 1698431365
transform 1 0 1313 0 1 15613
box 0 0 1 1
use M2_M1_CDNS_40661956134141  M2_M1_CDNS_40661956134141_6
timestamp 1698431365
transform 1 0 11649 0 1 15613
box 0 0 1 1
use M2_M1_CDNS_40661956134141  M2_M1_CDNS_40661956134141_7
timestamp 1698431365
transform 1 0 11649 0 1 21485
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_0
timestamp 1698431365
transform 1 0 7078 0 1 7301
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_1
timestamp 1698431365
transform 1 0 7078 0 1 7789
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_2
timestamp 1698431365
transform 1 0 7078 0 1 8277
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_3
timestamp 1698431365
transform 1 0 7078 0 1 8765
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_4
timestamp 1698431365
transform 1 0 7078 0 1 9253
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_5
timestamp 1698431365
transform 1 0 7078 0 1 12181
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_6
timestamp 1698431365
transform 1 0 7078 0 1 9741
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_7
timestamp 1698431365
transform 1 0 7078 0 1 10229
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_8
timestamp 1698431365
transform 1 0 7078 0 1 10717
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_9
timestamp 1698431365
transform 1 0 7078 0 1 11205
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_10
timestamp 1698431365
transform 1 0 7078 0 1 11693
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_11
timestamp 1698431365
transform 1 0 7078 0 1 6309
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_12
timestamp 1698431365
transform 1 0 7078 0 1 1429
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_13
timestamp 1698431365
transform 1 0 7078 0 1 1917
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_14
timestamp 1698431365
transform 1 0 7078 0 1 2405
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_15
timestamp 1698431365
transform 1 0 7078 0 1 2893
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_16
timestamp 1698431365
transform 1 0 7078 0 1 3381
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_17
timestamp 1698431365
transform 1 0 7078 0 1 3869
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_18
timestamp 1698431365
transform 1 0 7078 0 1 4357
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_19
timestamp 1698431365
transform 1 0 7078 0 1 4845
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_20
timestamp 1698431365
transform 1 0 7078 0 1 5333
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_21
timestamp 1698431365
transform 1 0 7078 0 1 5821
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_22
timestamp 1698431365
transform 1 0 5884 0 1 7545
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_23
timestamp 1698431365
transform 1 0 5884 0 1 8033
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_24
timestamp 1698431365
transform 1 0 5884 0 1 8521
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_25
timestamp 1698431365
transform 1 0 5884 0 1 9009
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_26
timestamp 1698431365
transform 1 0 5884 0 1 9985
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_27
timestamp 1698431365
transform 1 0 5884 0 1 10473
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_28
timestamp 1698431365
transform 1 0 5884 0 1 10961
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_29
timestamp 1698431365
transform 1 0 5884 0 1 11449
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_30
timestamp 1698431365
transform 1 0 5884 0 1 11937
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_31
timestamp 1698431365
transform 1 0 5884 0 1 9497
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_32
timestamp 1698431365
transform 1 0 5884 0 1 1673
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_33
timestamp 1698431365
transform 1 0 5884 0 1 2161
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_34
timestamp 1698431365
transform 1 0 5884 0 1 2649
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_35
timestamp 1698431365
transform 1 0 5884 0 1 3137
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_36
timestamp 1698431365
transform 1 0 5884 0 1 3625
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_37
timestamp 1698431365
transform 1 0 5884 0 1 4113
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_38
timestamp 1698431365
transform 1 0 5884 0 1 4601
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_39
timestamp 1698431365
transform 1 0 5884 0 1 5089
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_40
timestamp 1698431365
transform 1 0 5884 0 1 5577
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_41
timestamp 1698431365
transform 1 0 5884 0 1 6065
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_42
timestamp 1698431365
transform 1 0 5884 0 1 19289
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_43
timestamp 1698431365
transform 1 0 5884 0 1 19777
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_44
timestamp 1698431365
transform 1 0 5884 0 1 20265
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_45
timestamp 1698431365
transform 1 0 5884 0 1 20753
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_46
timestamp 1698431365
transform 1 0 5884 0 1 21729
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_47
timestamp 1698431365
transform 1 0 5884 0 1 22217
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_48
timestamp 1698431365
transform 1 0 5884 0 1 22705
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_49
timestamp 1698431365
transform 1 0 5884 0 1 23193
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_50
timestamp 1698431365
transform 1 0 5884 0 1 23681
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_51
timestamp 1698431365
transform 1 0 5884 0 1 21241
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_52
timestamp 1698431365
transform 1 0 5884 0 1 13417
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_53
timestamp 1698431365
transform 1 0 5884 0 1 13905
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_54
timestamp 1698431365
transform 1 0 5884 0 1 14393
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_55
timestamp 1698431365
transform 1 0 5884 0 1 14881
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_56
timestamp 1698431365
transform 1 0 5884 0 1 15369
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_57
timestamp 1698431365
transform 1 0 5884 0 1 15857
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_58
timestamp 1698431365
transform 1 0 5884 0 1 16345
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_59
timestamp 1698431365
transform 1 0 5884 0 1 16833
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_60
timestamp 1698431365
transform 1 0 5884 0 1 17321
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_61
timestamp 1698431365
transform 1 0 5884 0 1 17809
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_62
timestamp 1698431365
transform 1 0 7078 0 1 19045
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_63
timestamp 1698431365
transform 1 0 7078 0 1 19533
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_64
timestamp 1698431365
transform 1 0 7078 0 1 20021
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_65
timestamp 1698431365
transform 1 0 7078 0 1 20509
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_66
timestamp 1698431365
transform 1 0 7078 0 1 20997
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_67
timestamp 1698431365
transform 1 0 7078 0 1 18053
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_68
timestamp 1698431365
transform 1 0 7078 0 1 21485
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_69
timestamp 1698431365
transform 1 0 7078 0 1 21973
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_70
timestamp 1698431365
transform 1 0 7078 0 1 22461
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_71
timestamp 1698431365
transform 1 0 7078 0 1 22949
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_72
timestamp 1698431365
transform 1 0 7078 0 1 23437
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_73
timestamp 1698431365
transform 1 0 7078 0 1 13173
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_74
timestamp 1698431365
transform 1 0 7078 0 1 23925
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_75
timestamp 1698431365
transform 1 0 7078 0 1 13661
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_76
timestamp 1698431365
transform 1 0 7078 0 1 14149
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_77
timestamp 1698431365
transform 1 0 7078 0 1 14637
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_78
timestamp 1698431365
transform 1 0 7078 0 1 15125
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_79
timestamp 1698431365
transform 1 0 7078 0 1 15613
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_80
timestamp 1698431365
transform 1 0 7078 0 1 16101
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_81
timestamp 1698431365
transform 1 0 7078 0 1 16589
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_82
timestamp 1698431365
transform 1 0 7078 0 1 17077
box 0 0 1 1
use M2_M1_CDNS_40661956134142  M2_M1_CDNS_40661956134142_83
timestamp 1698431365
transform 1 0 7078 0 1 17565
box 0 0 1 1
use M2_M1_CDNS_40661956134143  M2_M1_CDNS_40661956134143_0
timestamp 1698431365
transform 1 0 8639 0 1 6805
box 0 0 1 1
use M2_M1_CDNS_40661956134143  M2_M1_CDNS_40661956134143_1
timestamp 1698431365
transform 1 0 2395 0 1 6805
box 0 0 1 1
use M2_M1_CDNS_40661956134143  M2_M1_CDNS_40661956134143_2
timestamp 1698431365
transform 1 0 2395 0 1 18549
box 0 0 1 1
use M2_M1_CDNS_40661956134143  M2_M1_CDNS_40661956134143_3
timestamp 1698431365
transform 1 0 8639 0 1 18549
box 0 0 1 1
use M2_M1_CDNS_40661956134143  M2_M1_CDNS_40661956134143_4
timestamp 1698431365
transform 1 0 8639 0 1 12677
box 0 0 1 1
use M2_M1_CDNS_40661956134143  M2_M1_CDNS_40661956134143_5
timestamp 1698431365
transform 1 0 2395 0 1 12677
box 0 0 1 1
use M2_M1_CDNS_40661956134144  M2_M1_CDNS_40661956134144_0
timestamp 1698431365
transform 1 0 8639 0 1 827
box 0 0 1 1
use M2_M1_CDNS_40661956134144  M2_M1_CDNS_40661956134144_1
timestamp 1698431365
transform 1 0 10567 0 1 227
box 0 0 1 1
use M2_M1_CDNS_40661956134144  M2_M1_CDNS_40661956134144_2
timestamp 1698431365
transform 1 0 2395 0 1 827
box 0 0 1 1
use M2_M1_CDNS_40661956134144  M2_M1_CDNS_40661956134144_3
timestamp 1698431365
transform 1 0 4323 0 1 227
box 0 0 1 1
use M2_M1_CDNS_40661956134144  M2_M1_CDNS_40661956134144_4
timestamp 1698431365
transform 1 0 4323 0 1 25127
box 0 0 1 1
use M2_M1_CDNS_40661956134144  M2_M1_CDNS_40661956134144_5
timestamp 1698431365
transform 1 0 2395 0 1 24527
box 0 0 1 1
use M2_M1_CDNS_40661956134144  M2_M1_CDNS_40661956134144_6
timestamp 1698431365
transform 1 0 8639 0 1 24527
box 0 0 1 1
use M2_M1_CDNS_40661956134144  M2_M1_CDNS_40661956134144_7
timestamp 1698431365
transform 1 0 10567 0 1 25127
box 0 0 1 1
use M2_M1_CDNS_40661956134145  M2_M1_CDNS_40661956134145_0
timestamp 1698431365
transform 1 0 7078 0 1 227
box 0 0 1 1
use M2_M1_CDNS_40661956134145  M2_M1_CDNS_40661956134145_1
timestamp 1698431365
transform 1 0 5884 0 1 827
box 0 0 1 1
use M2_M1_CDNS_40661956134145  M2_M1_CDNS_40661956134145_2
timestamp 1698431365
transform 1 0 594 0 1 227
box 0 0 1 1
use M2_M1_CDNS_40661956134145  M2_M1_CDNS_40661956134145_3
timestamp 1698431365
transform 1 0 594 0 1 25127
box 0 0 1 1
use M2_M1_CDNS_40661956134145  M2_M1_CDNS_40661956134145_4
timestamp 1698431365
transform 1 0 5884 0 1 24527
box 0 0 1 1
use M2_M1_CDNS_40661956134145  M2_M1_CDNS_40661956134145_5
timestamp 1698431365
transform 1 0 7078 0 1 25127
box 0 0 1 1
use M2_M1_CDNS_40661956134146  M2_M1_CDNS_40661956134146_0
timestamp 1698431365
transform 1 0 12185 0 1 12677
box 0 0 1 1
use M2_M1_CDNS_40661956134147  M2_M1_CDNS_40661956134147_0
timestamp 1698431365
transform 1 0 5884 0 1 6805
box 0 0 1 1
use M2_M1_CDNS_40661956134147  M2_M1_CDNS_40661956134147_1
timestamp 1698431365
transform 1 0 5884 0 1 18549
box 0 0 1 1
use M2_M1_CDNS_40661956134147  M2_M1_CDNS_40661956134147_2
timestamp 1698431365
transform 1 0 5884 0 1 12677
box 0 0 1 1
use M2_M1_CDNS_40661956134148  M2_M1_CDNS_40661956134148_0
timestamp 1698431365
transform 1 0 227 0 1 12677
box 0 0 1 1
use nmos_6p0_CDNS_406619561341  nmos_6p0_CDNS_406619561341_0
timestamp 1698431365
transform 0 -1 11481 1 0 13225
box 0 0 1 1
use nmos_6p0_CDNS_406619561341  nmos_6p0_CDNS_406619561341_1
timestamp 1698431365
transform 0 -1 11481 1 0 7353
box 0 0 1 1
use nmos_6p0_CDNS_406619561341  nmos_6p0_CDNS_406619561341_2
timestamp 1698431365
transform 0 -1 11481 1 0 1481
box 0 0 1 1
use nmos_6p0_CDNS_406619561341  nmos_6p0_CDNS_406619561341_3
timestamp 1698431365
transform 0 -1 11481 1 0 19097
box 0 0 1 1
<< properties >>
string GDS_END 4688652
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 4654626
string path 309.200 1.075 309.200 640.425 
<< end >>
