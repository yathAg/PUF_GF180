magic
tech gf180mcuA
magscale 1 10
timestamp 1698431365
use pnp_05p00x00p42_0  pnp_05p00x00p42_0_0
timestamp 1698431365
transform 1 0 400 0 1 840
box -338 -796 338 796
<< labels >>
flabel metal1 s 363 345 363 345 0 FreeSans 200 0 0 0 I1_default_E
port 3 nsew
flabel metal1 s 67 49 67 49 0 FreeSans 200 0 0 0 I1_default_C
port 1 nsew
flabel metal1 s 67 49 67 49 0 FreeSans 200 0 0 0 I1_default_C
port 1 nsew
flabel metal1 s 659 49 659 49 0 FreeSans 200 0 0 0 I1_default_C
port 1 nsew
flabel metal1 s 67 1557 67 1557 0 FreeSans 200 0 0 0 I1_default_C
port 1 nsew
flabel metal1 s 215 197 215 197 0 FreeSans 200 0 0 0 I1_default_B
port 2 nsew
flabel metal1 s 215 197 215 197 0 FreeSans 200 0 0 0 I1_default_B
port 2 nsew
flabel metal1 s 511 197 511 197 0 FreeSans 200 0 0 0 I1_default_B
port 2 nsew
flabel metal1 s 215 1409 215 1409 0 FreeSans 200 0 0 0 I1_default_B
port 2 nsew
<< properties >>
string GDS_END 8168
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_pr/gds/pnp_05p00x00p42.gds
string GDS_START 7474
string device primitive
<< end >>
