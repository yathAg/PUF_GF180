magic
tech gf180mcuA
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 453 2102 1094
<< pwell >>
rect -86 -86 2102 453
<< mvnmos >>
rect 124 69 244 333
rect 348 69 468 333
rect 572 69 692 333
rect 796 69 916 333
rect 1020 69 1140 333
rect 1244 69 1364 333
rect 1468 69 1588 333
rect 1692 69 1812 333
<< mvpmos >>
rect 144 573 244 939
rect 348 573 448 939
rect 582 573 682 939
rect 796 573 896 939
rect 1040 573 1140 939
rect 1254 573 1354 939
rect 1478 573 1578 939
rect 1692 573 1792 939
<< mvndiff >>
rect 36 294 124 333
rect 36 154 49 294
rect 95 154 124 294
rect 36 69 124 154
rect 244 294 348 333
rect 244 154 273 294
rect 319 154 348 294
rect 244 69 348 154
rect 468 314 572 333
rect 468 268 497 314
rect 543 268 572 314
rect 468 69 572 268
rect 692 200 796 333
rect 692 154 721 200
rect 767 154 796 200
rect 692 69 796 154
rect 916 294 1020 333
rect 916 154 945 294
rect 991 154 1020 294
rect 916 69 1020 154
rect 1140 285 1244 333
rect 1140 239 1169 285
rect 1215 239 1244 285
rect 1140 69 1244 239
rect 1364 294 1468 333
rect 1364 154 1393 294
rect 1439 154 1468 294
rect 1364 69 1468 154
rect 1588 285 1692 333
rect 1588 239 1617 285
rect 1663 239 1692 285
rect 1588 69 1692 239
rect 1812 294 1900 333
rect 1812 154 1841 294
rect 1887 154 1900 294
rect 1812 69 1900 154
<< mvpdiff >>
rect 56 923 144 939
rect 56 783 69 923
rect 115 783 144 923
rect 56 573 144 783
rect 244 573 348 939
rect 448 861 582 939
rect 448 721 507 861
rect 553 721 582 861
rect 448 573 582 721
rect 682 573 796 939
rect 896 923 1040 939
rect 896 783 925 923
rect 971 783 1040 923
rect 896 573 1040 783
rect 1140 573 1254 939
rect 1354 861 1478 939
rect 1354 721 1383 861
rect 1429 721 1478 861
rect 1354 573 1478 721
rect 1578 573 1692 939
rect 1792 923 1880 939
rect 1792 783 1821 923
rect 1867 783 1880 923
rect 1792 573 1880 783
<< mvndiffc >>
rect 49 154 95 294
rect 273 154 319 294
rect 497 268 543 314
rect 721 154 767 200
rect 945 154 991 294
rect 1169 239 1215 285
rect 1393 154 1439 294
rect 1617 239 1663 285
rect 1841 154 1887 294
<< mvpdiffc >>
rect 69 783 115 923
rect 507 721 553 861
rect 925 783 971 923
rect 1383 721 1429 861
rect 1821 783 1867 923
<< polysilicon >>
rect 144 939 244 983
rect 348 939 448 983
rect 582 939 682 983
rect 796 939 896 983
rect 1040 939 1140 983
rect 1254 939 1354 983
rect 1478 939 1578 983
rect 1692 939 1792 983
rect 144 500 244 573
rect 144 454 185 500
rect 231 454 244 500
rect 144 377 244 454
rect 124 333 244 377
rect 348 513 448 573
rect 582 513 682 573
rect 348 500 682 513
rect 348 454 361 500
rect 407 454 682 500
rect 348 441 682 454
rect 348 333 468 441
rect 572 377 682 441
rect 796 500 896 573
rect 796 454 809 500
rect 855 454 896 500
rect 796 377 896 454
rect 1040 500 1140 573
rect 1040 454 1081 500
rect 1127 454 1140 500
rect 1040 377 1140 454
rect 1254 513 1354 573
rect 1478 513 1578 573
rect 1254 500 1578 513
rect 1254 454 1267 500
rect 1313 454 1578 500
rect 1254 441 1578 454
rect 1254 377 1364 441
rect 572 333 692 377
rect 796 333 916 377
rect 1020 333 1140 377
rect 1244 333 1364 377
rect 1468 377 1578 441
rect 1692 500 1792 573
rect 1692 454 1705 500
rect 1751 454 1792 500
rect 1692 377 1792 454
rect 1468 333 1588 377
rect 1692 333 1812 377
rect 124 25 244 69
rect 348 25 468 69
rect 572 25 692 69
rect 796 25 916 69
rect 1020 25 1140 69
rect 1244 25 1364 69
rect 1468 25 1588 69
rect 1692 25 1812 69
<< polycontact >>
rect 185 454 231 500
rect 361 454 407 500
rect 809 454 855 500
rect 1081 454 1127 500
rect 1267 454 1313 500
rect 1705 454 1751 500
<< metal1 >>
rect 0 923 2016 1098
rect 0 918 69 923
rect 115 918 925 923
rect 69 772 115 783
rect 507 861 553 872
rect 971 918 1821 923
rect 925 772 971 783
rect 1383 861 1429 872
rect 553 721 1383 726
rect 1867 918 2016 923
rect 1821 772 1867 783
rect 1429 721 1843 726
rect 507 680 1843 721
rect 174 588 866 634
rect 174 500 242 588
rect 174 454 185 500
rect 231 454 242 500
rect 350 500 418 542
rect 350 454 361 500
rect 407 454 418 500
rect 478 500 866 588
rect 478 454 809 500
rect 855 454 866 500
rect 1070 588 1751 634
rect 1070 500 1138 588
rect 1070 454 1081 500
rect 1127 454 1138 500
rect 1256 500 1324 542
rect 1256 454 1267 500
rect 1313 454 1324 500
rect 1374 500 1751 588
rect 1374 454 1705 500
rect 1374 443 1751 454
rect 1797 397 1843 680
rect 49 351 991 397
rect 49 294 95 351
rect 497 314 991 351
rect 49 143 95 154
rect 273 294 319 305
rect 543 294 991 314
rect 543 268 945 294
rect 497 257 945 268
rect 273 90 319 154
rect 721 200 767 211
rect 721 90 767 154
rect 1169 351 1843 397
rect 1169 285 1215 351
rect 1169 228 1215 239
rect 1393 294 1439 305
rect 991 154 1393 182
rect 1598 285 1663 351
rect 1598 239 1617 285
rect 1598 228 1663 239
rect 1841 294 1887 305
rect 1439 154 1841 182
rect 945 136 1887 154
rect 0 -90 2016 90
<< labels >>
flabel metal1 s 1256 454 1324 542 0 FreeSans 200 0 0 0 A1
port 1 nsew default input
flabel metal1 s 1070 588 1751 634 0 FreeSans 200 0 0 0 A2
port 2 nsew default input
flabel metal1 s 350 454 418 542 0 FreeSans 200 0 0 0 B1
port 3 nsew default input
flabel metal1 s 174 588 866 634 0 FreeSans 200 0 0 0 B2
port 4 nsew default input
flabel metal1 s 0 918 2016 1098 0 FreeSans 200 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 273 211 319 305 0 FreeSans 200 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel metal1 s 1383 726 1429 872 0 FreeSans 200 0 0 0 ZN
port 5 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 7 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 8 nsew ground bidirectional
rlabel metal1 s 1374 454 1751 588 1 A2
port 2 nsew default input
rlabel metal1 s 1070 454 1138 588 1 A2
port 2 nsew default input
rlabel metal1 s 1374 443 1751 454 1 A2
port 2 nsew default input
rlabel metal1 s 478 454 866 588 1 B2
port 4 nsew default input
rlabel metal1 s 174 454 242 588 1 B2
port 4 nsew default input
rlabel metal1 s 507 726 553 872 1 ZN
port 5 nsew default output
rlabel metal1 s 507 680 1843 726 1 ZN
port 5 nsew default output
rlabel metal1 s 1797 397 1843 680 1 ZN
port 5 nsew default output
rlabel metal1 s 1169 351 1843 397 1 ZN
port 5 nsew default output
rlabel metal1 s 1598 228 1663 351 1 ZN
port 5 nsew default output
rlabel metal1 s 1169 228 1215 351 1 ZN
port 5 nsew default output
rlabel metal1 s 1821 772 1867 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 925 772 971 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 69 772 115 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 721 90 767 211 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 211 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 2016 90 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2016 1008
string GDS_END 137490
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 132498
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
