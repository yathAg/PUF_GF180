magic
tech gf180mcuB
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 377 3670 870
rect -86 352 2046 377
rect 3170 352 3670 377
<< pwell >>
rect 2046 352 3170 377
rect -86 -86 3670 352
<< mvnmos >>
rect 124 68 244 232
rect 308 68 428 232
rect 532 68 652 232
rect 716 68 836 232
rect 940 68 1060 232
rect 1124 68 1244 232
rect 1348 68 1468 232
rect 1542 68 1662 232
rect 1746 68 1866 232
rect 1940 68 2060 232
rect 2252 68 2372 232
rect 2436 68 2556 232
rect 2660 68 2780 232
rect 2844 68 2964 232
rect 3156 68 3276 232
rect 3340 68 3460 232
<< mvpmos >>
rect 124 547 224 716
rect 328 547 428 716
rect 532 547 632 716
rect 736 547 836 716
rect 940 547 1040 716
rect 1144 547 1244 716
rect 1348 547 1448 716
rect 1552 547 1652 716
rect 1756 547 1856 716
rect 1960 547 2060 716
rect 2252 547 2352 716
rect 2456 547 2556 716
rect 2660 547 2760 716
rect 2864 547 2964 716
rect 3156 547 3256 716
rect 3360 547 3460 716
<< mvndiff >>
rect 2120 244 2192 257
rect 2120 232 2133 244
rect 36 219 124 232
rect 36 173 49 219
rect 95 173 124 219
rect 36 68 124 173
rect 244 68 308 232
rect 428 127 532 232
rect 428 81 457 127
rect 503 81 532 127
rect 428 68 532 81
rect 652 68 716 232
rect 836 190 940 232
rect 836 144 865 190
rect 911 144 940 190
rect 836 68 940 144
rect 1060 68 1124 232
rect 1244 127 1348 232
rect 1244 81 1273 127
rect 1319 81 1348 127
rect 1244 68 1348 81
rect 1468 68 1542 232
rect 1662 68 1746 232
rect 1866 68 1940 232
rect 2060 198 2133 232
rect 2179 232 2192 244
rect 3024 244 3096 257
rect 3024 232 3037 244
rect 2179 198 2252 232
rect 2060 68 2252 198
rect 2372 68 2436 232
rect 2556 152 2660 232
rect 2556 106 2585 152
rect 2631 106 2660 152
rect 2556 68 2660 106
rect 2780 68 2844 232
rect 2964 198 3037 232
rect 3083 232 3096 244
rect 3083 198 3156 232
rect 2964 68 3156 198
rect 3276 68 3340 232
rect 3460 152 3548 232
rect 3460 106 3489 152
rect 3535 106 3548 152
rect 3460 68 3548 106
<< mvpdiff >>
rect 36 654 124 716
rect 36 608 49 654
rect 95 608 124 654
rect 36 547 124 608
rect 224 639 328 716
rect 224 593 253 639
rect 299 593 328 639
rect 224 547 328 593
rect 428 654 532 716
rect 428 608 457 654
rect 503 608 532 654
rect 428 547 532 608
rect 632 639 736 716
rect 632 593 661 639
rect 707 593 736 639
rect 632 547 736 593
rect 836 654 940 716
rect 836 608 865 654
rect 911 608 940 654
rect 836 547 940 608
rect 1040 639 1144 716
rect 1040 593 1069 639
rect 1115 593 1144 639
rect 1040 547 1144 593
rect 1244 654 1348 716
rect 1244 608 1273 654
rect 1319 608 1348 654
rect 1244 547 1348 608
rect 1448 639 1552 716
rect 1448 593 1477 639
rect 1523 593 1552 639
rect 1448 547 1552 593
rect 1652 654 1756 716
rect 1652 608 1681 654
rect 1727 608 1756 654
rect 1652 547 1756 608
rect 1856 639 1960 716
rect 1856 593 1885 639
rect 1931 593 1960 639
rect 1856 547 1960 593
rect 2060 654 2252 716
rect 2060 608 2177 654
rect 2223 608 2252 654
rect 2060 547 2252 608
rect 2352 639 2456 716
rect 2352 593 2381 639
rect 2427 593 2456 639
rect 2352 547 2456 593
rect 2556 654 2660 716
rect 2556 608 2585 654
rect 2631 608 2660 654
rect 2556 547 2660 608
rect 2760 639 2864 716
rect 2760 593 2789 639
rect 2835 593 2864 639
rect 2760 547 2864 593
rect 2964 654 3156 716
rect 2964 608 3081 654
rect 3127 608 3156 654
rect 2964 547 3156 608
rect 3256 639 3360 716
rect 3256 593 3285 639
rect 3331 593 3360 639
rect 3256 547 3360 593
rect 3460 654 3548 716
rect 3460 608 3489 654
rect 3535 608 3548 654
rect 3460 547 3548 608
<< mvndiffc >>
rect 49 173 95 219
rect 457 81 503 127
rect 865 144 911 190
rect 1273 81 1319 127
rect 2133 198 2179 244
rect 2585 106 2631 152
rect 3037 198 3083 244
rect 3489 106 3535 152
<< mvpdiffc >>
rect 49 608 95 654
rect 253 593 299 639
rect 457 608 503 654
rect 661 593 707 639
rect 865 608 911 654
rect 1069 593 1115 639
rect 1273 608 1319 654
rect 1477 593 1523 639
rect 1681 608 1727 654
rect 1885 593 1931 639
rect 2177 608 2223 654
rect 2381 593 2427 639
rect 2585 608 2631 654
rect 2789 593 2835 639
rect 3081 608 3127 654
rect 3285 593 3331 639
rect 3489 608 3535 654
<< polysilicon >>
rect 124 716 224 760
rect 328 716 428 760
rect 532 716 632 760
rect 736 716 836 760
rect 940 716 1040 760
rect 1144 716 1244 760
rect 1348 716 1448 760
rect 1552 716 1652 760
rect 1756 716 1856 760
rect 1960 716 2060 760
rect 2252 716 2352 760
rect 2456 716 2556 760
rect 2660 716 2760 760
rect 2864 716 2964 760
rect 3156 716 3256 760
rect 3360 716 3460 760
rect 124 415 224 547
rect 124 369 153 415
rect 199 369 224 415
rect 124 288 224 369
rect 328 394 428 547
rect 532 394 632 547
rect 328 348 632 394
rect 328 311 428 348
rect 328 288 357 311
rect 124 232 244 288
rect 308 265 357 288
rect 403 265 428 311
rect 308 232 428 265
rect 532 311 632 348
rect 532 265 557 311
rect 603 288 632 311
rect 736 415 836 547
rect 736 369 763 415
rect 809 394 836 415
rect 940 415 1040 547
rect 940 394 966 415
rect 809 369 966 394
rect 1012 369 1040 415
rect 736 348 1040 369
rect 736 288 836 348
rect 603 265 652 288
rect 532 232 652 265
rect 716 232 836 288
rect 940 288 1040 348
rect 1144 394 1244 547
rect 1348 394 1448 547
rect 1144 348 1448 394
rect 1144 311 1244 348
rect 1144 288 1170 311
rect 940 232 1060 288
rect 1124 265 1170 288
rect 1216 265 1244 311
rect 1124 232 1244 265
rect 1348 311 1448 348
rect 1348 265 1371 311
rect 1417 288 1448 311
rect 1552 415 1652 547
rect 1552 369 1577 415
rect 1623 369 1652 415
rect 1552 288 1652 369
rect 1756 428 1856 547
rect 1756 382 1783 428
rect 1829 382 1856 428
rect 1756 288 1856 382
rect 1960 394 2060 547
rect 2252 394 2352 547
rect 1960 348 2352 394
rect 1960 336 2060 348
rect 1960 290 2001 336
rect 2047 290 2060 336
rect 1960 288 2060 290
rect 1417 265 1468 288
rect 1348 232 1468 265
rect 1542 232 1662 288
rect 1746 232 1866 288
rect 1940 232 2060 288
rect 2252 336 2352 348
rect 2252 290 2282 336
rect 2328 290 2352 336
rect 2252 288 2352 290
rect 2456 428 2556 547
rect 2456 382 2482 428
rect 2528 394 2556 428
rect 2660 428 2760 547
rect 2660 394 2692 428
rect 2528 382 2692 394
rect 2738 382 2760 428
rect 2456 348 2760 382
rect 2456 288 2556 348
rect 2252 232 2372 288
rect 2436 232 2556 288
rect 2660 288 2760 348
rect 2864 394 2964 547
rect 3156 394 3256 547
rect 3360 428 3460 547
rect 3360 394 3384 428
rect 2864 348 3256 394
rect 2864 336 2964 348
rect 2864 290 2890 336
rect 2936 290 2964 336
rect 2864 288 2964 290
rect 2660 232 2780 288
rect 2844 232 2964 288
rect 3156 336 3256 348
rect 3156 290 3169 336
rect 3215 290 3256 336
rect 3156 288 3256 290
rect 3340 382 3384 394
rect 3430 382 3460 428
rect 3156 232 3276 288
rect 3340 232 3460 382
rect 124 24 244 68
rect 308 24 428 68
rect 532 24 652 68
rect 716 24 836 68
rect 940 24 1060 68
rect 1124 24 1244 68
rect 1348 24 1468 68
rect 1542 24 1662 68
rect 1746 24 1866 68
rect 1940 24 2060 68
rect 2252 24 2372 68
rect 2436 24 2556 68
rect 2660 24 2780 68
rect 2844 24 2964 68
rect 3156 24 3276 68
rect 3340 24 3460 68
<< polycontact >>
rect 153 369 199 415
rect 357 265 403 311
rect 557 265 603 311
rect 763 369 809 415
rect 966 369 1012 415
rect 1170 265 1216 311
rect 1371 265 1417 311
rect 1577 369 1623 415
rect 1783 382 1829 428
rect 2001 290 2047 336
rect 2282 290 2328 336
rect 2482 382 2528 428
rect 2692 382 2738 428
rect 2890 290 2936 336
rect 3169 290 3215 336
rect 3384 382 3430 428
<< metal1 >>
rect 0 724 3584 844
rect 49 654 95 724
rect 49 568 95 608
rect 253 639 299 662
rect 253 531 299 593
rect 457 654 503 724
rect 457 587 503 608
rect 661 639 707 662
rect 661 531 707 593
rect 865 654 911 724
rect 865 587 911 608
rect 1069 639 1115 662
rect 1069 531 1115 593
rect 1273 654 1319 724
rect 1273 587 1319 608
rect 1477 639 1523 662
rect 1477 531 1523 593
rect 1681 654 1727 724
rect 1681 587 1727 608
rect 1885 639 1931 662
rect 1885 531 1931 593
rect 2177 654 2223 724
rect 2177 587 2223 608
rect 2381 639 2427 662
rect 2381 531 2427 593
rect 2585 654 2631 724
rect 2585 587 2631 608
rect 2789 639 2835 662
rect 2789 531 2835 593
rect 3081 654 3127 724
rect 3081 587 3127 608
rect 3285 639 3331 662
rect 3285 531 3331 593
rect 3489 654 3535 724
rect 3489 587 3535 608
rect 253 476 3555 531
rect 1690 428 3454 430
rect 124 415 1640 419
rect 124 369 153 415
rect 199 369 763 415
rect 809 369 966 415
rect 1012 369 1577 415
rect 1623 369 1640 415
rect 124 365 1640 369
rect 1690 382 1783 428
rect 1829 382 2482 428
rect 2528 382 2692 428
rect 2738 382 3384 428
rect 3430 382 3454 428
rect 1690 365 1894 382
rect 3277 350 3454 382
rect 346 265 357 311
rect 403 265 557 311
rect 603 265 1170 311
rect 1216 265 1371 311
rect 1417 265 1436 311
rect 1990 307 2001 336
rect 1690 290 2001 307
rect 2047 290 2282 336
rect 2328 290 2890 336
rect 2936 290 3169 336
rect 3215 290 3231 336
rect 669 242 1102 265
rect 1690 253 2060 290
rect 3501 244 3555 476
rect 36 173 49 219
rect 95 196 608 219
rect 1168 196 1527 219
rect 2120 198 2133 244
rect 2179 198 3037 244
rect 3083 198 3555 244
rect 95 190 1527 196
rect 95 173 865 190
rect 562 144 865 173
rect 911 173 1527 190
rect 911 144 1214 173
rect 562 138 1214 144
rect 1481 152 1527 173
rect 444 81 457 127
rect 503 81 516 127
rect 444 60 516 81
rect 1260 81 1273 127
rect 1319 81 1332 127
rect 1481 106 2585 152
rect 2631 106 3489 152
rect 3535 106 3546 152
rect 1260 60 1332 81
rect 0 -60 3584 60
<< labels >>
flabel metal1 s 124 365 1640 419 0 FreeSans 400 0 0 0 A3
port 3 nsew default input
flabel metal1 s 346 265 1436 311 0 FreeSans 400 0 0 0 A4
port 4 nsew default input
flabel metal1 s 0 724 3584 844 0 FreeSans 400 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 1260 60 1332 127 0 FreeSans 400 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel metal1 s 3285 531 3331 662 0 FreeSans 400 0 0 0 ZN
port 5 nsew default output
flabel metal1 s 1990 307 3231 336 0 FreeSans 400 0 0 0 A1
port 1 nsew default input
flabel metal1 s 1690 382 3454 430 0 FreeSans 400 0 0 0 A2
port 2 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 7 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 8 nsew ground bidirectional
rlabel metal1 s 1690 290 3231 307 1 A1
port 1 nsew default input
rlabel metal1 s 1690 253 2060 290 1 A1
port 1 nsew default input
rlabel metal1 s 3277 365 3454 382 1 A2
port 2 nsew default input
rlabel metal1 s 1690 365 1894 382 1 A2
port 2 nsew default input
rlabel metal1 s 3277 350 3454 365 1 A2
port 2 nsew default input
rlabel metal1 s 669 242 1102 265 1 A4
port 4 nsew default input
rlabel metal1 s 2789 531 2835 662 1 ZN
port 5 nsew default output
rlabel metal1 s 2381 531 2427 662 1 ZN
port 5 nsew default output
rlabel metal1 s 1885 531 1931 662 1 ZN
port 5 nsew default output
rlabel metal1 s 1477 531 1523 662 1 ZN
port 5 nsew default output
rlabel metal1 s 1069 531 1115 662 1 ZN
port 5 nsew default output
rlabel metal1 s 661 531 707 662 1 ZN
port 5 nsew default output
rlabel metal1 s 253 531 299 662 1 ZN
port 5 nsew default output
rlabel metal1 s 253 476 3555 531 1 ZN
port 5 nsew default output
rlabel metal1 s 3501 244 3555 476 1 ZN
port 5 nsew default output
rlabel metal1 s 2120 198 3555 244 1 ZN
port 5 nsew default output
rlabel metal1 s 3489 587 3535 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3081 587 3127 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2585 587 2631 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2177 587 2223 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1681 587 1727 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1273 587 1319 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 865 587 911 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 457 587 503 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 49 587 95 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 49 568 95 587 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 444 60 516 127 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3584 60 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3584 784
string GDS_END 737418
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 730492
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
