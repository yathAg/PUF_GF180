magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 453 1318 1094
<< pwell >>
rect -86 -86 1318 453
<< metal1 >>
rect 0 918 1232 1098
rect 264 775 310 918
rect 672 775 718 918
rect 1116 775 1162 918
rect 23 430 194 542
rect 242 430 418 542
rect 478 458 642 542
rect 672 90 718 233
rect 896 169 978 737
rect 1120 90 1166 233
rect 0 -90 1232 90
<< obsm1 >>
rect 468 706 514 822
rect 49 660 842 706
rect 796 384 842 660
rect 60 338 842 384
rect 60 169 106 338
<< labels >>
rlabel metal1 s 23 430 194 542 6 A1
port 1 nsew default input
rlabel metal1 s 242 430 418 542 6 A2
port 2 nsew default input
rlabel metal1 s 478 458 642 542 6 A3
port 3 nsew default input
rlabel metal1 s 896 169 978 737 6 Z
port 4 nsew default output
rlabel metal1 s 1116 775 1162 918 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 672 775 718 918 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 264 775 310 918 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 918 1232 1098 6 VDD
port 5 nsew power bidirectional abutment
rlabel nwell s -86 453 1318 1094 6 VNW
port 6 nsew power bidirectional
rlabel pwell s -86 -86 1318 453 6 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 0 -90 1232 90 8 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1120 90 1166 233 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 672 90 718 233 6 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1232 1008
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1144468
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1140418
<< end >>
