magic
tech gf180mcuD
magscale 1 10
timestamp 1698431365
<< metal1 >>
rect 2203 55545 88011 55557
rect 2203 55493 27130 55545
rect 27182 55493 27254 55545
rect 27306 55493 27378 55545
rect 27430 55493 27502 55545
rect 27554 55493 27626 55545
rect 27678 55493 27750 55545
rect 27802 55493 27874 55545
rect 27926 55493 27998 55545
rect 28050 55493 35986 55545
rect 36038 55493 36110 55545
rect 36162 55493 36234 55545
rect 36286 55493 36358 55545
rect 36410 55493 36482 55545
rect 36534 55493 36606 55545
rect 36658 55493 36730 55545
rect 36782 55493 36854 55545
rect 36906 55493 41828 55545
rect 41880 55493 41952 55545
rect 42004 55493 42076 55545
rect 42128 55493 42200 55545
rect 42252 55493 42324 55545
rect 42376 55493 42448 55545
rect 42500 55493 42572 55545
rect 42624 55493 42696 55545
rect 42748 55493 45659 55545
rect 45711 55493 45783 55545
rect 45835 55493 45907 55545
rect 45959 55493 46031 55545
rect 46083 55493 46155 55545
rect 46207 55493 46279 55545
rect 46331 55493 46403 55545
rect 46455 55493 46527 55545
rect 46579 55493 52411 55545
rect 52463 55493 52535 55545
rect 52587 55493 52659 55545
rect 52711 55493 52783 55545
rect 52835 55493 52907 55545
rect 52959 55493 53031 55545
rect 53083 55493 53155 55545
rect 53207 55493 53279 55545
rect 53331 55493 57936 55545
rect 57988 55493 58060 55545
rect 58112 55493 58184 55545
rect 58236 55493 58308 55545
rect 58360 55493 58432 55545
rect 58484 55493 58556 55545
rect 58608 55493 58680 55545
rect 58732 55493 58804 55545
rect 58856 55493 60737 55545
rect 60789 55493 60861 55545
rect 60913 55493 60985 55545
rect 61037 55493 61109 55545
rect 61161 55493 61233 55545
rect 61285 55493 61357 55545
rect 61409 55493 61481 55545
rect 61533 55493 61605 55545
rect 61657 55493 88011 55545
rect 2203 55421 88011 55493
rect 2203 55369 27130 55421
rect 27182 55369 27254 55421
rect 27306 55369 27378 55421
rect 27430 55369 27502 55421
rect 27554 55369 27626 55421
rect 27678 55369 27750 55421
rect 27802 55369 27874 55421
rect 27926 55369 27998 55421
rect 28050 55369 35986 55421
rect 36038 55369 36110 55421
rect 36162 55369 36234 55421
rect 36286 55369 36358 55421
rect 36410 55369 36482 55421
rect 36534 55369 36606 55421
rect 36658 55369 36730 55421
rect 36782 55369 36854 55421
rect 36906 55369 41828 55421
rect 41880 55369 41952 55421
rect 42004 55369 42076 55421
rect 42128 55369 42200 55421
rect 42252 55369 42324 55421
rect 42376 55369 42448 55421
rect 42500 55369 42572 55421
rect 42624 55369 42696 55421
rect 42748 55369 45659 55421
rect 45711 55369 45783 55421
rect 45835 55369 45907 55421
rect 45959 55369 46031 55421
rect 46083 55369 46155 55421
rect 46207 55369 46279 55421
rect 46331 55369 46403 55421
rect 46455 55369 46527 55421
rect 46579 55369 52411 55421
rect 52463 55369 52535 55421
rect 52587 55369 52659 55421
rect 52711 55369 52783 55421
rect 52835 55369 52907 55421
rect 52959 55369 53031 55421
rect 53083 55369 53155 55421
rect 53207 55369 53279 55421
rect 53331 55369 57936 55421
rect 57988 55369 58060 55421
rect 58112 55369 58184 55421
rect 58236 55369 58308 55421
rect 58360 55369 58432 55421
rect 58484 55369 58556 55421
rect 58608 55369 58680 55421
rect 58732 55369 58804 55421
rect 58856 55369 60737 55421
rect 60789 55369 60861 55421
rect 60913 55369 60985 55421
rect 61037 55369 61109 55421
rect 61161 55369 61233 55421
rect 61285 55369 61357 55421
rect 61409 55369 61481 55421
rect 61533 55369 61605 55421
rect 61657 55369 88011 55421
rect 2203 55297 88011 55369
rect 2203 55245 27130 55297
rect 27182 55245 27254 55297
rect 27306 55245 27378 55297
rect 27430 55245 27502 55297
rect 27554 55245 27626 55297
rect 27678 55245 27750 55297
rect 27802 55245 27874 55297
rect 27926 55245 27998 55297
rect 28050 55245 35986 55297
rect 36038 55245 36110 55297
rect 36162 55245 36234 55297
rect 36286 55245 36358 55297
rect 36410 55245 36482 55297
rect 36534 55245 36606 55297
rect 36658 55245 36730 55297
rect 36782 55245 36854 55297
rect 36906 55245 41828 55297
rect 41880 55245 41952 55297
rect 42004 55245 42076 55297
rect 42128 55245 42200 55297
rect 42252 55245 42324 55297
rect 42376 55245 42448 55297
rect 42500 55245 42572 55297
rect 42624 55245 42696 55297
rect 42748 55245 45659 55297
rect 45711 55245 45783 55297
rect 45835 55245 45907 55297
rect 45959 55245 46031 55297
rect 46083 55245 46155 55297
rect 46207 55245 46279 55297
rect 46331 55245 46403 55297
rect 46455 55245 46527 55297
rect 46579 55245 52411 55297
rect 52463 55245 52535 55297
rect 52587 55245 52659 55297
rect 52711 55245 52783 55297
rect 52835 55245 52907 55297
rect 52959 55245 53031 55297
rect 53083 55245 53155 55297
rect 53207 55245 53279 55297
rect 53331 55245 57936 55297
rect 57988 55245 58060 55297
rect 58112 55245 58184 55297
rect 58236 55245 58308 55297
rect 58360 55245 58432 55297
rect 58484 55245 58556 55297
rect 58608 55245 58680 55297
rect 58732 55245 58804 55297
rect 58856 55245 60737 55297
rect 60789 55245 60861 55297
rect 60913 55245 60985 55297
rect 61037 55245 61109 55297
rect 61161 55245 61233 55297
rect 61285 55245 61357 55297
rect 61409 55245 61481 55297
rect 61533 55245 61605 55297
rect 61657 55245 88011 55297
rect 2203 54557 88011 55245
rect 35945 53519 36945 54557
rect 42135 53477 42444 54557
rect 45745 53475 46606 54557
rect 59270 4787 59594 4799
rect 59270 4735 59282 4787
rect 59334 4735 59406 4787
rect 59458 4735 59530 4787
rect 59582 4735 59594 4787
rect 59270 4663 59594 4735
rect 59270 4611 59282 4663
rect 59334 4611 59406 4663
rect 59458 4611 59530 4663
rect 59582 4611 59594 4663
rect 59270 4539 59594 4611
rect 59270 4487 59282 4539
rect 59334 4487 59406 4539
rect 59458 4487 59530 4539
rect 59582 4487 59594 4539
rect 59270 4415 59594 4487
rect 59270 4363 59282 4415
rect 59334 4363 59406 4415
rect 59458 4363 59530 4415
rect 59582 4363 59594 4415
rect 28753 4280 29077 4292
rect 59270 4291 59594 4363
rect 28753 4228 28765 4280
rect 28817 4228 28889 4280
rect 28941 4228 29013 4280
rect 29065 4228 29077 4280
rect 28753 4156 29077 4228
rect 28753 4104 28765 4156
rect 28817 4104 28889 4156
rect 28941 4104 29013 4156
rect 29065 4104 29077 4156
rect 28753 4032 29077 4104
rect 28753 3980 28765 4032
rect 28817 3980 28889 4032
rect 28941 3980 29013 4032
rect 29065 3980 29077 4032
rect 28753 3908 29077 3980
rect 28753 3856 28765 3908
rect 28817 3856 28889 3908
rect 28941 3856 29013 3908
rect 29065 3856 29077 3908
rect 28753 3844 29077 3856
rect 29362 4273 29686 4285
rect 29362 4221 29374 4273
rect 29426 4221 29498 4273
rect 29550 4221 29622 4273
rect 29674 4221 29686 4273
rect 29362 4149 29686 4221
rect 29362 4097 29374 4149
rect 29426 4097 29498 4149
rect 29550 4097 29622 4149
rect 29674 4097 29686 4149
rect 29362 4025 29686 4097
rect 29362 3973 29374 4025
rect 29426 3973 29498 4025
rect 29550 3973 29622 4025
rect 29674 3973 29686 4025
rect 29362 3901 29686 3973
rect 29362 3849 29374 3901
rect 29426 3849 29498 3901
rect 29550 3849 29622 3901
rect 29674 3849 29686 3901
rect 29362 3777 29686 3849
rect 29362 3725 29374 3777
rect 29426 3725 29498 3777
rect 29550 3725 29622 3777
rect 29674 3725 29686 3777
rect 29362 3653 29686 3725
rect 29362 3601 29374 3653
rect 29426 3601 29498 3653
rect 29550 3601 29622 3653
rect 29674 3601 29686 3653
rect 29362 3529 29686 3601
rect 29362 3477 29374 3529
rect 29426 3477 29498 3529
rect 29550 3477 29622 3529
rect 29674 3477 29686 3529
rect 29362 3405 29686 3477
rect 29362 3353 29374 3405
rect 29426 3353 29498 3405
rect 29550 3353 29622 3405
rect 29674 3353 29686 3405
rect 29362 3345 29686 3353
rect 59270 4239 59282 4291
rect 59334 4239 59406 4291
rect 59458 4239 59530 4291
rect 59582 4239 59594 4291
rect 59270 4167 59594 4239
rect 59270 4115 59282 4167
rect 59334 4115 59406 4167
rect 59458 4115 59530 4167
rect 59582 4115 59594 4167
rect 59270 4043 59594 4115
rect 59270 3991 59282 4043
rect 59334 3991 59406 4043
rect 59458 3991 59530 4043
rect 59582 3991 59594 4043
rect 59270 3919 59594 3991
rect 59270 3867 59282 3919
rect 59334 3867 59406 3919
rect 59458 3867 59530 3919
rect 59582 3867 59594 3919
rect 59270 3795 59594 3867
rect 59890 4280 60214 4292
rect 59890 4228 59902 4280
rect 59954 4228 60026 4280
rect 60078 4228 60150 4280
rect 60202 4228 60214 4280
rect 59890 4156 60214 4228
rect 59890 4104 59902 4156
rect 59954 4104 60026 4156
rect 60078 4104 60150 4156
rect 60202 4104 60214 4156
rect 59890 4032 60214 4104
rect 59890 3980 59902 4032
rect 59954 3980 60026 4032
rect 60078 3980 60150 4032
rect 60202 3980 60214 4032
rect 59890 3908 60214 3980
rect 59890 3856 59902 3908
rect 59954 3856 60026 3908
rect 60078 3856 60150 3908
rect 60202 3856 60214 3908
rect 59890 3844 60214 3856
rect 59270 3743 59282 3795
rect 59334 3743 59406 3795
rect 59458 3743 59530 3795
rect 59582 3743 59594 3795
rect 59270 3671 59594 3743
rect 59270 3619 59282 3671
rect 59334 3619 59406 3671
rect 59458 3619 59530 3671
rect 59582 3619 59594 3671
rect 59270 3547 59594 3619
rect 59270 3495 59282 3547
rect 59334 3495 59406 3547
rect 59458 3495 59530 3547
rect 59582 3495 59594 3547
rect 59270 3423 59594 3495
rect 59270 3371 59282 3423
rect 59334 3371 59406 3423
rect 59458 3371 59530 3423
rect 59582 3371 59594 3423
rect 59270 3345 59594 3371
rect 87011 3345 88011 54557
rect 2203 3299 88011 3345
rect 2203 3281 59282 3299
rect 2203 3229 29374 3281
rect 29426 3229 29498 3281
rect 29550 3229 29622 3281
rect 29674 3247 59282 3281
rect 59334 3247 59406 3299
rect 59458 3247 59530 3299
rect 59582 3247 88011 3299
rect 29674 3229 88011 3247
rect 2203 3175 88011 3229
rect 2203 3157 59282 3175
rect 2203 3105 29374 3157
rect 29426 3105 29498 3157
rect 29550 3105 29622 3157
rect 29674 3123 59282 3157
rect 59334 3123 59406 3175
rect 59458 3123 59530 3175
rect 59582 3123 88011 3175
rect 29674 3105 88011 3123
rect 2203 3051 88011 3105
rect 2203 3033 59282 3051
rect 2203 2981 29374 3033
rect 29426 2981 29498 3033
rect 29550 2981 29622 3033
rect 29674 2999 59282 3033
rect 59334 2999 59406 3051
rect 59458 2999 59530 3051
rect 59582 2999 88011 3051
rect 29674 2981 88011 2999
rect 2203 2927 88011 2981
rect 2203 2909 59282 2927
rect 2203 2857 29374 2909
rect 29426 2857 29498 2909
rect 29550 2857 29622 2909
rect 29674 2875 59282 2909
rect 59334 2875 59406 2927
rect 59458 2875 59530 2927
rect 59582 2875 88011 2927
rect 29674 2857 88011 2875
rect 2203 2803 88011 2857
rect 2203 2785 59282 2803
rect 2203 2733 29374 2785
rect 29426 2733 29498 2785
rect 29550 2733 29622 2785
rect 29674 2751 59282 2785
rect 59334 2751 59406 2803
rect 59458 2751 59530 2803
rect 59582 2751 88011 2803
rect 29674 2733 88011 2751
rect 2203 2679 88011 2733
rect 2203 2661 59282 2679
rect 2203 2609 29374 2661
rect 29426 2609 29498 2661
rect 29550 2609 29622 2661
rect 29674 2627 59282 2661
rect 59334 2627 59406 2679
rect 59458 2627 59530 2679
rect 59582 2627 88011 2679
rect 29674 2609 88011 2627
rect 2203 2555 88011 2609
rect 2203 2537 59282 2555
rect 2203 2485 29374 2537
rect 29426 2485 29498 2537
rect 29550 2485 29622 2537
rect 29674 2503 59282 2537
rect 59334 2503 59406 2555
rect 59458 2503 59530 2555
rect 59582 2503 88011 2555
rect 29674 2485 88011 2503
rect 2203 2431 88011 2485
rect 2203 2413 59282 2431
rect 2203 2361 29374 2413
rect 29426 2361 29498 2413
rect 29550 2361 29622 2413
rect 29674 2379 59282 2413
rect 59334 2379 59406 2431
rect 59458 2379 59530 2431
rect 59582 2379 88011 2431
rect 29674 2361 88011 2379
rect 2203 2345 88011 2361
<< via1 >>
rect 27130 55493 27182 55545
rect 27254 55493 27306 55545
rect 27378 55493 27430 55545
rect 27502 55493 27554 55545
rect 27626 55493 27678 55545
rect 27750 55493 27802 55545
rect 27874 55493 27926 55545
rect 27998 55493 28050 55545
rect 35986 55493 36038 55545
rect 36110 55493 36162 55545
rect 36234 55493 36286 55545
rect 36358 55493 36410 55545
rect 36482 55493 36534 55545
rect 36606 55493 36658 55545
rect 36730 55493 36782 55545
rect 36854 55493 36906 55545
rect 41828 55493 41880 55545
rect 41952 55493 42004 55545
rect 42076 55493 42128 55545
rect 42200 55493 42252 55545
rect 42324 55493 42376 55545
rect 42448 55493 42500 55545
rect 42572 55493 42624 55545
rect 42696 55493 42748 55545
rect 45659 55493 45711 55545
rect 45783 55493 45835 55545
rect 45907 55493 45959 55545
rect 46031 55493 46083 55545
rect 46155 55493 46207 55545
rect 46279 55493 46331 55545
rect 46403 55493 46455 55545
rect 46527 55493 46579 55545
rect 52411 55493 52463 55545
rect 52535 55493 52587 55545
rect 52659 55493 52711 55545
rect 52783 55493 52835 55545
rect 52907 55493 52959 55545
rect 53031 55493 53083 55545
rect 53155 55493 53207 55545
rect 53279 55493 53331 55545
rect 57936 55493 57988 55545
rect 58060 55493 58112 55545
rect 58184 55493 58236 55545
rect 58308 55493 58360 55545
rect 58432 55493 58484 55545
rect 58556 55493 58608 55545
rect 58680 55493 58732 55545
rect 58804 55493 58856 55545
rect 60737 55493 60789 55545
rect 60861 55493 60913 55545
rect 60985 55493 61037 55545
rect 61109 55493 61161 55545
rect 61233 55493 61285 55545
rect 61357 55493 61409 55545
rect 61481 55493 61533 55545
rect 61605 55493 61657 55545
rect 27130 55369 27182 55421
rect 27254 55369 27306 55421
rect 27378 55369 27430 55421
rect 27502 55369 27554 55421
rect 27626 55369 27678 55421
rect 27750 55369 27802 55421
rect 27874 55369 27926 55421
rect 27998 55369 28050 55421
rect 35986 55369 36038 55421
rect 36110 55369 36162 55421
rect 36234 55369 36286 55421
rect 36358 55369 36410 55421
rect 36482 55369 36534 55421
rect 36606 55369 36658 55421
rect 36730 55369 36782 55421
rect 36854 55369 36906 55421
rect 41828 55369 41880 55421
rect 41952 55369 42004 55421
rect 42076 55369 42128 55421
rect 42200 55369 42252 55421
rect 42324 55369 42376 55421
rect 42448 55369 42500 55421
rect 42572 55369 42624 55421
rect 42696 55369 42748 55421
rect 45659 55369 45711 55421
rect 45783 55369 45835 55421
rect 45907 55369 45959 55421
rect 46031 55369 46083 55421
rect 46155 55369 46207 55421
rect 46279 55369 46331 55421
rect 46403 55369 46455 55421
rect 46527 55369 46579 55421
rect 52411 55369 52463 55421
rect 52535 55369 52587 55421
rect 52659 55369 52711 55421
rect 52783 55369 52835 55421
rect 52907 55369 52959 55421
rect 53031 55369 53083 55421
rect 53155 55369 53207 55421
rect 53279 55369 53331 55421
rect 57936 55369 57988 55421
rect 58060 55369 58112 55421
rect 58184 55369 58236 55421
rect 58308 55369 58360 55421
rect 58432 55369 58484 55421
rect 58556 55369 58608 55421
rect 58680 55369 58732 55421
rect 58804 55369 58856 55421
rect 60737 55369 60789 55421
rect 60861 55369 60913 55421
rect 60985 55369 61037 55421
rect 61109 55369 61161 55421
rect 61233 55369 61285 55421
rect 61357 55369 61409 55421
rect 61481 55369 61533 55421
rect 61605 55369 61657 55421
rect 27130 55245 27182 55297
rect 27254 55245 27306 55297
rect 27378 55245 27430 55297
rect 27502 55245 27554 55297
rect 27626 55245 27678 55297
rect 27750 55245 27802 55297
rect 27874 55245 27926 55297
rect 27998 55245 28050 55297
rect 35986 55245 36038 55297
rect 36110 55245 36162 55297
rect 36234 55245 36286 55297
rect 36358 55245 36410 55297
rect 36482 55245 36534 55297
rect 36606 55245 36658 55297
rect 36730 55245 36782 55297
rect 36854 55245 36906 55297
rect 41828 55245 41880 55297
rect 41952 55245 42004 55297
rect 42076 55245 42128 55297
rect 42200 55245 42252 55297
rect 42324 55245 42376 55297
rect 42448 55245 42500 55297
rect 42572 55245 42624 55297
rect 42696 55245 42748 55297
rect 45659 55245 45711 55297
rect 45783 55245 45835 55297
rect 45907 55245 45959 55297
rect 46031 55245 46083 55297
rect 46155 55245 46207 55297
rect 46279 55245 46331 55297
rect 46403 55245 46455 55297
rect 46527 55245 46579 55297
rect 52411 55245 52463 55297
rect 52535 55245 52587 55297
rect 52659 55245 52711 55297
rect 52783 55245 52835 55297
rect 52907 55245 52959 55297
rect 53031 55245 53083 55297
rect 53155 55245 53207 55297
rect 53279 55245 53331 55297
rect 57936 55245 57988 55297
rect 58060 55245 58112 55297
rect 58184 55245 58236 55297
rect 58308 55245 58360 55297
rect 58432 55245 58484 55297
rect 58556 55245 58608 55297
rect 58680 55245 58732 55297
rect 58804 55245 58856 55297
rect 60737 55245 60789 55297
rect 60861 55245 60913 55297
rect 60985 55245 61037 55297
rect 61109 55245 61161 55297
rect 61233 55245 61285 55297
rect 61357 55245 61409 55297
rect 61481 55245 61533 55297
rect 61605 55245 61657 55297
rect 59282 4735 59334 4787
rect 59406 4735 59458 4787
rect 59530 4735 59582 4787
rect 59282 4611 59334 4663
rect 59406 4611 59458 4663
rect 59530 4611 59582 4663
rect 59282 4487 59334 4539
rect 59406 4487 59458 4539
rect 59530 4487 59582 4539
rect 59282 4363 59334 4415
rect 59406 4363 59458 4415
rect 59530 4363 59582 4415
rect 28765 4228 28817 4280
rect 28889 4228 28941 4280
rect 29013 4228 29065 4280
rect 28765 4104 28817 4156
rect 28889 4104 28941 4156
rect 29013 4104 29065 4156
rect 28765 3980 28817 4032
rect 28889 3980 28941 4032
rect 29013 3980 29065 4032
rect 28765 3856 28817 3908
rect 28889 3856 28941 3908
rect 29013 3856 29065 3908
rect 29374 4221 29426 4273
rect 29498 4221 29550 4273
rect 29622 4221 29674 4273
rect 29374 4097 29426 4149
rect 29498 4097 29550 4149
rect 29622 4097 29674 4149
rect 29374 3973 29426 4025
rect 29498 3973 29550 4025
rect 29622 3973 29674 4025
rect 29374 3849 29426 3901
rect 29498 3849 29550 3901
rect 29622 3849 29674 3901
rect 29374 3725 29426 3777
rect 29498 3725 29550 3777
rect 29622 3725 29674 3777
rect 29374 3601 29426 3653
rect 29498 3601 29550 3653
rect 29622 3601 29674 3653
rect 29374 3477 29426 3529
rect 29498 3477 29550 3529
rect 29622 3477 29674 3529
rect 29374 3353 29426 3405
rect 29498 3353 29550 3405
rect 29622 3353 29674 3405
rect 59282 4239 59334 4291
rect 59406 4239 59458 4291
rect 59530 4239 59582 4291
rect 59282 4115 59334 4167
rect 59406 4115 59458 4167
rect 59530 4115 59582 4167
rect 59282 3991 59334 4043
rect 59406 3991 59458 4043
rect 59530 3991 59582 4043
rect 59282 3867 59334 3919
rect 59406 3867 59458 3919
rect 59530 3867 59582 3919
rect 59902 4228 59954 4280
rect 60026 4228 60078 4280
rect 60150 4228 60202 4280
rect 59902 4104 59954 4156
rect 60026 4104 60078 4156
rect 60150 4104 60202 4156
rect 59902 3980 59954 4032
rect 60026 3980 60078 4032
rect 60150 3980 60202 4032
rect 59902 3856 59954 3908
rect 60026 3856 60078 3908
rect 60150 3856 60202 3908
rect 59282 3743 59334 3795
rect 59406 3743 59458 3795
rect 59530 3743 59582 3795
rect 59282 3619 59334 3671
rect 59406 3619 59458 3671
rect 59530 3619 59582 3671
rect 59282 3495 59334 3547
rect 59406 3495 59458 3547
rect 59530 3495 59582 3547
rect 59282 3371 59334 3423
rect 59406 3371 59458 3423
rect 59530 3371 59582 3423
rect 29374 3229 29426 3281
rect 29498 3229 29550 3281
rect 29622 3229 29674 3281
rect 59282 3247 59334 3299
rect 59406 3247 59458 3299
rect 59530 3247 59582 3299
rect 29374 3105 29426 3157
rect 29498 3105 29550 3157
rect 29622 3105 29674 3157
rect 59282 3123 59334 3175
rect 59406 3123 59458 3175
rect 59530 3123 59582 3175
rect 29374 2981 29426 3033
rect 29498 2981 29550 3033
rect 29622 2981 29674 3033
rect 59282 2999 59334 3051
rect 59406 2999 59458 3051
rect 59530 2999 59582 3051
rect 29374 2857 29426 2909
rect 29498 2857 29550 2909
rect 29622 2857 29674 2909
rect 59282 2875 59334 2927
rect 59406 2875 59458 2927
rect 59530 2875 59582 2927
rect 29374 2733 29426 2785
rect 29498 2733 29550 2785
rect 29622 2733 29674 2785
rect 59282 2751 59334 2803
rect 59406 2751 59458 2803
rect 59530 2751 59582 2803
rect 29374 2609 29426 2661
rect 29498 2609 29550 2661
rect 29622 2609 29674 2661
rect 59282 2627 59334 2679
rect 59406 2627 59458 2679
rect 59530 2627 59582 2679
rect 29374 2485 29426 2537
rect 29498 2485 29550 2537
rect 29622 2485 29674 2537
rect 59282 2503 59334 2555
rect 59406 2503 59458 2555
rect 59530 2503 59582 2555
rect 29374 2361 29426 2413
rect 29498 2361 29550 2413
rect 29622 2361 29674 2413
rect 59282 2379 59334 2431
rect 59406 2379 59458 2431
rect 59530 2379 59582 2431
<< metal2 >>
rect 27118 55547 28062 55557
rect 27118 55491 27128 55547
rect 27184 55491 27252 55547
rect 27308 55491 27376 55547
rect 27432 55491 27500 55547
rect 27556 55491 27624 55547
rect 27680 55491 27748 55547
rect 27804 55491 27872 55547
rect 27928 55491 27996 55547
rect 28052 55491 28062 55547
rect 27118 55423 28062 55491
rect 27118 55367 27128 55423
rect 27184 55367 27252 55423
rect 27308 55367 27376 55423
rect 27432 55367 27500 55423
rect 27556 55367 27624 55423
rect 27680 55367 27748 55423
rect 27804 55367 27872 55423
rect 27928 55367 27996 55423
rect 28052 55367 28062 55423
rect 27118 55299 28062 55367
rect 27118 55243 27128 55299
rect 27184 55243 27252 55299
rect 27308 55243 27376 55299
rect 27432 55243 27500 55299
rect 27556 55243 27624 55299
rect 27680 55243 27748 55299
rect 27804 55243 27872 55299
rect 27928 55243 27996 55299
rect 28052 55243 28062 55299
rect 27118 55233 28062 55243
rect 35974 55547 36918 55557
rect 35974 55491 35984 55547
rect 36040 55491 36108 55547
rect 36164 55491 36232 55547
rect 36288 55491 36356 55547
rect 36412 55491 36480 55547
rect 36536 55491 36604 55547
rect 36660 55491 36728 55547
rect 36784 55491 36852 55547
rect 36908 55491 36918 55547
rect 35974 55423 36918 55491
rect 35974 55367 35984 55423
rect 36040 55367 36108 55423
rect 36164 55367 36232 55423
rect 36288 55367 36356 55423
rect 36412 55367 36480 55423
rect 36536 55367 36604 55423
rect 36660 55367 36728 55423
rect 36784 55367 36852 55423
rect 36908 55367 36918 55423
rect 35974 55299 36918 55367
rect 35974 55243 35984 55299
rect 36040 55243 36108 55299
rect 36164 55243 36232 55299
rect 36288 55243 36356 55299
rect 36412 55243 36480 55299
rect 36536 55243 36604 55299
rect 36660 55243 36728 55299
rect 36784 55243 36852 55299
rect 36908 55243 36918 55299
rect 35974 55233 36918 55243
rect 41816 55547 42760 55557
rect 41816 55491 41826 55547
rect 41882 55491 41950 55547
rect 42006 55491 42074 55547
rect 42130 55491 42198 55547
rect 42254 55491 42322 55547
rect 42378 55491 42446 55547
rect 42502 55491 42570 55547
rect 42626 55491 42694 55547
rect 42750 55491 42760 55547
rect 41816 55423 42760 55491
rect 41816 55367 41826 55423
rect 41882 55367 41950 55423
rect 42006 55367 42074 55423
rect 42130 55367 42198 55423
rect 42254 55367 42322 55423
rect 42378 55367 42446 55423
rect 42502 55367 42570 55423
rect 42626 55367 42694 55423
rect 42750 55367 42760 55423
rect 41816 55299 42760 55367
rect 41816 55243 41826 55299
rect 41882 55243 41950 55299
rect 42006 55243 42074 55299
rect 42130 55243 42198 55299
rect 42254 55243 42322 55299
rect 42378 55243 42446 55299
rect 42502 55243 42570 55299
rect 42626 55243 42694 55299
rect 42750 55243 42760 55299
rect 41816 55233 42760 55243
rect 45647 55547 46591 55557
rect 45647 55491 45657 55547
rect 45713 55491 45781 55547
rect 45837 55491 45905 55547
rect 45961 55491 46029 55547
rect 46085 55491 46153 55547
rect 46209 55491 46277 55547
rect 46333 55491 46401 55547
rect 46457 55491 46525 55547
rect 46581 55491 46591 55547
rect 45647 55423 46591 55491
rect 45647 55367 45657 55423
rect 45713 55367 45781 55423
rect 45837 55367 45905 55423
rect 45961 55367 46029 55423
rect 46085 55367 46153 55423
rect 46209 55367 46277 55423
rect 46333 55367 46401 55423
rect 46457 55367 46525 55423
rect 46581 55367 46591 55423
rect 45647 55299 46591 55367
rect 45647 55243 45657 55299
rect 45713 55243 45781 55299
rect 45837 55243 45905 55299
rect 45961 55243 46029 55299
rect 46085 55243 46153 55299
rect 46209 55243 46277 55299
rect 46333 55243 46401 55299
rect 46457 55243 46525 55299
rect 46581 55243 46591 55299
rect 45647 55233 46591 55243
rect 52399 55547 53343 55557
rect 52399 55491 52409 55547
rect 52465 55491 52533 55547
rect 52589 55491 52657 55547
rect 52713 55491 52781 55547
rect 52837 55491 52905 55547
rect 52961 55491 53029 55547
rect 53085 55491 53153 55547
rect 53209 55491 53277 55547
rect 53333 55491 53343 55547
rect 52399 55423 53343 55491
rect 52399 55367 52409 55423
rect 52465 55367 52533 55423
rect 52589 55367 52657 55423
rect 52713 55367 52781 55423
rect 52837 55367 52905 55423
rect 52961 55367 53029 55423
rect 53085 55367 53153 55423
rect 53209 55367 53277 55423
rect 53333 55367 53343 55423
rect 52399 55299 53343 55367
rect 52399 55243 52409 55299
rect 52465 55243 52533 55299
rect 52589 55243 52657 55299
rect 52713 55243 52781 55299
rect 52837 55243 52905 55299
rect 52961 55243 53029 55299
rect 53085 55243 53153 55299
rect 53209 55243 53277 55299
rect 53333 55243 53343 55299
rect 52399 55233 53343 55243
rect 57924 55547 58868 55557
rect 57924 55491 57934 55547
rect 57990 55491 58058 55547
rect 58114 55491 58182 55547
rect 58238 55491 58306 55547
rect 58362 55491 58430 55547
rect 58486 55491 58554 55547
rect 58610 55491 58678 55547
rect 58734 55491 58802 55547
rect 58858 55491 58868 55547
rect 57924 55423 58868 55491
rect 57924 55367 57934 55423
rect 57990 55367 58058 55423
rect 58114 55367 58182 55423
rect 58238 55367 58306 55423
rect 58362 55367 58430 55423
rect 58486 55367 58554 55423
rect 58610 55367 58678 55423
rect 58734 55367 58802 55423
rect 58858 55367 58868 55423
rect 57924 55299 58868 55367
rect 57924 55243 57934 55299
rect 57990 55243 58058 55299
rect 58114 55243 58182 55299
rect 58238 55243 58306 55299
rect 58362 55243 58430 55299
rect 58486 55243 58554 55299
rect 58610 55243 58678 55299
rect 58734 55243 58802 55299
rect 58858 55243 58868 55299
rect 57924 55233 58868 55243
rect 60725 55547 61669 55557
rect 60725 55491 60735 55547
rect 60791 55491 60859 55547
rect 60915 55491 60983 55547
rect 61039 55491 61107 55547
rect 61163 55491 61231 55547
rect 61287 55491 61355 55547
rect 61411 55491 61479 55547
rect 61535 55491 61603 55547
rect 61659 55491 61669 55547
rect 60725 55423 61669 55491
rect 60725 55367 60735 55423
rect 60791 55367 60859 55423
rect 60915 55367 60983 55423
rect 61039 55367 61107 55423
rect 61163 55367 61231 55423
rect 61287 55367 61355 55423
rect 61411 55367 61479 55423
rect 61535 55367 61603 55423
rect 61659 55367 61669 55423
rect 60725 55299 61669 55367
rect 60725 55243 60735 55299
rect 60791 55243 60859 55299
rect 60915 55243 60983 55299
rect 61039 55243 61107 55299
rect 61163 55243 61231 55299
rect 61287 55243 61355 55299
rect 61411 55243 61479 55299
rect 61535 55243 61603 55299
rect 61659 55243 61669 55299
rect 60725 55233 61669 55243
rect 28523 54998 29467 55008
rect 28523 54942 28533 54998
rect 28589 54942 28657 54998
rect 28713 54942 28781 54998
rect 28837 54942 28905 54998
rect 28961 54942 29029 54998
rect 29085 54942 29153 54998
rect 29209 54942 29277 54998
rect 29333 54942 29401 54998
rect 29457 54942 29467 54998
rect 28523 54874 29467 54942
rect 28523 54818 28533 54874
rect 28589 54818 28657 54874
rect 28713 54818 28781 54874
rect 28837 54818 28905 54874
rect 28961 54818 29029 54874
rect 29085 54818 29153 54874
rect 29209 54818 29277 54874
rect 29333 54818 29401 54874
rect 29457 54818 29467 54874
rect 28523 54750 29467 54818
rect 28523 54694 28533 54750
rect 28589 54694 28657 54750
rect 28713 54694 28781 54750
rect 28837 54694 28905 54750
rect 28961 54694 29029 54750
rect 29085 54694 29153 54750
rect 29209 54694 29277 54750
rect 29333 54694 29401 54750
rect 29457 54694 29467 54750
rect 28523 54626 29467 54694
rect 28523 54570 28533 54626
rect 28589 54570 28657 54626
rect 28713 54570 28781 54626
rect 28837 54570 28905 54626
rect 28961 54570 29029 54626
rect 29085 54570 29153 54626
rect 29209 54570 29277 54626
rect 29333 54570 29401 54626
rect 29457 54570 29467 54626
rect 28523 54502 29467 54570
rect 28523 54446 28533 54502
rect 28589 54446 28657 54502
rect 28713 54446 28781 54502
rect 28837 54446 28905 54502
rect 28961 54446 29029 54502
rect 29085 54446 29153 54502
rect 29209 54446 29277 54502
rect 29333 54446 29401 54502
rect 29457 54446 29467 54502
rect 28523 54378 29467 54446
rect 28523 54322 28533 54378
rect 28589 54322 28657 54378
rect 28713 54322 28781 54378
rect 28837 54322 28905 54378
rect 28961 54322 29029 54378
rect 29085 54322 29153 54378
rect 29209 54322 29277 54378
rect 29333 54322 29401 54378
rect 29457 54322 29467 54378
rect 28523 54254 29467 54322
rect 28523 54198 28533 54254
rect 28589 54198 28657 54254
rect 28713 54198 28781 54254
rect 28837 54198 28905 54254
rect 28961 54198 29029 54254
rect 29085 54198 29153 54254
rect 29209 54198 29277 54254
rect 29333 54198 29401 54254
rect 29457 54198 29467 54254
rect 28523 54130 29467 54198
rect 28523 54074 28533 54130
rect 28589 54074 28657 54130
rect 28713 54074 28781 54130
rect 28837 54074 28905 54130
rect 28961 54074 29029 54130
rect 29085 54074 29153 54130
rect 29209 54074 29277 54130
rect 29333 54074 29401 54130
rect 29457 54074 29467 54130
rect 28523 54064 29467 54074
rect 31407 55003 34809 55039
rect 31407 54947 31566 55003
rect 31622 54947 31690 55003
rect 31746 54947 31814 55003
rect 31870 54947 31938 55003
rect 31994 54947 32062 55003
rect 32118 54947 32186 55003
rect 32242 54947 32310 55003
rect 32366 54947 32715 55003
rect 32771 54947 32839 55003
rect 32895 54947 32963 55003
rect 33019 54947 33087 55003
rect 33143 54947 33211 55003
rect 33267 54947 33335 55003
rect 33391 54947 33459 55003
rect 33515 54947 33850 55003
rect 33906 54947 33974 55003
rect 34030 54947 34098 55003
rect 34154 54947 34222 55003
rect 34278 54947 34346 55003
rect 34402 54947 34470 55003
rect 34526 54947 34594 55003
rect 34650 54947 34809 55003
rect 31407 54879 34809 54947
rect 31407 54823 31566 54879
rect 31622 54823 31690 54879
rect 31746 54823 31814 54879
rect 31870 54823 31938 54879
rect 31994 54823 32062 54879
rect 32118 54823 32186 54879
rect 32242 54823 32310 54879
rect 32366 54823 32715 54879
rect 32771 54823 32839 54879
rect 32895 54823 32963 54879
rect 33019 54823 33087 54879
rect 33143 54823 33211 54879
rect 33267 54823 33335 54879
rect 33391 54823 33459 54879
rect 33515 54823 33850 54879
rect 33906 54823 33974 54879
rect 34030 54823 34098 54879
rect 34154 54823 34222 54879
rect 34278 54823 34346 54879
rect 34402 54823 34470 54879
rect 34526 54823 34594 54879
rect 34650 54823 34809 54879
rect 31407 54755 34809 54823
rect 31407 54699 31566 54755
rect 31622 54699 31690 54755
rect 31746 54699 31814 54755
rect 31870 54699 31938 54755
rect 31994 54699 32062 54755
rect 32118 54699 32186 54755
rect 32242 54699 32310 54755
rect 32366 54699 32715 54755
rect 32771 54699 32839 54755
rect 32895 54699 32963 54755
rect 33019 54699 33087 54755
rect 33143 54699 33211 54755
rect 33267 54699 33335 54755
rect 33391 54699 33459 54755
rect 33515 54699 33850 54755
rect 33906 54699 33974 54755
rect 34030 54699 34098 54755
rect 34154 54699 34222 54755
rect 34278 54699 34346 54755
rect 34402 54699 34470 54755
rect 34526 54699 34594 54755
rect 34650 54699 34809 54755
rect 31407 54631 34809 54699
rect 31407 54575 31566 54631
rect 31622 54575 31690 54631
rect 31746 54575 31814 54631
rect 31870 54575 31938 54631
rect 31994 54575 32062 54631
rect 32118 54575 32186 54631
rect 32242 54575 32310 54631
rect 32366 54575 32715 54631
rect 32771 54575 32839 54631
rect 32895 54575 32963 54631
rect 33019 54575 33087 54631
rect 33143 54575 33211 54631
rect 33267 54575 33335 54631
rect 33391 54575 33459 54631
rect 33515 54575 33850 54631
rect 33906 54575 33974 54631
rect 34030 54575 34098 54631
rect 34154 54575 34222 54631
rect 34278 54575 34346 54631
rect 34402 54575 34470 54631
rect 34526 54575 34594 54631
rect 34650 54575 34809 54631
rect 31407 54507 34809 54575
rect 31407 54451 31566 54507
rect 31622 54451 31690 54507
rect 31746 54451 31814 54507
rect 31870 54451 31938 54507
rect 31994 54451 32062 54507
rect 32118 54451 32186 54507
rect 32242 54451 32310 54507
rect 32366 54451 32715 54507
rect 32771 54451 32839 54507
rect 32895 54451 32963 54507
rect 33019 54451 33087 54507
rect 33143 54451 33211 54507
rect 33267 54451 33335 54507
rect 33391 54451 33459 54507
rect 33515 54451 33850 54507
rect 33906 54451 33974 54507
rect 34030 54451 34098 54507
rect 34154 54451 34222 54507
rect 34278 54451 34346 54507
rect 34402 54451 34470 54507
rect 34526 54451 34594 54507
rect 34650 54451 34809 54507
rect 31407 54383 34809 54451
rect 31407 54327 31566 54383
rect 31622 54327 31690 54383
rect 31746 54327 31814 54383
rect 31870 54327 31938 54383
rect 31994 54327 32062 54383
rect 32118 54327 32186 54383
rect 32242 54327 32310 54383
rect 32366 54327 32715 54383
rect 32771 54327 32839 54383
rect 32895 54327 32963 54383
rect 33019 54327 33087 54383
rect 33143 54327 33211 54383
rect 33267 54327 33335 54383
rect 33391 54327 33459 54383
rect 33515 54327 33850 54383
rect 33906 54327 33974 54383
rect 34030 54327 34098 54383
rect 34154 54327 34222 54383
rect 34278 54327 34346 54383
rect 34402 54327 34470 54383
rect 34526 54327 34594 54383
rect 34650 54327 34809 54383
rect 31407 54259 34809 54327
rect 31407 54203 31566 54259
rect 31622 54203 31690 54259
rect 31746 54203 31814 54259
rect 31870 54203 31938 54259
rect 31994 54203 32062 54259
rect 32118 54203 32186 54259
rect 32242 54203 32310 54259
rect 32366 54203 32715 54259
rect 32771 54203 32839 54259
rect 32895 54203 32963 54259
rect 33019 54203 33087 54259
rect 33143 54203 33211 54259
rect 33267 54203 33335 54259
rect 33391 54203 33459 54259
rect 33515 54203 33850 54259
rect 33906 54203 33974 54259
rect 34030 54203 34098 54259
rect 34154 54203 34222 54259
rect 34278 54203 34346 54259
rect 34402 54203 34470 54259
rect 34526 54203 34594 54259
rect 34650 54203 34809 54259
rect 31407 54135 34809 54203
rect 31407 54079 31566 54135
rect 31622 54079 31690 54135
rect 31746 54079 31814 54135
rect 31870 54079 31938 54135
rect 31994 54079 32062 54135
rect 32118 54079 32186 54135
rect 32242 54079 32310 54135
rect 32366 54079 32715 54135
rect 32771 54079 32839 54135
rect 32895 54079 32963 54135
rect 33019 54079 33087 54135
rect 33143 54079 33211 54135
rect 33267 54079 33335 54135
rect 33391 54079 33459 54135
rect 33515 54079 33850 54135
rect 33906 54079 33974 54135
rect 34030 54079 34098 54135
rect 34154 54079 34222 54135
rect 34278 54079 34346 54135
rect 34402 54079 34470 54135
rect 34526 54079 34594 54135
rect 34650 54079 34809 54135
rect 31407 53974 34809 54079
rect 37049 54984 38336 55039
rect 37049 54928 37087 54984
rect 37143 54928 37211 54984
rect 37267 54928 37335 54984
rect 37391 54928 37459 54984
rect 37515 54928 37583 54984
rect 37639 54928 37707 54984
rect 37763 54928 37831 54984
rect 37887 54928 37955 54984
rect 38011 54928 38079 54984
rect 38135 54928 38203 54984
rect 38259 54928 38336 54984
rect 37049 54860 38336 54928
rect 37049 54804 37087 54860
rect 37143 54804 37211 54860
rect 37267 54804 37335 54860
rect 37391 54804 37459 54860
rect 37515 54804 37583 54860
rect 37639 54804 37707 54860
rect 37763 54804 37831 54860
rect 37887 54804 37955 54860
rect 38011 54804 38079 54860
rect 38135 54804 38203 54860
rect 38259 54804 38336 54860
rect 37049 54736 38336 54804
rect 37049 54680 37087 54736
rect 37143 54680 37211 54736
rect 37267 54680 37335 54736
rect 37391 54680 37459 54736
rect 37515 54680 37583 54736
rect 37639 54680 37707 54736
rect 37763 54680 37831 54736
rect 37887 54680 37955 54736
rect 38011 54680 38079 54736
rect 38135 54680 38203 54736
rect 38259 54680 38336 54736
rect 37049 54612 38336 54680
rect 37049 54556 37087 54612
rect 37143 54556 37211 54612
rect 37267 54556 37335 54612
rect 37391 54556 37459 54612
rect 37515 54556 37583 54612
rect 37639 54556 37707 54612
rect 37763 54556 37831 54612
rect 37887 54556 37955 54612
rect 38011 54556 38079 54612
rect 38135 54556 38203 54612
rect 38259 54556 38336 54612
rect 37049 54488 38336 54556
rect 37049 54432 37087 54488
rect 37143 54432 37211 54488
rect 37267 54432 37335 54488
rect 37391 54432 37459 54488
rect 37515 54432 37583 54488
rect 37639 54432 37707 54488
rect 37763 54432 37831 54488
rect 37887 54432 37955 54488
rect 38011 54432 38079 54488
rect 38135 54432 38203 54488
rect 38259 54432 38336 54488
rect 37049 54364 38336 54432
rect 37049 54308 37087 54364
rect 37143 54308 37211 54364
rect 37267 54308 37335 54364
rect 37391 54308 37459 54364
rect 37515 54308 37583 54364
rect 37639 54308 37707 54364
rect 37763 54308 37831 54364
rect 37887 54308 37955 54364
rect 38011 54308 38079 54364
rect 38135 54308 38203 54364
rect 38259 54308 38336 54364
rect 37049 54240 38336 54308
rect 37049 54184 37087 54240
rect 37143 54184 37211 54240
rect 37267 54184 37335 54240
rect 37391 54184 37459 54240
rect 37515 54184 37583 54240
rect 37639 54184 37707 54240
rect 37763 54184 37831 54240
rect 37887 54184 37955 54240
rect 38011 54184 38079 54240
rect 38135 54184 38203 54240
rect 38259 54184 38336 54240
rect 37049 54116 38336 54184
rect 37049 54060 37087 54116
rect 37143 54060 37211 54116
rect 37267 54060 37335 54116
rect 37391 54060 37459 54116
rect 37515 54060 37583 54116
rect 37639 54060 37707 54116
rect 37763 54060 37831 54116
rect 37887 54060 37955 54116
rect 38011 54060 38079 54116
rect 38135 54060 38203 54116
rect 38259 54060 38336 54116
rect 37049 53974 38336 54060
rect 40506 54984 41539 55039
rect 40506 54928 40544 54984
rect 40600 54928 40668 54984
rect 40724 54928 40792 54984
rect 40848 54928 40916 54984
rect 40972 54928 41040 54984
rect 41096 54928 41164 54984
rect 41220 54928 41288 54984
rect 41344 54928 41412 54984
rect 41468 54928 41539 54984
rect 40506 54860 41539 54928
rect 40506 54804 40544 54860
rect 40600 54804 40668 54860
rect 40724 54804 40792 54860
rect 40848 54804 40916 54860
rect 40972 54804 41040 54860
rect 41096 54804 41164 54860
rect 41220 54804 41288 54860
rect 41344 54804 41412 54860
rect 41468 54804 41539 54860
rect 40506 54736 41539 54804
rect 40506 54680 40544 54736
rect 40600 54680 40668 54736
rect 40724 54680 40792 54736
rect 40848 54680 40916 54736
rect 40972 54680 41040 54736
rect 41096 54680 41164 54736
rect 41220 54680 41288 54736
rect 41344 54680 41412 54736
rect 41468 54680 41539 54736
rect 40506 54612 41539 54680
rect 40506 54556 40544 54612
rect 40600 54556 40668 54612
rect 40724 54556 40792 54612
rect 40848 54556 40916 54612
rect 40972 54556 41040 54612
rect 41096 54556 41164 54612
rect 41220 54556 41288 54612
rect 41344 54556 41412 54612
rect 41468 54556 41539 54612
rect 40506 54488 41539 54556
rect 40506 54432 40544 54488
rect 40600 54432 40668 54488
rect 40724 54432 40792 54488
rect 40848 54432 40916 54488
rect 40972 54432 41040 54488
rect 41096 54432 41164 54488
rect 41220 54432 41288 54488
rect 41344 54432 41412 54488
rect 41468 54432 41539 54488
rect 40506 54364 41539 54432
rect 40506 54308 40544 54364
rect 40600 54308 40668 54364
rect 40724 54308 40792 54364
rect 40848 54308 40916 54364
rect 40972 54308 41040 54364
rect 41096 54308 41164 54364
rect 41220 54308 41288 54364
rect 41344 54308 41412 54364
rect 41468 54308 41539 54364
rect 40506 54240 41539 54308
rect 40506 54184 40544 54240
rect 40600 54184 40668 54240
rect 40724 54184 40792 54240
rect 40848 54184 40916 54240
rect 40972 54184 41040 54240
rect 41096 54184 41164 54240
rect 41220 54184 41288 54240
rect 41344 54184 41412 54240
rect 41468 54184 41539 54240
rect 40506 54116 41539 54184
rect 40506 54060 40544 54116
rect 40600 54060 40668 54116
rect 40724 54060 40792 54116
rect 40848 54060 40916 54116
rect 40972 54060 41040 54116
rect 41096 54060 41164 54116
rect 41220 54060 41288 54116
rect 41344 54060 41412 54116
rect 41468 54060 41539 54116
rect 40506 54039 41539 54060
rect 50710 54984 51911 55039
rect 50710 54928 50860 54984
rect 50916 54928 50984 54984
rect 51040 54928 51108 54984
rect 51164 54928 51232 54984
rect 51288 54928 51356 54984
rect 51412 54928 51480 54984
rect 51536 54928 51604 54984
rect 51660 54928 51728 54984
rect 51784 54928 51911 54984
rect 50710 54860 51911 54928
rect 50710 54804 50860 54860
rect 50916 54804 50984 54860
rect 51040 54804 51108 54860
rect 51164 54804 51232 54860
rect 51288 54804 51356 54860
rect 51412 54804 51480 54860
rect 51536 54804 51604 54860
rect 51660 54804 51728 54860
rect 51784 54804 51911 54860
rect 50710 54736 51911 54804
rect 50710 54680 50860 54736
rect 50916 54680 50984 54736
rect 51040 54680 51108 54736
rect 51164 54680 51232 54736
rect 51288 54680 51356 54736
rect 51412 54680 51480 54736
rect 51536 54680 51604 54736
rect 51660 54680 51728 54736
rect 51784 54680 51911 54736
rect 50710 54612 51911 54680
rect 50710 54556 50860 54612
rect 50916 54556 50984 54612
rect 51040 54556 51108 54612
rect 51164 54556 51232 54612
rect 51288 54556 51356 54612
rect 51412 54556 51480 54612
rect 51536 54556 51604 54612
rect 51660 54556 51728 54612
rect 51784 54556 51911 54612
rect 50710 54488 51911 54556
rect 50710 54432 50860 54488
rect 50916 54432 50984 54488
rect 51040 54432 51108 54488
rect 51164 54432 51232 54488
rect 51288 54432 51356 54488
rect 51412 54432 51480 54488
rect 51536 54432 51604 54488
rect 51660 54432 51728 54488
rect 51784 54432 51911 54488
rect 50710 54364 51911 54432
rect 50710 54308 50860 54364
rect 50916 54308 50984 54364
rect 51040 54308 51108 54364
rect 51164 54308 51232 54364
rect 51288 54308 51356 54364
rect 51412 54308 51480 54364
rect 51536 54308 51604 54364
rect 51660 54308 51728 54364
rect 51784 54308 51911 54364
rect 50710 54240 51911 54308
rect 50710 54184 50860 54240
rect 50916 54184 50984 54240
rect 51040 54184 51108 54240
rect 51164 54184 51232 54240
rect 51288 54184 51356 54240
rect 51412 54184 51480 54240
rect 51536 54184 51604 54240
rect 51660 54184 51728 54240
rect 51784 54184 51911 54240
rect 50710 54116 51911 54184
rect 50710 54060 50860 54116
rect 50916 54060 50984 54116
rect 51040 54060 51108 54116
rect 51164 54060 51232 54116
rect 51288 54060 51356 54116
rect 51412 54060 51480 54116
rect 51536 54060 51604 54116
rect 51660 54060 51728 54116
rect 51784 54060 51911 54116
rect 50710 53974 51911 54060
rect 54147 54984 57559 55039
rect 54147 54928 54528 54984
rect 54584 54928 54652 54984
rect 54708 54928 54776 54984
rect 54832 54928 54900 54984
rect 54956 54928 55024 54984
rect 55080 54928 55148 54984
rect 55204 54928 55272 54984
rect 55328 54928 55396 54984
rect 55452 54928 56221 54984
rect 56277 54928 56345 54984
rect 56401 54928 56469 54984
rect 56525 54928 56593 54984
rect 56649 54928 56717 54984
rect 56773 54928 56841 54984
rect 56897 54928 56965 54984
rect 57021 54928 57089 54984
rect 57145 54928 57559 54984
rect 54147 54860 57559 54928
rect 54147 54804 54528 54860
rect 54584 54804 54652 54860
rect 54708 54804 54776 54860
rect 54832 54804 54900 54860
rect 54956 54804 55024 54860
rect 55080 54804 55148 54860
rect 55204 54804 55272 54860
rect 55328 54804 55396 54860
rect 55452 54804 56221 54860
rect 56277 54804 56345 54860
rect 56401 54804 56469 54860
rect 56525 54804 56593 54860
rect 56649 54804 56717 54860
rect 56773 54804 56841 54860
rect 56897 54804 56965 54860
rect 57021 54804 57089 54860
rect 57145 54804 57559 54860
rect 54147 54736 57559 54804
rect 54147 54680 54528 54736
rect 54584 54680 54652 54736
rect 54708 54680 54776 54736
rect 54832 54680 54900 54736
rect 54956 54680 55024 54736
rect 55080 54680 55148 54736
rect 55204 54680 55272 54736
rect 55328 54680 55396 54736
rect 55452 54680 56221 54736
rect 56277 54680 56345 54736
rect 56401 54680 56469 54736
rect 56525 54680 56593 54736
rect 56649 54680 56717 54736
rect 56773 54680 56841 54736
rect 56897 54680 56965 54736
rect 57021 54680 57089 54736
rect 57145 54680 57559 54736
rect 54147 54612 57559 54680
rect 54147 54556 54528 54612
rect 54584 54556 54652 54612
rect 54708 54556 54776 54612
rect 54832 54556 54900 54612
rect 54956 54556 55024 54612
rect 55080 54556 55148 54612
rect 55204 54556 55272 54612
rect 55328 54556 55396 54612
rect 55452 54556 56221 54612
rect 56277 54556 56345 54612
rect 56401 54556 56469 54612
rect 56525 54556 56593 54612
rect 56649 54556 56717 54612
rect 56773 54556 56841 54612
rect 56897 54556 56965 54612
rect 57021 54556 57089 54612
rect 57145 54556 57559 54612
rect 54147 54488 57559 54556
rect 54147 54432 54528 54488
rect 54584 54432 54652 54488
rect 54708 54432 54776 54488
rect 54832 54432 54900 54488
rect 54956 54432 55024 54488
rect 55080 54432 55148 54488
rect 55204 54432 55272 54488
rect 55328 54432 55396 54488
rect 55452 54432 56221 54488
rect 56277 54432 56345 54488
rect 56401 54432 56469 54488
rect 56525 54432 56593 54488
rect 56649 54432 56717 54488
rect 56773 54432 56841 54488
rect 56897 54432 56965 54488
rect 57021 54432 57089 54488
rect 57145 54432 57559 54488
rect 54147 54364 57559 54432
rect 54147 54308 54528 54364
rect 54584 54308 54652 54364
rect 54708 54308 54776 54364
rect 54832 54308 54900 54364
rect 54956 54308 55024 54364
rect 55080 54308 55148 54364
rect 55204 54308 55272 54364
rect 55328 54308 55396 54364
rect 55452 54308 56221 54364
rect 56277 54308 56345 54364
rect 56401 54308 56469 54364
rect 56525 54308 56593 54364
rect 56649 54308 56717 54364
rect 56773 54308 56841 54364
rect 56897 54308 56965 54364
rect 57021 54308 57089 54364
rect 57145 54308 57559 54364
rect 54147 54240 57559 54308
rect 54147 54184 54528 54240
rect 54584 54184 54652 54240
rect 54708 54184 54776 54240
rect 54832 54184 54900 54240
rect 54956 54184 55024 54240
rect 55080 54184 55148 54240
rect 55204 54184 55272 54240
rect 55328 54184 55396 54240
rect 55452 54184 56221 54240
rect 56277 54184 56345 54240
rect 56401 54184 56469 54240
rect 56525 54184 56593 54240
rect 56649 54184 56717 54240
rect 56773 54184 56841 54240
rect 56897 54184 56965 54240
rect 57021 54184 57089 54240
rect 57145 54184 57559 54240
rect 54147 54116 57559 54184
rect 54147 54060 54528 54116
rect 54584 54060 54652 54116
rect 54708 54060 54776 54116
rect 54832 54060 54900 54116
rect 54956 54060 55024 54116
rect 55080 54060 55148 54116
rect 55204 54060 55272 54116
rect 55328 54060 55396 54116
rect 55452 54060 56221 54116
rect 56277 54060 56345 54116
rect 56401 54060 56469 54116
rect 56525 54060 56593 54116
rect 56649 54060 56717 54116
rect 56773 54060 56841 54116
rect 56897 54060 56965 54116
rect 57021 54060 57089 54116
rect 57145 54060 57559 54116
rect 54147 53974 57559 54060
rect 59496 54984 60440 54994
rect 59496 54928 59506 54984
rect 59562 54928 59630 54984
rect 59686 54928 59754 54984
rect 59810 54928 59878 54984
rect 59934 54928 60002 54984
rect 60058 54928 60126 54984
rect 60182 54928 60250 54984
rect 60306 54928 60374 54984
rect 60430 54928 60440 54984
rect 59496 54860 60440 54928
rect 59496 54804 59506 54860
rect 59562 54804 59630 54860
rect 59686 54804 59754 54860
rect 59810 54804 59878 54860
rect 59934 54804 60002 54860
rect 60058 54804 60126 54860
rect 60182 54804 60250 54860
rect 60306 54804 60374 54860
rect 60430 54804 60440 54860
rect 59496 54736 60440 54804
rect 59496 54680 59506 54736
rect 59562 54680 59630 54736
rect 59686 54680 59754 54736
rect 59810 54680 59878 54736
rect 59934 54680 60002 54736
rect 60058 54680 60126 54736
rect 60182 54680 60250 54736
rect 60306 54680 60374 54736
rect 60430 54680 60440 54736
rect 59496 54612 60440 54680
rect 59496 54556 59506 54612
rect 59562 54556 59630 54612
rect 59686 54556 59754 54612
rect 59810 54556 59878 54612
rect 59934 54556 60002 54612
rect 60058 54556 60126 54612
rect 60182 54556 60250 54612
rect 60306 54556 60374 54612
rect 60430 54556 60440 54612
rect 59496 54488 60440 54556
rect 59496 54432 59506 54488
rect 59562 54432 59630 54488
rect 59686 54432 59754 54488
rect 59810 54432 59878 54488
rect 59934 54432 60002 54488
rect 60058 54432 60126 54488
rect 60182 54432 60250 54488
rect 60306 54432 60374 54488
rect 60430 54432 60440 54488
rect 59496 54364 60440 54432
rect 59496 54308 59506 54364
rect 59562 54308 59630 54364
rect 59686 54308 59754 54364
rect 59810 54308 59878 54364
rect 59934 54308 60002 54364
rect 60058 54308 60126 54364
rect 60182 54308 60250 54364
rect 60306 54308 60374 54364
rect 60430 54308 60440 54364
rect 59496 54240 60440 54308
rect 59496 54184 59506 54240
rect 59562 54184 59630 54240
rect 59686 54184 59754 54240
rect 59810 54184 59878 54240
rect 59934 54184 60002 54240
rect 60058 54184 60126 54240
rect 60182 54184 60250 54240
rect 60306 54184 60374 54240
rect 60430 54184 60440 54240
rect 59496 54116 60440 54184
rect 59496 54060 59506 54116
rect 59562 54060 59630 54116
rect 59686 54060 59754 54116
rect 59810 54060 59878 54116
rect 59934 54060 60002 54116
rect 60058 54060 60126 54116
rect 60182 54060 60250 54116
rect 60306 54060 60374 54116
rect 60430 54060 60440 54116
rect 59496 54050 60440 54060
rect 59830 53974 60272 54050
rect 59216 4787 59658 4835
rect 59216 4735 59282 4787
rect 59334 4735 59406 4787
rect 59458 4735 59530 4787
rect 59582 4735 59658 4787
rect 59216 4663 59658 4735
rect 59216 4611 59282 4663
rect 59334 4611 59406 4663
rect 59458 4611 59530 4663
rect 59582 4611 59658 4663
rect 59216 4539 59658 4611
rect 59216 4487 59282 4539
rect 59334 4487 59406 4539
rect 59458 4487 59530 4539
rect 59582 4487 59658 4539
rect 59216 4415 59658 4487
rect 59216 4363 59282 4415
rect 59334 4363 59406 4415
rect 59458 4363 59530 4415
rect 59582 4363 59658 4415
rect 28693 4282 29135 4295
rect 28693 4226 28763 4282
rect 28819 4226 28887 4282
rect 28943 4226 29011 4282
rect 29067 4226 29135 4282
rect 28693 4158 29135 4226
rect 28693 4102 28763 4158
rect 28819 4102 28887 4158
rect 28943 4102 29011 4158
rect 29067 4102 29135 4158
rect 28693 4034 29135 4102
rect 28693 3978 28763 4034
rect 28819 3978 28887 4034
rect 28943 3978 29011 4034
rect 29067 3978 29135 4034
rect 28693 3910 29135 3978
rect 28693 3854 28763 3910
rect 28819 3854 28887 3910
rect 28943 3854 29011 3910
rect 29067 3854 29135 3910
rect 28693 3786 29135 3854
rect 28693 3730 28763 3786
rect 28819 3730 28887 3786
rect 28943 3730 29011 3786
rect 29067 3730 29135 3786
rect 28693 3662 29135 3730
rect 28693 3606 28763 3662
rect 28819 3606 28887 3662
rect 28943 3606 29011 3662
rect 29067 3606 29135 3662
rect 28693 3538 29135 3606
rect 28693 3482 28763 3538
rect 28819 3482 28887 3538
rect 28943 3482 29011 3538
rect 29067 3482 29135 3538
rect 28693 3414 29135 3482
rect 28693 3358 28763 3414
rect 28819 3358 28887 3414
rect 28943 3358 29011 3414
rect 29067 3358 29135 3414
rect 28693 2345 29135 3358
rect 29308 4273 29750 4295
rect 29308 4221 29374 4273
rect 29426 4221 29498 4273
rect 29550 4221 29622 4273
rect 29674 4221 29750 4273
rect 29308 4149 29750 4221
rect 29308 4097 29374 4149
rect 29426 4097 29498 4149
rect 29550 4097 29622 4149
rect 29674 4097 29750 4149
rect 29308 4025 29750 4097
rect 29308 3973 29374 4025
rect 29426 3973 29498 4025
rect 29550 3973 29622 4025
rect 29674 3973 29750 4025
rect 29308 3901 29750 3973
rect 29308 3849 29374 3901
rect 29426 3849 29498 3901
rect 29550 3849 29622 3901
rect 29674 3849 29750 3901
rect 29308 3777 29750 3849
rect 29308 3725 29374 3777
rect 29426 3725 29498 3777
rect 29550 3725 29622 3777
rect 29674 3725 29750 3777
rect 29308 3653 29750 3725
rect 29308 3601 29374 3653
rect 29426 3601 29498 3653
rect 29550 3601 29622 3653
rect 29674 3601 29750 3653
rect 29308 3529 29750 3601
rect 29308 3477 29374 3529
rect 29426 3477 29498 3529
rect 29550 3477 29622 3529
rect 29674 3477 29750 3529
rect 29308 3405 29750 3477
rect 29308 3353 29374 3405
rect 29426 3353 29498 3405
rect 29550 3353 29622 3405
rect 29674 3353 29750 3405
rect 29308 3281 29750 3353
rect 29308 3229 29374 3281
rect 29426 3229 29498 3281
rect 29550 3229 29622 3281
rect 29674 3229 29750 3281
rect 29308 3157 29750 3229
rect 29308 3105 29374 3157
rect 29426 3105 29498 3157
rect 29550 3105 29622 3157
rect 29674 3105 29750 3157
rect 29308 3033 29750 3105
rect 29308 2981 29374 3033
rect 29426 2981 29498 3033
rect 29550 2981 29622 3033
rect 29674 2981 29750 3033
rect 29308 2909 29750 2981
rect 29308 2857 29374 2909
rect 29426 2857 29498 2909
rect 29550 2857 29622 2909
rect 29674 2857 29750 2909
rect 29308 2785 29750 2857
rect 29308 2733 29374 2785
rect 29426 2733 29498 2785
rect 29550 2733 29622 2785
rect 29674 2733 29750 2785
rect 29308 2661 29750 2733
rect 29308 2609 29374 2661
rect 29426 2609 29498 2661
rect 29550 2609 29622 2661
rect 29674 2609 29750 2661
rect 29308 2537 29750 2609
rect 29308 2485 29374 2537
rect 29426 2485 29498 2537
rect 29550 2485 29622 2537
rect 29674 2485 29750 2537
rect 29308 2413 29750 2485
rect 29308 2361 29374 2413
rect 29426 2361 29498 2413
rect 29550 2361 29622 2413
rect 29674 2361 29750 2413
rect 29308 2345 29750 2361
rect 59216 4291 59658 4363
rect 59216 4239 59282 4291
rect 59334 4239 59406 4291
rect 59458 4239 59530 4291
rect 59582 4239 59658 4291
rect 59216 4167 59658 4239
rect 59216 4115 59282 4167
rect 59334 4115 59406 4167
rect 59458 4115 59530 4167
rect 59582 4115 59658 4167
rect 59216 4043 59658 4115
rect 59216 3991 59282 4043
rect 59334 3991 59406 4043
rect 59458 3991 59530 4043
rect 59582 3991 59658 4043
rect 59216 3919 59658 3991
rect 59216 3867 59282 3919
rect 59334 3867 59406 3919
rect 59458 3867 59530 3919
rect 59582 3867 59658 3919
rect 59216 3795 59658 3867
rect 59216 3743 59282 3795
rect 59334 3743 59406 3795
rect 59458 3743 59530 3795
rect 59582 3743 59658 3795
rect 59216 3671 59658 3743
rect 59216 3619 59282 3671
rect 59334 3619 59406 3671
rect 59458 3619 59530 3671
rect 59582 3619 59658 3671
rect 59216 3547 59658 3619
rect 59216 3495 59282 3547
rect 59334 3495 59406 3547
rect 59458 3495 59530 3547
rect 59582 3495 59658 3547
rect 59216 3423 59658 3495
rect 59216 3371 59282 3423
rect 59334 3371 59406 3423
rect 59458 3371 59530 3423
rect 59582 3371 59658 3423
rect 59216 3299 59658 3371
rect 59216 3247 59282 3299
rect 59334 3247 59406 3299
rect 59458 3247 59530 3299
rect 59582 3247 59658 3299
rect 59830 4282 60272 4295
rect 59830 4226 59900 4282
rect 59956 4226 60024 4282
rect 60080 4226 60148 4282
rect 60204 4226 60272 4282
rect 59830 4158 60272 4226
rect 59830 4102 59900 4158
rect 59956 4102 60024 4158
rect 60080 4102 60148 4158
rect 60204 4102 60272 4158
rect 59830 4034 60272 4102
rect 59830 3978 59900 4034
rect 59956 3978 60024 4034
rect 60080 3978 60148 4034
rect 60204 3978 60272 4034
rect 59830 3910 60272 3978
rect 59830 3854 59900 3910
rect 59956 3854 60024 3910
rect 60080 3854 60148 3910
rect 60204 3854 60272 3910
rect 59830 3786 60272 3854
rect 59830 3730 59900 3786
rect 59956 3730 60024 3786
rect 60080 3730 60148 3786
rect 60204 3730 60272 3786
rect 59830 3662 60272 3730
rect 59830 3606 59900 3662
rect 59956 3606 60024 3662
rect 60080 3606 60148 3662
rect 60204 3606 60272 3662
rect 59830 3538 60272 3606
rect 59830 3482 59900 3538
rect 59956 3482 60024 3538
rect 60080 3482 60148 3538
rect 60204 3482 60272 3538
rect 59830 3414 60272 3482
rect 59830 3358 59900 3414
rect 59956 3358 60024 3414
rect 60080 3358 60148 3414
rect 60204 3358 60272 3414
rect 59830 3295 60272 3358
rect 59216 3175 59658 3247
rect 59216 3123 59282 3175
rect 59334 3123 59406 3175
rect 59458 3123 59530 3175
rect 59582 3123 59658 3175
rect 59216 3051 59658 3123
rect 59216 2999 59282 3051
rect 59334 2999 59406 3051
rect 59458 2999 59530 3051
rect 59582 2999 59658 3051
rect 59216 2927 59658 2999
rect 59216 2875 59282 2927
rect 59334 2875 59406 2927
rect 59458 2875 59530 2927
rect 59582 2875 59658 2927
rect 59216 2803 59658 2875
rect 59216 2751 59282 2803
rect 59334 2751 59406 2803
rect 59458 2751 59530 2803
rect 59582 2751 59658 2803
rect 59216 2679 59658 2751
rect 59216 2627 59282 2679
rect 59334 2627 59406 2679
rect 59458 2627 59530 2679
rect 59582 2627 59658 2679
rect 59216 2555 59658 2627
rect 59216 2503 59282 2555
rect 59334 2503 59406 2555
rect 59458 2503 59530 2555
rect 59582 2503 59658 2555
rect 59216 2431 59658 2503
rect 59216 2379 59282 2431
rect 59334 2379 59406 2431
rect 59458 2379 59530 2431
rect 59582 2379 59658 2431
rect 59216 2345 59658 2379
rect 86587 2345 87587 55029
<< via2 >>
rect 27128 55545 27184 55547
rect 27128 55493 27130 55545
rect 27130 55493 27182 55545
rect 27182 55493 27184 55545
rect 27128 55491 27184 55493
rect 27252 55545 27308 55547
rect 27252 55493 27254 55545
rect 27254 55493 27306 55545
rect 27306 55493 27308 55545
rect 27252 55491 27308 55493
rect 27376 55545 27432 55547
rect 27376 55493 27378 55545
rect 27378 55493 27430 55545
rect 27430 55493 27432 55545
rect 27376 55491 27432 55493
rect 27500 55545 27556 55547
rect 27500 55493 27502 55545
rect 27502 55493 27554 55545
rect 27554 55493 27556 55545
rect 27500 55491 27556 55493
rect 27624 55545 27680 55547
rect 27624 55493 27626 55545
rect 27626 55493 27678 55545
rect 27678 55493 27680 55545
rect 27624 55491 27680 55493
rect 27748 55545 27804 55547
rect 27748 55493 27750 55545
rect 27750 55493 27802 55545
rect 27802 55493 27804 55545
rect 27748 55491 27804 55493
rect 27872 55545 27928 55547
rect 27872 55493 27874 55545
rect 27874 55493 27926 55545
rect 27926 55493 27928 55545
rect 27872 55491 27928 55493
rect 27996 55545 28052 55547
rect 27996 55493 27998 55545
rect 27998 55493 28050 55545
rect 28050 55493 28052 55545
rect 27996 55491 28052 55493
rect 27128 55421 27184 55423
rect 27128 55369 27130 55421
rect 27130 55369 27182 55421
rect 27182 55369 27184 55421
rect 27128 55367 27184 55369
rect 27252 55421 27308 55423
rect 27252 55369 27254 55421
rect 27254 55369 27306 55421
rect 27306 55369 27308 55421
rect 27252 55367 27308 55369
rect 27376 55421 27432 55423
rect 27376 55369 27378 55421
rect 27378 55369 27430 55421
rect 27430 55369 27432 55421
rect 27376 55367 27432 55369
rect 27500 55421 27556 55423
rect 27500 55369 27502 55421
rect 27502 55369 27554 55421
rect 27554 55369 27556 55421
rect 27500 55367 27556 55369
rect 27624 55421 27680 55423
rect 27624 55369 27626 55421
rect 27626 55369 27678 55421
rect 27678 55369 27680 55421
rect 27624 55367 27680 55369
rect 27748 55421 27804 55423
rect 27748 55369 27750 55421
rect 27750 55369 27802 55421
rect 27802 55369 27804 55421
rect 27748 55367 27804 55369
rect 27872 55421 27928 55423
rect 27872 55369 27874 55421
rect 27874 55369 27926 55421
rect 27926 55369 27928 55421
rect 27872 55367 27928 55369
rect 27996 55421 28052 55423
rect 27996 55369 27998 55421
rect 27998 55369 28050 55421
rect 28050 55369 28052 55421
rect 27996 55367 28052 55369
rect 27128 55297 27184 55299
rect 27128 55245 27130 55297
rect 27130 55245 27182 55297
rect 27182 55245 27184 55297
rect 27128 55243 27184 55245
rect 27252 55297 27308 55299
rect 27252 55245 27254 55297
rect 27254 55245 27306 55297
rect 27306 55245 27308 55297
rect 27252 55243 27308 55245
rect 27376 55297 27432 55299
rect 27376 55245 27378 55297
rect 27378 55245 27430 55297
rect 27430 55245 27432 55297
rect 27376 55243 27432 55245
rect 27500 55297 27556 55299
rect 27500 55245 27502 55297
rect 27502 55245 27554 55297
rect 27554 55245 27556 55297
rect 27500 55243 27556 55245
rect 27624 55297 27680 55299
rect 27624 55245 27626 55297
rect 27626 55245 27678 55297
rect 27678 55245 27680 55297
rect 27624 55243 27680 55245
rect 27748 55297 27804 55299
rect 27748 55245 27750 55297
rect 27750 55245 27802 55297
rect 27802 55245 27804 55297
rect 27748 55243 27804 55245
rect 27872 55297 27928 55299
rect 27872 55245 27874 55297
rect 27874 55245 27926 55297
rect 27926 55245 27928 55297
rect 27872 55243 27928 55245
rect 27996 55297 28052 55299
rect 27996 55245 27998 55297
rect 27998 55245 28050 55297
rect 28050 55245 28052 55297
rect 27996 55243 28052 55245
rect 35984 55545 36040 55547
rect 35984 55493 35986 55545
rect 35986 55493 36038 55545
rect 36038 55493 36040 55545
rect 35984 55491 36040 55493
rect 36108 55545 36164 55547
rect 36108 55493 36110 55545
rect 36110 55493 36162 55545
rect 36162 55493 36164 55545
rect 36108 55491 36164 55493
rect 36232 55545 36288 55547
rect 36232 55493 36234 55545
rect 36234 55493 36286 55545
rect 36286 55493 36288 55545
rect 36232 55491 36288 55493
rect 36356 55545 36412 55547
rect 36356 55493 36358 55545
rect 36358 55493 36410 55545
rect 36410 55493 36412 55545
rect 36356 55491 36412 55493
rect 36480 55545 36536 55547
rect 36480 55493 36482 55545
rect 36482 55493 36534 55545
rect 36534 55493 36536 55545
rect 36480 55491 36536 55493
rect 36604 55545 36660 55547
rect 36604 55493 36606 55545
rect 36606 55493 36658 55545
rect 36658 55493 36660 55545
rect 36604 55491 36660 55493
rect 36728 55545 36784 55547
rect 36728 55493 36730 55545
rect 36730 55493 36782 55545
rect 36782 55493 36784 55545
rect 36728 55491 36784 55493
rect 36852 55545 36908 55547
rect 36852 55493 36854 55545
rect 36854 55493 36906 55545
rect 36906 55493 36908 55545
rect 36852 55491 36908 55493
rect 35984 55421 36040 55423
rect 35984 55369 35986 55421
rect 35986 55369 36038 55421
rect 36038 55369 36040 55421
rect 35984 55367 36040 55369
rect 36108 55421 36164 55423
rect 36108 55369 36110 55421
rect 36110 55369 36162 55421
rect 36162 55369 36164 55421
rect 36108 55367 36164 55369
rect 36232 55421 36288 55423
rect 36232 55369 36234 55421
rect 36234 55369 36286 55421
rect 36286 55369 36288 55421
rect 36232 55367 36288 55369
rect 36356 55421 36412 55423
rect 36356 55369 36358 55421
rect 36358 55369 36410 55421
rect 36410 55369 36412 55421
rect 36356 55367 36412 55369
rect 36480 55421 36536 55423
rect 36480 55369 36482 55421
rect 36482 55369 36534 55421
rect 36534 55369 36536 55421
rect 36480 55367 36536 55369
rect 36604 55421 36660 55423
rect 36604 55369 36606 55421
rect 36606 55369 36658 55421
rect 36658 55369 36660 55421
rect 36604 55367 36660 55369
rect 36728 55421 36784 55423
rect 36728 55369 36730 55421
rect 36730 55369 36782 55421
rect 36782 55369 36784 55421
rect 36728 55367 36784 55369
rect 36852 55421 36908 55423
rect 36852 55369 36854 55421
rect 36854 55369 36906 55421
rect 36906 55369 36908 55421
rect 36852 55367 36908 55369
rect 35984 55297 36040 55299
rect 35984 55245 35986 55297
rect 35986 55245 36038 55297
rect 36038 55245 36040 55297
rect 35984 55243 36040 55245
rect 36108 55297 36164 55299
rect 36108 55245 36110 55297
rect 36110 55245 36162 55297
rect 36162 55245 36164 55297
rect 36108 55243 36164 55245
rect 36232 55297 36288 55299
rect 36232 55245 36234 55297
rect 36234 55245 36286 55297
rect 36286 55245 36288 55297
rect 36232 55243 36288 55245
rect 36356 55297 36412 55299
rect 36356 55245 36358 55297
rect 36358 55245 36410 55297
rect 36410 55245 36412 55297
rect 36356 55243 36412 55245
rect 36480 55297 36536 55299
rect 36480 55245 36482 55297
rect 36482 55245 36534 55297
rect 36534 55245 36536 55297
rect 36480 55243 36536 55245
rect 36604 55297 36660 55299
rect 36604 55245 36606 55297
rect 36606 55245 36658 55297
rect 36658 55245 36660 55297
rect 36604 55243 36660 55245
rect 36728 55297 36784 55299
rect 36728 55245 36730 55297
rect 36730 55245 36782 55297
rect 36782 55245 36784 55297
rect 36728 55243 36784 55245
rect 36852 55297 36908 55299
rect 36852 55245 36854 55297
rect 36854 55245 36906 55297
rect 36906 55245 36908 55297
rect 36852 55243 36908 55245
rect 41826 55545 41882 55547
rect 41826 55493 41828 55545
rect 41828 55493 41880 55545
rect 41880 55493 41882 55545
rect 41826 55491 41882 55493
rect 41950 55545 42006 55547
rect 41950 55493 41952 55545
rect 41952 55493 42004 55545
rect 42004 55493 42006 55545
rect 41950 55491 42006 55493
rect 42074 55545 42130 55547
rect 42074 55493 42076 55545
rect 42076 55493 42128 55545
rect 42128 55493 42130 55545
rect 42074 55491 42130 55493
rect 42198 55545 42254 55547
rect 42198 55493 42200 55545
rect 42200 55493 42252 55545
rect 42252 55493 42254 55545
rect 42198 55491 42254 55493
rect 42322 55545 42378 55547
rect 42322 55493 42324 55545
rect 42324 55493 42376 55545
rect 42376 55493 42378 55545
rect 42322 55491 42378 55493
rect 42446 55545 42502 55547
rect 42446 55493 42448 55545
rect 42448 55493 42500 55545
rect 42500 55493 42502 55545
rect 42446 55491 42502 55493
rect 42570 55545 42626 55547
rect 42570 55493 42572 55545
rect 42572 55493 42624 55545
rect 42624 55493 42626 55545
rect 42570 55491 42626 55493
rect 42694 55545 42750 55547
rect 42694 55493 42696 55545
rect 42696 55493 42748 55545
rect 42748 55493 42750 55545
rect 42694 55491 42750 55493
rect 41826 55421 41882 55423
rect 41826 55369 41828 55421
rect 41828 55369 41880 55421
rect 41880 55369 41882 55421
rect 41826 55367 41882 55369
rect 41950 55421 42006 55423
rect 41950 55369 41952 55421
rect 41952 55369 42004 55421
rect 42004 55369 42006 55421
rect 41950 55367 42006 55369
rect 42074 55421 42130 55423
rect 42074 55369 42076 55421
rect 42076 55369 42128 55421
rect 42128 55369 42130 55421
rect 42074 55367 42130 55369
rect 42198 55421 42254 55423
rect 42198 55369 42200 55421
rect 42200 55369 42252 55421
rect 42252 55369 42254 55421
rect 42198 55367 42254 55369
rect 42322 55421 42378 55423
rect 42322 55369 42324 55421
rect 42324 55369 42376 55421
rect 42376 55369 42378 55421
rect 42322 55367 42378 55369
rect 42446 55421 42502 55423
rect 42446 55369 42448 55421
rect 42448 55369 42500 55421
rect 42500 55369 42502 55421
rect 42446 55367 42502 55369
rect 42570 55421 42626 55423
rect 42570 55369 42572 55421
rect 42572 55369 42624 55421
rect 42624 55369 42626 55421
rect 42570 55367 42626 55369
rect 42694 55421 42750 55423
rect 42694 55369 42696 55421
rect 42696 55369 42748 55421
rect 42748 55369 42750 55421
rect 42694 55367 42750 55369
rect 41826 55297 41882 55299
rect 41826 55245 41828 55297
rect 41828 55245 41880 55297
rect 41880 55245 41882 55297
rect 41826 55243 41882 55245
rect 41950 55297 42006 55299
rect 41950 55245 41952 55297
rect 41952 55245 42004 55297
rect 42004 55245 42006 55297
rect 41950 55243 42006 55245
rect 42074 55297 42130 55299
rect 42074 55245 42076 55297
rect 42076 55245 42128 55297
rect 42128 55245 42130 55297
rect 42074 55243 42130 55245
rect 42198 55297 42254 55299
rect 42198 55245 42200 55297
rect 42200 55245 42252 55297
rect 42252 55245 42254 55297
rect 42198 55243 42254 55245
rect 42322 55297 42378 55299
rect 42322 55245 42324 55297
rect 42324 55245 42376 55297
rect 42376 55245 42378 55297
rect 42322 55243 42378 55245
rect 42446 55297 42502 55299
rect 42446 55245 42448 55297
rect 42448 55245 42500 55297
rect 42500 55245 42502 55297
rect 42446 55243 42502 55245
rect 42570 55297 42626 55299
rect 42570 55245 42572 55297
rect 42572 55245 42624 55297
rect 42624 55245 42626 55297
rect 42570 55243 42626 55245
rect 42694 55297 42750 55299
rect 42694 55245 42696 55297
rect 42696 55245 42748 55297
rect 42748 55245 42750 55297
rect 42694 55243 42750 55245
rect 45657 55545 45713 55547
rect 45657 55493 45659 55545
rect 45659 55493 45711 55545
rect 45711 55493 45713 55545
rect 45657 55491 45713 55493
rect 45781 55545 45837 55547
rect 45781 55493 45783 55545
rect 45783 55493 45835 55545
rect 45835 55493 45837 55545
rect 45781 55491 45837 55493
rect 45905 55545 45961 55547
rect 45905 55493 45907 55545
rect 45907 55493 45959 55545
rect 45959 55493 45961 55545
rect 45905 55491 45961 55493
rect 46029 55545 46085 55547
rect 46029 55493 46031 55545
rect 46031 55493 46083 55545
rect 46083 55493 46085 55545
rect 46029 55491 46085 55493
rect 46153 55545 46209 55547
rect 46153 55493 46155 55545
rect 46155 55493 46207 55545
rect 46207 55493 46209 55545
rect 46153 55491 46209 55493
rect 46277 55545 46333 55547
rect 46277 55493 46279 55545
rect 46279 55493 46331 55545
rect 46331 55493 46333 55545
rect 46277 55491 46333 55493
rect 46401 55545 46457 55547
rect 46401 55493 46403 55545
rect 46403 55493 46455 55545
rect 46455 55493 46457 55545
rect 46401 55491 46457 55493
rect 46525 55545 46581 55547
rect 46525 55493 46527 55545
rect 46527 55493 46579 55545
rect 46579 55493 46581 55545
rect 46525 55491 46581 55493
rect 45657 55421 45713 55423
rect 45657 55369 45659 55421
rect 45659 55369 45711 55421
rect 45711 55369 45713 55421
rect 45657 55367 45713 55369
rect 45781 55421 45837 55423
rect 45781 55369 45783 55421
rect 45783 55369 45835 55421
rect 45835 55369 45837 55421
rect 45781 55367 45837 55369
rect 45905 55421 45961 55423
rect 45905 55369 45907 55421
rect 45907 55369 45959 55421
rect 45959 55369 45961 55421
rect 45905 55367 45961 55369
rect 46029 55421 46085 55423
rect 46029 55369 46031 55421
rect 46031 55369 46083 55421
rect 46083 55369 46085 55421
rect 46029 55367 46085 55369
rect 46153 55421 46209 55423
rect 46153 55369 46155 55421
rect 46155 55369 46207 55421
rect 46207 55369 46209 55421
rect 46153 55367 46209 55369
rect 46277 55421 46333 55423
rect 46277 55369 46279 55421
rect 46279 55369 46331 55421
rect 46331 55369 46333 55421
rect 46277 55367 46333 55369
rect 46401 55421 46457 55423
rect 46401 55369 46403 55421
rect 46403 55369 46455 55421
rect 46455 55369 46457 55421
rect 46401 55367 46457 55369
rect 46525 55421 46581 55423
rect 46525 55369 46527 55421
rect 46527 55369 46579 55421
rect 46579 55369 46581 55421
rect 46525 55367 46581 55369
rect 45657 55297 45713 55299
rect 45657 55245 45659 55297
rect 45659 55245 45711 55297
rect 45711 55245 45713 55297
rect 45657 55243 45713 55245
rect 45781 55297 45837 55299
rect 45781 55245 45783 55297
rect 45783 55245 45835 55297
rect 45835 55245 45837 55297
rect 45781 55243 45837 55245
rect 45905 55297 45961 55299
rect 45905 55245 45907 55297
rect 45907 55245 45959 55297
rect 45959 55245 45961 55297
rect 45905 55243 45961 55245
rect 46029 55297 46085 55299
rect 46029 55245 46031 55297
rect 46031 55245 46083 55297
rect 46083 55245 46085 55297
rect 46029 55243 46085 55245
rect 46153 55297 46209 55299
rect 46153 55245 46155 55297
rect 46155 55245 46207 55297
rect 46207 55245 46209 55297
rect 46153 55243 46209 55245
rect 46277 55297 46333 55299
rect 46277 55245 46279 55297
rect 46279 55245 46331 55297
rect 46331 55245 46333 55297
rect 46277 55243 46333 55245
rect 46401 55297 46457 55299
rect 46401 55245 46403 55297
rect 46403 55245 46455 55297
rect 46455 55245 46457 55297
rect 46401 55243 46457 55245
rect 46525 55297 46581 55299
rect 46525 55245 46527 55297
rect 46527 55245 46579 55297
rect 46579 55245 46581 55297
rect 46525 55243 46581 55245
rect 52409 55545 52465 55547
rect 52409 55493 52411 55545
rect 52411 55493 52463 55545
rect 52463 55493 52465 55545
rect 52409 55491 52465 55493
rect 52533 55545 52589 55547
rect 52533 55493 52535 55545
rect 52535 55493 52587 55545
rect 52587 55493 52589 55545
rect 52533 55491 52589 55493
rect 52657 55545 52713 55547
rect 52657 55493 52659 55545
rect 52659 55493 52711 55545
rect 52711 55493 52713 55545
rect 52657 55491 52713 55493
rect 52781 55545 52837 55547
rect 52781 55493 52783 55545
rect 52783 55493 52835 55545
rect 52835 55493 52837 55545
rect 52781 55491 52837 55493
rect 52905 55545 52961 55547
rect 52905 55493 52907 55545
rect 52907 55493 52959 55545
rect 52959 55493 52961 55545
rect 52905 55491 52961 55493
rect 53029 55545 53085 55547
rect 53029 55493 53031 55545
rect 53031 55493 53083 55545
rect 53083 55493 53085 55545
rect 53029 55491 53085 55493
rect 53153 55545 53209 55547
rect 53153 55493 53155 55545
rect 53155 55493 53207 55545
rect 53207 55493 53209 55545
rect 53153 55491 53209 55493
rect 53277 55545 53333 55547
rect 53277 55493 53279 55545
rect 53279 55493 53331 55545
rect 53331 55493 53333 55545
rect 53277 55491 53333 55493
rect 52409 55421 52465 55423
rect 52409 55369 52411 55421
rect 52411 55369 52463 55421
rect 52463 55369 52465 55421
rect 52409 55367 52465 55369
rect 52533 55421 52589 55423
rect 52533 55369 52535 55421
rect 52535 55369 52587 55421
rect 52587 55369 52589 55421
rect 52533 55367 52589 55369
rect 52657 55421 52713 55423
rect 52657 55369 52659 55421
rect 52659 55369 52711 55421
rect 52711 55369 52713 55421
rect 52657 55367 52713 55369
rect 52781 55421 52837 55423
rect 52781 55369 52783 55421
rect 52783 55369 52835 55421
rect 52835 55369 52837 55421
rect 52781 55367 52837 55369
rect 52905 55421 52961 55423
rect 52905 55369 52907 55421
rect 52907 55369 52959 55421
rect 52959 55369 52961 55421
rect 52905 55367 52961 55369
rect 53029 55421 53085 55423
rect 53029 55369 53031 55421
rect 53031 55369 53083 55421
rect 53083 55369 53085 55421
rect 53029 55367 53085 55369
rect 53153 55421 53209 55423
rect 53153 55369 53155 55421
rect 53155 55369 53207 55421
rect 53207 55369 53209 55421
rect 53153 55367 53209 55369
rect 53277 55421 53333 55423
rect 53277 55369 53279 55421
rect 53279 55369 53331 55421
rect 53331 55369 53333 55421
rect 53277 55367 53333 55369
rect 52409 55297 52465 55299
rect 52409 55245 52411 55297
rect 52411 55245 52463 55297
rect 52463 55245 52465 55297
rect 52409 55243 52465 55245
rect 52533 55297 52589 55299
rect 52533 55245 52535 55297
rect 52535 55245 52587 55297
rect 52587 55245 52589 55297
rect 52533 55243 52589 55245
rect 52657 55297 52713 55299
rect 52657 55245 52659 55297
rect 52659 55245 52711 55297
rect 52711 55245 52713 55297
rect 52657 55243 52713 55245
rect 52781 55297 52837 55299
rect 52781 55245 52783 55297
rect 52783 55245 52835 55297
rect 52835 55245 52837 55297
rect 52781 55243 52837 55245
rect 52905 55297 52961 55299
rect 52905 55245 52907 55297
rect 52907 55245 52959 55297
rect 52959 55245 52961 55297
rect 52905 55243 52961 55245
rect 53029 55297 53085 55299
rect 53029 55245 53031 55297
rect 53031 55245 53083 55297
rect 53083 55245 53085 55297
rect 53029 55243 53085 55245
rect 53153 55297 53209 55299
rect 53153 55245 53155 55297
rect 53155 55245 53207 55297
rect 53207 55245 53209 55297
rect 53153 55243 53209 55245
rect 53277 55297 53333 55299
rect 53277 55245 53279 55297
rect 53279 55245 53331 55297
rect 53331 55245 53333 55297
rect 53277 55243 53333 55245
rect 57934 55545 57990 55547
rect 57934 55493 57936 55545
rect 57936 55493 57988 55545
rect 57988 55493 57990 55545
rect 57934 55491 57990 55493
rect 58058 55545 58114 55547
rect 58058 55493 58060 55545
rect 58060 55493 58112 55545
rect 58112 55493 58114 55545
rect 58058 55491 58114 55493
rect 58182 55545 58238 55547
rect 58182 55493 58184 55545
rect 58184 55493 58236 55545
rect 58236 55493 58238 55545
rect 58182 55491 58238 55493
rect 58306 55545 58362 55547
rect 58306 55493 58308 55545
rect 58308 55493 58360 55545
rect 58360 55493 58362 55545
rect 58306 55491 58362 55493
rect 58430 55545 58486 55547
rect 58430 55493 58432 55545
rect 58432 55493 58484 55545
rect 58484 55493 58486 55545
rect 58430 55491 58486 55493
rect 58554 55545 58610 55547
rect 58554 55493 58556 55545
rect 58556 55493 58608 55545
rect 58608 55493 58610 55545
rect 58554 55491 58610 55493
rect 58678 55545 58734 55547
rect 58678 55493 58680 55545
rect 58680 55493 58732 55545
rect 58732 55493 58734 55545
rect 58678 55491 58734 55493
rect 58802 55545 58858 55547
rect 58802 55493 58804 55545
rect 58804 55493 58856 55545
rect 58856 55493 58858 55545
rect 58802 55491 58858 55493
rect 57934 55421 57990 55423
rect 57934 55369 57936 55421
rect 57936 55369 57988 55421
rect 57988 55369 57990 55421
rect 57934 55367 57990 55369
rect 58058 55421 58114 55423
rect 58058 55369 58060 55421
rect 58060 55369 58112 55421
rect 58112 55369 58114 55421
rect 58058 55367 58114 55369
rect 58182 55421 58238 55423
rect 58182 55369 58184 55421
rect 58184 55369 58236 55421
rect 58236 55369 58238 55421
rect 58182 55367 58238 55369
rect 58306 55421 58362 55423
rect 58306 55369 58308 55421
rect 58308 55369 58360 55421
rect 58360 55369 58362 55421
rect 58306 55367 58362 55369
rect 58430 55421 58486 55423
rect 58430 55369 58432 55421
rect 58432 55369 58484 55421
rect 58484 55369 58486 55421
rect 58430 55367 58486 55369
rect 58554 55421 58610 55423
rect 58554 55369 58556 55421
rect 58556 55369 58608 55421
rect 58608 55369 58610 55421
rect 58554 55367 58610 55369
rect 58678 55421 58734 55423
rect 58678 55369 58680 55421
rect 58680 55369 58732 55421
rect 58732 55369 58734 55421
rect 58678 55367 58734 55369
rect 58802 55421 58858 55423
rect 58802 55369 58804 55421
rect 58804 55369 58856 55421
rect 58856 55369 58858 55421
rect 58802 55367 58858 55369
rect 57934 55297 57990 55299
rect 57934 55245 57936 55297
rect 57936 55245 57988 55297
rect 57988 55245 57990 55297
rect 57934 55243 57990 55245
rect 58058 55297 58114 55299
rect 58058 55245 58060 55297
rect 58060 55245 58112 55297
rect 58112 55245 58114 55297
rect 58058 55243 58114 55245
rect 58182 55297 58238 55299
rect 58182 55245 58184 55297
rect 58184 55245 58236 55297
rect 58236 55245 58238 55297
rect 58182 55243 58238 55245
rect 58306 55297 58362 55299
rect 58306 55245 58308 55297
rect 58308 55245 58360 55297
rect 58360 55245 58362 55297
rect 58306 55243 58362 55245
rect 58430 55297 58486 55299
rect 58430 55245 58432 55297
rect 58432 55245 58484 55297
rect 58484 55245 58486 55297
rect 58430 55243 58486 55245
rect 58554 55297 58610 55299
rect 58554 55245 58556 55297
rect 58556 55245 58608 55297
rect 58608 55245 58610 55297
rect 58554 55243 58610 55245
rect 58678 55297 58734 55299
rect 58678 55245 58680 55297
rect 58680 55245 58732 55297
rect 58732 55245 58734 55297
rect 58678 55243 58734 55245
rect 58802 55297 58858 55299
rect 58802 55245 58804 55297
rect 58804 55245 58856 55297
rect 58856 55245 58858 55297
rect 58802 55243 58858 55245
rect 60735 55545 60791 55547
rect 60735 55493 60737 55545
rect 60737 55493 60789 55545
rect 60789 55493 60791 55545
rect 60735 55491 60791 55493
rect 60859 55545 60915 55547
rect 60859 55493 60861 55545
rect 60861 55493 60913 55545
rect 60913 55493 60915 55545
rect 60859 55491 60915 55493
rect 60983 55545 61039 55547
rect 60983 55493 60985 55545
rect 60985 55493 61037 55545
rect 61037 55493 61039 55545
rect 60983 55491 61039 55493
rect 61107 55545 61163 55547
rect 61107 55493 61109 55545
rect 61109 55493 61161 55545
rect 61161 55493 61163 55545
rect 61107 55491 61163 55493
rect 61231 55545 61287 55547
rect 61231 55493 61233 55545
rect 61233 55493 61285 55545
rect 61285 55493 61287 55545
rect 61231 55491 61287 55493
rect 61355 55545 61411 55547
rect 61355 55493 61357 55545
rect 61357 55493 61409 55545
rect 61409 55493 61411 55545
rect 61355 55491 61411 55493
rect 61479 55545 61535 55547
rect 61479 55493 61481 55545
rect 61481 55493 61533 55545
rect 61533 55493 61535 55545
rect 61479 55491 61535 55493
rect 61603 55545 61659 55547
rect 61603 55493 61605 55545
rect 61605 55493 61657 55545
rect 61657 55493 61659 55545
rect 61603 55491 61659 55493
rect 60735 55421 60791 55423
rect 60735 55369 60737 55421
rect 60737 55369 60789 55421
rect 60789 55369 60791 55421
rect 60735 55367 60791 55369
rect 60859 55421 60915 55423
rect 60859 55369 60861 55421
rect 60861 55369 60913 55421
rect 60913 55369 60915 55421
rect 60859 55367 60915 55369
rect 60983 55421 61039 55423
rect 60983 55369 60985 55421
rect 60985 55369 61037 55421
rect 61037 55369 61039 55421
rect 60983 55367 61039 55369
rect 61107 55421 61163 55423
rect 61107 55369 61109 55421
rect 61109 55369 61161 55421
rect 61161 55369 61163 55421
rect 61107 55367 61163 55369
rect 61231 55421 61287 55423
rect 61231 55369 61233 55421
rect 61233 55369 61285 55421
rect 61285 55369 61287 55421
rect 61231 55367 61287 55369
rect 61355 55421 61411 55423
rect 61355 55369 61357 55421
rect 61357 55369 61409 55421
rect 61409 55369 61411 55421
rect 61355 55367 61411 55369
rect 61479 55421 61535 55423
rect 61479 55369 61481 55421
rect 61481 55369 61533 55421
rect 61533 55369 61535 55421
rect 61479 55367 61535 55369
rect 61603 55421 61659 55423
rect 61603 55369 61605 55421
rect 61605 55369 61657 55421
rect 61657 55369 61659 55421
rect 61603 55367 61659 55369
rect 60735 55297 60791 55299
rect 60735 55245 60737 55297
rect 60737 55245 60789 55297
rect 60789 55245 60791 55297
rect 60735 55243 60791 55245
rect 60859 55297 60915 55299
rect 60859 55245 60861 55297
rect 60861 55245 60913 55297
rect 60913 55245 60915 55297
rect 60859 55243 60915 55245
rect 60983 55297 61039 55299
rect 60983 55245 60985 55297
rect 60985 55245 61037 55297
rect 61037 55245 61039 55297
rect 60983 55243 61039 55245
rect 61107 55297 61163 55299
rect 61107 55245 61109 55297
rect 61109 55245 61161 55297
rect 61161 55245 61163 55297
rect 61107 55243 61163 55245
rect 61231 55297 61287 55299
rect 61231 55245 61233 55297
rect 61233 55245 61285 55297
rect 61285 55245 61287 55297
rect 61231 55243 61287 55245
rect 61355 55297 61411 55299
rect 61355 55245 61357 55297
rect 61357 55245 61409 55297
rect 61409 55245 61411 55297
rect 61355 55243 61411 55245
rect 61479 55297 61535 55299
rect 61479 55245 61481 55297
rect 61481 55245 61533 55297
rect 61533 55245 61535 55297
rect 61479 55243 61535 55245
rect 61603 55297 61659 55299
rect 61603 55245 61605 55297
rect 61605 55245 61657 55297
rect 61657 55245 61659 55297
rect 61603 55243 61659 55245
rect 28533 54942 28589 54998
rect 28657 54942 28713 54998
rect 28781 54942 28837 54998
rect 28905 54942 28961 54998
rect 29029 54942 29085 54998
rect 29153 54942 29209 54998
rect 29277 54942 29333 54998
rect 29401 54942 29457 54998
rect 28533 54818 28589 54874
rect 28657 54818 28713 54874
rect 28781 54818 28837 54874
rect 28905 54818 28961 54874
rect 29029 54818 29085 54874
rect 29153 54818 29209 54874
rect 29277 54818 29333 54874
rect 29401 54818 29457 54874
rect 28533 54694 28589 54750
rect 28657 54694 28713 54750
rect 28781 54694 28837 54750
rect 28905 54694 28961 54750
rect 29029 54694 29085 54750
rect 29153 54694 29209 54750
rect 29277 54694 29333 54750
rect 29401 54694 29457 54750
rect 28533 54570 28589 54626
rect 28657 54570 28713 54626
rect 28781 54570 28837 54626
rect 28905 54570 28961 54626
rect 29029 54570 29085 54626
rect 29153 54570 29209 54626
rect 29277 54570 29333 54626
rect 29401 54570 29457 54626
rect 28533 54446 28589 54502
rect 28657 54446 28713 54502
rect 28781 54446 28837 54502
rect 28905 54446 28961 54502
rect 29029 54446 29085 54502
rect 29153 54446 29209 54502
rect 29277 54446 29333 54502
rect 29401 54446 29457 54502
rect 28533 54322 28589 54378
rect 28657 54322 28713 54378
rect 28781 54322 28837 54378
rect 28905 54322 28961 54378
rect 29029 54322 29085 54378
rect 29153 54322 29209 54378
rect 29277 54322 29333 54378
rect 29401 54322 29457 54378
rect 28533 54198 28589 54254
rect 28657 54198 28713 54254
rect 28781 54198 28837 54254
rect 28905 54198 28961 54254
rect 29029 54198 29085 54254
rect 29153 54198 29209 54254
rect 29277 54198 29333 54254
rect 29401 54198 29457 54254
rect 28533 54074 28589 54130
rect 28657 54074 28713 54130
rect 28781 54074 28837 54130
rect 28905 54074 28961 54130
rect 29029 54074 29085 54130
rect 29153 54074 29209 54130
rect 29277 54074 29333 54130
rect 29401 54074 29457 54130
rect 31566 54947 31622 55003
rect 31690 54947 31746 55003
rect 31814 54947 31870 55003
rect 31938 54947 31994 55003
rect 32062 54947 32118 55003
rect 32186 54947 32242 55003
rect 32310 54947 32366 55003
rect 32715 54947 32771 55003
rect 32839 54947 32895 55003
rect 32963 54947 33019 55003
rect 33087 54947 33143 55003
rect 33211 54947 33267 55003
rect 33335 54947 33391 55003
rect 33459 54947 33515 55003
rect 33850 54947 33906 55003
rect 33974 54947 34030 55003
rect 34098 54947 34154 55003
rect 34222 54947 34278 55003
rect 34346 54947 34402 55003
rect 34470 54947 34526 55003
rect 34594 54947 34650 55003
rect 31566 54823 31622 54879
rect 31690 54823 31746 54879
rect 31814 54823 31870 54879
rect 31938 54823 31994 54879
rect 32062 54823 32118 54879
rect 32186 54823 32242 54879
rect 32310 54823 32366 54879
rect 32715 54823 32771 54879
rect 32839 54823 32895 54879
rect 32963 54823 33019 54879
rect 33087 54823 33143 54879
rect 33211 54823 33267 54879
rect 33335 54823 33391 54879
rect 33459 54823 33515 54879
rect 33850 54823 33906 54879
rect 33974 54823 34030 54879
rect 34098 54823 34154 54879
rect 34222 54823 34278 54879
rect 34346 54823 34402 54879
rect 34470 54823 34526 54879
rect 34594 54823 34650 54879
rect 31566 54699 31622 54755
rect 31690 54699 31746 54755
rect 31814 54699 31870 54755
rect 31938 54699 31994 54755
rect 32062 54699 32118 54755
rect 32186 54699 32242 54755
rect 32310 54699 32366 54755
rect 32715 54699 32771 54755
rect 32839 54699 32895 54755
rect 32963 54699 33019 54755
rect 33087 54699 33143 54755
rect 33211 54699 33267 54755
rect 33335 54699 33391 54755
rect 33459 54699 33515 54755
rect 33850 54699 33906 54755
rect 33974 54699 34030 54755
rect 34098 54699 34154 54755
rect 34222 54699 34278 54755
rect 34346 54699 34402 54755
rect 34470 54699 34526 54755
rect 34594 54699 34650 54755
rect 31566 54575 31622 54631
rect 31690 54575 31746 54631
rect 31814 54575 31870 54631
rect 31938 54575 31994 54631
rect 32062 54575 32118 54631
rect 32186 54575 32242 54631
rect 32310 54575 32366 54631
rect 32715 54575 32771 54631
rect 32839 54575 32895 54631
rect 32963 54575 33019 54631
rect 33087 54575 33143 54631
rect 33211 54575 33267 54631
rect 33335 54575 33391 54631
rect 33459 54575 33515 54631
rect 33850 54575 33906 54631
rect 33974 54575 34030 54631
rect 34098 54575 34154 54631
rect 34222 54575 34278 54631
rect 34346 54575 34402 54631
rect 34470 54575 34526 54631
rect 34594 54575 34650 54631
rect 31566 54451 31622 54507
rect 31690 54451 31746 54507
rect 31814 54451 31870 54507
rect 31938 54451 31994 54507
rect 32062 54451 32118 54507
rect 32186 54451 32242 54507
rect 32310 54451 32366 54507
rect 32715 54451 32771 54507
rect 32839 54451 32895 54507
rect 32963 54451 33019 54507
rect 33087 54451 33143 54507
rect 33211 54451 33267 54507
rect 33335 54451 33391 54507
rect 33459 54451 33515 54507
rect 33850 54451 33906 54507
rect 33974 54451 34030 54507
rect 34098 54451 34154 54507
rect 34222 54451 34278 54507
rect 34346 54451 34402 54507
rect 34470 54451 34526 54507
rect 34594 54451 34650 54507
rect 31566 54327 31622 54383
rect 31690 54327 31746 54383
rect 31814 54327 31870 54383
rect 31938 54327 31994 54383
rect 32062 54327 32118 54383
rect 32186 54327 32242 54383
rect 32310 54327 32366 54383
rect 32715 54327 32771 54383
rect 32839 54327 32895 54383
rect 32963 54327 33019 54383
rect 33087 54327 33143 54383
rect 33211 54327 33267 54383
rect 33335 54327 33391 54383
rect 33459 54327 33515 54383
rect 33850 54327 33906 54383
rect 33974 54327 34030 54383
rect 34098 54327 34154 54383
rect 34222 54327 34278 54383
rect 34346 54327 34402 54383
rect 34470 54327 34526 54383
rect 34594 54327 34650 54383
rect 31566 54203 31622 54259
rect 31690 54203 31746 54259
rect 31814 54203 31870 54259
rect 31938 54203 31994 54259
rect 32062 54203 32118 54259
rect 32186 54203 32242 54259
rect 32310 54203 32366 54259
rect 32715 54203 32771 54259
rect 32839 54203 32895 54259
rect 32963 54203 33019 54259
rect 33087 54203 33143 54259
rect 33211 54203 33267 54259
rect 33335 54203 33391 54259
rect 33459 54203 33515 54259
rect 33850 54203 33906 54259
rect 33974 54203 34030 54259
rect 34098 54203 34154 54259
rect 34222 54203 34278 54259
rect 34346 54203 34402 54259
rect 34470 54203 34526 54259
rect 34594 54203 34650 54259
rect 31566 54079 31622 54135
rect 31690 54079 31746 54135
rect 31814 54079 31870 54135
rect 31938 54079 31994 54135
rect 32062 54079 32118 54135
rect 32186 54079 32242 54135
rect 32310 54079 32366 54135
rect 32715 54079 32771 54135
rect 32839 54079 32895 54135
rect 32963 54079 33019 54135
rect 33087 54079 33143 54135
rect 33211 54079 33267 54135
rect 33335 54079 33391 54135
rect 33459 54079 33515 54135
rect 33850 54079 33906 54135
rect 33974 54079 34030 54135
rect 34098 54079 34154 54135
rect 34222 54079 34278 54135
rect 34346 54079 34402 54135
rect 34470 54079 34526 54135
rect 34594 54079 34650 54135
rect 37087 54928 37143 54984
rect 37211 54928 37267 54984
rect 37335 54928 37391 54984
rect 37459 54928 37515 54984
rect 37583 54928 37639 54984
rect 37707 54928 37763 54984
rect 37831 54928 37887 54984
rect 37955 54928 38011 54984
rect 38079 54928 38135 54984
rect 38203 54928 38259 54984
rect 37087 54804 37143 54860
rect 37211 54804 37267 54860
rect 37335 54804 37391 54860
rect 37459 54804 37515 54860
rect 37583 54804 37639 54860
rect 37707 54804 37763 54860
rect 37831 54804 37887 54860
rect 37955 54804 38011 54860
rect 38079 54804 38135 54860
rect 38203 54804 38259 54860
rect 37087 54680 37143 54736
rect 37211 54680 37267 54736
rect 37335 54680 37391 54736
rect 37459 54680 37515 54736
rect 37583 54680 37639 54736
rect 37707 54680 37763 54736
rect 37831 54680 37887 54736
rect 37955 54680 38011 54736
rect 38079 54680 38135 54736
rect 38203 54680 38259 54736
rect 37087 54556 37143 54612
rect 37211 54556 37267 54612
rect 37335 54556 37391 54612
rect 37459 54556 37515 54612
rect 37583 54556 37639 54612
rect 37707 54556 37763 54612
rect 37831 54556 37887 54612
rect 37955 54556 38011 54612
rect 38079 54556 38135 54612
rect 38203 54556 38259 54612
rect 37087 54432 37143 54488
rect 37211 54432 37267 54488
rect 37335 54432 37391 54488
rect 37459 54432 37515 54488
rect 37583 54432 37639 54488
rect 37707 54432 37763 54488
rect 37831 54432 37887 54488
rect 37955 54432 38011 54488
rect 38079 54432 38135 54488
rect 38203 54432 38259 54488
rect 37087 54308 37143 54364
rect 37211 54308 37267 54364
rect 37335 54308 37391 54364
rect 37459 54308 37515 54364
rect 37583 54308 37639 54364
rect 37707 54308 37763 54364
rect 37831 54308 37887 54364
rect 37955 54308 38011 54364
rect 38079 54308 38135 54364
rect 38203 54308 38259 54364
rect 37087 54184 37143 54240
rect 37211 54184 37267 54240
rect 37335 54184 37391 54240
rect 37459 54184 37515 54240
rect 37583 54184 37639 54240
rect 37707 54184 37763 54240
rect 37831 54184 37887 54240
rect 37955 54184 38011 54240
rect 38079 54184 38135 54240
rect 38203 54184 38259 54240
rect 37087 54060 37143 54116
rect 37211 54060 37267 54116
rect 37335 54060 37391 54116
rect 37459 54060 37515 54116
rect 37583 54060 37639 54116
rect 37707 54060 37763 54116
rect 37831 54060 37887 54116
rect 37955 54060 38011 54116
rect 38079 54060 38135 54116
rect 38203 54060 38259 54116
rect 40544 54928 40600 54984
rect 40668 54928 40724 54984
rect 40792 54928 40848 54984
rect 40916 54928 40972 54984
rect 41040 54928 41096 54984
rect 41164 54928 41220 54984
rect 41288 54928 41344 54984
rect 41412 54928 41468 54984
rect 40544 54804 40600 54860
rect 40668 54804 40724 54860
rect 40792 54804 40848 54860
rect 40916 54804 40972 54860
rect 41040 54804 41096 54860
rect 41164 54804 41220 54860
rect 41288 54804 41344 54860
rect 41412 54804 41468 54860
rect 40544 54680 40600 54736
rect 40668 54680 40724 54736
rect 40792 54680 40848 54736
rect 40916 54680 40972 54736
rect 41040 54680 41096 54736
rect 41164 54680 41220 54736
rect 41288 54680 41344 54736
rect 41412 54680 41468 54736
rect 40544 54556 40600 54612
rect 40668 54556 40724 54612
rect 40792 54556 40848 54612
rect 40916 54556 40972 54612
rect 41040 54556 41096 54612
rect 41164 54556 41220 54612
rect 41288 54556 41344 54612
rect 41412 54556 41468 54612
rect 40544 54432 40600 54488
rect 40668 54432 40724 54488
rect 40792 54432 40848 54488
rect 40916 54432 40972 54488
rect 41040 54432 41096 54488
rect 41164 54432 41220 54488
rect 41288 54432 41344 54488
rect 41412 54432 41468 54488
rect 40544 54308 40600 54364
rect 40668 54308 40724 54364
rect 40792 54308 40848 54364
rect 40916 54308 40972 54364
rect 41040 54308 41096 54364
rect 41164 54308 41220 54364
rect 41288 54308 41344 54364
rect 41412 54308 41468 54364
rect 40544 54184 40600 54240
rect 40668 54184 40724 54240
rect 40792 54184 40848 54240
rect 40916 54184 40972 54240
rect 41040 54184 41096 54240
rect 41164 54184 41220 54240
rect 41288 54184 41344 54240
rect 41412 54184 41468 54240
rect 40544 54060 40600 54116
rect 40668 54060 40724 54116
rect 40792 54060 40848 54116
rect 40916 54060 40972 54116
rect 41040 54060 41096 54116
rect 41164 54060 41220 54116
rect 41288 54060 41344 54116
rect 41412 54060 41468 54116
rect 50860 54928 50916 54984
rect 50984 54928 51040 54984
rect 51108 54928 51164 54984
rect 51232 54928 51288 54984
rect 51356 54928 51412 54984
rect 51480 54928 51536 54984
rect 51604 54928 51660 54984
rect 51728 54928 51784 54984
rect 50860 54804 50916 54860
rect 50984 54804 51040 54860
rect 51108 54804 51164 54860
rect 51232 54804 51288 54860
rect 51356 54804 51412 54860
rect 51480 54804 51536 54860
rect 51604 54804 51660 54860
rect 51728 54804 51784 54860
rect 50860 54680 50916 54736
rect 50984 54680 51040 54736
rect 51108 54680 51164 54736
rect 51232 54680 51288 54736
rect 51356 54680 51412 54736
rect 51480 54680 51536 54736
rect 51604 54680 51660 54736
rect 51728 54680 51784 54736
rect 50860 54556 50916 54612
rect 50984 54556 51040 54612
rect 51108 54556 51164 54612
rect 51232 54556 51288 54612
rect 51356 54556 51412 54612
rect 51480 54556 51536 54612
rect 51604 54556 51660 54612
rect 51728 54556 51784 54612
rect 50860 54432 50916 54488
rect 50984 54432 51040 54488
rect 51108 54432 51164 54488
rect 51232 54432 51288 54488
rect 51356 54432 51412 54488
rect 51480 54432 51536 54488
rect 51604 54432 51660 54488
rect 51728 54432 51784 54488
rect 50860 54308 50916 54364
rect 50984 54308 51040 54364
rect 51108 54308 51164 54364
rect 51232 54308 51288 54364
rect 51356 54308 51412 54364
rect 51480 54308 51536 54364
rect 51604 54308 51660 54364
rect 51728 54308 51784 54364
rect 50860 54184 50916 54240
rect 50984 54184 51040 54240
rect 51108 54184 51164 54240
rect 51232 54184 51288 54240
rect 51356 54184 51412 54240
rect 51480 54184 51536 54240
rect 51604 54184 51660 54240
rect 51728 54184 51784 54240
rect 50860 54060 50916 54116
rect 50984 54060 51040 54116
rect 51108 54060 51164 54116
rect 51232 54060 51288 54116
rect 51356 54060 51412 54116
rect 51480 54060 51536 54116
rect 51604 54060 51660 54116
rect 51728 54060 51784 54116
rect 54528 54928 54584 54984
rect 54652 54928 54708 54984
rect 54776 54928 54832 54984
rect 54900 54928 54956 54984
rect 55024 54928 55080 54984
rect 55148 54928 55204 54984
rect 55272 54928 55328 54984
rect 55396 54928 55452 54984
rect 56221 54928 56277 54984
rect 56345 54928 56401 54984
rect 56469 54928 56525 54984
rect 56593 54928 56649 54984
rect 56717 54928 56773 54984
rect 56841 54928 56897 54984
rect 56965 54928 57021 54984
rect 57089 54928 57145 54984
rect 54528 54804 54584 54860
rect 54652 54804 54708 54860
rect 54776 54804 54832 54860
rect 54900 54804 54956 54860
rect 55024 54804 55080 54860
rect 55148 54804 55204 54860
rect 55272 54804 55328 54860
rect 55396 54804 55452 54860
rect 56221 54804 56277 54860
rect 56345 54804 56401 54860
rect 56469 54804 56525 54860
rect 56593 54804 56649 54860
rect 56717 54804 56773 54860
rect 56841 54804 56897 54860
rect 56965 54804 57021 54860
rect 57089 54804 57145 54860
rect 54528 54680 54584 54736
rect 54652 54680 54708 54736
rect 54776 54680 54832 54736
rect 54900 54680 54956 54736
rect 55024 54680 55080 54736
rect 55148 54680 55204 54736
rect 55272 54680 55328 54736
rect 55396 54680 55452 54736
rect 56221 54680 56277 54736
rect 56345 54680 56401 54736
rect 56469 54680 56525 54736
rect 56593 54680 56649 54736
rect 56717 54680 56773 54736
rect 56841 54680 56897 54736
rect 56965 54680 57021 54736
rect 57089 54680 57145 54736
rect 54528 54556 54584 54612
rect 54652 54556 54708 54612
rect 54776 54556 54832 54612
rect 54900 54556 54956 54612
rect 55024 54556 55080 54612
rect 55148 54556 55204 54612
rect 55272 54556 55328 54612
rect 55396 54556 55452 54612
rect 56221 54556 56277 54612
rect 56345 54556 56401 54612
rect 56469 54556 56525 54612
rect 56593 54556 56649 54612
rect 56717 54556 56773 54612
rect 56841 54556 56897 54612
rect 56965 54556 57021 54612
rect 57089 54556 57145 54612
rect 54528 54432 54584 54488
rect 54652 54432 54708 54488
rect 54776 54432 54832 54488
rect 54900 54432 54956 54488
rect 55024 54432 55080 54488
rect 55148 54432 55204 54488
rect 55272 54432 55328 54488
rect 55396 54432 55452 54488
rect 56221 54432 56277 54488
rect 56345 54432 56401 54488
rect 56469 54432 56525 54488
rect 56593 54432 56649 54488
rect 56717 54432 56773 54488
rect 56841 54432 56897 54488
rect 56965 54432 57021 54488
rect 57089 54432 57145 54488
rect 54528 54308 54584 54364
rect 54652 54308 54708 54364
rect 54776 54308 54832 54364
rect 54900 54308 54956 54364
rect 55024 54308 55080 54364
rect 55148 54308 55204 54364
rect 55272 54308 55328 54364
rect 55396 54308 55452 54364
rect 56221 54308 56277 54364
rect 56345 54308 56401 54364
rect 56469 54308 56525 54364
rect 56593 54308 56649 54364
rect 56717 54308 56773 54364
rect 56841 54308 56897 54364
rect 56965 54308 57021 54364
rect 57089 54308 57145 54364
rect 54528 54184 54584 54240
rect 54652 54184 54708 54240
rect 54776 54184 54832 54240
rect 54900 54184 54956 54240
rect 55024 54184 55080 54240
rect 55148 54184 55204 54240
rect 55272 54184 55328 54240
rect 55396 54184 55452 54240
rect 56221 54184 56277 54240
rect 56345 54184 56401 54240
rect 56469 54184 56525 54240
rect 56593 54184 56649 54240
rect 56717 54184 56773 54240
rect 56841 54184 56897 54240
rect 56965 54184 57021 54240
rect 57089 54184 57145 54240
rect 54528 54060 54584 54116
rect 54652 54060 54708 54116
rect 54776 54060 54832 54116
rect 54900 54060 54956 54116
rect 55024 54060 55080 54116
rect 55148 54060 55204 54116
rect 55272 54060 55328 54116
rect 55396 54060 55452 54116
rect 56221 54060 56277 54116
rect 56345 54060 56401 54116
rect 56469 54060 56525 54116
rect 56593 54060 56649 54116
rect 56717 54060 56773 54116
rect 56841 54060 56897 54116
rect 56965 54060 57021 54116
rect 57089 54060 57145 54116
rect 59506 54928 59562 54984
rect 59630 54928 59686 54984
rect 59754 54928 59810 54984
rect 59878 54928 59934 54984
rect 60002 54928 60058 54984
rect 60126 54928 60182 54984
rect 60250 54928 60306 54984
rect 60374 54928 60430 54984
rect 59506 54804 59562 54860
rect 59630 54804 59686 54860
rect 59754 54804 59810 54860
rect 59878 54804 59934 54860
rect 60002 54804 60058 54860
rect 60126 54804 60182 54860
rect 60250 54804 60306 54860
rect 60374 54804 60430 54860
rect 59506 54680 59562 54736
rect 59630 54680 59686 54736
rect 59754 54680 59810 54736
rect 59878 54680 59934 54736
rect 60002 54680 60058 54736
rect 60126 54680 60182 54736
rect 60250 54680 60306 54736
rect 60374 54680 60430 54736
rect 59506 54556 59562 54612
rect 59630 54556 59686 54612
rect 59754 54556 59810 54612
rect 59878 54556 59934 54612
rect 60002 54556 60058 54612
rect 60126 54556 60182 54612
rect 60250 54556 60306 54612
rect 60374 54556 60430 54612
rect 59506 54432 59562 54488
rect 59630 54432 59686 54488
rect 59754 54432 59810 54488
rect 59878 54432 59934 54488
rect 60002 54432 60058 54488
rect 60126 54432 60182 54488
rect 60250 54432 60306 54488
rect 60374 54432 60430 54488
rect 59506 54308 59562 54364
rect 59630 54308 59686 54364
rect 59754 54308 59810 54364
rect 59878 54308 59934 54364
rect 60002 54308 60058 54364
rect 60126 54308 60182 54364
rect 60250 54308 60306 54364
rect 60374 54308 60430 54364
rect 59506 54184 59562 54240
rect 59630 54184 59686 54240
rect 59754 54184 59810 54240
rect 59878 54184 59934 54240
rect 60002 54184 60058 54240
rect 60126 54184 60182 54240
rect 60250 54184 60306 54240
rect 60374 54184 60430 54240
rect 59506 54060 59562 54116
rect 59630 54060 59686 54116
rect 59754 54060 59810 54116
rect 59878 54060 59934 54116
rect 60002 54060 60058 54116
rect 60126 54060 60182 54116
rect 60250 54060 60306 54116
rect 60374 54060 60430 54116
rect 28763 4280 28819 4282
rect 28763 4228 28765 4280
rect 28765 4228 28817 4280
rect 28817 4228 28819 4280
rect 28763 4226 28819 4228
rect 28887 4280 28943 4282
rect 28887 4228 28889 4280
rect 28889 4228 28941 4280
rect 28941 4228 28943 4280
rect 28887 4226 28943 4228
rect 29011 4280 29067 4282
rect 29011 4228 29013 4280
rect 29013 4228 29065 4280
rect 29065 4228 29067 4280
rect 29011 4226 29067 4228
rect 28763 4156 28819 4158
rect 28763 4104 28765 4156
rect 28765 4104 28817 4156
rect 28817 4104 28819 4156
rect 28763 4102 28819 4104
rect 28887 4156 28943 4158
rect 28887 4104 28889 4156
rect 28889 4104 28941 4156
rect 28941 4104 28943 4156
rect 28887 4102 28943 4104
rect 29011 4156 29067 4158
rect 29011 4104 29013 4156
rect 29013 4104 29065 4156
rect 29065 4104 29067 4156
rect 29011 4102 29067 4104
rect 28763 4032 28819 4034
rect 28763 3980 28765 4032
rect 28765 3980 28817 4032
rect 28817 3980 28819 4032
rect 28763 3978 28819 3980
rect 28887 4032 28943 4034
rect 28887 3980 28889 4032
rect 28889 3980 28941 4032
rect 28941 3980 28943 4032
rect 28887 3978 28943 3980
rect 29011 4032 29067 4034
rect 29011 3980 29013 4032
rect 29013 3980 29065 4032
rect 29065 3980 29067 4032
rect 29011 3978 29067 3980
rect 28763 3908 28819 3910
rect 28763 3856 28765 3908
rect 28765 3856 28817 3908
rect 28817 3856 28819 3908
rect 28763 3854 28819 3856
rect 28887 3908 28943 3910
rect 28887 3856 28889 3908
rect 28889 3856 28941 3908
rect 28941 3856 28943 3908
rect 28887 3854 28943 3856
rect 29011 3908 29067 3910
rect 29011 3856 29013 3908
rect 29013 3856 29065 3908
rect 29065 3856 29067 3908
rect 29011 3854 29067 3856
rect 28763 3730 28819 3786
rect 28887 3730 28943 3786
rect 29011 3730 29067 3786
rect 28763 3606 28819 3662
rect 28887 3606 28943 3662
rect 29011 3606 29067 3662
rect 28763 3482 28819 3538
rect 28887 3482 28943 3538
rect 29011 3482 29067 3538
rect 28763 3358 28819 3414
rect 28887 3358 28943 3414
rect 29011 3358 29067 3414
rect 59900 4280 59956 4282
rect 59900 4228 59902 4280
rect 59902 4228 59954 4280
rect 59954 4228 59956 4280
rect 59900 4226 59956 4228
rect 60024 4280 60080 4282
rect 60024 4228 60026 4280
rect 60026 4228 60078 4280
rect 60078 4228 60080 4280
rect 60024 4226 60080 4228
rect 60148 4280 60204 4282
rect 60148 4228 60150 4280
rect 60150 4228 60202 4280
rect 60202 4228 60204 4280
rect 60148 4226 60204 4228
rect 59900 4156 59956 4158
rect 59900 4104 59902 4156
rect 59902 4104 59954 4156
rect 59954 4104 59956 4156
rect 59900 4102 59956 4104
rect 60024 4156 60080 4158
rect 60024 4104 60026 4156
rect 60026 4104 60078 4156
rect 60078 4104 60080 4156
rect 60024 4102 60080 4104
rect 60148 4156 60204 4158
rect 60148 4104 60150 4156
rect 60150 4104 60202 4156
rect 60202 4104 60204 4156
rect 60148 4102 60204 4104
rect 59900 4032 59956 4034
rect 59900 3980 59902 4032
rect 59902 3980 59954 4032
rect 59954 3980 59956 4032
rect 59900 3978 59956 3980
rect 60024 4032 60080 4034
rect 60024 3980 60026 4032
rect 60026 3980 60078 4032
rect 60078 3980 60080 4032
rect 60024 3978 60080 3980
rect 60148 4032 60204 4034
rect 60148 3980 60150 4032
rect 60150 3980 60202 4032
rect 60202 3980 60204 4032
rect 60148 3978 60204 3980
rect 59900 3908 59956 3910
rect 59900 3856 59902 3908
rect 59902 3856 59954 3908
rect 59954 3856 59956 3908
rect 59900 3854 59956 3856
rect 60024 3908 60080 3910
rect 60024 3856 60026 3908
rect 60026 3856 60078 3908
rect 60078 3856 60080 3908
rect 60024 3854 60080 3856
rect 60148 3908 60204 3910
rect 60148 3856 60150 3908
rect 60150 3856 60202 3908
rect 60202 3856 60204 3908
rect 60148 3854 60204 3856
rect 59900 3730 59956 3786
rect 60024 3730 60080 3786
rect 60148 3730 60204 3786
rect 59900 3606 59956 3662
rect 60024 3606 60080 3662
rect 60148 3606 60204 3662
rect 59900 3482 59956 3538
rect 60024 3482 60080 3538
rect 60148 3482 60204 3538
rect 59900 3358 59956 3414
rect 60024 3358 60080 3414
rect 60148 3358 60204 3414
<< metal3 >>
rect 27079 55547 28079 55839
rect 27079 55491 27128 55547
rect 27184 55491 27252 55547
rect 27308 55491 27376 55547
rect 27432 55491 27500 55547
rect 27556 55491 27624 55547
rect 27680 55491 27748 55547
rect 27804 55491 27872 55547
rect 27928 55491 27996 55547
rect 28052 55491 28079 55547
rect 27079 55423 28079 55491
rect 27079 55367 27128 55423
rect 27184 55367 27252 55423
rect 27308 55367 27376 55423
rect 27432 55367 27500 55423
rect 27556 55367 27624 55423
rect 27680 55367 27748 55423
rect 27804 55367 27872 55423
rect 27928 55367 27996 55423
rect 28052 55367 28079 55423
rect 27079 55299 28079 55367
rect 27079 55243 27128 55299
rect 27184 55243 27252 55299
rect 27308 55243 27376 55299
rect 27432 55243 27500 55299
rect 27556 55243 27624 55299
rect 27680 55243 27748 55299
rect 27804 55243 27872 55299
rect 27928 55243 27996 55299
rect 28052 55243 28079 55299
rect 27079 55231 28079 55243
rect 28493 55039 29493 55839
rect 32631 55039 33631 55839
rect 35945 55547 36945 55839
rect 35945 55491 35984 55547
rect 36040 55491 36108 55547
rect 36164 55491 36232 55547
rect 36288 55491 36356 55547
rect 36412 55491 36480 55547
rect 36536 55491 36604 55547
rect 36660 55491 36728 55547
rect 36784 55491 36852 55547
rect 36908 55491 36945 55547
rect 35945 55423 36945 55491
rect 35945 55367 35984 55423
rect 36040 55367 36108 55423
rect 36164 55367 36232 55423
rect 36288 55367 36356 55423
rect 36412 55367 36480 55423
rect 36536 55367 36604 55423
rect 36660 55367 36728 55423
rect 36784 55367 36852 55423
rect 36908 55367 36945 55423
rect 35945 55299 36945 55367
rect 35945 55243 35984 55299
rect 36040 55243 36108 55299
rect 36164 55243 36232 55299
rect 36288 55243 36356 55299
rect 36412 55243 36480 55299
rect 36536 55243 36604 55299
rect 36660 55243 36728 55299
rect 36784 55243 36852 55299
rect 36908 55243 36945 55299
rect 35945 55231 36945 55243
rect 37336 55039 38336 55839
rect 40506 55039 41506 55839
rect 41803 55547 42803 55839
rect 41803 55491 41826 55547
rect 41882 55491 41950 55547
rect 42006 55491 42074 55547
rect 42130 55491 42198 55547
rect 42254 55491 42322 55547
rect 42378 55491 42446 55547
rect 42502 55491 42570 55547
rect 42626 55491 42694 55547
rect 42750 55491 42803 55547
rect 41803 55423 42803 55491
rect 41803 55367 41826 55423
rect 41882 55367 41950 55423
rect 42006 55367 42074 55423
rect 42130 55367 42198 55423
rect 42254 55367 42322 55423
rect 42378 55367 42446 55423
rect 42502 55367 42570 55423
rect 42626 55367 42694 55423
rect 42750 55367 42803 55423
rect 41803 55299 42803 55367
rect 41803 55243 41826 55299
rect 41882 55243 41950 55299
rect 42006 55243 42074 55299
rect 42130 55243 42198 55299
rect 42254 55243 42322 55299
rect 42378 55243 42446 55299
rect 42502 55243 42570 55299
rect 42626 55243 42694 55299
rect 42750 55243 42803 55299
rect 41803 55231 42803 55243
rect 45634 55547 46634 55839
rect 45634 55491 45657 55547
rect 45713 55491 45781 55547
rect 45837 55491 45905 55547
rect 45961 55491 46029 55547
rect 46085 55491 46153 55547
rect 46209 55491 46277 55547
rect 46333 55491 46401 55547
rect 46457 55491 46525 55547
rect 46581 55491 46634 55547
rect 45634 55423 46634 55491
rect 45634 55367 45657 55423
rect 45713 55367 45781 55423
rect 45837 55367 45905 55423
rect 45961 55367 46029 55423
rect 46085 55367 46153 55423
rect 46209 55367 46277 55423
rect 46333 55367 46401 55423
rect 46457 55367 46525 55423
rect 46581 55367 46634 55423
rect 45634 55299 46634 55367
rect 45634 55243 45657 55299
rect 45713 55243 45781 55299
rect 45837 55243 45905 55299
rect 45961 55243 46029 55299
rect 46085 55243 46153 55299
rect 46209 55243 46277 55299
rect 46333 55243 46401 55299
rect 46457 55243 46525 55299
rect 46581 55243 46634 55299
rect 45634 55231 46634 55243
rect 50822 55039 51822 55839
rect 52386 55547 53386 55839
rect 52386 55491 52409 55547
rect 52465 55491 52533 55547
rect 52589 55491 52657 55547
rect 52713 55491 52781 55547
rect 52837 55491 52905 55547
rect 52961 55491 53029 55547
rect 53085 55491 53153 55547
rect 53209 55491 53277 55547
rect 53333 55491 53386 55547
rect 52386 55423 53386 55491
rect 52386 55367 52409 55423
rect 52465 55367 52533 55423
rect 52589 55367 52657 55423
rect 52713 55367 52781 55423
rect 52837 55367 52905 55423
rect 52961 55367 53029 55423
rect 53085 55367 53153 55423
rect 53209 55367 53277 55423
rect 53333 55367 53386 55423
rect 52386 55299 53386 55367
rect 52386 55243 52409 55299
rect 52465 55243 52533 55299
rect 52589 55243 52657 55299
rect 52713 55243 52781 55299
rect 52837 55243 52905 55299
rect 52961 55243 53029 55299
rect 53085 55243 53153 55299
rect 53209 55243 53277 55299
rect 53333 55243 53386 55299
rect 52386 55231 53386 55243
rect 54490 55039 55490 55839
rect 56183 55039 57183 55839
rect 57911 55547 58911 55839
rect 57911 55491 57934 55547
rect 57990 55491 58058 55547
rect 58114 55491 58182 55547
rect 58238 55491 58306 55547
rect 58362 55491 58430 55547
rect 58486 55491 58554 55547
rect 58610 55491 58678 55547
rect 58734 55491 58802 55547
rect 58858 55491 58911 55547
rect 57911 55423 58911 55491
rect 57911 55367 57934 55423
rect 57990 55367 58058 55423
rect 58114 55367 58182 55423
rect 58238 55367 58306 55423
rect 58362 55367 58430 55423
rect 58486 55367 58554 55423
rect 58610 55367 58678 55423
rect 58734 55367 58802 55423
rect 58858 55367 58911 55423
rect 57911 55299 58911 55367
rect 57911 55243 57934 55299
rect 57990 55243 58058 55299
rect 58114 55243 58182 55299
rect 58238 55243 58306 55299
rect 58362 55243 58430 55299
rect 58486 55243 58554 55299
rect 58610 55243 58678 55299
rect 58734 55243 58802 55299
rect 58858 55243 58911 55299
rect 57911 55231 58911 55243
rect 59468 55039 60468 55839
rect 60712 55547 61712 55839
rect 60712 55491 60735 55547
rect 60791 55491 60859 55547
rect 60915 55491 60983 55547
rect 61039 55491 61107 55547
rect 61163 55491 61231 55547
rect 61287 55491 61355 55547
rect 61411 55491 61479 55547
rect 61535 55491 61603 55547
rect 61659 55491 61712 55547
rect 60712 55423 61712 55491
rect 60712 55367 60735 55423
rect 60791 55367 60859 55423
rect 60915 55367 60983 55423
rect 61039 55367 61107 55423
rect 61163 55367 61231 55423
rect 61287 55367 61355 55423
rect 61411 55367 61479 55423
rect 61535 55367 61603 55423
rect 61659 55367 61712 55423
rect 60712 55299 61712 55367
rect 60712 55243 60735 55299
rect 60791 55243 60859 55299
rect 60915 55243 60983 55299
rect 61039 55243 61107 55299
rect 61163 55243 61231 55299
rect 61287 55243 61355 55299
rect 61411 55243 61479 55299
rect 61535 55243 61603 55299
rect 61659 55243 61712 55299
rect 60712 55231 61712 55243
rect 2203 55003 88293 55039
rect 2203 54998 31566 55003
rect 2203 54942 28533 54998
rect 28589 54942 28657 54998
rect 28713 54942 28781 54998
rect 28837 54942 28905 54998
rect 28961 54942 29029 54998
rect 29085 54942 29153 54998
rect 29209 54942 29277 54998
rect 29333 54942 29401 54998
rect 29457 54947 31566 54998
rect 31622 54947 31690 55003
rect 31746 54947 31814 55003
rect 31870 54947 31938 55003
rect 31994 54947 32062 55003
rect 32118 54947 32186 55003
rect 32242 54947 32310 55003
rect 32366 54947 32715 55003
rect 32771 54947 32839 55003
rect 32895 54947 32963 55003
rect 33019 54947 33087 55003
rect 33143 54947 33211 55003
rect 33267 54947 33335 55003
rect 33391 54947 33459 55003
rect 33515 54947 33850 55003
rect 33906 54947 33974 55003
rect 34030 54947 34098 55003
rect 34154 54947 34222 55003
rect 34278 54947 34346 55003
rect 34402 54947 34470 55003
rect 34526 54947 34594 55003
rect 34650 54984 88293 55003
rect 34650 54947 37087 54984
rect 29457 54942 37087 54947
rect 2203 54928 37087 54942
rect 37143 54928 37211 54984
rect 37267 54928 37335 54984
rect 37391 54928 37459 54984
rect 37515 54928 37583 54984
rect 37639 54928 37707 54984
rect 37763 54928 37831 54984
rect 37887 54928 37955 54984
rect 38011 54928 38079 54984
rect 38135 54928 38203 54984
rect 38259 54928 40544 54984
rect 40600 54928 40668 54984
rect 40724 54928 40792 54984
rect 40848 54928 40916 54984
rect 40972 54928 41040 54984
rect 41096 54928 41164 54984
rect 41220 54928 41288 54984
rect 41344 54928 41412 54984
rect 41468 54928 50860 54984
rect 50916 54928 50984 54984
rect 51040 54928 51108 54984
rect 51164 54928 51232 54984
rect 51288 54928 51356 54984
rect 51412 54928 51480 54984
rect 51536 54928 51604 54984
rect 51660 54928 51728 54984
rect 51784 54928 54528 54984
rect 54584 54928 54652 54984
rect 54708 54928 54776 54984
rect 54832 54928 54900 54984
rect 54956 54928 55024 54984
rect 55080 54928 55148 54984
rect 55204 54928 55272 54984
rect 55328 54928 55396 54984
rect 55452 54928 56221 54984
rect 56277 54928 56345 54984
rect 56401 54928 56469 54984
rect 56525 54928 56593 54984
rect 56649 54928 56717 54984
rect 56773 54928 56841 54984
rect 56897 54928 56965 54984
rect 57021 54928 57089 54984
rect 57145 54928 59506 54984
rect 59562 54928 59630 54984
rect 59686 54928 59754 54984
rect 59810 54928 59878 54984
rect 59934 54928 60002 54984
rect 60058 54928 60126 54984
rect 60182 54928 60250 54984
rect 60306 54928 60374 54984
rect 60430 54928 88293 54984
rect 2203 54879 88293 54928
rect 2203 54874 31566 54879
rect 2203 54818 28533 54874
rect 28589 54818 28657 54874
rect 28713 54818 28781 54874
rect 28837 54818 28905 54874
rect 28961 54818 29029 54874
rect 29085 54818 29153 54874
rect 29209 54818 29277 54874
rect 29333 54818 29401 54874
rect 29457 54823 31566 54874
rect 31622 54823 31690 54879
rect 31746 54823 31814 54879
rect 31870 54823 31938 54879
rect 31994 54823 32062 54879
rect 32118 54823 32186 54879
rect 32242 54823 32310 54879
rect 32366 54823 32715 54879
rect 32771 54823 32839 54879
rect 32895 54823 32963 54879
rect 33019 54823 33087 54879
rect 33143 54823 33211 54879
rect 33267 54823 33335 54879
rect 33391 54823 33459 54879
rect 33515 54823 33850 54879
rect 33906 54823 33974 54879
rect 34030 54823 34098 54879
rect 34154 54823 34222 54879
rect 34278 54823 34346 54879
rect 34402 54823 34470 54879
rect 34526 54823 34594 54879
rect 34650 54860 88293 54879
rect 34650 54823 37087 54860
rect 29457 54818 37087 54823
rect 2203 54804 37087 54818
rect 37143 54804 37211 54860
rect 37267 54804 37335 54860
rect 37391 54804 37459 54860
rect 37515 54804 37583 54860
rect 37639 54804 37707 54860
rect 37763 54804 37831 54860
rect 37887 54804 37955 54860
rect 38011 54804 38079 54860
rect 38135 54804 38203 54860
rect 38259 54804 40544 54860
rect 40600 54804 40668 54860
rect 40724 54804 40792 54860
rect 40848 54804 40916 54860
rect 40972 54804 41040 54860
rect 41096 54804 41164 54860
rect 41220 54804 41288 54860
rect 41344 54804 41412 54860
rect 41468 54804 50860 54860
rect 50916 54804 50984 54860
rect 51040 54804 51108 54860
rect 51164 54804 51232 54860
rect 51288 54804 51356 54860
rect 51412 54804 51480 54860
rect 51536 54804 51604 54860
rect 51660 54804 51728 54860
rect 51784 54804 54528 54860
rect 54584 54804 54652 54860
rect 54708 54804 54776 54860
rect 54832 54804 54900 54860
rect 54956 54804 55024 54860
rect 55080 54804 55148 54860
rect 55204 54804 55272 54860
rect 55328 54804 55396 54860
rect 55452 54804 56221 54860
rect 56277 54804 56345 54860
rect 56401 54804 56469 54860
rect 56525 54804 56593 54860
rect 56649 54804 56717 54860
rect 56773 54804 56841 54860
rect 56897 54804 56965 54860
rect 57021 54804 57089 54860
rect 57145 54804 59506 54860
rect 59562 54804 59630 54860
rect 59686 54804 59754 54860
rect 59810 54804 59878 54860
rect 59934 54804 60002 54860
rect 60058 54804 60126 54860
rect 60182 54804 60250 54860
rect 60306 54804 60374 54860
rect 60430 54804 88293 54860
rect 2203 54755 88293 54804
rect 2203 54750 31566 54755
rect 2203 54694 28533 54750
rect 28589 54694 28657 54750
rect 28713 54694 28781 54750
rect 28837 54694 28905 54750
rect 28961 54694 29029 54750
rect 29085 54694 29153 54750
rect 29209 54694 29277 54750
rect 29333 54694 29401 54750
rect 29457 54699 31566 54750
rect 31622 54699 31690 54755
rect 31746 54699 31814 54755
rect 31870 54699 31938 54755
rect 31994 54699 32062 54755
rect 32118 54699 32186 54755
rect 32242 54699 32310 54755
rect 32366 54699 32715 54755
rect 32771 54699 32839 54755
rect 32895 54699 32963 54755
rect 33019 54699 33087 54755
rect 33143 54699 33211 54755
rect 33267 54699 33335 54755
rect 33391 54699 33459 54755
rect 33515 54699 33850 54755
rect 33906 54699 33974 54755
rect 34030 54699 34098 54755
rect 34154 54699 34222 54755
rect 34278 54699 34346 54755
rect 34402 54699 34470 54755
rect 34526 54699 34594 54755
rect 34650 54736 88293 54755
rect 34650 54699 37087 54736
rect 29457 54694 37087 54699
rect 2203 54680 37087 54694
rect 37143 54680 37211 54736
rect 37267 54680 37335 54736
rect 37391 54680 37459 54736
rect 37515 54680 37583 54736
rect 37639 54680 37707 54736
rect 37763 54680 37831 54736
rect 37887 54680 37955 54736
rect 38011 54680 38079 54736
rect 38135 54680 38203 54736
rect 38259 54680 40544 54736
rect 40600 54680 40668 54736
rect 40724 54680 40792 54736
rect 40848 54680 40916 54736
rect 40972 54680 41040 54736
rect 41096 54680 41164 54736
rect 41220 54680 41288 54736
rect 41344 54680 41412 54736
rect 41468 54680 50860 54736
rect 50916 54680 50984 54736
rect 51040 54680 51108 54736
rect 51164 54680 51232 54736
rect 51288 54680 51356 54736
rect 51412 54680 51480 54736
rect 51536 54680 51604 54736
rect 51660 54680 51728 54736
rect 51784 54680 54528 54736
rect 54584 54680 54652 54736
rect 54708 54680 54776 54736
rect 54832 54680 54900 54736
rect 54956 54680 55024 54736
rect 55080 54680 55148 54736
rect 55204 54680 55272 54736
rect 55328 54680 55396 54736
rect 55452 54680 56221 54736
rect 56277 54680 56345 54736
rect 56401 54680 56469 54736
rect 56525 54680 56593 54736
rect 56649 54680 56717 54736
rect 56773 54680 56841 54736
rect 56897 54680 56965 54736
rect 57021 54680 57089 54736
rect 57145 54680 59506 54736
rect 59562 54680 59630 54736
rect 59686 54680 59754 54736
rect 59810 54680 59878 54736
rect 59934 54680 60002 54736
rect 60058 54680 60126 54736
rect 60182 54680 60250 54736
rect 60306 54680 60374 54736
rect 60430 54680 88293 54736
rect 2203 54631 88293 54680
rect 2203 54626 31566 54631
rect 2203 54570 28533 54626
rect 28589 54570 28657 54626
rect 28713 54570 28781 54626
rect 28837 54570 28905 54626
rect 28961 54570 29029 54626
rect 29085 54570 29153 54626
rect 29209 54570 29277 54626
rect 29333 54570 29401 54626
rect 29457 54575 31566 54626
rect 31622 54575 31690 54631
rect 31746 54575 31814 54631
rect 31870 54575 31938 54631
rect 31994 54575 32062 54631
rect 32118 54575 32186 54631
rect 32242 54575 32310 54631
rect 32366 54575 32715 54631
rect 32771 54575 32839 54631
rect 32895 54575 32963 54631
rect 33019 54575 33087 54631
rect 33143 54575 33211 54631
rect 33267 54575 33335 54631
rect 33391 54575 33459 54631
rect 33515 54575 33850 54631
rect 33906 54575 33974 54631
rect 34030 54575 34098 54631
rect 34154 54575 34222 54631
rect 34278 54575 34346 54631
rect 34402 54575 34470 54631
rect 34526 54575 34594 54631
rect 34650 54612 88293 54631
rect 34650 54575 37087 54612
rect 29457 54570 37087 54575
rect 2203 54556 37087 54570
rect 37143 54556 37211 54612
rect 37267 54556 37335 54612
rect 37391 54556 37459 54612
rect 37515 54556 37583 54612
rect 37639 54556 37707 54612
rect 37763 54556 37831 54612
rect 37887 54556 37955 54612
rect 38011 54556 38079 54612
rect 38135 54556 38203 54612
rect 38259 54556 40544 54612
rect 40600 54556 40668 54612
rect 40724 54556 40792 54612
rect 40848 54556 40916 54612
rect 40972 54556 41040 54612
rect 41096 54556 41164 54612
rect 41220 54556 41288 54612
rect 41344 54556 41412 54612
rect 41468 54556 50860 54612
rect 50916 54556 50984 54612
rect 51040 54556 51108 54612
rect 51164 54556 51232 54612
rect 51288 54556 51356 54612
rect 51412 54556 51480 54612
rect 51536 54556 51604 54612
rect 51660 54556 51728 54612
rect 51784 54556 54528 54612
rect 54584 54556 54652 54612
rect 54708 54556 54776 54612
rect 54832 54556 54900 54612
rect 54956 54556 55024 54612
rect 55080 54556 55148 54612
rect 55204 54556 55272 54612
rect 55328 54556 55396 54612
rect 55452 54556 56221 54612
rect 56277 54556 56345 54612
rect 56401 54556 56469 54612
rect 56525 54556 56593 54612
rect 56649 54556 56717 54612
rect 56773 54556 56841 54612
rect 56897 54556 56965 54612
rect 57021 54556 57089 54612
rect 57145 54556 59506 54612
rect 59562 54556 59630 54612
rect 59686 54556 59754 54612
rect 59810 54556 59878 54612
rect 59934 54556 60002 54612
rect 60058 54556 60126 54612
rect 60182 54556 60250 54612
rect 60306 54556 60374 54612
rect 60430 54556 88293 54612
rect 2203 54507 88293 54556
rect 2203 54502 31566 54507
rect 2203 54446 28533 54502
rect 28589 54446 28657 54502
rect 28713 54446 28781 54502
rect 28837 54446 28905 54502
rect 28961 54446 29029 54502
rect 29085 54446 29153 54502
rect 29209 54446 29277 54502
rect 29333 54446 29401 54502
rect 29457 54451 31566 54502
rect 31622 54451 31690 54507
rect 31746 54451 31814 54507
rect 31870 54451 31938 54507
rect 31994 54451 32062 54507
rect 32118 54451 32186 54507
rect 32242 54451 32310 54507
rect 32366 54451 32715 54507
rect 32771 54451 32839 54507
rect 32895 54451 32963 54507
rect 33019 54451 33087 54507
rect 33143 54451 33211 54507
rect 33267 54451 33335 54507
rect 33391 54451 33459 54507
rect 33515 54451 33850 54507
rect 33906 54451 33974 54507
rect 34030 54451 34098 54507
rect 34154 54451 34222 54507
rect 34278 54451 34346 54507
rect 34402 54451 34470 54507
rect 34526 54451 34594 54507
rect 34650 54488 88293 54507
rect 34650 54451 37087 54488
rect 29457 54446 37087 54451
rect 2203 54432 37087 54446
rect 37143 54432 37211 54488
rect 37267 54432 37335 54488
rect 37391 54432 37459 54488
rect 37515 54432 37583 54488
rect 37639 54432 37707 54488
rect 37763 54432 37831 54488
rect 37887 54432 37955 54488
rect 38011 54432 38079 54488
rect 38135 54432 38203 54488
rect 38259 54432 40544 54488
rect 40600 54432 40668 54488
rect 40724 54432 40792 54488
rect 40848 54432 40916 54488
rect 40972 54432 41040 54488
rect 41096 54432 41164 54488
rect 41220 54432 41288 54488
rect 41344 54432 41412 54488
rect 41468 54432 50860 54488
rect 50916 54432 50984 54488
rect 51040 54432 51108 54488
rect 51164 54432 51232 54488
rect 51288 54432 51356 54488
rect 51412 54432 51480 54488
rect 51536 54432 51604 54488
rect 51660 54432 51728 54488
rect 51784 54432 54528 54488
rect 54584 54432 54652 54488
rect 54708 54432 54776 54488
rect 54832 54432 54900 54488
rect 54956 54432 55024 54488
rect 55080 54432 55148 54488
rect 55204 54432 55272 54488
rect 55328 54432 55396 54488
rect 55452 54432 56221 54488
rect 56277 54432 56345 54488
rect 56401 54432 56469 54488
rect 56525 54432 56593 54488
rect 56649 54432 56717 54488
rect 56773 54432 56841 54488
rect 56897 54432 56965 54488
rect 57021 54432 57089 54488
rect 57145 54432 59506 54488
rect 59562 54432 59630 54488
rect 59686 54432 59754 54488
rect 59810 54432 59878 54488
rect 59934 54432 60002 54488
rect 60058 54432 60126 54488
rect 60182 54432 60250 54488
rect 60306 54432 60374 54488
rect 60430 54432 88293 54488
rect 2203 54383 88293 54432
rect 2203 54378 31566 54383
rect 2203 54322 28533 54378
rect 28589 54322 28657 54378
rect 28713 54322 28781 54378
rect 28837 54322 28905 54378
rect 28961 54322 29029 54378
rect 29085 54322 29153 54378
rect 29209 54322 29277 54378
rect 29333 54322 29401 54378
rect 29457 54327 31566 54378
rect 31622 54327 31690 54383
rect 31746 54327 31814 54383
rect 31870 54327 31938 54383
rect 31994 54327 32062 54383
rect 32118 54327 32186 54383
rect 32242 54327 32310 54383
rect 32366 54327 32715 54383
rect 32771 54327 32839 54383
rect 32895 54327 32963 54383
rect 33019 54327 33087 54383
rect 33143 54327 33211 54383
rect 33267 54327 33335 54383
rect 33391 54327 33459 54383
rect 33515 54327 33850 54383
rect 33906 54327 33974 54383
rect 34030 54327 34098 54383
rect 34154 54327 34222 54383
rect 34278 54327 34346 54383
rect 34402 54327 34470 54383
rect 34526 54327 34594 54383
rect 34650 54364 88293 54383
rect 34650 54327 37087 54364
rect 29457 54322 37087 54327
rect 2203 54308 37087 54322
rect 37143 54308 37211 54364
rect 37267 54308 37335 54364
rect 37391 54308 37459 54364
rect 37515 54308 37583 54364
rect 37639 54308 37707 54364
rect 37763 54308 37831 54364
rect 37887 54308 37955 54364
rect 38011 54308 38079 54364
rect 38135 54308 38203 54364
rect 38259 54308 40544 54364
rect 40600 54308 40668 54364
rect 40724 54308 40792 54364
rect 40848 54308 40916 54364
rect 40972 54308 41040 54364
rect 41096 54308 41164 54364
rect 41220 54308 41288 54364
rect 41344 54308 41412 54364
rect 41468 54308 50860 54364
rect 50916 54308 50984 54364
rect 51040 54308 51108 54364
rect 51164 54308 51232 54364
rect 51288 54308 51356 54364
rect 51412 54308 51480 54364
rect 51536 54308 51604 54364
rect 51660 54308 51728 54364
rect 51784 54308 54528 54364
rect 54584 54308 54652 54364
rect 54708 54308 54776 54364
rect 54832 54308 54900 54364
rect 54956 54308 55024 54364
rect 55080 54308 55148 54364
rect 55204 54308 55272 54364
rect 55328 54308 55396 54364
rect 55452 54308 56221 54364
rect 56277 54308 56345 54364
rect 56401 54308 56469 54364
rect 56525 54308 56593 54364
rect 56649 54308 56717 54364
rect 56773 54308 56841 54364
rect 56897 54308 56965 54364
rect 57021 54308 57089 54364
rect 57145 54308 59506 54364
rect 59562 54308 59630 54364
rect 59686 54308 59754 54364
rect 59810 54308 59878 54364
rect 59934 54308 60002 54364
rect 60058 54308 60126 54364
rect 60182 54308 60250 54364
rect 60306 54308 60374 54364
rect 60430 54308 88293 54364
rect 2203 54259 88293 54308
rect 2203 54254 31566 54259
rect 2203 54198 28533 54254
rect 28589 54198 28657 54254
rect 28713 54198 28781 54254
rect 28837 54198 28905 54254
rect 28961 54198 29029 54254
rect 29085 54198 29153 54254
rect 29209 54198 29277 54254
rect 29333 54198 29401 54254
rect 29457 54203 31566 54254
rect 31622 54203 31690 54259
rect 31746 54203 31814 54259
rect 31870 54203 31938 54259
rect 31994 54203 32062 54259
rect 32118 54203 32186 54259
rect 32242 54203 32310 54259
rect 32366 54203 32715 54259
rect 32771 54203 32839 54259
rect 32895 54203 32963 54259
rect 33019 54203 33087 54259
rect 33143 54203 33211 54259
rect 33267 54203 33335 54259
rect 33391 54203 33459 54259
rect 33515 54203 33850 54259
rect 33906 54203 33974 54259
rect 34030 54203 34098 54259
rect 34154 54203 34222 54259
rect 34278 54203 34346 54259
rect 34402 54203 34470 54259
rect 34526 54203 34594 54259
rect 34650 54240 88293 54259
rect 34650 54203 37087 54240
rect 29457 54198 37087 54203
rect 2203 54184 37087 54198
rect 37143 54184 37211 54240
rect 37267 54184 37335 54240
rect 37391 54184 37459 54240
rect 37515 54184 37583 54240
rect 37639 54184 37707 54240
rect 37763 54184 37831 54240
rect 37887 54184 37955 54240
rect 38011 54184 38079 54240
rect 38135 54184 38203 54240
rect 38259 54184 40544 54240
rect 40600 54184 40668 54240
rect 40724 54184 40792 54240
rect 40848 54184 40916 54240
rect 40972 54184 41040 54240
rect 41096 54184 41164 54240
rect 41220 54184 41288 54240
rect 41344 54184 41412 54240
rect 41468 54184 50860 54240
rect 50916 54184 50984 54240
rect 51040 54184 51108 54240
rect 51164 54184 51232 54240
rect 51288 54184 51356 54240
rect 51412 54184 51480 54240
rect 51536 54184 51604 54240
rect 51660 54184 51728 54240
rect 51784 54184 54528 54240
rect 54584 54184 54652 54240
rect 54708 54184 54776 54240
rect 54832 54184 54900 54240
rect 54956 54184 55024 54240
rect 55080 54184 55148 54240
rect 55204 54184 55272 54240
rect 55328 54184 55396 54240
rect 55452 54184 56221 54240
rect 56277 54184 56345 54240
rect 56401 54184 56469 54240
rect 56525 54184 56593 54240
rect 56649 54184 56717 54240
rect 56773 54184 56841 54240
rect 56897 54184 56965 54240
rect 57021 54184 57089 54240
rect 57145 54184 59506 54240
rect 59562 54184 59630 54240
rect 59686 54184 59754 54240
rect 59810 54184 59878 54240
rect 59934 54184 60002 54240
rect 60058 54184 60126 54240
rect 60182 54184 60250 54240
rect 60306 54184 60374 54240
rect 60430 54184 88293 54240
rect 2203 54135 88293 54184
rect 2203 54130 31566 54135
rect 2203 54074 28533 54130
rect 28589 54074 28657 54130
rect 28713 54074 28781 54130
rect 28837 54074 28905 54130
rect 28961 54074 29029 54130
rect 29085 54074 29153 54130
rect 29209 54074 29277 54130
rect 29333 54074 29401 54130
rect 29457 54079 31566 54130
rect 31622 54079 31690 54135
rect 31746 54079 31814 54135
rect 31870 54079 31938 54135
rect 31994 54079 32062 54135
rect 32118 54079 32186 54135
rect 32242 54079 32310 54135
rect 32366 54079 32715 54135
rect 32771 54079 32839 54135
rect 32895 54079 32963 54135
rect 33019 54079 33087 54135
rect 33143 54079 33211 54135
rect 33267 54079 33335 54135
rect 33391 54079 33459 54135
rect 33515 54079 33850 54135
rect 33906 54079 33974 54135
rect 34030 54079 34098 54135
rect 34154 54079 34222 54135
rect 34278 54079 34346 54135
rect 34402 54079 34470 54135
rect 34526 54079 34594 54135
rect 34650 54116 88293 54135
rect 34650 54079 37087 54116
rect 29457 54074 37087 54079
rect 2203 54060 37087 54074
rect 37143 54060 37211 54116
rect 37267 54060 37335 54116
rect 37391 54060 37459 54116
rect 37515 54060 37583 54116
rect 37639 54060 37707 54116
rect 37763 54060 37831 54116
rect 37887 54060 37955 54116
rect 38011 54060 38079 54116
rect 38135 54060 38203 54116
rect 38259 54060 40544 54116
rect 40600 54060 40668 54116
rect 40724 54060 40792 54116
rect 40848 54060 40916 54116
rect 40972 54060 41040 54116
rect 41096 54060 41164 54116
rect 41220 54060 41288 54116
rect 41344 54060 41412 54116
rect 41468 54060 50860 54116
rect 50916 54060 50984 54116
rect 51040 54060 51108 54116
rect 51164 54060 51232 54116
rect 51288 54060 51356 54116
rect 51412 54060 51480 54116
rect 51536 54060 51604 54116
rect 51660 54060 51728 54116
rect 51784 54060 54528 54116
rect 54584 54060 54652 54116
rect 54708 54060 54776 54116
rect 54832 54060 54900 54116
rect 54956 54060 55024 54116
rect 55080 54060 55148 54116
rect 55204 54060 55272 54116
rect 55328 54060 55396 54116
rect 55452 54060 56221 54116
rect 56277 54060 56345 54116
rect 56401 54060 56469 54116
rect 56525 54060 56593 54116
rect 56649 54060 56717 54116
rect 56773 54060 56841 54116
rect 56897 54060 56965 54116
rect 57021 54060 57089 54116
rect 57145 54060 59506 54116
rect 59562 54060 59630 54116
rect 59686 54060 59754 54116
rect 59810 54060 59878 54116
rect 59934 54060 60002 54116
rect 60058 54060 60126 54116
rect 60182 54060 60250 54116
rect 60306 54060 60374 54116
rect 60430 54060 88293 54116
rect 2203 54039 88293 54060
rect 28753 4282 29077 4292
rect 28753 4226 28763 4282
rect 28819 4226 28887 4282
rect 28943 4226 29011 4282
rect 29067 4226 29077 4282
rect 28753 4158 29077 4226
rect 28753 4102 28763 4158
rect 28819 4102 28887 4158
rect 28943 4102 29011 4158
rect 29067 4102 29077 4158
rect 28753 4034 29077 4102
rect 28753 3978 28763 4034
rect 28819 3978 28887 4034
rect 28943 3978 29011 4034
rect 29067 3978 29077 4034
rect 28753 3910 29077 3978
rect 28753 3854 28763 3910
rect 28819 3854 28887 3910
rect 28943 3854 29011 3910
rect 29067 3854 29077 3910
rect 28753 3786 29077 3854
rect 28753 3730 28763 3786
rect 28819 3730 28887 3786
rect 28943 3730 29011 3786
rect 29067 3730 29077 3786
rect 28753 3662 29077 3730
rect 28753 3606 28763 3662
rect 28819 3606 28887 3662
rect 28943 3606 29011 3662
rect 29067 3606 29077 3662
rect 28753 3538 29077 3606
rect 28753 3482 28763 3538
rect 28819 3482 28887 3538
rect 28943 3482 29011 3538
rect 29067 3482 29077 3538
rect 28753 3414 29077 3482
rect 28753 3358 28763 3414
rect 28819 3358 28887 3414
rect 28943 3358 29011 3414
rect 29067 3358 29077 3414
rect 28753 3348 29077 3358
rect 59890 4282 60214 4292
rect 59890 4226 59900 4282
rect 59956 4226 60024 4282
rect 60080 4226 60148 4282
rect 60204 4226 60214 4282
rect 59890 4158 60214 4226
rect 59890 4102 59900 4158
rect 59956 4102 60024 4158
rect 60080 4102 60148 4158
rect 60204 4102 60214 4158
rect 59890 4034 60214 4102
rect 59890 3978 59900 4034
rect 59956 3978 60024 4034
rect 60080 3978 60148 4034
rect 60204 3978 60214 4034
rect 59890 3910 60214 3978
rect 59890 3854 59900 3910
rect 59956 3854 60024 3910
rect 60080 3854 60148 3910
rect 60204 3854 60214 3910
rect 59890 3786 60214 3854
rect 59890 3730 59900 3786
rect 59956 3730 60024 3786
rect 60080 3730 60148 3786
rect 60204 3730 60214 3786
rect 59890 3662 60214 3730
rect 59890 3606 59900 3662
rect 59956 3606 60024 3662
rect 60080 3606 60148 3662
rect 60204 3606 60214 3662
rect 59890 3538 60214 3606
rect 59890 3482 59900 3538
rect 59956 3482 60024 3538
rect 60080 3482 60148 3538
rect 60204 3482 60214 3538
rect 59890 3414 60214 3482
rect 59890 3358 59900 3414
rect 59956 3358 60024 3414
rect 60080 3358 60148 3414
rect 60204 3358 60214 3414
rect 59890 3348 60214 3358
use M2_M14310590548777_128x8m81  M2_M14310590548777_128x8m81_0
timestamp 1698431365
transform 1 0 59432 0 1 3583
box 0 0 1 1
use M2_M14310590548778_128x8m81  M2_M14310590548778_128x8m81_0
timestamp 1698431365
transform 1 0 60052 0 1 4068
box 0 0 1 1
use M2_M14310590548778_128x8m81  M2_M14310590548778_128x8m81_1
timestamp 1698431365
transform 1 0 28915 0 1 4068
box 0 0 1 1
use M2_M14310590548782_128x8m81  M2_M14310590548782_128x8m81_0
timestamp 1698431365
transform 1 0 29524 0 1 3317
box 0 0 1 1
use M2_M14310590548783_128x8m81  M2_M14310590548783_128x8m81_0
timestamp 1698431365
transform 1 0 27590 0 1 55395
box 0 0 1 1
use M2_M14310590548783_128x8m81  M2_M14310590548783_128x8m81_1
timestamp 1698431365
transform 1 0 46119 0 1 55395
box 0 0 1 1
use M2_M14310590548783_128x8m81  M2_M14310590548783_128x8m81_2
timestamp 1698431365
transform 1 0 36446 0 1 55395
box 0 0 1 1
use M2_M14310590548783_128x8m81  M2_M14310590548783_128x8m81_3
timestamp 1698431365
transform 1 0 42288 0 1 55395
box 0 0 1 1
use M2_M14310590548783_128x8m81  M2_M14310590548783_128x8m81_4
timestamp 1698431365
transform 1 0 61197 0 1 55395
box 0 0 1 1
use M2_M14310590548783_128x8m81  M2_M14310590548783_128x8m81_5
timestamp 1698431365
transform 1 0 52871 0 1 55395
box 0 0 1 1
use M2_M14310590548783_128x8m81  M2_M14310590548783_128x8m81_6
timestamp 1698431365
transform 1 0 58396 0 1 55395
box 0 0 1 1
use M3_M2431059054879_128x8m81  M3_M2431059054879_128x8m81_0
timestamp 1698431365
transform 1 0 60052 0 1 3820
box 0 0 1 1
use M3_M2431059054879_128x8m81  M3_M2431059054879_128x8m81_1
timestamp 1698431365
transform 1 0 28915 0 1 3820
box 0 0 1 1
use M3_M24310590548776_128x8m81  M3_M24310590548776_128x8m81_0
timestamp 1698431365
transform 1 0 46119 0 1 55395
box 0 0 1 1
use M3_M24310590548776_128x8m81  M3_M24310590548776_128x8m81_1
timestamp 1698431365
transform 1 0 61197 0 1 55395
box 0 0 1 1
use M3_M24310590548776_128x8m81  M3_M24310590548776_128x8m81_2
timestamp 1698431365
transform 1 0 36446 0 1 55395
box 0 0 1 1
use M3_M24310590548776_128x8m81  M3_M24310590548776_128x8m81_3
timestamp 1698431365
transform 1 0 42288 0 1 55395
box 0 0 1 1
use M3_M24310590548776_128x8m81  M3_M24310590548776_128x8m81_4
timestamp 1698431365
transform 1 0 52871 0 1 55395
box 0 0 1 1
use M3_M24310590548776_128x8m81  M3_M24310590548776_128x8m81_5
timestamp 1698431365
transform 1 0 58396 0 1 55395
box 0 0 1 1
use M3_M24310590548776_128x8m81  M3_M24310590548776_128x8m81_6
timestamp 1698431365
transform 1 0 27590 0 1 55395
box 0 0 1 1
use M3_M24310590548779_128x8m81  M3_M24310590548779_128x8m81_0
timestamp 1698431365
transform 1 0 37673 0 1 54522
box 0 0 1 1
use M3_M24310590548780_128x8m81  M3_M24310590548780_128x8m81_0
timestamp 1698431365
transform 1 0 34250 0 1 54541
box 0 0 1 1
use M3_M24310590548780_128x8m81  M3_M24310590548780_128x8m81_1
timestamp 1698431365
transform 1 0 31966 0 1 54541
box 0 0 1 1
use M3_M24310590548780_128x8m81  M3_M24310590548780_128x8m81_2
timestamp 1698431365
transform 1 0 33115 0 1 54541
box 0 0 1 1
use M3_M24310590548781_128x8m81  M3_M24310590548781_128x8m81_0
timestamp 1698431365
transform 1 0 56683 0 1 54522
box 0 0 1 1
use M3_M24310590548781_128x8m81  M3_M24310590548781_128x8m81_1
timestamp 1698431365
transform 1 0 28995 0 1 54536
box 0 0 1 1
use M3_M24310590548781_128x8m81  M3_M24310590548781_128x8m81_2
timestamp 1698431365
transform 1 0 59968 0 1 54522
box 0 0 1 1
use M3_M24310590548781_128x8m81  M3_M24310590548781_128x8m81_3
timestamp 1698431365
transform 1 0 51322 0 1 54522
box 0 0 1 1
use M3_M24310590548781_128x8m81  M3_M24310590548781_128x8m81_4
timestamp 1698431365
transform 1 0 54990 0 1 54522
box 0 0 1 1
use M3_M24310590548781_128x8m81  M3_M24310590548781_128x8m81_5
timestamp 1698431365
transform 1 0 41006 0 1 54522
box 0 0 1 1
use M3_M24310590548784_128x8m81  M3_M24310590548784_128x8m81_0
timestamp 1698431365
transform 1 0 60052 0 1 4068
box 0 0 1 1
use M3_M24310590548784_128x8m81  M3_M24310590548784_128x8m81_1
timestamp 1698431365
transform 1 0 28915 0 1 4068
box 0 0 1 1
use power_route_01_128x8m81  power_route_01_128x8m81_0
timestamp 1698431365
transform -1 0 85469 0 1 53414
box -511 0 1714 2425
use power_route_01_128x8m81  power_route_01_128x8m81_1
timestamp 1698431365
transform -1 0 25893 0 1 53414
box -511 0 1714 2425
use power_route_01_128x8m81  power_route_01_128x8m81_2
timestamp 1698431365
transform 1 0 9233 0 1 53414
box -511 0 1714 2425
use power_route_01_128x8m81  power_route_01_128x8m81_3
timestamp 1698431365
transform 1 0 20033 0 1 53414
box -511 0 1714 2425
use power_route_01_128x8m81  power_route_01_128x8m81_4
timestamp 1698431365
transform 1 0 14633 0 1 53414
box -511 0 1714 2425
use power_route_01_128x8m81  power_route_01_128x8m81_5
timestamp 1698431365
transform 1 0 63409 0 1 53414
box -511 0 1714 2425
use power_route_01_128x8m81  power_route_01_128x8m81_6
timestamp 1698431365
transform 1 0 79609 0 1 53414
box -511 0 1714 2425
use power_route_01_128x8m81  power_route_01_128x8m81_7
timestamp 1698431365
transform 1 0 74209 0 1 53414
box -511 0 1714 2425
use power_route_01_128x8m81  power_route_01_128x8m81_8
timestamp 1698431365
transform 1 0 68809 0 1 53414
box -511 0 1714 2425
use power_route_01_128x8m81  power_route_01_128x8m81_9
timestamp 1698431365
transform 1 0 3833 0 1 53414
box -511 0 1714 2425
use power_route_02_a_128x8m81  power_route_02_a_128x8m81_0
timestamp 1698431365
transform 1 0 -1418 0 1 50689
box 3339 -250 30611 1350
use power_route_02_a_128x8m81  power_route_02_a_128x8m81_1
timestamp 1698431365
transform 1 0 -1418 0 1 47089
box 3339 -250 30611 1350
use power_route_02_a_128x8m81  power_route_02_a_128x8m81_2
timestamp 1698431365
transform 1 0 -1418 0 1 48889
box 3339 -250 30611 1350
use power_route_02_a_128x8m81  power_route_02_a_128x8m81_3
timestamp 1698431365
transform 1 0 -1418 0 1 39889
box 3339 -250 30611 1350
use power_route_02_a_128x8m81  power_route_02_a_128x8m81_4
timestamp 1698431365
transform 1 0 -1418 0 1 41689
box 3339 -250 30611 1350
use power_route_02_a_128x8m81  power_route_02_a_128x8m81_5
timestamp 1698431365
transform 1 0 -1418 0 1 45289
box 3339 -250 30611 1350
use power_route_02_a_128x8m81  power_route_02_a_128x8m81_6
timestamp 1698431365
transform 1 0 -1418 0 1 43489
box 3339 -250 30611 1350
use power_route_02_a_128x8m81  power_route_02_a_128x8m81_7
timestamp 1698431365
transform 1 0 -1418 0 1 38089
box 3339 -250 30611 1350
use power_route_02_a_128x8m81  power_route_02_a_128x8m81_8
timestamp 1698431365
transform 1 0 -1418 0 1 52489
box 3339 -250 30611 1350
use power_route_02_b_128x8m81  power_route_02_b_128x8m81_0
timestamp 1698431365
transform -1 0 91632 0 1 39889
box 3339 -250 30290 1350
use power_route_02_b_128x8m81  power_route_02_b_128x8m81_1
timestamp 1698431365
transform -1 0 91632 0 1 41689
box 3339 -250 30290 1350
use power_route_02_b_128x8m81  power_route_02_b_128x8m81_2
timestamp 1698431365
transform -1 0 91632 0 1 43489
box 3339 -250 30290 1350
use power_route_02_b_128x8m81  power_route_02_b_128x8m81_3
timestamp 1698431365
transform -1 0 91632 0 1 45289
box 3339 -250 30290 1350
use power_route_02_b_128x8m81  power_route_02_b_128x8m81_4
timestamp 1698431365
transform -1 0 91632 0 1 47089
box 3339 -250 30290 1350
use power_route_02_b_128x8m81  power_route_02_b_128x8m81_5
timestamp 1698431365
transform -1 0 91632 0 1 48889
box 3339 -250 30290 1350
use power_route_02_b_128x8m81  power_route_02_b_128x8m81_6
timestamp 1698431365
transform -1 0 91632 0 1 50689
box 3339 -250 30290 1350
use power_route_02_b_128x8m81  power_route_02_b_128x8m81_7
timestamp 1698431365
transform -1 0 91632 0 1 52489
box 3339 -250 30290 1350
use power_route_02_b_128x8m81  power_route_02_b_128x8m81_8
timestamp 1698431365
transform -1 0 91632 0 1 38089
box 3339 -250 30290 1350
use power_route_04_128x8m81  power_route_04_128x8m81_0
timestamp 1698431365
transform -1 0 91632 0 1 244
box 3339 2101 6632 52645
use power_route_04_128x8m81  power_route_04_128x8m81_1
timestamp 1698431365
transform 1 0 -1418 0 1 244
box 3339 2101 6632 52645
use power_route_05_128x8m81  power_route_05_128x8m81_0
timestamp 1698431365
transform 1 0 19656 0 1 230
box -8 2115 1235 7462
use power_route_05_128x8m81  power_route_05_128x8m81_1
timestamp 1698431365
transform 1 0 68432 0 1 230
box -8 2115 1235 7462
use power_route_05_128x8m81  power_route_05_128x8m81_2
timestamp 1698431365
transform 1 0 79232 0 1 230
box -8 2115 1235 7462
use power_route_05_128x8m81  power_route_05_128x8m81_3
timestamp 1698431365
transform 1 0 8856 0 1 230
box -8 2115 1235 7462
use power_route_06_128x8m81  power_route_06_128x8m81_0
timestamp 1698431365
transform 1 0 61241 0 1 230
box -7 2115 1234 18431
use power_route_06_128x8m81  power_route_06_128x8m81_1
timestamp 1698431365
transform 1 0 26784 0 1 230
box -7 2115 1234 18431
use power_route_07_128x8m81  power_route_07_128x8m81_0
timestamp 1698431365
transform 1 0 40746 0 1 230
box -8 3065 1235 7462
use power_route_07_128x8m81  power_route_07_128x8m81_1
timestamp 1698431365
transform 1 0 38926 0 1 230
box -8 3065 1235 7462
<< properties >>
string GDS_END 2287280
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 2281564
string path 274.950 279.195 274.950 270.195 
<< end >>
