magic
tech gf180mcuB
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 453 2550 1094
<< pwell >>
rect -86 -86 2550 453
<< mvnmos >>
rect 124 69 244 279
rect 348 69 468 279
rect 572 69 692 279
rect 796 69 916 279
rect 1020 69 1140 279
rect 1244 69 1364 279
rect 1504 69 1624 333
rect 1728 69 1848 333
rect 1952 69 2072 333
rect 2176 69 2296 333
<< mvpmos >>
rect 144 573 244 939
rect 358 573 458 939
rect 582 573 682 939
rect 806 573 906 939
rect 1030 573 1130 939
rect 1244 573 1344 939
rect 1524 573 1624 939
rect 1738 573 1838 939
rect 1962 573 2062 939
rect 2176 573 2276 939
<< mvndiff >>
rect 1424 279 1504 333
rect 36 266 124 279
rect 36 126 49 266
rect 95 126 124 266
rect 36 69 124 126
rect 244 193 348 279
rect 244 147 273 193
rect 319 147 348 193
rect 244 69 348 147
rect 468 172 572 279
rect 468 126 497 172
rect 543 126 572 172
rect 468 69 572 126
rect 692 193 796 279
rect 692 147 721 193
rect 767 147 796 193
rect 692 69 796 147
rect 916 172 1020 279
rect 916 126 945 172
rect 991 126 1020 172
rect 916 69 1020 126
rect 1140 193 1244 279
rect 1140 147 1169 193
rect 1215 147 1244 193
rect 1140 69 1244 147
rect 1364 172 1504 279
rect 1364 126 1393 172
rect 1439 126 1504 172
rect 1364 69 1504 126
rect 1624 287 1728 333
rect 1624 147 1653 287
rect 1699 147 1728 287
rect 1624 69 1728 147
rect 1848 172 1952 333
rect 1848 126 1877 172
rect 1923 126 1952 172
rect 1848 69 1952 126
rect 2072 287 2176 333
rect 2072 147 2101 287
rect 2147 147 2176 287
rect 2072 69 2176 147
rect 2296 266 2384 333
rect 2296 126 2325 266
rect 2371 126 2384 266
rect 2296 69 2384 126
<< mvpdiff >>
rect 56 923 144 939
rect 56 783 69 923
rect 115 783 144 923
rect 56 573 144 783
rect 244 573 358 939
rect 458 573 582 939
rect 682 861 806 939
rect 682 721 731 861
rect 777 721 806 861
rect 682 573 806 721
rect 906 573 1030 939
rect 1130 573 1244 939
rect 1344 923 1524 939
rect 1344 783 1373 923
rect 1419 783 1524 923
rect 1344 573 1524 783
rect 1624 861 1738 939
rect 1624 721 1663 861
rect 1709 721 1738 861
rect 1624 573 1738 721
rect 1838 923 1962 939
rect 1838 783 1867 923
rect 1913 783 1962 923
rect 1838 573 1962 783
rect 2062 861 2176 939
rect 2062 721 2091 861
rect 2137 721 2176 861
rect 2062 573 2176 721
rect 2276 923 2364 939
rect 2276 783 2305 923
rect 2351 783 2364 923
rect 2276 573 2364 783
<< mvndiffc >>
rect 49 126 95 266
rect 273 147 319 193
rect 497 126 543 172
rect 721 147 767 193
rect 945 126 991 172
rect 1169 147 1215 193
rect 1393 126 1439 172
rect 1653 147 1699 287
rect 1877 126 1923 172
rect 2101 147 2147 287
rect 2325 126 2371 266
<< mvpdiffc >>
rect 69 783 115 923
rect 731 721 777 861
rect 1373 783 1419 923
rect 1663 721 1709 861
rect 1867 783 1913 923
rect 2091 721 2137 861
rect 2305 783 2351 923
<< polysilicon >>
rect 144 939 244 983
rect 358 939 458 983
rect 582 939 682 983
rect 806 939 906 983
rect 1030 939 1130 983
rect 1244 939 1344 983
rect 1524 939 1624 983
rect 1738 939 1838 983
rect 1962 939 2062 983
rect 2176 939 2276 983
rect 144 500 244 573
rect 144 454 157 500
rect 203 454 244 500
rect 144 323 244 454
rect 358 500 458 573
rect 358 454 377 500
rect 423 454 458 500
rect 358 323 458 454
rect 582 513 682 573
rect 806 513 906 573
rect 582 500 906 513
rect 582 454 595 500
rect 641 454 906 500
rect 582 441 906 454
rect 582 323 692 441
rect 124 279 244 323
rect 348 279 468 323
rect 572 279 692 323
rect 796 323 906 441
rect 1030 500 1130 573
rect 1030 454 1043 500
rect 1089 454 1130 500
rect 1030 323 1130 454
rect 1244 500 1344 573
rect 1244 454 1257 500
rect 1303 454 1344 500
rect 1244 323 1344 454
rect 1524 513 1624 573
rect 1738 513 1838 573
rect 1962 513 2062 573
rect 2176 513 2276 573
rect 1524 500 2276 513
rect 1524 454 1653 500
rect 1699 454 1877 500
rect 1923 454 2276 500
rect 1524 441 2276 454
rect 1524 377 1624 441
rect 1504 333 1624 377
rect 1728 333 1848 441
rect 1952 333 2072 441
rect 2176 377 2276 441
rect 2176 333 2296 377
rect 796 279 916 323
rect 1020 279 1140 323
rect 1244 279 1364 323
rect 124 25 244 69
rect 348 25 468 69
rect 572 25 692 69
rect 796 25 916 69
rect 1020 25 1140 69
rect 1244 25 1364 69
rect 1504 25 1624 69
rect 1728 25 1848 69
rect 1952 25 2072 69
rect 2176 25 2296 69
<< polycontact >>
rect 157 454 203 500
rect 377 454 423 500
rect 595 454 641 500
rect 1043 454 1089 500
rect 1257 454 1303 500
rect 1653 454 1699 500
rect 1877 454 1923 500
<< metal1 >>
rect 0 923 2464 1098
rect 0 918 69 923
rect 115 918 1373 923
rect 69 772 115 783
rect 731 861 777 872
rect 1419 918 1867 923
rect 1373 772 1419 783
rect 1663 861 1709 872
rect 777 721 1406 726
rect 731 680 1406 721
rect 1913 918 2305 923
rect 1867 772 1913 783
rect 2091 861 2137 872
rect 1709 721 2091 726
rect 2351 918 2464 923
rect 2305 772 2351 783
rect 1663 680 2137 721
rect 142 588 1314 634
rect 142 500 214 588
rect 584 500 652 542
rect 1246 500 1314 588
rect 142 454 157 500
rect 203 454 214 500
rect 366 454 377 500
rect 423 454 434 500
rect 584 454 595 500
rect 641 454 652 500
rect 698 454 1043 500
rect 1089 454 1100 500
rect 1246 454 1257 500
rect 1303 454 1314 500
rect 1360 500 1406 680
rect 1360 454 1653 500
rect 1699 454 1877 500
rect 1923 454 1934 500
rect 366 400 434 454
rect 698 400 744 454
rect 366 354 744 400
rect 49 266 95 277
rect 1360 275 1406 454
rect 1980 318 2026 680
rect 273 229 1406 275
rect 1653 298 2026 318
rect 1653 287 2147 298
rect 273 193 319 229
rect 721 193 767 229
rect 273 136 319 147
rect 497 172 543 183
rect 49 90 95 126
rect 1169 193 1215 229
rect 721 136 767 147
rect 945 172 991 183
rect 497 90 543 126
rect 1169 136 1215 147
rect 1393 172 1439 183
rect 945 90 991 126
rect 1699 242 2101 287
rect 1653 136 1699 147
rect 1877 172 1923 183
rect 1393 90 1439 126
rect 2101 136 2147 147
rect 2325 266 2371 277
rect 1877 90 1923 126
rect 2325 90 2371 126
rect 0 -90 2464 90
<< labels >>
flabel metal1 s 584 454 652 542 0 FreeSans 200 0 0 0 A1
port 1 nsew default input
flabel metal1 s 698 454 1100 500 0 FreeSans 200 0 0 0 A2
port 2 nsew default input
flabel metal1 s 142 588 1314 634 0 FreeSans 200 0 0 0 A3
port 3 nsew default input
flabel metal1 s 0 918 2464 1098 0 FreeSans 200 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 2325 183 2371 277 0 FreeSans 200 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel metal1 s 2091 726 2137 872 0 FreeSans 200 0 0 0 Z
port 4 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 6 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 366 454 434 500 1 A2
port 2 nsew default input
rlabel metal1 s 698 400 744 454 1 A2
port 2 nsew default input
rlabel metal1 s 366 400 434 454 1 A2
port 2 nsew default input
rlabel metal1 s 366 354 744 400 1 A2
port 2 nsew default input
rlabel metal1 s 1246 454 1314 588 1 A3
port 3 nsew default input
rlabel metal1 s 142 454 214 588 1 A3
port 3 nsew default input
rlabel metal1 s 1663 726 1709 872 1 Z
port 4 nsew default output
rlabel metal1 s 1663 680 2137 726 1 Z
port 4 nsew default output
rlabel metal1 s 1980 318 2026 680 1 Z
port 4 nsew default output
rlabel metal1 s 1653 298 2026 318 1 Z
port 4 nsew default output
rlabel metal1 s 1653 242 2147 298 1 Z
port 4 nsew default output
rlabel metal1 s 2101 136 2147 242 1 Z
port 4 nsew default output
rlabel metal1 s 1653 136 1699 242 1 Z
port 4 nsew default output
rlabel metal1 s 2305 772 2351 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1867 772 1913 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1373 772 1419 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 69 772 115 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 49 183 95 277 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2325 90 2371 183 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1877 90 1923 183 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1393 90 1439 183 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 945 90 991 183 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 497 90 543 183 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 49 90 95 183 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 2464 90 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2464 1008
string GDS_END 288486
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 282820
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
