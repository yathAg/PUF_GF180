magic
tech gf180mcuA
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 352 2326 870
<< pwell >>
rect -86 -86 2326 352
<< metal1 >>
rect 0 724 2240 844
rect 253 532 299 724
rect 354 424 430 550
rect 165 360 430 424
rect 697 617 743 724
rect 273 60 319 163
rect 670 248 886 312
rect 677 60 723 165
rect 800 110 886 248
rect 1553 531 1599 724
rect 1553 60 1599 179
rect 1921 106 1992 676
rect 2125 506 2171 724
rect 2145 60 2191 232
rect 0 -60 2240 60
<< obsm1 >>
rect 38 278 106 678
rect 522 417 579 678
rect 1020 628 1301 674
rect 625 467 1020 513
rect 1151 417 1197 562
rect 522 371 1197 417
rect 38 232 472 278
rect 38 106 106 232
rect 522 106 590 371
rect 957 202 1003 371
rect 1255 295 1301 628
rect 1757 461 1807 645
rect 1405 415 1834 461
rect 1255 249 1716 295
rect 1255 152 1301 249
rect 1040 106 1301 152
rect 1766 106 1834 415
<< labels >>
rlabel metal1 s 800 110 886 248 6 D
port 1 nsew default input
rlabel metal1 s 670 248 886 312 6 D
port 1 nsew default input
rlabel metal1 s 165 360 430 424 6 E
port 2 nsew clock input
rlabel metal1 s 354 424 430 550 6 E
port 2 nsew clock input
rlabel metal1 s 1921 106 1992 676 6 Q
port 3 nsew default output
rlabel metal1 s 2125 506 2171 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1553 531 1599 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 697 617 743 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 253 532 299 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 724 2240 844 6 VDD
port 4 nsew power bidirectional abutment
rlabel nwell s -86 352 2326 870 6 VNW
port 5 nsew power bidirectional
rlabel pwell s -86 -86 2326 352 6 VPW
port 6 nsew ground bidirectional
rlabel metal1 s 0 -60 2240 60 8 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2145 60 2191 232 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1553 60 1599 179 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 677 60 723 165 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 60 319 163 6 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2240 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 585744
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 580238
<< end >>
