magic
tech gf180mcuD
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 453 758 1094
<< pwell >>
rect -86 -86 758 453
<< metal1 >>
rect 0 918 672 1098
rect 49 710 95 918
rect 279 766 325 872
rect 279 690 474 766
rect 520 710 566 918
rect 126 454 382 542
rect 428 370 474 690
rect 366 334 474 370
rect 366 298 457 334
rect 49 90 95 298
rect 279 242 457 298
rect 279 136 325 242
rect 503 90 549 298
rect 0 -90 672 90
<< labels >>
rlabel metal1 s 126 454 382 542 6 I
port 1 nsew default input
rlabel metal1 s 279 136 325 242 6 ZN
port 2 nsew default output
rlabel metal1 s 279 242 457 298 6 ZN
port 2 nsew default output
rlabel metal1 s 366 298 457 334 6 ZN
port 2 nsew default output
rlabel metal1 s 366 334 474 370 6 ZN
port 2 nsew default output
rlabel metal1 s 428 370 474 690 6 ZN
port 2 nsew default output
rlabel metal1 s 279 690 474 766 6 ZN
port 2 nsew default output
rlabel metal1 s 279 766 325 872 6 ZN
port 2 nsew default output
rlabel metal1 s 520 710 566 918 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 710 95 918 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 918 672 1098 6 VDD
port 3 nsew power bidirectional abutment
rlabel nwell s -86 453 758 1094 6 VNW
port 4 nsew power bidirectional
rlabel pwell s -86 -86 758 453 6 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 0 -90 672 90 8 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 503 90 549 298 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 49 90 95 298 6 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 672 1008
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 874092
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 871222
<< end >>
