************************************************************************
* auCdl Netlist:
* 
* Library Name:  TCG_Library
* Top Cell Name: rm1
* View Name:     schematic
* Netlisted on:  Nov 24 10:16:24 2021
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: TCG_Library
* Cell Name:    rm1
* View Name:    schematic
************************************************************************

.SUBCKT rm1 I1_0_0_R0_MINUS I1_0_0_R0_PLUS I1_0_1_R0_MINUS I1_0_1_R0_PLUS 
+ I1_0_2_R0_MINUS I1_0_2_R0_PLUS I1_1_0_R0_MINUS I1_1_0_R0_PLUS 
+ I1_1_1_R0_MINUS I1_1_1_R0_PLUS I1_1_2_R0_MINUS I1_1_2_R0_PLUS 
+ I1_2_0_R0_MINUS I1_2_0_R0_PLUS I1_2_1_R0_MINUS I1_2_1_R0_PLUS 
+ I1_2_2_R0_MINUS I1_2_2_R0_PLUS I1_default_MINUS I1_default_PLUS
*.PININFO I1_0_0_R0_MINUS:I I1_0_0_R0_PLUS:I I1_0_1_R0_MINUS:I 
*.PININFO I1_0_1_R0_PLUS:I I1_0_2_R0_MINUS:I I1_0_2_R0_PLUS:I 
*.PININFO I1_1_0_R0_MINUS:I I1_1_0_R0_PLUS:I I1_1_1_R0_MINUS:I 
*.PININFO I1_1_1_R0_PLUS:I I1_1_2_R0_MINUS:I I1_1_2_R0_PLUS:I 
*.PININFO I1_2_0_R0_MINUS:I I1_2_0_R0_PLUS:I I1_2_1_R0_MINUS:I 
*.PININFO I1_2_1_R0_PLUS:I I1_2_2_R0_MINUS:I I1_2_2_R0_PLUS:I 
*.PININFO I1_default_MINUS:I I1_default_PLUS:I
RI1_2_2_R0 I1_2_2_R0_PLUS I1_2_2_R0_MINUS rm1 W=50u L=50u m=1 r=90m 
+ dtemp=0
RI1_2_1_R0 I1_2_1_R0_PLUS I1_2_1_R0_MINUS rm1 W=50u L=13.5u m=1 r=24.3m 
+ dtemp=0
RI1_2_0_R0 I1_2_0_R0_PLUS I1_2_0_R0_MINUS rm1 W=50u L=230n m=1 r=414u 
+ dtemp=0
RI1_1_2_R0 I1_1_2_R0_PLUS I1_1_2_R0_MINUS rm1 W=13.5u L=50u m=1 
+ r=333.333m dtemp=0
RI1_1_1_R0 I1_1_1_R0_PLUS I1_1_1_R0_MINUS rm1 W=13.5u L=13.5u m=1 r=90m 
+ dtemp=0
RI1_1_0_R0 I1_1_0_R0_PLUS I1_1_0_R0_MINUS rm1 W=13.5u L=230n m=1 
+ r=1.53333m dtemp=0
RI1_0_2_R0 I1_0_2_R0_PLUS I1_0_2_R0_MINUS rm1 W=230n L=50u m=1 r=19.5652 
+ dtemp=0
RI1_0_1_R0 I1_0_1_R0_PLUS I1_0_1_R0_MINUS rm1 W=230n L=13.5u m=1 
+ r=5.28261 dtemp=0
RI1_0_0_R0 I1_0_0_R0_PLUS I1_0_0_R0_MINUS rm1 W=230n L=230n m=1 r=90m 
+ dtemp=0
RI1_default I1_default_PLUS I1_default_MINUS rm1 W=230.00n L=230.00n m=1 
+ r=90.00m dtemp=0
.ENDS

