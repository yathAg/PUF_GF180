magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 352 1542 870
<< pwell >>
rect -86 -86 1542 352
<< metal1 >>
rect 0 724 1456 844
rect 26 130 115 654
rect 273 552 319 724
rect 1062 621 1130 724
rect 273 60 319 173
rect 466 242 542 542
rect 588 472 1218 557
rect 588 289 659 472
rect 802 354 1214 424
rect 1093 60 1139 176
rect 0 -60 1456 60
<< obsm1 >>
rect 365 622 778 668
rect 365 325 411 622
rect 168 278 411 325
rect 365 163 411 278
rect 1270 275 1363 676
rect 825 229 1363 275
rect 365 115 776 163
rect 1270 106 1363 229
<< labels >>
rlabel metal1 s 802 354 1214 424 6 I0
port 1 nsew default input
rlabel metal1 s 466 242 542 542 6 I1
port 2 nsew default input
rlabel metal1 s 588 289 659 472 6 S
port 3 nsew default input
rlabel metal1 s 588 472 1218 557 6 S
port 3 nsew default input
rlabel metal1 s 26 130 115 654 6 Z
port 4 nsew default output
rlabel metal1 s 1062 621 1130 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 552 319 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 724 1456 844 6 VDD
port 5 nsew power bidirectional abutment
rlabel nwell s -86 352 1542 870 6 VNW
port 6 nsew power bidirectional
rlabel pwell s -86 -86 1542 352 6 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 0 -60 1456 60 8 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1093 60 1139 176 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 60 319 173 6 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1456 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 664396
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 660396
<< end >>
