magic
tech gf180mcuB
magscale 1 10
timestamp 1698431365
<< psubdiff >>
rect 13097 70975 69968 71000
rect 13097 70929 13119 70975
rect 13165 70929 13223 70975
rect 13269 70929 13377 70975
rect 13423 70929 13481 70975
rect 13527 70929 13585 70975
rect 13631 70929 13689 70975
rect 13735 70929 13793 70975
rect 13839 70929 13897 70975
rect 13943 70929 14001 70975
rect 14047 70929 14105 70975
rect 14151 70929 14209 70975
rect 14255 70929 14313 70975
rect 14359 70929 14417 70975
rect 14463 70929 14521 70975
rect 14567 70929 14625 70975
rect 14671 70929 14729 70975
rect 14775 70929 14833 70975
rect 14879 70929 14937 70975
rect 14983 70929 15041 70975
rect 15087 70929 15145 70975
rect 15191 70929 15249 70975
rect 15295 70929 15353 70975
rect 15399 70929 15457 70975
rect 15503 70929 15561 70975
rect 15607 70929 15665 70975
rect 15711 70929 15769 70975
rect 15815 70929 15873 70975
rect 15919 70929 15977 70975
rect 16023 70929 16081 70975
rect 16127 70929 16185 70975
rect 16231 70929 16289 70975
rect 16335 70929 16393 70975
rect 16439 70929 16497 70975
rect 16543 70929 16601 70975
rect 16647 70929 16705 70975
rect 16751 70929 16809 70975
rect 16855 70929 16913 70975
rect 16959 70929 17017 70975
rect 17063 70929 17121 70975
rect 17167 70929 17225 70975
rect 17271 70929 17329 70975
rect 17375 70929 17433 70975
rect 17479 70929 17537 70975
rect 17583 70929 17641 70975
rect 17687 70929 17745 70975
rect 17791 70929 17849 70975
rect 17895 70929 17953 70975
rect 17999 70929 18057 70975
rect 18103 70929 18161 70975
rect 18207 70929 18265 70975
rect 18311 70929 18369 70975
rect 18415 70929 18473 70975
rect 18519 70929 18577 70975
rect 18623 70929 18681 70975
rect 18727 70929 18785 70975
rect 18831 70929 18889 70975
rect 18935 70929 18993 70975
rect 19039 70929 19097 70975
rect 19143 70929 19201 70975
rect 19247 70929 19305 70975
rect 19351 70929 19409 70975
rect 19455 70929 19513 70975
rect 19559 70929 19617 70975
rect 19663 70929 19721 70975
rect 19767 70929 19825 70975
rect 19871 70929 19929 70975
rect 19975 70929 20033 70975
rect 20079 70929 20137 70975
rect 20183 70929 20241 70975
rect 20287 70929 20345 70975
rect 20391 70929 20449 70975
rect 20495 70929 20553 70975
rect 20599 70929 20657 70975
rect 20703 70929 20761 70975
rect 20807 70929 20865 70975
rect 20911 70929 20969 70975
rect 21015 70929 21073 70975
rect 21119 70929 21177 70975
rect 21223 70929 21281 70975
rect 21327 70929 21385 70975
rect 21431 70929 21489 70975
rect 21535 70929 21593 70975
rect 21639 70929 21697 70975
rect 21743 70929 21801 70975
rect 21847 70929 21905 70975
rect 21951 70929 22009 70975
rect 22055 70929 22113 70975
rect 22159 70929 22217 70975
rect 22263 70929 22321 70975
rect 22367 70929 22425 70975
rect 22471 70929 22529 70975
rect 22575 70929 22633 70975
rect 22679 70929 22737 70975
rect 22783 70929 22841 70975
rect 22887 70929 22945 70975
rect 22991 70929 23049 70975
rect 23095 70929 23153 70975
rect 23199 70929 23257 70975
rect 23303 70929 23361 70975
rect 23407 70929 23465 70975
rect 23511 70929 23569 70975
rect 23615 70929 23673 70975
rect 23719 70929 23777 70975
rect 23823 70929 23881 70975
rect 23927 70929 23985 70975
rect 24031 70929 24089 70975
rect 24135 70929 24193 70975
rect 24239 70929 24297 70975
rect 24343 70929 24401 70975
rect 24447 70929 24505 70975
rect 24551 70929 24609 70975
rect 24655 70929 24713 70975
rect 24759 70929 24817 70975
rect 24863 70929 24921 70975
rect 24967 70929 25025 70975
rect 25071 70929 25129 70975
rect 25175 70929 25233 70975
rect 25279 70929 25337 70975
rect 25383 70929 25441 70975
rect 25487 70929 25545 70975
rect 25591 70929 25649 70975
rect 25695 70929 25753 70975
rect 25799 70929 25857 70975
rect 25903 70929 25961 70975
rect 26007 70929 26065 70975
rect 26111 70929 26169 70975
rect 26215 70929 26273 70975
rect 26319 70929 26377 70975
rect 26423 70929 26481 70975
rect 26527 70929 26585 70975
rect 26631 70929 26689 70975
rect 26735 70929 26793 70975
rect 26839 70929 26897 70975
rect 26943 70929 27001 70975
rect 27047 70929 27105 70975
rect 27151 70929 27209 70975
rect 27255 70929 27313 70975
rect 27359 70929 27417 70975
rect 27463 70929 27521 70975
rect 27567 70929 27625 70975
rect 27671 70929 27729 70975
rect 27775 70929 27833 70975
rect 27879 70929 27937 70975
rect 27983 70929 28041 70975
rect 28087 70929 28145 70975
rect 28191 70929 28249 70975
rect 28295 70929 28353 70975
rect 28399 70929 28457 70975
rect 28503 70929 28561 70975
rect 28607 70929 28665 70975
rect 28711 70929 28769 70975
rect 28815 70929 28873 70975
rect 28919 70929 28977 70975
rect 29023 70929 29081 70975
rect 29127 70929 29185 70975
rect 29231 70929 29289 70975
rect 29335 70929 29393 70975
rect 29439 70929 29497 70975
rect 29543 70929 29601 70975
rect 29647 70929 29705 70975
rect 29751 70929 29809 70975
rect 29855 70929 29913 70975
rect 29959 70929 30017 70975
rect 30063 70929 30121 70975
rect 30167 70929 30225 70975
rect 30271 70929 30329 70975
rect 30375 70929 30433 70975
rect 30479 70929 30537 70975
rect 30583 70929 30641 70975
rect 30687 70929 30745 70975
rect 30791 70929 30849 70975
rect 30895 70929 30953 70975
rect 30999 70929 31057 70975
rect 31103 70929 31161 70975
rect 31207 70929 31265 70975
rect 31311 70929 31369 70975
rect 31415 70929 31473 70975
rect 31519 70929 31577 70975
rect 31623 70929 31681 70975
rect 31727 70929 31785 70975
rect 31831 70929 31889 70975
rect 31935 70929 31993 70975
rect 32039 70929 32097 70975
rect 32143 70929 32201 70975
rect 32247 70929 32305 70975
rect 32351 70929 32409 70975
rect 32455 70929 32513 70975
rect 32559 70929 32617 70975
rect 32663 70929 32721 70975
rect 32767 70929 32825 70975
rect 32871 70929 32929 70975
rect 32975 70929 33033 70975
rect 33079 70929 33137 70975
rect 33183 70929 33241 70975
rect 33287 70929 33345 70975
rect 33391 70929 33449 70975
rect 33495 70929 33553 70975
rect 33599 70929 33657 70975
rect 33703 70929 33761 70975
rect 33807 70929 33865 70975
rect 33911 70929 33969 70975
rect 34015 70929 34073 70975
rect 34119 70929 34177 70975
rect 34223 70929 34281 70975
rect 34327 70929 34385 70975
rect 34431 70929 34489 70975
rect 34535 70929 34593 70975
rect 34639 70929 34697 70975
rect 34743 70929 34801 70975
rect 34847 70929 34905 70975
rect 34951 70929 35009 70975
rect 35055 70929 35113 70975
rect 35159 70929 35217 70975
rect 35263 70929 35321 70975
rect 35367 70929 35425 70975
rect 35471 70929 35529 70975
rect 35575 70929 35633 70975
rect 35679 70929 35737 70975
rect 35783 70929 35841 70975
rect 35887 70929 35945 70975
rect 35991 70929 36049 70975
rect 36095 70929 36153 70975
rect 36199 70929 36257 70975
rect 36303 70929 36361 70975
rect 36407 70929 36465 70975
rect 36511 70929 36569 70975
rect 36615 70929 36673 70975
rect 36719 70929 36777 70975
rect 36823 70929 36881 70975
rect 36927 70929 36985 70975
rect 37031 70929 37089 70975
rect 37135 70929 37193 70975
rect 37239 70929 37297 70975
rect 37343 70929 37401 70975
rect 37447 70929 37505 70975
rect 37551 70929 37609 70975
rect 37655 70929 37713 70975
rect 37759 70929 37817 70975
rect 37863 70929 37921 70975
rect 37967 70929 38025 70975
rect 38071 70929 38129 70975
rect 38175 70929 38233 70975
rect 38279 70929 38337 70975
rect 38383 70929 38441 70975
rect 38487 70929 38545 70975
rect 38591 70929 38649 70975
rect 38695 70929 38753 70975
rect 38799 70929 38857 70975
rect 38903 70929 38961 70975
rect 39007 70929 39065 70975
rect 39111 70929 39169 70975
rect 39215 70929 39273 70975
rect 39319 70929 39377 70975
rect 39423 70929 39481 70975
rect 39527 70929 39585 70975
rect 39631 70929 39689 70975
rect 39735 70929 39793 70975
rect 39839 70929 39897 70975
rect 39943 70929 40001 70975
rect 40047 70929 40105 70975
rect 40151 70929 40209 70975
rect 40255 70929 40313 70975
rect 40359 70929 40417 70975
rect 40463 70929 40521 70975
rect 40567 70929 40625 70975
rect 40671 70929 40729 70975
rect 40775 70929 40833 70975
rect 40879 70929 40937 70975
rect 40983 70929 41041 70975
rect 41087 70929 41145 70975
rect 41191 70929 41249 70975
rect 41295 70929 41353 70975
rect 41399 70929 41457 70975
rect 41503 70929 41561 70975
rect 41607 70929 41665 70975
rect 41711 70929 41769 70975
rect 41815 70929 41873 70975
rect 41919 70929 41977 70975
rect 42023 70929 42081 70975
rect 42127 70929 42185 70975
rect 42231 70929 42289 70975
rect 42335 70929 42393 70975
rect 42439 70929 42497 70975
rect 42543 70929 42601 70975
rect 42647 70929 42705 70975
rect 42751 70929 42809 70975
rect 42855 70929 42913 70975
rect 42959 70929 43017 70975
rect 43063 70929 43121 70975
rect 43167 70929 43225 70975
rect 43271 70929 43329 70975
rect 43375 70929 43433 70975
rect 43479 70929 43537 70975
rect 43583 70929 43641 70975
rect 43687 70929 43745 70975
rect 43791 70929 43849 70975
rect 43895 70929 43953 70975
rect 43999 70929 44057 70975
rect 44103 70929 44161 70975
rect 44207 70929 44265 70975
rect 44311 70929 44369 70975
rect 44415 70929 44473 70975
rect 44519 70929 44577 70975
rect 44623 70929 44681 70975
rect 44727 70929 44785 70975
rect 44831 70929 44889 70975
rect 44935 70929 44993 70975
rect 45039 70929 45097 70975
rect 45143 70929 45201 70975
rect 45247 70929 45305 70975
rect 45351 70929 45409 70975
rect 45455 70929 45513 70975
rect 45559 70929 45617 70975
rect 45663 70929 45721 70975
rect 45767 70929 45825 70975
rect 45871 70929 45929 70975
rect 45975 70929 46033 70975
rect 46079 70929 46137 70975
rect 46183 70929 46241 70975
rect 46287 70929 46345 70975
rect 46391 70929 46449 70975
rect 46495 70929 46553 70975
rect 46599 70929 46657 70975
rect 46703 70929 46761 70975
rect 46807 70929 46865 70975
rect 46911 70929 46969 70975
rect 47015 70929 47073 70975
rect 47119 70929 47177 70975
rect 47223 70929 47281 70975
rect 47327 70929 47385 70975
rect 47431 70929 47489 70975
rect 47535 70929 47593 70975
rect 47639 70929 47697 70975
rect 47743 70929 47801 70975
rect 47847 70929 47905 70975
rect 47951 70929 48009 70975
rect 48055 70929 48113 70975
rect 48159 70929 48217 70975
rect 48263 70929 48321 70975
rect 48367 70929 48425 70975
rect 48471 70929 48529 70975
rect 48575 70929 48633 70975
rect 48679 70929 48737 70975
rect 48783 70929 48841 70975
rect 48887 70929 48945 70975
rect 48991 70929 49049 70975
rect 49095 70929 49153 70975
rect 49199 70929 49257 70975
rect 49303 70929 49361 70975
rect 49407 70929 49465 70975
rect 49511 70929 49569 70975
rect 49615 70929 49673 70975
rect 49719 70929 49777 70975
rect 49823 70929 49881 70975
rect 49927 70929 49985 70975
rect 50031 70929 50089 70975
rect 50135 70929 50193 70975
rect 50239 70929 50297 70975
rect 50343 70929 50401 70975
rect 50447 70929 50505 70975
rect 50551 70929 50609 70975
rect 50655 70929 50713 70975
rect 50759 70929 50817 70975
rect 50863 70929 50921 70975
rect 50967 70929 51025 70975
rect 51071 70929 51129 70975
rect 51175 70929 51233 70975
rect 51279 70929 51337 70975
rect 51383 70929 51441 70975
rect 51487 70929 51545 70975
rect 51591 70929 51649 70975
rect 51695 70929 51753 70975
rect 51799 70929 51857 70975
rect 51903 70929 51961 70975
rect 52007 70929 52065 70975
rect 52111 70929 52169 70975
rect 52215 70929 52273 70975
rect 52319 70929 52377 70975
rect 52423 70929 52481 70975
rect 52527 70929 52585 70975
rect 52631 70929 52689 70975
rect 52735 70929 52793 70975
rect 52839 70929 52897 70975
rect 52943 70929 53001 70975
rect 53047 70929 53105 70975
rect 53151 70929 53209 70975
rect 53255 70929 53313 70975
rect 53359 70929 53417 70975
rect 53463 70929 53521 70975
rect 53567 70929 53625 70975
rect 53671 70929 53729 70975
rect 53775 70929 53833 70975
rect 53879 70929 53937 70975
rect 53983 70929 54041 70975
rect 54087 70929 54145 70975
rect 54191 70929 54249 70975
rect 54295 70929 54353 70975
rect 54399 70929 54457 70975
rect 54503 70929 54561 70975
rect 54607 70929 54665 70975
rect 54711 70929 54769 70975
rect 54815 70929 54873 70975
rect 54919 70929 54977 70975
rect 55023 70929 55081 70975
rect 55127 70929 55185 70975
rect 55231 70929 55289 70975
rect 55335 70929 55393 70975
rect 55439 70929 55497 70975
rect 55543 70929 55601 70975
rect 55647 70929 55705 70975
rect 55751 70929 55809 70975
rect 55855 70929 55913 70975
rect 55959 70929 56017 70975
rect 56063 70929 56121 70975
rect 56167 70929 56225 70975
rect 56271 70929 56329 70975
rect 56375 70929 56433 70975
rect 56479 70929 56537 70975
rect 56583 70929 56641 70975
rect 56687 70929 56745 70975
rect 56791 70929 56849 70975
rect 56895 70929 56953 70975
rect 56999 70929 57057 70975
rect 57103 70929 57161 70975
rect 57207 70929 57265 70975
rect 57311 70929 57369 70975
rect 57415 70929 57473 70975
rect 57519 70929 57577 70975
rect 57623 70929 57681 70975
rect 57727 70929 57785 70975
rect 57831 70929 57889 70975
rect 57935 70929 57993 70975
rect 58039 70929 58097 70975
rect 58143 70929 58201 70975
rect 58247 70929 58305 70975
rect 58351 70929 58409 70975
rect 58455 70929 58513 70975
rect 58559 70929 58617 70975
rect 58663 70929 58721 70975
rect 58767 70929 58825 70975
rect 58871 70929 58929 70975
rect 58975 70929 59033 70975
rect 59079 70929 59137 70975
rect 59183 70929 59241 70975
rect 59287 70929 59345 70975
rect 59391 70929 59449 70975
rect 59495 70929 59553 70975
rect 59599 70929 59657 70975
rect 59703 70929 59761 70975
rect 59807 70929 59865 70975
rect 59911 70929 59969 70975
rect 60015 70929 60073 70975
rect 60119 70929 60177 70975
rect 60223 70929 60281 70975
rect 60327 70929 60385 70975
rect 60431 70929 60489 70975
rect 60535 70929 60593 70975
rect 60639 70929 60697 70975
rect 60743 70929 60801 70975
rect 60847 70929 60905 70975
rect 60951 70929 61009 70975
rect 61055 70929 61113 70975
rect 61159 70929 61217 70975
rect 61263 70929 61321 70975
rect 61367 70929 61425 70975
rect 61471 70929 61529 70975
rect 61575 70929 61633 70975
rect 61679 70929 61737 70975
rect 61783 70929 61841 70975
rect 61887 70929 61945 70975
rect 61991 70929 62049 70975
rect 62095 70929 62153 70975
rect 62199 70929 62257 70975
rect 62303 70929 62361 70975
rect 62407 70929 62465 70975
rect 62511 70929 62569 70975
rect 62615 70929 62673 70975
rect 62719 70929 62777 70975
rect 62823 70929 62881 70975
rect 62927 70929 62985 70975
rect 63031 70929 63089 70975
rect 63135 70929 63193 70975
rect 63239 70929 63297 70975
rect 63343 70929 63401 70975
rect 63447 70929 63505 70975
rect 63551 70929 63609 70975
rect 63655 70929 63713 70975
rect 63759 70929 63817 70975
rect 63863 70929 63921 70975
rect 63967 70929 64025 70975
rect 64071 70929 64129 70975
rect 64175 70929 64233 70975
rect 64279 70929 64337 70975
rect 64383 70929 64441 70975
rect 64487 70929 64545 70975
rect 64591 70929 64649 70975
rect 64695 70929 64753 70975
rect 64799 70929 64857 70975
rect 64903 70929 64961 70975
rect 65007 70929 65065 70975
rect 65111 70929 65169 70975
rect 65215 70929 65273 70975
rect 65319 70929 65377 70975
rect 65423 70929 65481 70975
rect 65527 70929 65585 70975
rect 65631 70929 65689 70975
rect 65735 70929 65793 70975
rect 65839 70929 65897 70975
rect 65943 70929 66001 70975
rect 66047 70929 66105 70975
rect 66151 70929 66209 70975
rect 66255 70929 66313 70975
rect 66359 70929 66417 70975
rect 66463 70929 66521 70975
rect 66567 70929 66625 70975
rect 66671 70929 66729 70975
rect 66775 70929 66833 70975
rect 66879 70929 66937 70975
rect 66983 70929 67041 70975
rect 67087 70929 67145 70975
rect 67191 70929 67249 70975
rect 67295 70929 67353 70975
rect 67399 70929 67457 70975
rect 67503 70929 67561 70975
rect 67607 70929 67665 70975
rect 67711 70929 67769 70975
rect 67815 70929 67873 70975
rect 67919 70929 67977 70975
rect 68023 70929 68081 70975
rect 68127 70929 68185 70975
rect 68231 70929 68289 70975
rect 68335 70929 68393 70975
rect 68439 70929 68497 70975
rect 68543 70929 68601 70975
rect 68647 70929 68705 70975
rect 68751 70929 68809 70975
rect 68855 70929 68913 70975
rect 68959 70929 69017 70975
rect 69063 70929 69121 70975
rect 69167 70929 69225 70975
rect 69271 70929 69329 70975
rect 69375 70929 69433 70975
rect 69479 70929 69537 70975
rect 69583 70929 69641 70975
rect 69687 70929 69745 70975
rect 69791 70929 69849 70975
rect 69895 70929 69968 70975
rect 13097 70871 69968 70929
rect 13097 70825 13119 70871
rect 13165 70825 13223 70871
rect 13269 70825 13377 70871
rect 13423 70825 13481 70871
rect 13527 70825 13585 70871
rect 13631 70825 13689 70871
rect 13735 70825 13793 70871
rect 13839 70825 13897 70871
rect 13943 70825 14001 70871
rect 14047 70825 14105 70871
rect 14151 70825 14209 70871
rect 14255 70825 14313 70871
rect 14359 70825 14417 70871
rect 14463 70825 14521 70871
rect 14567 70825 14625 70871
rect 14671 70825 14729 70871
rect 14775 70825 14833 70871
rect 14879 70825 14937 70871
rect 14983 70825 15041 70871
rect 15087 70825 15145 70871
rect 15191 70825 15249 70871
rect 15295 70825 15353 70871
rect 15399 70825 15457 70871
rect 15503 70825 15561 70871
rect 15607 70825 15665 70871
rect 15711 70825 15769 70871
rect 15815 70825 15873 70871
rect 15919 70825 15977 70871
rect 16023 70825 16081 70871
rect 16127 70825 16185 70871
rect 16231 70825 16289 70871
rect 16335 70825 16393 70871
rect 16439 70825 16497 70871
rect 16543 70825 16601 70871
rect 16647 70825 16705 70871
rect 16751 70825 16809 70871
rect 16855 70825 16913 70871
rect 16959 70825 17017 70871
rect 17063 70825 17121 70871
rect 17167 70825 17225 70871
rect 17271 70825 17329 70871
rect 17375 70825 17433 70871
rect 17479 70825 17537 70871
rect 17583 70825 17641 70871
rect 17687 70825 17745 70871
rect 17791 70825 17849 70871
rect 17895 70825 17953 70871
rect 17999 70825 18057 70871
rect 18103 70825 18161 70871
rect 18207 70825 18265 70871
rect 18311 70825 18369 70871
rect 18415 70825 18473 70871
rect 18519 70825 18577 70871
rect 18623 70825 18681 70871
rect 18727 70825 18785 70871
rect 18831 70825 18889 70871
rect 18935 70825 18993 70871
rect 19039 70825 19097 70871
rect 19143 70825 19201 70871
rect 19247 70825 19305 70871
rect 19351 70825 19409 70871
rect 19455 70825 19513 70871
rect 19559 70825 19617 70871
rect 19663 70825 19721 70871
rect 19767 70825 19825 70871
rect 19871 70825 19929 70871
rect 19975 70825 20033 70871
rect 20079 70825 20137 70871
rect 20183 70825 20241 70871
rect 20287 70825 20345 70871
rect 20391 70825 20449 70871
rect 20495 70825 20553 70871
rect 20599 70825 20657 70871
rect 20703 70825 20761 70871
rect 20807 70825 20865 70871
rect 20911 70825 20969 70871
rect 21015 70825 21073 70871
rect 21119 70825 21177 70871
rect 21223 70825 21281 70871
rect 21327 70825 21385 70871
rect 21431 70825 21489 70871
rect 21535 70825 21593 70871
rect 21639 70825 21697 70871
rect 21743 70825 21801 70871
rect 21847 70825 21905 70871
rect 21951 70825 22009 70871
rect 22055 70825 22113 70871
rect 22159 70825 22217 70871
rect 22263 70825 22321 70871
rect 22367 70825 22425 70871
rect 22471 70825 22529 70871
rect 22575 70825 22633 70871
rect 22679 70825 22737 70871
rect 22783 70825 22841 70871
rect 22887 70825 22945 70871
rect 22991 70825 23049 70871
rect 23095 70825 23153 70871
rect 23199 70825 23257 70871
rect 23303 70825 23361 70871
rect 23407 70825 23465 70871
rect 23511 70825 23569 70871
rect 23615 70825 23673 70871
rect 23719 70825 23777 70871
rect 23823 70825 23881 70871
rect 23927 70825 23985 70871
rect 24031 70825 24089 70871
rect 24135 70825 24193 70871
rect 24239 70825 24297 70871
rect 24343 70825 24401 70871
rect 24447 70825 24505 70871
rect 24551 70825 24609 70871
rect 24655 70825 24713 70871
rect 24759 70825 24817 70871
rect 24863 70825 24921 70871
rect 24967 70825 25025 70871
rect 25071 70825 25129 70871
rect 25175 70825 25233 70871
rect 25279 70825 25337 70871
rect 25383 70825 25441 70871
rect 25487 70825 25545 70871
rect 25591 70825 25649 70871
rect 25695 70825 25753 70871
rect 25799 70825 25857 70871
rect 25903 70825 25961 70871
rect 26007 70825 26065 70871
rect 26111 70825 26169 70871
rect 26215 70825 26273 70871
rect 26319 70825 26377 70871
rect 26423 70825 26481 70871
rect 26527 70825 26585 70871
rect 26631 70825 26689 70871
rect 26735 70825 26793 70871
rect 26839 70825 26897 70871
rect 26943 70825 27001 70871
rect 27047 70825 27105 70871
rect 27151 70825 27209 70871
rect 27255 70825 27313 70871
rect 27359 70825 27417 70871
rect 27463 70825 27521 70871
rect 27567 70825 27625 70871
rect 27671 70825 27729 70871
rect 27775 70825 27833 70871
rect 27879 70825 27937 70871
rect 27983 70825 28041 70871
rect 28087 70825 28145 70871
rect 28191 70825 28249 70871
rect 28295 70825 28353 70871
rect 28399 70825 28457 70871
rect 28503 70825 28561 70871
rect 28607 70825 28665 70871
rect 28711 70825 28769 70871
rect 28815 70825 28873 70871
rect 28919 70825 28977 70871
rect 29023 70825 29081 70871
rect 29127 70825 29185 70871
rect 29231 70825 29289 70871
rect 29335 70825 29393 70871
rect 29439 70825 29497 70871
rect 29543 70825 29601 70871
rect 29647 70825 29705 70871
rect 29751 70825 29809 70871
rect 29855 70825 29913 70871
rect 29959 70825 30017 70871
rect 30063 70825 30121 70871
rect 30167 70825 30225 70871
rect 30271 70825 30329 70871
rect 30375 70825 30433 70871
rect 30479 70825 30537 70871
rect 30583 70825 30641 70871
rect 30687 70825 30745 70871
rect 30791 70825 30849 70871
rect 30895 70825 30953 70871
rect 30999 70825 31057 70871
rect 31103 70825 31161 70871
rect 31207 70825 31265 70871
rect 31311 70825 31369 70871
rect 31415 70825 31473 70871
rect 31519 70825 31577 70871
rect 31623 70825 31681 70871
rect 31727 70825 31785 70871
rect 31831 70825 31889 70871
rect 31935 70825 31993 70871
rect 32039 70825 32097 70871
rect 32143 70825 32201 70871
rect 32247 70825 32305 70871
rect 32351 70825 32409 70871
rect 32455 70825 32513 70871
rect 32559 70825 32617 70871
rect 32663 70825 32721 70871
rect 32767 70825 32825 70871
rect 32871 70825 32929 70871
rect 32975 70825 33033 70871
rect 33079 70825 33137 70871
rect 33183 70825 33241 70871
rect 33287 70825 33345 70871
rect 33391 70825 33449 70871
rect 33495 70825 33553 70871
rect 33599 70825 33657 70871
rect 33703 70825 33761 70871
rect 33807 70825 33865 70871
rect 33911 70825 33969 70871
rect 34015 70825 34073 70871
rect 34119 70825 34177 70871
rect 34223 70825 34281 70871
rect 34327 70825 34385 70871
rect 34431 70825 34489 70871
rect 34535 70825 34593 70871
rect 34639 70825 34697 70871
rect 34743 70825 34801 70871
rect 34847 70825 34905 70871
rect 34951 70825 35009 70871
rect 35055 70825 35113 70871
rect 35159 70825 35217 70871
rect 35263 70825 35321 70871
rect 35367 70825 35425 70871
rect 35471 70825 35529 70871
rect 35575 70825 35633 70871
rect 35679 70825 35737 70871
rect 35783 70825 35841 70871
rect 35887 70825 35945 70871
rect 35991 70825 36049 70871
rect 36095 70825 36153 70871
rect 36199 70825 36257 70871
rect 36303 70825 36361 70871
rect 36407 70825 36465 70871
rect 36511 70825 36569 70871
rect 36615 70825 36673 70871
rect 36719 70825 36777 70871
rect 36823 70825 36881 70871
rect 36927 70825 36985 70871
rect 37031 70825 37089 70871
rect 37135 70825 37193 70871
rect 37239 70825 37297 70871
rect 37343 70825 37401 70871
rect 37447 70825 37505 70871
rect 37551 70825 37609 70871
rect 37655 70825 37713 70871
rect 37759 70825 37817 70871
rect 37863 70825 37921 70871
rect 37967 70825 38025 70871
rect 38071 70825 38129 70871
rect 38175 70825 38233 70871
rect 38279 70825 38337 70871
rect 38383 70825 38441 70871
rect 38487 70825 38545 70871
rect 38591 70825 38649 70871
rect 38695 70825 38753 70871
rect 38799 70825 38857 70871
rect 38903 70825 38961 70871
rect 39007 70825 39065 70871
rect 39111 70825 39169 70871
rect 39215 70825 39273 70871
rect 39319 70825 39377 70871
rect 39423 70825 39481 70871
rect 39527 70825 39585 70871
rect 39631 70825 39689 70871
rect 39735 70825 39793 70871
rect 39839 70825 39897 70871
rect 39943 70825 40001 70871
rect 40047 70825 40105 70871
rect 40151 70825 40209 70871
rect 40255 70825 40313 70871
rect 40359 70825 40417 70871
rect 40463 70825 40521 70871
rect 40567 70825 40625 70871
rect 40671 70825 40729 70871
rect 40775 70825 40833 70871
rect 40879 70825 40937 70871
rect 40983 70825 41041 70871
rect 41087 70825 41145 70871
rect 41191 70825 41249 70871
rect 41295 70825 41353 70871
rect 41399 70825 41457 70871
rect 41503 70825 41561 70871
rect 41607 70825 41665 70871
rect 41711 70825 41769 70871
rect 41815 70825 41873 70871
rect 41919 70825 41977 70871
rect 42023 70825 42081 70871
rect 42127 70825 42185 70871
rect 42231 70825 42289 70871
rect 42335 70825 42393 70871
rect 42439 70825 42497 70871
rect 42543 70825 42601 70871
rect 42647 70825 42705 70871
rect 42751 70825 42809 70871
rect 42855 70825 42913 70871
rect 42959 70825 43017 70871
rect 43063 70825 43121 70871
rect 43167 70825 43225 70871
rect 43271 70825 43329 70871
rect 43375 70825 43433 70871
rect 43479 70825 43537 70871
rect 43583 70825 43641 70871
rect 43687 70825 43745 70871
rect 43791 70825 43849 70871
rect 43895 70825 43953 70871
rect 43999 70825 44057 70871
rect 44103 70825 44161 70871
rect 44207 70825 44265 70871
rect 44311 70825 44369 70871
rect 44415 70825 44473 70871
rect 44519 70825 44577 70871
rect 44623 70825 44681 70871
rect 44727 70825 44785 70871
rect 44831 70825 44889 70871
rect 44935 70825 44993 70871
rect 45039 70825 45097 70871
rect 45143 70825 45201 70871
rect 45247 70825 45305 70871
rect 45351 70825 45409 70871
rect 45455 70825 45513 70871
rect 45559 70825 45617 70871
rect 45663 70825 45721 70871
rect 45767 70825 45825 70871
rect 45871 70825 45929 70871
rect 45975 70825 46033 70871
rect 46079 70825 46137 70871
rect 46183 70825 46241 70871
rect 46287 70825 46345 70871
rect 46391 70825 46449 70871
rect 46495 70825 46553 70871
rect 46599 70825 46657 70871
rect 46703 70825 46761 70871
rect 46807 70825 46865 70871
rect 46911 70825 46969 70871
rect 47015 70825 47073 70871
rect 47119 70825 47177 70871
rect 47223 70825 47281 70871
rect 47327 70825 47385 70871
rect 47431 70825 47489 70871
rect 47535 70825 47593 70871
rect 47639 70825 47697 70871
rect 47743 70825 47801 70871
rect 47847 70825 47905 70871
rect 47951 70825 48009 70871
rect 48055 70825 48113 70871
rect 48159 70825 48217 70871
rect 48263 70825 48321 70871
rect 48367 70825 48425 70871
rect 48471 70825 48529 70871
rect 48575 70825 48633 70871
rect 48679 70825 48737 70871
rect 48783 70825 48841 70871
rect 48887 70825 48945 70871
rect 48991 70825 49049 70871
rect 49095 70825 49153 70871
rect 49199 70825 49257 70871
rect 49303 70825 49361 70871
rect 49407 70825 49465 70871
rect 49511 70825 49569 70871
rect 49615 70825 49673 70871
rect 49719 70825 49777 70871
rect 49823 70825 49881 70871
rect 49927 70825 49985 70871
rect 50031 70825 50089 70871
rect 50135 70825 50193 70871
rect 50239 70825 50297 70871
rect 50343 70825 50401 70871
rect 50447 70825 50505 70871
rect 50551 70825 50609 70871
rect 50655 70825 50713 70871
rect 50759 70825 50817 70871
rect 50863 70825 50921 70871
rect 50967 70825 51025 70871
rect 51071 70825 51129 70871
rect 51175 70825 51233 70871
rect 51279 70825 51337 70871
rect 51383 70825 51441 70871
rect 51487 70825 51545 70871
rect 51591 70825 51649 70871
rect 51695 70825 51753 70871
rect 51799 70825 51857 70871
rect 51903 70825 51961 70871
rect 52007 70825 52065 70871
rect 52111 70825 52169 70871
rect 52215 70825 52273 70871
rect 52319 70825 52377 70871
rect 52423 70825 52481 70871
rect 52527 70825 52585 70871
rect 52631 70825 52689 70871
rect 52735 70825 52793 70871
rect 52839 70825 52897 70871
rect 52943 70825 53001 70871
rect 53047 70825 53105 70871
rect 53151 70825 53209 70871
rect 53255 70825 53313 70871
rect 53359 70825 53417 70871
rect 53463 70825 53521 70871
rect 53567 70825 53625 70871
rect 53671 70825 53729 70871
rect 53775 70825 53833 70871
rect 53879 70825 53937 70871
rect 53983 70825 54041 70871
rect 54087 70825 54145 70871
rect 54191 70825 54249 70871
rect 54295 70825 54353 70871
rect 54399 70825 54457 70871
rect 54503 70825 54561 70871
rect 54607 70825 54665 70871
rect 54711 70825 54769 70871
rect 54815 70825 54873 70871
rect 54919 70825 54977 70871
rect 55023 70825 55081 70871
rect 55127 70825 55185 70871
rect 55231 70825 55289 70871
rect 55335 70825 55393 70871
rect 55439 70825 55497 70871
rect 55543 70825 55601 70871
rect 55647 70825 55705 70871
rect 55751 70825 55809 70871
rect 55855 70825 55913 70871
rect 55959 70825 56017 70871
rect 56063 70825 56121 70871
rect 56167 70825 56225 70871
rect 56271 70825 56329 70871
rect 56375 70825 56433 70871
rect 56479 70825 56537 70871
rect 56583 70825 56641 70871
rect 56687 70825 56745 70871
rect 56791 70825 56849 70871
rect 56895 70825 56953 70871
rect 56999 70825 57057 70871
rect 57103 70825 57161 70871
rect 57207 70825 57265 70871
rect 57311 70825 57369 70871
rect 57415 70825 57473 70871
rect 57519 70825 57577 70871
rect 57623 70825 57681 70871
rect 57727 70825 57785 70871
rect 57831 70825 57889 70871
rect 57935 70825 57993 70871
rect 58039 70825 58097 70871
rect 58143 70825 58201 70871
rect 58247 70825 58305 70871
rect 58351 70825 58409 70871
rect 58455 70825 58513 70871
rect 58559 70825 58617 70871
rect 58663 70825 58721 70871
rect 58767 70825 58825 70871
rect 58871 70825 58929 70871
rect 58975 70825 59033 70871
rect 59079 70825 59137 70871
rect 59183 70825 59241 70871
rect 59287 70825 59345 70871
rect 59391 70825 59449 70871
rect 59495 70825 59553 70871
rect 59599 70825 59657 70871
rect 59703 70825 59761 70871
rect 59807 70825 59865 70871
rect 59911 70825 59969 70871
rect 60015 70825 60073 70871
rect 60119 70825 60177 70871
rect 60223 70825 60281 70871
rect 60327 70825 60385 70871
rect 60431 70825 60489 70871
rect 60535 70825 60593 70871
rect 60639 70825 60697 70871
rect 60743 70825 60801 70871
rect 60847 70825 60905 70871
rect 60951 70825 61009 70871
rect 61055 70825 61113 70871
rect 61159 70825 61217 70871
rect 61263 70825 61321 70871
rect 61367 70825 61425 70871
rect 61471 70825 61529 70871
rect 61575 70825 61633 70871
rect 61679 70825 61737 70871
rect 61783 70825 61841 70871
rect 61887 70825 61945 70871
rect 61991 70825 62049 70871
rect 62095 70825 62153 70871
rect 62199 70825 62257 70871
rect 62303 70825 62361 70871
rect 62407 70825 62465 70871
rect 62511 70825 62569 70871
rect 62615 70825 62673 70871
rect 62719 70825 62777 70871
rect 62823 70825 62881 70871
rect 62927 70825 62985 70871
rect 63031 70825 63089 70871
rect 63135 70825 63193 70871
rect 63239 70825 63297 70871
rect 63343 70825 63401 70871
rect 63447 70825 63505 70871
rect 63551 70825 63609 70871
rect 63655 70825 63713 70871
rect 63759 70825 63817 70871
rect 63863 70825 63921 70871
rect 63967 70825 64025 70871
rect 64071 70825 64129 70871
rect 64175 70825 64233 70871
rect 64279 70825 64337 70871
rect 64383 70825 64441 70871
rect 64487 70825 64545 70871
rect 64591 70825 64649 70871
rect 64695 70825 64753 70871
rect 64799 70825 64857 70871
rect 64903 70825 64961 70871
rect 65007 70825 65065 70871
rect 65111 70825 65169 70871
rect 65215 70825 65273 70871
rect 65319 70825 65377 70871
rect 65423 70825 65481 70871
rect 65527 70825 65585 70871
rect 65631 70825 65689 70871
rect 65735 70825 65793 70871
rect 65839 70825 65897 70871
rect 65943 70825 66001 70871
rect 66047 70825 66105 70871
rect 66151 70825 66209 70871
rect 66255 70825 66313 70871
rect 66359 70825 66417 70871
rect 66463 70825 66521 70871
rect 66567 70825 66625 70871
rect 66671 70825 66729 70871
rect 66775 70825 66833 70871
rect 66879 70825 66937 70871
rect 66983 70825 67041 70871
rect 67087 70825 67145 70871
rect 67191 70825 67249 70871
rect 67295 70825 67353 70871
rect 67399 70825 67457 70871
rect 67503 70825 67561 70871
rect 67607 70825 67665 70871
rect 67711 70825 67769 70871
rect 67815 70825 67873 70871
rect 67919 70825 67977 70871
rect 68023 70825 68081 70871
rect 68127 70825 68185 70871
rect 68231 70825 68289 70871
rect 68335 70825 68393 70871
rect 68439 70825 68497 70871
rect 68543 70825 68601 70871
rect 68647 70825 68705 70871
rect 68751 70825 68809 70871
rect 68855 70825 68913 70871
rect 68959 70825 69017 70871
rect 69063 70825 69121 70871
rect 69167 70825 69225 70871
rect 69271 70825 69329 70871
rect 69375 70825 69433 70871
rect 69479 70825 69537 70871
rect 69583 70825 69641 70871
rect 69687 70825 69745 70871
rect 69791 70825 69849 70871
rect 69895 70825 69968 70871
rect 13097 70803 69968 70825
rect 13097 70767 13291 70803
rect 13097 70721 13119 70767
rect 13165 70721 13223 70767
rect 13269 70721 13291 70767
rect 13097 70663 13291 70721
rect 13097 70617 13119 70663
rect 13165 70617 13223 70663
rect 13269 70617 13291 70663
rect 13097 70559 13291 70617
rect 13097 70513 13119 70559
rect 13165 70513 13223 70559
rect 13269 70513 13291 70559
rect 13097 70455 13291 70513
rect 13097 70409 13119 70455
rect 13165 70409 13223 70455
rect 13269 70409 13291 70455
rect 13097 70351 13291 70409
rect 13097 70305 13119 70351
rect 13165 70305 13223 70351
rect 13269 70305 13291 70351
rect 13097 70247 13291 70305
rect 13097 70201 13119 70247
rect 13165 70201 13223 70247
rect 13269 70201 13291 70247
rect 13097 70143 13291 70201
rect 13097 70097 13119 70143
rect 13165 70097 13223 70143
rect 13269 70097 13291 70143
rect 13097 70039 13291 70097
rect 13097 69993 13119 70039
rect 13165 69993 13223 70039
rect 13269 69993 13291 70039
rect 13097 69935 13291 69993
rect 13097 69889 13119 69935
rect 13165 69889 13223 69935
rect 13269 69889 13291 69935
rect 13097 69831 13291 69889
rect 13097 69785 13119 69831
rect 13165 69785 13223 69831
rect 13269 69785 13291 69831
rect 13097 69727 13291 69785
rect 69774 70720 69968 70803
rect 69774 70674 69796 70720
rect 69842 70674 69900 70720
rect 69946 70674 69968 70720
rect 69774 70616 69968 70674
rect 69774 70570 69796 70616
rect 69842 70570 69900 70616
rect 69946 70570 69968 70616
rect 69774 70512 69968 70570
rect 69774 70466 69796 70512
rect 69842 70466 69900 70512
rect 69946 70466 69968 70512
rect 69774 70408 69968 70466
rect 69774 70362 69796 70408
rect 69842 70362 69900 70408
rect 69946 70362 69968 70408
rect 69774 70304 69968 70362
rect 69774 70258 69796 70304
rect 69842 70258 69900 70304
rect 69946 70258 69968 70304
rect 69774 70200 69968 70258
rect 69774 70154 69796 70200
rect 69842 70154 69900 70200
rect 69946 70154 69968 70200
rect 69774 70096 69968 70154
rect 69774 70050 69796 70096
rect 69842 70050 69900 70096
rect 69946 70050 69968 70096
rect 69774 69968 69968 70050
rect 69774 69946 71000 69968
rect 69774 69900 69796 69946
rect 69842 69900 69900 69946
rect 69946 69900 70004 69946
rect 70050 69900 70108 69946
rect 70154 69900 70212 69946
rect 70258 69900 70316 69946
rect 70362 69900 70420 69946
rect 70466 69900 70524 69946
rect 70570 69900 70628 69946
rect 70674 69908 71000 69946
rect 70674 69900 70824 69908
rect 69774 69862 70824 69900
rect 70870 69862 70928 69908
rect 70974 69862 71000 69908
rect 69774 69842 71000 69862
rect 69774 69796 69796 69842
rect 69842 69796 69900 69842
rect 69946 69796 70004 69842
rect 70050 69796 70108 69842
rect 70154 69796 70212 69842
rect 70258 69796 70316 69842
rect 70362 69796 70420 69842
rect 70466 69796 70524 69842
rect 70570 69796 70628 69842
rect 70674 69804 71000 69842
rect 70674 69796 70824 69804
rect 69774 69774 70824 69796
rect 13097 69681 13119 69727
rect 13165 69681 13223 69727
rect 13269 69681 13291 69727
rect 13097 69623 13291 69681
rect 13097 69577 13119 69623
rect 13165 69577 13223 69623
rect 13269 69577 13291 69623
rect 13097 69519 13291 69577
rect 13097 69473 13119 69519
rect 13165 69473 13223 69519
rect 13269 69473 13291 69519
rect 13097 69415 13291 69473
rect 13097 69369 13119 69415
rect 13165 69369 13223 69415
rect 13269 69369 13291 69415
rect 13097 69311 13291 69369
rect 13097 69265 13119 69311
rect 13165 69265 13223 69311
rect 13269 69265 13291 69311
rect 13097 69207 13291 69265
rect 13097 69161 13119 69207
rect 13165 69161 13223 69207
rect 13269 69161 13291 69207
rect 13097 69103 13291 69161
rect 13097 69057 13119 69103
rect 13165 69057 13223 69103
rect 13269 69057 13291 69103
rect 13097 68999 13291 69057
rect 13097 68953 13119 68999
rect 13165 68953 13223 68999
rect 13269 68953 13291 68999
rect 13097 68895 13291 68953
rect 13097 68849 13119 68895
rect 13165 68849 13223 68895
rect 13269 68849 13291 68895
rect 13097 68791 13291 68849
rect 13097 68745 13119 68791
rect 13165 68745 13223 68791
rect 13269 68745 13291 68791
rect 13097 68687 13291 68745
rect 13097 68641 13119 68687
rect 13165 68641 13223 68687
rect 13269 68641 13291 68687
rect 13097 68583 13291 68641
rect 13097 68537 13119 68583
rect 13165 68537 13223 68583
rect 13269 68537 13291 68583
rect 13097 68479 13291 68537
rect 13097 68433 13119 68479
rect 13165 68433 13223 68479
rect 13269 68433 13291 68479
rect 13097 68375 13291 68433
rect 13097 68329 13119 68375
rect 13165 68329 13223 68375
rect 13269 68329 13291 68375
rect 13097 68271 13291 68329
rect 13097 68225 13119 68271
rect 13165 68225 13223 68271
rect 13269 68225 13291 68271
rect 13097 68167 13291 68225
rect 13097 68121 13119 68167
rect 13165 68121 13223 68167
rect 13269 68121 13291 68167
rect 13097 68063 13291 68121
rect 13097 68017 13119 68063
rect 13165 68017 13223 68063
rect 13269 68017 13291 68063
rect 13097 67959 13291 68017
rect 13097 67913 13119 67959
rect 13165 67913 13223 67959
rect 13269 67913 13291 67959
rect 13097 67855 13291 67913
rect 13097 67809 13119 67855
rect 13165 67809 13223 67855
rect 13269 67809 13291 67855
rect 13097 67751 13291 67809
rect 13097 67705 13119 67751
rect 13165 67705 13223 67751
rect 13269 67705 13291 67751
rect 13097 67647 13291 67705
rect 13097 67601 13119 67647
rect 13165 67601 13223 67647
rect 13269 67601 13291 67647
rect 13097 67543 13291 67601
rect 13097 67497 13119 67543
rect 13165 67497 13223 67543
rect 13269 67497 13291 67543
rect 13097 67439 13291 67497
rect 13097 67393 13119 67439
rect 13165 67393 13223 67439
rect 13269 67393 13291 67439
rect 13097 67335 13291 67393
rect 13097 67289 13119 67335
rect 13165 67289 13223 67335
rect 13269 67289 13291 67335
rect 13097 67231 13291 67289
rect 13097 67185 13119 67231
rect 13165 67185 13223 67231
rect 13269 67185 13291 67231
rect 13097 67127 13291 67185
rect 13097 67081 13119 67127
rect 13165 67081 13223 67127
rect 13269 67081 13291 67127
rect 13097 67023 13291 67081
rect 13097 66977 13119 67023
rect 13165 66977 13223 67023
rect 13269 66977 13291 67023
rect 13097 66919 13291 66977
rect 13097 66873 13119 66919
rect 13165 66873 13223 66919
rect 13269 66873 13291 66919
rect 13097 66815 13291 66873
rect 13097 66769 13119 66815
rect 13165 66769 13223 66815
rect 13269 66769 13291 66815
rect 13097 66711 13291 66769
rect 13097 66665 13119 66711
rect 13165 66665 13223 66711
rect 13269 66665 13291 66711
rect 13097 66607 13291 66665
rect 13097 66561 13119 66607
rect 13165 66561 13223 66607
rect 13269 66561 13291 66607
rect 13097 66503 13291 66561
rect 13097 66457 13119 66503
rect 13165 66457 13223 66503
rect 13269 66457 13291 66503
rect 13097 66399 13291 66457
rect 13097 66353 13119 66399
rect 13165 66353 13223 66399
rect 13269 66353 13291 66399
rect 13097 66295 13291 66353
rect 13097 66249 13119 66295
rect 13165 66249 13223 66295
rect 13269 66249 13291 66295
rect 13097 66191 13291 66249
rect 13097 66145 13119 66191
rect 13165 66145 13223 66191
rect 13269 66145 13291 66191
rect 13097 66087 13291 66145
rect 13097 66041 13119 66087
rect 13165 66041 13223 66087
rect 13269 66041 13291 66087
rect 13097 65983 13291 66041
rect 13097 65937 13119 65983
rect 13165 65937 13223 65983
rect 13269 65937 13291 65983
rect 13097 65879 13291 65937
rect 13097 65833 13119 65879
rect 13165 65833 13223 65879
rect 13269 65833 13291 65879
rect 13097 65775 13291 65833
rect 13097 65729 13119 65775
rect 13165 65729 13223 65775
rect 13269 65729 13291 65775
rect 13097 65671 13291 65729
rect 13097 65625 13119 65671
rect 13165 65625 13223 65671
rect 13269 65625 13291 65671
rect 13097 65567 13291 65625
rect 13097 65521 13119 65567
rect 13165 65521 13223 65567
rect 13269 65521 13291 65567
rect 13097 65463 13291 65521
rect 13097 65417 13119 65463
rect 13165 65417 13223 65463
rect 13269 65417 13291 65463
rect 13097 65359 13291 65417
rect 13097 65313 13119 65359
rect 13165 65313 13223 65359
rect 13269 65313 13291 65359
rect 13097 65255 13291 65313
rect 13097 65209 13119 65255
rect 13165 65209 13223 65255
rect 13269 65209 13291 65255
rect 13097 65151 13291 65209
rect 13097 65105 13119 65151
rect 13165 65105 13223 65151
rect 13269 65105 13291 65151
rect 13097 65047 13291 65105
rect 13097 65001 13119 65047
rect 13165 65001 13223 65047
rect 13269 65001 13291 65047
rect 13097 64943 13291 65001
rect 13097 64897 13119 64943
rect 13165 64897 13223 64943
rect 13269 64897 13291 64943
rect 13097 64839 13291 64897
rect 13097 64793 13119 64839
rect 13165 64793 13223 64839
rect 13269 64793 13291 64839
rect 13097 64735 13291 64793
rect 13097 64689 13119 64735
rect 13165 64689 13223 64735
rect 13269 64689 13291 64735
rect 13097 64631 13291 64689
rect 13097 64585 13119 64631
rect 13165 64585 13223 64631
rect 13269 64585 13291 64631
rect 13097 64527 13291 64585
rect 13097 64481 13119 64527
rect 13165 64481 13223 64527
rect 13269 64481 13291 64527
rect 13097 64423 13291 64481
rect 13097 64377 13119 64423
rect 13165 64377 13223 64423
rect 13269 64377 13291 64423
rect 13097 64319 13291 64377
rect 13097 64273 13119 64319
rect 13165 64273 13223 64319
rect 13269 64273 13291 64319
rect 13097 64215 13291 64273
rect 13097 64169 13119 64215
rect 13165 64169 13223 64215
rect 13269 64169 13291 64215
rect 13097 64111 13291 64169
rect 13097 64065 13119 64111
rect 13165 64065 13223 64111
rect 13269 64065 13291 64111
rect 13097 64007 13291 64065
rect 13097 63961 13119 64007
rect 13165 63961 13223 64007
rect 13269 63961 13291 64007
rect 13097 63903 13291 63961
rect 13097 63857 13119 63903
rect 13165 63857 13223 63903
rect 13269 63857 13291 63903
rect 13097 63799 13291 63857
rect 13097 63753 13119 63799
rect 13165 63753 13223 63799
rect 13269 63753 13291 63799
rect 13097 63695 13291 63753
rect 13097 63649 13119 63695
rect 13165 63649 13223 63695
rect 13269 63649 13291 63695
rect 13097 63591 13291 63649
rect 13097 63545 13119 63591
rect 13165 63545 13223 63591
rect 13269 63545 13291 63591
rect 13097 63487 13291 63545
rect 13097 63441 13119 63487
rect 13165 63441 13223 63487
rect 13269 63441 13291 63487
rect 13097 63383 13291 63441
rect 13097 63337 13119 63383
rect 13165 63337 13223 63383
rect 13269 63337 13291 63383
rect 13097 63279 13291 63337
rect 13097 63233 13119 63279
rect 13165 63233 13223 63279
rect 13269 63233 13291 63279
rect 13097 63175 13291 63233
rect 13097 63129 13119 63175
rect 13165 63129 13223 63175
rect 13269 63129 13291 63175
rect 13097 63071 13291 63129
rect 13097 63025 13119 63071
rect 13165 63025 13223 63071
rect 13269 63025 13291 63071
rect 13097 62967 13291 63025
rect 13097 62921 13119 62967
rect 13165 62921 13223 62967
rect 13269 62921 13291 62967
rect 13097 62863 13291 62921
rect 13097 62817 13119 62863
rect 13165 62817 13223 62863
rect 13269 62817 13291 62863
rect 13097 62759 13291 62817
rect 13097 62713 13119 62759
rect 13165 62713 13223 62759
rect 13269 62713 13291 62759
rect 13097 62655 13291 62713
rect 13097 62609 13119 62655
rect 13165 62609 13223 62655
rect 13269 62609 13291 62655
rect 13097 62551 13291 62609
rect 13097 62505 13119 62551
rect 13165 62505 13223 62551
rect 13269 62505 13291 62551
rect 13097 62447 13291 62505
rect 13097 62401 13119 62447
rect 13165 62401 13223 62447
rect 13269 62401 13291 62447
rect 13097 62343 13291 62401
rect 13097 62297 13119 62343
rect 13165 62297 13223 62343
rect 13269 62297 13291 62343
rect 13097 62239 13291 62297
rect 13097 62193 13119 62239
rect 13165 62193 13223 62239
rect 13269 62193 13291 62239
rect 13097 62135 13291 62193
rect 13097 62089 13119 62135
rect 13165 62089 13223 62135
rect 13269 62089 13291 62135
rect 13097 62031 13291 62089
rect 13097 61985 13119 62031
rect 13165 61985 13223 62031
rect 13269 61985 13291 62031
rect 13097 61927 13291 61985
rect 13097 61881 13119 61927
rect 13165 61881 13223 61927
rect 13269 61881 13291 61927
rect 13097 61823 13291 61881
rect 13097 61777 13119 61823
rect 13165 61777 13223 61823
rect 13269 61777 13291 61823
rect 13097 61719 13291 61777
rect 13097 61673 13119 61719
rect 13165 61673 13223 61719
rect 13269 61673 13291 61719
rect 13097 61615 13291 61673
rect 13097 61569 13119 61615
rect 13165 61569 13223 61615
rect 13269 61569 13291 61615
rect 13097 61511 13291 61569
rect 13097 61465 13119 61511
rect 13165 61465 13223 61511
rect 13269 61465 13291 61511
rect 13097 61407 13291 61465
rect 13097 61361 13119 61407
rect 13165 61361 13223 61407
rect 13269 61361 13291 61407
rect 13097 61303 13291 61361
rect 13097 61257 13119 61303
rect 13165 61257 13223 61303
rect 13269 61257 13291 61303
rect 13097 61199 13291 61257
rect 13097 61153 13119 61199
rect 13165 61153 13223 61199
rect 13269 61153 13291 61199
rect 13097 61095 13291 61153
rect 13097 61049 13119 61095
rect 13165 61049 13223 61095
rect 13269 61049 13291 61095
rect 13097 60991 13291 61049
rect 13097 60945 13119 60991
rect 13165 60945 13223 60991
rect 13269 60945 13291 60991
rect 13097 60887 13291 60945
rect 13097 60841 13119 60887
rect 13165 60841 13223 60887
rect 13269 60841 13291 60887
rect 13097 60783 13291 60841
rect 13097 60737 13119 60783
rect 13165 60737 13223 60783
rect 13269 60737 13291 60783
rect 13097 60679 13291 60737
rect 13097 60633 13119 60679
rect 13165 60633 13223 60679
rect 13269 60633 13291 60679
rect 13097 60575 13291 60633
rect 13097 60529 13119 60575
rect 13165 60529 13223 60575
rect 13269 60529 13291 60575
rect 13097 60471 13291 60529
rect 13097 60425 13119 60471
rect 13165 60425 13223 60471
rect 13269 60425 13291 60471
rect 13097 60367 13291 60425
rect 13097 60321 13119 60367
rect 13165 60321 13223 60367
rect 13269 60321 13291 60367
rect 13097 60263 13291 60321
rect 13097 60217 13119 60263
rect 13165 60217 13223 60263
rect 13269 60217 13291 60263
rect 13097 60159 13291 60217
rect 13097 60113 13119 60159
rect 13165 60113 13223 60159
rect 13269 60113 13291 60159
rect 13097 60055 13291 60113
rect 13097 60009 13119 60055
rect 13165 60009 13223 60055
rect 13269 60009 13291 60055
rect 13097 59951 13291 60009
rect 13097 59905 13119 59951
rect 13165 59905 13223 59951
rect 13269 59905 13291 59951
rect 13097 59847 13291 59905
rect 13097 59801 13119 59847
rect 13165 59801 13223 59847
rect 13269 59801 13291 59847
rect 13097 59743 13291 59801
rect 13097 59697 13119 59743
rect 13165 59697 13223 59743
rect 13269 59697 13291 59743
rect 13097 59639 13291 59697
rect 13097 59593 13119 59639
rect 13165 59593 13223 59639
rect 13269 59593 13291 59639
rect 13097 59535 13291 59593
rect 13097 59489 13119 59535
rect 13165 59489 13223 59535
rect 13269 59489 13291 59535
rect 13097 59431 13291 59489
rect 13097 59385 13119 59431
rect 13165 59385 13223 59431
rect 13269 59385 13291 59431
rect 13097 59327 13291 59385
rect 13097 59281 13119 59327
rect 13165 59281 13223 59327
rect 13269 59281 13291 59327
rect 13097 59223 13291 59281
rect 13097 59177 13119 59223
rect 13165 59177 13223 59223
rect 13269 59177 13291 59223
rect 13097 59119 13291 59177
rect 13097 59073 13119 59119
rect 13165 59073 13223 59119
rect 13269 59073 13291 59119
rect 13097 59015 13291 59073
rect 13097 58969 13119 59015
rect 13165 58969 13223 59015
rect 13269 58969 13291 59015
rect 13097 58911 13291 58969
rect 13097 58865 13119 58911
rect 13165 58865 13223 58911
rect 13269 58865 13291 58911
rect 13097 58807 13291 58865
rect 13097 58761 13119 58807
rect 13165 58761 13223 58807
rect 13269 58761 13291 58807
rect 13097 58703 13291 58761
rect 13097 58657 13119 58703
rect 13165 58657 13223 58703
rect 13269 58657 13291 58703
rect 13097 58599 13291 58657
rect 13097 58553 13119 58599
rect 13165 58553 13223 58599
rect 13269 58553 13291 58599
rect 13097 58495 13291 58553
rect 13097 58449 13119 58495
rect 13165 58449 13223 58495
rect 13269 58449 13291 58495
rect 13097 58391 13291 58449
rect 13097 58345 13119 58391
rect 13165 58345 13223 58391
rect 13269 58345 13291 58391
rect 13097 58287 13291 58345
rect 13097 58241 13119 58287
rect 13165 58241 13223 58287
rect 13269 58241 13291 58287
rect 13097 58183 13291 58241
rect 13097 58137 13119 58183
rect 13165 58137 13223 58183
rect 13269 58137 13291 58183
rect 13097 58079 13291 58137
rect 13097 58033 13119 58079
rect 13165 58033 13223 58079
rect 13269 58033 13291 58079
rect 13097 57975 13291 58033
rect 13097 57929 13119 57975
rect 13165 57929 13223 57975
rect 13269 57929 13291 57975
rect 13097 57871 13291 57929
rect 13097 57825 13119 57871
rect 13165 57825 13223 57871
rect 13269 57825 13291 57871
rect 13097 57767 13291 57825
rect 13097 57721 13119 57767
rect 13165 57721 13223 57767
rect 13269 57721 13291 57767
rect 13097 57663 13291 57721
rect 13097 57617 13119 57663
rect 13165 57617 13223 57663
rect 13269 57617 13291 57663
rect 13097 57559 13291 57617
rect 13097 57513 13119 57559
rect 13165 57513 13223 57559
rect 13269 57513 13291 57559
rect 13097 57455 13291 57513
rect 13097 57409 13119 57455
rect 13165 57409 13223 57455
rect 13269 57409 13291 57455
rect 13097 57351 13291 57409
rect 13097 57305 13119 57351
rect 13165 57305 13223 57351
rect 13269 57305 13291 57351
rect 13097 57247 13291 57305
rect 13097 57201 13119 57247
rect 13165 57201 13223 57247
rect 13269 57201 13291 57247
rect 13097 57143 13291 57201
rect 13097 57097 13119 57143
rect 13165 57097 13223 57143
rect 13269 57097 13291 57143
rect 13097 57039 13291 57097
rect 13097 56993 13119 57039
rect 13165 56993 13223 57039
rect 13269 56993 13291 57039
rect 13097 56935 13291 56993
rect 13097 56889 13119 56935
rect 13165 56889 13223 56935
rect 13269 56889 13291 56935
rect 13097 56831 13291 56889
rect 13097 56785 13119 56831
rect 13165 56785 13223 56831
rect 13269 56785 13291 56831
rect 13097 56727 13291 56785
rect 13097 56681 13119 56727
rect 13165 56681 13223 56727
rect 13269 56681 13291 56727
rect 13097 56623 13291 56681
rect 13097 56577 13119 56623
rect 13165 56577 13223 56623
rect 13269 56577 13291 56623
rect 13097 56519 13291 56577
rect 13097 56473 13119 56519
rect 13165 56473 13223 56519
rect 13269 56473 13291 56519
rect 13097 56415 13291 56473
rect 13097 56369 13119 56415
rect 13165 56369 13223 56415
rect 13269 56369 13291 56415
rect 13097 56311 13291 56369
rect 13097 56265 13119 56311
rect 13165 56265 13223 56311
rect 13269 56265 13291 56311
rect 13097 56207 13291 56265
rect 13097 56161 13119 56207
rect 13165 56161 13223 56207
rect 13269 56161 13291 56207
rect 13097 56103 13291 56161
rect 13097 56057 13119 56103
rect 13165 56057 13223 56103
rect 13269 56057 13291 56103
rect 13097 55999 13291 56057
rect 13097 55953 13119 55999
rect 13165 55953 13223 55999
rect 13269 55953 13291 55999
rect 13097 55895 13291 55953
rect 13097 55849 13119 55895
rect 13165 55849 13223 55895
rect 13269 55849 13291 55895
rect 13097 55791 13291 55849
rect 13097 55745 13119 55791
rect 13165 55745 13223 55791
rect 13269 55745 13291 55791
rect 13097 55687 13291 55745
rect 13097 55641 13119 55687
rect 13165 55641 13223 55687
rect 13269 55641 13291 55687
rect 13097 55583 13291 55641
rect 13097 55537 13119 55583
rect 13165 55537 13223 55583
rect 13269 55537 13291 55583
rect 13097 55479 13291 55537
rect 13097 55433 13119 55479
rect 13165 55433 13223 55479
rect 13269 55433 13291 55479
rect 13097 55375 13291 55433
rect 13097 55329 13119 55375
rect 13165 55329 13223 55375
rect 13269 55329 13291 55375
rect 13097 55271 13291 55329
rect 13097 55225 13119 55271
rect 13165 55225 13223 55271
rect 13269 55225 13291 55271
rect 13097 55167 13291 55225
rect 13097 55121 13119 55167
rect 13165 55121 13223 55167
rect 13269 55121 13291 55167
rect 13097 55063 13291 55121
rect 13097 55017 13119 55063
rect 13165 55017 13223 55063
rect 13269 55017 13291 55063
rect 13097 54959 13291 55017
rect 13097 54913 13119 54959
rect 13165 54913 13223 54959
rect 13269 54913 13291 54959
rect 13097 54855 13291 54913
rect 13097 54809 13119 54855
rect 13165 54809 13223 54855
rect 13269 54809 13291 54855
rect 13097 54751 13291 54809
rect 13097 54705 13119 54751
rect 13165 54705 13223 54751
rect 13269 54705 13291 54751
rect 13097 54647 13291 54705
rect 13097 54601 13119 54647
rect 13165 54601 13223 54647
rect 13269 54601 13291 54647
rect 13097 54543 13291 54601
rect 13097 54497 13119 54543
rect 13165 54497 13223 54543
rect 13269 54497 13291 54543
rect 13097 54439 13291 54497
rect 13097 54393 13119 54439
rect 13165 54393 13223 54439
rect 13269 54393 13291 54439
rect 13097 54335 13291 54393
rect 13097 54289 13119 54335
rect 13165 54289 13223 54335
rect 13269 54289 13291 54335
rect 13097 54231 13291 54289
rect 13097 54185 13119 54231
rect 13165 54185 13223 54231
rect 13269 54185 13291 54231
rect 13097 54127 13291 54185
rect 13097 54081 13119 54127
rect 13165 54081 13223 54127
rect 13269 54081 13291 54127
rect 13097 54023 13291 54081
rect 13097 53977 13119 54023
rect 13165 53977 13223 54023
rect 13269 53977 13291 54023
rect 13097 53919 13291 53977
rect 13097 53873 13119 53919
rect 13165 53873 13223 53919
rect 13269 53873 13291 53919
rect 13097 53815 13291 53873
rect 13097 53769 13119 53815
rect 13165 53769 13223 53815
rect 13269 53769 13291 53815
rect 13097 53711 13291 53769
rect 13097 53665 13119 53711
rect 13165 53665 13223 53711
rect 13269 53665 13291 53711
rect 13097 53607 13291 53665
rect 13097 53561 13119 53607
rect 13165 53561 13223 53607
rect 13269 53561 13291 53607
rect 13097 53503 13291 53561
rect 13097 53457 13119 53503
rect 13165 53457 13223 53503
rect 13269 53457 13291 53503
rect 13097 53399 13291 53457
rect 13097 53353 13119 53399
rect 13165 53353 13223 53399
rect 13269 53353 13291 53399
rect 13097 53295 13291 53353
rect 13097 53249 13119 53295
rect 13165 53249 13223 53295
rect 13269 53249 13291 53295
rect 13097 53191 13291 53249
rect 13097 53145 13119 53191
rect 13165 53145 13223 53191
rect 13269 53145 13291 53191
rect 13097 53087 13291 53145
rect 13097 53041 13119 53087
rect 13165 53041 13223 53087
rect 13269 53041 13291 53087
rect 13097 52983 13291 53041
rect 13097 52937 13119 52983
rect 13165 52937 13223 52983
rect 13269 52937 13291 52983
rect 13097 52879 13291 52937
rect 13097 52833 13119 52879
rect 13165 52833 13223 52879
rect 13269 52833 13291 52879
rect 13097 52775 13291 52833
rect 13097 52729 13119 52775
rect 13165 52729 13223 52775
rect 13269 52729 13291 52775
rect 13097 52671 13291 52729
rect 13097 52625 13119 52671
rect 13165 52625 13223 52671
rect 13269 52625 13291 52671
rect 13097 52567 13291 52625
rect 13097 52521 13119 52567
rect 13165 52521 13223 52567
rect 13269 52521 13291 52567
rect 13097 52463 13291 52521
rect 13097 52417 13119 52463
rect 13165 52417 13223 52463
rect 13269 52417 13291 52463
rect 13097 52359 13291 52417
rect 13097 52313 13119 52359
rect 13165 52313 13223 52359
rect 13269 52313 13291 52359
rect 13097 52255 13291 52313
rect 13097 52209 13119 52255
rect 13165 52209 13223 52255
rect 13269 52209 13291 52255
rect 13097 52151 13291 52209
rect 13097 52105 13119 52151
rect 13165 52105 13223 52151
rect 13269 52105 13291 52151
rect 13097 52047 13291 52105
rect 13097 52001 13119 52047
rect 13165 52001 13223 52047
rect 13269 52001 13291 52047
rect 13097 51943 13291 52001
rect 13097 51897 13119 51943
rect 13165 51897 13223 51943
rect 13269 51897 13291 51943
rect 13097 51839 13291 51897
rect 13097 51793 13119 51839
rect 13165 51793 13223 51839
rect 13269 51793 13291 51839
rect 13097 51735 13291 51793
rect 13097 51689 13119 51735
rect 13165 51689 13223 51735
rect 13269 51689 13291 51735
rect 13097 51631 13291 51689
rect 13097 51585 13119 51631
rect 13165 51585 13223 51631
rect 13269 51585 13291 51631
rect 13097 51527 13291 51585
rect 13097 51481 13119 51527
rect 13165 51481 13223 51527
rect 13269 51481 13291 51527
rect 13097 51423 13291 51481
rect 13097 51377 13119 51423
rect 13165 51377 13223 51423
rect 13269 51377 13291 51423
rect 13097 51319 13291 51377
rect 13097 51273 13119 51319
rect 13165 51273 13223 51319
rect 13269 51273 13291 51319
rect 13097 51215 13291 51273
rect 13097 51169 13119 51215
rect 13165 51169 13223 51215
rect 13269 51169 13291 51215
rect 13097 51111 13291 51169
rect 13097 51065 13119 51111
rect 13165 51065 13223 51111
rect 13269 51065 13291 51111
rect 13097 51007 13291 51065
rect 13097 50961 13119 51007
rect 13165 50961 13223 51007
rect 13269 50961 13291 51007
rect 13097 50903 13291 50961
rect 13097 50857 13119 50903
rect 13165 50857 13223 50903
rect 13269 50857 13291 50903
rect 13097 50799 13291 50857
rect 13097 50753 13119 50799
rect 13165 50753 13223 50799
rect 13269 50753 13291 50799
rect 13097 50695 13291 50753
rect 13097 50649 13119 50695
rect 13165 50649 13223 50695
rect 13269 50649 13291 50695
rect 13097 50591 13291 50649
rect 13097 50545 13119 50591
rect 13165 50545 13223 50591
rect 13269 50545 13291 50591
rect 13097 50487 13291 50545
rect 13097 50441 13119 50487
rect 13165 50441 13223 50487
rect 13269 50441 13291 50487
rect 13097 50383 13291 50441
rect 13097 50337 13119 50383
rect 13165 50337 13223 50383
rect 13269 50337 13291 50383
rect 13097 50279 13291 50337
rect 13097 50233 13119 50279
rect 13165 50233 13223 50279
rect 13269 50233 13291 50279
rect 13097 50175 13291 50233
rect 13097 50129 13119 50175
rect 13165 50129 13223 50175
rect 13269 50129 13291 50175
rect 13097 50071 13291 50129
rect 13097 50025 13119 50071
rect 13165 50025 13223 50071
rect 13269 50025 13291 50071
rect 13097 49967 13291 50025
rect 13097 49921 13119 49967
rect 13165 49921 13223 49967
rect 13269 49921 13291 49967
rect 13097 49863 13291 49921
rect 13097 49817 13119 49863
rect 13165 49817 13223 49863
rect 13269 49817 13291 49863
rect 13097 49759 13291 49817
rect 13097 49713 13119 49759
rect 13165 49713 13223 49759
rect 13269 49713 13291 49759
rect 13097 49655 13291 49713
rect 13097 49609 13119 49655
rect 13165 49609 13223 49655
rect 13269 49609 13291 49655
rect 13097 49551 13291 49609
rect 13097 49505 13119 49551
rect 13165 49505 13223 49551
rect 13269 49505 13291 49551
rect 13097 49447 13291 49505
rect 13097 49401 13119 49447
rect 13165 49401 13223 49447
rect 13269 49401 13291 49447
rect 13097 49343 13291 49401
rect 13097 49297 13119 49343
rect 13165 49297 13223 49343
rect 13269 49297 13291 49343
rect 13097 49239 13291 49297
rect 13097 49193 13119 49239
rect 13165 49193 13223 49239
rect 13269 49193 13291 49239
rect 13097 49135 13291 49193
rect 13097 49089 13119 49135
rect 13165 49089 13223 49135
rect 13269 49089 13291 49135
rect 13097 49031 13291 49089
rect 13097 48985 13119 49031
rect 13165 48985 13223 49031
rect 13269 48985 13291 49031
rect 13097 48927 13291 48985
rect 13097 48881 13119 48927
rect 13165 48881 13223 48927
rect 13269 48881 13291 48927
rect 13097 48823 13291 48881
rect 13097 48777 13119 48823
rect 13165 48777 13223 48823
rect 13269 48777 13291 48823
rect 13097 48719 13291 48777
rect 13097 48673 13119 48719
rect 13165 48673 13223 48719
rect 13269 48673 13291 48719
rect 13097 48615 13291 48673
rect 13097 48569 13119 48615
rect 13165 48569 13223 48615
rect 13269 48569 13291 48615
rect 13097 48511 13291 48569
rect 13097 48465 13119 48511
rect 13165 48465 13223 48511
rect 13269 48465 13291 48511
rect 13097 48407 13291 48465
rect 13097 48361 13119 48407
rect 13165 48361 13223 48407
rect 13269 48361 13291 48407
rect 13097 48303 13291 48361
rect 13097 48257 13119 48303
rect 13165 48257 13223 48303
rect 13269 48257 13291 48303
rect 13097 48199 13291 48257
rect 13097 48153 13119 48199
rect 13165 48153 13223 48199
rect 13269 48153 13291 48199
rect 13097 48095 13291 48153
rect 13097 48049 13119 48095
rect 13165 48049 13223 48095
rect 13269 48049 13291 48095
rect 13097 47991 13291 48049
rect 13097 47945 13119 47991
rect 13165 47945 13223 47991
rect 13269 47945 13291 47991
rect 13097 47887 13291 47945
rect 13097 47841 13119 47887
rect 13165 47841 13223 47887
rect 13269 47841 13291 47887
rect 13097 47783 13291 47841
rect 13097 47737 13119 47783
rect 13165 47737 13223 47783
rect 13269 47737 13291 47783
rect 13097 47679 13291 47737
rect 13097 47633 13119 47679
rect 13165 47633 13223 47679
rect 13269 47633 13291 47679
rect 13097 47575 13291 47633
rect 13097 47529 13119 47575
rect 13165 47529 13223 47575
rect 13269 47529 13291 47575
rect 13097 47471 13291 47529
rect 13097 47425 13119 47471
rect 13165 47425 13223 47471
rect 13269 47425 13291 47471
rect 13097 47367 13291 47425
rect 13097 47321 13119 47367
rect 13165 47321 13223 47367
rect 13269 47321 13291 47367
rect 13097 47263 13291 47321
rect 13097 47217 13119 47263
rect 13165 47217 13223 47263
rect 13269 47217 13291 47263
rect 13097 47159 13291 47217
rect 13097 47113 13119 47159
rect 13165 47113 13223 47159
rect 13269 47113 13291 47159
rect 13097 47055 13291 47113
rect 13097 47009 13119 47055
rect 13165 47009 13223 47055
rect 13269 47009 13291 47055
rect 13097 46951 13291 47009
rect 13097 46905 13119 46951
rect 13165 46905 13223 46951
rect 13269 46905 13291 46951
rect 13097 46847 13291 46905
rect 13097 46801 13119 46847
rect 13165 46801 13223 46847
rect 13269 46801 13291 46847
rect 13097 46743 13291 46801
rect 13097 46697 13119 46743
rect 13165 46697 13223 46743
rect 13269 46697 13291 46743
rect 13097 46639 13291 46697
rect 13097 46593 13119 46639
rect 13165 46593 13223 46639
rect 13269 46593 13291 46639
rect 13097 46535 13291 46593
rect 13097 46489 13119 46535
rect 13165 46489 13223 46535
rect 13269 46489 13291 46535
rect 13097 46431 13291 46489
rect 13097 46385 13119 46431
rect 13165 46385 13223 46431
rect 13269 46385 13291 46431
rect 13097 46327 13291 46385
rect 13097 46281 13119 46327
rect 13165 46281 13223 46327
rect 13269 46281 13291 46327
rect 13097 46223 13291 46281
rect 13097 46177 13119 46223
rect 13165 46177 13223 46223
rect 13269 46177 13291 46223
rect 13097 46119 13291 46177
rect 13097 46073 13119 46119
rect 13165 46073 13223 46119
rect 13269 46073 13291 46119
rect 13097 46015 13291 46073
rect 13097 45969 13119 46015
rect 13165 45969 13223 46015
rect 13269 45969 13291 46015
rect 13097 45911 13291 45969
rect 13097 45865 13119 45911
rect 13165 45865 13223 45911
rect 13269 45865 13291 45911
rect 13097 45807 13291 45865
rect 13097 45761 13119 45807
rect 13165 45761 13223 45807
rect 13269 45761 13291 45807
rect 13097 45703 13291 45761
rect 13097 45657 13119 45703
rect 13165 45657 13223 45703
rect 13269 45657 13291 45703
rect 13097 45599 13291 45657
rect 13097 45553 13119 45599
rect 13165 45553 13223 45599
rect 13269 45553 13291 45599
rect 13097 45495 13291 45553
rect 13097 45449 13119 45495
rect 13165 45449 13223 45495
rect 13269 45449 13291 45495
rect 13097 45391 13291 45449
rect 13097 45345 13119 45391
rect 13165 45345 13223 45391
rect 13269 45345 13291 45391
rect 13097 45287 13291 45345
rect 13097 45241 13119 45287
rect 13165 45241 13223 45287
rect 13269 45241 13291 45287
rect 13097 45183 13291 45241
rect 13097 45137 13119 45183
rect 13165 45137 13223 45183
rect 13269 45137 13291 45183
rect 13097 45079 13291 45137
rect 13097 45033 13119 45079
rect 13165 45033 13223 45079
rect 13269 45033 13291 45079
rect 13097 44892 13291 45033
rect 70802 69758 70824 69774
rect 70870 69758 70928 69804
rect 70974 69758 71000 69804
rect 70802 69700 71000 69758
rect 70802 69654 70824 69700
rect 70870 69654 70928 69700
rect 70974 69654 71000 69700
rect 70802 69596 71000 69654
rect 70802 69550 70824 69596
rect 70870 69550 70928 69596
rect 70974 69550 71000 69596
rect 70802 69492 71000 69550
rect 70802 69446 70824 69492
rect 70870 69446 70928 69492
rect 70974 69446 71000 69492
rect 70802 69388 71000 69446
rect 70802 69342 70824 69388
rect 70870 69342 70928 69388
rect 70974 69342 71000 69388
rect 70802 69284 71000 69342
rect 70802 69238 70824 69284
rect 70870 69238 70928 69284
rect 70974 69238 71000 69284
rect 70802 69180 71000 69238
rect 70802 69134 70824 69180
rect 70870 69134 70928 69180
rect 70974 69134 71000 69180
rect 70802 69076 71000 69134
rect 70802 69030 70824 69076
rect 70870 69030 70928 69076
rect 70974 69030 71000 69076
rect 70802 68972 71000 69030
rect 70802 68926 70824 68972
rect 70870 68926 70928 68972
rect 70974 68926 71000 68972
rect 70802 68868 71000 68926
rect 70802 68822 70824 68868
rect 70870 68822 70928 68868
rect 70974 68822 71000 68868
rect 70802 68764 71000 68822
rect 70802 68718 70824 68764
rect 70870 68718 70928 68764
rect 70974 68718 71000 68764
rect 70802 68660 71000 68718
rect 70802 68614 70824 68660
rect 70870 68614 70928 68660
rect 70974 68614 71000 68660
rect 70802 68556 71000 68614
rect 70802 68510 70824 68556
rect 70870 68510 70928 68556
rect 70974 68510 71000 68556
rect 70802 68452 71000 68510
rect 70802 68406 70824 68452
rect 70870 68406 70928 68452
rect 70974 68406 71000 68452
rect 70802 68348 71000 68406
rect 70802 68302 70824 68348
rect 70870 68302 70928 68348
rect 70974 68302 71000 68348
rect 70802 68244 71000 68302
rect 70802 68198 70824 68244
rect 70870 68198 70928 68244
rect 70974 68198 71000 68244
rect 70802 68140 71000 68198
rect 70802 68094 70824 68140
rect 70870 68094 70928 68140
rect 70974 68094 71000 68140
rect 70802 68036 71000 68094
rect 70802 67990 70824 68036
rect 70870 67990 70928 68036
rect 70974 67990 71000 68036
rect 70802 67932 71000 67990
rect 70802 67886 70824 67932
rect 70870 67886 70928 67932
rect 70974 67886 71000 67932
rect 70802 67828 71000 67886
rect 70802 67782 70824 67828
rect 70870 67782 70928 67828
rect 70974 67782 71000 67828
rect 70802 67724 71000 67782
rect 70802 67678 70824 67724
rect 70870 67678 70928 67724
rect 70974 67678 71000 67724
rect 70802 67620 71000 67678
rect 70802 67574 70824 67620
rect 70870 67574 70928 67620
rect 70974 67574 71000 67620
rect 70802 67516 71000 67574
rect 70802 67470 70824 67516
rect 70870 67470 70928 67516
rect 70974 67470 71000 67516
rect 70802 67412 71000 67470
rect 70802 67366 70824 67412
rect 70870 67366 70928 67412
rect 70974 67366 71000 67412
rect 70802 67308 71000 67366
rect 70802 67262 70824 67308
rect 70870 67262 70928 67308
rect 70974 67262 71000 67308
rect 70802 67204 71000 67262
rect 70802 67158 70824 67204
rect 70870 67158 70928 67204
rect 70974 67158 71000 67204
rect 70802 67100 71000 67158
rect 70802 67054 70824 67100
rect 70870 67054 70928 67100
rect 70974 67054 71000 67100
rect 70802 66996 71000 67054
rect 70802 66950 70824 66996
rect 70870 66950 70928 66996
rect 70974 66950 71000 66996
rect 70802 66892 71000 66950
rect 70802 66846 70824 66892
rect 70870 66846 70928 66892
rect 70974 66846 71000 66892
rect 70802 66788 71000 66846
rect 70802 66742 70824 66788
rect 70870 66742 70928 66788
rect 70974 66742 71000 66788
rect 70802 66684 71000 66742
rect 70802 66638 70824 66684
rect 70870 66638 70928 66684
rect 70974 66638 71000 66684
rect 70802 66580 71000 66638
rect 70802 66534 70824 66580
rect 70870 66534 70928 66580
rect 70974 66534 71000 66580
rect 70802 66476 71000 66534
rect 70802 66430 70824 66476
rect 70870 66430 70928 66476
rect 70974 66430 71000 66476
rect 70802 66372 71000 66430
rect 70802 66326 70824 66372
rect 70870 66326 70928 66372
rect 70974 66326 71000 66372
rect 70802 66268 71000 66326
rect 70802 66222 70824 66268
rect 70870 66222 70928 66268
rect 70974 66222 71000 66268
rect 70802 66164 71000 66222
rect 70802 66118 70824 66164
rect 70870 66118 70928 66164
rect 70974 66118 71000 66164
rect 70802 66060 71000 66118
rect 70802 66014 70824 66060
rect 70870 66014 70928 66060
rect 70974 66014 71000 66060
rect 70802 65956 71000 66014
rect 70802 65910 70824 65956
rect 70870 65910 70928 65956
rect 70974 65910 71000 65956
rect 70802 65852 71000 65910
rect 70802 65806 70824 65852
rect 70870 65806 70928 65852
rect 70974 65806 71000 65852
rect 70802 65748 71000 65806
rect 70802 65702 70824 65748
rect 70870 65702 70928 65748
rect 70974 65702 71000 65748
rect 70802 65644 71000 65702
rect 70802 65598 70824 65644
rect 70870 65598 70928 65644
rect 70974 65598 71000 65644
rect 70802 65540 71000 65598
rect 70802 65494 70824 65540
rect 70870 65494 70928 65540
rect 70974 65494 71000 65540
rect 70802 65436 71000 65494
rect 70802 65390 70824 65436
rect 70870 65390 70928 65436
rect 70974 65390 71000 65436
rect 70802 65332 71000 65390
rect 70802 65286 70824 65332
rect 70870 65286 70928 65332
rect 70974 65286 71000 65332
rect 70802 65228 71000 65286
rect 70802 65182 70824 65228
rect 70870 65182 70928 65228
rect 70974 65182 71000 65228
rect 70802 65124 71000 65182
rect 70802 65078 70824 65124
rect 70870 65078 70928 65124
rect 70974 65078 71000 65124
rect 70802 65020 71000 65078
rect 70802 64974 70824 65020
rect 70870 64974 70928 65020
rect 70974 64974 71000 65020
rect 70802 64916 71000 64974
rect 70802 64870 70824 64916
rect 70870 64870 70928 64916
rect 70974 64870 71000 64916
rect 70802 64812 71000 64870
rect 70802 64766 70824 64812
rect 70870 64766 70928 64812
rect 70974 64766 71000 64812
rect 70802 64708 71000 64766
rect 70802 64662 70824 64708
rect 70870 64662 70928 64708
rect 70974 64662 71000 64708
rect 70802 64604 71000 64662
rect 70802 64558 70824 64604
rect 70870 64558 70928 64604
rect 70974 64558 71000 64604
rect 70802 64500 71000 64558
rect 70802 64454 70824 64500
rect 70870 64454 70928 64500
rect 70974 64454 71000 64500
rect 70802 64396 71000 64454
rect 70802 64350 70824 64396
rect 70870 64350 70928 64396
rect 70974 64350 71000 64396
rect 70802 64292 71000 64350
rect 70802 64246 70824 64292
rect 70870 64246 70928 64292
rect 70974 64246 71000 64292
rect 70802 64188 71000 64246
rect 70802 64142 70824 64188
rect 70870 64142 70928 64188
rect 70974 64142 71000 64188
rect 70802 64084 71000 64142
rect 70802 64038 70824 64084
rect 70870 64038 70928 64084
rect 70974 64038 71000 64084
rect 70802 63980 71000 64038
rect 70802 63934 70824 63980
rect 70870 63934 70928 63980
rect 70974 63934 71000 63980
rect 70802 63876 71000 63934
rect 70802 63830 70824 63876
rect 70870 63830 70928 63876
rect 70974 63830 71000 63876
rect 70802 63772 71000 63830
rect 70802 63726 70824 63772
rect 70870 63726 70928 63772
rect 70974 63726 71000 63772
rect 70802 63668 71000 63726
rect 70802 63622 70824 63668
rect 70870 63622 70928 63668
rect 70974 63622 71000 63668
rect 70802 63564 71000 63622
rect 70802 63518 70824 63564
rect 70870 63518 70928 63564
rect 70974 63518 71000 63564
rect 70802 63460 71000 63518
rect 70802 63414 70824 63460
rect 70870 63414 70928 63460
rect 70974 63414 71000 63460
rect 70802 63356 71000 63414
rect 70802 63310 70824 63356
rect 70870 63310 70928 63356
rect 70974 63310 71000 63356
rect 70802 63252 71000 63310
rect 70802 63206 70824 63252
rect 70870 63206 70928 63252
rect 70974 63206 71000 63252
rect 70802 63148 71000 63206
rect 70802 63102 70824 63148
rect 70870 63102 70928 63148
rect 70974 63102 71000 63148
rect 70802 63044 71000 63102
rect 70802 62998 70824 63044
rect 70870 62998 70928 63044
rect 70974 62998 71000 63044
rect 70802 62940 71000 62998
rect 70802 62894 70824 62940
rect 70870 62894 70928 62940
rect 70974 62894 71000 62940
rect 70802 62836 71000 62894
rect 70802 62790 70824 62836
rect 70870 62790 70928 62836
rect 70974 62790 71000 62836
rect 70802 62732 71000 62790
rect 70802 62686 70824 62732
rect 70870 62686 70928 62732
rect 70974 62686 71000 62732
rect 70802 62628 71000 62686
rect 70802 62582 70824 62628
rect 70870 62582 70928 62628
rect 70974 62582 71000 62628
rect 70802 62524 71000 62582
rect 70802 62478 70824 62524
rect 70870 62478 70928 62524
rect 70974 62478 71000 62524
rect 70802 62420 71000 62478
rect 70802 62374 70824 62420
rect 70870 62374 70928 62420
rect 70974 62374 71000 62420
rect 70802 62316 71000 62374
rect 70802 62270 70824 62316
rect 70870 62270 70928 62316
rect 70974 62270 71000 62316
rect 70802 62212 71000 62270
rect 70802 62166 70824 62212
rect 70870 62166 70928 62212
rect 70974 62166 71000 62212
rect 70802 62108 71000 62166
rect 70802 62062 70824 62108
rect 70870 62062 70928 62108
rect 70974 62062 71000 62108
rect 70802 62004 71000 62062
rect 70802 61958 70824 62004
rect 70870 61958 70928 62004
rect 70974 61958 71000 62004
rect 70802 61900 71000 61958
rect 70802 61854 70824 61900
rect 70870 61854 70928 61900
rect 70974 61854 71000 61900
rect 70802 61796 71000 61854
rect 70802 61750 70824 61796
rect 70870 61750 70928 61796
rect 70974 61750 71000 61796
rect 70802 61692 71000 61750
rect 70802 61646 70824 61692
rect 70870 61646 70928 61692
rect 70974 61646 71000 61692
rect 70802 61588 71000 61646
rect 70802 61542 70824 61588
rect 70870 61542 70928 61588
rect 70974 61542 71000 61588
rect 70802 61484 71000 61542
rect 70802 61438 70824 61484
rect 70870 61438 70928 61484
rect 70974 61438 71000 61484
rect 70802 61380 71000 61438
rect 70802 61334 70824 61380
rect 70870 61334 70928 61380
rect 70974 61334 71000 61380
rect 70802 61276 71000 61334
rect 70802 61230 70824 61276
rect 70870 61230 70928 61276
rect 70974 61230 71000 61276
rect 70802 61172 71000 61230
rect 70802 61126 70824 61172
rect 70870 61126 70928 61172
rect 70974 61126 71000 61172
rect 70802 61068 71000 61126
rect 70802 61022 70824 61068
rect 70870 61022 70928 61068
rect 70974 61022 71000 61068
rect 70802 60964 71000 61022
rect 70802 60918 70824 60964
rect 70870 60918 70928 60964
rect 70974 60918 71000 60964
rect 70802 60860 71000 60918
rect 70802 60814 70824 60860
rect 70870 60814 70928 60860
rect 70974 60814 71000 60860
rect 70802 60756 71000 60814
rect 70802 60710 70824 60756
rect 70870 60710 70928 60756
rect 70974 60710 71000 60756
rect 70802 60652 71000 60710
rect 70802 60606 70824 60652
rect 70870 60606 70928 60652
rect 70974 60606 71000 60652
rect 70802 60548 71000 60606
rect 70802 60502 70824 60548
rect 70870 60502 70928 60548
rect 70974 60502 71000 60548
rect 70802 60444 71000 60502
rect 70802 60398 70824 60444
rect 70870 60398 70928 60444
rect 70974 60398 71000 60444
rect 70802 60340 71000 60398
rect 70802 60294 70824 60340
rect 70870 60294 70928 60340
rect 70974 60294 71000 60340
rect 70802 60236 71000 60294
rect 70802 60190 70824 60236
rect 70870 60190 70928 60236
rect 70974 60190 71000 60236
rect 70802 60132 71000 60190
rect 70802 60086 70824 60132
rect 70870 60086 70928 60132
rect 70974 60086 71000 60132
rect 70802 60028 71000 60086
rect 70802 59982 70824 60028
rect 70870 59982 70928 60028
rect 70974 59982 71000 60028
rect 70802 59924 71000 59982
rect 70802 59878 70824 59924
rect 70870 59878 70928 59924
rect 70974 59878 71000 59924
rect 70802 59820 71000 59878
rect 70802 59774 70824 59820
rect 70870 59774 70928 59820
rect 70974 59774 71000 59820
rect 70802 59716 71000 59774
rect 70802 59670 70824 59716
rect 70870 59670 70928 59716
rect 70974 59670 71000 59716
rect 70802 59612 71000 59670
rect 70802 59566 70824 59612
rect 70870 59566 70928 59612
rect 70974 59566 71000 59612
rect 70802 59508 71000 59566
rect 70802 59462 70824 59508
rect 70870 59462 70928 59508
rect 70974 59462 71000 59508
rect 70802 59404 71000 59462
rect 70802 59358 70824 59404
rect 70870 59358 70928 59404
rect 70974 59358 71000 59404
rect 70802 59300 71000 59358
rect 70802 59254 70824 59300
rect 70870 59254 70928 59300
rect 70974 59254 71000 59300
rect 70802 59196 71000 59254
rect 70802 59150 70824 59196
rect 70870 59150 70928 59196
rect 70974 59150 71000 59196
rect 70802 59092 71000 59150
rect 70802 59046 70824 59092
rect 70870 59046 70928 59092
rect 70974 59046 71000 59092
rect 70802 58988 71000 59046
rect 70802 58942 70824 58988
rect 70870 58942 70928 58988
rect 70974 58942 71000 58988
rect 70802 58884 71000 58942
rect 70802 58838 70824 58884
rect 70870 58838 70928 58884
rect 70974 58838 71000 58884
rect 70802 58780 71000 58838
rect 70802 58734 70824 58780
rect 70870 58734 70928 58780
rect 70974 58734 71000 58780
rect 70802 58676 71000 58734
rect 70802 58630 70824 58676
rect 70870 58630 70928 58676
rect 70974 58630 71000 58676
rect 70802 58572 71000 58630
rect 70802 58526 70824 58572
rect 70870 58526 70928 58572
rect 70974 58526 71000 58572
rect 70802 58468 71000 58526
rect 70802 58422 70824 58468
rect 70870 58422 70928 58468
rect 70974 58422 71000 58468
rect 70802 58364 71000 58422
rect 70802 58318 70824 58364
rect 70870 58318 70928 58364
rect 70974 58318 71000 58364
rect 70802 58260 71000 58318
rect 70802 58214 70824 58260
rect 70870 58214 70928 58260
rect 70974 58214 71000 58260
rect 70802 58156 71000 58214
rect 70802 58110 70824 58156
rect 70870 58110 70928 58156
rect 70974 58110 71000 58156
rect 70802 58052 71000 58110
rect 70802 58006 70824 58052
rect 70870 58006 70928 58052
rect 70974 58006 71000 58052
rect 70802 57948 71000 58006
rect 70802 57902 70824 57948
rect 70870 57902 70928 57948
rect 70974 57902 71000 57948
rect 70802 57844 71000 57902
rect 70802 57798 70824 57844
rect 70870 57798 70928 57844
rect 70974 57798 71000 57844
rect 70802 57740 71000 57798
rect 70802 57694 70824 57740
rect 70870 57694 70928 57740
rect 70974 57694 71000 57740
rect 70802 57636 71000 57694
rect 70802 57590 70824 57636
rect 70870 57590 70928 57636
rect 70974 57590 71000 57636
rect 70802 57532 71000 57590
rect 70802 57486 70824 57532
rect 70870 57486 70928 57532
rect 70974 57486 71000 57532
rect 70802 57428 71000 57486
rect 70802 57382 70824 57428
rect 70870 57382 70928 57428
rect 70974 57382 71000 57428
rect 70802 57324 71000 57382
rect 70802 57278 70824 57324
rect 70870 57278 70928 57324
rect 70974 57278 71000 57324
rect 70802 57220 71000 57278
rect 70802 57174 70824 57220
rect 70870 57174 70928 57220
rect 70974 57174 71000 57220
rect 70802 57116 71000 57174
rect 70802 57070 70824 57116
rect 70870 57070 70928 57116
rect 70974 57070 71000 57116
rect 70802 57012 71000 57070
rect 70802 56966 70824 57012
rect 70870 56966 70928 57012
rect 70974 56966 71000 57012
rect 70802 56908 71000 56966
rect 70802 56862 70824 56908
rect 70870 56862 70928 56908
rect 70974 56862 71000 56908
rect 70802 56804 71000 56862
rect 70802 56758 70824 56804
rect 70870 56758 70928 56804
rect 70974 56758 71000 56804
rect 70802 56700 71000 56758
rect 70802 56654 70824 56700
rect 70870 56654 70928 56700
rect 70974 56654 71000 56700
rect 70802 56596 71000 56654
rect 70802 56550 70824 56596
rect 70870 56550 70928 56596
rect 70974 56550 71000 56596
rect 70802 56492 71000 56550
rect 70802 56446 70824 56492
rect 70870 56446 70928 56492
rect 70974 56446 71000 56492
rect 70802 56388 71000 56446
rect 70802 56342 70824 56388
rect 70870 56342 70928 56388
rect 70974 56342 71000 56388
rect 70802 56284 71000 56342
rect 70802 56238 70824 56284
rect 70870 56238 70928 56284
rect 70974 56238 71000 56284
rect 70802 56180 71000 56238
rect 70802 56134 70824 56180
rect 70870 56134 70928 56180
rect 70974 56134 71000 56180
rect 70802 56076 71000 56134
rect 70802 56030 70824 56076
rect 70870 56030 70928 56076
rect 70974 56030 71000 56076
rect 70802 55972 71000 56030
rect 70802 55926 70824 55972
rect 70870 55926 70928 55972
rect 70974 55926 71000 55972
rect 70802 55868 71000 55926
rect 70802 55822 70824 55868
rect 70870 55822 70928 55868
rect 70974 55822 71000 55868
rect 70802 55764 71000 55822
rect 70802 55718 70824 55764
rect 70870 55718 70928 55764
rect 70974 55718 71000 55764
rect 70802 55660 71000 55718
rect 70802 55614 70824 55660
rect 70870 55614 70928 55660
rect 70974 55614 71000 55660
rect 70802 55556 71000 55614
rect 70802 55510 70824 55556
rect 70870 55510 70928 55556
rect 70974 55510 71000 55556
rect 70802 55452 71000 55510
rect 70802 55406 70824 55452
rect 70870 55406 70928 55452
rect 70974 55406 71000 55452
rect 70802 55348 71000 55406
rect 70802 55302 70824 55348
rect 70870 55302 70928 55348
rect 70974 55302 71000 55348
rect 70802 55244 71000 55302
rect 70802 55198 70824 55244
rect 70870 55198 70928 55244
rect 70974 55198 71000 55244
rect 70802 55140 71000 55198
rect 70802 55094 70824 55140
rect 70870 55094 70928 55140
rect 70974 55094 71000 55140
rect 70802 55036 71000 55094
rect 70802 54990 70824 55036
rect 70870 54990 70928 55036
rect 70974 54990 71000 55036
rect 70802 54932 71000 54990
rect 70802 54886 70824 54932
rect 70870 54886 70928 54932
rect 70974 54886 71000 54932
rect 70802 54828 71000 54886
rect 70802 54782 70824 54828
rect 70870 54782 70928 54828
rect 70974 54782 71000 54828
rect 70802 54724 71000 54782
rect 70802 54678 70824 54724
rect 70870 54678 70928 54724
rect 70974 54678 71000 54724
rect 70802 54620 71000 54678
rect 70802 54574 70824 54620
rect 70870 54574 70928 54620
rect 70974 54574 71000 54620
rect 70802 54516 71000 54574
rect 70802 54470 70824 54516
rect 70870 54470 70928 54516
rect 70974 54470 71000 54516
rect 70802 54412 71000 54470
rect 70802 54366 70824 54412
rect 70870 54366 70928 54412
rect 70974 54366 71000 54412
rect 70802 54308 71000 54366
rect 70802 54262 70824 54308
rect 70870 54262 70928 54308
rect 70974 54262 71000 54308
rect 70802 54204 71000 54262
rect 70802 54158 70824 54204
rect 70870 54158 70928 54204
rect 70974 54158 71000 54204
rect 70802 54100 71000 54158
rect 70802 54054 70824 54100
rect 70870 54054 70928 54100
rect 70974 54054 71000 54100
rect 70802 53996 71000 54054
rect 70802 53950 70824 53996
rect 70870 53950 70928 53996
rect 70974 53950 71000 53996
rect 70802 53892 71000 53950
rect 70802 53846 70824 53892
rect 70870 53846 70928 53892
rect 70974 53846 71000 53892
rect 70802 53788 71000 53846
rect 70802 53742 70824 53788
rect 70870 53742 70928 53788
rect 70974 53742 71000 53788
rect 70802 53684 71000 53742
rect 70802 53638 70824 53684
rect 70870 53638 70928 53684
rect 70974 53638 71000 53684
rect 70802 53580 71000 53638
rect 70802 53534 70824 53580
rect 70870 53534 70928 53580
rect 70974 53534 71000 53580
rect 70802 53476 71000 53534
rect 70802 53430 70824 53476
rect 70870 53430 70928 53476
rect 70974 53430 71000 53476
rect 70802 53372 71000 53430
rect 70802 53326 70824 53372
rect 70870 53326 70928 53372
rect 70974 53326 71000 53372
rect 70802 53268 71000 53326
rect 70802 53222 70824 53268
rect 70870 53222 70928 53268
rect 70974 53222 71000 53268
rect 70802 53164 71000 53222
rect 70802 53118 70824 53164
rect 70870 53118 70928 53164
rect 70974 53118 71000 53164
rect 70802 53060 71000 53118
rect 70802 53014 70824 53060
rect 70870 53014 70928 53060
rect 70974 53014 71000 53060
rect 70802 52956 71000 53014
rect 70802 52910 70824 52956
rect 70870 52910 70928 52956
rect 70974 52910 71000 52956
rect 70802 52852 71000 52910
rect 70802 52806 70824 52852
rect 70870 52806 70928 52852
rect 70974 52806 71000 52852
rect 70802 52748 71000 52806
rect 70802 52702 70824 52748
rect 70870 52702 70928 52748
rect 70974 52702 71000 52748
rect 70802 52644 71000 52702
rect 70802 52598 70824 52644
rect 70870 52598 70928 52644
rect 70974 52598 71000 52644
rect 70802 52540 71000 52598
rect 70802 52494 70824 52540
rect 70870 52494 70928 52540
rect 70974 52494 71000 52540
rect 70802 52436 71000 52494
rect 70802 52390 70824 52436
rect 70870 52390 70928 52436
rect 70974 52390 71000 52436
rect 70802 52332 71000 52390
rect 70802 52286 70824 52332
rect 70870 52286 70928 52332
rect 70974 52286 71000 52332
rect 70802 52228 71000 52286
rect 70802 52182 70824 52228
rect 70870 52182 70928 52228
rect 70974 52182 71000 52228
rect 70802 52124 71000 52182
rect 70802 52078 70824 52124
rect 70870 52078 70928 52124
rect 70974 52078 71000 52124
rect 70802 52020 71000 52078
rect 70802 51974 70824 52020
rect 70870 51974 70928 52020
rect 70974 51974 71000 52020
rect 70802 51916 71000 51974
rect 70802 51870 70824 51916
rect 70870 51870 70928 51916
rect 70974 51870 71000 51916
rect 70802 51812 71000 51870
rect 70802 51766 70824 51812
rect 70870 51766 70928 51812
rect 70974 51766 71000 51812
rect 70802 51708 71000 51766
rect 70802 51662 70824 51708
rect 70870 51662 70928 51708
rect 70974 51662 71000 51708
rect 70802 51604 71000 51662
rect 70802 51558 70824 51604
rect 70870 51558 70928 51604
rect 70974 51558 71000 51604
rect 70802 51500 71000 51558
rect 70802 51454 70824 51500
rect 70870 51454 70928 51500
rect 70974 51454 71000 51500
rect 70802 51396 71000 51454
rect 70802 51350 70824 51396
rect 70870 51350 70928 51396
rect 70974 51350 71000 51396
rect 70802 51292 71000 51350
rect 70802 51246 70824 51292
rect 70870 51246 70928 51292
rect 70974 51246 71000 51292
rect 70802 51188 71000 51246
rect 70802 51142 70824 51188
rect 70870 51142 70928 51188
rect 70974 51142 71000 51188
rect 70802 51084 71000 51142
rect 70802 51038 70824 51084
rect 70870 51038 70928 51084
rect 70974 51038 71000 51084
rect 70802 50980 71000 51038
rect 70802 50934 70824 50980
rect 70870 50934 70928 50980
rect 70974 50934 71000 50980
rect 70802 50876 71000 50934
rect 70802 50830 70824 50876
rect 70870 50830 70928 50876
rect 70974 50830 71000 50876
rect 70802 50772 71000 50830
rect 70802 50726 70824 50772
rect 70870 50726 70928 50772
rect 70974 50726 71000 50772
rect 70802 50668 71000 50726
rect 70802 50622 70824 50668
rect 70870 50622 70928 50668
rect 70974 50622 71000 50668
rect 70802 50564 71000 50622
rect 70802 50518 70824 50564
rect 70870 50518 70928 50564
rect 70974 50518 71000 50564
rect 70802 50460 71000 50518
rect 70802 50414 70824 50460
rect 70870 50414 70928 50460
rect 70974 50414 71000 50460
rect 70802 50356 71000 50414
rect 70802 50310 70824 50356
rect 70870 50310 70928 50356
rect 70974 50310 71000 50356
rect 70802 50252 71000 50310
rect 70802 50206 70824 50252
rect 70870 50206 70928 50252
rect 70974 50206 71000 50252
rect 70802 50148 71000 50206
rect 70802 50102 70824 50148
rect 70870 50102 70928 50148
rect 70974 50102 71000 50148
rect 70802 50044 71000 50102
rect 70802 49998 70824 50044
rect 70870 49998 70928 50044
rect 70974 49998 71000 50044
rect 70802 49940 71000 49998
rect 70802 49894 70824 49940
rect 70870 49894 70928 49940
rect 70974 49894 71000 49940
rect 70802 49836 71000 49894
rect 70802 49790 70824 49836
rect 70870 49790 70928 49836
rect 70974 49790 71000 49836
rect 70802 49732 71000 49790
rect 70802 49686 70824 49732
rect 70870 49686 70928 49732
rect 70974 49686 71000 49732
rect 70802 49628 71000 49686
rect 70802 49582 70824 49628
rect 70870 49582 70928 49628
rect 70974 49582 71000 49628
rect 70802 49524 71000 49582
rect 70802 49478 70824 49524
rect 70870 49478 70928 49524
rect 70974 49478 71000 49524
rect 70802 49420 71000 49478
rect 70802 49374 70824 49420
rect 70870 49374 70928 49420
rect 70974 49374 71000 49420
rect 70802 49316 71000 49374
rect 70802 49270 70824 49316
rect 70870 49270 70928 49316
rect 70974 49270 71000 49316
rect 70802 49212 71000 49270
rect 70802 49166 70824 49212
rect 70870 49166 70928 49212
rect 70974 49166 71000 49212
rect 70802 49108 71000 49166
rect 70802 49062 70824 49108
rect 70870 49062 70928 49108
rect 70974 49062 71000 49108
rect 70802 49004 71000 49062
rect 70802 48958 70824 49004
rect 70870 48958 70928 49004
rect 70974 48958 71000 49004
rect 70802 48900 71000 48958
rect 70802 48854 70824 48900
rect 70870 48854 70928 48900
rect 70974 48854 71000 48900
rect 70802 48796 71000 48854
rect 70802 48750 70824 48796
rect 70870 48750 70928 48796
rect 70974 48750 71000 48796
rect 70802 48692 71000 48750
rect 70802 48646 70824 48692
rect 70870 48646 70928 48692
rect 70974 48646 71000 48692
rect 70802 48588 71000 48646
rect 70802 48542 70824 48588
rect 70870 48542 70928 48588
rect 70974 48542 71000 48588
rect 70802 48484 71000 48542
rect 70802 48438 70824 48484
rect 70870 48438 70928 48484
rect 70974 48438 71000 48484
rect 70802 48380 71000 48438
rect 70802 48334 70824 48380
rect 70870 48334 70928 48380
rect 70974 48334 71000 48380
rect 70802 48276 71000 48334
rect 70802 48230 70824 48276
rect 70870 48230 70928 48276
rect 70974 48230 71000 48276
rect 70802 48172 71000 48230
rect 70802 48126 70824 48172
rect 70870 48126 70928 48172
rect 70974 48126 71000 48172
rect 70802 48068 71000 48126
rect 70802 48022 70824 48068
rect 70870 48022 70928 48068
rect 70974 48022 71000 48068
rect 70802 47964 71000 48022
rect 70802 47918 70824 47964
rect 70870 47918 70928 47964
rect 70974 47918 71000 47964
rect 70802 47860 71000 47918
rect 70802 47814 70824 47860
rect 70870 47814 70928 47860
rect 70974 47814 71000 47860
rect 70802 47756 71000 47814
rect 70802 47710 70824 47756
rect 70870 47710 70928 47756
rect 70974 47710 71000 47756
rect 70802 47652 71000 47710
rect 70802 47606 70824 47652
rect 70870 47606 70928 47652
rect 70974 47606 71000 47652
rect 70802 47548 71000 47606
rect 70802 47502 70824 47548
rect 70870 47502 70928 47548
rect 70974 47502 71000 47548
rect 70802 47444 71000 47502
rect 70802 47398 70824 47444
rect 70870 47398 70928 47444
rect 70974 47398 71000 47444
rect 70802 47340 71000 47398
rect 70802 47294 70824 47340
rect 70870 47294 70928 47340
rect 70974 47294 71000 47340
rect 70802 47236 71000 47294
rect 70802 47190 70824 47236
rect 70870 47190 70928 47236
rect 70974 47190 71000 47236
rect 70802 47132 71000 47190
rect 70802 47086 70824 47132
rect 70870 47086 70928 47132
rect 70974 47086 71000 47132
rect 70802 47028 71000 47086
rect 70802 46982 70824 47028
rect 70870 46982 70928 47028
rect 70974 46982 71000 47028
rect 70802 46924 71000 46982
rect 70802 46878 70824 46924
rect 70870 46878 70928 46924
rect 70974 46878 71000 46924
rect 70802 46820 71000 46878
rect 70802 46774 70824 46820
rect 70870 46774 70928 46820
rect 70974 46774 71000 46820
rect 70802 46716 71000 46774
rect 70802 46670 70824 46716
rect 70870 46670 70928 46716
rect 70974 46670 71000 46716
rect 70802 46612 71000 46670
rect 70802 46566 70824 46612
rect 70870 46566 70928 46612
rect 70974 46566 71000 46612
rect 70802 46508 71000 46566
rect 70802 46462 70824 46508
rect 70870 46462 70928 46508
rect 70974 46462 71000 46508
rect 70802 46404 71000 46462
rect 70802 46358 70824 46404
rect 70870 46358 70928 46404
rect 70974 46358 71000 46404
rect 70802 46300 71000 46358
rect 70802 46254 70824 46300
rect 70870 46254 70928 46300
rect 70974 46254 71000 46300
rect 70802 46196 71000 46254
rect 70802 46150 70824 46196
rect 70870 46150 70928 46196
rect 70974 46150 71000 46196
rect 70802 46092 71000 46150
rect 70802 46046 70824 46092
rect 70870 46046 70928 46092
rect 70974 46046 71000 46092
rect 70802 45988 71000 46046
rect 70802 45942 70824 45988
rect 70870 45942 70928 45988
rect 70974 45942 71000 45988
rect 70802 45884 71000 45942
rect 70802 45838 70824 45884
rect 70870 45838 70928 45884
rect 70974 45838 71000 45884
rect 70802 45780 71000 45838
rect 70802 45734 70824 45780
rect 70870 45734 70928 45780
rect 70974 45734 71000 45780
rect 70802 45676 71000 45734
rect 70802 45630 70824 45676
rect 70870 45630 70928 45676
rect 70974 45630 71000 45676
rect 70802 45572 71000 45630
rect 70802 45526 70824 45572
rect 70870 45526 70928 45572
rect 70974 45526 71000 45572
rect 70802 45468 71000 45526
rect 70802 45422 70824 45468
rect 70870 45422 70928 45468
rect 70974 45422 71000 45468
rect 70802 45364 71000 45422
rect 70802 45318 70824 45364
rect 70870 45318 70928 45364
rect 70974 45318 71000 45364
rect 70802 45260 71000 45318
rect 70802 45214 70824 45260
rect 70870 45214 70928 45260
rect 70974 45214 71000 45260
rect 70802 45156 71000 45214
rect 70802 45110 70824 45156
rect 70870 45110 70928 45156
rect 70974 45110 71000 45156
rect 70802 45052 71000 45110
rect 70802 45006 70824 45052
rect 70870 45006 70928 45052
rect 70974 45006 71000 45052
rect 70802 44948 71000 45006
tri 13291 44892 13323 44924 sw
rect 70802 44902 70824 44948
rect 70870 44902 70928 44948
rect 70974 44902 71000 44948
rect 13097 44878 13323 44892
tri 13323 44878 13337 44892 sw
rect 13097 44847 13337 44878
tri 13337 44847 13368 44878 sw
rect 13097 44846 13368 44847
tri 13368 44846 13369 44847 sw
rect 13097 44844 13369 44846
tri 13097 44831 13110 44844 ne
rect 13110 44833 13369 44844
tri 13369 44833 13382 44846 sw
rect 70802 44844 71000 44902
rect 13110 44831 13382 44833
tri 13110 44785 13155 44831 ne
rect 13155 44824 13382 44831
rect 13155 44785 13254 44824
tri 13155 44769 13172 44785 ne
rect 13172 44778 13254 44785
rect 13300 44801 13382 44824
tri 13382 44801 13414 44833 sw
rect 13300 44778 13414 44801
rect 13172 44769 13414 44778
tri 13172 44756 13185 44769 ne
rect 13185 44756 13414 44769
tri 13414 44756 13459 44801 sw
rect 70802 44798 70824 44844
rect 70870 44798 70928 44844
rect 70974 44798 71000 44844
tri 13185 44724 13217 44756 ne
rect 13217 44746 13459 44756
tri 13459 44746 13469 44756 sw
rect 13217 44724 13469 44746
tri 13217 44714 13227 44724 ne
rect 13227 44714 13469 44724
tri 13469 44714 13501 44746 sw
rect 70802 44740 71000 44798
tri 13227 44696 13245 44714 ne
rect 13245 44701 13501 44714
tri 13501 44701 13514 44714 sw
rect 13245 44696 13514 44701
tri 13514 44696 13519 44701 sw
tri 13245 44651 13290 44696 ne
rect 13290 44692 13519 44696
rect 13290 44651 13386 44692
tri 13290 44637 13304 44651 ne
rect 13304 44646 13386 44651
rect 13432 44651 13519 44692
tri 13519 44651 13565 44696 sw
rect 70802 44694 70824 44740
rect 70870 44694 70928 44740
rect 70974 44694 71000 44740
rect 13432 44646 13565 44651
rect 13304 44637 13565 44646
tri 13304 44624 13317 44637 ne
rect 13317 44624 13565 44637
tri 13565 44624 13591 44651 sw
rect 70802 44636 71000 44694
tri 13317 44592 13349 44624 ne
rect 13349 44614 13591 44624
tri 13591 44614 13601 44624 sw
rect 13349 44592 13601 44614
tri 13349 44573 13368 44592 ne
rect 13368 44582 13601 44592
tri 13601 44582 13633 44614 sw
rect 70802 44590 70824 44636
rect 70870 44590 70928 44636
rect 70974 44590 71000 44636
rect 13368 44573 13633 44582
tri 13633 44573 13643 44582 sw
tri 13368 44527 13413 44573 ne
rect 13413 44569 13643 44573
tri 13643 44569 13646 44573 sw
rect 13413 44560 13646 44569
rect 13413 44527 13518 44560
tri 13413 44505 13436 44527 ne
rect 13436 44514 13518 44527
rect 13564 44537 13646 44560
tri 13646 44537 13678 44569 sw
rect 13564 44514 13678 44537
rect 13436 44505 13678 44514
tri 13436 44492 13449 44505 ne
rect 13449 44492 13678 44505
tri 13678 44492 13723 44537 sw
rect 70802 44532 71000 44590
tri 13449 44460 13481 44492 ne
rect 13481 44482 13723 44492
tri 13723 44482 13733 44492 sw
rect 70802 44486 70824 44532
rect 70870 44486 70928 44532
rect 70974 44486 71000 44532
rect 13481 44460 13733 44482
tri 13481 44450 13491 44460 ne
rect 13491 44450 13733 44460
tri 13733 44450 13765 44482 sw
tri 13491 44405 13536 44450 ne
rect 13536 44437 13765 44450
tri 13765 44437 13778 44450 sw
rect 13536 44428 13778 44437
rect 13536 44405 13650 44428
tri 13536 44376 13565 44405 ne
rect 13565 44382 13650 44405
rect 13696 44405 13778 44428
tri 13778 44405 13810 44437 sw
rect 70802 44428 71000 44486
rect 13696 44382 13810 44405
rect 13565 44376 13810 44382
tri 13565 44360 13581 44376 ne
rect 13581 44360 13810 44376
tri 13810 44360 13855 44405 sw
rect 70802 44382 70824 44428
rect 70870 44382 70928 44428
rect 70974 44382 71000 44428
tri 13581 44328 13613 44360 ne
rect 13613 44350 13855 44360
tri 13855 44350 13865 44360 sw
rect 13613 44328 13865 44350
tri 13613 44298 13643 44328 ne
rect 13643 44318 13865 44328
tri 13865 44318 13897 44350 sw
rect 70802 44324 71000 44382
rect 13643 44298 13897 44318
tri 13897 44298 13917 44318 sw
tri 13643 44253 13688 44298 ne
rect 13688 44296 13917 44298
rect 13688 44253 13782 44296
tri 13688 44241 13700 44253 ne
rect 13700 44250 13782 44253
rect 13828 44286 13917 44296
tri 13917 44286 13929 44298 sw
rect 13828 44273 13929 44286
tri 13929 44273 13942 44286 sw
rect 70802 44278 70824 44324
rect 70870 44278 70928 44324
rect 70974 44278 71000 44324
rect 13828 44250 13942 44273
rect 13700 44241 13942 44250
tri 13700 44228 13713 44241 ne
rect 13713 44228 13942 44241
tri 13942 44228 13987 44273 sw
tri 13713 44196 13745 44228 ne
rect 13745 44218 13987 44228
tri 13987 44218 13997 44228 sw
rect 70802 44220 71000 44278
rect 13745 44196 13997 44218
tri 13745 44186 13755 44196 ne
rect 13755 44186 13997 44196
tri 13997 44186 14029 44218 sw
tri 13755 44141 13800 44186 ne
rect 13800 44173 14029 44186
tri 14029 44173 14042 44186 sw
rect 70802 44174 70824 44220
rect 70870 44174 70928 44220
rect 70974 44174 71000 44220
rect 13800 44164 14042 44173
rect 13800 44141 13914 44164
tri 13800 44109 13832 44141 ne
rect 13832 44118 13914 44141
rect 13960 44141 14042 44164
tri 14042 44141 14074 44173 sw
rect 13960 44118 14074 44141
rect 13832 44109 14074 44118
tri 13832 44096 13845 44109 ne
rect 13845 44096 14074 44109
tri 14074 44096 14119 44141 sw
rect 70802 44116 71000 44174
tri 13845 44064 13877 44096 ne
rect 13877 44086 14119 44096
tri 14119 44086 14129 44096 sw
rect 13877 44064 14129 44086
tri 13877 44024 13917 44064 ne
rect 13917 44054 14129 44064
tri 14129 44054 14161 44086 sw
rect 70802 44070 70824 44116
rect 70870 44070 70928 44116
rect 70974 44070 71000 44116
rect 13917 44041 14161 44054
tri 14161 44041 14174 44054 sw
rect 13917 44032 14174 44041
rect 13917 44024 14046 44032
tri 13917 44011 13929 44024 ne
rect 13929 44011 14046 44024
tri 13929 43966 13975 44011 ne
rect 13975 43986 14046 44011
rect 14092 44024 14174 44032
tri 14174 44024 14191 44041 sw
rect 14092 44011 14191 44024
tri 14191 44011 14204 44024 sw
rect 70802 44012 71000 44070
rect 14092 43986 14204 44011
rect 13975 43966 14204 43986
tri 14204 43966 14249 44011 sw
rect 70802 43966 70824 44012
rect 70870 43966 70928 44012
rect 70974 43966 71000 44012
tri 13975 43964 13977 43966 ne
rect 13977 43964 14249 43966
tri 14249 43964 14251 43966 sw
tri 13977 43932 14009 43964 ne
rect 14009 43932 14251 43964
tri 14009 43922 14019 43932 ne
rect 14019 43922 14251 43932
tri 14251 43922 14293 43964 sw
tri 14019 43877 14064 43922 ne
rect 14064 43909 14293 43922
tri 14293 43909 14306 43922 sw
rect 14064 43900 14306 43909
rect 14064 43877 14178 43900
tri 14064 43845 14096 43877 ne
rect 14096 43854 14178 43877
rect 14224 43877 14306 43900
tri 14306 43877 14338 43909 sw
rect 70802 43908 71000 43966
rect 14224 43854 14338 43877
rect 14096 43845 14338 43854
tri 14096 43832 14109 43845 ne
rect 14109 43832 14338 43845
tri 14338 43832 14383 43877 sw
rect 70802 43862 70824 43908
rect 70870 43862 70928 43908
rect 70974 43862 71000 43908
tri 14109 43800 14141 43832 ne
rect 14141 43822 14383 43832
tri 14383 43822 14393 43832 sw
rect 14141 43800 14393 43822
tri 14141 43755 14186 43800 ne
rect 14186 43790 14393 43800
tri 14393 43790 14425 43822 sw
rect 70802 43804 71000 43862
rect 14186 43777 14425 43790
tri 14425 43777 14438 43790 sw
rect 14186 43768 14438 43777
rect 14186 43755 14310 43768
tri 14186 43749 14191 43755 ne
rect 14191 43749 14310 43755
tri 14191 43713 14228 43749 ne
rect 14228 43722 14310 43749
rect 14356 43749 14438 43768
tri 14438 43749 14466 43777 sw
rect 70802 43758 70824 43804
rect 70870 43758 70928 43804
rect 70974 43758 71000 43804
rect 14356 43745 14466 43749
tri 14466 43745 14470 43749 sw
rect 14356 43722 14470 43745
rect 14228 43713 14470 43722
tri 14228 43700 14241 43713 ne
rect 14241 43700 14470 43713
tri 14470 43700 14515 43745 sw
rect 70802 43700 71000 43758
tri 14241 43668 14273 43700 ne
rect 14273 43690 14515 43700
tri 14515 43690 14525 43700 sw
rect 14273 43668 14525 43690
tri 14273 43658 14283 43668 ne
rect 14283 43658 14525 43668
tri 14525 43658 14557 43690 sw
tri 14283 43647 14294 43658 ne
rect 14294 43647 14557 43658
tri 14294 43601 14339 43647 ne
rect 14339 43645 14557 43647
tri 14557 43645 14570 43658 sw
rect 70802 43654 70824 43700
rect 70870 43654 70928 43700
rect 70974 43654 71000 43700
rect 14339 43636 14570 43645
rect 14339 43601 14442 43636
tri 14339 43581 14360 43601 ne
rect 14360 43590 14442 43601
rect 14488 43601 14570 43636
tri 14570 43601 14614 43645 sw
rect 14488 43590 14614 43601
rect 14360 43581 14614 43590
tri 14360 43568 14373 43581 ne
rect 14373 43568 14614 43581
tri 14614 43568 14647 43601 sw
rect 70802 43596 71000 43654
tri 14373 43536 14405 43568 ne
rect 14405 43558 14647 43568
tri 14647 43558 14657 43568 sw
rect 14405 43536 14657 43558
tri 14405 43491 14450 43536 ne
rect 14450 43526 14657 43536
tri 14657 43526 14689 43558 sw
rect 70802 43550 70824 43596
rect 70870 43550 70928 43596
rect 70974 43550 71000 43596
rect 14450 43513 14689 43526
tri 14689 43513 14702 43526 sw
rect 14450 43504 14702 43513
rect 14450 43491 14574 43504
tri 14450 43475 14466 43491 ne
rect 14466 43475 14574 43491
tri 14466 43449 14492 43475 ne
rect 14492 43458 14574 43475
rect 14620 43475 14702 43504
tri 14702 43475 14740 43513 sw
rect 70802 43492 71000 43550
rect 14620 43458 14740 43475
rect 14492 43449 14740 43458
tri 14492 43436 14505 43449 ne
rect 14505 43436 14740 43449
tri 14740 43436 14779 43475 sw
rect 70802 43446 70824 43492
rect 70870 43446 70928 43492
rect 70974 43446 71000 43492
tri 14505 43404 14537 43436 ne
rect 14537 43426 14779 43436
tri 14779 43426 14789 43436 sw
rect 14537 43404 14789 43426
tri 14537 43394 14547 43404 ne
rect 14547 43394 14789 43404
tri 14789 43394 14821 43426 sw
tri 14547 43349 14592 43394 ne
rect 14592 43381 14821 43394
tri 14821 43381 14834 43394 sw
rect 70802 43388 71000 43446
rect 14592 43372 14834 43381
rect 14592 43349 14706 43372
tri 14592 43317 14624 43349 ne
rect 14624 43326 14706 43349
rect 14752 43349 14834 43372
tri 14834 43349 14866 43381 sw
rect 14752 43326 14866 43349
rect 14624 43317 14866 43326
tri 14624 43304 14637 43317 ne
rect 14637 43304 14866 43317
tri 14866 43304 14911 43349 sw
rect 70802 43342 70824 43388
rect 70870 43342 70928 43388
rect 70974 43342 71000 43388
tri 14637 43272 14669 43304 ne
rect 14669 43294 14911 43304
tri 14911 43294 14921 43304 sw
rect 14669 43272 14921 43294
tri 14669 43237 14704 43272 ne
rect 14704 43262 14921 43272
tri 14921 43262 14953 43294 sw
rect 70802 43284 71000 43342
rect 14704 43249 14953 43262
tri 14953 43249 14966 43262 sw
rect 14704 43240 14966 43249
rect 14704 43237 14838 43240
tri 14704 43201 14740 43237 ne
rect 14740 43201 14838 43237
tri 14740 43185 14756 43201 ne
rect 14756 43194 14838 43201
rect 14884 43237 14966 43240
tri 14966 43237 14979 43249 sw
rect 70802 43238 70824 43284
rect 70870 43238 70928 43284
rect 70974 43238 71000 43284
rect 14884 43201 14979 43237
tri 14979 43201 15015 43237 sw
rect 14884 43194 15015 43201
rect 14756 43191 15015 43194
tri 15015 43191 15024 43201 sw
rect 14756 43185 15024 43191
tri 14756 43172 14769 43185 ne
rect 14769 43172 15024 43185
tri 15024 43172 15043 43191 sw
rect 70802 43180 71000 43238
tri 14769 43140 14801 43172 ne
rect 14801 43162 15043 43172
tri 15043 43162 15053 43172 sw
rect 14801 43140 15053 43162
tri 14801 43130 14811 43140 ne
rect 14811 43130 15053 43140
tri 15053 43130 15085 43162 sw
rect 70802 43134 70824 43180
rect 70870 43134 70928 43180
rect 70974 43134 71000 43180
tri 14811 43085 14856 43130 ne
rect 14856 43117 15085 43130
tri 15085 43117 15098 43130 sw
rect 14856 43108 15098 43117
rect 14856 43085 14970 43108
tri 14856 43053 14888 43085 ne
rect 14888 43062 14970 43085
rect 15016 43085 15098 43108
tri 15098 43085 15130 43117 sw
rect 15016 43062 15130 43085
rect 14888 43053 15130 43062
tri 14888 43040 14901 43053 ne
rect 14901 43040 15130 43053
tri 15130 43040 15175 43085 sw
rect 70802 43076 71000 43134
tri 14901 43008 14933 43040 ne
rect 14933 43030 15175 43040
tri 15175 43030 15185 43040 sw
rect 70802 43030 70824 43076
rect 70870 43030 70928 43076
rect 70974 43030 71000 43076
rect 14933 43008 15185 43030
tri 14933 42963 14978 43008 ne
rect 14978 42998 15185 43008
tri 15185 42998 15217 43030 sw
rect 14978 42985 15217 42998
tri 15217 42985 15230 42998 sw
rect 14978 42976 15230 42985
rect 14978 42963 15102 42976
tri 14978 42926 15015 42963 ne
rect 15015 42930 15102 42963
rect 15148 42971 15230 42976
tri 15230 42971 15244 42985 sw
rect 70802 42972 71000 43030
rect 15148 42930 15244 42971
rect 15015 42926 15244 42930
tri 15244 42926 15289 42971 sw
rect 70802 42926 70824 42972
rect 70870 42926 70928 42972
rect 70974 42926 71000 42972
tri 15015 42917 15024 42926 ne
rect 15024 42917 15289 42926
tri 15024 42908 15033 42917 ne
rect 15033 42908 15289 42917
tri 15289 42908 15307 42926 sw
tri 15033 42872 15069 42908 ne
rect 15069 42898 15307 42908
tri 15307 42898 15317 42908 sw
rect 15069 42872 15317 42898
tri 15069 42866 15075 42872 ne
rect 15075 42866 15317 42872
tri 15317 42866 15349 42898 sw
rect 70802 42868 71000 42926
tri 15075 42821 15120 42866 ne
rect 15120 42844 15349 42866
rect 15120 42821 15234 42844
tri 15120 42789 15152 42821 ne
rect 15152 42798 15234 42821
rect 15280 42827 15349 42844
tri 15349 42827 15389 42866 sw
rect 15280 42821 15389 42827
tri 15389 42821 15394 42827 sw
rect 70802 42822 70824 42868
rect 70870 42822 70928 42868
rect 70974 42822 71000 42868
rect 15280 42798 15394 42821
rect 15152 42789 15394 42798
tri 15152 42776 15165 42789 ne
rect 15165 42776 15394 42789
tri 15394 42776 15439 42821 sw
tri 15165 42744 15197 42776 ne
rect 15197 42766 15439 42776
tri 15439 42766 15449 42776 sw
rect 15197 42744 15449 42766
tri 15197 42699 15242 42744 ne
rect 15242 42734 15449 42744
tri 15449 42734 15481 42766 sw
rect 70802 42764 71000 42822
rect 15242 42721 15481 42734
tri 15481 42721 15494 42734 sw
rect 15242 42712 15494 42721
rect 15242 42699 15366 42712
tri 15242 42657 15284 42699 ne
rect 15284 42666 15366 42699
rect 15412 42697 15494 42712
tri 15494 42697 15518 42721 sw
rect 70802 42718 70824 42764
rect 70870 42718 70928 42764
rect 70974 42718 71000 42764
rect 15412 42666 15518 42697
rect 15284 42657 15518 42666
tri 15284 42652 15289 42657 ne
rect 15289 42652 15518 42657
tri 15518 42652 15563 42697 sw
rect 70802 42660 71000 42718
tri 15289 42644 15297 42652 ne
rect 15297 42644 15563 42652
tri 15563 42644 15571 42652 sw
tri 15297 42612 15329 42644 ne
rect 15329 42634 15571 42644
tri 15571 42634 15581 42644 sw
rect 15329 42612 15581 42634
tri 15329 42602 15339 42612 ne
rect 15339 42602 15581 42612
tri 15581 42602 15613 42634 sw
rect 70802 42614 70824 42660
rect 70870 42614 70928 42660
rect 70974 42614 71000 42660
tri 15339 42557 15384 42602 ne
rect 15384 42589 15613 42602
tri 15613 42589 15626 42602 sw
rect 15384 42580 15626 42589
rect 15384 42557 15498 42580
tri 15384 42552 15389 42557 ne
rect 15389 42552 15498 42557
tri 15389 42512 15429 42552 ne
rect 15429 42534 15498 42552
rect 15544 42557 15626 42580
tri 15626 42557 15658 42589 sw
rect 15544 42534 15658 42557
rect 15429 42512 15658 42534
tri 15658 42512 15703 42557 sw
rect 70802 42556 71000 42614
tri 15429 42480 15461 42512 ne
rect 15461 42507 15703 42512
tri 15703 42507 15708 42512 sw
rect 70802 42510 70824 42556
rect 70870 42510 70928 42556
rect 70974 42510 71000 42556
rect 15461 42480 15708 42507
tri 15461 42435 15506 42480 ne
rect 15506 42470 15708 42480
tri 15708 42470 15745 42507 sw
rect 15506 42457 15745 42470
tri 15745 42457 15758 42470 sw
rect 15506 42448 15758 42457
rect 15506 42435 15630 42448
tri 15506 42393 15548 42435 ne
rect 15548 42402 15630 42435
rect 15676 42425 15758 42448
tri 15758 42425 15790 42457 sw
rect 70802 42452 71000 42510
rect 15676 42402 15790 42425
rect 15548 42393 15790 42402
tri 15548 42377 15563 42393 ne
rect 15563 42380 15790 42393
tri 15790 42380 15835 42425 sw
rect 70802 42406 70824 42452
rect 70870 42406 70928 42452
rect 70974 42406 71000 42452
rect 15563 42377 15835 42380
tri 15835 42377 15838 42380 sw
tri 15563 42348 15593 42377 ne
rect 15593 42370 15838 42377
tri 15838 42370 15845 42377 sw
rect 15593 42348 15845 42370
tri 15593 42338 15603 42348 ne
rect 15603 42338 15845 42348
tri 15845 42338 15877 42370 sw
rect 70802 42348 71000 42406
tri 15603 42293 15648 42338 ne
rect 15648 42325 15877 42338
tri 15877 42325 15890 42338 sw
rect 15648 42316 15890 42325
rect 15648 42293 15762 42316
tri 15648 42261 15680 42293 ne
rect 15680 42270 15762 42293
rect 15808 42293 15890 42316
tri 15890 42293 15922 42325 sw
rect 70802 42302 70824 42348
rect 70870 42302 70928 42348
rect 70974 42302 71000 42348
rect 15808 42270 15922 42293
rect 15680 42261 15922 42270
tri 15680 42248 15693 42261 ne
rect 15693 42248 15922 42261
tri 15922 42248 15967 42293 sw
tri 15693 42216 15725 42248 ne
rect 15725 42238 15967 42248
tri 15967 42238 15977 42248 sw
rect 70802 42244 71000 42302
rect 15725 42216 15977 42238
tri 15725 42187 15753 42216 ne
rect 15753 42206 15977 42216
tri 15977 42206 16009 42238 sw
rect 15753 42193 16009 42206
tri 16009 42193 16022 42206 sw
rect 70802 42198 70824 42244
rect 70870 42198 70928 42244
rect 70974 42198 71000 42244
rect 15753 42187 16022 42193
tri 16022 42187 16028 42193 sw
tri 15753 42142 15799 42187 ne
rect 15799 42184 16028 42187
rect 15799 42142 15894 42184
tri 15799 42129 15812 42142 ne
rect 15812 42138 15894 42142
rect 15940 42142 16028 42184
tri 16028 42142 16073 42187 sw
rect 15940 42138 16073 42142
rect 15812 42129 16073 42138
tri 15812 42103 15838 42129 ne
rect 15838 42116 16073 42129
tri 16073 42116 16099 42142 sw
rect 70802 42140 71000 42198
rect 15838 42103 16099 42116
tri 16099 42103 16112 42116 sw
tri 15838 42084 15857 42103 ne
rect 15857 42084 16112 42103
tri 15857 42074 15867 42084 ne
rect 15867 42074 16112 42084
tri 16112 42074 16141 42103 sw
rect 70802 42094 70824 42140
rect 70870 42094 70928 42140
rect 70974 42094 71000 42140
tri 15867 42029 15912 42074 ne
rect 15912 42061 16141 42074
tri 16141 42061 16154 42074 sw
rect 15912 42052 16154 42061
rect 15912 42029 16026 42052
tri 15912 41997 15944 42029 ne
rect 15944 42006 16026 42029
rect 16072 42029 16154 42052
tri 16154 42029 16186 42061 sw
rect 70802 42036 71000 42094
rect 16072 42006 16186 42029
rect 15944 41997 16186 42006
tri 15944 41984 15957 41997 ne
rect 15957 41984 16186 41997
tri 16186 41984 16231 42029 sw
rect 70802 41990 70824 42036
rect 70870 41990 70928 42036
rect 70974 41990 71000 42036
tri 15957 41952 15989 41984 ne
rect 15989 41974 16231 41984
tri 16231 41974 16241 41984 sw
rect 15989 41952 16241 41974
tri 15989 41907 16034 41952 ne
rect 16034 41942 16241 41952
tri 16241 41942 16273 41974 sw
rect 16034 41929 16273 41942
tri 16273 41929 16286 41942 sw
rect 70802 41932 71000 41990
rect 16034 41920 16286 41929
rect 16034 41907 16158 41920
tri 16034 41865 16076 41907 ne
rect 16076 41874 16158 41907
rect 16204 41897 16286 41920
tri 16286 41897 16318 41929 sw
rect 16204 41874 16318 41897
rect 16076 41865 16318 41874
tri 16076 41829 16112 41865 ne
rect 16112 41852 16318 41865
tri 16318 41852 16363 41897 sw
rect 70802 41886 70824 41932
rect 70870 41886 70928 41932
rect 70974 41886 71000 41932
rect 16112 41842 16363 41852
tri 16363 41842 16373 41852 sw
rect 16112 41829 16373 41842
tri 16373 41829 16387 41842 sw
tri 16112 41820 16121 41829 ne
rect 16121 41820 16387 41829
tri 16121 41810 16131 41820 ne
rect 16131 41810 16387 41820
tri 16387 41810 16405 41829 sw
rect 70802 41828 71000 41886
tri 16131 41777 16163 41810 ne
rect 16163 41797 16405 41810
tri 16405 41797 16418 41810 sw
rect 16163 41788 16418 41797
rect 16163 41777 16290 41788
tri 16163 41733 16208 41777 ne
rect 16208 41742 16290 41777
rect 16336 41777 16418 41788
tri 16418 41777 16438 41797 sw
rect 70802 41782 70824 41828
rect 70870 41782 70928 41828
rect 70974 41782 71000 41828
rect 16336 41742 16438 41777
rect 16208 41733 16438 41742
tri 16208 41720 16221 41733 ne
rect 16221 41732 16438 41733
tri 16438 41732 16483 41777 sw
rect 16221 41720 16483 41732
tri 16483 41720 16495 41732 sw
rect 70802 41724 71000 41782
tri 16221 41688 16253 41720 ne
rect 16253 41710 16495 41720
tri 16495 41710 16505 41720 sw
rect 16253 41688 16505 41710
tri 16253 41643 16298 41688 ne
rect 16298 41678 16505 41688
tri 16505 41678 16537 41710 sw
rect 70802 41678 70824 41724
rect 70870 41678 70928 41724
rect 70974 41678 71000 41724
rect 16298 41665 16537 41678
tri 16537 41665 16550 41678 sw
rect 16298 41656 16550 41665
rect 16298 41643 16422 41656
tri 16298 41601 16340 41643 ne
rect 16340 41610 16422 41643
rect 16468 41633 16550 41656
tri 16550 41633 16582 41665 sw
rect 16468 41610 16582 41633
rect 16340 41601 16582 41610
tri 16340 41556 16385 41601 ne
rect 16385 41588 16582 41601
tri 16582 41588 16627 41633 sw
rect 70802 41620 71000 41678
rect 16385 41578 16627 41588
tri 16627 41578 16637 41588 sw
rect 16385 41556 16637 41578
tri 16385 41554 16387 41556 ne
rect 16387 41554 16637 41556
tri 16637 41554 16661 41578 sw
rect 70802 41574 70824 41620
rect 70870 41574 70928 41620
rect 70974 41574 71000 41620
tri 16387 41546 16395 41554 ne
rect 16395 41546 16661 41554
tri 16661 41546 16669 41554 sw
tri 16395 41501 16440 41546 ne
rect 16440 41533 16669 41546
tri 16669 41533 16682 41546 sw
rect 16440 41524 16682 41533
rect 16440 41501 16554 41524
tri 16440 41458 16483 41501 ne
rect 16483 41478 16554 41501
rect 16600 41501 16682 41524
tri 16682 41501 16714 41533 sw
rect 70802 41516 71000 41574
rect 16600 41478 16714 41501
rect 16483 41458 16714 41478
tri 16483 41456 16485 41458 ne
rect 16485 41456 16714 41458
tri 16714 41456 16759 41501 sw
rect 70802 41470 70824 41516
rect 70870 41470 70928 41516
rect 70974 41470 71000 41516
tri 16485 41413 16528 41456 ne
rect 16528 41446 16759 41456
tri 16759 41446 16769 41456 sw
rect 16528 41414 16769 41446
tri 16769 41414 16801 41446 sw
rect 16528 41413 16801 41414
tri 16801 41413 16803 41414 sw
tri 16528 41367 16573 41413 ne
rect 16573 41392 16803 41413
rect 16573 41367 16686 41392
tri 16573 41337 16604 41367 ne
rect 16604 41346 16686 41367
rect 16732 41367 16803 41392
tri 16803 41367 16848 41413 sw
rect 70802 41412 71000 41470
rect 16732 41346 16848 41367
rect 16604 41337 16848 41346
tri 16604 41292 16649 41337 ne
rect 16649 41324 16848 41337
tri 16848 41324 16891 41367 sw
rect 70802 41366 70824 41412
rect 70870 41366 70928 41412
rect 70974 41366 71000 41412
rect 16649 41314 16891 41324
tri 16891 41314 16901 41324 sw
rect 16649 41292 16901 41314
tri 16649 41280 16661 41292 ne
rect 16661 41282 16901 41292
tri 16901 41282 16933 41314 sw
rect 70802 41308 71000 41366
rect 16661 41280 16933 41282
tri 16933 41280 16935 41282 sw
tri 16661 41235 16706 41280 ne
rect 16706 41269 16935 41280
tri 16935 41269 16946 41280 sw
rect 16706 41260 16946 41269
rect 16706 41235 16818 41260
tri 16706 41205 16736 41235 ne
rect 16736 41214 16818 41235
rect 16864 41237 16946 41260
tri 16946 41237 16978 41269 sw
rect 70802 41262 70824 41308
rect 70870 41262 70928 41308
rect 70974 41262 71000 41308
rect 16864 41214 16978 41237
rect 16736 41205 16978 41214
tri 16736 41192 16749 41205 ne
rect 16749 41192 16978 41205
tri 16978 41192 17023 41237 sw
rect 70802 41204 71000 41262
tri 16749 41160 16781 41192 ne
rect 16781 41182 17023 41192
tri 17023 41182 17033 41192 sw
rect 16781 41160 17033 41182
tri 16781 41150 16791 41160 ne
rect 16791 41150 17033 41160
tri 17033 41150 17065 41182 sw
rect 70802 41158 70824 41204
rect 70870 41158 70928 41204
rect 70974 41158 71000 41204
tri 16791 41105 16836 41150 ne
rect 16836 41137 17065 41150
tri 17065 41137 17078 41150 sw
rect 16836 41128 17078 41137
rect 16836 41105 16950 41128
tri 16836 41093 16848 41105 ne
rect 16848 41093 16950 41105
tri 16848 41060 16881 41093 ne
rect 16881 41082 16950 41093
rect 16996 41105 17078 41128
tri 17078 41105 17110 41137 sw
rect 16996 41082 17110 41105
rect 16881 41060 17110 41082
tri 17110 41060 17155 41105 sw
rect 70802 41100 71000 41158
tri 16881 41028 16913 41060 ne
rect 16913 41050 17155 41060
tri 17155 41050 17165 41060 sw
rect 70802 41054 70824 41100
rect 70870 41054 70928 41100
rect 70974 41054 71000 41100
rect 16913 41028 17165 41050
tri 16913 41005 16935 41028 ne
rect 16935 41018 17165 41028
tri 17165 41018 17197 41050 sw
rect 16935 41005 17197 41018
tri 17197 41005 17210 41018 sw
tri 16935 40960 16981 41005 ne
rect 16981 41003 17210 41005
tri 17210 41003 17213 41005 sw
rect 16981 40996 17213 41003
rect 16981 40960 17082 40996
tri 16981 40941 17000 40960 ne
rect 17000 40950 17082 40960
rect 17128 40973 17213 40996
tri 17213 40973 17242 41003 sw
rect 70802 40996 71000 41054
rect 17128 40950 17242 40973
rect 17000 40941 17242 40950
tri 17000 40928 17013 40941 ne
rect 17013 40928 17242 40941
tri 17242 40928 17287 40973 sw
rect 70802 40950 70824 40996
rect 70870 40950 70928 40996
rect 70974 40950 71000 40996
tri 17013 40896 17045 40928 ne
rect 17045 40918 17287 40928
tri 17287 40918 17297 40928 sw
rect 17045 40896 17297 40918
tri 17045 40886 17055 40896 ne
rect 17055 40886 17297 40896
tri 17297 40886 17329 40918 sw
rect 70802 40892 71000 40950
tri 17055 40841 17100 40886 ne
rect 17100 40873 17329 40886
tri 17329 40873 17342 40886 sw
rect 17100 40864 17342 40873
rect 17100 40841 17214 40864
tri 17100 40809 17132 40841 ne
rect 17132 40818 17214 40841
rect 17260 40841 17342 40864
tri 17342 40841 17374 40873 sw
rect 70802 40846 70824 40892
rect 70870 40846 70928 40892
rect 70974 40846 71000 40892
rect 17260 40818 17374 40841
rect 17132 40809 17374 40818
tri 17132 40796 17145 40809 ne
rect 17145 40796 17374 40809
tri 17374 40796 17419 40841 sw
tri 17145 40764 17177 40796 ne
rect 17177 40786 17419 40796
tri 17419 40786 17429 40796 sw
rect 70802 40788 71000 40846
rect 17177 40764 17429 40786
tri 17177 40731 17210 40764 ne
rect 17210 40754 17429 40764
tri 17429 40754 17461 40786 sw
rect 17210 40741 17461 40754
tri 17461 40741 17474 40754 sw
rect 70802 40742 70824 40788
rect 70870 40742 70928 40788
rect 70974 40742 71000 40788
rect 17210 40732 17474 40741
rect 17210 40731 17346 40732
tri 17210 40728 17213 40731 ne
rect 17213 40728 17346 40731
tri 17213 40683 17258 40728 ne
rect 17258 40686 17346 40728
rect 17392 40731 17474 40732
tri 17474 40731 17484 40741 sw
rect 17392 40728 17484 40731
tri 17484 40728 17487 40731 sw
rect 17392 40686 17487 40728
rect 17258 40683 17487 40686
tri 17487 40683 17532 40728 sw
rect 70802 40684 71000 40742
tri 17258 40677 17264 40683 ne
rect 17264 40677 17532 40683
tri 17264 40664 17277 40677 ne
rect 17277 40664 17532 40677
tri 17532 40664 17551 40683 sw
tri 17277 40632 17309 40664 ne
rect 17309 40654 17551 40664
tri 17551 40654 17561 40664 sw
rect 17309 40632 17561 40654
tri 17309 40622 17319 40632 ne
rect 17319 40622 17561 40632
tri 17561 40622 17593 40654 sw
rect 70802 40638 70824 40684
rect 70870 40638 70928 40684
rect 70974 40638 71000 40684
tri 17319 40577 17364 40622 ne
rect 17364 40609 17593 40622
tri 17593 40609 17606 40622 sw
rect 17364 40600 17606 40609
rect 17364 40577 17478 40600
tri 17364 40545 17396 40577 ne
rect 17396 40554 17478 40577
rect 17524 40577 17606 40600
tri 17606 40577 17638 40609 sw
rect 70802 40580 71000 40638
rect 17524 40554 17638 40577
rect 17396 40545 17638 40554
tri 17396 40532 17409 40545 ne
rect 17409 40532 17638 40545
tri 17638 40532 17683 40577 sw
rect 70802 40534 70824 40580
rect 70870 40534 70928 40580
rect 70974 40534 71000 40580
tri 17409 40500 17441 40532 ne
rect 17441 40522 17683 40532
tri 17683 40522 17693 40532 sw
rect 17441 40500 17693 40522
tri 17441 40457 17484 40500 ne
rect 17484 40490 17693 40500
tri 17693 40490 17725 40522 sw
rect 17484 40477 17725 40490
tri 17725 40477 17738 40490 sw
rect 17484 40468 17738 40477
rect 17484 40457 17610 40468
tri 17484 40413 17528 40457 ne
rect 17528 40422 17610 40457
rect 17656 40457 17738 40468
tri 17738 40457 17759 40477 sw
rect 70802 40476 71000 40534
rect 17656 40445 17759 40457
tri 17759 40445 17770 40457 sw
rect 17656 40422 17770 40445
rect 17528 40413 17770 40422
tri 17528 40400 17541 40413 ne
rect 17541 40400 17770 40413
tri 17770 40400 17815 40445 sw
rect 70802 40430 70824 40476
rect 70870 40430 70928 40476
rect 70974 40430 71000 40476
tri 17541 40368 17573 40400 ne
rect 17573 40390 17815 40400
tri 17815 40390 17825 40400 sw
rect 17573 40368 17825 40390
tri 17573 40363 17577 40368 ne
rect 17577 40363 17825 40368
tri 17577 40358 17583 40363 ne
rect 17583 40358 17825 40363
tri 17825 40358 17857 40390 sw
rect 70802 40372 71000 40430
tri 17583 40318 17623 40358 ne
rect 17623 40345 17857 40358
tri 17857 40345 17870 40358 sw
rect 17623 40336 17870 40345
rect 17623 40318 17742 40336
tri 17623 40281 17660 40318 ne
rect 17660 40290 17742 40318
rect 17788 40318 17870 40336
tri 17870 40318 17897 40345 sw
rect 70802 40326 70824 40372
rect 70870 40326 70928 40372
rect 70974 40326 71000 40372
rect 17788 40290 17897 40318
rect 17660 40281 17897 40290
tri 17660 40268 17673 40281 ne
rect 17673 40273 17897 40281
tri 17897 40273 17942 40318 sw
rect 17673 40268 17942 40273
tri 17942 40268 17947 40273 sw
rect 70802 40268 71000 40326
tri 17673 40236 17705 40268 ne
rect 17705 40258 17947 40268
tri 17947 40258 17957 40268 sw
rect 17705 40236 17957 40258
tri 17705 40191 17750 40236 ne
rect 17750 40226 17957 40236
tri 17957 40226 17989 40258 sw
rect 17750 40213 17989 40226
tri 17989 40213 18002 40226 sw
rect 70802 40222 70824 40268
rect 70870 40222 70928 40268
rect 70974 40222 71000 40268
rect 17750 40204 18002 40213
rect 17750 40191 17874 40204
tri 17750 40182 17759 40191 ne
rect 17759 40182 17874 40191
tri 17759 40149 17792 40182 ne
rect 17792 40158 17874 40182
rect 17920 40182 18002 40204
tri 18002 40182 18033 40213 sw
rect 17920 40181 18033 40182
tri 18033 40181 18034 40182 sw
rect 17920 40158 18034 40181
rect 17792 40149 18034 40158
tri 17792 40136 17805 40149 ne
rect 17805 40136 18034 40149
tri 18034 40136 18079 40181 sw
rect 70802 40164 71000 40222
tri 17805 40104 17837 40136 ne
rect 17837 40126 18079 40136
tri 18079 40126 18089 40136 sw
rect 17837 40104 18089 40126
tri 17837 40094 17847 40104 ne
rect 17847 40094 18089 40104
tri 18089 40094 18121 40126 sw
rect 70802 40118 70824 40164
rect 70870 40118 70928 40164
rect 70974 40118 71000 40164
tri 17847 40049 17892 40094 ne
rect 17892 40081 18121 40094
tri 18121 40081 18134 40094 sw
rect 17892 40072 18134 40081
rect 17892 40049 18006 40072
tri 17892 40004 17937 40049 ne
rect 17937 40026 18006 40049
rect 18052 40049 18134 40072
tri 18134 40049 18166 40081 sw
rect 70802 40060 71000 40118
rect 18052 40026 18166 40049
rect 17937 40004 18166 40026
tri 18166 40004 18211 40049 sw
rect 70802 40014 70824 40060
rect 70870 40014 70928 40060
rect 70974 40014 71000 40060
tri 17937 39999 17942 40004 ne
rect 17942 39999 18211 40004
tri 17942 39953 17987 39999 ne
rect 17987 39994 18211 39999
tri 18211 39994 18221 40004 sw
rect 17987 39962 18221 39994
tri 18221 39962 18253 39994 sw
rect 17987 39953 18253 39962
tri 18253 39953 18262 39962 sw
rect 70802 39956 71000 40014
tri 17987 39908 18033 39953 ne
rect 18033 39940 18262 39953
rect 18033 39908 18138 39940
tri 18033 39885 18056 39908 ne
rect 18056 39894 18138 39908
rect 18184 39908 18262 39940
tri 18262 39908 18307 39953 sw
rect 70802 39910 70824 39956
rect 70870 39910 70928 39956
rect 70974 39910 71000 39956
rect 18184 39894 18307 39908
rect 18056 39885 18307 39894
tri 18056 39872 18069 39885 ne
rect 18069 39872 18307 39885
tri 18307 39872 18343 39908 sw
tri 18069 39840 18101 39872 ne
rect 18101 39862 18343 39872
tri 18343 39862 18353 39872 sw
rect 18101 39840 18353 39862
tri 18101 39830 18111 39840 ne
rect 18111 39830 18353 39840
tri 18353 39830 18385 39862 sw
rect 70802 39852 71000 39910
tri 18111 39785 18156 39830 ne
rect 18156 39817 18385 39830
tri 18385 39817 18398 39830 sw
rect 18156 39808 18398 39817
rect 18156 39785 18270 39808
tri 18156 39753 18188 39785 ne
rect 18188 39762 18270 39785
rect 18316 39785 18398 39808
tri 18398 39785 18430 39817 sw
rect 70802 39806 70824 39852
rect 70870 39806 70928 39852
rect 70974 39806 71000 39852
rect 18316 39762 18430 39785
rect 18188 39753 18430 39762
tri 18188 39740 18201 39753 ne
rect 18201 39740 18430 39753
tri 18430 39740 18475 39785 sw
rect 70802 39748 71000 39806
tri 18201 39708 18233 39740 ne
rect 18233 39730 18475 39740
tri 18475 39730 18485 39740 sw
rect 18233 39708 18485 39730
tri 18233 39663 18278 39708 ne
rect 18278 39698 18485 39708
tri 18485 39698 18517 39730 sw
rect 70802 39702 70824 39748
rect 70870 39702 70928 39748
rect 70974 39702 71000 39748
rect 18278 39685 18517 39698
tri 18517 39685 18530 39698 sw
rect 18278 39679 18530 39685
tri 18530 39679 18537 39685 sw
rect 18278 39676 18537 39679
rect 18278 39663 18402 39676
tri 18278 39634 18307 39663 ne
rect 18307 39633 18402 39663
tri 18307 39608 18333 39633 ne
rect 18333 39630 18402 39633
rect 18448 39633 18537 39676
tri 18537 39633 18582 39679 sw
rect 70802 39644 71000 39702
rect 18448 39630 18582 39633
rect 18333 39608 18582 39630
tri 18582 39608 18607 39633 sw
tri 18333 39576 18365 39608 ne
rect 18365 39598 18607 39608
tri 18607 39598 18617 39608 sw
rect 70802 39598 70824 39644
rect 70870 39598 70928 39644
rect 70974 39598 71000 39644
rect 18365 39576 18617 39598
tri 18365 39566 18375 39576 ne
rect 18375 39566 18617 39576
tri 18617 39566 18649 39598 sw
tri 18375 39521 18420 39566 ne
rect 18420 39544 18649 39566
rect 18420 39521 18534 39544
tri 18420 39489 18452 39521 ne
rect 18452 39498 18534 39521
rect 18580 39543 18649 39544
tri 18649 39543 18672 39566 sw
rect 18580 39521 18672 39543
tri 18672 39521 18694 39543 sw
rect 70802 39540 71000 39598
rect 18580 39498 18694 39521
rect 18452 39489 18694 39498
tri 18452 39476 18465 39489 ne
rect 18465 39476 18694 39489
tri 18694 39476 18739 39521 sw
rect 70802 39494 70824 39540
rect 70870 39494 70928 39540
rect 70974 39494 71000 39540
tri 18465 39444 18497 39476 ne
rect 18497 39466 18739 39476
tri 18739 39466 18749 39476 sw
rect 18497 39444 18749 39466
tri 18497 39399 18542 39444 ne
rect 18542 39434 18749 39444
tri 18749 39434 18781 39466 sw
rect 70802 39436 71000 39494
rect 18542 39421 18781 39434
tri 18781 39421 18794 39434 sw
rect 18542 39412 18794 39421
rect 18542 39399 18666 39412
tri 18542 39359 18582 39399 ne
rect 18582 39366 18666 39399
rect 18712 39404 18794 39412
tri 18794 39404 18811 39421 sw
rect 18712 39366 18811 39404
rect 18582 39359 18811 39366
tri 18811 39359 18856 39404 sw
rect 70802 39390 70824 39436
rect 70870 39390 70928 39436
rect 70974 39390 71000 39436
tri 18582 39357 18584 39359 ne
rect 18584 39357 18856 39359
tri 18584 39344 18597 39357 ne
rect 18597 39344 18856 39357
tri 18856 39344 18871 39359 sw
tri 18597 39312 18629 39344 ne
rect 18629 39334 18871 39344
tri 18871 39334 18881 39344 sw
rect 18629 39312 18881 39334
tri 18629 39302 18639 39312 ne
rect 18639 39302 18881 39312
tri 18881 39302 18913 39334 sw
rect 70802 39332 71000 39390
tri 18639 39269 18672 39302 ne
rect 18672 39289 18913 39302
tri 18913 39289 18926 39302 sw
rect 18672 39280 18926 39289
rect 18672 39269 18798 39280
tri 18672 39224 18717 39269 ne
rect 18717 39234 18798 39269
rect 18844 39269 18926 39280
tri 18926 39269 18946 39289 sw
rect 70802 39286 70824 39332
rect 70870 39286 70928 39332
rect 70974 39286 71000 39332
rect 18844 39234 18946 39269
rect 18717 39224 18946 39234
tri 18946 39224 18991 39269 sw
rect 70802 39228 71000 39286
tri 18717 39212 18729 39224 ne
rect 18729 39212 18991 39224
tri 18991 39212 19003 39224 sw
tri 18729 39180 18761 39212 ne
rect 18761 39202 19003 39212
tri 19003 39202 19013 39212 sw
rect 18761 39180 19013 39202
tri 18761 39135 18806 39180 ne
rect 18806 39170 19013 39180
tri 19013 39170 19045 39202 sw
rect 70802 39182 70824 39228
rect 70870 39182 70928 39228
rect 70974 39182 71000 39228
rect 18806 39157 19045 39170
tri 19045 39157 19058 39170 sw
rect 18806 39148 19058 39157
rect 18806 39135 18930 39148
tri 18806 39093 18848 39135 ne
rect 18848 39102 18930 39135
rect 18976 39130 19058 39148
tri 19058 39130 19085 39157 sw
rect 18976 39102 19085 39130
rect 18848 39093 19085 39102
tri 18848 39085 18856 39093 ne
rect 18856 39085 19085 39093
tri 19085 39085 19131 39130 sw
rect 70802 39124 71000 39182
tri 18856 39080 18861 39085 ne
rect 18861 39080 19131 39085
tri 19131 39080 19135 39085 sw
tri 18861 39048 18893 39080 ne
rect 18893 39070 19135 39080
tri 19135 39070 19145 39080 sw
rect 70802 39078 70824 39124
rect 70870 39078 70928 39124
rect 70974 39078 71000 39124
rect 18893 39048 19145 39070
tri 18893 39038 18903 39048 ne
rect 18903 39038 19145 39048
tri 19145 39038 19177 39070 sw
tri 18903 38993 18948 39038 ne
rect 18948 39025 19177 39038
tri 19177 39025 19190 39038 sw
rect 18948 39016 19190 39025
rect 18948 38993 19062 39016
tri 18948 38961 18980 38993 ne
rect 18980 38970 19062 38993
rect 19108 38993 19190 39016
tri 19190 38993 19222 39025 sw
rect 70802 39020 71000 39078
rect 19108 38970 19222 38993
rect 18980 38961 19222 38970
tri 18980 38948 18993 38961 ne
rect 18993 38948 19222 38961
tri 19222 38948 19267 38993 sw
rect 70802 38974 70824 39020
rect 70870 38974 70928 39020
rect 70974 38974 71000 39020
tri 18993 38916 19025 38948 ne
rect 19025 38938 19267 38948
tri 19267 38938 19277 38948 sw
rect 19025 38916 19277 38938
tri 19025 38904 19037 38916 ne
rect 19037 38906 19277 38916
tri 19277 38906 19309 38938 sw
rect 70802 38916 71000 38974
rect 19037 38904 19309 38906
tri 19037 38859 19082 38904 ne
rect 19082 38893 19309 38904
tri 19309 38893 19322 38906 sw
rect 19082 38884 19322 38893
rect 19082 38859 19194 38884
tri 19082 38829 19112 38859 ne
rect 19112 38838 19194 38859
rect 19240 38859 19322 38884
tri 19322 38859 19356 38893 sw
rect 70802 38870 70824 38916
rect 70870 38870 70928 38916
rect 70974 38870 71000 38916
rect 19240 38838 19356 38859
rect 19112 38829 19356 38838
tri 19112 38810 19131 38829 ne
rect 19131 38816 19356 38829
tri 19356 38816 19399 38859 sw
rect 19131 38814 19399 38816
tri 19399 38814 19401 38816 sw
rect 19131 38810 19401 38814
tri 19401 38810 19405 38814 sw
rect 70802 38812 71000 38870
tri 19131 38784 19157 38810 ne
rect 19157 38806 19405 38810
tri 19405 38806 19409 38810 sw
rect 19157 38784 19409 38806
tri 19157 38774 19167 38784 ne
rect 19167 38774 19409 38784
tri 19409 38774 19441 38806 sw
tri 19167 38729 19212 38774 ne
rect 19212 38761 19441 38774
tri 19441 38761 19454 38774 sw
rect 70802 38766 70824 38812
rect 70870 38766 70928 38812
rect 70974 38766 71000 38812
rect 19212 38752 19454 38761
rect 19212 38729 19326 38752
tri 19212 38697 19244 38729 ne
rect 19244 38706 19326 38729
rect 19372 38729 19454 38752
tri 19454 38729 19486 38761 sw
rect 19372 38706 19486 38729
rect 19244 38697 19486 38706
tri 19244 38684 19257 38697 ne
rect 19257 38684 19486 38697
tri 19486 38684 19531 38729 sw
rect 70802 38708 71000 38766
tri 19257 38652 19289 38684 ne
rect 19289 38674 19531 38684
tri 19531 38674 19541 38684 sw
rect 19289 38652 19541 38674
tri 19289 38607 19334 38652 ne
rect 19334 38642 19541 38652
tri 19541 38642 19573 38674 sw
rect 70802 38662 70824 38708
rect 70870 38662 70928 38708
rect 70974 38662 71000 38708
rect 19334 38629 19573 38642
tri 19573 38629 19586 38642 sw
rect 19334 38620 19586 38629
rect 19334 38607 19458 38620
tri 19334 38585 19356 38607 ne
rect 19356 38585 19458 38607
tri 19356 38539 19401 38585 ne
rect 19401 38574 19458 38585
rect 19504 38597 19586 38620
tri 19586 38597 19618 38629 sw
rect 70802 38604 71000 38662
rect 19504 38574 19618 38597
rect 19401 38552 19618 38574
tri 19618 38552 19663 38597 sw
rect 70802 38558 70824 38604
rect 70870 38558 70928 38604
rect 70974 38558 71000 38604
rect 19401 38542 19663 38552
tri 19663 38542 19673 38552 sw
rect 19401 38539 19673 38542
tri 19401 38536 19405 38539 ne
rect 19405 38536 19673 38539
tri 19673 38536 19679 38542 sw
tri 19405 38510 19431 38536 ne
rect 19431 38510 19679 38536
tri 19679 38510 19705 38536 sw
tri 19431 38494 19447 38510 ne
rect 19447 38497 19705 38510
tri 19705 38497 19718 38510 sw
rect 70802 38500 71000 38558
rect 19447 38494 19718 38497
tri 19718 38494 19721 38497 sw
tri 19447 38449 19492 38494 ne
rect 19492 38488 19721 38494
rect 19492 38449 19590 38488
tri 19492 38433 19508 38449 ne
rect 19508 38442 19590 38449
rect 19636 38449 19721 38488
tri 19721 38449 19766 38494 sw
rect 70802 38454 70824 38500
rect 70870 38454 70928 38500
rect 70974 38454 71000 38500
rect 19636 38442 19766 38449
rect 19508 38433 19766 38442
tri 19508 38420 19521 38433 ne
rect 19521 38420 19766 38433
tri 19766 38420 19795 38449 sw
tri 19521 38388 19553 38420 ne
rect 19553 38410 19795 38420
tri 19795 38410 19805 38420 sw
rect 19553 38388 19805 38410
tri 19553 38343 19598 38388 ne
rect 19598 38378 19805 38388
tri 19805 38378 19837 38410 sw
rect 70802 38396 71000 38454
rect 19598 38365 19837 38378
tri 19837 38365 19850 38378 sw
rect 19598 38356 19850 38365
rect 19598 38343 19722 38356
tri 19598 38301 19640 38343 ne
rect 19640 38310 19722 38343
rect 19768 38333 19850 38356
tri 19850 38333 19882 38365 sw
rect 70802 38350 70824 38396
rect 70870 38350 70928 38396
rect 70974 38350 71000 38396
rect 19768 38310 19882 38333
rect 19640 38301 19882 38310
tri 19640 38261 19679 38301 ne
rect 19679 38288 19882 38301
tri 19882 38288 19927 38333 sw
rect 70802 38292 71000 38350
rect 19679 38278 19927 38288
tri 19927 38278 19937 38288 sw
rect 19679 38261 19937 38278
tri 19937 38261 19954 38278 sw
tri 19679 38256 19685 38261 ne
rect 19685 38256 19954 38261
tri 19685 38246 19695 38256 ne
rect 19695 38246 19954 38256
tri 19954 38246 19969 38261 sw
rect 70802 38246 70824 38292
rect 70870 38246 70928 38292
rect 70974 38246 71000 38292
tri 19695 38201 19740 38246 ne
rect 19740 38233 19969 38246
tri 19969 38233 19982 38246 sw
rect 19740 38224 19982 38233
rect 19740 38201 19854 38224
tri 19740 38175 19766 38201 ne
rect 19766 38178 19854 38201
rect 19900 38201 19982 38224
tri 19982 38201 20014 38233 sw
rect 19900 38178 20014 38201
rect 19766 38175 20014 38178
tri 19766 38156 19785 38175 ne
rect 19785 38156 20014 38175
tri 20014 38156 20059 38201 sw
rect 70802 38188 71000 38246
tri 19785 38124 19817 38156 ne
rect 19817 38146 20059 38156
tri 20059 38146 20069 38156 sw
rect 19817 38124 20069 38146
tri 19817 38079 19862 38124 ne
rect 19862 38114 20069 38124
tri 20069 38114 20101 38146 sw
rect 70802 38142 70824 38188
rect 70870 38142 70928 38188
rect 70974 38142 71000 38188
rect 19862 38092 20101 38114
rect 19862 38079 19986 38092
tri 19862 38037 19904 38079 ne
rect 19904 38046 19986 38079
rect 20032 38084 20101 38092
tri 20101 38084 20131 38114 sw
rect 70802 38084 71000 38142
rect 20032 38069 20131 38084
tri 20131 38069 20146 38084 sw
rect 20032 38046 20146 38069
rect 19904 38037 20146 38046
tri 19904 37992 19949 38037 ne
rect 19949 38024 20146 38037
tri 20146 38024 20191 38069 sw
rect 70802 38038 70824 38084
rect 70870 38038 70928 38084
rect 70974 38038 71000 38084
rect 19949 38014 20191 38024
tri 20191 38014 20201 38024 sw
rect 19949 37992 20201 38014
tri 19949 37987 19954 37992 ne
rect 19954 37987 20201 37992
tri 20201 37987 20228 38014 sw
tri 19954 37982 19959 37987 ne
rect 19959 37982 20228 37987
tri 20228 37982 20233 37987 sw
tri 19959 37937 20004 37982 ne
rect 20004 37969 20233 37982
tri 20233 37969 20246 37982 sw
rect 70802 37980 71000 38038
rect 20004 37960 20246 37969
rect 20004 37937 20118 37960
tri 20004 37905 20036 37937 ne
rect 20036 37914 20118 37937
rect 20164 37937 20246 37960
tri 20246 37937 20278 37969 sw
rect 20164 37914 20278 37937
rect 20036 37905 20278 37914
tri 20036 37892 20049 37905 ne
rect 20049 37892 20278 37905
tri 20278 37892 20323 37937 sw
rect 70802 37934 70824 37980
rect 70870 37934 70928 37980
rect 70974 37934 71000 37980
tri 20049 37860 20081 37892 ne
rect 20081 37882 20323 37892
tri 20323 37882 20333 37892 sw
rect 20081 37860 20333 37882
tri 20081 37850 20091 37860 ne
rect 20091 37850 20333 37860
tri 20333 37850 20365 37882 sw
rect 70802 37876 71000 37934
tri 20091 37810 20131 37850 ne
rect 20131 37837 20365 37850
tri 20365 37837 20378 37850 sw
rect 20131 37828 20378 37837
rect 20131 37810 20250 37828
tri 20131 37765 20176 37810 ne
rect 20176 37782 20250 37810
rect 20296 37810 20378 37828
tri 20378 37810 20405 37837 sw
rect 70802 37830 70824 37876
rect 70870 37830 70928 37876
rect 70974 37830 71000 37876
rect 20296 37782 20405 37810
rect 20176 37765 20405 37782
tri 20405 37765 20451 37810 sw
rect 70802 37772 71000 37830
tri 20176 37760 20181 37765 ne
rect 20181 37760 20451 37765
tri 20451 37760 20455 37765 sw
tri 20181 37728 20213 37760 ne
rect 20213 37750 20455 37760
tri 20455 37750 20465 37760 sw
rect 20213 37728 20465 37750
tri 20213 37713 20228 37728 ne
rect 20228 37718 20465 37728
tri 20465 37718 20497 37750 sw
rect 70802 37726 70824 37772
rect 70870 37726 70928 37772
rect 70974 37726 71000 37772
rect 20228 37713 20497 37718
tri 20497 37713 20503 37718 sw
tri 20228 37667 20273 37713 ne
rect 20273 37705 20503 37713
tri 20503 37705 20510 37713 sw
rect 20273 37696 20510 37705
rect 20273 37667 20382 37696
tri 20273 37641 20300 37667 ne
rect 20300 37650 20382 37667
rect 20428 37673 20510 37696
tri 20510 37673 20542 37705 sw
rect 20428 37650 20542 37673
rect 20300 37641 20542 37650
tri 20300 37628 20313 37641 ne
rect 20313 37628 20542 37641
tri 20542 37628 20587 37673 sw
rect 70802 37668 71000 37726
tri 20313 37596 20345 37628 ne
rect 20345 37618 20587 37628
tri 20587 37618 20597 37628 sw
rect 70802 37622 70824 37668
rect 70870 37622 70928 37668
rect 70974 37622 71000 37668
rect 20345 37596 20597 37618
tri 20345 37586 20355 37596 ne
rect 20355 37586 20597 37596
tri 20597 37586 20629 37618 sw
tri 20355 37541 20400 37586 ne
rect 20400 37573 20629 37586
tri 20629 37573 20642 37586 sw
rect 20400 37564 20642 37573
rect 20400 37541 20514 37564
tri 20400 37509 20432 37541 ne
rect 20432 37518 20514 37541
rect 20560 37541 20642 37564
tri 20642 37541 20674 37573 sw
rect 70802 37564 71000 37622
rect 20560 37518 20674 37541
rect 20432 37509 20674 37518
tri 20432 37496 20445 37509 ne
rect 20445 37496 20674 37509
tri 20674 37496 20719 37541 sw
rect 70802 37518 70824 37564
rect 70870 37518 70928 37564
rect 70974 37518 71000 37564
tri 20445 37464 20477 37496 ne
rect 20477 37486 20719 37496
tri 20719 37486 20729 37496 sw
rect 20477 37464 20729 37486
tri 20477 37445 20496 37464 ne
rect 20496 37454 20729 37464
tri 20729 37454 20761 37486 sw
rect 70802 37460 71000 37518
rect 20496 37445 20761 37454
tri 20496 37438 20503 37445 ne
rect 20503 37441 20761 37445
tri 20761 37441 20774 37454 sw
rect 20503 37438 20774 37441
tri 20774 37438 20777 37441 sw
tri 20503 37400 20541 37438 ne
rect 20541 37432 20777 37438
rect 20541 37400 20646 37432
tri 20541 37377 20564 37400 ne
rect 20564 37386 20646 37400
rect 20692 37400 20777 37432
tri 20777 37400 20815 37438 sw
rect 70802 37414 70824 37460
rect 70870 37414 70928 37460
rect 70974 37414 71000 37460
rect 20692 37386 20815 37400
rect 20564 37377 20815 37386
tri 20564 37364 20577 37377 ne
rect 20577 37364 20815 37377
tri 20815 37364 20851 37400 sw
tri 20577 37332 20609 37364 ne
rect 20609 37355 20851 37364
tri 20851 37355 20861 37364 sw
rect 20609 37332 20861 37355
rect 70802 37356 71000 37414
tri 20609 37322 20619 37332 ne
rect 20619 37322 20861 37332
tri 20861 37322 20893 37354 sw
tri 20619 37277 20664 37322 ne
rect 20664 37309 20893 37322
tri 20893 37309 20906 37322 sw
rect 70802 37310 70824 37356
rect 70870 37310 70928 37356
rect 70974 37310 71000 37356
rect 20664 37300 20906 37309
rect 20664 37277 20778 37300
tri 20664 37245 20696 37277 ne
rect 20696 37254 20778 37277
rect 20824 37277 20906 37300
tri 20906 37277 20938 37309 sw
rect 20824 37254 20938 37277
rect 20696 37245 20938 37254
tri 20696 37232 20709 37245 ne
rect 20709 37232 20938 37245
tri 20938 37232 20983 37277 sw
rect 70802 37252 71000 37310
tri 20709 37200 20741 37232 ne
rect 20741 37222 20983 37232
tri 20983 37222 20993 37232 sw
rect 20741 37200 20993 37222
tri 20741 37164 20777 37200 ne
rect 20777 37190 20993 37200
tri 20993 37190 21025 37222 sw
rect 70802 37206 70824 37252
rect 70870 37206 70928 37252
rect 70974 37206 71000 37252
rect 20777 37177 21025 37190
tri 21025 37177 21038 37190 sw
rect 20777 37168 21038 37177
rect 20777 37164 20910 37168
tri 20777 37119 20822 37164 ne
rect 20822 37122 20910 37164
rect 20956 37164 21038 37168
tri 21038 37164 21051 37177 sw
rect 20956 37145 21051 37164
tri 21051 37145 21070 37164 sw
rect 70802 37148 71000 37206
rect 20956 37122 21070 37145
rect 20822 37119 21070 37122
tri 20822 37113 20828 37119 ne
rect 20828 37113 21070 37119
tri 20828 37100 20841 37113 ne
rect 20841 37100 21070 37113
tri 21070 37100 21115 37145 sw
rect 70802 37102 70824 37148
rect 70870 37102 70928 37148
rect 70974 37102 71000 37148
tri 20841 37068 20873 37100 ne
rect 20873 37090 21115 37100
tri 21115 37090 21125 37100 sw
rect 20873 37068 21125 37090
tri 20873 37058 20883 37068 ne
rect 20883 37058 21125 37068
tri 21125 37058 21157 37090 sw
tri 20883 37035 20906 37058 ne
rect 20906 37045 21157 37058
tri 21157 37045 21170 37058 sw
rect 20906 37036 21170 37045
rect 20906 37035 21042 37036
tri 20906 36990 20951 37035 ne
rect 20951 36990 21042 37035
rect 21088 37035 21170 37036
tri 21170 37035 21180 37045 sw
rect 70802 37044 71000 37102
rect 21088 36990 21180 37035
tri 21180 36990 21225 37035 sw
rect 70802 36998 70824 37044
rect 70870 36998 70928 37044
rect 70974 36998 71000 37044
tri 20951 36981 20960 36990 ne
rect 20960 36981 21225 36990
tri 20960 36968 20973 36981 ne
rect 20973 36968 21225 36981
tri 21225 36968 21247 36990 sw
tri 20973 36936 21005 36968 ne
rect 21005 36958 21247 36968
tri 21247 36958 21257 36968 sw
rect 21005 36936 21257 36958
tri 21005 36891 21050 36936 ne
rect 21050 36926 21257 36936
tri 21257 36926 21289 36958 sw
rect 70802 36940 71000 36998
rect 21050 36913 21289 36926
tri 21289 36913 21302 36926 sw
rect 21050 36904 21302 36913
rect 21050 36891 21174 36904
tri 21050 36889 21051 36891 ne
rect 21051 36889 21174 36891
tri 21051 36849 21092 36889 ne
rect 21092 36858 21174 36889
rect 21220 36889 21302 36904
tri 21302 36889 21326 36913 sw
rect 70802 36894 70824 36940
rect 70870 36894 70928 36940
rect 70974 36894 71000 36940
rect 21220 36881 21326 36889
tri 21326 36881 21334 36889 sw
rect 21220 36858 21334 36881
rect 21092 36849 21334 36858
tri 21092 36836 21105 36849 ne
rect 21105 36836 21334 36849
tri 21334 36836 21379 36881 sw
rect 70802 36836 71000 36894
tri 21105 36804 21137 36836 ne
rect 21137 36826 21379 36836
tri 21379 36826 21389 36836 sw
rect 21137 36804 21389 36826
tri 21137 36794 21147 36804 ne
rect 21147 36794 21389 36804
tri 21389 36794 21421 36826 sw
tri 21147 36749 21192 36794 ne
rect 21192 36781 21421 36794
tri 21421 36781 21434 36794 sw
rect 70802 36790 70824 36836
rect 70870 36790 70928 36836
rect 70974 36790 71000 36836
rect 21192 36772 21434 36781
rect 21192 36749 21306 36772
tri 21192 36715 21225 36749 ne
rect 21225 36726 21306 36749
rect 21352 36749 21434 36772
tri 21434 36749 21466 36781 sw
rect 21352 36726 21466 36749
rect 21225 36715 21466 36726
tri 21225 36704 21237 36715 ne
rect 21237 36704 21466 36715
tri 21466 36704 21511 36749 sw
rect 70802 36732 71000 36790
tri 21237 36670 21271 36704 ne
rect 21271 36694 21511 36704
tri 21511 36694 21521 36704 sw
rect 21271 36670 21521 36694
tri 21271 36625 21316 36670 ne
rect 21316 36662 21521 36670
tri 21521 36662 21553 36694 sw
rect 70802 36686 70824 36732
rect 70870 36686 70928 36732
rect 70974 36686 71000 36732
rect 21316 36640 21553 36662
rect 21316 36625 21438 36640
tri 21316 36615 21326 36625 ne
rect 21326 36615 21438 36625
tri 21326 36585 21356 36615 ne
rect 21356 36594 21438 36615
rect 21484 36625 21553 36640
tri 21553 36625 21590 36662 sw
rect 70802 36628 71000 36686
rect 21484 36615 21590 36625
tri 21590 36615 21600 36625 sw
rect 21484 36594 21600 36615
rect 21356 36585 21600 36594
tri 21356 36572 21369 36585 ne
rect 21369 36572 21600 36585
tri 21600 36572 21643 36615 sw
rect 70802 36582 70824 36628
rect 70870 36582 70928 36628
rect 70974 36582 71000 36628
tri 21369 36540 21401 36572 ne
rect 21401 36562 21643 36572
tri 21643 36562 21653 36572 sw
rect 21401 36540 21653 36562
tri 21401 36530 21411 36540 ne
rect 21411 36530 21653 36540
tri 21653 36530 21685 36562 sw
tri 21411 36485 21456 36530 ne
rect 21456 36517 21685 36530
tri 21685 36517 21698 36530 sw
rect 70802 36524 71000 36582
rect 21456 36508 21698 36517
rect 21456 36485 21570 36508
tri 21456 36453 21488 36485 ne
rect 21488 36462 21570 36485
rect 21616 36485 21698 36508
tri 21698 36485 21730 36517 sw
rect 21616 36462 21730 36485
rect 21488 36453 21730 36462
tri 21488 36440 21501 36453 ne
rect 21501 36440 21730 36453
tri 21730 36440 21775 36485 sw
rect 70802 36478 70824 36524
rect 70870 36478 70928 36524
rect 70974 36478 71000 36524
tri 21501 36408 21533 36440 ne
rect 21533 36430 21775 36440
tri 21775 36430 21785 36440 sw
rect 21533 36408 21785 36430
tri 21533 36363 21578 36408 ne
rect 21578 36398 21785 36408
tri 21785 36398 21817 36430 sw
rect 70802 36420 71000 36478
rect 21578 36385 21817 36398
tri 21817 36385 21830 36398 sw
rect 21578 36376 21830 36385
rect 21578 36363 21702 36376
tri 21578 36351 21590 36363 ne
rect 21590 36351 21702 36363
tri 21590 36341 21600 36351 ne
rect 21600 36341 21702 36351
tri 21600 36308 21633 36341 ne
rect 21633 36330 21702 36341
rect 21748 36341 21830 36376
tri 21830 36341 21875 36385 sw
rect 70802 36374 70824 36420
rect 70870 36374 70928 36420
rect 70974 36374 71000 36420
rect 21748 36330 21875 36341
rect 21633 36308 21875 36330
tri 21875 36308 21907 36341 sw
rect 70802 36316 71000 36374
tri 21633 36276 21665 36308 ne
rect 21665 36305 21907 36308
tri 21907 36305 21910 36308 sw
rect 21665 36276 21910 36305
tri 21665 36266 21675 36276 ne
rect 21675 36266 21910 36276
tri 21910 36266 21949 36305 sw
rect 70802 36270 70824 36316
rect 70870 36270 70928 36316
rect 70974 36270 71000 36316
tri 21675 36221 21720 36266 ne
rect 21720 36253 21949 36266
tri 21949 36253 21962 36266 sw
rect 21720 36244 21962 36253
rect 21720 36221 21834 36244
tri 21720 36189 21752 36221 ne
rect 21752 36198 21834 36221
rect 21880 36221 21962 36244
tri 21962 36221 21994 36253 sw
rect 21880 36198 21994 36221
rect 21752 36189 21994 36198
tri 21752 36176 21765 36189 ne
rect 21765 36176 21994 36189
tri 21994 36176 22039 36221 sw
rect 70802 36212 71000 36270
tri 21765 36144 21797 36176 ne
rect 21797 36166 22039 36176
tri 22039 36166 22049 36176 sw
rect 70802 36166 70824 36212
rect 70870 36166 70928 36212
rect 70974 36166 71000 36212
rect 21797 36144 22049 36166
tri 21797 36099 21842 36144 ne
rect 21842 36134 22049 36144
tri 22049 36134 22081 36166 sw
rect 21842 36121 22081 36134
tri 22081 36121 22094 36134 sw
rect 21842 36112 22094 36121
rect 21842 36099 21966 36112
tri 21842 36066 21875 36099 ne
rect 21875 36066 21966 36099
rect 22012 36111 22094 36112
tri 22094 36111 22104 36121 sw
rect 22012 36066 22104 36111
tri 22104 36066 22149 36111 sw
rect 70802 36108 71000 36166
tri 21875 36057 21884 36066 ne
rect 21884 36057 22149 36066
tri 21884 36044 21897 36057 ne
rect 21897 36044 22149 36057
tri 22149 36044 22171 36066 sw
rect 70802 36062 70824 36108
rect 70870 36062 70928 36108
rect 70974 36062 71000 36108
tri 21897 36012 21929 36044 ne
rect 21929 36034 22171 36044
tri 22171 36034 22181 36044 sw
rect 21929 36012 22181 36034
tri 21929 36002 21939 36012 ne
rect 21939 36002 22181 36012
tri 22181 36002 22213 36034 sw
rect 70802 36004 71000 36062
tri 21939 35986 21955 36002 ne
rect 21955 35989 22213 36002
tri 22213 35989 22226 36002 sw
rect 21955 35986 22226 35989
tri 22226 35986 22229 35989 sw
tri 21955 35941 22000 35986 ne
rect 22000 35980 22229 35986
rect 22000 35941 22098 35980
tri 22000 35925 22016 35941 ne
rect 22016 35934 22098 35941
rect 22144 35941 22229 35980
tri 22229 35941 22275 35986 sw
rect 70802 35958 70824 36004
rect 70870 35958 70928 36004
rect 70974 35958 71000 36004
rect 22144 35934 22275 35941
rect 22016 35925 22275 35934
tri 22016 35912 22029 35925 ne
rect 22029 35912 22275 35925
tri 22275 35912 22303 35941 sw
tri 22029 35880 22061 35912 ne
rect 22061 35902 22303 35912
tri 22303 35902 22313 35912 sw
rect 22061 35880 22313 35902
tri 22061 35835 22106 35880 ne
rect 22106 35870 22313 35880
tri 22313 35870 22345 35902 sw
rect 70802 35900 71000 35958
rect 22106 35857 22345 35870
tri 22345 35857 22358 35870 sw
rect 22106 35848 22358 35857
rect 22106 35835 22230 35848
tri 22106 35793 22148 35835 ne
rect 22148 35802 22230 35835
rect 22276 35837 22358 35848
tri 22358 35837 22378 35857 sw
rect 70802 35854 70824 35900
rect 70870 35854 70928 35900
rect 70974 35854 71000 35900
rect 22276 35802 22378 35837
rect 22148 35793 22378 35802
tri 22148 35792 22149 35793 ne
rect 22149 35792 22378 35793
tri 22378 35792 22423 35837 sw
rect 70802 35796 71000 35854
tri 22149 35780 22161 35792 ne
rect 22161 35780 22423 35792
tri 22423 35780 22435 35792 sw
tri 22161 35748 22193 35780 ne
rect 22193 35770 22435 35780
tri 22435 35770 22445 35780 sw
rect 22193 35748 22445 35770
tri 22193 35738 22203 35748 ne
rect 22203 35738 22445 35748
tri 22445 35738 22477 35770 sw
rect 70802 35750 70824 35796
rect 70870 35750 70928 35796
rect 70974 35750 71000 35796
tri 22203 35693 22248 35738 ne
rect 22248 35725 22477 35738
tri 22477 35725 22490 35738 sw
rect 22248 35716 22490 35725
rect 22248 35693 22362 35716
tri 22248 35661 22280 35693 ne
rect 22280 35670 22362 35693
rect 22408 35693 22490 35716
tri 22490 35693 22522 35725 sw
rect 22408 35670 22522 35693
rect 22280 35661 22522 35670
tri 22280 35648 22293 35661 ne
rect 22293 35648 22522 35661
tri 22522 35648 22567 35693 sw
rect 70802 35692 71000 35750
tri 22293 35616 22325 35648 ne
rect 22325 35638 22567 35648
tri 22567 35638 22577 35648 sw
rect 70802 35646 70824 35692
rect 70870 35646 70928 35692
rect 70974 35646 71000 35692
rect 22325 35616 22577 35638
tri 22325 35576 22365 35616 ne
rect 22365 35606 22577 35616
tri 22577 35606 22609 35638 sw
rect 22365 35593 22609 35606
tri 22609 35593 22622 35606 sw
rect 22365 35584 22622 35593
rect 22365 35576 22494 35584
tri 22365 35531 22410 35576 ne
rect 22410 35538 22494 35576
rect 22540 35576 22622 35584
tri 22622 35576 22639 35593 sw
rect 70802 35588 71000 35646
rect 22540 35538 22639 35576
rect 22410 35531 22639 35538
tri 22639 35531 22685 35576 sw
rect 70802 35542 70824 35588
rect 70870 35542 70928 35588
rect 70974 35542 71000 35588
tri 22410 35529 22412 35531 ne
rect 22412 35529 22685 35531
tri 22412 35517 22423 35529 ne
rect 22423 35517 22685 35529
tri 22685 35517 22698 35531 sw
tri 22423 35516 22425 35517 ne
rect 22425 35516 22698 35517
tri 22698 35516 22699 35517 sw
tri 22425 35484 22457 35516 ne
rect 22457 35506 22699 35516
tri 22699 35506 22709 35516 sw
rect 22457 35484 22709 35506
tri 22457 35474 22467 35484 ne
rect 22467 35474 22709 35484
tri 22709 35474 22741 35506 sw
rect 70802 35484 71000 35542
tri 22467 35429 22512 35474 ne
rect 22512 35461 22741 35474
tri 22741 35461 22754 35474 sw
rect 22512 35452 22754 35461
rect 22512 35429 22626 35452
tri 22512 35397 22544 35429 ne
rect 22544 35406 22626 35429
rect 22672 35429 22754 35452
tri 22754 35429 22786 35461 sw
rect 70802 35438 70824 35484
rect 70870 35438 70928 35484
rect 70974 35438 71000 35484
rect 22672 35406 22786 35429
rect 22544 35397 22786 35406
tri 22544 35384 22557 35397 ne
rect 22557 35384 22786 35397
tri 22786 35384 22831 35429 sw
tri 22557 35352 22589 35384 ne
rect 22589 35374 22831 35384
tri 22831 35374 22841 35384 sw
rect 70802 35380 71000 35438
rect 22589 35352 22841 35374
tri 22589 35307 22634 35352 ne
rect 22634 35342 22841 35352
tri 22841 35342 22873 35374 sw
rect 22634 35329 22873 35342
tri 22873 35329 22886 35342 sw
rect 70802 35334 70824 35380
rect 70870 35334 70928 35380
rect 70974 35334 71000 35380
rect 22634 35320 22886 35329
rect 22634 35307 22758 35320
tri 22634 35301 22639 35307 ne
rect 22639 35301 22758 35307
tri 22639 35256 22685 35301 ne
rect 22685 35274 22758 35301
rect 22804 35297 22886 35320
tri 22886 35297 22918 35329 sw
rect 22804 35274 22918 35297
rect 22685 35256 22918 35274
tri 22685 35243 22698 35256 ne
rect 22698 35252 22918 35256
tri 22918 35252 22963 35297 sw
rect 70802 35276 71000 35334
rect 22698 35243 22963 35252
tri 22963 35243 22972 35252 sw
tri 22698 35211 22730 35243 ne
rect 22730 35242 22972 35243
tri 22972 35242 22973 35243 sw
rect 22730 35211 22973 35242
tri 22730 35210 22731 35211 ne
rect 22731 35210 22973 35211
tri 22973 35210 23005 35242 sw
rect 70802 35230 70824 35276
rect 70870 35230 70928 35276
rect 70974 35230 71000 35276
tri 22731 35165 22776 35210 ne
rect 22776 35188 23005 35210
rect 22776 35165 22890 35188
tri 22776 35133 22808 35165 ne
rect 22808 35142 22890 35165
rect 22936 35166 23005 35188
tri 23005 35166 23049 35210 sw
rect 70802 35172 71000 35230
rect 22936 35165 23049 35166
tri 23049 35165 23050 35166 sw
rect 22936 35142 23050 35165
rect 22808 35133 23050 35142
tri 22808 35120 22821 35133 ne
rect 22821 35120 23050 35133
tri 23050 35120 23095 35165 sw
rect 70802 35126 70824 35172
rect 70870 35126 70928 35172
rect 70974 35126 71000 35172
tri 22821 35088 22853 35120 ne
rect 22853 35110 23095 35120
tri 23095 35110 23105 35120 sw
rect 22853 35088 23105 35110
tri 22853 35043 22898 35088 ne
rect 22898 35078 23105 35088
tri 23105 35078 23137 35110 sw
rect 22898 35065 23137 35078
tri 23137 35065 23150 35078 sw
rect 70802 35068 71000 35126
rect 22898 35056 23150 35065
rect 22898 35043 23022 35056
tri 22898 35001 22940 35043 ne
rect 22940 35010 23022 35043
rect 23068 35033 23150 35056
tri 23150 35033 23182 35065 sw
rect 23068 35010 23182 35033
rect 22940 35001 23182 35010
tri 22940 34969 22972 35001 ne
rect 22972 34988 23182 35001
tri 23182 34988 23227 35033 sw
rect 70802 35022 70824 35068
rect 70870 35022 70928 35068
rect 70974 35022 71000 35068
rect 22972 34978 23227 34988
tri 23227 34978 23237 34988 sw
rect 22972 34969 23237 34978
tri 23237 34969 23247 34978 sw
tri 22972 34956 22985 34969 ne
rect 22985 34956 23247 34969
tri 22985 34946 22995 34956 ne
rect 22995 34946 23247 34956
tri 23247 34946 23269 34969 sw
rect 70802 34964 71000 35022
tri 22995 34901 23040 34946 ne
rect 23040 34933 23269 34946
tri 23269 34933 23282 34946 sw
rect 23040 34924 23282 34933
rect 23040 34901 23154 34924
tri 23040 34891 23049 34901 ne
rect 23049 34891 23154 34901
tri 23049 34856 23085 34891 ne
rect 23085 34878 23154 34891
rect 23200 34901 23282 34924
tri 23282 34901 23314 34933 sw
rect 70802 34918 70824 34964
rect 70870 34918 70928 34964
rect 70974 34918 71000 34964
rect 23200 34878 23314 34901
rect 23085 34856 23314 34878
tri 23314 34856 23359 34901 sw
rect 70802 34860 71000 34918
tri 23085 34824 23117 34856 ne
rect 23117 34846 23359 34856
tri 23359 34846 23369 34856 sw
rect 23117 34824 23369 34846
tri 23117 34779 23162 34824 ne
rect 23162 34814 23369 34824
tri 23369 34814 23401 34846 sw
rect 70802 34814 70824 34860
rect 70870 34814 70928 34860
rect 70974 34814 71000 34860
rect 23162 34801 23401 34814
tri 23401 34801 23414 34814 sw
rect 23162 34792 23414 34801
rect 23162 34779 23286 34792
tri 23162 34737 23204 34779 ne
rect 23204 34746 23286 34779
rect 23332 34769 23414 34792
tri 23414 34769 23446 34801 sw
rect 23332 34746 23446 34769
rect 23204 34737 23446 34746
tri 23204 34694 23247 34737 ne
rect 23247 34724 23446 34737
tri 23446 34724 23491 34769 sw
rect 70802 34756 71000 34814
rect 23247 34714 23491 34724
tri 23491 34714 23501 34724 sw
rect 23247 34694 23501 34714
tri 23501 34694 23521 34714 sw
rect 70802 34710 70824 34756
rect 70870 34710 70928 34756
rect 70974 34710 71000 34756
tri 23247 34692 23249 34694 ne
rect 23249 34692 23521 34694
tri 23249 34682 23259 34692 ne
rect 23259 34682 23521 34692
tri 23521 34682 23533 34694 sw
tri 23259 34637 23304 34682 ne
rect 23304 34669 23533 34682
tri 23533 34669 23546 34682 sw
rect 23304 34660 23546 34669
rect 23304 34637 23418 34660
tri 23304 34605 23336 34637 ne
rect 23336 34614 23418 34637
rect 23464 34637 23546 34660
tri 23546 34637 23578 34669 sw
rect 70802 34652 71000 34710
rect 23464 34614 23578 34637
rect 23336 34605 23578 34614
tri 23336 34592 23349 34605 ne
rect 23349 34592 23578 34605
tri 23578 34592 23623 34637 sw
rect 70802 34606 70824 34652
rect 70870 34606 70928 34652
rect 70974 34606 71000 34652
tri 23349 34560 23381 34592 ne
rect 23381 34582 23623 34592
tri 23623 34582 23633 34592 sw
rect 23381 34560 23633 34582
tri 23381 34527 23414 34560 ne
rect 23414 34550 23633 34560
tri 23633 34550 23665 34582 sw
rect 23414 34537 23665 34550
tri 23665 34537 23678 34550 sw
rect 70802 34548 71000 34606
rect 23414 34528 23678 34537
rect 23414 34527 23550 34528
tri 23414 34481 23459 34527 ne
rect 23459 34482 23550 34527
rect 23596 34527 23678 34528
tri 23678 34527 23689 34537 sw
rect 23596 34482 23689 34527
rect 23459 34481 23689 34482
tri 23689 34481 23734 34527 sw
rect 70802 34502 70824 34548
rect 70870 34502 70928 34548
rect 70974 34502 71000 34548
tri 23459 34473 23468 34481 ne
rect 23468 34473 23734 34481
tri 23468 34428 23513 34473 ne
rect 23513 34460 23734 34473
tri 23734 34460 23755 34481 sw
rect 23513 34450 23755 34460
tri 23755 34450 23765 34460 sw
rect 23513 34428 23765 34450
tri 23513 34420 23521 34428 ne
rect 23521 34420 23765 34428
tri 23765 34420 23795 34450 sw
rect 70802 34444 71000 34502
tri 23521 34418 23523 34420 ne
rect 23523 34418 23795 34420
tri 23795 34418 23797 34420 sw
tri 23523 34373 23568 34418 ne
rect 23568 34405 23797 34418
tri 23797 34405 23810 34418 sw
rect 23568 34396 23810 34405
rect 23568 34373 23682 34396
tri 23568 34341 23600 34373 ne
rect 23600 34350 23682 34373
rect 23728 34373 23810 34396
tri 23810 34373 23842 34405 sw
rect 70802 34398 70824 34444
rect 70870 34398 70928 34444
rect 70974 34398 71000 34444
rect 23728 34350 23842 34373
rect 23600 34341 23842 34350
tri 23600 34328 23613 34341 ne
rect 23613 34328 23842 34341
tri 23842 34328 23887 34373 sw
rect 70802 34340 71000 34398
tri 23613 34296 23645 34328 ne
rect 23645 34318 23887 34328
tri 23887 34318 23897 34328 sw
rect 23645 34296 23897 34318
tri 23645 34286 23655 34296 ne
rect 23655 34286 23897 34296
tri 23897 34286 23929 34318 sw
rect 70802 34294 70824 34340
rect 70870 34294 70928 34340
rect 70974 34294 71000 34340
tri 23655 34241 23700 34286 ne
rect 23700 34273 23929 34286
tri 23929 34273 23942 34286 sw
rect 23700 34264 23942 34273
rect 23700 34241 23814 34264
tri 23700 34209 23732 34241 ne
rect 23732 34218 23814 34241
rect 23860 34241 23942 34264
tri 23942 34241 23974 34273 sw
rect 23860 34218 23974 34241
rect 23732 34209 23974 34218
tri 23732 34196 23745 34209 ne
rect 23745 34196 23974 34209
tri 23974 34196 24019 34241 sw
rect 70802 34236 71000 34294
tri 23745 34164 23777 34196 ne
rect 23777 34186 24019 34196
tri 24019 34186 24029 34196 sw
rect 70802 34190 70824 34236
rect 70870 34190 70928 34236
rect 70974 34190 71000 34236
rect 23777 34164 24029 34186
tri 23777 34162 23779 34164 ne
rect 23779 34162 24029 34164
tri 23779 34145 23795 34162 ne
rect 23795 34154 24029 34162
tri 24029 34154 24061 34186 sw
rect 23795 34145 24061 34154
tri 24061 34145 24070 34154 sw
tri 23795 34117 23824 34145 ne
rect 23824 34141 24070 34145
tri 24070 34141 24074 34145 sw
rect 23824 34132 24074 34141
rect 23824 34117 23946 34132
tri 23824 34077 23864 34117 ne
rect 23864 34086 23946 34117
rect 23992 34117 24074 34132
tri 24074 34117 24099 34141 sw
rect 70802 34132 71000 34190
rect 23992 34086 24099 34117
rect 23864 34077 24099 34086
tri 23864 34064 23877 34077 ne
rect 23877 34071 24099 34077
tri 24099 34071 24144 34117 sw
rect 70802 34086 70824 34132
rect 70870 34086 70928 34132
rect 70974 34086 71000 34132
rect 23877 34064 24144 34071
tri 24144 34064 24151 34071 sw
tri 23877 34032 23909 34064 ne
rect 23909 34054 24151 34064
tri 24151 34054 24161 34064 sw
rect 23909 34032 24161 34054
tri 23909 34022 23919 34032 ne
rect 23919 34022 24161 34032
tri 24161 34022 24193 34054 sw
rect 70802 34028 71000 34086
tri 23919 33977 23964 34022 ne
rect 23964 34009 24193 34022
tri 24193 34009 24206 34022 sw
rect 23964 34000 24206 34009
rect 23964 33977 24078 34000
tri 23964 33945 23996 33977 ne
rect 23996 33954 24078 33977
rect 24124 33977 24206 34000
tri 24206 33977 24238 34009 sw
rect 70802 33982 70824 34028
rect 70870 33982 70928 34028
rect 70974 33982 71000 34028
rect 24124 33954 24238 33977
rect 23996 33945 24238 33954
tri 23996 33932 24009 33945 ne
rect 24009 33932 24238 33945
tri 24238 33932 24283 33977 sw
tri 24009 33900 24041 33932 ne
rect 24041 33922 24283 33932
tri 24283 33922 24293 33932 sw
rect 70802 33924 71000 33982
rect 24041 33900 24293 33922
tri 24041 33871 24070 33900 ne
rect 24070 33890 24293 33900
tri 24293 33890 24325 33922 sw
rect 24070 33877 24325 33890
tri 24325 33877 24338 33890 sw
rect 70802 33878 70824 33924
rect 70870 33878 70928 33924
rect 70974 33878 71000 33924
rect 24070 33871 24338 33877
tri 24338 33871 24344 33877 sw
tri 24070 33826 24115 33871 ne
rect 24115 33868 24344 33871
rect 24115 33826 24210 33868
tri 24115 33800 24141 33826 ne
rect 24141 33822 24210 33826
rect 24256 33845 24344 33868
tri 24344 33845 24370 33871 sw
rect 24256 33822 24370 33845
rect 24141 33800 24370 33822
tri 24370 33800 24415 33845 sw
rect 70802 33820 71000 33878
tri 24141 33797 24144 33800 ne
rect 24144 33797 24415 33800
tri 24144 33758 24183 33797 ne
rect 24183 33790 24415 33797
tri 24415 33790 24425 33800 sw
rect 24183 33758 24425 33790
tri 24425 33758 24457 33790 sw
rect 70802 33774 70824 33820
rect 70870 33774 70928 33820
rect 70974 33774 71000 33820
tri 24183 33752 24189 33758 ne
rect 24189 33752 24457 33758
tri 24457 33752 24463 33758 sw
tri 24189 33707 24234 33752 ne
rect 24234 33736 24463 33752
rect 24234 33707 24342 33736
tri 24234 33681 24260 33707 ne
rect 24260 33690 24342 33707
rect 24388 33707 24463 33736
tri 24463 33707 24509 33752 sw
rect 70802 33716 71000 33774
rect 24388 33690 24509 33707
rect 24260 33681 24509 33690
tri 24260 33668 24273 33681 ne
rect 24273 33668 24509 33681
tri 24509 33668 24547 33707 sw
rect 70802 33670 70824 33716
rect 70870 33670 70928 33716
rect 70974 33670 71000 33716
tri 24273 33636 24305 33668 ne
rect 24305 33658 24547 33668
tri 24547 33658 24557 33668 sw
rect 24305 33636 24557 33658
tri 24305 33597 24344 33636 ne
rect 24344 33626 24557 33636
tri 24557 33626 24589 33658 sw
rect 24344 33613 24589 33626
tri 24589 33613 24602 33626 sw
rect 24344 33604 24602 33613
rect 24344 33597 24474 33604
tri 24344 33551 24389 33597 ne
rect 24389 33558 24474 33597
rect 24520 33597 24602 33604
tri 24602 33597 24619 33613 sw
rect 70802 33612 71000 33670
rect 24520 33581 24619 33597
tri 24619 33581 24634 33597 sw
rect 24520 33558 24634 33581
rect 24389 33551 24634 33558
tri 24389 33549 24392 33551 ne
rect 24392 33549 24634 33551
tri 24392 33536 24405 33549 ne
rect 24405 33536 24634 33549
tri 24634 33536 24679 33581 sw
rect 70802 33566 70824 33612
rect 70870 33566 70928 33612
rect 70974 33566 71000 33612
tri 24405 33504 24437 33536 ne
rect 24437 33526 24679 33536
tri 24679 33526 24689 33536 sw
rect 24437 33504 24689 33526
tri 24437 33494 24447 33504 ne
rect 24447 33494 24689 33504
tri 24689 33494 24721 33526 sw
rect 70802 33508 71000 33566
tri 24447 33449 24492 33494 ne
rect 24492 33481 24721 33494
tri 24721 33481 24734 33494 sw
rect 24492 33472 24734 33481
rect 24492 33449 24606 33472
tri 24492 33432 24509 33449 ne
rect 24509 33432 24606 33449
tri 24509 33404 24537 33432 ne
rect 24537 33426 24606 33432
rect 24652 33449 24734 33472
tri 24734 33449 24766 33481 sw
rect 70802 33462 70824 33508
rect 70870 33462 70928 33508
rect 70974 33462 71000 33508
rect 24652 33426 24766 33449
rect 24537 33404 24766 33426
tri 24766 33404 24811 33449 sw
rect 70802 33404 71000 33462
tri 24537 33372 24569 33404 ne
rect 24569 33394 24811 33404
tri 24811 33394 24821 33404 sw
rect 24569 33372 24821 33394
tri 24569 33327 24614 33372 ne
rect 24614 33362 24821 33372
tri 24821 33362 24853 33394 sw
rect 24614 33342 24853 33362
tri 24853 33342 24873 33362 sw
rect 70802 33358 70824 33404
rect 70870 33358 70928 33404
rect 70974 33358 71000 33404
rect 24614 33340 24873 33342
rect 24614 33327 24738 33340
tri 24614 33322 24619 33327 ne
rect 24619 33322 24738 33327
tri 24619 33285 24656 33322 ne
rect 24656 33294 24738 33322
rect 24784 33322 24873 33340
tri 24873 33322 24893 33342 sw
rect 24784 33317 24893 33322
tri 24893 33317 24898 33322 sw
rect 24784 33294 24898 33317
rect 24656 33285 24898 33294
tri 24656 33272 24669 33285 ne
rect 24669 33272 24898 33285
tri 24898 33272 24943 33317 sw
rect 70802 33300 71000 33358
tri 24669 33240 24701 33272 ne
rect 24701 33262 24943 33272
tri 24943 33262 24953 33272 sw
rect 24701 33240 24953 33262
tri 24701 33230 24711 33240 ne
rect 24711 33230 24953 33240
tri 24953 33230 24985 33262 sw
rect 70802 33254 70824 33300
rect 70870 33254 70928 33300
rect 70974 33254 71000 33300
tri 24711 33185 24756 33230 ne
rect 24756 33217 24985 33230
tri 24985 33217 24998 33230 sw
rect 24756 33208 24998 33217
rect 24756 33185 24870 33208
tri 24756 33153 24788 33185 ne
rect 24788 33162 24870 33185
rect 24916 33185 24998 33208
tri 24998 33185 25030 33217 sw
rect 70802 33196 71000 33254
rect 24916 33162 25030 33185
rect 24788 33153 25030 33162
tri 24788 33140 24801 33153 ne
rect 24801 33140 25030 33153
tri 25030 33140 25075 33185 sw
rect 70802 33150 70824 33196
rect 70870 33150 70928 33196
rect 70974 33150 71000 33196
tri 24801 33108 24833 33140 ne
rect 24833 33130 25075 33140
tri 25075 33130 25085 33140 sw
rect 24833 33108 25085 33130
tri 24833 33067 24873 33108 ne
rect 24873 33098 25085 33108
tri 25085 33098 25117 33130 sw
rect 24873 33085 25117 33098
tri 25117 33085 25130 33098 sw
rect 70802 33092 71000 33150
rect 24873 33076 25130 33085
rect 24873 33067 25002 33076
tri 24873 33048 24893 33067 ne
rect 24893 33048 25002 33067
tri 24893 33022 24919 33048 ne
rect 24919 33030 25002 33048
rect 25048 33048 25130 33076
tri 25130 33048 25167 33085 sw
rect 25048 33030 25167 33048
rect 24919 33022 25167 33030
tri 25167 33022 25193 33048 sw
rect 70802 33046 70824 33092
rect 70870 33046 70928 33092
rect 70974 33046 71000 33092
tri 24919 33021 24920 33022 ne
rect 24920 33021 25193 33022
tri 24920 33008 24933 33021 ne
rect 24933 33008 25193 33021
tri 25193 33008 25207 33022 sw
tri 24933 32976 24965 33008 ne
rect 24965 32998 25207 33008
tri 25207 32998 25217 33008 sw
rect 24965 32976 25217 32998
tri 24965 32966 24975 32976 ne
rect 24975 32966 25217 32976
tri 25217 32966 25249 32998 sw
rect 70802 32988 71000 33046
tri 24975 32921 25020 32966 ne
rect 25020 32953 25249 32966
tri 25249 32953 25262 32966 sw
rect 25020 32944 25262 32953
rect 25020 32921 25134 32944
tri 25020 32889 25052 32921 ne
rect 25052 32898 25134 32921
rect 25180 32921 25262 32944
tri 25262 32921 25294 32953 sw
rect 70802 32942 70824 32988
rect 70870 32942 70928 32988
rect 70974 32942 71000 32988
rect 25180 32898 25294 32921
rect 25052 32889 25294 32898
tri 25052 32876 25065 32889 ne
rect 25065 32876 25294 32889
tri 25294 32876 25339 32921 sw
rect 70802 32884 71000 32942
tri 25065 32844 25097 32876 ne
rect 25097 32866 25339 32876
tri 25339 32866 25349 32876 sw
rect 25097 32844 25349 32866
tri 25097 32799 25142 32844 ne
rect 25142 32834 25349 32844
tri 25349 32834 25381 32866 sw
rect 70802 32838 70824 32884
rect 70870 32838 70928 32884
rect 70974 32838 71000 32884
rect 25142 32821 25381 32834
tri 25381 32821 25394 32834 sw
rect 25142 32819 25394 32821
tri 25394 32819 25397 32821 sw
rect 25142 32812 25397 32819
rect 25142 32799 25266 32812
tri 25142 32773 25167 32799 ne
rect 25167 32773 25266 32799
tri 25167 32757 25184 32773 ne
rect 25184 32766 25266 32773
rect 25312 32773 25397 32812
tri 25397 32773 25442 32819 sw
rect 70802 32780 71000 32838
rect 25312 32766 25442 32773
rect 25184 32757 25442 32766
tri 25184 32744 25197 32757 ne
rect 25197 32744 25442 32757
tri 25442 32744 25471 32773 sw
tri 25197 32712 25229 32744 ne
rect 25229 32734 25471 32744
tri 25471 32734 25481 32744 sw
rect 70802 32734 70824 32780
rect 70870 32734 70928 32780
rect 70974 32734 71000 32780
rect 25229 32712 25481 32734
tri 25229 32703 25238 32712 ne
rect 25238 32703 25481 32712
tri 25238 32702 25239 32703 ne
rect 25239 32702 25481 32703
tri 25481 32702 25513 32734 sw
tri 25239 32657 25283 32702 ne
rect 25283 32689 25513 32702
tri 25513 32689 25526 32702 sw
rect 25283 32680 25526 32689
rect 25283 32657 25398 32680
tri 25283 32625 25316 32657 ne
rect 25316 32634 25398 32657
rect 25444 32657 25526 32680
tri 25526 32657 25558 32689 sw
rect 70802 32676 71000 32734
rect 25444 32634 25558 32657
rect 25316 32625 25558 32634
tri 25316 32612 25329 32625 ne
rect 25329 32612 25558 32625
tri 25558 32612 25603 32657 sw
rect 70802 32630 70824 32676
rect 70870 32630 70928 32676
rect 70974 32630 71000 32676
tri 25329 32580 25361 32612 ne
rect 25361 32602 25603 32612
tri 25603 32602 25613 32612 sw
rect 25361 32580 25613 32602
tri 25361 32535 25406 32580 ne
rect 25406 32570 25613 32580
tri 25613 32570 25645 32602 sw
rect 70802 32572 71000 32630
rect 25406 32557 25645 32570
tri 25645 32557 25658 32570 sw
rect 25406 32548 25658 32557
rect 25406 32535 25530 32548
tri 25406 32499 25442 32535 ne
rect 25442 32502 25530 32535
rect 25576 32544 25658 32548
tri 25658 32544 25671 32557 sw
rect 25576 32502 25671 32544
rect 25442 32499 25671 32502
tri 25671 32499 25716 32544 sw
rect 70802 32526 70824 32572
rect 70870 32526 70928 32572
rect 70974 32526 71000 32572
tri 25442 32493 25448 32499 ne
rect 25448 32493 25716 32499
tri 25448 32480 25461 32493 ne
rect 25461 32480 25716 32493
tri 25716 32480 25735 32499 sw
tri 25461 32448 25493 32480 ne
rect 25493 32470 25735 32480
tri 25735 32470 25745 32480 sw
rect 25493 32448 25745 32470
tri 25493 32438 25503 32448 ne
rect 25503 32438 25745 32448
tri 25745 32438 25777 32470 sw
rect 70802 32468 71000 32526
tri 25503 32393 25548 32438 ne
rect 25548 32425 25777 32438
tri 25777 32425 25790 32438 sw
rect 25548 32416 25790 32425
rect 25548 32393 25662 32416
tri 25548 32348 25593 32393 ne
rect 25593 32370 25662 32393
rect 25708 32393 25790 32416
tri 25790 32393 25822 32425 sw
rect 70802 32422 70824 32468
rect 70870 32422 70928 32468
rect 70974 32422 71000 32468
rect 25708 32370 25822 32393
rect 25593 32348 25822 32370
tri 25822 32348 25867 32393 sw
rect 70802 32364 71000 32422
tri 25593 32338 25603 32348 ne
rect 25603 32338 25867 32348
tri 25867 32338 25877 32348 sw
tri 25603 32293 25648 32338 ne
rect 25648 32306 25877 32338
tri 25877 32306 25909 32338 sw
rect 70802 32318 70824 32364
rect 70870 32318 70928 32364
rect 70974 32318 71000 32364
rect 25648 32293 25909 32306
tri 25909 32293 25922 32306 sw
tri 25648 32247 25693 32293 ne
rect 25693 32284 25923 32293
rect 25693 32247 25794 32284
tri 25693 32229 25712 32247 ne
rect 25712 32238 25794 32247
rect 25840 32247 25923 32284
tri 25923 32247 25968 32293 sw
rect 70802 32260 71000 32318
rect 25840 32238 25968 32247
rect 25712 32229 25968 32238
tri 25712 32225 25716 32229 ne
rect 25716 32225 25968 32229
tri 25968 32225 25991 32247 sw
tri 25716 32216 25725 32225 ne
rect 25725 32216 25991 32225
tri 25991 32216 25999 32225 sw
tri 25725 32184 25757 32216 ne
rect 25757 32206 25999 32216
tri 25999 32206 26009 32216 sw
rect 70802 32214 70824 32260
rect 70870 32214 70928 32260
rect 70974 32214 71000 32260
rect 25757 32184 26009 32206
tri 25757 32174 25767 32184 ne
rect 25767 32174 26009 32184
tri 26009 32174 26041 32206 sw
tri 25767 32129 25812 32174 ne
rect 25812 32161 26041 32174
tri 26041 32161 26054 32174 sw
rect 25812 32152 26054 32161
rect 25812 32129 25926 32152
tri 25812 32097 25844 32129 ne
rect 25844 32106 25926 32129
rect 25972 32129 26054 32152
tri 26054 32129 26086 32161 sw
rect 70802 32156 71000 32214
rect 25972 32106 26086 32129
rect 25844 32097 26086 32106
tri 25844 32084 25857 32097 ne
rect 25857 32084 26086 32097
tri 26086 32084 26131 32129 sw
rect 70802 32110 70824 32156
rect 70870 32110 70928 32156
rect 70974 32110 71000 32156
tri 25857 32052 25889 32084 ne
rect 25889 32074 26131 32084
tri 26131 32074 26141 32084 sw
rect 25889 32052 26141 32074
tri 25889 32007 25934 32052 ne
rect 25934 32042 26141 32052
tri 26141 32042 26173 32074 sw
rect 70802 32052 71000 32110
rect 25934 32029 26173 32042
tri 26173 32029 26186 32042 sw
rect 25934 32020 26186 32029
rect 25934 32007 26058 32020
tri 25934 31973 25968 32007 ne
rect 25968 31974 26058 32007
rect 26104 31997 26186 32020
tri 26186 31997 26218 32029 sw
rect 70802 32006 70824 32052
rect 70870 32006 70928 32052
rect 70974 32006 71000 32052
rect 26104 31974 26218 31997
rect 25968 31973 26218 31974
tri 25968 31950 25991 31973 ne
rect 25991 31952 26218 31973
tri 26218 31952 26263 31997 sw
rect 25991 31950 26263 31952
tri 26263 31950 26265 31952 sw
tri 25991 31920 26021 31950 ne
rect 26021 31942 26265 31950
tri 26265 31942 26273 31950 sw
rect 70802 31948 71000 32006
rect 26021 31920 26273 31942
tri 26021 31910 26031 31920 ne
rect 26031 31910 26273 31920
tri 26273 31910 26305 31942 sw
tri 26031 31865 26076 31910 ne
rect 26076 31888 26305 31910
rect 26076 31865 26190 31888
tri 26076 31833 26108 31865 ne
rect 26108 31842 26190 31865
rect 26236 31883 26305 31888
tri 26305 31883 26333 31910 sw
rect 70802 31902 70824 31948
rect 70870 31902 70928 31948
rect 70974 31902 71000 31948
rect 26236 31865 26333 31883
tri 26333 31865 26350 31883 sw
rect 26236 31842 26350 31865
rect 26108 31833 26350 31842
tri 26108 31820 26121 31833 ne
rect 26121 31820 26350 31833
tri 26350 31820 26395 31865 sw
rect 70802 31844 71000 31902
tri 26121 31788 26153 31820 ne
rect 26153 31810 26395 31820
tri 26395 31810 26405 31820 sw
rect 26153 31788 26405 31810
tri 26153 31743 26198 31788 ne
rect 26198 31778 26405 31788
tri 26405 31778 26437 31810 sw
rect 70802 31798 70824 31844
rect 70870 31798 70928 31844
rect 70974 31798 71000 31844
rect 26198 31765 26437 31778
tri 26437 31765 26450 31778 sw
rect 26198 31756 26450 31765
rect 26198 31743 26322 31756
tri 26198 31701 26240 31743 ne
rect 26240 31710 26322 31743
rect 26368 31733 26450 31756
tri 26450 31733 26482 31765 sw
rect 70802 31740 71000 31798
rect 26368 31710 26482 31733
rect 26240 31701 26482 31710
tri 26240 31676 26265 31701 ne
rect 26265 31688 26482 31701
tri 26482 31688 26527 31733 sw
rect 70802 31694 70824 31740
rect 70870 31694 70928 31740
rect 70974 31694 71000 31740
rect 26265 31678 26527 31688
tri 26527 31678 26537 31688 sw
rect 26265 31676 26537 31678
tri 26537 31676 26539 31678 sw
tri 26265 31656 26285 31676 ne
rect 26285 31656 26539 31676
tri 26285 31646 26295 31656 ne
rect 26295 31646 26539 31656
tri 26539 31646 26569 31676 sw
tri 26295 31608 26333 31646 ne
rect 26333 31633 26569 31646
tri 26569 31633 26582 31646 sw
rect 70802 31636 71000 31694
rect 26333 31624 26582 31633
rect 26333 31608 26454 31624
tri 26333 31563 26378 31608 ne
rect 26378 31578 26454 31608
rect 26500 31608 26582 31624
tri 26582 31608 26607 31633 sw
rect 26500 31578 26607 31608
rect 26378 31563 26607 31578
tri 26607 31563 26652 31608 sw
rect 70802 31590 70824 31636
rect 70870 31590 70928 31636
rect 70974 31590 71000 31636
tri 26378 31556 26385 31563 ne
rect 26385 31556 26652 31563
tri 26652 31556 26659 31563 sw
tri 26385 31524 26417 31556 ne
rect 26417 31546 26659 31556
tri 26659 31546 26669 31556 sw
rect 26417 31524 26669 31546
tri 26417 31479 26462 31524 ne
rect 26462 31514 26669 31524
tri 26669 31514 26701 31546 sw
rect 70802 31532 71000 31590
rect 26462 31501 26701 31514
tri 26701 31501 26714 31514 sw
rect 26462 31492 26714 31501
rect 26462 31479 26586 31492
tri 26462 31437 26504 31479 ne
rect 26504 31446 26586 31479
rect 26632 31469 26714 31492
tri 26714 31469 26746 31501 sw
rect 70802 31486 70824 31532
rect 70870 31486 70928 31532
rect 70974 31486 71000 31532
rect 26632 31446 26746 31469
rect 26504 31437 26746 31446
tri 26504 31401 26539 31437 ne
rect 26539 31424 26746 31437
tri 26746 31424 26791 31469 sw
rect 70802 31428 71000 31486
rect 26539 31414 26791 31424
tri 26791 31414 26801 31424 sw
rect 26539 31401 26801 31414
tri 26801 31401 26814 31414 sw
tri 26539 31392 26549 31401 ne
rect 26549 31392 26814 31401
tri 26549 31382 26559 31392 ne
rect 26559 31382 26814 31392
tri 26814 31382 26833 31401 sw
rect 70802 31382 70824 31428
rect 70870 31382 70928 31428
rect 70974 31382 71000 31428
tri 26559 31337 26604 31382 ne
rect 26604 31369 26833 31382
tri 26833 31369 26846 31382 sw
rect 26604 31360 26846 31369
rect 26604 31337 26718 31360
tri 26604 31305 26636 31337 ne
rect 26636 31314 26718 31337
rect 26764 31337 26846 31360
tri 26846 31337 26878 31369 sw
rect 26764 31314 26878 31337
rect 26636 31305 26878 31314
tri 26636 31292 26649 31305 ne
rect 26649 31292 26878 31305
tri 26878 31292 26923 31337 sw
rect 70802 31324 71000 31382
tri 26649 31260 26681 31292 ne
rect 26681 31282 26923 31292
tri 26923 31282 26933 31292 sw
rect 26681 31260 26933 31282
tri 26681 31243 26697 31260 ne
rect 26697 31250 26933 31260
tri 26933 31250 26965 31282 sw
rect 70802 31278 70824 31324
rect 70870 31278 70928 31324
rect 70974 31278 71000 31324
rect 26697 31243 26965 31250
tri 26697 31198 26743 31243 ne
rect 26743 31237 26965 31243
tri 26965 31237 26978 31250 sw
rect 26743 31228 26978 31237
rect 26743 31198 26850 31228
tri 26743 31173 26768 31198 ne
rect 26768 31182 26850 31198
rect 26896 31198 26978 31228
tri 26978 31198 27017 31237 sw
rect 70802 31220 71000 31278
rect 26896 31182 27017 31198
rect 26768 31173 27017 31182
tri 26768 31128 26813 31173 ne
rect 26813 31160 27017 31173
tri 27017 31160 27055 31198 sw
rect 70802 31174 70824 31220
rect 70870 31174 70928 31220
rect 70974 31174 71000 31220
rect 26813 31153 27055 31160
tri 27055 31153 27062 31160 sw
rect 26813 31150 27062 31153
tri 27062 31150 27065 31153 sw
rect 26813 31128 27065 31150
tri 26813 31127 26814 31128 ne
rect 26814 31127 27065 31128
tri 27065 31127 27088 31150 sw
tri 26814 31118 26823 31127 ne
rect 26823 31118 27088 31127
tri 27088 31118 27097 31127 sw
tri 26823 31073 26868 31118 ne
rect 26868 31105 27097 31118
tri 27097 31105 27110 31118 sw
rect 70802 31116 71000 31174
rect 26868 31096 27110 31105
rect 26868 31073 26982 31096
tri 26868 31041 26900 31073 ne
rect 26900 31050 26982 31073
rect 27028 31073 27110 31096
tri 27110 31073 27142 31105 sw
rect 27028 31050 27142 31073
rect 26900 31041 27142 31050
tri 26900 31028 26913 31041 ne
rect 26913 31028 27142 31041
tri 27142 31028 27187 31073 sw
rect 70802 31070 70824 31116
rect 70870 31070 70928 31116
rect 70974 31070 71000 31116
tri 26913 30996 26945 31028 ne
rect 26945 31018 27187 31028
tri 27187 31018 27197 31028 sw
rect 26945 30996 27197 31018
tri 26945 30951 26990 30996 ne
rect 26990 30986 27197 30996
tri 27197 30986 27229 31018 sw
rect 70802 31012 71000 31070
rect 26990 30973 27229 30986
tri 27229 30973 27242 30986 sw
rect 26990 30964 27242 30973
rect 26990 30951 27114 30964
tri 26990 30909 27032 30951 ne
rect 27032 30918 27114 30951
rect 27160 30941 27242 30964
tri 27242 30941 27274 30973 sw
rect 70802 30966 70824 31012
rect 70870 30966 70928 31012
rect 70974 30966 71000 31012
rect 27160 30918 27274 30941
rect 27032 30909 27274 30918
tri 27032 30864 27077 30909 ne
rect 27077 30896 27274 30909
tri 27274 30896 27319 30941 sw
rect 70802 30908 71000 30966
rect 27077 30886 27319 30896
tri 27319 30886 27329 30896 sw
rect 27077 30864 27329 30886
tri 27077 30853 27088 30864 ne
rect 27088 30854 27329 30864
tri 27329 30854 27361 30886 sw
rect 70802 30862 70824 30908
rect 70870 30862 70928 30908
rect 70974 30862 71000 30908
rect 27088 30853 27361 30854
tri 27361 30853 27363 30854 sw
tri 27088 30833 27107 30853 ne
rect 27107 30841 27363 30853
tri 27363 30841 27374 30853 sw
rect 27107 30833 27374 30841
tri 27374 30833 27382 30841 sw
tri 27107 30788 27153 30833 ne
rect 27153 30832 27382 30833
rect 27153 30788 27246 30832
tri 27153 30777 27164 30788 ne
rect 27164 30786 27246 30788
rect 27292 30788 27382 30832
tri 27382 30788 27427 30833 sw
rect 70802 30804 71000 30862
rect 27292 30786 27427 30788
rect 27164 30777 27427 30786
tri 27164 30764 27177 30777 ne
rect 27177 30764 27427 30777
tri 27427 30764 27451 30788 sw
tri 27177 30732 27209 30764 ne
rect 27209 30754 27451 30764
tri 27451 30754 27461 30764 sw
rect 70802 30758 70824 30804
rect 70870 30758 70928 30804
rect 70974 30758 71000 30804
rect 27209 30732 27461 30754
tri 27209 30722 27219 30732 ne
rect 27219 30722 27461 30732
tri 27461 30722 27493 30754 sw
tri 27219 30677 27264 30722 ne
rect 27264 30709 27493 30722
tri 27493 30709 27506 30722 sw
rect 27264 30700 27506 30709
rect 27264 30677 27378 30700
tri 27264 30645 27296 30677 ne
rect 27296 30654 27378 30677
rect 27424 30677 27506 30700
tri 27506 30677 27538 30709 sw
rect 70802 30700 71000 30758
rect 27424 30654 27538 30677
rect 27296 30645 27538 30654
tri 27296 30632 27309 30645 ne
rect 27309 30632 27538 30645
tri 27538 30632 27583 30677 sw
rect 70802 30654 70824 30700
rect 70870 30654 70928 30700
rect 70974 30654 71000 30700
tri 27309 30600 27341 30632 ne
rect 27341 30622 27583 30632
tri 27583 30622 27593 30632 sw
rect 27341 30600 27593 30622
tri 27341 30578 27363 30600 ne
rect 27363 30590 27593 30600
tri 27593 30590 27625 30622 sw
rect 70802 30596 71000 30654
rect 27363 30578 27625 30590
tri 27625 30578 27637 30590 sw
tri 27363 30533 27408 30578 ne
rect 27408 30577 27637 30578
tri 27637 30577 27638 30578 sw
rect 27408 30568 27638 30577
rect 27408 30533 27510 30568
tri 27408 30514 27427 30533 ne
rect 27427 30522 27510 30533
rect 27556 30545 27638 30568
tri 27638 30545 27670 30577 sw
rect 70802 30550 70824 30596
rect 70870 30550 70928 30596
rect 70974 30550 71000 30596
rect 27556 30522 27670 30545
rect 27427 30514 27670 30522
tri 27427 30500 27441 30514 ne
rect 27441 30500 27670 30514
tri 27670 30500 27715 30545 sw
tri 27441 30468 27473 30500 ne
rect 27473 30490 27715 30500
tri 27715 30490 27725 30500 sw
rect 70802 30492 71000 30550
rect 27473 30468 27725 30490
tri 27473 30458 27483 30468 ne
rect 27483 30458 27725 30468
tri 27725 30458 27757 30490 sw
tri 27483 30413 27528 30458 ne
rect 27528 30436 27757 30458
rect 27528 30413 27642 30436
tri 27528 30381 27560 30413 ne
rect 27560 30390 27642 30413
rect 27688 30423 27757 30436
tri 27757 30423 27792 30458 sw
rect 70802 30446 70824 30492
rect 70870 30446 70928 30492
rect 70974 30446 71000 30492
rect 27688 30413 27792 30423
tri 27792 30413 27802 30423 sw
rect 27688 30390 27802 30413
rect 27560 30381 27802 30390
tri 27560 30368 27573 30381 ne
rect 27573 30368 27802 30381
tri 27802 30368 27847 30413 sw
rect 70802 30388 71000 30446
tri 27573 30336 27605 30368 ne
rect 27605 30358 27847 30368
tri 27847 30358 27857 30368 sw
rect 27605 30336 27857 30358
tri 27605 30304 27637 30336 ne
rect 27637 30326 27857 30336
tri 27857 30326 27889 30358 sw
rect 70802 30342 70824 30388
rect 70870 30342 70928 30388
rect 70974 30342 71000 30388
rect 27637 30313 27889 30326
tri 27889 30313 27902 30326 sw
rect 27637 30304 27902 30313
tri 27902 30304 27911 30313 sw
tri 27637 30259 27682 30304 ne
rect 27682 30259 27774 30304
tri 27682 30249 27692 30259 ne
rect 27692 30258 27774 30259
rect 27820 30281 27911 30304
tri 27911 30281 27934 30304 sw
rect 70802 30284 71000 30342
rect 27820 30258 27934 30281
rect 27692 30249 27934 30258
tri 27692 30236 27705 30249 ne
rect 27705 30236 27934 30249
tri 27934 30236 27979 30281 sw
rect 70802 30238 70824 30284
rect 70870 30238 70928 30284
rect 70974 30238 71000 30284
tri 27705 30204 27737 30236 ne
rect 27737 30226 27979 30236
tri 27979 30226 27989 30236 sw
rect 27737 30204 27989 30226
tri 27737 30194 27747 30204 ne
rect 27747 30194 27989 30204
tri 27989 30194 28021 30226 sw
tri 27747 30149 27792 30194 ne
rect 27792 30181 28021 30194
tri 28021 30181 28034 30194 sw
rect 27792 30172 28034 30181
rect 27792 30149 27906 30172
tri 27792 30104 27837 30149 ne
rect 27837 30126 27906 30149
rect 27952 30149 28034 30172
tri 28034 30149 28066 30181 sw
rect 70802 30180 71000 30238
rect 27952 30126 28066 30149
rect 27837 30104 28066 30126
tri 28066 30104 28111 30149 sw
rect 70802 30134 70824 30180
rect 70870 30134 70928 30180
rect 70974 30134 71000 30180
tri 27837 30072 27869 30104 ne
rect 27869 30072 28111 30104
tri 27869 30029 27911 30072 ne
rect 27911 30062 28111 30072
tri 28111 30062 28153 30104 sw
rect 70802 30076 71000 30134
rect 27911 30049 28153 30062
tri 28153 30049 28166 30062 sw
rect 27911 30040 28166 30049
rect 27911 30029 28038 30040
tri 27911 29985 27956 30029 ne
rect 27956 29994 28038 30029
rect 28084 30029 28166 30040
tri 28166 30029 28186 30049 sw
rect 70802 30030 70824 30076
rect 70870 30030 70928 30076
rect 70974 30030 71000 30076
rect 28084 30017 28186 30029
tri 28186 30017 28198 30029 sw
rect 28084 29994 28198 30017
rect 27956 29985 28198 29994
tri 27956 29972 27969 29985 ne
rect 27969 29972 28198 29985
tri 28198 29972 28243 30017 sw
rect 70802 29972 71000 30030
tri 27969 29940 28001 29972 ne
rect 28001 29962 28243 29972
tri 28243 29962 28253 29972 sw
rect 28001 29940 28253 29962
tri 28001 29930 28011 29940 ne
rect 28011 29930 28253 29940
tri 28253 29930 28285 29962 sw
tri 28011 29885 28056 29930 ne
rect 28056 29917 28285 29930
tri 28285 29917 28298 29930 sw
rect 70802 29926 70824 29972
rect 70870 29926 70928 29972
rect 70974 29926 71000 29972
rect 28056 29908 28298 29917
rect 28056 29885 28170 29908
tri 28056 29853 28088 29885 ne
rect 28088 29862 28170 29885
rect 28216 29885 28298 29908
tri 28298 29885 28330 29917 sw
rect 28216 29862 28330 29885
rect 28088 29853 28330 29862
tri 28088 29840 28101 29853 ne
rect 28101 29840 28330 29853
tri 28330 29840 28375 29885 sw
rect 70802 29868 71000 29926
tri 28101 29808 28133 29840 ne
rect 28133 29830 28375 29840
tri 28375 29830 28385 29840 sw
rect 28133 29808 28385 29830
tri 28133 29784 28157 29808 ne
rect 28157 29798 28385 29808
tri 28385 29798 28417 29830 sw
rect 70802 29822 70824 29868
rect 70870 29822 70928 29868
rect 70974 29822 71000 29868
rect 28157 29785 28417 29798
tri 28417 29785 28430 29798 sw
rect 28157 29784 28430 29785
tri 28157 29755 28186 29784 ne
rect 28186 29776 28430 29784
rect 28186 29755 28302 29776
tri 28186 29739 28202 29755 ne
rect 28202 29739 28302 29755
tri 28202 29721 28220 29739 ne
rect 28220 29730 28302 29739
rect 28348 29755 28430 29776
tri 28430 29755 28460 29785 sw
rect 70802 29764 71000 29822
rect 28348 29739 28460 29755
tri 28460 29739 28476 29755 sw
rect 28348 29730 28476 29739
rect 28220 29721 28476 29730
tri 28220 29708 28233 29721 ne
rect 28233 29708 28476 29721
tri 28476 29708 28507 29739 sw
rect 70802 29718 70824 29764
rect 70870 29718 70928 29764
rect 70974 29718 71000 29764
tri 28233 29676 28265 29708 ne
rect 28265 29698 28507 29708
tri 28507 29698 28517 29708 sw
rect 28265 29676 28517 29698
tri 28265 29666 28275 29676 ne
rect 28275 29666 28517 29676
tri 28517 29666 28549 29698 sw
tri 28275 29621 28320 29666 ne
rect 28320 29653 28549 29666
tri 28549 29653 28562 29666 sw
rect 70802 29660 71000 29718
rect 28320 29644 28562 29653
rect 28320 29621 28434 29644
tri 28320 29589 28352 29621 ne
rect 28352 29598 28434 29621
rect 28480 29621 28562 29644
tri 28562 29621 28594 29653 sw
rect 28480 29598 28594 29621
rect 28352 29589 28594 29598
tri 28352 29576 28365 29589 ne
rect 28365 29576 28594 29589
tri 28594 29576 28639 29621 sw
rect 70802 29614 70824 29660
rect 70870 29614 70928 29660
rect 70974 29614 71000 29660
tri 28365 29544 28397 29576 ne
rect 28397 29566 28639 29576
tri 28639 29566 28649 29576 sw
rect 28397 29544 28649 29566
tri 28397 29499 28442 29544 ne
rect 28442 29534 28649 29544
tri 28649 29534 28681 29566 sw
rect 70802 29556 71000 29614
rect 28442 29521 28681 29534
tri 28681 29521 28694 29534 sw
rect 28442 29512 28694 29521
rect 28442 29499 28566 29512
tri 28442 29481 28460 29499 ne
rect 28460 29481 28566 29499
tri 28460 29457 28484 29481 ne
rect 28484 29466 28566 29481
rect 28612 29481 28694 29512
tri 28694 29481 28735 29521 sw
rect 70802 29510 70824 29556
rect 70870 29510 70928 29556
rect 70974 29510 71000 29556
rect 28612 29466 28735 29481
rect 28484 29457 28735 29466
tri 28484 29444 28497 29457 ne
rect 28497 29444 28735 29457
tri 28735 29444 28771 29481 sw
rect 70802 29452 71000 29510
tri 28497 29412 28529 29444 ne
rect 28529 29434 28771 29444
tri 28771 29434 28781 29444 sw
rect 28529 29412 28781 29434
tri 28529 29402 28539 29412 ne
rect 28539 29402 28781 29412
tri 28781 29402 28813 29434 sw
rect 70802 29406 70824 29452
rect 70870 29406 70928 29452
rect 70974 29406 71000 29452
tri 28539 29374 28567 29402 ne
rect 28567 29389 28813 29402
tri 28813 29389 28826 29402 sw
rect 28567 29380 28826 29389
rect 28567 29374 28698 29380
tri 28567 29329 28612 29374 ne
rect 28612 29334 28698 29374
rect 28744 29374 28826 29380
tri 28826 29374 28841 29389 sw
rect 28744 29334 28841 29374
rect 28612 29329 28841 29334
tri 28841 29329 28886 29374 sw
rect 70802 29348 71000 29406
tri 28612 29325 28616 29329 ne
rect 28616 29325 28886 29329
tri 28616 29312 28629 29325 ne
rect 28629 29312 28886 29325
tri 28886 29312 28903 29329 sw
tri 28629 29280 28661 29312 ne
rect 28661 29302 28903 29312
tri 28903 29302 28913 29312 sw
rect 70802 29302 70824 29348
rect 70870 29302 70928 29348
rect 70974 29302 71000 29348
rect 28661 29280 28913 29302
tri 28661 29235 28706 29280 ne
rect 28706 29270 28913 29280
tri 28913 29270 28945 29302 sw
rect 28706 29257 28945 29270
tri 28945 29257 28958 29270 sw
rect 28706 29251 28958 29257
tri 28958 29251 28964 29257 sw
rect 28706 29248 28964 29251
rect 28706 29235 28830 29248
tri 28706 29206 28735 29235 ne
rect 28735 29206 28830 29235
tri 28735 29193 28748 29206 ne
rect 28748 29202 28830 29206
rect 28876 29206 28964 29248
tri 28964 29206 29009 29251 sw
rect 70802 29244 71000 29302
rect 28876 29202 29009 29206
rect 28748 29193 29009 29202
tri 28748 29180 28761 29193 ne
rect 28761 29180 29009 29193
tri 29009 29180 29035 29206 sw
rect 70802 29198 70824 29244
rect 70870 29198 70928 29244
rect 70974 29198 71000 29244
tri 28761 29148 28793 29180 ne
rect 28793 29170 29035 29180
tri 29035 29170 29045 29180 sw
rect 28793 29148 29045 29170
tri 28793 29138 28803 29148 ne
rect 28803 29138 29045 29148
tri 29045 29138 29077 29170 sw
rect 70802 29140 71000 29198
tri 28803 29093 28848 29138 ne
rect 28848 29125 29077 29138
tri 29077 29125 29090 29138 sw
rect 28848 29116 29090 29125
rect 28848 29093 28962 29116
tri 28848 29055 28886 29093 ne
rect 28886 29070 28962 29093
rect 29008 29093 29090 29116
tri 29090 29093 29122 29125 sw
rect 70802 29094 70824 29140
rect 70870 29094 70928 29140
rect 70974 29094 71000 29140
rect 29008 29070 29122 29093
rect 28886 29055 29122 29070
tri 28886 29048 28893 29055 ne
rect 28893 29048 29122 29055
tri 29122 29048 29167 29093 sw
tri 28893 29009 28931 29048 ne
rect 28931 29038 29167 29048
tri 29167 29038 29177 29048 sw
rect 28931 29009 29177 29038
tri 28931 28964 28977 29009 ne
rect 28977 29006 29177 29009
tri 29177 29006 29209 29038 sw
rect 70802 29036 71000 29094
rect 28977 28984 29209 29006
rect 28977 28964 29094 28984
tri 28977 28932 29009 28964 ne
rect 29009 28938 29094 28964
rect 29140 28964 29209 28984
tri 29209 28964 29251 29006 sw
rect 70802 28990 70824 29036
rect 70870 28990 70928 29036
rect 70974 28990 71000 29036
rect 29140 28938 29251 28964
rect 29009 28932 29251 28938
tri 29251 28932 29283 28964 sw
rect 70802 28932 71000 28990
tri 29009 28929 29012 28932 ne
rect 29012 28929 29283 28932
tri 29012 28916 29025 28929 ne
rect 29025 28916 29283 28929
tri 29283 28916 29299 28932 sw
tri 29025 28884 29057 28916 ne
rect 29057 28906 29299 28916
tri 29299 28906 29309 28916 sw
rect 29057 28884 29309 28906
tri 29057 28874 29067 28884 ne
rect 29067 28874 29309 28884
tri 29309 28874 29341 28906 sw
rect 70802 28886 70824 28932
rect 70870 28886 70928 28932
rect 70974 28886 71000 28932
tri 29067 28829 29112 28874 ne
rect 29112 28861 29341 28874
tri 29341 28861 29354 28874 sw
rect 29112 28852 29354 28861
rect 29112 28829 29226 28852
tri 29112 28797 29144 28829 ne
rect 29144 28806 29226 28829
rect 29272 28829 29354 28852
tri 29354 28829 29386 28861 sw
rect 29272 28806 29386 28829
rect 29144 28797 29386 28806
tri 29144 28784 29157 28797 ne
rect 29157 28784 29386 28797
tri 29386 28784 29431 28829 sw
rect 70802 28828 71000 28886
tri 29157 28752 29189 28784 ne
rect 29189 28774 29431 28784
tri 29431 28774 29441 28784 sw
rect 70802 28782 70824 28828
rect 70870 28782 70928 28828
rect 70974 28782 71000 28828
rect 29189 28752 29441 28774
tri 29189 28707 29234 28752 ne
rect 29234 28742 29441 28752
tri 29441 28742 29473 28774 sw
rect 29234 28729 29473 28742
tri 29473 28729 29486 28742 sw
rect 29234 28720 29486 28729
rect 29234 28707 29358 28720
tri 29234 28690 29251 28707 ne
rect 29251 28690 29358 28707
tri 29251 28657 29283 28690 ne
rect 29283 28674 29358 28690
rect 29404 28703 29486 28720
tri 29486 28703 29513 28729 sw
rect 70802 28724 71000 28782
rect 29404 28674 29513 28703
rect 29283 28657 29513 28674
tri 29513 28657 29558 28703 sw
rect 70802 28678 70824 28724
rect 70870 28678 70928 28724
rect 70974 28678 71000 28724
tri 29283 28652 29289 28657 ne
rect 29289 28652 29558 28657
tri 29558 28652 29563 28657 sw
tri 29289 28620 29321 28652 ne
rect 29321 28645 29563 28652
tri 29563 28645 29571 28652 sw
rect 29321 28620 29571 28645
tri 29321 28610 29331 28620 ne
rect 29331 28610 29571 28620
tri 29571 28610 29605 28645 sw
rect 70802 28620 71000 28678
tri 29331 28565 29376 28610 ne
rect 29376 28597 29605 28610
tri 29605 28597 29618 28610 sw
rect 29376 28588 29618 28597
rect 29376 28565 29490 28588
tri 29376 28533 29408 28565 ne
rect 29408 28542 29490 28565
rect 29536 28565 29618 28588
tri 29618 28565 29650 28597 sw
rect 70802 28574 70824 28620
rect 70870 28574 70928 28620
rect 70974 28574 71000 28620
rect 29536 28542 29650 28565
rect 29408 28533 29650 28542
tri 29408 28520 29421 28533 ne
rect 29421 28520 29650 28533
tri 29650 28520 29695 28565 sw
tri 29421 28488 29453 28520 ne
rect 29453 28510 29695 28520
tri 29695 28510 29705 28520 sw
rect 70802 28516 71000 28574
rect 29453 28488 29705 28510
tri 29453 28443 29498 28488 ne
rect 29498 28478 29705 28488
tri 29705 28478 29737 28510 sw
rect 29498 28465 29737 28478
tri 29737 28465 29750 28478 sw
rect 70802 28470 70824 28516
rect 70870 28470 70928 28516
rect 70974 28470 71000 28516
rect 29498 28456 29750 28465
rect 29498 28443 29622 28456
tri 29498 28401 29540 28443 ne
rect 29540 28410 29622 28443
rect 29668 28433 29750 28456
tri 29750 28433 29782 28465 sw
rect 29668 28410 29782 28433
rect 29540 28401 29782 28410
tri 29540 28383 29558 28401 ne
rect 29558 28388 29782 28401
tri 29782 28388 29827 28433 sw
rect 70802 28412 71000 28470
rect 29558 28383 29827 28388
tri 29827 28383 29832 28388 sw
tri 29558 28356 29585 28383 ne
rect 29585 28378 29832 28383
tri 29832 28378 29837 28383 sw
rect 29585 28356 29837 28378
tri 29585 28346 29595 28356 ne
rect 29595 28346 29837 28356
tri 29837 28346 29869 28378 sw
rect 70802 28366 70824 28412
rect 70870 28366 70928 28412
rect 70974 28366 71000 28412
tri 29595 28325 29616 28346 ne
rect 29616 28333 29869 28346
tri 29869 28333 29882 28346 sw
rect 29616 28325 29882 28333
tri 29882 28325 29890 28333 sw
tri 29616 28280 29661 28325 ne
rect 29661 28324 29890 28325
rect 29661 28280 29754 28324
tri 29661 28269 29672 28280 ne
rect 29672 28278 29754 28280
rect 29800 28280 29890 28324
tri 29890 28280 29935 28325 sw
rect 70802 28308 71000 28366
rect 29800 28278 29935 28280
rect 29672 28269 29935 28278
tri 29672 28256 29685 28269 ne
rect 29685 28256 29935 28269
tri 29935 28256 29959 28280 sw
rect 70802 28262 70824 28308
rect 70870 28262 70928 28308
rect 70974 28262 71000 28308
tri 29685 28224 29717 28256 ne
rect 29717 28246 29959 28256
tri 29959 28246 29969 28256 sw
rect 29717 28224 29969 28246
tri 29717 28179 29762 28224 ne
rect 29762 28214 29969 28224
tri 29969 28214 30001 28246 sw
rect 29762 28201 30001 28214
tri 30001 28201 30014 28214 sw
rect 70802 28204 71000 28262
rect 29762 28192 30014 28201
rect 29762 28179 29886 28192
tri 29762 28137 29804 28179 ne
rect 29804 28146 29886 28179
rect 29932 28169 30014 28192
tri 30014 28169 30046 28201 sw
rect 29932 28146 30046 28169
rect 29804 28137 30046 28146
tri 29804 28109 29832 28137 ne
rect 29832 28124 30046 28137
tri 30046 28124 30091 28169 sw
rect 70802 28158 70824 28204
rect 70870 28158 70928 28204
rect 70974 28158 71000 28204
rect 29832 28114 30091 28124
tri 30091 28114 30101 28124 sw
rect 29832 28109 30101 28114
tri 30101 28109 30107 28114 sw
tri 29832 28092 29849 28109 ne
rect 29849 28092 30107 28109
tri 29849 28082 29859 28092 ne
rect 29859 28082 30107 28092
tri 30107 28082 30133 28109 sw
rect 70802 28100 71000 28158
tri 29859 28037 29904 28082 ne
rect 29904 28069 30133 28082
tri 30133 28069 30146 28082 sw
rect 29904 28060 30146 28069
rect 29904 28037 30018 28060
tri 29904 28005 29936 28037 ne
rect 29936 28014 30018 28037
rect 30064 28037 30146 28060
tri 30146 28037 30178 28069 sw
rect 70802 28054 70824 28100
rect 70870 28054 70928 28100
rect 70974 28054 71000 28100
rect 30064 28014 30178 28037
rect 29936 28005 30178 28014
tri 29936 27992 29949 28005 ne
rect 29949 27992 30178 28005
tri 30178 27992 30223 28037 sw
rect 70802 27996 71000 28054
tri 29949 27960 29981 27992 ne
rect 29981 27982 30223 27992
tri 30223 27982 30233 27992 sw
rect 29981 27960 30233 27982
tri 29981 27915 30026 27960 ne
rect 30026 27950 30233 27960
tri 30233 27950 30265 27982 sw
rect 70802 27950 70824 27996
rect 70870 27950 70928 27996
rect 70974 27950 71000 27996
rect 30026 27937 30265 27950
tri 30265 27937 30278 27950 sw
rect 30026 27928 30278 27937
rect 30026 27915 30150 27928
tri 30026 27873 30068 27915 ne
rect 30068 27882 30150 27915
rect 30196 27915 30278 27928
tri 30278 27915 30300 27937 sw
rect 30196 27882 30300 27915
rect 30068 27873 30300 27882
tri 30068 27834 30107 27873 ne
rect 30107 27870 30300 27873
tri 30300 27870 30345 27915 sw
rect 70802 27892 71000 27950
rect 30107 27860 30345 27870
tri 30345 27860 30355 27870 sw
rect 30107 27850 30355 27860
tri 30355 27850 30365 27860 sw
rect 30107 27834 30365 27850
tri 30365 27834 30381 27850 sw
rect 70802 27846 70824 27892
rect 70870 27846 70928 27892
rect 70974 27846 71000 27892
tri 30107 27828 30113 27834 ne
rect 30113 27828 30381 27834
tri 30113 27818 30123 27828 ne
rect 30123 27818 30381 27828
tri 30381 27818 30397 27834 sw
tri 30123 27773 30168 27818 ne
rect 30168 27805 30397 27818
tri 30397 27805 30410 27818 sw
rect 30168 27796 30410 27805
rect 30168 27773 30282 27796
tri 30168 27741 30200 27773 ne
rect 30200 27750 30282 27773
rect 30328 27773 30410 27796
tri 30410 27773 30442 27805 sw
rect 70802 27788 71000 27846
rect 30328 27750 30442 27773
rect 30200 27741 30442 27750
tri 30200 27728 30213 27741 ne
rect 30213 27728 30442 27741
tri 30442 27728 30487 27773 sw
rect 70802 27742 70824 27788
rect 70870 27742 70928 27788
rect 70974 27742 71000 27788
tri 30213 27696 30245 27728 ne
rect 30245 27718 30487 27728
tri 30487 27718 30497 27728 sw
rect 30245 27696 30497 27718
tri 30245 27651 30290 27696 ne
rect 30290 27686 30497 27696
tri 30497 27686 30529 27718 sw
rect 30290 27673 30529 27686
tri 30529 27673 30542 27686 sw
rect 70802 27684 71000 27742
rect 30290 27664 30542 27673
rect 30290 27651 30414 27664
tri 30290 27641 30300 27651 ne
rect 30300 27641 30414 27651
tri 30300 27595 30345 27641 ne
rect 30345 27618 30414 27641
rect 30460 27641 30542 27664
tri 30542 27641 30574 27673 sw
rect 30460 27618 30574 27641
rect 30345 27596 30574 27618
tri 30574 27596 30619 27641 sw
rect 70802 27638 70824 27684
rect 70870 27638 70928 27684
rect 70974 27638 71000 27684
rect 30345 27595 30619 27596
tri 30345 27560 30381 27595 ne
rect 30381 27586 30619 27595
tri 30619 27586 30629 27596 sw
rect 30381 27560 30629 27586
tri 30629 27560 30655 27586 sw
rect 70802 27580 71000 27638
tri 30381 27554 30387 27560 ne
rect 30387 27554 30655 27560
tri 30655 27554 30661 27560 sw
tri 30387 27550 30391 27554 ne
rect 30391 27550 30661 27554
tri 30661 27550 30665 27554 sw
tri 30391 27505 30436 27550 ne
rect 30436 27532 30665 27550
rect 30436 27505 30546 27532
tri 30436 27477 30464 27505 ne
rect 30464 27486 30546 27505
rect 30592 27505 30665 27532
tri 30665 27505 30710 27550 sw
rect 70802 27534 70824 27580
rect 70870 27534 70928 27580
rect 70974 27534 71000 27580
rect 30592 27486 30710 27505
rect 30464 27477 30710 27486
tri 30464 27464 30477 27477 ne
rect 30477 27464 30710 27477
tri 30710 27464 30751 27505 sw
rect 70802 27476 71000 27534
tri 30477 27432 30509 27464 ne
rect 30509 27454 30751 27464
tri 30751 27454 30761 27464 sw
rect 30509 27432 30761 27454
tri 30509 27387 30554 27432 ne
rect 30554 27422 30761 27432
tri 30761 27422 30793 27454 sw
rect 70802 27430 70824 27476
rect 70870 27430 70928 27476
rect 70974 27430 71000 27476
rect 30554 27409 30793 27422
tri 30793 27409 30806 27422 sw
rect 30554 27400 30806 27409
rect 30554 27387 30678 27400
tri 30554 27345 30596 27387 ne
rect 30596 27354 30678 27387
rect 30724 27377 30806 27400
tri 30806 27377 30838 27409 sw
rect 30724 27354 30838 27377
rect 30596 27345 30838 27354
tri 30596 27300 30641 27345 ne
rect 30641 27332 30838 27345
tri 30838 27332 30883 27377 sw
rect 70802 27372 71000 27430
rect 30641 27322 30883 27332
tri 30883 27322 30893 27332 sw
rect 70802 27326 70824 27372
rect 70870 27326 70928 27372
rect 70974 27326 71000 27372
rect 30641 27300 30893 27322
tri 30641 27285 30655 27300 ne
rect 30655 27290 30893 27300
tri 30893 27290 30925 27322 sw
rect 30655 27285 30925 27290
tri 30925 27285 30930 27290 sw
tri 30655 27240 30701 27285 ne
rect 30701 27277 30930 27285
tri 30930 27277 30938 27285 sw
rect 30701 27268 30938 27277
rect 30701 27240 30810 27268
tri 30701 27231 30710 27240 ne
rect 30710 27231 30810 27240
tri 30710 27200 30741 27231 ne
rect 30741 27222 30810 27231
rect 30856 27245 30938 27268
tri 30938 27245 30970 27277 sw
rect 70802 27268 71000 27326
rect 30856 27222 30970 27245
rect 30741 27200 30970 27222
tri 30970 27200 31015 27245 sw
rect 70802 27222 70824 27268
rect 70870 27222 70928 27268
rect 70974 27222 71000 27268
tri 30741 27168 30773 27200 ne
rect 30773 27190 31015 27200
tri 31015 27190 31025 27200 sw
rect 30773 27168 31025 27190
tri 30773 27158 30783 27168 ne
rect 30783 27158 31025 27168
tri 31025 27158 31057 27190 sw
rect 70802 27164 71000 27222
tri 30783 27113 30828 27158 ne
rect 30828 27140 31057 27158
tri 31057 27140 31075 27158 sw
rect 30828 27136 31075 27140
rect 30828 27113 30942 27136
tri 30828 27081 30860 27113 ne
rect 30860 27090 30942 27113
rect 30988 27113 31075 27136
tri 31075 27113 31102 27140 sw
rect 70802 27118 70824 27164
rect 70870 27118 70928 27164
rect 70974 27118 71000 27164
rect 30988 27090 31102 27113
rect 30860 27081 31102 27090
tri 30860 27068 30873 27081 ne
rect 30873 27068 31102 27081
tri 31102 27068 31147 27113 sw
tri 30873 27036 30905 27068 ne
rect 30905 27058 31147 27068
tri 31147 27058 31157 27068 sw
rect 70802 27060 71000 27118
rect 30905 27036 31157 27058
tri 30905 27011 30930 27036 ne
rect 30930 27026 31157 27036
tri 31157 27026 31189 27058 sw
rect 30930 27013 31189 27026
tri 31189 27013 31202 27026 sw
rect 70802 27014 70824 27060
rect 70870 27014 70928 27060
rect 70974 27014 71000 27060
rect 30930 27011 31202 27013
tri 31202 27011 31204 27013 sw
tri 30930 26966 30975 27011 ne
rect 30975 27004 31204 27011
rect 30975 26966 31074 27004
tri 30975 26949 30992 26966 ne
rect 30992 26958 31074 26966
rect 31120 26981 31204 27004
tri 31204 26981 31234 27011 sw
rect 31120 26958 31234 26981
rect 30992 26949 31234 26958
tri 30992 26936 31005 26949 ne
rect 31005 26936 31234 26949
tri 31234 26936 31279 26981 sw
rect 70802 26956 71000 27014
tri 31005 26904 31037 26936 ne
rect 31037 26926 31279 26936
tri 31279 26926 31289 26936 sw
rect 31037 26904 31289 26926
tri 31037 26894 31047 26904 ne
rect 31047 26894 31289 26904
tri 31289 26894 31321 26926 sw
rect 70802 26910 70824 26956
rect 70870 26910 70928 26956
rect 70974 26910 71000 26956
tri 31047 26866 31075 26894 ne
rect 31075 26881 31321 26894
tri 31321 26881 31334 26894 sw
rect 31075 26872 31334 26881
rect 31075 26866 31206 26872
tri 31075 26821 31120 26866 ne
rect 31120 26826 31206 26866
rect 31252 26866 31334 26872
tri 31334 26866 31349 26881 sw
rect 31252 26826 31349 26866
rect 31120 26821 31349 26826
tri 31349 26821 31395 26866 sw
rect 70802 26852 71000 26910
tri 31120 26817 31124 26821 ne
rect 31124 26817 31395 26821
tri 31124 26804 31137 26817 ne
rect 31137 26804 31395 26817
tri 31395 26804 31411 26821 sw
rect 70802 26806 70824 26852
rect 70870 26806 70928 26852
rect 70974 26806 71000 26852
tri 31137 26772 31169 26804 ne
rect 31169 26794 31411 26804
tri 31411 26794 31421 26804 sw
rect 31169 26772 31421 26794
tri 31169 26737 31204 26772 ne
rect 31204 26762 31421 26772
tri 31421 26762 31453 26794 sw
rect 31204 26749 31453 26762
tri 31453 26749 31466 26762 sw
rect 31204 26740 31466 26749
rect 31204 26737 31338 26740
tri 31204 26691 31249 26737 ne
rect 31249 26694 31338 26737
rect 31384 26737 31466 26740
tri 31466 26737 31479 26749 sw
rect 70802 26748 71000 26806
rect 31384 26717 31479 26737
tri 31479 26717 31498 26737 sw
rect 31384 26694 31498 26717
rect 31249 26691 31498 26694
tri 31249 26685 31256 26691 ne
rect 31256 26685 31498 26691
tri 31256 26672 31269 26685 ne
rect 31269 26672 31498 26685
tri 31498 26672 31543 26717 sw
rect 70802 26702 70824 26748
rect 70870 26702 70928 26748
rect 70974 26702 71000 26748
tri 31269 26640 31301 26672 ne
rect 31301 26662 31543 26672
tri 31543 26662 31553 26672 sw
rect 31301 26640 31553 26662
tri 31301 26630 31311 26640 ne
rect 31311 26630 31553 26640
tri 31553 26630 31585 26662 sw
rect 70802 26644 71000 26702
tri 31311 26585 31356 26630 ne
rect 31356 26617 31585 26630
tri 31585 26617 31598 26630 sw
rect 31356 26608 31598 26617
rect 31356 26585 31470 26608
tri 31356 26553 31388 26585 ne
rect 31388 26562 31470 26585
rect 31516 26585 31598 26608
tri 31598 26585 31630 26617 sw
rect 70802 26598 70824 26644
rect 70870 26598 70928 26644
rect 70974 26598 71000 26644
rect 31516 26562 31630 26585
rect 31388 26553 31630 26562
tri 31388 26540 31401 26553 ne
rect 31401 26540 31630 26553
tri 31630 26540 31675 26585 sw
rect 70802 26540 71000 26598
tri 31401 26508 31433 26540 ne
rect 31433 26530 31675 26540
tri 31675 26530 31685 26540 sw
rect 31433 26508 31685 26530
tri 31433 26501 31440 26508 ne
rect 31440 26501 31685 26508
tri 31440 26462 31479 26501 ne
rect 31479 26498 31685 26501
tri 31685 26498 31717 26530 sw
rect 31479 26485 31717 26498
tri 31717 26485 31730 26498 sw
rect 70802 26494 70824 26540
rect 70870 26494 70928 26540
rect 70974 26494 71000 26540
rect 31479 26476 31730 26485
rect 31479 26462 31602 26476
tri 31479 26456 31485 26462 ne
rect 31485 26456 31602 26462
tri 31485 26421 31520 26456 ne
rect 31520 26430 31602 26456
rect 31648 26462 31730 26476
tri 31730 26462 31753 26485 sw
rect 31648 26456 31753 26462
tri 31753 26456 31759 26462 sw
rect 31648 26430 31759 26456
rect 31520 26421 31759 26430
tri 31520 26408 31533 26421 ne
rect 31533 26411 31759 26421
tri 31759 26411 31805 26456 sw
rect 70802 26436 71000 26494
rect 31533 26408 31805 26411
tri 31805 26408 31807 26411 sw
tri 31533 26376 31565 26408 ne
rect 31565 26398 31807 26408
tri 31807 26398 31817 26408 sw
rect 31565 26376 31817 26398
tri 31565 26366 31575 26376 ne
rect 31575 26366 31817 26376
tri 31817 26366 31849 26398 sw
rect 70802 26390 70824 26436
rect 70870 26390 70928 26436
rect 70974 26390 71000 26436
tri 31575 26321 31620 26366 ne
rect 31620 26353 31849 26366
tri 31849 26353 31862 26366 sw
rect 31620 26344 31862 26353
rect 31620 26321 31734 26344
tri 31620 26289 31652 26321 ne
rect 31652 26298 31734 26321
rect 31780 26321 31862 26344
tri 31862 26321 31894 26353 sw
rect 70802 26332 71000 26390
rect 31780 26298 31894 26321
rect 31652 26289 31894 26298
tri 31652 26276 31665 26289 ne
rect 31665 26276 31894 26289
tri 31894 26276 31939 26321 sw
rect 70802 26286 70824 26332
rect 70870 26286 70928 26332
rect 70974 26286 71000 26332
tri 31665 26244 31697 26276 ne
rect 31697 26266 31939 26276
tri 31939 26266 31949 26276 sw
rect 31697 26244 31949 26266
tri 31697 26199 31742 26244 ne
rect 31742 26234 31949 26244
tri 31949 26234 31981 26266 sw
rect 31742 26221 31981 26234
tri 31981 26221 31994 26234 sw
rect 70802 26228 71000 26286
rect 31742 26212 31994 26221
rect 31742 26199 31866 26212
tri 31742 26188 31753 26199 ne
rect 31753 26188 31866 26199
tri 31753 26144 31797 26188 ne
rect 31797 26166 31866 26188
rect 31912 26188 31994 26212
tri 31994 26188 32027 26221 sw
rect 31912 26166 32027 26188
rect 31797 26144 32027 26166
tri 32027 26144 32071 26188 sw
rect 70802 26182 70824 26228
rect 70870 26182 70928 26228
rect 70974 26182 71000 26228
tri 31797 26136 31805 26144 ne
rect 31805 26136 32071 26144
tri 31805 26102 31839 26136 ne
rect 31839 26134 32071 26136
tri 32071 26134 32081 26144 sw
rect 31839 26102 32081 26134
tri 32081 26102 32113 26134 sw
rect 70802 26124 71000 26182
tri 31839 26091 31850 26102 ne
rect 31850 26091 32113 26102
tri 32113 26091 32124 26102 sw
tri 31850 26046 31895 26091 ne
rect 31895 26080 32124 26091
rect 31895 26046 31998 26080
tri 31895 26025 31916 26046 ne
rect 31916 26034 31998 26046
rect 32044 26046 32124 26080
tri 32124 26046 32169 26091 sw
rect 70802 26078 70824 26124
rect 70870 26078 70928 26124
rect 70974 26078 71000 26124
rect 32044 26034 32169 26046
rect 31916 26025 32169 26034
tri 31916 26012 31929 26025 ne
rect 31929 26012 32169 26025
tri 32169 26012 32203 26046 sw
rect 70802 26020 71000 26078
tri 31929 25980 31961 26012 ne
rect 31961 26002 32203 26012
tri 32203 26002 32213 26012 sw
rect 31961 25980 32213 26002
tri 31961 25935 32006 25980 ne
rect 32006 25970 32213 25980
tri 32213 25970 32245 26002 sw
rect 70802 25974 70824 26020
rect 70870 25974 70928 26020
rect 70974 25974 71000 26020
rect 32006 25957 32245 25970
tri 32245 25957 32258 25970 sw
rect 32006 25948 32258 25957
rect 32006 25935 32130 25948
tri 32006 25913 32027 25935 ne
rect 32027 25913 32130 25935
tri 32027 25893 32048 25913 ne
rect 32048 25902 32130 25913
rect 32176 25913 32258 25948
tri 32258 25913 32302 25957 sw
rect 70802 25916 71000 25974
rect 32176 25902 32302 25913
rect 32048 25893 32302 25902
tri 32048 25880 32061 25893 ne
rect 32061 25880 32302 25893
tri 32302 25880 32335 25913 sw
tri 32061 25848 32093 25880 ne
rect 32093 25870 32335 25880
tri 32335 25870 32345 25880 sw
rect 70802 25870 70824 25916
rect 70870 25870 70928 25916
rect 70974 25870 71000 25916
rect 32093 25848 32345 25870
tri 32093 25838 32103 25848 ne
rect 32103 25838 32345 25848
tri 32345 25838 32377 25870 sw
tri 32103 25793 32148 25838 ne
rect 32148 25825 32377 25838
tri 32377 25825 32390 25838 sw
rect 32148 25816 32390 25825
rect 32148 25793 32262 25816
tri 32148 25771 32169 25793 ne
rect 32169 25771 32262 25793
tri 32169 25748 32193 25771 ne
rect 32193 25770 32262 25771
rect 32308 25793 32390 25816
tri 32390 25793 32422 25825 sw
rect 70802 25812 71000 25870
rect 32308 25770 32422 25793
rect 32193 25748 32422 25770
tri 32422 25748 32467 25793 sw
rect 70802 25766 70824 25812
rect 70870 25766 70928 25812
rect 70974 25766 71000 25812
tri 32193 25716 32225 25748 ne
rect 32225 25738 32467 25748
tri 32467 25738 32477 25748 sw
rect 32225 25716 32477 25738
tri 32225 25671 32270 25716 ne
rect 32270 25706 32477 25716
tri 32477 25706 32509 25738 sw
rect 70802 25708 71000 25766
rect 32270 25684 32509 25706
rect 32270 25671 32394 25684
tri 32270 25639 32302 25671 ne
rect 32302 25639 32394 25671
tri 32302 25629 32312 25639 ne
rect 32312 25638 32394 25639
rect 32440 25681 32509 25684
tri 32509 25681 32534 25706 sw
rect 32440 25639 32534 25681
tri 32534 25639 32576 25681 sw
rect 70802 25662 70824 25708
rect 70870 25662 70928 25708
rect 70974 25662 71000 25708
rect 32440 25638 32576 25639
rect 32312 25629 32576 25638
tri 32312 25616 32325 25629 ne
rect 32325 25616 32576 25629
tri 32576 25616 32599 25639 sw
tri 32325 25584 32357 25616 ne
rect 32357 25606 32599 25616
tri 32599 25606 32609 25616 sw
rect 32357 25584 32609 25606
tri 32357 25574 32367 25584 ne
rect 32367 25574 32609 25584
tri 32609 25574 32641 25606 sw
rect 70802 25604 71000 25662
tri 32367 25529 32412 25574 ne
rect 32412 25561 32641 25574
tri 32641 25561 32654 25574 sw
rect 32412 25552 32654 25561
rect 32412 25529 32526 25552
tri 32412 25497 32444 25529 ne
rect 32444 25506 32526 25529
rect 32572 25529 32654 25552
tri 32654 25529 32686 25561 sw
rect 70802 25558 70824 25604
rect 70870 25558 70928 25604
rect 70974 25558 71000 25604
rect 32572 25506 32686 25529
rect 32444 25497 32686 25506
tri 32444 25484 32457 25497 ne
rect 32457 25484 32686 25497
tri 32686 25484 32731 25529 sw
rect 70802 25500 71000 25558
tri 32457 25452 32489 25484 ne
rect 32489 25474 32731 25484
tri 32731 25474 32741 25484 sw
rect 32489 25452 32741 25474
tri 32489 25407 32534 25452 ne
rect 32534 25442 32741 25452
tri 32741 25442 32773 25474 sw
rect 70802 25454 70824 25500
rect 70870 25454 70928 25500
rect 70974 25454 71000 25500
rect 32534 25429 32773 25442
tri 32773 25429 32786 25442 sw
rect 32534 25420 32786 25429
rect 32534 25407 32658 25420
tri 32534 25365 32576 25407 ne
rect 32576 25374 32658 25407
rect 32704 25410 32786 25420
tri 32786 25410 32805 25429 sw
rect 32704 25374 32805 25410
rect 32576 25365 32805 25374
tri 32805 25365 32851 25410 sw
rect 70802 25396 71000 25454
tri 32576 25352 32589 25365 ne
rect 32589 25361 32851 25365
tri 32851 25361 32854 25365 sw
rect 32589 25352 32854 25361
tri 32854 25352 32863 25361 sw
tri 32589 25320 32621 25352 ne
rect 32621 25342 32863 25352
tri 32863 25342 32873 25352 sw
rect 70802 25350 70824 25396
rect 70870 25350 70928 25396
rect 70974 25350 71000 25396
rect 32621 25320 32873 25342
tri 32621 25310 32631 25320 ne
rect 32631 25310 32873 25320
tri 32873 25310 32905 25342 sw
tri 32631 25265 32676 25310 ne
rect 32676 25297 32905 25310
tri 32905 25297 32918 25310 sw
rect 32676 25288 32918 25297
rect 32676 25265 32790 25288
tri 32676 25233 32708 25265 ne
rect 32708 25242 32790 25265
rect 32836 25265 32918 25288
tri 32918 25265 32950 25297 sw
rect 70802 25292 71000 25350
rect 32836 25242 32950 25265
rect 32708 25233 32950 25242
tri 32708 25220 32721 25233 ne
rect 32721 25220 32950 25233
tri 32950 25220 32995 25265 sw
rect 70802 25246 70824 25292
rect 70870 25246 70928 25292
rect 70974 25246 71000 25292
tri 32721 25188 32753 25220 ne
rect 32753 25210 32995 25220
tri 32995 25210 33005 25220 sw
rect 32753 25188 33005 25210
tri 32753 25143 32798 25188 ne
rect 32798 25178 33005 25188
tri 33005 25178 33037 25210 sw
rect 70802 25188 71000 25246
rect 32798 25165 33037 25178
tri 33037 25165 33050 25178 sw
rect 32798 25156 33050 25165
rect 32798 25143 32922 25156
tri 32798 25101 32840 25143 ne
rect 32840 25110 32922 25143
rect 32968 25135 33050 25156
tri 33050 25135 33080 25165 sw
rect 70802 25142 70824 25188
rect 70870 25142 70928 25188
rect 70974 25142 71000 25188
rect 32968 25110 33080 25135
rect 32840 25101 33080 25110
tri 32840 25090 32851 25101 ne
rect 32851 25090 33080 25101
tri 33080 25090 33125 25135 sw
tri 32851 25088 32853 25090 ne
rect 32853 25088 33125 25090
tri 33125 25088 33127 25090 sw
tri 32853 25056 32885 25088 ne
rect 32885 25078 33127 25088
tri 33127 25078 33137 25088 sw
rect 70802 25084 71000 25142
rect 32885 25056 33137 25078
tri 32885 25046 32895 25056 ne
rect 32895 25046 33137 25056
tri 33137 25046 33169 25078 sw
tri 32895 25042 32899 25046 ne
rect 32899 25042 33169 25046
tri 32899 24997 32944 25042 ne
rect 32944 25033 33169 25042
tri 33169 25033 33182 25046 sw
rect 70802 25038 70824 25084
rect 70870 25038 70928 25084
rect 70974 25038 71000 25084
rect 32944 25024 33182 25033
rect 32944 24997 33054 25024
tri 32944 24969 32972 24997 ne
rect 32972 24978 33054 24997
rect 33100 24997 33182 25024
tri 33182 24997 33219 25033 sw
rect 33100 24978 33219 24997
rect 32972 24969 33219 24978
tri 32972 24956 32985 24969 ne
rect 32985 24956 33219 24969
tri 33219 24956 33259 24997 sw
rect 70802 24980 71000 25038
tri 32985 24924 33017 24956 ne
rect 33017 24951 33259 24956
tri 33259 24951 33264 24956 sw
rect 33017 24946 33264 24951
tri 33264 24946 33269 24951 sw
rect 33017 24924 33269 24946
tri 33017 24879 33062 24924 ne
rect 33062 24914 33269 24924
tri 33269 24914 33301 24946 sw
rect 70802 24934 70824 24980
rect 70870 24934 70928 24980
rect 70974 24934 71000 24980
rect 33062 24901 33301 24914
tri 33301 24901 33314 24914 sw
rect 33062 24892 33314 24901
rect 33062 24879 33186 24892
tri 33062 24837 33104 24879 ne
rect 33104 24846 33186 24879
rect 33232 24869 33314 24892
tri 33314 24869 33346 24901 sw
rect 70802 24876 71000 24934
rect 33232 24846 33346 24869
rect 33104 24837 33346 24846
tri 33104 24816 33125 24837 ne
rect 33125 24824 33346 24837
tri 33346 24824 33391 24869 sw
rect 70802 24830 70824 24876
rect 70870 24830 70928 24876
rect 70974 24830 71000 24876
rect 33125 24816 33391 24824
tri 33391 24816 33399 24824 sw
tri 33125 24792 33149 24816 ne
rect 33149 24814 33399 24816
tri 33399 24814 33401 24816 sw
rect 33149 24792 33401 24814
tri 33149 24782 33159 24792 ne
rect 33159 24782 33401 24792
tri 33401 24782 33433 24814 sw
tri 33159 24737 33204 24782 ne
rect 33204 24769 33433 24782
tri 33433 24769 33446 24782 sw
rect 70802 24772 71000 24830
rect 33204 24760 33446 24769
rect 33204 24737 33318 24760
tri 33204 24692 33249 24737 ne
rect 33249 24714 33318 24737
rect 33364 24737 33446 24760
tri 33446 24737 33478 24769 sw
rect 33364 24714 33478 24737
rect 33249 24692 33478 24714
tri 33478 24692 33523 24737 sw
rect 70802 24726 70824 24772
rect 70870 24726 70928 24772
rect 70974 24726 71000 24772
tri 33249 24677 33264 24692 ne
rect 33264 24682 33523 24692
tri 33523 24682 33533 24692 sw
rect 33264 24677 33533 24682
tri 33264 24632 33309 24677 ne
rect 33309 24650 33533 24677
tri 33533 24650 33565 24682 sw
rect 70802 24668 71000 24726
rect 33309 24637 33565 24650
tri 33565 24637 33578 24650 sw
rect 33309 24632 33578 24637
tri 33578 24632 33583 24637 sw
tri 33309 24587 33354 24632 ne
rect 33354 24628 33583 24632
rect 33354 24587 33450 24628
tri 33354 24573 33368 24587 ne
rect 33368 24582 33450 24587
rect 33496 24587 33583 24628
tri 33583 24587 33629 24632 sw
rect 70802 24622 70824 24668
rect 70870 24622 70928 24668
rect 70974 24622 71000 24668
rect 33496 24582 33629 24587
rect 33368 24573 33629 24582
tri 33368 24541 33399 24573 ne
rect 33399 24560 33629 24573
tri 33629 24560 33655 24587 sw
rect 70802 24564 71000 24622
rect 33399 24550 33655 24560
tri 33655 24550 33665 24560 sw
rect 33399 24541 33665 24550
tri 33665 24541 33674 24550 sw
tri 33399 24528 33413 24541 ne
rect 33413 24528 33674 24541
tri 33413 24518 33423 24528 ne
rect 33423 24518 33674 24528
tri 33674 24518 33697 24541 sw
rect 70802 24518 70824 24564
rect 70870 24518 70928 24564
rect 70974 24518 71000 24564
tri 33423 24473 33468 24518 ne
rect 33468 24505 33697 24518
tri 33697 24505 33710 24518 sw
rect 33468 24496 33710 24505
rect 33468 24473 33582 24496
tri 33468 24441 33500 24473 ne
rect 33500 24450 33582 24473
rect 33628 24473 33710 24496
tri 33710 24473 33742 24505 sw
rect 33628 24450 33742 24473
rect 33500 24441 33742 24450
tri 33500 24428 33513 24441 ne
rect 33513 24428 33742 24441
tri 33742 24428 33787 24473 sw
rect 70802 24460 71000 24518
tri 33513 24396 33545 24428 ne
rect 33545 24418 33787 24428
tri 33787 24418 33797 24428 sw
rect 33545 24396 33797 24418
tri 33545 24351 33590 24396 ne
rect 33590 24386 33797 24396
tri 33797 24386 33829 24418 sw
rect 70802 24414 70824 24460
rect 70870 24414 70928 24460
rect 70974 24414 71000 24460
rect 33590 24373 33829 24386
tri 33829 24373 33842 24386 sw
rect 33590 24364 33842 24373
rect 33590 24351 33714 24364
tri 33590 24312 33629 24351 ne
rect 33629 24318 33714 24351
rect 33760 24341 33842 24364
tri 33842 24341 33874 24373 sw
rect 70802 24356 71000 24414
rect 33760 24318 33874 24341
rect 33629 24312 33874 24318
tri 33629 24267 33674 24312 ne
rect 33674 24296 33874 24312
tri 33874 24296 33919 24341 sw
rect 70802 24310 70824 24356
rect 70870 24310 70928 24356
rect 70974 24310 71000 24356
rect 33674 24286 33919 24296
tri 33919 24286 33929 24296 sw
rect 33674 24267 33929 24286
tri 33929 24267 33948 24286 sw
tri 33674 24264 33677 24267 ne
rect 33677 24264 33948 24267
tri 33677 24254 33687 24264 ne
rect 33687 24254 33948 24264
tri 33948 24254 33961 24267 sw
tri 33687 24209 33732 24254 ne
rect 33732 24232 33961 24254
rect 33732 24209 33846 24232
tri 33732 24177 33764 24209 ne
rect 33764 24186 33846 24209
rect 33892 24222 33961 24232
tri 33961 24222 33993 24254 sw
rect 70802 24252 71000 24310
rect 33892 24209 33993 24222
tri 33993 24209 34006 24222 sw
rect 33892 24186 34006 24209
rect 33764 24177 34006 24186
tri 33764 24164 33777 24177 ne
rect 33777 24164 34006 24177
tri 34006 24164 34051 24209 sw
rect 70802 24206 70824 24252
rect 70870 24206 70928 24252
rect 70974 24206 71000 24252
tri 33777 24132 33809 24164 ne
rect 33809 24154 34051 24164
tri 34051 24154 34061 24164 sw
rect 33809 24132 34061 24154
tri 33809 24087 33854 24132 ne
rect 33854 24122 34061 24132
tri 34061 24122 34093 24154 sw
rect 70802 24148 71000 24206
rect 33854 24109 34093 24122
tri 34093 24109 34106 24122 sw
rect 33854 24100 34106 24109
rect 33854 24087 33978 24100
tri 33854 24045 33896 24087 ne
rect 33896 24054 33978 24087
rect 34024 24077 34106 24100
tri 34106 24077 34138 24109 sw
rect 70802 24102 70824 24148
rect 70870 24102 70928 24148
rect 70974 24102 71000 24148
rect 34024 24054 34138 24077
rect 33896 24045 34138 24054
tri 33896 24000 33941 24045 ne
rect 33941 24032 34138 24045
tri 34138 24032 34183 24077 sw
rect 70802 24044 71000 24102
rect 33941 24022 34183 24032
tri 34183 24022 34193 24032 sw
rect 33941 24000 34193 24022
tri 33941 23993 33948 24000 ne
rect 33948 23993 34193 24000
tri 34193 23993 34223 24022 sw
rect 70802 23998 70824 24044
rect 70870 23998 70928 24044
rect 70974 23998 71000 24044
tri 33948 23990 33951 23993 ne
rect 33951 23990 34223 23993
tri 34223 23990 34225 23993 sw
tri 33951 23947 33993 23990 ne
rect 33993 23977 34225 23990
tri 34225 23977 34238 23990 sw
rect 33993 23968 34238 23977
rect 33993 23947 34110 23968
tri 33993 23902 34039 23947 ne
rect 34039 23922 34110 23947
rect 34156 23947 34238 23968
tri 34238 23947 34268 23977 sw
rect 34156 23922 34268 23947
rect 34039 23902 34268 23922
tri 34268 23902 34313 23947 sw
rect 70802 23940 71000 23998
tri 34039 23900 34041 23902 ne
rect 34041 23900 34313 23902
tri 34313 23900 34315 23902 sw
tri 34041 23868 34073 23900 ne
rect 34073 23868 34315 23900
tri 34073 23858 34083 23868 ne
rect 34083 23858 34315 23868
tri 34315 23858 34357 23900 sw
rect 70802 23894 70824 23940
rect 70870 23894 70928 23940
rect 70974 23894 71000 23940
tri 34083 23813 34128 23858 ne
rect 34128 23845 34357 23858
tri 34357 23845 34370 23858 sw
rect 34128 23836 34370 23845
rect 34128 23813 34242 23836
tri 34128 23781 34160 23813 ne
rect 34160 23790 34242 23813
rect 34288 23813 34370 23836
tri 34370 23813 34402 23845 sw
rect 70802 23836 71000 23894
rect 34288 23790 34402 23813
rect 34160 23781 34402 23790
tri 34160 23768 34173 23781 ne
rect 34173 23768 34402 23781
tri 34402 23768 34447 23813 sw
rect 70802 23790 70824 23836
rect 70870 23790 70928 23836
rect 70974 23790 71000 23836
tri 34173 23736 34205 23768 ne
rect 34205 23758 34447 23768
tri 34447 23758 34457 23768 sw
rect 34205 23736 34457 23758
tri 34205 23718 34223 23736 ne
rect 34223 23726 34457 23736
tri 34457 23726 34489 23758 sw
rect 70802 23732 71000 23790
rect 34223 23718 34489 23726
tri 34489 23718 34497 23726 sw
tri 34223 23673 34268 23718 ne
rect 34268 23713 34497 23718
tri 34497 23713 34502 23718 sw
rect 34268 23704 34502 23713
rect 34268 23673 34374 23704
tri 34268 23649 34292 23673 ne
rect 34292 23658 34374 23673
rect 34420 23681 34502 23704
tri 34502 23681 34534 23713 sw
rect 70802 23686 70824 23732
rect 70870 23686 70928 23732
rect 70974 23686 71000 23732
rect 34420 23658 34534 23681
rect 34292 23649 34534 23658
tri 34292 23636 34305 23649 ne
rect 34305 23636 34534 23649
tri 34534 23636 34579 23681 sw
tri 34305 23604 34337 23636 ne
rect 34337 23626 34579 23636
tri 34579 23626 34589 23636 sw
rect 70802 23628 71000 23686
rect 34337 23604 34589 23626
tri 34337 23594 34347 23604 ne
rect 34347 23594 34589 23604
tri 34589 23594 34621 23626 sw
tri 34347 23583 34358 23594 ne
rect 34358 23583 34621 23594
tri 34358 23537 34403 23583 ne
rect 34403 23581 34621 23583
tri 34621 23581 34634 23594 sw
rect 70802 23582 70824 23628
rect 70870 23582 70928 23628
rect 70974 23582 71000 23628
rect 34403 23572 34634 23581
rect 34403 23537 34506 23572
tri 34403 23517 34424 23537 ne
rect 34424 23526 34506 23537
rect 34552 23537 34634 23572
tri 34634 23537 34678 23581 sw
rect 34552 23526 34678 23537
rect 34424 23517 34678 23526
tri 34424 23504 34437 23517 ne
rect 34437 23504 34678 23517
tri 34678 23504 34711 23537 sw
rect 70802 23524 71000 23582
tri 34437 23472 34469 23504 ne
rect 34469 23494 34711 23504
tri 34711 23494 34721 23504 sw
rect 34469 23472 34721 23494
tri 34469 23444 34497 23472 ne
rect 34497 23462 34721 23472
tri 34721 23462 34753 23494 sw
rect 70802 23478 70824 23524
rect 70870 23478 70928 23524
rect 70974 23478 71000 23524
rect 34497 23449 34753 23462
tri 34753 23449 34766 23462 sw
rect 34497 23444 34766 23449
tri 34766 23444 34771 23449 sw
tri 34497 23399 34542 23444 ne
rect 34542 23440 34771 23444
rect 34542 23399 34638 23440
tri 34542 23385 34556 23399 ne
rect 34556 23394 34638 23399
rect 34684 23417 34771 23440
tri 34771 23417 34798 23444 sw
rect 70802 23420 71000 23478
rect 34684 23394 34798 23417
rect 34556 23385 34798 23394
tri 34556 23372 34569 23385 ne
rect 34569 23372 34798 23385
tri 34798 23372 34843 23417 sw
rect 70802 23374 70824 23420
rect 70870 23374 70928 23420
rect 70974 23374 71000 23420
tri 34569 23340 34601 23372 ne
rect 34601 23362 34843 23372
tri 34843 23362 34853 23372 sw
rect 34601 23340 34853 23362
tri 34601 23330 34611 23340 ne
rect 34611 23330 34853 23340
tri 34853 23330 34885 23362 sw
tri 34611 23285 34656 23330 ne
rect 34656 23317 34885 23330
tri 34885 23317 34898 23330 sw
rect 34656 23308 34898 23317
rect 34656 23285 34770 23308
tri 34656 23253 34688 23285 ne
rect 34688 23262 34770 23285
rect 34816 23285 34898 23308
tri 34898 23285 34930 23317 sw
rect 70802 23316 71000 23374
rect 34816 23262 34930 23285
rect 34688 23253 34930 23262
tri 34688 23240 34701 23253 ne
rect 34701 23240 34930 23253
tri 34930 23240 34975 23285 sw
rect 70802 23270 70824 23316
rect 70870 23270 70928 23316
rect 70974 23270 71000 23316
tri 34701 23208 34733 23240 ne
rect 34733 23230 34975 23240
tri 34975 23230 34985 23240 sw
rect 34733 23208 34985 23230
tri 34733 23173 34768 23208 ne
rect 34768 23198 34985 23208
tri 34985 23198 35017 23230 sw
rect 70802 23212 71000 23270
rect 34768 23185 35017 23198
tri 35017 23185 35030 23198 sw
rect 34768 23176 35030 23185
rect 34768 23173 34902 23176
tri 34768 23169 34771 23173 ne
rect 34771 23169 34902 23173
tri 34771 23124 34817 23169 ne
rect 34817 23130 34902 23169
rect 34948 23173 35030 23176
tri 35030 23173 35043 23185 sw
rect 34948 23169 35043 23173
tri 35043 23169 35046 23173 sw
rect 34948 23130 35046 23169
rect 34817 23127 35046 23130
tri 35046 23127 35088 23169 sw
rect 70802 23166 70824 23212
rect 70870 23166 70928 23212
rect 70974 23166 71000 23212
rect 34817 23124 35088 23127
tri 34817 23121 34820 23124 ne
rect 34820 23121 35088 23124
tri 34820 23108 34833 23121 ne
rect 34833 23108 35088 23121
tri 35088 23108 35107 23127 sw
rect 70802 23108 71000 23166
tri 34833 23076 34865 23108 ne
rect 34865 23098 35107 23108
tri 35107 23098 35117 23108 sw
rect 34865 23076 35117 23098
tri 34865 23066 34875 23076 ne
rect 34875 23066 35117 23076
tri 35117 23066 35149 23098 sw
tri 34875 23021 34920 23066 ne
rect 34920 23053 35149 23066
tri 35149 23053 35162 23066 sw
rect 70802 23062 70824 23108
rect 70870 23062 70928 23108
rect 70974 23062 71000 23108
rect 34920 23044 35162 23053
rect 34920 23021 35034 23044
tri 34920 22989 34952 23021 ne
rect 34952 22998 35034 23021
rect 35080 23021 35162 23044
tri 35162 23021 35194 23053 sw
rect 35080 22998 35194 23021
rect 34952 22989 35194 22998
tri 34952 22976 34965 22989 ne
rect 34965 22976 35194 22989
tri 35194 22976 35239 23021 sw
rect 70802 23004 71000 23062
tri 34965 22944 34997 22976 ne
rect 34997 22966 35239 22976
tri 35239 22966 35249 22976 sw
rect 34997 22944 35249 22966
tri 34997 22899 35042 22944 ne
rect 35042 22934 35249 22944
tri 35249 22934 35281 22966 sw
rect 70802 22958 70824 23004
rect 70870 22958 70928 23004
rect 70974 22958 71000 23004
rect 35042 22921 35281 22934
tri 35281 22921 35294 22934 sw
rect 35042 22912 35294 22921
rect 35042 22899 35166 22912
tri 35042 22895 35046 22899 ne
rect 35046 22895 35166 22899
tri 35046 22853 35088 22895 ne
rect 35088 22866 35166 22895
rect 35212 22895 35294 22912
tri 35294 22895 35320 22921 sw
rect 70802 22900 71000 22958
rect 35212 22889 35320 22895
tri 35320 22889 35326 22895 sw
rect 35212 22866 35326 22889
rect 35088 22853 35326 22866
tri 35088 22844 35097 22853 ne
rect 35097 22844 35326 22853
tri 35326 22844 35371 22889 sw
rect 70802 22854 70824 22900
rect 70870 22854 70928 22900
rect 70974 22854 71000 22900
tri 35097 22808 35133 22844 ne
rect 35133 22834 35371 22844
tri 35371 22834 35381 22844 sw
rect 35133 22808 35381 22834
tri 35133 22802 35139 22808 ne
rect 35139 22802 35381 22808
tri 35381 22802 35413 22834 sw
tri 35139 22757 35184 22802 ne
rect 35184 22780 35413 22802
rect 35184 22757 35298 22780
tri 35184 22725 35216 22757 ne
rect 35216 22734 35298 22757
rect 35344 22763 35413 22780
tri 35413 22763 35453 22802 sw
rect 70802 22796 71000 22854
rect 35344 22757 35453 22763
tri 35453 22757 35458 22763 sw
rect 35344 22734 35458 22757
rect 35216 22725 35458 22734
tri 35216 22712 35229 22725 ne
rect 35229 22712 35458 22725
tri 35458 22712 35503 22757 sw
rect 70802 22750 70824 22796
rect 70870 22750 70928 22796
rect 70974 22750 71000 22796
tri 35229 22680 35261 22712 ne
rect 35261 22702 35503 22712
tri 35503 22702 35513 22712 sw
rect 35261 22680 35513 22702
tri 35261 22635 35306 22680 ne
rect 35306 22670 35513 22680
tri 35513 22670 35545 22702 sw
rect 70802 22692 71000 22750
rect 35306 22657 35545 22670
tri 35545 22657 35558 22670 sw
rect 35306 22648 35558 22657
rect 35306 22635 35430 22648
tri 35306 22621 35320 22635 ne
rect 35320 22621 35430 22635
tri 35320 22593 35348 22621 ne
rect 35348 22602 35430 22621
rect 35476 22621 35558 22648
tri 35558 22621 35595 22657 sw
rect 70802 22646 70824 22692
rect 70870 22646 70928 22692
rect 70974 22646 71000 22692
rect 35476 22602 35595 22621
rect 35348 22593 35595 22602
tri 35348 22580 35361 22593 ne
rect 35361 22580 35595 22593
tri 35595 22580 35635 22621 sw
rect 70802 22588 71000 22646
tri 35361 22548 35393 22580 ne
rect 35393 22570 35635 22580
tri 35635 22570 35645 22580 sw
rect 35393 22548 35645 22570
tri 35393 22538 35403 22548 ne
rect 35403 22538 35645 22548
tri 35645 22538 35677 22570 sw
rect 70802 22542 70824 22588
rect 70870 22542 70928 22588
rect 70974 22542 71000 22588
tri 35403 22493 35448 22538 ne
rect 35448 22525 35677 22538
tri 35677 22525 35690 22538 sw
rect 35448 22516 35690 22525
rect 35448 22493 35562 22516
tri 35448 22488 35453 22493 ne
rect 35453 22488 35562 22493
tri 35453 22448 35493 22488 ne
rect 35493 22470 35562 22488
rect 35608 22493 35690 22516
tri 35690 22493 35722 22525 sw
rect 35608 22470 35722 22493
rect 35493 22448 35722 22470
tri 35722 22448 35767 22493 sw
rect 70802 22484 71000 22542
tri 35493 22416 35525 22448 ne
rect 35525 22443 35767 22448
tri 35767 22443 35772 22448 sw
rect 35525 22416 35772 22443
tri 35525 22371 35570 22416 ne
rect 35570 22406 35772 22416
tri 35772 22406 35809 22443 sw
rect 70802 22438 70824 22484
rect 70870 22438 70928 22484
rect 70974 22438 71000 22484
rect 35570 22393 35809 22406
tri 35809 22393 35822 22406 sw
rect 35570 22391 35822 22393
tri 35822 22391 35824 22393 sw
rect 35570 22384 35824 22391
rect 35570 22371 35694 22384
tri 35570 22346 35595 22371 ne
rect 35595 22346 35694 22371
tri 35595 22329 35612 22346 ne
rect 35612 22338 35694 22346
rect 35740 22346 35824 22384
tri 35824 22346 35869 22391 sw
rect 70802 22380 71000 22438
rect 35740 22338 35869 22346
rect 35612 22329 35869 22338
tri 35612 22316 35625 22329 ne
rect 35625 22316 35869 22329
tri 35869 22316 35899 22346 sw
rect 70802 22334 70824 22380
rect 70870 22334 70928 22380
rect 70974 22334 71000 22380
tri 35625 22284 35657 22316 ne
rect 35657 22306 35899 22316
tri 35899 22306 35909 22316 sw
rect 35657 22284 35909 22306
tri 35657 22274 35667 22284 ne
rect 35667 22274 35909 22284
tri 35909 22274 35941 22306 sw
rect 70802 22276 71000 22334
tri 35667 22229 35712 22274 ne
rect 35712 22261 35941 22274
tri 35941 22261 35954 22274 sw
rect 35712 22252 35954 22261
rect 35712 22229 35826 22252
tri 35712 22197 35744 22229 ne
rect 35744 22206 35826 22229
rect 35872 22229 35954 22252
tri 35954 22229 35986 22261 sw
rect 70802 22230 70824 22276
rect 70870 22230 70928 22276
rect 70974 22230 71000 22276
rect 35872 22206 35986 22229
rect 35744 22197 35986 22206
tri 35744 22184 35757 22197 ne
rect 35757 22184 35986 22197
tri 35986 22184 36031 22229 sw
tri 35757 22152 35789 22184 ne
rect 35789 22174 36031 22184
tri 36031 22174 36041 22184 sw
rect 35789 22152 36041 22174
tri 35789 22123 35817 22152 ne
rect 35817 22142 36041 22152
tri 36041 22142 36073 22174 sw
rect 70802 22172 71000 22230
rect 35817 22129 36073 22142
tri 36073 22129 36086 22142 sw
rect 35817 22123 36086 22129
tri 36086 22123 36092 22129 sw
rect 70802 22126 70824 22172
rect 70870 22126 70928 22172
rect 70974 22126 71000 22172
tri 35817 22078 35863 22123 ne
rect 35863 22120 36092 22123
rect 35863 22078 35958 22120
tri 35863 22072 35869 22078 ne
rect 35869 22074 35958 22078
rect 36004 22078 36092 22120
tri 36092 22078 36137 22123 sw
rect 36004 22074 36137 22078
rect 35869 22072 36137 22074
tri 36137 22072 36143 22078 sw
tri 35869 22065 35876 22072 ne
rect 35876 22065 36143 22072
tri 35876 22052 35889 22065 ne
rect 35889 22052 36143 22065
tri 36143 22052 36163 22072 sw
rect 70802 22068 71000 22126
tri 35889 22020 35921 22052 ne
rect 35921 22042 36163 22052
tri 36163 22042 36173 22052 sw
rect 35921 22020 36173 22042
tri 35921 22010 35931 22020 ne
rect 35931 22010 36173 22020
tri 36173 22010 36205 22042 sw
rect 70802 22022 70824 22068
rect 70870 22022 70928 22068
rect 70974 22022 71000 22068
tri 35931 21965 35976 22010 ne
rect 35976 21997 36205 22010
tri 36205 21997 36218 22010 sw
rect 35976 21988 36218 21997
rect 35976 21965 36090 21988
tri 35976 21933 36008 21965 ne
rect 36008 21942 36090 21965
rect 36136 21965 36218 21988
tri 36218 21965 36250 21997 sw
rect 36136 21942 36250 21965
rect 36008 21933 36250 21942
tri 36008 21920 36021 21933 ne
rect 36021 21920 36250 21933
tri 36250 21920 36295 21965 sw
rect 70802 21964 71000 22022
tri 36021 21888 36053 21920 ne
rect 36053 21910 36295 21920
tri 36295 21910 36305 21920 sw
rect 70802 21918 70824 21964
rect 70870 21918 70928 21964
rect 70974 21918 71000 21964
rect 36053 21888 36305 21910
tri 36053 21843 36098 21888 ne
rect 36098 21878 36305 21888
tri 36305 21878 36337 21910 sw
rect 36098 21865 36337 21878
tri 36337 21865 36350 21878 sw
rect 36098 21856 36350 21865
rect 36098 21843 36222 21856
tri 36098 21801 36140 21843 ne
rect 36140 21810 36222 21843
rect 36268 21843 36350 21856
tri 36350 21843 36373 21865 sw
rect 70802 21860 71000 21918
rect 36268 21810 36373 21843
rect 36140 21801 36373 21810
tri 36140 21797 36143 21801 ne
rect 36143 21797 36373 21801
tri 36373 21797 36418 21843 sw
rect 70802 21814 70824 21860
rect 70870 21814 70928 21860
rect 70974 21814 71000 21860
tri 36143 21788 36153 21797 ne
rect 36153 21788 36418 21797
tri 36418 21788 36427 21797 sw
tri 36153 21756 36185 21788 ne
rect 36185 21778 36427 21788
tri 36427 21778 36437 21788 sw
rect 36185 21756 36437 21778
tri 36185 21746 36195 21756 ne
rect 36195 21746 36437 21756
tri 36437 21746 36469 21778 sw
rect 70802 21756 71000 21814
tri 36195 21713 36227 21746 ne
rect 36227 21733 36469 21746
tri 36469 21733 36482 21746 sw
rect 36227 21724 36482 21733
rect 36227 21713 36354 21724
tri 36227 21669 36272 21713 ne
rect 36272 21678 36354 21713
rect 36400 21713 36482 21724
tri 36482 21713 36502 21733 sw
rect 36400 21678 36502 21713
rect 36272 21669 36502 21678
tri 36272 21656 36285 21669 ne
rect 36285 21668 36502 21669
tri 36502 21668 36547 21713 sw
rect 70802 21710 70824 21756
rect 70870 21710 70928 21756
rect 70974 21710 71000 21756
rect 36285 21656 36547 21668
tri 36547 21656 36559 21668 sw
tri 36285 21624 36317 21656 ne
rect 36317 21646 36559 21656
tri 36559 21646 36569 21656 sw
rect 70802 21652 71000 21710
rect 36317 21624 36569 21646
tri 36317 21579 36362 21624 ne
rect 36362 21614 36569 21624
tri 36569 21614 36601 21646 sw
rect 36362 21601 36601 21614
tri 36601 21601 36614 21614 sw
rect 70802 21606 70824 21652
rect 70870 21606 70928 21652
rect 70974 21606 71000 21652
rect 36362 21592 36614 21601
rect 36362 21579 36486 21592
tri 36362 21537 36404 21579 ne
rect 36404 21546 36486 21579
rect 36532 21569 36614 21592
tri 36614 21569 36646 21601 sw
rect 36532 21546 36646 21569
rect 36404 21537 36646 21546
tri 36404 21523 36418 21537 ne
rect 36418 21524 36646 21537
tri 36646 21524 36691 21569 sw
rect 70802 21548 71000 21606
rect 36418 21523 36691 21524
tri 36691 21523 36692 21524 sw
tri 36418 21492 36449 21523 ne
rect 36449 21514 36692 21523
tri 36692 21514 36701 21523 sw
rect 36449 21492 36701 21514
tri 36449 21482 36459 21492 ne
rect 36459 21482 36701 21492
tri 36701 21482 36733 21514 sw
rect 70802 21502 70824 21548
rect 70870 21502 70928 21548
rect 70974 21502 71000 21548
tri 36459 21437 36504 21482 ne
rect 36504 21469 36733 21482
tri 36733 21469 36746 21482 sw
rect 36504 21460 36746 21469
rect 36504 21437 36618 21460
tri 36504 21394 36547 21437 ne
rect 36547 21414 36618 21437
rect 36664 21437 36746 21460
tri 36746 21437 36778 21469 sw
rect 70802 21444 71000 21502
rect 36664 21414 36778 21437
rect 36547 21394 36778 21414
tri 36547 21392 36549 21394 ne
rect 36549 21392 36778 21394
tri 36778 21392 36823 21437 sw
rect 70802 21398 70824 21444
rect 70870 21398 70928 21444
rect 70974 21398 71000 21444
tri 36549 21349 36592 21392 ne
rect 36592 21382 36823 21392
tri 36823 21382 36833 21392 sw
rect 36592 21350 36833 21382
tri 36833 21350 36865 21382 sw
rect 36592 21349 36865 21350
tri 36865 21349 36867 21350 sw
tri 36592 21303 36637 21349 ne
rect 36637 21328 36867 21349
rect 36637 21303 36750 21328
tri 36637 21273 36668 21303 ne
rect 36668 21282 36750 21303
rect 36796 21303 36867 21328
tri 36867 21303 36912 21349 sw
rect 70802 21340 71000 21398
rect 36796 21282 36912 21303
rect 36668 21273 36912 21282
tri 36668 21249 36692 21273 ne
rect 36692 21260 36912 21273
tri 36912 21260 36955 21303 sw
rect 70802 21294 70824 21340
rect 70870 21294 70928 21340
rect 70974 21294 71000 21340
rect 36692 21250 36955 21260
tri 36955 21250 36965 21260 sw
rect 36692 21249 36965 21250
tri 36965 21249 36967 21250 sw
tri 36692 21228 36713 21249 ne
rect 36713 21228 36967 21249
tri 36713 21218 36723 21228 ne
rect 36723 21218 36967 21228
tri 36967 21218 36997 21249 sw
rect 70802 21236 71000 21294
tri 36723 21173 36768 21218 ne
rect 36768 21205 36997 21218
tri 36997 21205 37010 21218 sw
rect 36768 21196 37010 21205
rect 36768 21173 36882 21196
tri 36768 21141 36800 21173 ne
rect 36800 21150 36882 21173
rect 36928 21173 37010 21196
tri 37010 21173 37042 21205 sw
rect 70802 21190 70824 21236
rect 70870 21190 70928 21236
rect 70974 21190 71000 21236
rect 36928 21150 37042 21173
rect 36800 21141 37042 21150
tri 36800 21128 36813 21141 ne
rect 36813 21128 37042 21141
tri 37042 21128 37087 21173 sw
rect 70802 21132 71000 21190
tri 36813 21096 36845 21128 ne
rect 36845 21118 37087 21128
tri 37087 21118 37097 21128 sw
rect 36845 21096 37097 21118
tri 36845 21051 36890 21096 ne
rect 36890 21086 37097 21096
tri 37097 21086 37129 21118 sw
rect 70802 21086 70824 21132
rect 70870 21086 70928 21132
rect 70974 21086 71000 21132
rect 36890 21073 37129 21086
tri 37129 21073 37142 21086 sw
rect 36890 21064 37142 21073
rect 36890 21051 37014 21064
tri 36890 21029 36912 21051 ne
rect 36912 21029 37014 21051
tri 36912 20984 36957 21029 ne
rect 36957 21018 37014 21029
rect 37060 21041 37142 21064
tri 37142 21041 37174 21073 sw
rect 37060 21018 37174 21041
rect 36957 20996 37174 21018
tri 37174 20996 37219 21041 sw
rect 70802 21028 71000 21086
rect 36957 20986 37219 20996
tri 37219 20986 37229 20996 sw
rect 36957 20984 37229 20986
tri 36957 20974 36967 20984 ne
rect 36967 20974 37229 20984
tri 37229 20974 37241 20986 sw
rect 70802 20982 70824 21028
rect 70870 20982 70928 21028
rect 70974 20982 71000 21028
tri 36967 20964 36977 20974 ne
rect 36977 20964 37241 20974
tri 36977 20954 36987 20964 ne
rect 36987 20954 37241 20964
tri 37241 20954 37261 20974 sw
tri 36987 20909 37032 20954 ne
rect 37032 20939 37261 20954
tri 37261 20939 37277 20954 sw
rect 37032 20932 37277 20939
rect 37032 20909 37146 20932
tri 37032 20877 37064 20909 ne
rect 37064 20886 37146 20909
rect 37192 20909 37277 20932
tri 37277 20909 37306 20939 sw
rect 70802 20924 71000 20982
rect 37192 20886 37306 20909
rect 37064 20877 37306 20886
tri 37064 20864 37077 20877 ne
rect 37077 20864 37306 20877
tri 37306 20864 37351 20909 sw
rect 70802 20878 70824 20924
rect 70870 20878 70928 20924
rect 70974 20878 71000 20924
tri 37077 20832 37109 20864 ne
rect 37109 20854 37351 20864
tri 37351 20854 37361 20864 sw
rect 37109 20832 37361 20854
tri 37109 20787 37154 20832 ne
rect 37154 20822 37361 20832
tri 37361 20822 37393 20854 sw
rect 37154 20809 37393 20822
tri 37393 20809 37406 20822 sw
rect 70802 20820 71000 20878
rect 37154 20800 37406 20809
rect 37154 20787 37278 20800
tri 37154 20745 37196 20787 ne
rect 37196 20754 37278 20787
rect 37324 20777 37406 20800
tri 37406 20777 37438 20809 sw
rect 37324 20754 37438 20777
rect 37196 20745 37438 20754
tri 37196 20700 37241 20745 ne
rect 37241 20732 37438 20745
tri 37438 20732 37483 20777 sw
rect 70802 20774 70824 20820
rect 70870 20774 70928 20820
rect 70974 20774 71000 20820
rect 37241 20722 37483 20732
tri 37483 20722 37493 20732 sw
rect 37241 20700 37493 20722
tri 37493 20700 37515 20722 sw
rect 70802 20716 71000 20774
tri 37241 20690 37251 20700 ne
rect 37251 20690 37515 20700
tri 37515 20690 37525 20700 sw
tri 37251 20664 37277 20690 ne
rect 37277 20677 37525 20690
tri 37525 20677 37538 20690 sw
rect 37277 20668 37538 20677
rect 37277 20664 37410 20668
tri 37277 20619 37322 20664 ne
rect 37322 20622 37410 20664
rect 37456 20664 37538 20668
tri 37538 20664 37551 20677 sw
rect 70802 20670 70824 20716
rect 70870 20670 70928 20716
rect 70974 20670 71000 20716
rect 37456 20622 37551 20664
rect 37322 20619 37551 20622
tri 37551 20619 37596 20664 sw
tri 37322 20613 37328 20619 ne
rect 37328 20613 37596 20619
tri 37328 20600 37341 20613 ne
rect 37341 20600 37596 20613
tri 37596 20600 37615 20619 sw
rect 70802 20612 71000 20670
tri 37341 20568 37373 20600 ne
rect 37373 20590 37615 20600
tri 37615 20590 37625 20600 sw
rect 37373 20568 37625 20590
tri 37373 20523 37418 20568 ne
rect 37418 20558 37625 20568
tri 37625 20558 37657 20590 sw
rect 70802 20566 70824 20612
rect 70870 20566 70928 20612
rect 70974 20566 71000 20612
rect 37418 20545 37657 20558
tri 37657 20545 37670 20558 sw
rect 37418 20536 37670 20545
rect 37418 20523 37542 20536
tri 37418 20481 37460 20523 ne
rect 37460 20490 37542 20523
rect 37588 20513 37670 20536
tri 37670 20513 37702 20545 sw
rect 37588 20490 37702 20513
rect 37460 20481 37702 20490
tri 37460 20436 37505 20481 ne
rect 37505 20468 37702 20481
tri 37702 20468 37747 20513 sw
rect 70802 20508 71000 20566
rect 37505 20458 37747 20468
tri 37747 20458 37757 20468 sw
rect 70802 20462 70824 20508
rect 70870 20462 70928 20508
rect 70974 20462 71000 20508
rect 37505 20436 37757 20458
tri 37505 20425 37515 20436 ne
rect 37515 20426 37757 20436
tri 37757 20426 37789 20458 sw
rect 37515 20425 37789 20426
tri 37789 20425 37790 20426 sw
tri 37515 20380 37561 20425 ne
rect 37561 20413 37790 20425
tri 37790 20413 37802 20425 sw
rect 37561 20404 37802 20413
rect 37561 20380 37674 20404
tri 37561 20349 37592 20380 ne
rect 37592 20358 37674 20380
rect 37720 20381 37802 20404
tri 37802 20381 37834 20413 sw
rect 70802 20404 71000 20462
rect 37720 20358 37834 20381
rect 37592 20349 37834 20358
tri 37592 20336 37605 20349 ne
rect 37605 20336 37834 20349
tri 37834 20336 37879 20381 sw
rect 70802 20358 70824 20404
rect 70870 20358 70928 20404
rect 70974 20358 71000 20404
tri 37605 20304 37637 20336 ne
rect 37637 20326 37879 20336
tri 37879 20326 37889 20336 sw
rect 37637 20304 37889 20326
tri 37637 20299 37641 20304 ne
rect 37641 20299 37889 20304
tri 37641 20294 37647 20299 ne
rect 37647 20294 37889 20299
tri 37889 20294 37921 20326 sw
rect 70802 20300 71000 20358
tri 37647 20254 37687 20294 ne
rect 37687 20281 37921 20294
tri 37921 20281 37934 20294 sw
rect 37687 20272 37934 20281
rect 37687 20254 37806 20272
tri 37687 20217 37724 20254 ne
rect 37724 20226 37806 20254
rect 37852 20254 37934 20272
tri 37934 20254 37961 20281 sw
rect 70802 20254 70824 20300
rect 70870 20254 70928 20300
rect 70974 20254 71000 20300
rect 37852 20226 37961 20254
rect 37724 20217 37961 20226
tri 37724 20204 37737 20217 ne
rect 37737 20209 37961 20217
tri 37961 20209 38006 20254 sw
rect 37737 20204 38006 20209
tri 38006 20204 38011 20209 sw
tri 37737 20172 37769 20204 ne
rect 37769 20194 38011 20204
tri 38011 20194 38021 20204 sw
rect 70802 20196 71000 20254
rect 37769 20172 38021 20194
tri 37769 20151 37790 20172 ne
rect 37790 20162 38021 20172
tri 38021 20162 38053 20194 sw
rect 37790 20151 38053 20162
tri 38053 20151 38064 20162 sw
tri 37790 20106 37835 20151 ne
rect 37835 20149 38064 20151
tri 38064 20149 38066 20151 sw
rect 70802 20150 70824 20196
rect 70870 20150 70928 20196
rect 70974 20150 71000 20196
rect 37835 20140 38066 20149
rect 37835 20106 37938 20140
tri 37835 20085 37856 20106 ne
rect 37856 20094 37938 20106
rect 37984 20117 38066 20140
tri 38066 20117 38098 20149 sw
rect 37984 20094 38098 20117
rect 37856 20085 38098 20094
tri 37856 20072 37869 20085 ne
rect 37869 20072 38098 20085
tri 38098 20072 38143 20117 sw
rect 70802 20092 71000 20150
tri 37869 20040 37901 20072 ne
rect 37901 20062 38143 20072
tri 38143 20062 38153 20072 sw
rect 37901 20040 38153 20062
tri 37901 20030 37911 20040 ne
rect 37911 20030 38153 20040
tri 38153 20030 38185 20062 sw
rect 70802 20046 70824 20092
rect 70870 20046 70928 20092
rect 70974 20046 71000 20092
tri 37911 19985 37956 20030 ne
rect 37956 20017 38185 20030
tri 38185 20017 38198 20030 sw
rect 37956 20008 38198 20017
rect 37956 19985 38070 20008
tri 37956 19940 38001 19985 ne
rect 38001 19962 38070 19985
rect 38116 19985 38198 20008
tri 38198 19985 38230 20017 sw
rect 70802 19988 71000 20046
rect 38116 19962 38230 19985
rect 38001 19940 38230 19962
tri 38230 19940 38275 19985 sw
rect 70802 19942 70824 19988
rect 70870 19942 70928 19988
rect 70974 19942 71000 19988
tri 38001 19935 38006 19940 ne
rect 38006 19935 38275 19940
tri 38006 19889 38051 19935 ne
rect 38051 19930 38275 19935
tri 38275 19930 38285 19940 sw
rect 38051 19898 38285 19930
tri 38285 19898 38317 19930 sw
rect 38051 19889 38317 19898
tri 38317 19889 38326 19898 sw
tri 38051 19877 38064 19889 ne
rect 38064 19877 38326 19889
tri 38326 19877 38339 19889 sw
rect 70802 19884 71000 19942
tri 38064 19831 38109 19877 ne
rect 38109 19876 38339 19877
rect 38109 19831 38202 19876
tri 38109 19821 38120 19831 ne
rect 38120 19830 38202 19831
rect 38248 19844 38339 19876
tri 38339 19844 38371 19877 sw
rect 38248 19830 38371 19844
rect 38120 19821 38371 19830
tri 38120 19808 38133 19821 ne
rect 38133 19808 38371 19821
tri 38371 19808 38407 19844 sw
rect 70802 19838 70824 19884
rect 70870 19838 70928 19884
rect 70974 19838 71000 19884
tri 38133 19776 38165 19808 ne
rect 38165 19798 38407 19808
tri 38407 19798 38417 19808 sw
rect 38165 19776 38417 19798
tri 38165 19766 38175 19776 ne
rect 38175 19766 38417 19776
tri 38417 19766 38449 19798 sw
rect 70802 19780 71000 19838
tri 38175 19721 38220 19766 ne
rect 38220 19753 38449 19766
tri 38449 19753 38462 19766 sw
rect 38220 19744 38462 19753
rect 38220 19721 38334 19744
tri 38220 19689 38252 19721 ne
rect 38252 19698 38334 19721
rect 38380 19721 38462 19744
tri 38462 19721 38494 19753 sw
rect 70802 19734 70824 19780
rect 70870 19734 70928 19780
rect 70974 19734 71000 19780
rect 38380 19698 38494 19721
rect 38252 19689 38494 19698
tri 38252 19676 38265 19689 ne
rect 38265 19676 38494 19689
tri 38494 19676 38539 19721 sw
rect 70802 19676 71000 19734
tri 38265 19644 38297 19676 ne
rect 38297 19666 38539 19676
tri 38539 19666 38549 19676 sw
rect 38297 19644 38549 19666
tri 38297 19602 38339 19644 ne
rect 38339 19634 38549 19644
tri 38549 19634 38581 19666 sw
rect 38339 19621 38581 19634
tri 38581 19621 38594 19634 sw
rect 70802 19630 70824 19676
rect 70870 19630 70928 19676
rect 70974 19630 71000 19676
rect 38339 19612 38594 19621
rect 38339 19602 38466 19612
tri 38339 19570 38371 19602 ne
rect 38371 19570 38466 19602
tri 38371 19544 38397 19570 ne
rect 38397 19566 38466 19570
rect 38512 19602 38594 19612
tri 38594 19602 38613 19621 sw
rect 38512 19589 38613 19602
tri 38613 19589 38626 19602 sw
rect 38512 19566 38626 19589
rect 38397 19544 38626 19566
tri 38626 19544 38671 19589 sw
rect 70802 19572 71000 19630
tri 38397 19512 38429 19544 ne
rect 38429 19534 38671 19544
tri 38671 19534 38681 19544 sw
rect 38429 19512 38681 19534
tri 38429 19502 38439 19512 ne
rect 38439 19502 38681 19512
tri 38681 19502 38713 19534 sw
rect 70802 19526 70824 19572
rect 70870 19526 70928 19572
rect 70974 19526 71000 19572
tri 38439 19457 38484 19502 ne
rect 38484 19480 38713 19502
rect 38484 19457 38598 19480
tri 38484 19425 38516 19457 ne
rect 38516 19434 38598 19457
rect 38644 19479 38713 19480
tri 38713 19479 38736 19502 sw
rect 38644 19457 38736 19479
tri 38736 19457 38758 19479 sw
rect 70802 19468 71000 19526
rect 38644 19434 38758 19457
rect 38516 19425 38758 19434
tri 38516 19412 38529 19425 ne
rect 38529 19412 38758 19425
tri 38758 19412 38803 19457 sw
rect 70802 19422 70824 19468
rect 70870 19422 70928 19468
rect 70974 19422 71000 19468
tri 38529 19380 38561 19412 ne
rect 38561 19402 38803 19412
tri 38803 19402 38813 19412 sw
rect 38561 19380 38813 19402
tri 38561 19335 38606 19380 ne
rect 38606 19370 38813 19380
tri 38813 19370 38845 19402 sw
rect 38606 19357 38845 19370
tri 38845 19357 38858 19370 sw
rect 70802 19364 71000 19422
rect 38606 19348 38858 19357
rect 38606 19335 38730 19348
tri 38606 19328 38613 19335 ne
rect 38613 19328 38730 19335
tri 38613 19293 38648 19328 ne
rect 38648 19302 38730 19328
rect 38776 19328 38858 19348
tri 38858 19328 38887 19357 sw
rect 38776 19325 38887 19328
tri 38887 19325 38890 19328 sw
rect 38776 19302 38890 19325
rect 38648 19293 38890 19302
tri 38648 19280 38661 19293 ne
rect 38661 19280 38890 19293
tri 38890 19280 38935 19325 sw
rect 70802 19318 70824 19364
rect 70870 19318 70928 19364
rect 70974 19318 71000 19364
tri 38661 19248 38693 19280 ne
rect 38693 19270 38935 19280
tri 38935 19270 38945 19280 sw
rect 38693 19248 38945 19270
tri 38693 19238 38703 19248 ne
rect 38703 19238 38945 19248
tri 38945 19238 38977 19270 sw
rect 70802 19260 71000 19318
tri 38703 19205 38736 19238 ne
rect 38736 19225 38977 19238
tri 38977 19225 38990 19238 sw
rect 38736 19216 38990 19225
rect 38736 19205 38862 19216
tri 38736 19160 38781 19205 ne
rect 38781 19170 38862 19205
rect 38908 19205 38990 19216
tri 38990 19205 39010 19225 sw
rect 70802 19214 70824 19260
rect 70870 19214 70928 19260
rect 70974 19214 71000 19260
rect 38908 19170 39010 19205
rect 38781 19160 39010 19170
tri 39010 19160 39055 19205 sw
tri 38781 19148 38793 19160 ne
rect 38793 19148 39055 19160
tri 39055 19148 39067 19160 sw
rect 70802 19156 71000 19214
tri 38793 19116 38825 19148 ne
rect 38825 19138 39067 19148
tri 39067 19138 39077 19148 sw
rect 38825 19116 39077 19138
tri 38825 19071 38870 19116 ne
rect 38870 19106 39077 19116
tri 39077 19106 39109 19138 sw
rect 70802 19110 70824 19156
rect 70870 19110 70928 19156
rect 70974 19110 71000 19156
rect 38870 19093 39109 19106
tri 39109 19093 39122 19106 sw
rect 38870 19084 39122 19093
rect 38870 19071 38994 19084
tri 38870 19053 38887 19071 ne
rect 38887 19053 38994 19071
tri 38887 19029 38912 19053 ne
rect 38912 19038 38994 19053
rect 39040 19053 39122 19084
tri 39122 19053 39162 19093 sw
rect 39040 19038 39162 19053
rect 38912 19029 39162 19038
tri 38912 19016 38925 19029 ne
rect 38925 19016 39162 19029
tri 39162 19016 39199 19053 sw
rect 70802 19052 71000 19110
tri 38925 18984 38957 19016 ne
rect 38957 19006 39199 19016
tri 39199 19006 39209 19016 sw
rect 70802 19006 70824 19052
rect 70870 19006 70928 19052
rect 70974 19006 71000 19052
rect 38957 18984 39209 19006
tri 38957 18974 38967 18984 ne
rect 38967 18974 39209 18984
tri 39209 18974 39241 19006 sw
tri 38967 18929 39012 18974 ne
rect 39012 18961 39241 18974
tri 39241 18961 39254 18974 sw
rect 39012 18952 39254 18961
rect 39012 18929 39126 18952
tri 39012 18897 39044 18929 ne
rect 39044 18906 39126 18929
rect 39172 18929 39254 18952
tri 39254 18929 39286 18961 sw
rect 70802 18948 71000 19006
rect 39172 18906 39286 18929
rect 39044 18897 39286 18906
tri 39044 18884 39057 18897 ne
rect 39057 18884 39286 18897
tri 39286 18884 39331 18929 sw
rect 70802 18902 70824 18948
rect 70870 18902 70928 18948
rect 70974 18902 71000 18948
tri 39057 18852 39089 18884 ne
rect 39089 18874 39331 18884
tri 39331 18874 39341 18884 sw
rect 39089 18852 39341 18874
tri 39089 18840 39101 18852 ne
rect 39101 18842 39341 18852
tri 39341 18842 39373 18874 sw
rect 70802 18844 71000 18902
rect 39101 18840 39373 18842
tri 39101 18795 39146 18840 ne
rect 39146 18829 39373 18840
tri 39373 18829 39386 18842 sw
rect 39146 18820 39386 18829
rect 39146 18795 39258 18820
tri 39146 18779 39162 18795 ne
rect 39162 18779 39258 18795
tri 39162 18765 39176 18779 ne
rect 39176 18774 39258 18779
rect 39304 18795 39386 18820
tri 39386 18795 39420 18829 sw
rect 70802 18798 70824 18844
rect 70870 18798 70928 18844
rect 70974 18798 71000 18844
rect 39304 18779 39420 18795
tri 39420 18779 39436 18795 sw
rect 39304 18774 39436 18779
rect 39176 18765 39436 18774
tri 39176 18752 39189 18765 ne
rect 39189 18752 39436 18765
tri 39436 18752 39463 18779 sw
tri 39189 18720 39221 18752 ne
rect 39221 18750 39463 18752
tri 39463 18750 39465 18752 sw
rect 39221 18742 39465 18750
tri 39465 18742 39473 18750 sw
rect 39221 18720 39473 18742
tri 39221 18710 39231 18720 ne
rect 39231 18710 39473 18720
tri 39473 18710 39505 18742 sw
rect 70802 18740 71000 18798
tri 39231 18665 39276 18710 ne
rect 39276 18697 39505 18710
tri 39505 18697 39518 18710 sw
rect 39276 18688 39518 18697
rect 39276 18665 39390 18688
tri 39276 18633 39308 18665 ne
rect 39308 18642 39390 18665
rect 39436 18665 39518 18688
tri 39518 18665 39550 18697 sw
rect 70802 18694 70824 18740
rect 70870 18694 70928 18740
rect 70974 18694 71000 18740
rect 39436 18642 39550 18665
rect 39308 18633 39550 18642
tri 39308 18620 39321 18633 ne
rect 39321 18620 39550 18633
tri 39550 18620 39595 18665 sw
rect 70802 18636 71000 18694
tri 39321 18588 39353 18620 ne
rect 39353 18610 39595 18620
tri 39595 18610 39605 18620 sw
rect 39353 18588 39605 18610
tri 39353 18543 39398 18588 ne
rect 39398 18578 39605 18588
tri 39605 18578 39637 18610 sw
rect 70802 18590 70824 18636
rect 70870 18590 70928 18636
rect 70974 18590 71000 18636
rect 39398 18565 39637 18578
tri 39637 18565 39650 18578 sw
rect 39398 18556 39650 18565
rect 39398 18543 39522 18556
tri 39398 18505 39436 18543 ne
rect 39436 18510 39522 18543
rect 39568 18550 39650 18556
tri 39650 18550 39665 18565 sw
rect 39568 18510 39665 18550
rect 39436 18505 39665 18510
tri 39665 18505 39711 18550 sw
rect 70802 18532 71000 18590
tri 39436 18488 39453 18505 ne
rect 39453 18488 39711 18505
tri 39711 18488 39727 18505 sw
tri 39453 18475 39465 18488 ne
rect 39465 18478 39727 18488
tri 39727 18478 39737 18488 sw
rect 70802 18486 70824 18532
rect 70870 18486 70928 18532
rect 70974 18486 71000 18532
rect 39465 18475 39737 18478
tri 39465 18446 39495 18475 ne
rect 39495 18446 39737 18475
tri 39737 18446 39769 18478 sw
tri 39495 18430 39511 18446 ne
rect 39511 18433 39769 18446
tri 39769 18433 39782 18446 sw
rect 39511 18430 39782 18433
tri 39782 18430 39785 18433 sw
tri 39511 18385 39556 18430 ne
rect 39556 18424 39785 18430
rect 39556 18385 39654 18424
tri 39556 18369 39572 18385 ne
rect 39572 18378 39654 18385
rect 39700 18385 39785 18424
tri 39785 18385 39830 18430 sw
rect 70802 18428 71000 18486
rect 39700 18378 39830 18385
rect 39572 18369 39830 18378
tri 39572 18356 39585 18369 ne
rect 39585 18356 39830 18369
tri 39830 18356 39859 18385 sw
rect 70802 18382 70824 18428
rect 70870 18382 70928 18428
rect 70974 18382 71000 18428
tri 39585 18324 39617 18356 ne
rect 39617 18346 39859 18356
tri 39859 18346 39869 18356 sw
rect 39617 18324 39869 18346
tri 39617 18279 39662 18324 ne
rect 39662 18314 39869 18324
tri 39869 18314 39901 18346 sw
rect 70802 18324 71000 18382
rect 39662 18301 39901 18314
tri 39901 18301 39914 18314 sw
rect 39662 18292 39914 18301
rect 39662 18279 39786 18292
tri 39662 18237 39704 18279 ne
rect 39704 18246 39786 18279
rect 39832 18275 39914 18292
tri 39914 18275 39940 18301 sw
rect 70802 18278 70824 18324
rect 70870 18278 70928 18324
rect 70974 18278 71000 18324
rect 39832 18246 39940 18275
rect 39704 18237 39940 18246
tri 39704 18230 39711 18237 ne
rect 39711 18230 39940 18237
tri 39940 18230 39985 18275 sw
tri 39711 18224 39717 18230 ne
rect 39717 18224 39985 18230
tri 39985 18224 39991 18230 sw
tri 39717 18192 39749 18224 ne
rect 39749 18214 39991 18224
tri 39991 18214 40001 18224 sw
rect 70802 18220 71000 18278
rect 39749 18192 40001 18214
tri 39749 18182 39759 18192 ne
rect 39759 18182 40001 18192
tri 40001 18182 40033 18214 sw
tri 39759 18137 39804 18182 ne
rect 39804 18169 40033 18182
tri 40033 18169 40046 18182 sw
rect 70802 18174 70824 18220
rect 70870 18174 70928 18220
rect 70974 18174 71000 18220
rect 39804 18160 40046 18169
rect 39804 18137 39918 18160
tri 39804 18111 39830 18137 ne
rect 39830 18114 39918 18137
rect 39964 18137 40046 18160
tri 40046 18137 40078 18169 sw
rect 39964 18114 40078 18137
rect 39830 18111 40078 18114
tri 39830 18092 39849 18111 ne
rect 39849 18092 40078 18111
tri 40078 18092 40123 18137 sw
rect 70802 18116 71000 18174
tri 39849 18060 39881 18092 ne
rect 39881 18082 40123 18092
tri 40123 18082 40133 18092 sw
rect 39881 18060 40133 18082
tri 39881 18015 39926 18060 ne
rect 39926 18050 40133 18060
tri 40133 18050 40165 18082 sw
rect 70802 18070 70824 18116
rect 70870 18070 70928 18116
rect 70974 18070 71000 18116
rect 39926 18028 40165 18050
rect 39926 18015 40050 18028
tri 39926 17973 39968 18015 ne
rect 39968 17982 40050 18015
rect 40096 18020 40165 18028
tri 40165 18020 40195 18050 sw
rect 40096 18005 40195 18020
tri 40195 18005 40210 18020 sw
rect 70802 18012 71000 18070
rect 40096 17982 40210 18005
rect 39968 17973 40210 17982
tri 39968 17956 39985 17973 ne
rect 39985 17960 40210 17973
tri 40210 17960 40255 18005 sw
rect 70802 17966 70824 18012
rect 70870 17966 70928 18012
rect 70974 17966 71000 18012
rect 39985 17956 40255 17960
tri 40255 17956 40259 17960 sw
tri 39985 17928 40013 17956 ne
rect 40013 17950 40259 17956
tri 40259 17950 40265 17956 sw
rect 40013 17928 40265 17950
tri 40013 17918 40023 17928 ne
rect 40023 17918 40265 17928
tri 40265 17918 40297 17950 sw
tri 40023 17873 40068 17918 ne
rect 40068 17905 40297 17918
tri 40297 17905 40310 17918 sw
rect 70802 17908 71000 17966
rect 40068 17896 40310 17905
rect 40068 17873 40182 17896
tri 40068 17841 40100 17873 ne
rect 40100 17850 40182 17873
rect 40228 17873 40310 17896
tri 40310 17873 40342 17905 sw
rect 40228 17850 40342 17873
rect 40100 17841 40342 17850
tri 40100 17828 40113 17841 ne
rect 40113 17828 40342 17841
tri 40342 17828 40387 17873 sw
rect 70802 17862 70824 17908
rect 70870 17862 70928 17908
rect 70974 17862 71000 17908
tri 40113 17796 40145 17828 ne
rect 40145 17818 40387 17828
tri 40387 17818 40397 17828 sw
rect 40145 17796 40397 17818
tri 40145 17751 40190 17796 ne
rect 40190 17786 40397 17796
tri 40397 17786 40429 17818 sw
rect 70802 17804 71000 17862
rect 40190 17773 40429 17786
tri 40429 17773 40442 17786 sw
rect 40190 17764 40442 17773
rect 40190 17751 40314 17764
tri 40190 17746 40195 17751 ne
rect 40195 17746 40314 17751
tri 40195 17701 40240 17746 ne
rect 40240 17718 40314 17746
rect 40360 17746 40442 17764
tri 40442 17746 40469 17773 sw
rect 70802 17758 70824 17804
rect 70870 17758 70928 17804
rect 70974 17758 71000 17804
rect 40360 17718 40469 17746
rect 40240 17701 40469 17718
tri 40469 17701 40515 17746 sw
tri 40240 17681 40259 17701 ne
rect 40259 17696 40515 17701
tri 40515 17696 40519 17701 sw
rect 70802 17700 71000 17758
rect 40259 17681 40519 17696
tri 40519 17681 40534 17696 sw
tri 40259 17664 40277 17681 ne
rect 40277 17664 40534 17681
tri 40277 17654 40287 17664 ne
rect 40287 17654 40534 17664
tri 40534 17654 40561 17681 sw
rect 70802 17654 70824 17700
rect 70870 17654 70928 17700
rect 70974 17654 71000 17700
tri 40287 17609 40332 17654 ne
rect 40332 17641 40561 17654
tri 40561 17641 40574 17654 sw
rect 40332 17632 40574 17641
rect 40332 17609 40446 17632
tri 40332 17577 40364 17609 ne
rect 40364 17586 40446 17609
rect 40492 17609 40574 17632
tri 40574 17609 40606 17641 sw
rect 40492 17586 40606 17609
rect 40364 17577 40606 17586
tri 40364 17564 40377 17577 ne
rect 40377 17564 40606 17577
tri 40606 17564 40651 17609 sw
rect 70802 17596 71000 17654
tri 40377 17532 40409 17564 ne
rect 40409 17554 40651 17564
tri 40651 17554 40661 17564 sw
rect 40409 17532 40661 17554
tri 40409 17487 40454 17532 ne
rect 40454 17522 40661 17532
tri 40661 17522 40693 17554 sw
rect 70802 17550 70824 17596
rect 70870 17550 70928 17596
rect 70974 17550 71000 17596
rect 40454 17509 40693 17522
tri 40693 17509 40706 17522 sw
rect 40454 17500 40706 17509
rect 40454 17487 40578 17500
tri 40454 17445 40496 17487 ne
rect 40496 17454 40578 17487
rect 40624 17477 40706 17500
tri 40706 17477 40738 17509 sw
rect 70802 17492 71000 17550
rect 40624 17454 40738 17477
rect 40496 17445 40738 17454
tri 40496 17407 40534 17445 ne
rect 40534 17432 40738 17445
tri 40738 17432 40783 17477 sw
rect 70802 17446 70824 17492
rect 70870 17446 70928 17492
rect 70974 17446 71000 17492
rect 40534 17422 40783 17432
tri 40783 17422 40793 17432 sw
rect 40534 17407 40793 17422
tri 40793 17407 40808 17422 sw
tri 40534 17400 40541 17407 ne
rect 40541 17400 40808 17407
tri 40541 17390 40551 17400 ne
rect 40551 17390 40808 17400
tri 40808 17390 40825 17407 sw
tri 40551 17381 40560 17390 ne
rect 40560 17381 40825 17390
tri 40560 17336 40605 17381 ne
rect 40605 17377 40825 17381
tri 40825 17377 40838 17390 sw
rect 70802 17388 71000 17446
rect 40605 17368 40838 17377
rect 40605 17336 40710 17368
tri 40605 17313 40628 17336 ne
rect 40628 17322 40710 17336
rect 40756 17336 40838 17368
tri 40838 17336 40879 17377 sw
rect 70802 17342 70824 17388
rect 70870 17342 70928 17388
rect 70974 17342 71000 17388
rect 40756 17322 40879 17336
rect 40628 17313 40879 17322
tri 40628 17300 40641 17313 ne
rect 40641 17300 40879 17313
tri 40879 17300 40915 17336 sw
tri 40641 17268 40673 17300 ne
rect 40673 17291 40915 17300
tri 40915 17291 40925 17300 sw
rect 40673 17268 40925 17291
tri 40673 17223 40718 17268 ne
rect 40718 17258 40925 17268
tri 40925 17258 40957 17290 sw
rect 70802 17284 71000 17342
rect 40718 17245 40957 17258
tri 40957 17245 40970 17258 sw
rect 40718 17236 40970 17245
rect 40718 17223 40842 17236
tri 40718 17181 40760 17223 ne
rect 40760 17190 40842 17223
rect 40888 17213 40970 17236
tri 40970 17213 41002 17245 sw
rect 70802 17238 70824 17284
rect 70870 17238 70928 17284
rect 70974 17238 71000 17284
rect 40888 17190 41002 17213
rect 40760 17181 41002 17190
tri 40760 17136 40805 17181 ne
rect 40805 17168 41002 17181
tri 41002 17168 41047 17213 sw
rect 70802 17180 71000 17238
rect 40805 17158 41047 17168
tri 41047 17158 41057 17168 sw
rect 40805 17136 41057 17158
tri 40805 17133 40808 17136 ne
rect 40808 17133 41057 17136
tri 41057 17133 41083 17158 sw
rect 70802 17134 70824 17180
rect 70870 17134 70928 17180
rect 70974 17134 71000 17180
tri 40808 17126 40815 17133 ne
rect 40815 17126 41083 17133
tri 41083 17126 41089 17133 sw
tri 40815 17081 40860 17126 ne
rect 40860 17113 41089 17126
tri 41089 17113 41102 17126 sw
rect 40860 17104 41102 17113
rect 40860 17081 40974 17104
tri 40860 17049 40892 17081 ne
rect 40892 17058 40974 17081
rect 41020 17081 41102 17104
tri 41102 17081 41134 17113 sw
rect 41020 17058 41134 17081
rect 40892 17049 41134 17058
tri 40892 17036 40905 17049 ne
rect 40905 17036 41134 17049
tri 41134 17036 41179 17081 sw
rect 70802 17076 71000 17134
tri 40905 17004 40937 17036 ne
rect 40937 17026 41179 17036
tri 41179 17026 41189 17036 sw
rect 70802 17030 70824 17076
rect 70870 17030 70928 17076
rect 70974 17030 71000 17076
rect 40937 17004 41189 17026
tri 40937 16971 40970 17004 ne
rect 40970 16994 41189 17004
tri 41189 16994 41221 17026 sw
rect 40970 16981 41221 16994
tri 41221 16981 41234 16994 sw
rect 40970 16972 41234 16981
rect 40970 16971 41106 16972
tri 40970 16926 41015 16971 ne
rect 41015 16926 41106 16971
rect 41152 16971 41234 16972
tri 41234 16971 41244 16981 sw
rect 70802 16972 71000 17030
rect 41152 16926 41244 16971
tri 41244 16926 41289 16971 sw
rect 70802 16926 70824 16972
rect 70870 16926 70928 16972
rect 70974 16926 71000 16972
tri 41015 16917 41024 16926 ne
rect 41024 16917 41289 16926
tri 41024 16872 41069 16917 ne
rect 41069 16904 41289 16917
tri 41289 16904 41311 16926 sw
rect 41069 16894 41311 16904
tri 41311 16894 41321 16904 sw
rect 41069 16872 41321 16894
tri 41069 16858 41083 16872 ne
rect 41083 16862 41321 16872
tri 41321 16862 41353 16894 sw
rect 70802 16868 71000 16926
rect 41083 16858 41353 16862
tri 41353 16858 41357 16862 sw
tri 41083 16813 41128 16858 ne
rect 41128 16849 41357 16858
tri 41357 16849 41366 16858 sw
rect 41128 16840 41366 16849
rect 41128 16813 41238 16840
tri 41128 16785 41156 16813 ne
rect 41156 16794 41238 16813
rect 41284 16817 41366 16840
tri 41366 16817 41398 16849 sw
rect 70802 16822 70824 16868
rect 70870 16822 70928 16868
rect 70974 16822 71000 16868
rect 41284 16794 41398 16817
rect 41156 16785 41398 16794
tri 41156 16772 41169 16785 ne
rect 41169 16772 41398 16785
tri 41398 16772 41443 16817 sw
tri 41169 16740 41201 16772 ne
rect 41201 16762 41443 16772
tri 41443 16762 41453 16772 sw
rect 70802 16764 71000 16822
rect 41201 16740 41453 16762
tri 41201 16730 41211 16740 ne
rect 41211 16730 41453 16740
tri 41453 16730 41485 16762 sw
tri 41211 16685 41256 16730 ne
rect 41256 16717 41485 16730
tri 41485 16717 41498 16730 sw
rect 70802 16718 70824 16764
rect 70870 16718 70928 16764
rect 70974 16718 71000 16764
rect 41256 16708 41498 16717
rect 41256 16685 41370 16708
tri 41256 16651 41289 16685 ne
rect 41289 16662 41370 16685
rect 41416 16685 41498 16708
tri 41498 16685 41530 16717 sw
rect 41416 16662 41530 16685
rect 41289 16651 41530 16662
tri 41289 16640 41301 16651 ne
rect 41301 16640 41530 16651
tri 41530 16640 41575 16685 sw
rect 70802 16660 71000 16718
tri 41301 16606 41335 16640 ne
rect 41335 16630 41575 16640
tri 41575 16630 41585 16640 sw
rect 41335 16606 41585 16630
tri 41335 16584 41357 16606 ne
rect 41357 16598 41585 16606
tri 41585 16598 41617 16630 sw
rect 70802 16614 70824 16660
rect 70870 16614 70928 16660
rect 70974 16614 71000 16660
rect 41357 16584 41617 16598
tri 41617 16584 41631 16598 sw
tri 41357 16539 41402 16584 ne
rect 41402 16576 41631 16584
rect 41402 16539 41502 16576
tri 41402 16521 41420 16539 ne
rect 41420 16530 41502 16539
rect 41548 16561 41631 16576
tri 41631 16561 41654 16584 sw
rect 41548 16553 41654 16561
tri 41654 16553 41662 16561 sw
rect 70802 16556 71000 16614
rect 41548 16530 41662 16553
rect 41420 16521 41662 16530
tri 41420 16508 41433 16521 ne
rect 41433 16508 41662 16521
tri 41662 16508 41707 16553 sw
rect 70802 16510 70824 16556
rect 70870 16510 70928 16556
rect 70974 16510 71000 16556
tri 41433 16476 41465 16508 ne
rect 41465 16498 41707 16508
tri 41707 16498 41717 16508 sw
rect 41465 16476 41717 16498
tri 41465 16466 41475 16476 ne
rect 41475 16466 41717 16476
tri 41717 16466 41749 16498 sw
tri 41475 16421 41520 16466 ne
rect 41520 16453 41749 16466
tri 41749 16453 41762 16466 sw
rect 41520 16444 41762 16453
rect 41520 16421 41634 16444
tri 41520 16389 41552 16421 ne
rect 41552 16398 41634 16421
rect 41680 16421 41762 16444
tri 41762 16421 41794 16453 sw
rect 70802 16452 71000 16510
rect 41680 16398 41794 16421
rect 41552 16389 41794 16398
tri 41552 16376 41565 16389 ne
rect 41565 16376 41794 16389
tri 41794 16376 41839 16421 sw
rect 70802 16406 70824 16452
rect 70870 16406 70928 16452
rect 70974 16406 71000 16452
tri 41565 16344 41597 16376 ne
rect 41597 16366 41839 16376
tri 41839 16366 41849 16376 sw
rect 41597 16344 41849 16366
tri 41597 16309 41631 16344 ne
rect 41631 16334 41849 16344
tri 41849 16334 41881 16366 sw
rect 70802 16348 71000 16406
rect 41631 16321 41881 16334
tri 41881 16321 41894 16334 sw
rect 41631 16312 41894 16321
rect 41631 16309 41766 16312
tri 41631 16287 41654 16309 ne
rect 41654 16287 41766 16309
tri 41654 16244 41697 16287 ne
rect 41697 16266 41766 16287
rect 41812 16309 41894 16312
tri 41894 16309 41906 16321 sw
rect 41812 16289 41906 16309
tri 41906 16289 41926 16309 sw
rect 70802 16302 70824 16348
rect 70870 16302 70928 16348
rect 70974 16302 71000 16348
rect 41812 16266 41926 16289
rect 41697 16244 41926 16266
tri 41926 16244 41971 16289 sw
rect 70802 16244 71000 16302
tri 41697 16212 41729 16244 ne
rect 41729 16241 41971 16244
tri 41971 16241 41974 16244 sw
rect 41729 16212 41974 16241
tri 41729 16202 41739 16212 ne
rect 41739 16202 41974 16212
tri 41974 16202 42013 16241 sw
tri 41739 16157 41784 16202 ne
rect 41784 16189 42013 16202
tri 42013 16189 42026 16202 sw
rect 70802 16198 70824 16244
rect 70870 16198 70928 16244
rect 70974 16198 71000 16244
rect 41784 16180 42026 16189
rect 41784 16157 41898 16180
tri 41784 16125 41816 16157 ne
rect 41816 16134 41898 16157
rect 41944 16157 42026 16180
tri 42026 16157 42058 16189 sw
rect 41944 16134 42058 16157
rect 41816 16125 42058 16134
tri 41816 16112 41829 16125 ne
rect 41829 16112 42058 16125
tri 42058 16112 42103 16157 sw
rect 70802 16140 71000 16198
tri 41829 16080 41861 16112 ne
rect 41861 16102 42103 16112
tri 42103 16102 42113 16112 sw
rect 41861 16080 42113 16102
tri 41861 16035 41906 16080 ne
rect 41906 16070 42113 16080
tri 42113 16070 42145 16102 sw
rect 70802 16094 70824 16140
rect 70870 16094 70928 16140
rect 70974 16094 71000 16140
rect 41906 16057 42145 16070
tri 42145 16057 42158 16070 sw
rect 41906 16048 42158 16057
rect 41906 16035 42030 16048
tri 41906 15993 41948 16035 ne
rect 41948 16002 42030 16035
rect 42076 16035 42158 16048
tri 42158 16035 42180 16057 sw
rect 70802 16036 71000 16094
rect 42076 16025 42180 16035
tri 42180 16025 42190 16035 sw
rect 42076 16002 42190 16025
rect 41948 15993 42190 16002
tri 41948 15980 41961 15993 ne
rect 41961 15980 42190 15993
tri 42190 15980 42235 16025 sw
rect 70802 15990 70824 16036
rect 70870 15990 70928 16036
rect 70974 15990 71000 16036
tri 41961 15948 41993 15980 ne
rect 41993 15970 42235 15980
tri 42235 15970 42245 15980 sw
rect 41993 15948 42245 15970
tri 41993 15938 42003 15948 ne
rect 42003 15938 42245 15948
tri 42245 15938 42277 15970 sw
tri 42003 15922 42019 15938 ne
rect 42019 15925 42277 15938
tri 42277 15925 42290 15938 sw
rect 70802 15932 71000 15990
rect 42019 15922 42290 15925
tri 42290 15922 42293 15925 sw
tri 42019 15877 42064 15922 ne
rect 42064 15916 42293 15922
rect 42064 15877 42162 15916
tri 42064 15861 42080 15877 ne
rect 42080 15870 42162 15877
rect 42208 15877 42293 15916
tri 42293 15877 42339 15922 sw
rect 70802 15886 70824 15932
rect 70870 15886 70928 15932
rect 70974 15886 71000 15932
rect 42208 15870 42339 15877
rect 42080 15861 42339 15870
tri 42080 15848 42093 15861 ne
rect 42093 15848 42339 15861
tri 42339 15848 42367 15877 sw
tri 42093 15816 42125 15848 ne
rect 42125 15838 42367 15848
tri 42367 15838 42377 15848 sw
rect 42125 15816 42377 15838
tri 42125 15771 42170 15816 ne
rect 42170 15806 42377 15816
tri 42377 15806 42409 15838 sw
rect 70802 15828 71000 15886
rect 42170 15793 42409 15806
tri 42409 15793 42422 15806 sw
rect 42170 15784 42422 15793
rect 42170 15771 42294 15784
tri 42170 15761 42180 15771 ne
rect 42180 15761 42294 15771
tri 42180 15729 42212 15761 ne
rect 42212 15738 42294 15761
rect 42340 15761 42422 15784
tri 42422 15761 42455 15793 sw
rect 70802 15782 70824 15828
rect 70870 15782 70928 15828
rect 70974 15782 71000 15828
rect 42340 15738 42455 15761
rect 42212 15729 42455 15738
tri 42212 15716 42225 15729 ne
rect 42225 15716 42455 15729
tri 42455 15716 42499 15761 sw
rect 70802 15724 71000 15782
tri 42225 15684 42257 15716 ne
rect 42257 15706 42499 15716
tri 42499 15706 42509 15716 sw
rect 42257 15684 42509 15706
tri 42257 15674 42267 15684 ne
rect 42267 15674 42509 15684
tri 42509 15674 42541 15706 sw
rect 70802 15678 70824 15724
rect 70870 15678 70928 15724
rect 70974 15678 71000 15724
tri 42267 15629 42312 15674 ne
rect 42312 15661 42541 15674
tri 42541 15661 42554 15674 sw
rect 42312 15652 42554 15661
rect 42312 15629 42426 15652
tri 42312 15597 42344 15629 ne
rect 42344 15606 42426 15629
rect 42472 15629 42554 15652
tri 42554 15629 42586 15661 sw
rect 42472 15606 42586 15629
rect 42344 15597 42586 15606
tri 42344 15584 42357 15597 ne
rect 42357 15584 42586 15597
tri 42586 15584 42631 15629 sw
rect 70802 15620 71000 15678
tri 42357 15552 42389 15584 ne
rect 42389 15574 42631 15584
tri 42631 15574 42641 15584 sw
rect 70802 15574 70824 15620
rect 70870 15574 70928 15620
rect 70974 15574 71000 15620
rect 42389 15552 42641 15574
tri 42389 15512 42429 15552 ne
rect 42429 15542 42641 15552
tri 42641 15542 42673 15574 sw
rect 42429 15529 42673 15542
tri 42673 15529 42686 15542 sw
rect 42429 15520 42686 15529
rect 42429 15512 42558 15520
tri 42429 15486 42455 15512 ne
rect 42455 15486 42558 15512
tri 42455 15465 42476 15486 ne
rect 42476 15474 42558 15486
rect 42604 15512 42686 15520
tri 42686 15512 42703 15529 sw
rect 70802 15516 71000 15574
rect 42604 15486 42703 15512
tri 42703 15486 42729 15512 sw
rect 42604 15474 42729 15486
rect 42476 15467 42729 15474
tri 42729 15467 42749 15486 sw
rect 70802 15470 70824 15516
rect 70870 15470 70928 15516
rect 70974 15470 71000 15516
rect 42476 15465 42749 15467
tri 42476 15452 42489 15465 ne
rect 42489 15452 42749 15465
tri 42749 15452 42763 15467 sw
tri 42489 15420 42521 15452 ne
rect 42521 15442 42763 15452
tri 42763 15442 42773 15452 sw
rect 42521 15420 42773 15442
tri 42521 15410 42531 15420 ne
rect 42531 15410 42773 15420
tri 42773 15410 42805 15442 sw
rect 70802 15412 71000 15470
tri 42531 15365 42576 15410 ne
rect 42576 15397 42805 15410
tri 42805 15397 42818 15410 sw
rect 42576 15388 42818 15397
rect 42576 15365 42690 15388
tri 42576 15333 42608 15365 ne
rect 42608 15342 42690 15365
rect 42736 15365 42818 15388
tri 42818 15365 42850 15397 sw
rect 70802 15366 70824 15412
rect 70870 15366 70928 15412
rect 70974 15366 71000 15412
rect 42736 15342 42850 15365
rect 42608 15333 42850 15342
tri 42608 15320 42621 15333 ne
rect 42621 15320 42850 15333
tri 42850 15320 42895 15365 sw
tri 42621 15288 42653 15320 ne
rect 42653 15310 42895 15320
tri 42895 15310 42905 15320 sw
rect 42653 15288 42905 15310
tri 42653 15243 42698 15288 ne
rect 42698 15278 42905 15288
tri 42905 15278 42937 15310 sw
rect 70802 15308 71000 15366
rect 42698 15265 42937 15278
tri 42937 15265 42950 15278 sw
rect 42698 15257 42950 15265
tri 42950 15257 42958 15265 sw
rect 70802 15262 70824 15308
rect 70870 15262 70928 15308
rect 70974 15262 71000 15308
rect 42698 15256 42958 15257
rect 42698 15243 42822 15256
tri 42698 15212 42729 15243 ne
rect 42729 15212 42822 15243
tri 42729 15192 42749 15212 ne
rect 42749 15210 42822 15212
rect 42868 15212 42958 15256
tri 42958 15212 43003 15257 sw
rect 42868 15210 43003 15212
rect 42749 15192 43003 15210
tri 42749 15188 42753 15192 ne
rect 42753 15188 43003 15192
tri 43003 15188 43027 15212 sw
rect 70802 15204 71000 15262
tri 42753 15147 42794 15188 ne
rect 42794 15178 43027 15188
tri 43027 15178 43037 15188 sw
rect 42794 15147 43037 15178
tri 42794 15146 42795 15147 ne
rect 42795 15146 43037 15147
tri 43037 15146 43069 15178 sw
rect 70802 15158 70824 15204
rect 70870 15158 70928 15204
rect 70974 15158 71000 15204
tri 42795 15101 42840 15146 ne
rect 42840 15124 43069 15146
rect 42840 15101 42954 15124
tri 42840 15069 42872 15101 ne
rect 42872 15078 42954 15101
rect 43000 15102 43069 15124
tri 43069 15102 43113 15146 sw
rect 43000 15101 43113 15102
tri 43113 15101 43114 15102 sw
rect 43000 15078 43114 15101
rect 42872 15069 43114 15078
tri 42872 15056 42885 15069 ne
rect 42885 15056 43114 15069
tri 43114 15056 43159 15101 sw
rect 70802 15100 71000 15158
tri 42885 15024 42917 15056 ne
rect 42917 15046 43159 15056
tri 43159 15046 43169 15056 sw
rect 70802 15054 70824 15100
rect 70870 15054 70928 15100
rect 70974 15054 71000 15100
rect 42917 15024 43169 15046
tri 42917 14979 42962 15024 ne
rect 42962 15014 43169 15024
tri 43169 15014 43201 15046 sw
rect 42962 15001 43201 15014
tri 43201 15001 43214 15014 sw
rect 42962 14992 43214 15001
rect 42962 14979 43086 14992
tri 42962 14937 43003 14979 ne
rect 43003 14946 43086 14979
rect 43132 14983 43214 14992
tri 43214 14983 43233 15001 sw
rect 70802 14996 71000 15054
rect 43132 14946 43233 14983
rect 43003 14937 43233 14946
tri 43233 14937 43278 14983 sw
rect 70802 14950 70824 14996
rect 70870 14950 70928 14996
rect 70974 14950 71000 14996
tri 43004 14924 43017 14937 ne
rect 43017 14924 43278 14937
tri 43278 14924 43291 14937 sw
tri 43017 14892 43049 14924 ne
rect 43049 14914 43291 14924
tri 43291 14914 43301 14924 sw
rect 43049 14892 43301 14914
tri 43049 14882 43059 14892 ne
rect 43059 14882 43301 14892
tri 43301 14882 43333 14914 sw
rect 70802 14892 71000 14950
tri 43059 14837 43104 14882 ne
rect 43104 14869 43333 14882
tri 43333 14869 43346 14882 sw
rect 43104 14860 43346 14869
rect 43104 14837 43218 14860
tri 43104 14827 43113 14837 ne
rect 43113 14827 43218 14837
tri 43113 14792 43149 14827 ne
rect 43149 14814 43218 14827
rect 43264 14837 43346 14860
tri 43346 14837 43378 14869 sw
rect 70802 14846 70824 14892
rect 70870 14846 70928 14892
rect 70974 14846 71000 14892
rect 43264 14814 43378 14837
rect 43149 14792 43378 14814
tri 43378 14792 43423 14837 sw
tri 43149 14760 43181 14792 ne
rect 43181 14782 43423 14792
tri 43423 14782 43433 14792 sw
rect 70802 14788 71000 14846
rect 43181 14760 43433 14782
tri 43181 14715 43226 14760 ne
rect 43226 14750 43433 14760
tri 43433 14750 43465 14782 sw
rect 43226 14737 43465 14750
tri 43465 14737 43478 14750 sw
rect 70802 14742 70824 14788
rect 70870 14742 70928 14788
rect 70974 14742 71000 14788
rect 43226 14728 43478 14737
rect 43226 14715 43350 14728
tri 43226 14673 43268 14715 ne
rect 43268 14682 43350 14715
rect 43396 14708 43478 14728
tri 43478 14708 43507 14737 sw
rect 43396 14682 43507 14708
rect 43268 14673 43507 14682
tri 43268 14663 43278 14673 ne
rect 43278 14663 43507 14673
tri 43507 14663 43552 14708 sw
rect 70802 14684 71000 14742
tri 43278 14660 43281 14663 ne
rect 43281 14660 43552 14663
tri 43552 14660 43555 14663 sw
tri 43281 14628 43313 14660 ne
rect 43313 14650 43555 14660
tri 43555 14650 43565 14660 sw
rect 43313 14628 43565 14650
tri 43313 14618 43323 14628 ne
rect 43323 14618 43565 14628
tri 43565 14618 43597 14650 sw
rect 70802 14638 70824 14684
rect 70870 14638 70928 14684
rect 70974 14638 71000 14684
tri 43323 14573 43368 14618 ne
rect 43368 14605 43597 14618
tri 43597 14605 43610 14618 sw
rect 43368 14596 43610 14605
rect 43368 14573 43482 14596
tri 43368 14541 43400 14573 ne
rect 43400 14550 43482 14573
rect 43528 14573 43610 14596
tri 43610 14573 43642 14605 sw
rect 70802 14580 71000 14638
rect 43528 14550 43642 14573
rect 43400 14541 43642 14550
tri 43400 14528 43413 14541 ne
rect 43413 14528 43642 14541
tri 43642 14528 43687 14573 sw
rect 70802 14534 70824 14580
rect 70870 14534 70928 14580
rect 70974 14534 71000 14580
tri 43413 14496 43445 14528 ne
rect 43445 14518 43687 14528
tri 43687 14518 43697 14528 sw
rect 43445 14496 43697 14518
tri 43445 14463 43478 14496 ne
rect 43478 14486 43697 14496
tri 43697 14486 43729 14518 sw
rect 43478 14473 43729 14486
tri 43729 14473 43742 14486 sw
rect 70802 14476 71000 14534
rect 43478 14464 43742 14473
rect 43478 14463 43614 14464
tri 43478 14417 43523 14463 ne
rect 43523 14418 43614 14463
rect 43660 14463 43742 14464
tri 43742 14463 43753 14473 sw
rect 43660 14418 43753 14463
rect 43523 14417 43753 14418
tri 43753 14417 43798 14463 sw
rect 70802 14430 70824 14476
rect 70870 14430 70928 14476
rect 70974 14430 71000 14476
tri 43523 14409 43532 14417 ne
rect 43532 14409 43798 14417
tri 43532 14389 43552 14409 ne
rect 43552 14396 43798 14409
tri 43798 14396 43819 14417 sw
rect 43552 14389 43819 14396
tri 43819 14389 43827 14396 sw
tri 43552 14364 43577 14389 ne
rect 43577 14386 43827 14389
tri 43827 14386 43829 14389 sw
rect 43577 14364 43829 14386
tri 43577 14354 43587 14364 ne
rect 43587 14354 43829 14364
tri 43829 14354 43861 14386 sw
rect 70802 14372 71000 14430
tri 43587 14309 43632 14354 ne
rect 43632 14341 43861 14354
tri 43861 14341 43874 14354 sw
rect 43632 14332 43874 14341
rect 43632 14309 43746 14332
tri 43632 14277 43664 14309 ne
rect 43664 14286 43746 14309
rect 43792 14309 43874 14332
tri 43874 14309 43906 14341 sw
rect 70802 14326 70824 14372
rect 70870 14326 70928 14372
rect 70974 14326 71000 14372
rect 43792 14286 43906 14309
rect 43664 14277 43906 14286
tri 43664 14264 43677 14277 ne
rect 43677 14264 43906 14277
tri 43906 14264 43951 14309 sw
rect 70802 14268 71000 14326
tri 43677 14232 43709 14264 ne
rect 43709 14254 43951 14264
tri 43951 14254 43961 14264 sw
rect 43709 14232 43961 14254
tri 43709 14187 43754 14232 ne
rect 43754 14222 43961 14232
tri 43961 14222 43993 14254 sw
rect 70802 14222 70824 14268
rect 70870 14222 70928 14268
rect 70974 14222 71000 14268
rect 43754 14209 43993 14222
tri 43993 14209 44006 14222 sw
rect 43754 14200 44006 14209
rect 43754 14187 43878 14200
tri 43754 14145 43796 14187 ne
rect 43796 14154 43878 14187
rect 43924 14177 44006 14200
tri 44006 14177 44038 14209 sw
rect 43924 14154 44038 14177
rect 43796 14145 44038 14154
tri 43796 14114 43827 14145 ne
rect 43827 14132 44038 14145
tri 44038 14132 44083 14177 sw
rect 70802 14164 71000 14222
rect 43827 14122 44083 14132
tri 44083 14122 44093 14132 sw
rect 43827 14114 44093 14122
tri 44093 14114 44101 14122 sw
rect 70802 14118 70824 14164
rect 70870 14118 70928 14164
rect 70974 14118 71000 14164
tri 43827 14100 43841 14114 ne
rect 43841 14100 44101 14114
tri 43841 14098 43843 14100 ne
rect 43843 14098 44101 14100
tri 43843 14090 43851 14098 ne
rect 43851 14090 44101 14098
tri 44101 14090 44125 14114 sw
tri 43851 14053 43888 14090 ne
rect 43888 14077 44125 14090
tri 44125 14077 44138 14090 sw
rect 43888 14068 44138 14077
rect 43888 14053 44010 14068
tri 43888 14013 43928 14053 ne
rect 43928 14022 44010 14053
rect 44056 14053 44138 14068
tri 44138 14053 44163 14077 sw
rect 70802 14060 71000 14118
rect 44056 14022 44163 14053
rect 43928 14013 44163 14022
tri 43928 14000 43941 14013 ne
rect 43941 14007 44163 14013
tri 44163 14007 44208 14053 sw
rect 70802 14014 70824 14060
rect 70870 14014 70928 14060
rect 70974 14014 71000 14060
rect 43941 14000 44208 14007
tri 44208 14000 44215 14007 sw
tri 43941 13968 43973 14000 ne
rect 43973 13990 44215 14000
tri 44215 13990 44225 14000 sw
rect 43973 13968 44225 13990
tri 43973 13923 44018 13968 ne
rect 44018 13958 44225 13968
tri 44225 13958 44257 13990 sw
rect 44018 13945 44257 13958
tri 44257 13945 44270 13958 sw
rect 70802 13956 71000 14014
rect 44018 13936 44270 13945
rect 44018 13923 44142 13936
tri 44018 13881 44060 13923 ne
rect 44060 13890 44142 13923
rect 44188 13913 44270 13936
tri 44270 13913 44302 13945 sw
rect 44188 13890 44302 13913
rect 44060 13881 44302 13890
tri 44060 13840 44101 13881 ne
rect 44101 13868 44302 13881
tri 44302 13868 44347 13913 sw
rect 70802 13910 70824 13956
rect 70870 13910 70928 13956
rect 70974 13910 71000 13956
rect 44101 13858 44347 13868
tri 44347 13858 44357 13868 sw
rect 44101 13840 44357 13858
tri 44357 13840 44375 13858 sw
rect 70802 13852 71000 13910
tri 44101 13836 44105 13840 ne
rect 44105 13836 44375 13840
tri 44105 13826 44115 13836 ne
rect 44115 13826 44375 13836
tri 44375 13826 44389 13840 sw
tri 44115 13781 44160 13826 ne
rect 44160 13813 44389 13826
tri 44389 13813 44402 13826 sw
rect 44160 13804 44402 13813
rect 44160 13781 44274 13804
tri 44160 13736 44205 13781 ne
rect 44205 13758 44274 13781
rect 44320 13781 44402 13804
tri 44402 13781 44434 13813 sw
rect 70802 13806 70824 13852
rect 70870 13806 70928 13852
rect 70974 13806 71000 13852
rect 44320 13758 44434 13781
rect 44205 13736 44434 13758
tri 44434 13736 44479 13781 sw
rect 70802 13748 71000 13806
tri 44205 13733 44208 13736 ne
rect 44208 13733 44479 13736
tri 44208 13688 44253 13733 ne
rect 44253 13726 44479 13733
tri 44479 13726 44489 13736 sw
rect 44253 13694 44489 13726
tri 44489 13694 44521 13726 sw
rect 70802 13702 70824 13748
rect 70870 13702 70928 13748
rect 70974 13702 71000 13748
rect 44253 13688 44521 13694
tri 44521 13688 44527 13694 sw
tri 44253 13643 44298 13688 ne
rect 44298 13672 44527 13688
rect 44298 13643 44406 13672
tri 44298 13617 44324 13643 ne
rect 44324 13626 44406 13643
rect 44452 13643 44527 13672
tri 44527 13643 44573 13688 sw
rect 70802 13644 71000 13702
rect 44452 13626 44573 13643
rect 44324 13617 44573 13626
tri 44324 13572 44369 13617 ne
rect 44369 13604 44573 13617
tri 44573 13604 44611 13643 sw
rect 44369 13594 44611 13604
tri 44611 13594 44621 13604 sw
rect 70802 13598 70824 13644
rect 70870 13598 70928 13644
rect 70974 13598 71000 13644
rect 44369 13572 44621 13594
tri 44369 13565 44375 13572 ne
rect 44375 13565 44621 13572
tri 44621 13565 44650 13594 sw
tri 44375 13562 44379 13565 ne
rect 44379 13562 44650 13565
tri 44650 13562 44653 13565 sw
tri 44379 13517 44424 13562 ne
rect 44424 13549 44653 13562
tri 44653 13549 44666 13562 sw
rect 44424 13540 44666 13549
rect 44424 13517 44538 13540
tri 44424 13485 44456 13517 ne
rect 44456 13494 44538 13517
rect 44584 13517 44666 13540
tri 44666 13517 44698 13549 sw
rect 70802 13540 71000 13598
rect 44584 13494 44698 13517
rect 44456 13485 44698 13494
tri 44456 13472 44469 13485 ne
rect 44469 13472 44698 13485
tri 44698 13472 44743 13517 sw
rect 70802 13494 70824 13540
rect 70870 13494 70928 13540
rect 70974 13494 71000 13540
tri 44469 13440 44501 13472 ne
rect 44501 13462 44743 13472
tri 44743 13462 44753 13472 sw
rect 44501 13440 44753 13462
tri 44501 13430 44511 13440 ne
rect 44511 13430 44753 13440
tri 44753 13430 44785 13462 sw
rect 70802 13436 71000 13494
tri 44511 13385 44556 13430 ne
rect 44556 13417 44785 13430
tri 44785 13417 44798 13430 sw
rect 44556 13413 44798 13417
tri 44798 13413 44802 13417 sw
rect 44556 13408 44802 13413
rect 44556 13385 44670 13408
tri 44556 13368 44573 13385 ne
rect 44573 13368 44670 13385
tri 44573 13340 44601 13368 ne
rect 44601 13362 44670 13368
rect 44716 13368 44802 13408
tri 44802 13368 44847 13413 sw
rect 70802 13390 70824 13436
rect 70870 13390 70928 13436
rect 70974 13390 71000 13436
rect 44716 13362 44847 13368
rect 44601 13340 44847 13362
tri 44847 13340 44875 13368 sw
tri 44601 13308 44633 13340 ne
rect 44633 13336 44875 13340
tri 44875 13336 44879 13340 sw
rect 44633 13308 44879 13336
tri 44633 13291 44650 13308 ne
rect 44650 13291 44879 13308
tri 44879 13291 44924 13336 sw
rect 70802 13291 71000 13390
tri 44650 13278 44663 13291 ne
rect 44663 13278 71000 13291
tri 44663 13233 44708 13278 ne
rect 44708 13269 71000 13278
rect 44708 13256 45088 13269
rect 44708 13233 44850 13256
tri 44708 13201 44740 13233 ne
rect 44740 13210 44850 13233
rect 44896 13223 45088 13256
rect 45134 13223 45192 13269
rect 45238 13223 45296 13269
rect 45342 13223 45400 13269
rect 45446 13223 45504 13269
rect 45550 13223 45608 13269
rect 45654 13223 45712 13269
rect 45758 13223 45816 13269
rect 45862 13223 45920 13269
rect 45966 13223 46024 13269
rect 46070 13223 46128 13269
rect 46174 13223 46232 13269
rect 46278 13223 46336 13269
rect 46382 13223 46440 13269
rect 46486 13223 46544 13269
rect 46590 13223 46648 13269
rect 46694 13223 46752 13269
rect 46798 13223 46856 13269
rect 46902 13223 46960 13269
rect 47006 13223 47064 13269
rect 47110 13223 47168 13269
rect 47214 13223 47272 13269
rect 47318 13223 47376 13269
rect 47422 13223 47480 13269
rect 47526 13223 47584 13269
rect 47630 13223 47688 13269
rect 47734 13223 47792 13269
rect 47838 13223 47896 13269
rect 47942 13223 48000 13269
rect 48046 13223 48104 13269
rect 48150 13223 48208 13269
rect 48254 13223 48312 13269
rect 48358 13223 48416 13269
rect 48462 13223 48520 13269
rect 48566 13223 48624 13269
rect 48670 13223 48728 13269
rect 48774 13223 48832 13269
rect 48878 13223 48936 13269
rect 48982 13223 49040 13269
rect 49086 13223 49144 13269
rect 49190 13223 49248 13269
rect 49294 13223 49352 13269
rect 49398 13223 49456 13269
rect 49502 13223 49560 13269
rect 49606 13223 49664 13269
rect 49710 13223 49768 13269
rect 49814 13223 49872 13269
rect 49918 13223 49976 13269
rect 50022 13223 50080 13269
rect 50126 13223 50184 13269
rect 50230 13223 50288 13269
rect 50334 13223 50392 13269
rect 50438 13223 50496 13269
rect 50542 13223 50600 13269
rect 50646 13223 50704 13269
rect 50750 13223 50808 13269
rect 50854 13223 50912 13269
rect 50958 13223 51016 13269
rect 51062 13223 51120 13269
rect 51166 13223 51224 13269
rect 51270 13223 51328 13269
rect 51374 13223 51432 13269
rect 51478 13223 51536 13269
rect 51582 13223 51640 13269
rect 51686 13223 51744 13269
rect 51790 13223 51848 13269
rect 51894 13223 51952 13269
rect 51998 13223 52056 13269
rect 52102 13223 52160 13269
rect 52206 13223 52264 13269
rect 52310 13223 52368 13269
rect 52414 13223 52472 13269
rect 52518 13223 52576 13269
rect 52622 13223 52680 13269
rect 52726 13223 52784 13269
rect 52830 13223 52888 13269
rect 52934 13223 52992 13269
rect 53038 13223 53096 13269
rect 53142 13223 53200 13269
rect 53246 13223 53304 13269
rect 53350 13223 53408 13269
rect 53454 13223 53512 13269
rect 53558 13223 53616 13269
rect 53662 13223 53720 13269
rect 53766 13223 53824 13269
rect 53870 13223 53928 13269
rect 53974 13223 54032 13269
rect 54078 13223 54136 13269
rect 54182 13223 54240 13269
rect 54286 13223 54344 13269
rect 54390 13223 54448 13269
rect 54494 13223 54552 13269
rect 54598 13223 54656 13269
rect 54702 13223 54760 13269
rect 54806 13223 54864 13269
rect 54910 13223 54968 13269
rect 55014 13223 55072 13269
rect 55118 13223 55176 13269
rect 55222 13223 55280 13269
rect 55326 13223 55384 13269
rect 55430 13223 55488 13269
rect 55534 13223 55592 13269
rect 55638 13223 55696 13269
rect 55742 13223 55800 13269
rect 55846 13223 55904 13269
rect 55950 13223 56008 13269
rect 56054 13223 56112 13269
rect 56158 13223 56216 13269
rect 56262 13223 56320 13269
rect 56366 13223 56424 13269
rect 56470 13223 56528 13269
rect 56574 13223 56632 13269
rect 56678 13223 56736 13269
rect 56782 13223 56840 13269
rect 56886 13223 56944 13269
rect 56990 13223 57048 13269
rect 57094 13223 57152 13269
rect 57198 13223 57256 13269
rect 57302 13223 57360 13269
rect 57406 13223 57464 13269
rect 57510 13223 57568 13269
rect 57614 13223 57672 13269
rect 57718 13223 57776 13269
rect 57822 13223 57880 13269
rect 57926 13223 57984 13269
rect 58030 13223 58088 13269
rect 58134 13223 58192 13269
rect 58238 13223 58296 13269
rect 58342 13223 58400 13269
rect 58446 13223 58504 13269
rect 58550 13223 58608 13269
rect 58654 13223 58712 13269
rect 58758 13223 58816 13269
rect 58862 13223 58920 13269
rect 58966 13223 59024 13269
rect 59070 13223 59128 13269
rect 59174 13223 59232 13269
rect 59278 13223 59336 13269
rect 59382 13223 59440 13269
rect 59486 13223 59544 13269
rect 59590 13223 59648 13269
rect 59694 13223 59752 13269
rect 59798 13223 59856 13269
rect 59902 13223 59960 13269
rect 60006 13223 60064 13269
rect 60110 13223 60168 13269
rect 60214 13223 60272 13269
rect 60318 13223 60376 13269
rect 60422 13223 60480 13269
rect 60526 13223 60584 13269
rect 60630 13223 60688 13269
rect 60734 13223 60792 13269
rect 60838 13223 60896 13269
rect 60942 13223 61000 13269
rect 61046 13223 61104 13269
rect 61150 13223 61208 13269
rect 61254 13223 61312 13269
rect 61358 13223 61416 13269
rect 61462 13223 61520 13269
rect 61566 13223 61624 13269
rect 61670 13223 61728 13269
rect 61774 13223 61832 13269
rect 61878 13223 61936 13269
rect 61982 13223 62040 13269
rect 62086 13223 62144 13269
rect 62190 13223 62248 13269
rect 62294 13223 62352 13269
rect 62398 13223 62456 13269
rect 62502 13223 62560 13269
rect 62606 13223 62664 13269
rect 62710 13223 62768 13269
rect 62814 13223 62872 13269
rect 62918 13223 62976 13269
rect 63022 13223 63080 13269
rect 63126 13223 63184 13269
rect 63230 13223 63288 13269
rect 63334 13223 63392 13269
rect 63438 13223 63496 13269
rect 63542 13223 63600 13269
rect 63646 13223 63704 13269
rect 63750 13223 63808 13269
rect 63854 13223 63912 13269
rect 63958 13223 64016 13269
rect 64062 13223 64120 13269
rect 64166 13223 64224 13269
rect 64270 13223 64328 13269
rect 64374 13223 64432 13269
rect 64478 13223 64536 13269
rect 64582 13223 64640 13269
rect 64686 13223 64744 13269
rect 64790 13223 64848 13269
rect 64894 13223 64952 13269
rect 64998 13223 65056 13269
rect 65102 13223 65160 13269
rect 65206 13223 65264 13269
rect 65310 13223 65368 13269
rect 65414 13223 65472 13269
rect 65518 13223 65576 13269
rect 65622 13223 65680 13269
rect 65726 13223 65784 13269
rect 65830 13223 65888 13269
rect 65934 13223 65992 13269
rect 66038 13223 66096 13269
rect 66142 13223 66200 13269
rect 66246 13223 66304 13269
rect 66350 13223 66408 13269
rect 66454 13223 66512 13269
rect 66558 13223 66616 13269
rect 66662 13223 66720 13269
rect 66766 13223 66824 13269
rect 66870 13223 66928 13269
rect 66974 13223 67032 13269
rect 67078 13223 67136 13269
rect 67182 13223 67240 13269
rect 67286 13223 67344 13269
rect 67390 13223 67448 13269
rect 67494 13223 67552 13269
rect 67598 13223 67656 13269
rect 67702 13223 67760 13269
rect 67806 13223 67864 13269
rect 67910 13223 67968 13269
rect 68014 13223 68072 13269
rect 68118 13223 68176 13269
rect 68222 13223 68280 13269
rect 68326 13223 68384 13269
rect 68430 13223 68488 13269
rect 68534 13223 68592 13269
rect 68638 13223 68696 13269
rect 68742 13223 68800 13269
rect 68846 13223 68904 13269
rect 68950 13223 69008 13269
rect 69054 13223 69112 13269
rect 69158 13223 69216 13269
rect 69262 13223 69320 13269
rect 69366 13223 69424 13269
rect 69470 13223 69528 13269
rect 69574 13223 69632 13269
rect 69678 13223 69736 13269
rect 69782 13223 69840 13269
rect 69886 13223 69944 13269
rect 69990 13223 70048 13269
rect 70094 13223 70152 13269
rect 70198 13223 70256 13269
rect 70302 13223 70360 13269
rect 70406 13223 70464 13269
rect 70510 13223 70568 13269
rect 70614 13223 70672 13269
rect 70718 13223 70776 13269
rect 70822 13223 70880 13269
rect 70926 13223 71000 13269
rect 44896 13210 71000 13223
rect 44740 13201 71000 13210
tri 44740 13188 44753 13201 ne
rect 44753 13188 71000 13201
tri 44753 13156 44785 13188 ne
rect 44785 13165 71000 13188
rect 44785 13156 45088 13165
tri 44785 13111 44830 13156 ne
rect 44830 13119 45088 13156
rect 45134 13119 45192 13165
rect 45238 13119 45296 13165
rect 45342 13119 45400 13165
rect 45446 13119 45504 13165
rect 45550 13119 45608 13165
rect 45654 13119 45712 13165
rect 45758 13119 45816 13165
rect 45862 13119 45920 13165
rect 45966 13119 46024 13165
rect 46070 13119 46128 13165
rect 46174 13119 46232 13165
rect 46278 13119 46336 13165
rect 46382 13119 46440 13165
rect 46486 13119 46544 13165
rect 46590 13119 46648 13165
rect 46694 13119 46752 13165
rect 46798 13119 46856 13165
rect 46902 13119 46960 13165
rect 47006 13119 47064 13165
rect 47110 13119 47168 13165
rect 47214 13119 47272 13165
rect 47318 13119 47376 13165
rect 47422 13119 47480 13165
rect 47526 13119 47584 13165
rect 47630 13119 47688 13165
rect 47734 13119 47792 13165
rect 47838 13119 47896 13165
rect 47942 13119 48000 13165
rect 48046 13119 48104 13165
rect 48150 13119 48208 13165
rect 48254 13119 48312 13165
rect 48358 13119 48416 13165
rect 48462 13119 48520 13165
rect 48566 13119 48624 13165
rect 48670 13119 48728 13165
rect 48774 13119 48832 13165
rect 48878 13119 48936 13165
rect 48982 13119 49040 13165
rect 49086 13119 49144 13165
rect 49190 13119 49248 13165
rect 49294 13119 49352 13165
rect 49398 13119 49456 13165
rect 49502 13119 49560 13165
rect 49606 13119 49664 13165
rect 49710 13119 49768 13165
rect 49814 13119 49872 13165
rect 49918 13119 49976 13165
rect 50022 13119 50080 13165
rect 50126 13119 50184 13165
rect 50230 13119 50288 13165
rect 50334 13119 50392 13165
rect 50438 13119 50496 13165
rect 50542 13119 50600 13165
rect 50646 13119 50704 13165
rect 50750 13119 50808 13165
rect 50854 13119 50912 13165
rect 50958 13119 51016 13165
rect 51062 13119 51120 13165
rect 51166 13119 51224 13165
rect 51270 13119 51328 13165
rect 51374 13119 51432 13165
rect 51478 13119 51536 13165
rect 51582 13119 51640 13165
rect 51686 13119 51744 13165
rect 51790 13119 51848 13165
rect 51894 13119 51952 13165
rect 51998 13119 52056 13165
rect 52102 13119 52160 13165
rect 52206 13119 52264 13165
rect 52310 13119 52368 13165
rect 52414 13119 52472 13165
rect 52518 13119 52576 13165
rect 52622 13119 52680 13165
rect 52726 13119 52784 13165
rect 52830 13119 52888 13165
rect 52934 13119 52992 13165
rect 53038 13119 53096 13165
rect 53142 13119 53200 13165
rect 53246 13119 53304 13165
rect 53350 13119 53408 13165
rect 53454 13119 53512 13165
rect 53558 13119 53616 13165
rect 53662 13119 53720 13165
rect 53766 13119 53824 13165
rect 53870 13119 53928 13165
rect 53974 13119 54032 13165
rect 54078 13119 54136 13165
rect 54182 13119 54240 13165
rect 54286 13119 54344 13165
rect 54390 13119 54448 13165
rect 54494 13119 54552 13165
rect 54598 13119 54656 13165
rect 54702 13119 54760 13165
rect 54806 13119 54864 13165
rect 54910 13119 54968 13165
rect 55014 13119 55072 13165
rect 55118 13119 55176 13165
rect 55222 13119 55280 13165
rect 55326 13119 55384 13165
rect 55430 13119 55488 13165
rect 55534 13119 55592 13165
rect 55638 13119 55696 13165
rect 55742 13119 55800 13165
rect 55846 13119 55904 13165
rect 55950 13119 56008 13165
rect 56054 13119 56112 13165
rect 56158 13119 56216 13165
rect 56262 13119 56320 13165
rect 56366 13119 56424 13165
rect 56470 13119 56528 13165
rect 56574 13119 56632 13165
rect 56678 13119 56736 13165
rect 56782 13119 56840 13165
rect 56886 13119 56944 13165
rect 56990 13119 57048 13165
rect 57094 13119 57152 13165
rect 57198 13119 57256 13165
rect 57302 13119 57360 13165
rect 57406 13119 57464 13165
rect 57510 13119 57568 13165
rect 57614 13119 57672 13165
rect 57718 13119 57776 13165
rect 57822 13119 57880 13165
rect 57926 13119 57984 13165
rect 58030 13119 58088 13165
rect 58134 13119 58192 13165
rect 58238 13119 58296 13165
rect 58342 13119 58400 13165
rect 58446 13119 58504 13165
rect 58550 13119 58608 13165
rect 58654 13119 58712 13165
rect 58758 13119 58816 13165
rect 58862 13119 58920 13165
rect 58966 13119 59024 13165
rect 59070 13119 59128 13165
rect 59174 13119 59232 13165
rect 59278 13119 59336 13165
rect 59382 13119 59440 13165
rect 59486 13119 59544 13165
rect 59590 13119 59648 13165
rect 59694 13119 59752 13165
rect 59798 13119 59856 13165
rect 59902 13119 59960 13165
rect 60006 13119 60064 13165
rect 60110 13119 60168 13165
rect 60214 13119 60272 13165
rect 60318 13119 60376 13165
rect 60422 13119 60480 13165
rect 60526 13119 60584 13165
rect 60630 13119 60688 13165
rect 60734 13119 60792 13165
rect 60838 13119 60896 13165
rect 60942 13119 61000 13165
rect 61046 13119 61104 13165
rect 61150 13119 61208 13165
rect 61254 13119 61312 13165
rect 61358 13119 61416 13165
rect 61462 13119 61520 13165
rect 61566 13119 61624 13165
rect 61670 13119 61728 13165
rect 61774 13119 61832 13165
rect 61878 13119 61936 13165
rect 61982 13119 62040 13165
rect 62086 13119 62144 13165
rect 62190 13119 62248 13165
rect 62294 13119 62352 13165
rect 62398 13119 62456 13165
rect 62502 13119 62560 13165
rect 62606 13119 62664 13165
rect 62710 13119 62768 13165
rect 62814 13119 62872 13165
rect 62918 13119 62976 13165
rect 63022 13119 63080 13165
rect 63126 13119 63184 13165
rect 63230 13119 63288 13165
rect 63334 13119 63392 13165
rect 63438 13119 63496 13165
rect 63542 13119 63600 13165
rect 63646 13119 63704 13165
rect 63750 13119 63808 13165
rect 63854 13119 63912 13165
rect 63958 13119 64016 13165
rect 64062 13119 64120 13165
rect 64166 13119 64224 13165
rect 64270 13119 64328 13165
rect 64374 13119 64432 13165
rect 64478 13119 64536 13165
rect 64582 13119 64640 13165
rect 64686 13119 64744 13165
rect 64790 13119 64848 13165
rect 64894 13119 64952 13165
rect 64998 13119 65056 13165
rect 65102 13119 65160 13165
rect 65206 13119 65264 13165
rect 65310 13119 65368 13165
rect 65414 13119 65472 13165
rect 65518 13119 65576 13165
rect 65622 13119 65680 13165
rect 65726 13119 65784 13165
rect 65830 13119 65888 13165
rect 65934 13119 65992 13165
rect 66038 13119 66096 13165
rect 66142 13119 66200 13165
rect 66246 13119 66304 13165
rect 66350 13119 66408 13165
rect 66454 13119 66512 13165
rect 66558 13119 66616 13165
rect 66662 13119 66720 13165
rect 66766 13119 66824 13165
rect 66870 13119 66928 13165
rect 66974 13119 67032 13165
rect 67078 13119 67136 13165
rect 67182 13119 67240 13165
rect 67286 13119 67344 13165
rect 67390 13119 67448 13165
rect 67494 13119 67552 13165
rect 67598 13119 67656 13165
rect 67702 13119 67760 13165
rect 67806 13119 67864 13165
rect 67910 13119 67968 13165
rect 68014 13119 68072 13165
rect 68118 13119 68176 13165
rect 68222 13119 68280 13165
rect 68326 13119 68384 13165
rect 68430 13119 68488 13165
rect 68534 13119 68592 13165
rect 68638 13119 68696 13165
rect 68742 13119 68800 13165
rect 68846 13119 68904 13165
rect 68950 13119 69008 13165
rect 69054 13119 69112 13165
rect 69158 13119 69216 13165
rect 69262 13119 69320 13165
rect 69366 13119 69424 13165
rect 69470 13119 69528 13165
rect 69574 13119 69632 13165
rect 69678 13119 69736 13165
rect 69782 13119 69840 13165
rect 69886 13119 69944 13165
rect 69990 13119 70048 13165
rect 70094 13119 70152 13165
rect 70198 13119 70256 13165
rect 70302 13119 70360 13165
rect 70406 13119 70464 13165
rect 70510 13119 70568 13165
rect 70614 13119 70672 13165
rect 70718 13119 70776 13165
rect 70822 13119 70880 13165
rect 70926 13119 71000 13165
rect 44830 13111 71000 13119
tri 44830 13110 44831 13111 ne
rect 44831 13110 71000 13111
tri 44831 13097 44844 13110 ne
rect 44844 13097 71000 13110
<< psubdiffcont >>
rect 13119 70929 13165 70975
rect 13223 70929 13269 70975
rect 13377 70929 13423 70975
rect 13481 70929 13527 70975
rect 13585 70929 13631 70975
rect 13689 70929 13735 70975
rect 13793 70929 13839 70975
rect 13897 70929 13943 70975
rect 14001 70929 14047 70975
rect 14105 70929 14151 70975
rect 14209 70929 14255 70975
rect 14313 70929 14359 70975
rect 14417 70929 14463 70975
rect 14521 70929 14567 70975
rect 14625 70929 14671 70975
rect 14729 70929 14775 70975
rect 14833 70929 14879 70975
rect 14937 70929 14983 70975
rect 15041 70929 15087 70975
rect 15145 70929 15191 70975
rect 15249 70929 15295 70975
rect 15353 70929 15399 70975
rect 15457 70929 15503 70975
rect 15561 70929 15607 70975
rect 15665 70929 15711 70975
rect 15769 70929 15815 70975
rect 15873 70929 15919 70975
rect 15977 70929 16023 70975
rect 16081 70929 16127 70975
rect 16185 70929 16231 70975
rect 16289 70929 16335 70975
rect 16393 70929 16439 70975
rect 16497 70929 16543 70975
rect 16601 70929 16647 70975
rect 16705 70929 16751 70975
rect 16809 70929 16855 70975
rect 16913 70929 16959 70975
rect 17017 70929 17063 70975
rect 17121 70929 17167 70975
rect 17225 70929 17271 70975
rect 17329 70929 17375 70975
rect 17433 70929 17479 70975
rect 17537 70929 17583 70975
rect 17641 70929 17687 70975
rect 17745 70929 17791 70975
rect 17849 70929 17895 70975
rect 17953 70929 17999 70975
rect 18057 70929 18103 70975
rect 18161 70929 18207 70975
rect 18265 70929 18311 70975
rect 18369 70929 18415 70975
rect 18473 70929 18519 70975
rect 18577 70929 18623 70975
rect 18681 70929 18727 70975
rect 18785 70929 18831 70975
rect 18889 70929 18935 70975
rect 18993 70929 19039 70975
rect 19097 70929 19143 70975
rect 19201 70929 19247 70975
rect 19305 70929 19351 70975
rect 19409 70929 19455 70975
rect 19513 70929 19559 70975
rect 19617 70929 19663 70975
rect 19721 70929 19767 70975
rect 19825 70929 19871 70975
rect 19929 70929 19975 70975
rect 20033 70929 20079 70975
rect 20137 70929 20183 70975
rect 20241 70929 20287 70975
rect 20345 70929 20391 70975
rect 20449 70929 20495 70975
rect 20553 70929 20599 70975
rect 20657 70929 20703 70975
rect 20761 70929 20807 70975
rect 20865 70929 20911 70975
rect 20969 70929 21015 70975
rect 21073 70929 21119 70975
rect 21177 70929 21223 70975
rect 21281 70929 21327 70975
rect 21385 70929 21431 70975
rect 21489 70929 21535 70975
rect 21593 70929 21639 70975
rect 21697 70929 21743 70975
rect 21801 70929 21847 70975
rect 21905 70929 21951 70975
rect 22009 70929 22055 70975
rect 22113 70929 22159 70975
rect 22217 70929 22263 70975
rect 22321 70929 22367 70975
rect 22425 70929 22471 70975
rect 22529 70929 22575 70975
rect 22633 70929 22679 70975
rect 22737 70929 22783 70975
rect 22841 70929 22887 70975
rect 22945 70929 22991 70975
rect 23049 70929 23095 70975
rect 23153 70929 23199 70975
rect 23257 70929 23303 70975
rect 23361 70929 23407 70975
rect 23465 70929 23511 70975
rect 23569 70929 23615 70975
rect 23673 70929 23719 70975
rect 23777 70929 23823 70975
rect 23881 70929 23927 70975
rect 23985 70929 24031 70975
rect 24089 70929 24135 70975
rect 24193 70929 24239 70975
rect 24297 70929 24343 70975
rect 24401 70929 24447 70975
rect 24505 70929 24551 70975
rect 24609 70929 24655 70975
rect 24713 70929 24759 70975
rect 24817 70929 24863 70975
rect 24921 70929 24967 70975
rect 25025 70929 25071 70975
rect 25129 70929 25175 70975
rect 25233 70929 25279 70975
rect 25337 70929 25383 70975
rect 25441 70929 25487 70975
rect 25545 70929 25591 70975
rect 25649 70929 25695 70975
rect 25753 70929 25799 70975
rect 25857 70929 25903 70975
rect 25961 70929 26007 70975
rect 26065 70929 26111 70975
rect 26169 70929 26215 70975
rect 26273 70929 26319 70975
rect 26377 70929 26423 70975
rect 26481 70929 26527 70975
rect 26585 70929 26631 70975
rect 26689 70929 26735 70975
rect 26793 70929 26839 70975
rect 26897 70929 26943 70975
rect 27001 70929 27047 70975
rect 27105 70929 27151 70975
rect 27209 70929 27255 70975
rect 27313 70929 27359 70975
rect 27417 70929 27463 70975
rect 27521 70929 27567 70975
rect 27625 70929 27671 70975
rect 27729 70929 27775 70975
rect 27833 70929 27879 70975
rect 27937 70929 27983 70975
rect 28041 70929 28087 70975
rect 28145 70929 28191 70975
rect 28249 70929 28295 70975
rect 28353 70929 28399 70975
rect 28457 70929 28503 70975
rect 28561 70929 28607 70975
rect 28665 70929 28711 70975
rect 28769 70929 28815 70975
rect 28873 70929 28919 70975
rect 28977 70929 29023 70975
rect 29081 70929 29127 70975
rect 29185 70929 29231 70975
rect 29289 70929 29335 70975
rect 29393 70929 29439 70975
rect 29497 70929 29543 70975
rect 29601 70929 29647 70975
rect 29705 70929 29751 70975
rect 29809 70929 29855 70975
rect 29913 70929 29959 70975
rect 30017 70929 30063 70975
rect 30121 70929 30167 70975
rect 30225 70929 30271 70975
rect 30329 70929 30375 70975
rect 30433 70929 30479 70975
rect 30537 70929 30583 70975
rect 30641 70929 30687 70975
rect 30745 70929 30791 70975
rect 30849 70929 30895 70975
rect 30953 70929 30999 70975
rect 31057 70929 31103 70975
rect 31161 70929 31207 70975
rect 31265 70929 31311 70975
rect 31369 70929 31415 70975
rect 31473 70929 31519 70975
rect 31577 70929 31623 70975
rect 31681 70929 31727 70975
rect 31785 70929 31831 70975
rect 31889 70929 31935 70975
rect 31993 70929 32039 70975
rect 32097 70929 32143 70975
rect 32201 70929 32247 70975
rect 32305 70929 32351 70975
rect 32409 70929 32455 70975
rect 32513 70929 32559 70975
rect 32617 70929 32663 70975
rect 32721 70929 32767 70975
rect 32825 70929 32871 70975
rect 32929 70929 32975 70975
rect 33033 70929 33079 70975
rect 33137 70929 33183 70975
rect 33241 70929 33287 70975
rect 33345 70929 33391 70975
rect 33449 70929 33495 70975
rect 33553 70929 33599 70975
rect 33657 70929 33703 70975
rect 33761 70929 33807 70975
rect 33865 70929 33911 70975
rect 33969 70929 34015 70975
rect 34073 70929 34119 70975
rect 34177 70929 34223 70975
rect 34281 70929 34327 70975
rect 34385 70929 34431 70975
rect 34489 70929 34535 70975
rect 34593 70929 34639 70975
rect 34697 70929 34743 70975
rect 34801 70929 34847 70975
rect 34905 70929 34951 70975
rect 35009 70929 35055 70975
rect 35113 70929 35159 70975
rect 35217 70929 35263 70975
rect 35321 70929 35367 70975
rect 35425 70929 35471 70975
rect 35529 70929 35575 70975
rect 35633 70929 35679 70975
rect 35737 70929 35783 70975
rect 35841 70929 35887 70975
rect 35945 70929 35991 70975
rect 36049 70929 36095 70975
rect 36153 70929 36199 70975
rect 36257 70929 36303 70975
rect 36361 70929 36407 70975
rect 36465 70929 36511 70975
rect 36569 70929 36615 70975
rect 36673 70929 36719 70975
rect 36777 70929 36823 70975
rect 36881 70929 36927 70975
rect 36985 70929 37031 70975
rect 37089 70929 37135 70975
rect 37193 70929 37239 70975
rect 37297 70929 37343 70975
rect 37401 70929 37447 70975
rect 37505 70929 37551 70975
rect 37609 70929 37655 70975
rect 37713 70929 37759 70975
rect 37817 70929 37863 70975
rect 37921 70929 37967 70975
rect 38025 70929 38071 70975
rect 38129 70929 38175 70975
rect 38233 70929 38279 70975
rect 38337 70929 38383 70975
rect 38441 70929 38487 70975
rect 38545 70929 38591 70975
rect 38649 70929 38695 70975
rect 38753 70929 38799 70975
rect 38857 70929 38903 70975
rect 38961 70929 39007 70975
rect 39065 70929 39111 70975
rect 39169 70929 39215 70975
rect 39273 70929 39319 70975
rect 39377 70929 39423 70975
rect 39481 70929 39527 70975
rect 39585 70929 39631 70975
rect 39689 70929 39735 70975
rect 39793 70929 39839 70975
rect 39897 70929 39943 70975
rect 40001 70929 40047 70975
rect 40105 70929 40151 70975
rect 40209 70929 40255 70975
rect 40313 70929 40359 70975
rect 40417 70929 40463 70975
rect 40521 70929 40567 70975
rect 40625 70929 40671 70975
rect 40729 70929 40775 70975
rect 40833 70929 40879 70975
rect 40937 70929 40983 70975
rect 41041 70929 41087 70975
rect 41145 70929 41191 70975
rect 41249 70929 41295 70975
rect 41353 70929 41399 70975
rect 41457 70929 41503 70975
rect 41561 70929 41607 70975
rect 41665 70929 41711 70975
rect 41769 70929 41815 70975
rect 41873 70929 41919 70975
rect 41977 70929 42023 70975
rect 42081 70929 42127 70975
rect 42185 70929 42231 70975
rect 42289 70929 42335 70975
rect 42393 70929 42439 70975
rect 42497 70929 42543 70975
rect 42601 70929 42647 70975
rect 42705 70929 42751 70975
rect 42809 70929 42855 70975
rect 42913 70929 42959 70975
rect 43017 70929 43063 70975
rect 43121 70929 43167 70975
rect 43225 70929 43271 70975
rect 43329 70929 43375 70975
rect 43433 70929 43479 70975
rect 43537 70929 43583 70975
rect 43641 70929 43687 70975
rect 43745 70929 43791 70975
rect 43849 70929 43895 70975
rect 43953 70929 43999 70975
rect 44057 70929 44103 70975
rect 44161 70929 44207 70975
rect 44265 70929 44311 70975
rect 44369 70929 44415 70975
rect 44473 70929 44519 70975
rect 44577 70929 44623 70975
rect 44681 70929 44727 70975
rect 44785 70929 44831 70975
rect 44889 70929 44935 70975
rect 44993 70929 45039 70975
rect 45097 70929 45143 70975
rect 45201 70929 45247 70975
rect 45305 70929 45351 70975
rect 45409 70929 45455 70975
rect 45513 70929 45559 70975
rect 45617 70929 45663 70975
rect 45721 70929 45767 70975
rect 45825 70929 45871 70975
rect 45929 70929 45975 70975
rect 46033 70929 46079 70975
rect 46137 70929 46183 70975
rect 46241 70929 46287 70975
rect 46345 70929 46391 70975
rect 46449 70929 46495 70975
rect 46553 70929 46599 70975
rect 46657 70929 46703 70975
rect 46761 70929 46807 70975
rect 46865 70929 46911 70975
rect 46969 70929 47015 70975
rect 47073 70929 47119 70975
rect 47177 70929 47223 70975
rect 47281 70929 47327 70975
rect 47385 70929 47431 70975
rect 47489 70929 47535 70975
rect 47593 70929 47639 70975
rect 47697 70929 47743 70975
rect 47801 70929 47847 70975
rect 47905 70929 47951 70975
rect 48009 70929 48055 70975
rect 48113 70929 48159 70975
rect 48217 70929 48263 70975
rect 48321 70929 48367 70975
rect 48425 70929 48471 70975
rect 48529 70929 48575 70975
rect 48633 70929 48679 70975
rect 48737 70929 48783 70975
rect 48841 70929 48887 70975
rect 48945 70929 48991 70975
rect 49049 70929 49095 70975
rect 49153 70929 49199 70975
rect 49257 70929 49303 70975
rect 49361 70929 49407 70975
rect 49465 70929 49511 70975
rect 49569 70929 49615 70975
rect 49673 70929 49719 70975
rect 49777 70929 49823 70975
rect 49881 70929 49927 70975
rect 49985 70929 50031 70975
rect 50089 70929 50135 70975
rect 50193 70929 50239 70975
rect 50297 70929 50343 70975
rect 50401 70929 50447 70975
rect 50505 70929 50551 70975
rect 50609 70929 50655 70975
rect 50713 70929 50759 70975
rect 50817 70929 50863 70975
rect 50921 70929 50967 70975
rect 51025 70929 51071 70975
rect 51129 70929 51175 70975
rect 51233 70929 51279 70975
rect 51337 70929 51383 70975
rect 51441 70929 51487 70975
rect 51545 70929 51591 70975
rect 51649 70929 51695 70975
rect 51753 70929 51799 70975
rect 51857 70929 51903 70975
rect 51961 70929 52007 70975
rect 52065 70929 52111 70975
rect 52169 70929 52215 70975
rect 52273 70929 52319 70975
rect 52377 70929 52423 70975
rect 52481 70929 52527 70975
rect 52585 70929 52631 70975
rect 52689 70929 52735 70975
rect 52793 70929 52839 70975
rect 52897 70929 52943 70975
rect 53001 70929 53047 70975
rect 53105 70929 53151 70975
rect 53209 70929 53255 70975
rect 53313 70929 53359 70975
rect 53417 70929 53463 70975
rect 53521 70929 53567 70975
rect 53625 70929 53671 70975
rect 53729 70929 53775 70975
rect 53833 70929 53879 70975
rect 53937 70929 53983 70975
rect 54041 70929 54087 70975
rect 54145 70929 54191 70975
rect 54249 70929 54295 70975
rect 54353 70929 54399 70975
rect 54457 70929 54503 70975
rect 54561 70929 54607 70975
rect 54665 70929 54711 70975
rect 54769 70929 54815 70975
rect 54873 70929 54919 70975
rect 54977 70929 55023 70975
rect 55081 70929 55127 70975
rect 55185 70929 55231 70975
rect 55289 70929 55335 70975
rect 55393 70929 55439 70975
rect 55497 70929 55543 70975
rect 55601 70929 55647 70975
rect 55705 70929 55751 70975
rect 55809 70929 55855 70975
rect 55913 70929 55959 70975
rect 56017 70929 56063 70975
rect 56121 70929 56167 70975
rect 56225 70929 56271 70975
rect 56329 70929 56375 70975
rect 56433 70929 56479 70975
rect 56537 70929 56583 70975
rect 56641 70929 56687 70975
rect 56745 70929 56791 70975
rect 56849 70929 56895 70975
rect 56953 70929 56999 70975
rect 57057 70929 57103 70975
rect 57161 70929 57207 70975
rect 57265 70929 57311 70975
rect 57369 70929 57415 70975
rect 57473 70929 57519 70975
rect 57577 70929 57623 70975
rect 57681 70929 57727 70975
rect 57785 70929 57831 70975
rect 57889 70929 57935 70975
rect 57993 70929 58039 70975
rect 58097 70929 58143 70975
rect 58201 70929 58247 70975
rect 58305 70929 58351 70975
rect 58409 70929 58455 70975
rect 58513 70929 58559 70975
rect 58617 70929 58663 70975
rect 58721 70929 58767 70975
rect 58825 70929 58871 70975
rect 58929 70929 58975 70975
rect 59033 70929 59079 70975
rect 59137 70929 59183 70975
rect 59241 70929 59287 70975
rect 59345 70929 59391 70975
rect 59449 70929 59495 70975
rect 59553 70929 59599 70975
rect 59657 70929 59703 70975
rect 59761 70929 59807 70975
rect 59865 70929 59911 70975
rect 59969 70929 60015 70975
rect 60073 70929 60119 70975
rect 60177 70929 60223 70975
rect 60281 70929 60327 70975
rect 60385 70929 60431 70975
rect 60489 70929 60535 70975
rect 60593 70929 60639 70975
rect 60697 70929 60743 70975
rect 60801 70929 60847 70975
rect 60905 70929 60951 70975
rect 61009 70929 61055 70975
rect 61113 70929 61159 70975
rect 61217 70929 61263 70975
rect 61321 70929 61367 70975
rect 61425 70929 61471 70975
rect 61529 70929 61575 70975
rect 61633 70929 61679 70975
rect 61737 70929 61783 70975
rect 61841 70929 61887 70975
rect 61945 70929 61991 70975
rect 62049 70929 62095 70975
rect 62153 70929 62199 70975
rect 62257 70929 62303 70975
rect 62361 70929 62407 70975
rect 62465 70929 62511 70975
rect 62569 70929 62615 70975
rect 62673 70929 62719 70975
rect 62777 70929 62823 70975
rect 62881 70929 62927 70975
rect 62985 70929 63031 70975
rect 63089 70929 63135 70975
rect 63193 70929 63239 70975
rect 63297 70929 63343 70975
rect 63401 70929 63447 70975
rect 63505 70929 63551 70975
rect 63609 70929 63655 70975
rect 63713 70929 63759 70975
rect 63817 70929 63863 70975
rect 63921 70929 63967 70975
rect 64025 70929 64071 70975
rect 64129 70929 64175 70975
rect 64233 70929 64279 70975
rect 64337 70929 64383 70975
rect 64441 70929 64487 70975
rect 64545 70929 64591 70975
rect 64649 70929 64695 70975
rect 64753 70929 64799 70975
rect 64857 70929 64903 70975
rect 64961 70929 65007 70975
rect 65065 70929 65111 70975
rect 65169 70929 65215 70975
rect 65273 70929 65319 70975
rect 65377 70929 65423 70975
rect 65481 70929 65527 70975
rect 65585 70929 65631 70975
rect 65689 70929 65735 70975
rect 65793 70929 65839 70975
rect 65897 70929 65943 70975
rect 66001 70929 66047 70975
rect 66105 70929 66151 70975
rect 66209 70929 66255 70975
rect 66313 70929 66359 70975
rect 66417 70929 66463 70975
rect 66521 70929 66567 70975
rect 66625 70929 66671 70975
rect 66729 70929 66775 70975
rect 66833 70929 66879 70975
rect 66937 70929 66983 70975
rect 67041 70929 67087 70975
rect 67145 70929 67191 70975
rect 67249 70929 67295 70975
rect 67353 70929 67399 70975
rect 67457 70929 67503 70975
rect 67561 70929 67607 70975
rect 67665 70929 67711 70975
rect 67769 70929 67815 70975
rect 67873 70929 67919 70975
rect 67977 70929 68023 70975
rect 68081 70929 68127 70975
rect 68185 70929 68231 70975
rect 68289 70929 68335 70975
rect 68393 70929 68439 70975
rect 68497 70929 68543 70975
rect 68601 70929 68647 70975
rect 68705 70929 68751 70975
rect 68809 70929 68855 70975
rect 68913 70929 68959 70975
rect 69017 70929 69063 70975
rect 69121 70929 69167 70975
rect 69225 70929 69271 70975
rect 69329 70929 69375 70975
rect 69433 70929 69479 70975
rect 69537 70929 69583 70975
rect 69641 70929 69687 70975
rect 69745 70929 69791 70975
rect 69849 70929 69895 70975
rect 13119 70825 13165 70871
rect 13223 70825 13269 70871
rect 13377 70825 13423 70871
rect 13481 70825 13527 70871
rect 13585 70825 13631 70871
rect 13689 70825 13735 70871
rect 13793 70825 13839 70871
rect 13897 70825 13943 70871
rect 14001 70825 14047 70871
rect 14105 70825 14151 70871
rect 14209 70825 14255 70871
rect 14313 70825 14359 70871
rect 14417 70825 14463 70871
rect 14521 70825 14567 70871
rect 14625 70825 14671 70871
rect 14729 70825 14775 70871
rect 14833 70825 14879 70871
rect 14937 70825 14983 70871
rect 15041 70825 15087 70871
rect 15145 70825 15191 70871
rect 15249 70825 15295 70871
rect 15353 70825 15399 70871
rect 15457 70825 15503 70871
rect 15561 70825 15607 70871
rect 15665 70825 15711 70871
rect 15769 70825 15815 70871
rect 15873 70825 15919 70871
rect 15977 70825 16023 70871
rect 16081 70825 16127 70871
rect 16185 70825 16231 70871
rect 16289 70825 16335 70871
rect 16393 70825 16439 70871
rect 16497 70825 16543 70871
rect 16601 70825 16647 70871
rect 16705 70825 16751 70871
rect 16809 70825 16855 70871
rect 16913 70825 16959 70871
rect 17017 70825 17063 70871
rect 17121 70825 17167 70871
rect 17225 70825 17271 70871
rect 17329 70825 17375 70871
rect 17433 70825 17479 70871
rect 17537 70825 17583 70871
rect 17641 70825 17687 70871
rect 17745 70825 17791 70871
rect 17849 70825 17895 70871
rect 17953 70825 17999 70871
rect 18057 70825 18103 70871
rect 18161 70825 18207 70871
rect 18265 70825 18311 70871
rect 18369 70825 18415 70871
rect 18473 70825 18519 70871
rect 18577 70825 18623 70871
rect 18681 70825 18727 70871
rect 18785 70825 18831 70871
rect 18889 70825 18935 70871
rect 18993 70825 19039 70871
rect 19097 70825 19143 70871
rect 19201 70825 19247 70871
rect 19305 70825 19351 70871
rect 19409 70825 19455 70871
rect 19513 70825 19559 70871
rect 19617 70825 19663 70871
rect 19721 70825 19767 70871
rect 19825 70825 19871 70871
rect 19929 70825 19975 70871
rect 20033 70825 20079 70871
rect 20137 70825 20183 70871
rect 20241 70825 20287 70871
rect 20345 70825 20391 70871
rect 20449 70825 20495 70871
rect 20553 70825 20599 70871
rect 20657 70825 20703 70871
rect 20761 70825 20807 70871
rect 20865 70825 20911 70871
rect 20969 70825 21015 70871
rect 21073 70825 21119 70871
rect 21177 70825 21223 70871
rect 21281 70825 21327 70871
rect 21385 70825 21431 70871
rect 21489 70825 21535 70871
rect 21593 70825 21639 70871
rect 21697 70825 21743 70871
rect 21801 70825 21847 70871
rect 21905 70825 21951 70871
rect 22009 70825 22055 70871
rect 22113 70825 22159 70871
rect 22217 70825 22263 70871
rect 22321 70825 22367 70871
rect 22425 70825 22471 70871
rect 22529 70825 22575 70871
rect 22633 70825 22679 70871
rect 22737 70825 22783 70871
rect 22841 70825 22887 70871
rect 22945 70825 22991 70871
rect 23049 70825 23095 70871
rect 23153 70825 23199 70871
rect 23257 70825 23303 70871
rect 23361 70825 23407 70871
rect 23465 70825 23511 70871
rect 23569 70825 23615 70871
rect 23673 70825 23719 70871
rect 23777 70825 23823 70871
rect 23881 70825 23927 70871
rect 23985 70825 24031 70871
rect 24089 70825 24135 70871
rect 24193 70825 24239 70871
rect 24297 70825 24343 70871
rect 24401 70825 24447 70871
rect 24505 70825 24551 70871
rect 24609 70825 24655 70871
rect 24713 70825 24759 70871
rect 24817 70825 24863 70871
rect 24921 70825 24967 70871
rect 25025 70825 25071 70871
rect 25129 70825 25175 70871
rect 25233 70825 25279 70871
rect 25337 70825 25383 70871
rect 25441 70825 25487 70871
rect 25545 70825 25591 70871
rect 25649 70825 25695 70871
rect 25753 70825 25799 70871
rect 25857 70825 25903 70871
rect 25961 70825 26007 70871
rect 26065 70825 26111 70871
rect 26169 70825 26215 70871
rect 26273 70825 26319 70871
rect 26377 70825 26423 70871
rect 26481 70825 26527 70871
rect 26585 70825 26631 70871
rect 26689 70825 26735 70871
rect 26793 70825 26839 70871
rect 26897 70825 26943 70871
rect 27001 70825 27047 70871
rect 27105 70825 27151 70871
rect 27209 70825 27255 70871
rect 27313 70825 27359 70871
rect 27417 70825 27463 70871
rect 27521 70825 27567 70871
rect 27625 70825 27671 70871
rect 27729 70825 27775 70871
rect 27833 70825 27879 70871
rect 27937 70825 27983 70871
rect 28041 70825 28087 70871
rect 28145 70825 28191 70871
rect 28249 70825 28295 70871
rect 28353 70825 28399 70871
rect 28457 70825 28503 70871
rect 28561 70825 28607 70871
rect 28665 70825 28711 70871
rect 28769 70825 28815 70871
rect 28873 70825 28919 70871
rect 28977 70825 29023 70871
rect 29081 70825 29127 70871
rect 29185 70825 29231 70871
rect 29289 70825 29335 70871
rect 29393 70825 29439 70871
rect 29497 70825 29543 70871
rect 29601 70825 29647 70871
rect 29705 70825 29751 70871
rect 29809 70825 29855 70871
rect 29913 70825 29959 70871
rect 30017 70825 30063 70871
rect 30121 70825 30167 70871
rect 30225 70825 30271 70871
rect 30329 70825 30375 70871
rect 30433 70825 30479 70871
rect 30537 70825 30583 70871
rect 30641 70825 30687 70871
rect 30745 70825 30791 70871
rect 30849 70825 30895 70871
rect 30953 70825 30999 70871
rect 31057 70825 31103 70871
rect 31161 70825 31207 70871
rect 31265 70825 31311 70871
rect 31369 70825 31415 70871
rect 31473 70825 31519 70871
rect 31577 70825 31623 70871
rect 31681 70825 31727 70871
rect 31785 70825 31831 70871
rect 31889 70825 31935 70871
rect 31993 70825 32039 70871
rect 32097 70825 32143 70871
rect 32201 70825 32247 70871
rect 32305 70825 32351 70871
rect 32409 70825 32455 70871
rect 32513 70825 32559 70871
rect 32617 70825 32663 70871
rect 32721 70825 32767 70871
rect 32825 70825 32871 70871
rect 32929 70825 32975 70871
rect 33033 70825 33079 70871
rect 33137 70825 33183 70871
rect 33241 70825 33287 70871
rect 33345 70825 33391 70871
rect 33449 70825 33495 70871
rect 33553 70825 33599 70871
rect 33657 70825 33703 70871
rect 33761 70825 33807 70871
rect 33865 70825 33911 70871
rect 33969 70825 34015 70871
rect 34073 70825 34119 70871
rect 34177 70825 34223 70871
rect 34281 70825 34327 70871
rect 34385 70825 34431 70871
rect 34489 70825 34535 70871
rect 34593 70825 34639 70871
rect 34697 70825 34743 70871
rect 34801 70825 34847 70871
rect 34905 70825 34951 70871
rect 35009 70825 35055 70871
rect 35113 70825 35159 70871
rect 35217 70825 35263 70871
rect 35321 70825 35367 70871
rect 35425 70825 35471 70871
rect 35529 70825 35575 70871
rect 35633 70825 35679 70871
rect 35737 70825 35783 70871
rect 35841 70825 35887 70871
rect 35945 70825 35991 70871
rect 36049 70825 36095 70871
rect 36153 70825 36199 70871
rect 36257 70825 36303 70871
rect 36361 70825 36407 70871
rect 36465 70825 36511 70871
rect 36569 70825 36615 70871
rect 36673 70825 36719 70871
rect 36777 70825 36823 70871
rect 36881 70825 36927 70871
rect 36985 70825 37031 70871
rect 37089 70825 37135 70871
rect 37193 70825 37239 70871
rect 37297 70825 37343 70871
rect 37401 70825 37447 70871
rect 37505 70825 37551 70871
rect 37609 70825 37655 70871
rect 37713 70825 37759 70871
rect 37817 70825 37863 70871
rect 37921 70825 37967 70871
rect 38025 70825 38071 70871
rect 38129 70825 38175 70871
rect 38233 70825 38279 70871
rect 38337 70825 38383 70871
rect 38441 70825 38487 70871
rect 38545 70825 38591 70871
rect 38649 70825 38695 70871
rect 38753 70825 38799 70871
rect 38857 70825 38903 70871
rect 38961 70825 39007 70871
rect 39065 70825 39111 70871
rect 39169 70825 39215 70871
rect 39273 70825 39319 70871
rect 39377 70825 39423 70871
rect 39481 70825 39527 70871
rect 39585 70825 39631 70871
rect 39689 70825 39735 70871
rect 39793 70825 39839 70871
rect 39897 70825 39943 70871
rect 40001 70825 40047 70871
rect 40105 70825 40151 70871
rect 40209 70825 40255 70871
rect 40313 70825 40359 70871
rect 40417 70825 40463 70871
rect 40521 70825 40567 70871
rect 40625 70825 40671 70871
rect 40729 70825 40775 70871
rect 40833 70825 40879 70871
rect 40937 70825 40983 70871
rect 41041 70825 41087 70871
rect 41145 70825 41191 70871
rect 41249 70825 41295 70871
rect 41353 70825 41399 70871
rect 41457 70825 41503 70871
rect 41561 70825 41607 70871
rect 41665 70825 41711 70871
rect 41769 70825 41815 70871
rect 41873 70825 41919 70871
rect 41977 70825 42023 70871
rect 42081 70825 42127 70871
rect 42185 70825 42231 70871
rect 42289 70825 42335 70871
rect 42393 70825 42439 70871
rect 42497 70825 42543 70871
rect 42601 70825 42647 70871
rect 42705 70825 42751 70871
rect 42809 70825 42855 70871
rect 42913 70825 42959 70871
rect 43017 70825 43063 70871
rect 43121 70825 43167 70871
rect 43225 70825 43271 70871
rect 43329 70825 43375 70871
rect 43433 70825 43479 70871
rect 43537 70825 43583 70871
rect 43641 70825 43687 70871
rect 43745 70825 43791 70871
rect 43849 70825 43895 70871
rect 43953 70825 43999 70871
rect 44057 70825 44103 70871
rect 44161 70825 44207 70871
rect 44265 70825 44311 70871
rect 44369 70825 44415 70871
rect 44473 70825 44519 70871
rect 44577 70825 44623 70871
rect 44681 70825 44727 70871
rect 44785 70825 44831 70871
rect 44889 70825 44935 70871
rect 44993 70825 45039 70871
rect 45097 70825 45143 70871
rect 45201 70825 45247 70871
rect 45305 70825 45351 70871
rect 45409 70825 45455 70871
rect 45513 70825 45559 70871
rect 45617 70825 45663 70871
rect 45721 70825 45767 70871
rect 45825 70825 45871 70871
rect 45929 70825 45975 70871
rect 46033 70825 46079 70871
rect 46137 70825 46183 70871
rect 46241 70825 46287 70871
rect 46345 70825 46391 70871
rect 46449 70825 46495 70871
rect 46553 70825 46599 70871
rect 46657 70825 46703 70871
rect 46761 70825 46807 70871
rect 46865 70825 46911 70871
rect 46969 70825 47015 70871
rect 47073 70825 47119 70871
rect 47177 70825 47223 70871
rect 47281 70825 47327 70871
rect 47385 70825 47431 70871
rect 47489 70825 47535 70871
rect 47593 70825 47639 70871
rect 47697 70825 47743 70871
rect 47801 70825 47847 70871
rect 47905 70825 47951 70871
rect 48009 70825 48055 70871
rect 48113 70825 48159 70871
rect 48217 70825 48263 70871
rect 48321 70825 48367 70871
rect 48425 70825 48471 70871
rect 48529 70825 48575 70871
rect 48633 70825 48679 70871
rect 48737 70825 48783 70871
rect 48841 70825 48887 70871
rect 48945 70825 48991 70871
rect 49049 70825 49095 70871
rect 49153 70825 49199 70871
rect 49257 70825 49303 70871
rect 49361 70825 49407 70871
rect 49465 70825 49511 70871
rect 49569 70825 49615 70871
rect 49673 70825 49719 70871
rect 49777 70825 49823 70871
rect 49881 70825 49927 70871
rect 49985 70825 50031 70871
rect 50089 70825 50135 70871
rect 50193 70825 50239 70871
rect 50297 70825 50343 70871
rect 50401 70825 50447 70871
rect 50505 70825 50551 70871
rect 50609 70825 50655 70871
rect 50713 70825 50759 70871
rect 50817 70825 50863 70871
rect 50921 70825 50967 70871
rect 51025 70825 51071 70871
rect 51129 70825 51175 70871
rect 51233 70825 51279 70871
rect 51337 70825 51383 70871
rect 51441 70825 51487 70871
rect 51545 70825 51591 70871
rect 51649 70825 51695 70871
rect 51753 70825 51799 70871
rect 51857 70825 51903 70871
rect 51961 70825 52007 70871
rect 52065 70825 52111 70871
rect 52169 70825 52215 70871
rect 52273 70825 52319 70871
rect 52377 70825 52423 70871
rect 52481 70825 52527 70871
rect 52585 70825 52631 70871
rect 52689 70825 52735 70871
rect 52793 70825 52839 70871
rect 52897 70825 52943 70871
rect 53001 70825 53047 70871
rect 53105 70825 53151 70871
rect 53209 70825 53255 70871
rect 53313 70825 53359 70871
rect 53417 70825 53463 70871
rect 53521 70825 53567 70871
rect 53625 70825 53671 70871
rect 53729 70825 53775 70871
rect 53833 70825 53879 70871
rect 53937 70825 53983 70871
rect 54041 70825 54087 70871
rect 54145 70825 54191 70871
rect 54249 70825 54295 70871
rect 54353 70825 54399 70871
rect 54457 70825 54503 70871
rect 54561 70825 54607 70871
rect 54665 70825 54711 70871
rect 54769 70825 54815 70871
rect 54873 70825 54919 70871
rect 54977 70825 55023 70871
rect 55081 70825 55127 70871
rect 55185 70825 55231 70871
rect 55289 70825 55335 70871
rect 55393 70825 55439 70871
rect 55497 70825 55543 70871
rect 55601 70825 55647 70871
rect 55705 70825 55751 70871
rect 55809 70825 55855 70871
rect 55913 70825 55959 70871
rect 56017 70825 56063 70871
rect 56121 70825 56167 70871
rect 56225 70825 56271 70871
rect 56329 70825 56375 70871
rect 56433 70825 56479 70871
rect 56537 70825 56583 70871
rect 56641 70825 56687 70871
rect 56745 70825 56791 70871
rect 56849 70825 56895 70871
rect 56953 70825 56999 70871
rect 57057 70825 57103 70871
rect 57161 70825 57207 70871
rect 57265 70825 57311 70871
rect 57369 70825 57415 70871
rect 57473 70825 57519 70871
rect 57577 70825 57623 70871
rect 57681 70825 57727 70871
rect 57785 70825 57831 70871
rect 57889 70825 57935 70871
rect 57993 70825 58039 70871
rect 58097 70825 58143 70871
rect 58201 70825 58247 70871
rect 58305 70825 58351 70871
rect 58409 70825 58455 70871
rect 58513 70825 58559 70871
rect 58617 70825 58663 70871
rect 58721 70825 58767 70871
rect 58825 70825 58871 70871
rect 58929 70825 58975 70871
rect 59033 70825 59079 70871
rect 59137 70825 59183 70871
rect 59241 70825 59287 70871
rect 59345 70825 59391 70871
rect 59449 70825 59495 70871
rect 59553 70825 59599 70871
rect 59657 70825 59703 70871
rect 59761 70825 59807 70871
rect 59865 70825 59911 70871
rect 59969 70825 60015 70871
rect 60073 70825 60119 70871
rect 60177 70825 60223 70871
rect 60281 70825 60327 70871
rect 60385 70825 60431 70871
rect 60489 70825 60535 70871
rect 60593 70825 60639 70871
rect 60697 70825 60743 70871
rect 60801 70825 60847 70871
rect 60905 70825 60951 70871
rect 61009 70825 61055 70871
rect 61113 70825 61159 70871
rect 61217 70825 61263 70871
rect 61321 70825 61367 70871
rect 61425 70825 61471 70871
rect 61529 70825 61575 70871
rect 61633 70825 61679 70871
rect 61737 70825 61783 70871
rect 61841 70825 61887 70871
rect 61945 70825 61991 70871
rect 62049 70825 62095 70871
rect 62153 70825 62199 70871
rect 62257 70825 62303 70871
rect 62361 70825 62407 70871
rect 62465 70825 62511 70871
rect 62569 70825 62615 70871
rect 62673 70825 62719 70871
rect 62777 70825 62823 70871
rect 62881 70825 62927 70871
rect 62985 70825 63031 70871
rect 63089 70825 63135 70871
rect 63193 70825 63239 70871
rect 63297 70825 63343 70871
rect 63401 70825 63447 70871
rect 63505 70825 63551 70871
rect 63609 70825 63655 70871
rect 63713 70825 63759 70871
rect 63817 70825 63863 70871
rect 63921 70825 63967 70871
rect 64025 70825 64071 70871
rect 64129 70825 64175 70871
rect 64233 70825 64279 70871
rect 64337 70825 64383 70871
rect 64441 70825 64487 70871
rect 64545 70825 64591 70871
rect 64649 70825 64695 70871
rect 64753 70825 64799 70871
rect 64857 70825 64903 70871
rect 64961 70825 65007 70871
rect 65065 70825 65111 70871
rect 65169 70825 65215 70871
rect 65273 70825 65319 70871
rect 65377 70825 65423 70871
rect 65481 70825 65527 70871
rect 65585 70825 65631 70871
rect 65689 70825 65735 70871
rect 65793 70825 65839 70871
rect 65897 70825 65943 70871
rect 66001 70825 66047 70871
rect 66105 70825 66151 70871
rect 66209 70825 66255 70871
rect 66313 70825 66359 70871
rect 66417 70825 66463 70871
rect 66521 70825 66567 70871
rect 66625 70825 66671 70871
rect 66729 70825 66775 70871
rect 66833 70825 66879 70871
rect 66937 70825 66983 70871
rect 67041 70825 67087 70871
rect 67145 70825 67191 70871
rect 67249 70825 67295 70871
rect 67353 70825 67399 70871
rect 67457 70825 67503 70871
rect 67561 70825 67607 70871
rect 67665 70825 67711 70871
rect 67769 70825 67815 70871
rect 67873 70825 67919 70871
rect 67977 70825 68023 70871
rect 68081 70825 68127 70871
rect 68185 70825 68231 70871
rect 68289 70825 68335 70871
rect 68393 70825 68439 70871
rect 68497 70825 68543 70871
rect 68601 70825 68647 70871
rect 68705 70825 68751 70871
rect 68809 70825 68855 70871
rect 68913 70825 68959 70871
rect 69017 70825 69063 70871
rect 69121 70825 69167 70871
rect 69225 70825 69271 70871
rect 69329 70825 69375 70871
rect 69433 70825 69479 70871
rect 69537 70825 69583 70871
rect 69641 70825 69687 70871
rect 69745 70825 69791 70871
rect 69849 70825 69895 70871
rect 13119 70721 13165 70767
rect 13223 70721 13269 70767
rect 13119 70617 13165 70663
rect 13223 70617 13269 70663
rect 13119 70513 13165 70559
rect 13223 70513 13269 70559
rect 13119 70409 13165 70455
rect 13223 70409 13269 70455
rect 13119 70305 13165 70351
rect 13223 70305 13269 70351
rect 13119 70201 13165 70247
rect 13223 70201 13269 70247
rect 13119 70097 13165 70143
rect 13223 70097 13269 70143
rect 13119 69993 13165 70039
rect 13223 69993 13269 70039
rect 13119 69889 13165 69935
rect 13223 69889 13269 69935
rect 13119 69785 13165 69831
rect 13223 69785 13269 69831
rect 69796 70674 69842 70720
rect 69900 70674 69946 70720
rect 69796 70570 69842 70616
rect 69900 70570 69946 70616
rect 69796 70466 69842 70512
rect 69900 70466 69946 70512
rect 69796 70362 69842 70408
rect 69900 70362 69946 70408
rect 69796 70258 69842 70304
rect 69900 70258 69946 70304
rect 69796 70154 69842 70200
rect 69900 70154 69946 70200
rect 69796 70050 69842 70096
rect 69900 70050 69946 70096
rect 69796 69900 69842 69946
rect 69900 69900 69946 69946
rect 70004 69900 70050 69946
rect 70108 69900 70154 69946
rect 70212 69900 70258 69946
rect 70316 69900 70362 69946
rect 70420 69900 70466 69946
rect 70524 69900 70570 69946
rect 70628 69900 70674 69946
rect 70824 69862 70870 69908
rect 70928 69862 70974 69908
rect 69796 69796 69842 69842
rect 69900 69796 69946 69842
rect 70004 69796 70050 69842
rect 70108 69796 70154 69842
rect 70212 69796 70258 69842
rect 70316 69796 70362 69842
rect 70420 69796 70466 69842
rect 70524 69796 70570 69842
rect 70628 69796 70674 69842
rect 13119 69681 13165 69727
rect 13223 69681 13269 69727
rect 13119 69577 13165 69623
rect 13223 69577 13269 69623
rect 13119 69473 13165 69519
rect 13223 69473 13269 69519
rect 13119 69369 13165 69415
rect 13223 69369 13269 69415
rect 13119 69265 13165 69311
rect 13223 69265 13269 69311
rect 13119 69161 13165 69207
rect 13223 69161 13269 69207
rect 13119 69057 13165 69103
rect 13223 69057 13269 69103
rect 13119 68953 13165 68999
rect 13223 68953 13269 68999
rect 13119 68849 13165 68895
rect 13223 68849 13269 68895
rect 13119 68745 13165 68791
rect 13223 68745 13269 68791
rect 13119 68641 13165 68687
rect 13223 68641 13269 68687
rect 13119 68537 13165 68583
rect 13223 68537 13269 68583
rect 13119 68433 13165 68479
rect 13223 68433 13269 68479
rect 13119 68329 13165 68375
rect 13223 68329 13269 68375
rect 13119 68225 13165 68271
rect 13223 68225 13269 68271
rect 13119 68121 13165 68167
rect 13223 68121 13269 68167
rect 13119 68017 13165 68063
rect 13223 68017 13269 68063
rect 13119 67913 13165 67959
rect 13223 67913 13269 67959
rect 13119 67809 13165 67855
rect 13223 67809 13269 67855
rect 13119 67705 13165 67751
rect 13223 67705 13269 67751
rect 13119 67601 13165 67647
rect 13223 67601 13269 67647
rect 13119 67497 13165 67543
rect 13223 67497 13269 67543
rect 13119 67393 13165 67439
rect 13223 67393 13269 67439
rect 13119 67289 13165 67335
rect 13223 67289 13269 67335
rect 13119 67185 13165 67231
rect 13223 67185 13269 67231
rect 13119 67081 13165 67127
rect 13223 67081 13269 67127
rect 13119 66977 13165 67023
rect 13223 66977 13269 67023
rect 13119 66873 13165 66919
rect 13223 66873 13269 66919
rect 13119 66769 13165 66815
rect 13223 66769 13269 66815
rect 13119 66665 13165 66711
rect 13223 66665 13269 66711
rect 13119 66561 13165 66607
rect 13223 66561 13269 66607
rect 13119 66457 13165 66503
rect 13223 66457 13269 66503
rect 13119 66353 13165 66399
rect 13223 66353 13269 66399
rect 13119 66249 13165 66295
rect 13223 66249 13269 66295
rect 13119 66145 13165 66191
rect 13223 66145 13269 66191
rect 13119 66041 13165 66087
rect 13223 66041 13269 66087
rect 13119 65937 13165 65983
rect 13223 65937 13269 65983
rect 13119 65833 13165 65879
rect 13223 65833 13269 65879
rect 13119 65729 13165 65775
rect 13223 65729 13269 65775
rect 13119 65625 13165 65671
rect 13223 65625 13269 65671
rect 13119 65521 13165 65567
rect 13223 65521 13269 65567
rect 13119 65417 13165 65463
rect 13223 65417 13269 65463
rect 13119 65313 13165 65359
rect 13223 65313 13269 65359
rect 13119 65209 13165 65255
rect 13223 65209 13269 65255
rect 13119 65105 13165 65151
rect 13223 65105 13269 65151
rect 13119 65001 13165 65047
rect 13223 65001 13269 65047
rect 13119 64897 13165 64943
rect 13223 64897 13269 64943
rect 13119 64793 13165 64839
rect 13223 64793 13269 64839
rect 13119 64689 13165 64735
rect 13223 64689 13269 64735
rect 13119 64585 13165 64631
rect 13223 64585 13269 64631
rect 13119 64481 13165 64527
rect 13223 64481 13269 64527
rect 13119 64377 13165 64423
rect 13223 64377 13269 64423
rect 13119 64273 13165 64319
rect 13223 64273 13269 64319
rect 13119 64169 13165 64215
rect 13223 64169 13269 64215
rect 13119 64065 13165 64111
rect 13223 64065 13269 64111
rect 13119 63961 13165 64007
rect 13223 63961 13269 64007
rect 13119 63857 13165 63903
rect 13223 63857 13269 63903
rect 13119 63753 13165 63799
rect 13223 63753 13269 63799
rect 13119 63649 13165 63695
rect 13223 63649 13269 63695
rect 13119 63545 13165 63591
rect 13223 63545 13269 63591
rect 13119 63441 13165 63487
rect 13223 63441 13269 63487
rect 13119 63337 13165 63383
rect 13223 63337 13269 63383
rect 13119 63233 13165 63279
rect 13223 63233 13269 63279
rect 13119 63129 13165 63175
rect 13223 63129 13269 63175
rect 13119 63025 13165 63071
rect 13223 63025 13269 63071
rect 13119 62921 13165 62967
rect 13223 62921 13269 62967
rect 13119 62817 13165 62863
rect 13223 62817 13269 62863
rect 13119 62713 13165 62759
rect 13223 62713 13269 62759
rect 13119 62609 13165 62655
rect 13223 62609 13269 62655
rect 13119 62505 13165 62551
rect 13223 62505 13269 62551
rect 13119 62401 13165 62447
rect 13223 62401 13269 62447
rect 13119 62297 13165 62343
rect 13223 62297 13269 62343
rect 13119 62193 13165 62239
rect 13223 62193 13269 62239
rect 13119 62089 13165 62135
rect 13223 62089 13269 62135
rect 13119 61985 13165 62031
rect 13223 61985 13269 62031
rect 13119 61881 13165 61927
rect 13223 61881 13269 61927
rect 13119 61777 13165 61823
rect 13223 61777 13269 61823
rect 13119 61673 13165 61719
rect 13223 61673 13269 61719
rect 13119 61569 13165 61615
rect 13223 61569 13269 61615
rect 13119 61465 13165 61511
rect 13223 61465 13269 61511
rect 13119 61361 13165 61407
rect 13223 61361 13269 61407
rect 13119 61257 13165 61303
rect 13223 61257 13269 61303
rect 13119 61153 13165 61199
rect 13223 61153 13269 61199
rect 13119 61049 13165 61095
rect 13223 61049 13269 61095
rect 13119 60945 13165 60991
rect 13223 60945 13269 60991
rect 13119 60841 13165 60887
rect 13223 60841 13269 60887
rect 13119 60737 13165 60783
rect 13223 60737 13269 60783
rect 13119 60633 13165 60679
rect 13223 60633 13269 60679
rect 13119 60529 13165 60575
rect 13223 60529 13269 60575
rect 13119 60425 13165 60471
rect 13223 60425 13269 60471
rect 13119 60321 13165 60367
rect 13223 60321 13269 60367
rect 13119 60217 13165 60263
rect 13223 60217 13269 60263
rect 13119 60113 13165 60159
rect 13223 60113 13269 60159
rect 13119 60009 13165 60055
rect 13223 60009 13269 60055
rect 13119 59905 13165 59951
rect 13223 59905 13269 59951
rect 13119 59801 13165 59847
rect 13223 59801 13269 59847
rect 13119 59697 13165 59743
rect 13223 59697 13269 59743
rect 13119 59593 13165 59639
rect 13223 59593 13269 59639
rect 13119 59489 13165 59535
rect 13223 59489 13269 59535
rect 13119 59385 13165 59431
rect 13223 59385 13269 59431
rect 13119 59281 13165 59327
rect 13223 59281 13269 59327
rect 13119 59177 13165 59223
rect 13223 59177 13269 59223
rect 13119 59073 13165 59119
rect 13223 59073 13269 59119
rect 13119 58969 13165 59015
rect 13223 58969 13269 59015
rect 13119 58865 13165 58911
rect 13223 58865 13269 58911
rect 13119 58761 13165 58807
rect 13223 58761 13269 58807
rect 13119 58657 13165 58703
rect 13223 58657 13269 58703
rect 13119 58553 13165 58599
rect 13223 58553 13269 58599
rect 13119 58449 13165 58495
rect 13223 58449 13269 58495
rect 13119 58345 13165 58391
rect 13223 58345 13269 58391
rect 13119 58241 13165 58287
rect 13223 58241 13269 58287
rect 13119 58137 13165 58183
rect 13223 58137 13269 58183
rect 13119 58033 13165 58079
rect 13223 58033 13269 58079
rect 13119 57929 13165 57975
rect 13223 57929 13269 57975
rect 13119 57825 13165 57871
rect 13223 57825 13269 57871
rect 13119 57721 13165 57767
rect 13223 57721 13269 57767
rect 13119 57617 13165 57663
rect 13223 57617 13269 57663
rect 13119 57513 13165 57559
rect 13223 57513 13269 57559
rect 13119 57409 13165 57455
rect 13223 57409 13269 57455
rect 13119 57305 13165 57351
rect 13223 57305 13269 57351
rect 13119 57201 13165 57247
rect 13223 57201 13269 57247
rect 13119 57097 13165 57143
rect 13223 57097 13269 57143
rect 13119 56993 13165 57039
rect 13223 56993 13269 57039
rect 13119 56889 13165 56935
rect 13223 56889 13269 56935
rect 13119 56785 13165 56831
rect 13223 56785 13269 56831
rect 13119 56681 13165 56727
rect 13223 56681 13269 56727
rect 13119 56577 13165 56623
rect 13223 56577 13269 56623
rect 13119 56473 13165 56519
rect 13223 56473 13269 56519
rect 13119 56369 13165 56415
rect 13223 56369 13269 56415
rect 13119 56265 13165 56311
rect 13223 56265 13269 56311
rect 13119 56161 13165 56207
rect 13223 56161 13269 56207
rect 13119 56057 13165 56103
rect 13223 56057 13269 56103
rect 13119 55953 13165 55999
rect 13223 55953 13269 55999
rect 13119 55849 13165 55895
rect 13223 55849 13269 55895
rect 13119 55745 13165 55791
rect 13223 55745 13269 55791
rect 13119 55641 13165 55687
rect 13223 55641 13269 55687
rect 13119 55537 13165 55583
rect 13223 55537 13269 55583
rect 13119 55433 13165 55479
rect 13223 55433 13269 55479
rect 13119 55329 13165 55375
rect 13223 55329 13269 55375
rect 13119 55225 13165 55271
rect 13223 55225 13269 55271
rect 13119 55121 13165 55167
rect 13223 55121 13269 55167
rect 13119 55017 13165 55063
rect 13223 55017 13269 55063
rect 13119 54913 13165 54959
rect 13223 54913 13269 54959
rect 13119 54809 13165 54855
rect 13223 54809 13269 54855
rect 13119 54705 13165 54751
rect 13223 54705 13269 54751
rect 13119 54601 13165 54647
rect 13223 54601 13269 54647
rect 13119 54497 13165 54543
rect 13223 54497 13269 54543
rect 13119 54393 13165 54439
rect 13223 54393 13269 54439
rect 13119 54289 13165 54335
rect 13223 54289 13269 54335
rect 13119 54185 13165 54231
rect 13223 54185 13269 54231
rect 13119 54081 13165 54127
rect 13223 54081 13269 54127
rect 13119 53977 13165 54023
rect 13223 53977 13269 54023
rect 13119 53873 13165 53919
rect 13223 53873 13269 53919
rect 13119 53769 13165 53815
rect 13223 53769 13269 53815
rect 13119 53665 13165 53711
rect 13223 53665 13269 53711
rect 13119 53561 13165 53607
rect 13223 53561 13269 53607
rect 13119 53457 13165 53503
rect 13223 53457 13269 53503
rect 13119 53353 13165 53399
rect 13223 53353 13269 53399
rect 13119 53249 13165 53295
rect 13223 53249 13269 53295
rect 13119 53145 13165 53191
rect 13223 53145 13269 53191
rect 13119 53041 13165 53087
rect 13223 53041 13269 53087
rect 13119 52937 13165 52983
rect 13223 52937 13269 52983
rect 13119 52833 13165 52879
rect 13223 52833 13269 52879
rect 13119 52729 13165 52775
rect 13223 52729 13269 52775
rect 13119 52625 13165 52671
rect 13223 52625 13269 52671
rect 13119 52521 13165 52567
rect 13223 52521 13269 52567
rect 13119 52417 13165 52463
rect 13223 52417 13269 52463
rect 13119 52313 13165 52359
rect 13223 52313 13269 52359
rect 13119 52209 13165 52255
rect 13223 52209 13269 52255
rect 13119 52105 13165 52151
rect 13223 52105 13269 52151
rect 13119 52001 13165 52047
rect 13223 52001 13269 52047
rect 13119 51897 13165 51943
rect 13223 51897 13269 51943
rect 13119 51793 13165 51839
rect 13223 51793 13269 51839
rect 13119 51689 13165 51735
rect 13223 51689 13269 51735
rect 13119 51585 13165 51631
rect 13223 51585 13269 51631
rect 13119 51481 13165 51527
rect 13223 51481 13269 51527
rect 13119 51377 13165 51423
rect 13223 51377 13269 51423
rect 13119 51273 13165 51319
rect 13223 51273 13269 51319
rect 13119 51169 13165 51215
rect 13223 51169 13269 51215
rect 13119 51065 13165 51111
rect 13223 51065 13269 51111
rect 13119 50961 13165 51007
rect 13223 50961 13269 51007
rect 13119 50857 13165 50903
rect 13223 50857 13269 50903
rect 13119 50753 13165 50799
rect 13223 50753 13269 50799
rect 13119 50649 13165 50695
rect 13223 50649 13269 50695
rect 13119 50545 13165 50591
rect 13223 50545 13269 50591
rect 13119 50441 13165 50487
rect 13223 50441 13269 50487
rect 13119 50337 13165 50383
rect 13223 50337 13269 50383
rect 13119 50233 13165 50279
rect 13223 50233 13269 50279
rect 13119 50129 13165 50175
rect 13223 50129 13269 50175
rect 13119 50025 13165 50071
rect 13223 50025 13269 50071
rect 13119 49921 13165 49967
rect 13223 49921 13269 49967
rect 13119 49817 13165 49863
rect 13223 49817 13269 49863
rect 13119 49713 13165 49759
rect 13223 49713 13269 49759
rect 13119 49609 13165 49655
rect 13223 49609 13269 49655
rect 13119 49505 13165 49551
rect 13223 49505 13269 49551
rect 13119 49401 13165 49447
rect 13223 49401 13269 49447
rect 13119 49297 13165 49343
rect 13223 49297 13269 49343
rect 13119 49193 13165 49239
rect 13223 49193 13269 49239
rect 13119 49089 13165 49135
rect 13223 49089 13269 49135
rect 13119 48985 13165 49031
rect 13223 48985 13269 49031
rect 13119 48881 13165 48927
rect 13223 48881 13269 48927
rect 13119 48777 13165 48823
rect 13223 48777 13269 48823
rect 13119 48673 13165 48719
rect 13223 48673 13269 48719
rect 13119 48569 13165 48615
rect 13223 48569 13269 48615
rect 13119 48465 13165 48511
rect 13223 48465 13269 48511
rect 13119 48361 13165 48407
rect 13223 48361 13269 48407
rect 13119 48257 13165 48303
rect 13223 48257 13269 48303
rect 13119 48153 13165 48199
rect 13223 48153 13269 48199
rect 13119 48049 13165 48095
rect 13223 48049 13269 48095
rect 13119 47945 13165 47991
rect 13223 47945 13269 47991
rect 13119 47841 13165 47887
rect 13223 47841 13269 47887
rect 13119 47737 13165 47783
rect 13223 47737 13269 47783
rect 13119 47633 13165 47679
rect 13223 47633 13269 47679
rect 13119 47529 13165 47575
rect 13223 47529 13269 47575
rect 13119 47425 13165 47471
rect 13223 47425 13269 47471
rect 13119 47321 13165 47367
rect 13223 47321 13269 47367
rect 13119 47217 13165 47263
rect 13223 47217 13269 47263
rect 13119 47113 13165 47159
rect 13223 47113 13269 47159
rect 13119 47009 13165 47055
rect 13223 47009 13269 47055
rect 13119 46905 13165 46951
rect 13223 46905 13269 46951
rect 13119 46801 13165 46847
rect 13223 46801 13269 46847
rect 13119 46697 13165 46743
rect 13223 46697 13269 46743
rect 13119 46593 13165 46639
rect 13223 46593 13269 46639
rect 13119 46489 13165 46535
rect 13223 46489 13269 46535
rect 13119 46385 13165 46431
rect 13223 46385 13269 46431
rect 13119 46281 13165 46327
rect 13223 46281 13269 46327
rect 13119 46177 13165 46223
rect 13223 46177 13269 46223
rect 13119 46073 13165 46119
rect 13223 46073 13269 46119
rect 13119 45969 13165 46015
rect 13223 45969 13269 46015
rect 13119 45865 13165 45911
rect 13223 45865 13269 45911
rect 13119 45761 13165 45807
rect 13223 45761 13269 45807
rect 13119 45657 13165 45703
rect 13223 45657 13269 45703
rect 13119 45553 13165 45599
rect 13223 45553 13269 45599
rect 13119 45449 13165 45495
rect 13223 45449 13269 45495
rect 13119 45345 13165 45391
rect 13223 45345 13269 45391
rect 13119 45241 13165 45287
rect 13223 45241 13269 45287
rect 13119 45137 13165 45183
rect 13223 45137 13269 45183
rect 13119 45033 13165 45079
rect 13223 45033 13269 45079
rect 70824 69758 70870 69804
rect 70928 69758 70974 69804
rect 70824 69654 70870 69700
rect 70928 69654 70974 69700
rect 70824 69550 70870 69596
rect 70928 69550 70974 69596
rect 70824 69446 70870 69492
rect 70928 69446 70974 69492
rect 70824 69342 70870 69388
rect 70928 69342 70974 69388
rect 70824 69238 70870 69284
rect 70928 69238 70974 69284
rect 70824 69134 70870 69180
rect 70928 69134 70974 69180
rect 70824 69030 70870 69076
rect 70928 69030 70974 69076
rect 70824 68926 70870 68972
rect 70928 68926 70974 68972
rect 70824 68822 70870 68868
rect 70928 68822 70974 68868
rect 70824 68718 70870 68764
rect 70928 68718 70974 68764
rect 70824 68614 70870 68660
rect 70928 68614 70974 68660
rect 70824 68510 70870 68556
rect 70928 68510 70974 68556
rect 70824 68406 70870 68452
rect 70928 68406 70974 68452
rect 70824 68302 70870 68348
rect 70928 68302 70974 68348
rect 70824 68198 70870 68244
rect 70928 68198 70974 68244
rect 70824 68094 70870 68140
rect 70928 68094 70974 68140
rect 70824 67990 70870 68036
rect 70928 67990 70974 68036
rect 70824 67886 70870 67932
rect 70928 67886 70974 67932
rect 70824 67782 70870 67828
rect 70928 67782 70974 67828
rect 70824 67678 70870 67724
rect 70928 67678 70974 67724
rect 70824 67574 70870 67620
rect 70928 67574 70974 67620
rect 70824 67470 70870 67516
rect 70928 67470 70974 67516
rect 70824 67366 70870 67412
rect 70928 67366 70974 67412
rect 70824 67262 70870 67308
rect 70928 67262 70974 67308
rect 70824 67158 70870 67204
rect 70928 67158 70974 67204
rect 70824 67054 70870 67100
rect 70928 67054 70974 67100
rect 70824 66950 70870 66996
rect 70928 66950 70974 66996
rect 70824 66846 70870 66892
rect 70928 66846 70974 66892
rect 70824 66742 70870 66788
rect 70928 66742 70974 66788
rect 70824 66638 70870 66684
rect 70928 66638 70974 66684
rect 70824 66534 70870 66580
rect 70928 66534 70974 66580
rect 70824 66430 70870 66476
rect 70928 66430 70974 66476
rect 70824 66326 70870 66372
rect 70928 66326 70974 66372
rect 70824 66222 70870 66268
rect 70928 66222 70974 66268
rect 70824 66118 70870 66164
rect 70928 66118 70974 66164
rect 70824 66014 70870 66060
rect 70928 66014 70974 66060
rect 70824 65910 70870 65956
rect 70928 65910 70974 65956
rect 70824 65806 70870 65852
rect 70928 65806 70974 65852
rect 70824 65702 70870 65748
rect 70928 65702 70974 65748
rect 70824 65598 70870 65644
rect 70928 65598 70974 65644
rect 70824 65494 70870 65540
rect 70928 65494 70974 65540
rect 70824 65390 70870 65436
rect 70928 65390 70974 65436
rect 70824 65286 70870 65332
rect 70928 65286 70974 65332
rect 70824 65182 70870 65228
rect 70928 65182 70974 65228
rect 70824 65078 70870 65124
rect 70928 65078 70974 65124
rect 70824 64974 70870 65020
rect 70928 64974 70974 65020
rect 70824 64870 70870 64916
rect 70928 64870 70974 64916
rect 70824 64766 70870 64812
rect 70928 64766 70974 64812
rect 70824 64662 70870 64708
rect 70928 64662 70974 64708
rect 70824 64558 70870 64604
rect 70928 64558 70974 64604
rect 70824 64454 70870 64500
rect 70928 64454 70974 64500
rect 70824 64350 70870 64396
rect 70928 64350 70974 64396
rect 70824 64246 70870 64292
rect 70928 64246 70974 64292
rect 70824 64142 70870 64188
rect 70928 64142 70974 64188
rect 70824 64038 70870 64084
rect 70928 64038 70974 64084
rect 70824 63934 70870 63980
rect 70928 63934 70974 63980
rect 70824 63830 70870 63876
rect 70928 63830 70974 63876
rect 70824 63726 70870 63772
rect 70928 63726 70974 63772
rect 70824 63622 70870 63668
rect 70928 63622 70974 63668
rect 70824 63518 70870 63564
rect 70928 63518 70974 63564
rect 70824 63414 70870 63460
rect 70928 63414 70974 63460
rect 70824 63310 70870 63356
rect 70928 63310 70974 63356
rect 70824 63206 70870 63252
rect 70928 63206 70974 63252
rect 70824 63102 70870 63148
rect 70928 63102 70974 63148
rect 70824 62998 70870 63044
rect 70928 62998 70974 63044
rect 70824 62894 70870 62940
rect 70928 62894 70974 62940
rect 70824 62790 70870 62836
rect 70928 62790 70974 62836
rect 70824 62686 70870 62732
rect 70928 62686 70974 62732
rect 70824 62582 70870 62628
rect 70928 62582 70974 62628
rect 70824 62478 70870 62524
rect 70928 62478 70974 62524
rect 70824 62374 70870 62420
rect 70928 62374 70974 62420
rect 70824 62270 70870 62316
rect 70928 62270 70974 62316
rect 70824 62166 70870 62212
rect 70928 62166 70974 62212
rect 70824 62062 70870 62108
rect 70928 62062 70974 62108
rect 70824 61958 70870 62004
rect 70928 61958 70974 62004
rect 70824 61854 70870 61900
rect 70928 61854 70974 61900
rect 70824 61750 70870 61796
rect 70928 61750 70974 61796
rect 70824 61646 70870 61692
rect 70928 61646 70974 61692
rect 70824 61542 70870 61588
rect 70928 61542 70974 61588
rect 70824 61438 70870 61484
rect 70928 61438 70974 61484
rect 70824 61334 70870 61380
rect 70928 61334 70974 61380
rect 70824 61230 70870 61276
rect 70928 61230 70974 61276
rect 70824 61126 70870 61172
rect 70928 61126 70974 61172
rect 70824 61022 70870 61068
rect 70928 61022 70974 61068
rect 70824 60918 70870 60964
rect 70928 60918 70974 60964
rect 70824 60814 70870 60860
rect 70928 60814 70974 60860
rect 70824 60710 70870 60756
rect 70928 60710 70974 60756
rect 70824 60606 70870 60652
rect 70928 60606 70974 60652
rect 70824 60502 70870 60548
rect 70928 60502 70974 60548
rect 70824 60398 70870 60444
rect 70928 60398 70974 60444
rect 70824 60294 70870 60340
rect 70928 60294 70974 60340
rect 70824 60190 70870 60236
rect 70928 60190 70974 60236
rect 70824 60086 70870 60132
rect 70928 60086 70974 60132
rect 70824 59982 70870 60028
rect 70928 59982 70974 60028
rect 70824 59878 70870 59924
rect 70928 59878 70974 59924
rect 70824 59774 70870 59820
rect 70928 59774 70974 59820
rect 70824 59670 70870 59716
rect 70928 59670 70974 59716
rect 70824 59566 70870 59612
rect 70928 59566 70974 59612
rect 70824 59462 70870 59508
rect 70928 59462 70974 59508
rect 70824 59358 70870 59404
rect 70928 59358 70974 59404
rect 70824 59254 70870 59300
rect 70928 59254 70974 59300
rect 70824 59150 70870 59196
rect 70928 59150 70974 59196
rect 70824 59046 70870 59092
rect 70928 59046 70974 59092
rect 70824 58942 70870 58988
rect 70928 58942 70974 58988
rect 70824 58838 70870 58884
rect 70928 58838 70974 58884
rect 70824 58734 70870 58780
rect 70928 58734 70974 58780
rect 70824 58630 70870 58676
rect 70928 58630 70974 58676
rect 70824 58526 70870 58572
rect 70928 58526 70974 58572
rect 70824 58422 70870 58468
rect 70928 58422 70974 58468
rect 70824 58318 70870 58364
rect 70928 58318 70974 58364
rect 70824 58214 70870 58260
rect 70928 58214 70974 58260
rect 70824 58110 70870 58156
rect 70928 58110 70974 58156
rect 70824 58006 70870 58052
rect 70928 58006 70974 58052
rect 70824 57902 70870 57948
rect 70928 57902 70974 57948
rect 70824 57798 70870 57844
rect 70928 57798 70974 57844
rect 70824 57694 70870 57740
rect 70928 57694 70974 57740
rect 70824 57590 70870 57636
rect 70928 57590 70974 57636
rect 70824 57486 70870 57532
rect 70928 57486 70974 57532
rect 70824 57382 70870 57428
rect 70928 57382 70974 57428
rect 70824 57278 70870 57324
rect 70928 57278 70974 57324
rect 70824 57174 70870 57220
rect 70928 57174 70974 57220
rect 70824 57070 70870 57116
rect 70928 57070 70974 57116
rect 70824 56966 70870 57012
rect 70928 56966 70974 57012
rect 70824 56862 70870 56908
rect 70928 56862 70974 56908
rect 70824 56758 70870 56804
rect 70928 56758 70974 56804
rect 70824 56654 70870 56700
rect 70928 56654 70974 56700
rect 70824 56550 70870 56596
rect 70928 56550 70974 56596
rect 70824 56446 70870 56492
rect 70928 56446 70974 56492
rect 70824 56342 70870 56388
rect 70928 56342 70974 56388
rect 70824 56238 70870 56284
rect 70928 56238 70974 56284
rect 70824 56134 70870 56180
rect 70928 56134 70974 56180
rect 70824 56030 70870 56076
rect 70928 56030 70974 56076
rect 70824 55926 70870 55972
rect 70928 55926 70974 55972
rect 70824 55822 70870 55868
rect 70928 55822 70974 55868
rect 70824 55718 70870 55764
rect 70928 55718 70974 55764
rect 70824 55614 70870 55660
rect 70928 55614 70974 55660
rect 70824 55510 70870 55556
rect 70928 55510 70974 55556
rect 70824 55406 70870 55452
rect 70928 55406 70974 55452
rect 70824 55302 70870 55348
rect 70928 55302 70974 55348
rect 70824 55198 70870 55244
rect 70928 55198 70974 55244
rect 70824 55094 70870 55140
rect 70928 55094 70974 55140
rect 70824 54990 70870 55036
rect 70928 54990 70974 55036
rect 70824 54886 70870 54932
rect 70928 54886 70974 54932
rect 70824 54782 70870 54828
rect 70928 54782 70974 54828
rect 70824 54678 70870 54724
rect 70928 54678 70974 54724
rect 70824 54574 70870 54620
rect 70928 54574 70974 54620
rect 70824 54470 70870 54516
rect 70928 54470 70974 54516
rect 70824 54366 70870 54412
rect 70928 54366 70974 54412
rect 70824 54262 70870 54308
rect 70928 54262 70974 54308
rect 70824 54158 70870 54204
rect 70928 54158 70974 54204
rect 70824 54054 70870 54100
rect 70928 54054 70974 54100
rect 70824 53950 70870 53996
rect 70928 53950 70974 53996
rect 70824 53846 70870 53892
rect 70928 53846 70974 53892
rect 70824 53742 70870 53788
rect 70928 53742 70974 53788
rect 70824 53638 70870 53684
rect 70928 53638 70974 53684
rect 70824 53534 70870 53580
rect 70928 53534 70974 53580
rect 70824 53430 70870 53476
rect 70928 53430 70974 53476
rect 70824 53326 70870 53372
rect 70928 53326 70974 53372
rect 70824 53222 70870 53268
rect 70928 53222 70974 53268
rect 70824 53118 70870 53164
rect 70928 53118 70974 53164
rect 70824 53014 70870 53060
rect 70928 53014 70974 53060
rect 70824 52910 70870 52956
rect 70928 52910 70974 52956
rect 70824 52806 70870 52852
rect 70928 52806 70974 52852
rect 70824 52702 70870 52748
rect 70928 52702 70974 52748
rect 70824 52598 70870 52644
rect 70928 52598 70974 52644
rect 70824 52494 70870 52540
rect 70928 52494 70974 52540
rect 70824 52390 70870 52436
rect 70928 52390 70974 52436
rect 70824 52286 70870 52332
rect 70928 52286 70974 52332
rect 70824 52182 70870 52228
rect 70928 52182 70974 52228
rect 70824 52078 70870 52124
rect 70928 52078 70974 52124
rect 70824 51974 70870 52020
rect 70928 51974 70974 52020
rect 70824 51870 70870 51916
rect 70928 51870 70974 51916
rect 70824 51766 70870 51812
rect 70928 51766 70974 51812
rect 70824 51662 70870 51708
rect 70928 51662 70974 51708
rect 70824 51558 70870 51604
rect 70928 51558 70974 51604
rect 70824 51454 70870 51500
rect 70928 51454 70974 51500
rect 70824 51350 70870 51396
rect 70928 51350 70974 51396
rect 70824 51246 70870 51292
rect 70928 51246 70974 51292
rect 70824 51142 70870 51188
rect 70928 51142 70974 51188
rect 70824 51038 70870 51084
rect 70928 51038 70974 51084
rect 70824 50934 70870 50980
rect 70928 50934 70974 50980
rect 70824 50830 70870 50876
rect 70928 50830 70974 50876
rect 70824 50726 70870 50772
rect 70928 50726 70974 50772
rect 70824 50622 70870 50668
rect 70928 50622 70974 50668
rect 70824 50518 70870 50564
rect 70928 50518 70974 50564
rect 70824 50414 70870 50460
rect 70928 50414 70974 50460
rect 70824 50310 70870 50356
rect 70928 50310 70974 50356
rect 70824 50206 70870 50252
rect 70928 50206 70974 50252
rect 70824 50102 70870 50148
rect 70928 50102 70974 50148
rect 70824 49998 70870 50044
rect 70928 49998 70974 50044
rect 70824 49894 70870 49940
rect 70928 49894 70974 49940
rect 70824 49790 70870 49836
rect 70928 49790 70974 49836
rect 70824 49686 70870 49732
rect 70928 49686 70974 49732
rect 70824 49582 70870 49628
rect 70928 49582 70974 49628
rect 70824 49478 70870 49524
rect 70928 49478 70974 49524
rect 70824 49374 70870 49420
rect 70928 49374 70974 49420
rect 70824 49270 70870 49316
rect 70928 49270 70974 49316
rect 70824 49166 70870 49212
rect 70928 49166 70974 49212
rect 70824 49062 70870 49108
rect 70928 49062 70974 49108
rect 70824 48958 70870 49004
rect 70928 48958 70974 49004
rect 70824 48854 70870 48900
rect 70928 48854 70974 48900
rect 70824 48750 70870 48796
rect 70928 48750 70974 48796
rect 70824 48646 70870 48692
rect 70928 48646 70974 48692
rect 70824 48542 70870 48588
rect 70928 48542 70974 48588
rect 70824 48438 70870 48484
rect 70928 48438 70974 48484
rect 70824 48334 70870 48380
rect 70928 48334 70974 48380
rect 70824 48230 70870 48276
rect 70928 48230 70974 48276
rect 70824 48126 70870 48172
rect 70928 48126 70974 48172
rect 70824 48022 70870 48068
rect 70928 48022 70974 48068
rect 70824 47918 70870 47964
rect 70928 47918 70974 47964
rect 70824 47814 70870 47860
rect 70928 47814 70974 47860
rect 70824 47710 70870 47756
rect 70928 47710 70974 47756
rect 70824 47606 70870 47652
rect 70928 47606 70974 47652
rect 70824 47502 70870 47548
rect 70928 47502 70974 47548
rect 70824 47398 70870 47444
rect 70928 47398 70974 47444
rect 70824 47294 70870 47340
rect 70928 47294 70974 47340
rect 70824 47190 70870 47236
rect 70928 47190 70974 47236
rect 70824 47086 70870 47132
rect 70928 47086 70974 47132
rect 70824 46982 70870 47028
rect 70928 46982 70974 47028
rect 70824 46878 70870 46924
rect 70928 46878 70974 46924
rect 70824 46774 70870 46820
rect 70928 46774 70974 46820
rect 70824 46670 70870 46716
rect 70928 46670 70974 46716
rect 70824 46566 70870 46612
rect 70928 46566 70974 46612
rect 70824 46462 70870 46508
rect 70928 46462 70974 46508
rect 70824 46358 70870 46404
rect 70928 46358 70974 46404
rect 70824 46254 70870 46300
rect 70928 46254 70974 46300
rect 70824 46150 70870 46196
rect 70928 46150 70974 46196
rect 70824 46046 70870 46092
rect 70928 46046 70974 46092
rect 70824 45942 70870 45988
rect 70928 45942 70974 45988
rect 70824 45838 70870 45884
rect 70928 45838 70974 45884
rect 70824 45734 70870 45780
rect 70928 45734 70974 45780
rect 70824 45630 70870 45676
rect 70928 45630 70974 45676
rect 70824 45526 70870 45572
rect 70928 45526 70974 45572
rect 70824 45422 70870 45468
rect 70928 45422 70974 45468
rect 70824 45318 70870 45364
rect 70928 45318 70974 45364
rect 70824 45214 70870 45260
rect 70928 45214 70974 45260
rect 70824 45110 70870 45156
rect 70928 45110 70974 45156
rect 70824 45006 70870 45052
rect 70928 45006 70974 45052
rect 70824 44902 70870 44948
rect 70928 44902 70974 44948
rect 13254 44778 13300 44824
rect 70824 44798 70870 44844
rect 70928 44798 70974 44844
rect 13386 44646 13432 44692
rect 70824 44694 70870 44740
rect 70928 44694 70974 44740
rect 70824 44590 70870 44636
rect 70928 44590 70974 44636
rect 13518 44514 13564 44560
rect 70824 44486 70870 44532
rect 70928 44486 70974 44532
rect 13650 44382 13696 44428
rect 70824 44382 70870 44428
rect 70928 44382 70974 44428
rect 13782 44250 13828 44296
rect 70824 44278 70870 44324
rect 70928 44278 70974 44324
rect 70824 44174 70870 44220
rect 70928 44174 70974 44220
rect 13914 44118 13960 44164
rect 70824 44070 70870 44116
rect 70928 44070 70974 44116
rect 14046 43986 14092 44032
rect 70824 43966 70870 44012
rect 70928 43966 70974 44012
rect 14178 43854 14224 43900
rect 70824 43862 70870 43908
rect 70928 43862 70974 43908
rect 14310 43722 14356 43768
rect 70824 43758 70870 43804
rect 70928 43758 70974 43804
rect 70824 43654 70870 43700
rect 70928 43654 70974 43700
rect 14442 43590 14488 43636
rect 70824 43550 70870 43596
rect 70928 43550 70974 43596
rect 14574 43458 14620 43504
rect 70824 43446 70870 43492
rect 70928 43446 70974 43492
rect 14706 43326 14752 43372
rect 70824 43342 70870 43388
rect 70928 43342 70974 43388
rect 14838 43194 14884 43240
rect 70824 43238 70870 43284
rect 70928 43238 70974 43284
rect 70824 43134 70870 43180
rect 70928 43134 70974 43180
rect 14970 43062 15016 43108
rect 70824 43030 70870 43076
rect 70928 43030 70974 43076
rect 15102 42930 15148 42976
rect 70824 42926 70870 42972
rect 70928 42926 70974 42972
rect 15234 42798 15280 42844
rect 70824 42822 70870 42868
rect 70928 42822 70974 42868
rect 15366 42666 15412 42712
rect 70824 42718 70870 42764
rect 70928 42718 70974 42764
rect 70824 42614 70870 42660
rect 70928 42614 70974 42660
rect 15498 42534 15544 42580
rect 70824 42510 70870 42556
rect 70928 42510 70974 42556
rect 15630 42402 15676 42448
rect 70824 42406 70870 42452
rect 70928 42406 70974 42452
rect 15762 42270 15808 42316
rect 70824 42302 70870 42348
rect 70928 42302 70974 42348
rect 70824 42198 70870 42244
rect 70928 42198 70974 42244
rect 15894 42138 15940 42184
rect 70824 42094 70870 42140
rect 70928 42094 70974 42140
rect 16026 42006 16072 42052
rect 70824 41990 70870 42036
rect 70928 41990 70974 42036
rect 16158 41874 16204 41920
rect 70824 41886 70870 41932
rect 70928 41886 70974 41932
rect 16290 41742 16336 41788
rect 70824 41782 70870 41828
rect 70928 41782 70974 41828
rect 70824 41678 70870 41724
rect 70928 41678 70974 41724
rect 16422 41610 16468 41656
rect 70824 41574 70870 41620
rect 70928 41574 70974 41620
rect 16554 41478 16600 41524
rect 70824 41470 70870 41516
rect 70928 41470 70974 41516
rect 16686 41346 16732 41392
rect 70824 41366 70870 41412
rect 70928 41366 70974 41412
rect 16818 41214 16864 41260
rect 70824 41262 70870 41308
rect 70928 41262 70974 41308
rect 70824 41158 70870 41204
rect 70928 41158 70974 41204
rect 16950 41082 16996 41128
rect 70824 41054 70870 41100
rect 70928 41054 70974 41100
rect 17082 40950 17128 40996
rect 70824 40950 70870 40996
rect 70928 40950 70974 40996
rect 17214 40818 17260 40864
rect 70824 40846 70870 40892
rect 70928 40846 70974 40892
rect 70824 40742 70870 40788
rect 70928 40742 70974 40788
rect 17346 40686 17392 40732
rect 70824 40638 70870 40684
rect 70928 40638 70974 40684
rect 17478 40554 17524 40600
rect 70824 40534 70870 40580
rect 70928 40534 70974 40580
rect 17610 40422 17656 40468
rect 70824 40430 70870 40476
rect 70928 40430 70974 40476
rect 17742 40290 17788 40336
rect 70824 40326 70870 40372
rect 70928 40326 70974 40372
rect 70824 40222 70870 40268
rect 70928 40222 70974 40268
rect 17874 40158 17920 40204
rect 70824 40118 70870 40164
rect 70928 40118 70974 40164
rect 18006 40026 18052 40072
rect 70824 40014 70870 40060
rect 70928 40014 70974 40060
rect 18138 39894 18184 39940
rect 70824 39910 70870 39956
rect 70928 39910 70974 39956
rect 18270 39762 18316 39808
rect 70824 39806 70870 39852
rect 70928 39806 70974 39852
rect 70824 39702 70870 39748
rect 70928 39702 70974 39748
rect 18402 39630 18448 39676
rect 70824 39598 70870 39644
rect 70928 39598 70974 39644
rect 18534 39498 18580 39544
rect 70824 39494 70870 39540
rect 70928 39494 70974 39540
rect 18666 39366 18712 39412
rect 70824 39390 70870 39436
rect 70928 39390 70974 39436
rect 18798 39234 18844 39280
rect 70824 39286 70870 39332
rect 70928 39286 70974 39332
rect 70824 39182 70870 39228
rect 70928 39182 70974 39228
rect 18930 39102 18976 39148
rect 70824 39078 70870 39124
rect 70928 39078 70974 39124
rect 19062 38970 19108 39016
rect 70824 38974 70870 39020
rect 70928 38974 70974 39020
rect 19194 38838 19240 38884
rect 70824 38870 70870 38916
rect 70928 38870 70974 38916
rect 70824 38766 70870 38812
rect 70928 38766 70974 38812
rect 19326 38706 19372 38752
rect 70824 38662 70870 38708
rect 70928 38662 70974 38708
rect 19458 38574 19504 38620
rect 70824 38558 70870 38604
rect 70928 38558 70974 38604
rect 19590 38442 19636 38488
rect 70824 38454 70870 38500
rect 70928 38454 70974 38500
rect 19722 38310 19768 38356
rect 70824 38350 70870 38396
rect 70928 38350 70974 38396
rect 70824 38246 70870 38292
rect 70928 38246 70974 38292
rect 19854 38178 19900 38224
rect 70824 38142 70870 38188
rect 70928 38142 70974 38188
rect 19986 38046 20032 38092
rect 70824 38038 70870 38084
rect 70928 38038 70974 38084
rect 20118 37914 20164 37960
rect 70824 37934 70870 37980
rect 70928 37934 70974 37980
rect 20250 37782 20296 37828
rect 70824 37830 70870 37876
rect 70928 37830 70974 37876
rect 70824 37726 70870 37772
rect 70928 37726 70974 37772
rect 20382 37650 20428 37696
rect 70824 37622 70870 37668
rect 70928 37622 70974 37668
rect 20514 37518 20560 37564
rect 70824 37518 70870 37564
rect 70928 37518 70974 37564
rect 20646 37386 20692 37432
rect 70824 37414 70870 37460
rect 70928 37414 70974 37460
rect 70824 37310 70870 37356
rect 70928 37310 70974 37356
rect 20778 37254 20824 37300
rect 70824 37206 70870 37252
rect 70928 37206 70974 37252
rect 20910 37122 20956 37168
rect 70824 37102 70870 37148
rect 70928 37102 70974 37148
rect 21042 36990 21088 37036
rect 70824 36998 70870 37044
rect 70928 36998 70974 37044
rect 21174 36858 21220 36904
rect 70824 36894 70870 36940
rect 70928 36894 70974 36940
rect 70824 36790 70870 36836
rect 70928 36790 70974 36836
rect 21306 36726 21352 36772
rect 70824 36686 70870 36732
rect 70928 36686 70974 36732
rect 21438 36594 21484 36640
rect 70824 36582 70870 36628
rect 70928 36582 70974 36628
rect 21570 36462 21616 36508
rect 70824 36478 70870 36524
rect 70928 36478 70974 36524
rect 21702 36330 21748 36376
rect 70824 36374 70870 36420
rect 70928 36374 70974 36420
rect 70824 36270 70870 36316
rect 70928 36270 70974 36316
rect 21834 36198 21880 36244
rect 70824 36166 70870 36212
rect 70928 36166 70974 36212
rect 21966 36066 22012 36112
rect 70824 36062 70870 36108
rect 70928 36062 70974 36108
rect 22098 35934 22144 35980
rect 70824 35958 70870 36004
rect 70928 35958 70974 36004
rect 22230 35802 22276 35848
rect 70824 35854 70870 35900
rect 70928 35854 70974 35900
rect 70824 35750 70870 35796
rect 70928 35750 70974 35796
rect 22362 35670 22408 35716
rect 70824 35646 70870 35692
rect 70928 35646 70974 35692
rect 22494 35538 22540 35584
rect 70824 35542 70870 35588
rect 70928 35542 70974 35588
rect 22626 35406 22672 35452
rect 70824 35438 70870 35484
rect 70928 35438 70974 35484
rect 70824 35334 70870 35380
rect 70928 35334 70974 35380
rect 22758 35274 22804 35320
rect 70824 35230 70870 35276
rect 70928 35230 70974 35276
rect 22890 35142 22936 35188
rect 70824 35126 70870 35172
rect 70928 35126 70974 35172
rect 23022 35010 23068 35056
rect 70824 35022 70870 35068
rect 70928 35022 70974 35068
rect 23154 34878 23200 34924
rect 70824 34918 70870 34964
rect 70928 34918 70974 34964
rect 70824 34814 70870 34860
rect 70928 34814 70974 34860
rect 23286 34746 23332 34792
rect 70824 34710 70870 34756
rect 70928 34710 70974 34756
rect 23418 34614 23464 34660
rect 70824 34606 70870 34652
rect 70928 34606 70974 34652
rect 23550 34482 23596 34528
rect 70824 34502 70870 34548
rect 70928 34502 70974 34548
rect 23682 34350 23728 34396
rect 70824 34398 70870 34444
rect 70928 34398 70974 34444
rect 70824 34294 70870 34340
rect 70928 34294 70974 34340
rect 23814 34218 23860 34264
rect 70824 34190 70870 34236
rect 70928 34190 70974 34236
rect 23946 34086 23992 34132
rect 70824 34086 70870 34132
rect 70928 34086 70974 34132
rect 24078 33954 24124 34000
rect 70824 33982 70870 34028
rect 70928 33982 70974 34028
rect 70824 33878 70870 33924
rect 70928 33878 70974 33924
rect 24210 33822 24256 33868
rect 70824 33774 70870 33820
rect 70928 33774 70974 33820
rect 24342 33690 24388 33736
rect 70824 33670 70870 33716
rect 70928 33670 70974 33716
rect 24474 33558 24520 33604
rect 70824 33566 70870 33612
rect 70928 33566 70974 33612
rect 24606 33426 24652 33472
rect 70824 33462 70870 33508
rect 70928 33462 70974 33508
rect 70824 33358 70870 33404
rect 70928 33358 70974 33404
rect 24738 33294 24784 33340
rect 70824 33254 70870 33300
rect 70928 33254 70974 33300
rect 24870 33162 24916 33208
rect 70824 33150 70870 33196
rect 70928 33150 70974 33196
rect 25002 33030 25048 33076
rect 70824 33046 70870 33092
rect 70928 33046 70974 33092
rect 25134 32898 25180 32944
rect 70824 32942 70870 32988
rect 70928 32942 70974 32988
rect 70824 32838 70870 32884
rect 70928 32838 70974 32884
rect 25266 32766 25312 32812
rect 70824 32734 70870 32780
rect 70928 32734 70974 32780
rect 25398 32634 25444 32680
rect 70824 32630 70870 32676
rect 70928 32630 70974 32676
rect 25530 32502 25576 32548
rect 70824 32526 70870 32572
rect 70928 32526 70974 32572
rect 25662 32370 25708 32416
rect 70824 32422 70870 32468
rect 70928 32422 70974 32468
rect 70824 32318 70870 32364
rect 70928 32318 70974 32364
rect 25794 32238 25840 32284
rect 70824 32214 70870 32260
rect 70928 32214 70974 32260
rect 25926 32106 25972 32152
rect 70824 32110 70870 32156
rect 70928 32110 70974 32156
rect 26058 31974 26104 32020
rect 70824 32006 70870 32052
rect 70928 32006 70974 32052
rect 26190 31842 26236 31888
rect 70824 31902 70870 31948
rect 70928 31902 70974 31948
rect 70824 31798 70870 31844
rect 70928 31798 70974 31844
rect 26322 31710 26368 31756
rect 70824 31694 70870 31740
rect 70928 31694 70974 31740
rect 26454 31578 26500 31624
rect 70824 31590 70870 31636
rect 70928 31590 70974 31636
rect 26586 31446 26632 31492
rect 70824 31486 70870 31532
rect 70928 31486 70974 31532
rect 70824 31382 70870 31428
rect 70928 31382 70974 31428
rect 26718 31314 26764 31360
rect 70824 31278 70870 31324
rect 70928 31278 70974 31324
rect 26850 31182 26896 31228
rect 70824 31174 70870 31220
rect 70928 31174 70974 31220
rect 26982 31050 27028 31096
rect 70824 31070 70870 31116
rect 70928 31070 70974 31116
rect 27114 30918 27160 30964
rect 70824 30966 70870 31012
rect 70928 30966 70974 31012
rect 70824 30862 70870 30908
rect 70928 30862 70974 30908
rect 27246 30786 27292 30832
rect 70824 30758 70870 30804
rect 70928 30758 70974 30804
rect 27378 30654 27424 30700
rect 70824 30654 70870 30700
rect 70928 30654 70974 30700
rect 27510 30522 27556 30568
rect 70824 30550 70870 30596
rect 70928 30550 70974 30596
rect 27642 30390 27688 30436
rect 70824 30446 70870 30492
rect 70928 30446 70974 30492
rect 70824 30342 70870 30388
rect 70928 30342 70974 30388
rect 27774 30258 27820 30304
rect 70824 30238 70870 30284
rect 70928 30238 70974 30284
rect 27906 30126 27952 30172
rect 70824 30134 70870 30180
rect 70928 30134 70974 30180
rect 28038 29994 28084 30040
rect 70824 30030 70870 30076
rect 70928 30030 70974 30076
rect 70824 29926 70870 29972
rect 70928 29926 70974 29972
rect 28170 29862 28216 29908
rect 70824 29822 70870 29868
rect 70928 29822 70974 29868
rect 28302 29730 28348 29776
rect 70824 29718 70870 29764
rect 70928 29718 70974 29764
rect 28434 29598 28480 29644
rect 70824 29614 70870 29660
rect 70928 29614 70974 29660
rect 28566 29466 28612 29512
rect 70824 29510 70870 29556
rect 70928 29510 70974 29556
rect 70824 29406 70870 29452
rect 70928 29406 70974 29452
rect 28698 29334 28744 29380
rect 70824 29302 70870 29348
rect 70928 29302 70974 29348
rect 28830 29202 28876 29248
rect 70824 29198 70870 29244
rect 70928 29198 70974 29244
rect 28962 29070 29008 29116
rect 70824 29094 70870 29140
rect 70928 29094 70974 29140
rect 29094 28938 29140 28984
rect 70824 28990 70870 29036
rect 70928 28990 70974 29036
rect 70824 28886 70870 28932
rect 70928 28886 70974 28932
rect 29226 28806 29272 28852
rect 70824 28782 70870 28828
rect 70928 28782 70974 28828
rect 29358 28674 29404 28720
rect 70824 28678 70870 28724
rect 70928 28678 70974 28724
rect 29490 28542 29536 28588
rect 70824 28574 70870 28620
rect 70928 28574 70974 28620
rect 70824 28470 70870 28516
rect 70928 28470 70974 28516
rect 29622 28410 29668 28456
rect 70824 28366 70870 28412
rect 70928 28366 70974 28412
rect 29754 28278 29800 28324
rect 70824 28262 70870 28308
rect 70928 28262 70974 28308
rect 29886 28146 29932 28192
rect 70824 28158 70870 28204
rect 70928 28158 70974 28204
rect 30018 28014 30064 28060
rect 70824 28054 70870 28100
rect 70928 28054 70974 28100
rect 70824 27950 70870 27996
rect 70928 27950 70974 27996
rect 30150 27882 30196 27928
rect 70824 27846 70870 27892
rect 70928 27846 70974 27892
rect 30282 27750 30328 27796
rect 70824 27742 70870 27788
rect 70928 27742 70974 27788
rect 30414 27618 30460 27664
rect 70824 27638 70870 27684
rect 70928 27638 70974 27684
rect 30546 27486 30592 27532
rect 70824 27534 70870 27580
rect 70928 27534 70974 27580
rect 70824 27430 70870 27476
rect 70928 27430 70974 27476
rect 30678 27354 30724 27400
rect 70824 27326 70870 27372
rect 70928 27326 70974 27372
rect 30810 27222 30856 27268
rect 70824 27222 70870 27268
rect 70928 27222 70974 27268
rect 30942 27090 30988 27136
rect 70824 27118 70870 27164
rect 70928 27118 70974 27164
rect 70824 27014 70870 27060
rect 70928 27014 70974 27060
rect 31074 26958 31120 27004
rect 70824 26910 70870 26956
rect 70928 26910 70974 26956
rect 31206 26826 31252 26872
rect 70824 26806 70870 26852
rect 70928 26806 70974 26852
rect 31338 26694 31384 26740
rect 70824 26702 70870 26748
rect 70928 26702 70974 26748
rect 31470 26562 31516 26608
rect 70824 26598 70870 26644
rect 70928 26598 70974 26644
rect 70824 26494 70870 26540
rect 70928 26494 70974 26540
rect 31602 26430 31648 26476
rect 70824 26390 70870 26436
rect 70928 26390 70974 26436
rect 31734 26298 31780 26344
rect 70824 26286 70870 26332
rect 70928 26286 70974 26332
rect 31866 26166 31912 26212
rect 70824 26182 70870 26228
rect 70928 26182 70974 26228
rect 31998 26034 32044 26080
rect 70824 26078 70870 26124
rect 70928 26078 70974 26124
rect 70824 25974 70870 26020
rect 70928 25974 70974 26020
rect 32130 25902 32176 25948
rect 70824 25870 70870 25916
rect 70928 25870 70974 25916
rect 32262 25770 32308 25816
rect 70824 25766 70870 25812
rect 70928 25766 70974 25812
rect 32394 25638 32440 25684
rect 70824 25662 70870 25708
rect 70928 25662 70974 25708
rect 32526 25506 32572 25552
rect 70824 25558 70870 25604
rect 70928 25558 70974 25604
rect 70824 25454 70870 25500
rect 70928 25454 70974 25500
rect 32658 25374 32704 25420
rect 70824 25350 70870 25396
rect 70928 25350 70974 25396
rect 32790 25242 32836 25288
rect 70824 25246 70870 25292
rect 70928 25246 70974 25292
rect 32922 25110 32968 25156
rect 70824 25142 70870 25188
rect 70928 25142 70974 25188
rect 70824 25038 70870 25084
rect 70928 25038 70974 25084
rect 33054 24978 33100 25024
rect 70824 24934 70870 24980
rect 70928 24934 70974 24980
rect 33186 24846 33232 24892
rect 70824 24830 70870 24876
rect 70928 24830 70974 24876
rect 33318 24714 33364 24760
rect 70824 24726 70870 24772
rect 70928 24726 70974 24772
rect 33450 24582 33496 24628
rect 70824 24622 70870 24668
rect 70928 24622 70974 24668
rect 70824 24518 70870 24564
rect 70928 24518 70974 24564
rect 33582 24450 33628 24496
rect 70824 24414 70870 24460
rect 70928 24414 70974 24460
rect 33714 24318 33760 24364
rect 70824 24310 70870 24356
rect 70928 24310 70974 24356
rect 33846 24186 33892 24232
rect 70824 24206 70870 24252
rect 70928 24206 70974 24252
rect 33978 24054 34024 24100
rect 70824 24102 70870 24148
rect 70928 24102 70974 24148
rect 70824 23998 70870 24044
rect 70928 23998 70974 24044
rect 34110 23922 34156 23968
rect 70824 23894 70870 23940
rect 70928 23894 70974 23940
rect 34242 23790 34288 23836
rect 70824 23790 70870 23836
rect 70928 23790 70974 23836
rect 34374 23658 34420 23704
rect 70824 23686 70870 23732
rect 70928 23686 70974 23732
rect 70824 23582 70870 23628
rect 70928 23582 70974 23628
rect 34506 23526 34552 23572
rect 70824 23478 70870 23524
rect 70928 23478 70974 23524
rect 34638 23394 34684 23440
rect 70824 23374 70870 23420
rect 70928 23374 70974 23420
rect 34770 23262 34816 23308
rect 70824 23270 70870 23316
rect 70928 23270 70974 23316
rect 34902 23130 34948 23176
rect 70824 23166 70870 23212
rect 70928 23166 70974 23212
rect 70824 23062 70870 23108
rect 70928 23062 70974 23108
rect 35034 22998 35080 23044
rect 70824 22958 70870 23004
rect 70928 22958 70974 23004
rect 35166 22866 35212 22912
rect 70824 22854 70870 22900
rect 70928 22854 70974 22900
rect 35298 22734 35344 22780
rect 70824 22750 70870 22796
rect 70928 22750 70974 22796
rect 35430 22602 35476 22648
rect 70824 22646 70870 22692
rect 70928 22646 70974 22692
rect 70824 22542 70870 22588
rect 70928 22542 70974 22588
rect 35562 22470 35608 22516
rect 70824 22438 70870 22484
rect 70928 22438 70974 22484
rect 35694 22338 35740 22384
rect 70824 22334 70870 22380
rect 70928 22334 70974 22380
rect 35826 22206 35872 22252
rect 70824 22230 70870 22276
rect 70928 22230 70974 22276
rect 70824 22126 70870 22172
rect 70928 22126 70974 22172
rect 35958 22074 36004 22120
rect 70824 22022 70870 22068
rect 70928 22022 70974 22068
rect 36090 21942 36136 21988
rect 70824 21918 70870 21964
rect 70928 21918 70974 21964
rect 36222 21810 36268 21856
rect 70824 21814 70870 21860
rect 70928 21814 70974 21860
rect 36354 21678 36400 21724
rect 70824 21710 70870 21756
rect 70928 21710 70974 21756
rect 70824 21606 70870 21652
rect 70928 21606 70974 21652
rect 36486 21546 36532 21592
rect 70824 21502 70870 21548
rect 70928 21502 70974 21548
rect 36618 21414 36664 21460
rect 70824 21398 70870 21444
rect 70928 21398 70974 21444
rect 36750 21282 36796 21328
rect 70824 21294 70870 21340
rect 70928 21294 70974 21340
rect 36882 21150 36928 21196
rect 70824 21190 70870 21236
rect 70928 21190 70974 21236
rect 70824 21086 70870 21132
rect 70928 21086 70974 21132
rect 37014 21018 37060 21064
rect 70824 20982 70870 21028
rect 70928 20982 70974 21028
rect 37146 20886 37192 20932
rect 70824 20878 70870 20924
rect 70928 20878 70974 20924
rect 37278 20754 37324 20800
rect 70824 20774 70870 20820
rect 70928 20774 70974 20820
rect 37410 20622 37456 20668
rect 70824 20670 70870 20716
rect 70928 20670 70974 20716
rect 70824 20566 70870 20612
rect 70928 20566 70974 20612
rect 37542 20490 37588 20536
rect 70824 20462 70870 20508
rect 70928 20462 70974 20508
rect 37674 20358 37720 20404
rect 70824 20358 70870 20404
rect 70928 20358 70974 20404
rect 37806 20226 37852 20272
rect 70824 20254 70870 20300
rect 70928 20254 70974 20300
rect 70824 20150 70870 20196
rect 70928 20150 70974 20196
rect 37938 20094 37984 20140
rect 70824 20046 70870 20092
rect 70928 20046 70974 20092
rect 38070 19962 38116 20008
rect 70824 19942 70870 19988
rect 70928 19942 70974 19988
rect 38202 19830 38248 19876
rect 70824 19838 70870 19884
rect 70928 19838 70974 19884
rect 38334 19698 38380 19744
rect 70824 19734 70870 19780
rect 70928 19734 70974 19780
rect 70824 19630 70870 19676
rect 70928 19630 70974 19676
rect 38466 19566 38512 19612
rect 70824 19526 70870 19572
rect 70928 19526 70974 19572
rect 38598 19434 38644 19480
rect 70824 19422 70870 19468
rect 70928 19422 70974 19468
rect 38730 19302 38776 19348
rect 70824 19318 70870 19364
rect 70928 19318 70974 19364
rect 38862 19170 38908 19216
rect 70824 19214 70870 19260
rect 70928 19214 70974 19260
rect 70824 19110 70870 19156
rect 70928 19110 70974 19156
rect 38994 19038 39040 19084
rect 70824 19006 70870 19052
rect 70928 19006 70974 19052
rect 39126 18906 39172 18952
rect 70824 18902 70870 18948
rect 70928 18902 70974 18948
rect 39258 18774 39304 18820
rect 70824 18798 70870 18844
rect 70928 18798 70974 18844
rect 39390 18642 39436 18688
rect 70824 18694 70870 18740
rect 70928 18694 70974 18740
rect 70824 18590 70870 18636
rect 70928 18590 70974 18636
rect 39522 18510 39568 18556
rect 70824 18486 70870 18532
rect 70928 18486 70974 18532
rect 39654 18378 39700 18424
rect 70824 18382 70870 18428
rect 70928 18382 70974 18428
rect 39786 18246 39832 18292
rect 70824 18278 70870 18324
rect 70928 18278 70974 18324
rect 70824 18174 70870 18220
rect 70928 18174 70974 18220
rect 39918 18114 39964 18160
rect 70824 18070 70870 18116
rect 70928 18070 70974 18116
rect 40050 17982 40096 18028
rect 70824 17966 70870 18012
rect 70928 17966 70974 18012
rect 40182 17850 40228 17896
rect 70824 17862 70870 17908
rect 70928 17862 70974 17908
rect 40314 17718 40360 17764
rect 70824 17758 70870 17804
rect 70928 17758 70974 17804
rect 70824 17654 70870 17700
rect 70928 17654 70974 17700
rect 40446 17586 40492 17632
rect 70824 17550 70870 17596
rect 70928 17550 70974 17596
rect 40578 17454 40624 17500
rect 70824 17446 70870 17492
rect 70928 17446 70974 17492
rect 40710 17322 40756 17368
rect 70824 17342 70870 17388
rect 70928 17342 70974 17388
rect 40842 17190 40888 17236
rect 70824 17238 70870 17284
rect 70928 17238 70974 17284
rect 70824 17134 70870 17180
rect 70928 17134 70974 17180
rect 40974 17058 41020 17104
rect 70824 17030 70870 17076
rect 70928 17030 70974 17076
rect 41106 16926 41152 16972
rect 70824 16926 70870 16972
rect 70928 16926 70974 16972
rect 41238 16794 41284 16840
rect 70824 16822 70870 16868
rect 70928 16822 70974 16868
rect 70824 16718 70870 16764
rect 70928 16718 70974 16764
rect 41370 16662 41416 16708
rect 70824 16614 70870 16660
rect 70928 16614 70974 16660
rect 41502 16530 41548 16576
rect 70824 16510 70870 16556
rect 70928 16510 70974 16556
rect 41634 16398 41680 16444
rect 70824 16406 70870 16452
rect 70928 16406 70974 16452
rect 41766 16266 41812 16312
rect 70824 16302 70870 16348
rect 70928 16302 70974 16348
rect 70824 16198 70870 16244
rect 70928 16198 70974 16244
rect 41898 16134 41944 16180
rect 70824 16094 70870 16140
rect 70928 16094 70974 16140
rect 42030 16002 42076 16048
rect 70824 15990 70870 16036
rect 70928 15990 70974 16036
rect 42162 15870 42208 15916
rect 70824 15886 70870 15932
rect 70928 15886 70974 15932
rect 42294 15738 42340 15784
rect 70824 15782 70870 15828
rect 70928 15782 70974 15828
rect 70824 15678 70870 15724
rect 70928 15678 70974 15724
rect 42426 15606 42472 15652
rect 70824 15574 70870 15620
rect 70928 15574 70974 15620
rect 42558 15474 42604 15520
rect 70824 15470 70870 15516
rect 70928 15470 70974 15516
rect 42690 15342 42736 15388
rect 70824 15366 70870 15412
rect 70928 15366 70974 15412
rect 70824 15262 70870 15308
rect 70928 15262 70974 15308
rect 42822 15210 42868 15256
rect 70824 15158 70870 15204
rect 70928 15158 70974 15204
rect 42954 15078 43000 15124
rect 70824 15054 70870 15100
rect 70928 15054 70974 15100
rect 43086 14946 43132 14992
rect 70824 14950 70870 14996
rect 70928 14950 70974 14996
rect 43218 14814 43264 14860
rect 70824 14846 70870 14892
rect 70928 14846 70974 14892
rect 70824 14742 70870 14788
rect 70928 14742 70974 14788
rect 43350 14682 43396 14728
rect 70824 14638 70870 14684
rect 70928 14638 70974 14684
rect 43482 14550 43528 14596
rect 70824 14534 70870 14580
rect 70928 14534 70974 14580
rect 43614 14418 43660 14464
rect 70824 14430 70870 14476
rect 70928 14430 70974 14476
rect 43746 14286 43792 14332
rect 70824 14326 70870 14372
rect 70928 14326 70974 14372
rect 70824 14222 70870 14268
rect 70928 14222 70974 14268
rect 43878 14154 43924 14200
rect 70824 14118 70870 14164
rect 70928 14118 70974 14164
rect 44010 14022 44056 14068
rect 70824 14014 70870 14060
rect 70928 14014 70974 14060
rect 44142 13890 44188 13936
rect 70824 13910 70870 13956
rect 70928 13910 70974 13956
rect 44274 13758 44320 13804
rect 70824 13806 70870 13852
rect 70928 13806 70974 13852
rect 70824 13702 70870 13748
rect 70928 13702 70974 13748
rect 44406 13626 44452 13672
rect 70824 13598 70870 13644
rect 70928 13598 70974 13644
rect 44538 13494 44584 13540
rect 70824 13494 70870 13540
rect 70928 13494 70974 13540
rect 44670 13362 44716 13408
rect 70824 13390 70870 13436
rect 70928 13390 70974 13436
rect 44850 13210 44896 13256
rect 45088 13223 45134 13269
rect 45192 13223 45238 13269
rect 45296 13223 45342 13269
rect 45400 13223 45446 13269
rect 45504 13223 45550 13269
rect 45608 13223 45654 13269
rect 45712 13223 45758 13269
rect 45816 13223 45862 13269
rect 45920 13223 45966 13269
rect 46024 13223 46070 13269
rect 46128 13223 46174 13269
rect 46232 13223 46278 13269
rect 46336 13223 46382 13269
rect 46440 13223 46486 13269
rect 46544 13223 46590 13269
rect 46648 13223 46694 13269
rect 46752 13223 46798 13269
rect 46856 13223 46902 13269
rect 46960 13223 47006 13269
rect 47064 13223 47110 13269
rect 47168 13223 47214 13269
rect 47272 13223 47318 13269
rect 47376 13223 47422 13269
rect 47480 13223 47526 13269
rect 47584 13223 47630 13269
rect 47688 13223 47734 13269
rect 47792 13223 47838 13269
rect 47896 13223 47942 13269
rect 48000 13223 48046 13269
rect 48104 13223 48150 13269
rect 48208 13223 48254 13269
rect 48312 13223 48358 13269
rect 48416 13223 48462 13269
rect 48520 13223 48566 13269
rect 48624 13223 48670 13269
rect 48728 13223 48774 13269
rect 48832 13223 48878 13269
rect 48936 13223 48982 13269
rect 49040 13223 49086 13269
rect 49144 13223 49190 13269
rect 49248 13223 49294 13269
rect 49352 13223 49398 13269
rect 49456 13223 49502 13269
rect 49560 13223 49606 13269
rect 49664 13223 49710 13269
rect 49768 13223 49814 13269
rect 49872 13223 49918 13269
rect 49976 13223 50022 13269
rect 50080 13223 50126 13269
rect 50184 13223 50230 13269
rect 50288 13223 50334 13269
rect 50392 13223 50438 13269
rect 50496 13223 50542 13269
rect 50600 13223 50646 13269
rect 50704 13223 50750 13269
rect 50808 13223 50854 13269
rect 50912 13223 50958 13269
rect 51016 13223 51062 13269
rect 51120 13223 51166 13269
rect 51224 13223 51270 13269
rect 51328 13223 51374 13269
rect 51432 13223 51478 13269
rect 51536 13223 51582 13269
rect 51640 13223 51686 13269
rect 51744 13223 51790 13269
rect 51848 13223 51894 13269
rect 51952 13223 51998 13269
rect 52056 13223 52102 13269
rect 52160 13223 52206 13269
rect 52264 13223 52310 13269
rect 52368 13223 52414 13269
rect 52472 13223 52518 13269
rect 52576 13223 52622 13269
rect 52680 13223 52726 13269
rect 52784 13223 52830 13269
rect 52888 13223 52934 13269
rect 52992 13223 53038 13269
rect 53096 13223 53142 13269
rect 53200 13223 53246 13269
rect 53304 13223 53350 13269
rect 53408 13223 53454 13269
rect 53512 13223 53558 13269
rect 53616 13223 53662 13269
rect 53720 13223 53766 13269
rect 53824 13223 53870 13269
rect 53928 13223 53974 13269
rect 54032 13223 54078 13269
rect 54136 13223 54182 13269
rect 54240 13223 54286 13269
rect 54344 13223 54390 13269
rect 54448 13223 54494 13269
rect 54552 13223 54598 13269
rect 54656 13223 54702 13269
rect 54760 13223 54806 13269
rect 54864 13223 54910 13269
rect 54968 13223 55014 13269
rect 55072 13223 55118 13269
rect 55176 13223 55222 13269
rect 55280 13223 55326 13269
rect 55384 13223 55430 13269
rect 55488 13223 55534 13269
rect 55592 13223 55638 13269
rect 55696 13223 55742 13269
rect 55800 13223 55846 13269
rect 55904 13223 55950 13269
rect 56008 13223 56054 13269
rect 56112 13223 56158 13269
rect 56216 13223 56262 13269
rect 56320 13223 56366 13269
rect 56424 13223 56470 13269
rect 56528 13223 56574 13269
rect 56632 13223 56678 13269
rect 56736 13223 56782 13269
rect 56840 13223 56886 13269
rect 56944 13223 56990 13269
rect 57048 13223 57094 13269
rect 57152 13223 57198 13269
rect 57256 13223 57302 13269
rect 57360 13223 57406 13269
rect 57464 13223 57510 13269
rect 57568 13223 57614 13269
rect 57672 13223 57718 13269
rect 57776 13223 57822 13269
rect 57880 13223 57926 13269
rect 57984 13223 58030 13269
rect 58088 13223 58134 13269
rect 58192 13223 58238 13269
rect 58296 13223 58342 13269
rect 58400 13223 58446 13269
rect 58504 13223 58550 13269
rect 58608 13223 58654 13269
rect 58712 13223 58758 13269
rect 58816 13223 58862 13269
rect 58920 13223 58966 13269
rect 59024 13223 59070 13269
rect 59128 13223 59174 13269
rect 59232 13223 59278 13269
rect 59336 13223 59382 13269
rect 59440 13223 59486 13269
rect 59544 13223 59590 13269
rect 59648 13223 59694 13269
rect 59752 13223 59798 13269
rect 59856 13223 59902 13269
rect 59960 13223 60006 13269
rect 60064 13223 60110 13269
rect 60168 13223 60214 13269
rect 60272 13223 60318 13269
rect 60376 13223 60422 13269
rect 60480 13223 60526 13269
rect 60584 13223 60630 13269
rect 60688 13223 60734 13269
rect 60792 13223 60838 13269
rect 60896 13223 60942 13269
rect 61000 13223 61046 13269
rect 61104 13223 61150 13269
rect 61208 13223 61254 13269
rect 61312 13223 61358 13269
rect 61416 13223 61462 13269
rect 61520 13223 61566 13269
rect 61624 13223 61670 13269
rect 61728 13223 61774 13269
rect 61832 13223 61878 13269
rect 61936 13223 61982 13269
rect 62040 13223 62086 13269
rect 62144 13223 62190 13269
rect 62248 13223 62294 13269
rect 62352 13223 62398 13269
rect 62456 13223 62502 13269
rect 62560 13223 62606 13269
rect 62664 13223 62710 13269
rect 62768 13223 62814 13269
rect 62872 13223 62918 13269
rect 62976 13223 63022 13269
rect 63080 13223 63126 13269
rect 63184 13223 63230 13269
rect 63288 13223 63334 13269
rect 63392 13223 63438 13269
rect 63496 13223 63542 13269
rect 63600 13223 63646 13269
rect 63704 13223 63750 13269
rect 63808 13223 63854 13269
rect 63912 13223 63958 13269
rect 64016 13223 64062 13269
rect 64120 13223 64166 13269
rect 64224 13223 64270 13269
rect 64328 13223 64374 13269
rect 64432 13223 64478 13269
rect 64536 13223 64582 13269
rect 64640 13223 64686 13269
rect 64744 13223 64790 13269
rect 64848 13223 64894 13269
rect 64952 13223 64998 13269
rect 65056 13223 65102 13269
rect 65160 13223 65206 13269
rect 65264 13223 65310 13269
rect 65368 13223 65414 13269
rect 65472 13223 65518 13269
rect 65576 13223 65622 13269
rect 65680 13223 65726 13269
rect 65784 13223 65830 13269
rect 65888 13223 65934 13269
rect 65992 13223 66038 13269
rect 66096 13223 66142 13269
rect 66200 13223 66246 13269
rect 66304 13223 66350 13269
rect 66408 13223 66454 13269
rect 66512 13223 66558 13269
rect 66616 13223 66662 13269
rect 66720 13223 66766 13269
rect 66824 13223 66870 13269
rect 66928 13223 66974 13269
rect 67032 13223 67078 13269
rect 67136 13223 67182 13269
rect 67240 13223 67286 13269
rect 67344 13223 67390 13269
rect 67448 13223 67494 13269
rect 67552 13223 67598 13269
rect 67656 13223 67702 13269
rect 67760 13223 67806 13269
rect 67864 13223 67910 13269
rect 67968 13223 68014 13269
rect 68072 13223 68118 13269
rect 68176 13223 68222 13269
rect 68280 13223 68326 13269
rect 68384 13223 68430 13269
rect 68488 13223 68534 13269
rect 68592 13223 68638 13269
rect 68696 13223 68742 13269
rect 68800 13223 68846 13269
rect 68904 13223 68950 13269
rect 69008 13223 69054 13269
rect 69112 13223 69158 13269
rect 69216 13223 69262 13269
rect 69320 13223 69366 13269
rect 69424 13223 69470 13269
rect 69528 13223 69574 13269
rect 69632 13223 69678 13269
rect 69736 13223 69782 13269
rect 69840 13223 69886 13269
rect 69944 13223 69990 13269
rect 70048 13223 70094 13269
rect 70152 13223 70198 13269
rect 70256 13223 70302 13269
rect 70360 13223 70406 13269
rect 70464 13223 70510 13269
rect 70568 13223 70614 13269
rect 70672 13223 70718 13269
rect 70776 13223 70822 13269
rect 70880 13223 70926 13269
rect 45088 13119 45134 13165
rect 45192 13119 45238 13165
rect 45296 13119 45342 13165
rect 45400 13119 45446 13165
rect 45504 13119 45550 13165
rect 45608 13119 45654 13165
rect 45712 13119 45758 13165
rect 45816 13119 45862 13165
rect 45920 13119 45966 13165
rect 46024 13119 46070 13165
rect 46128 13119 46174 13165
rect 46232 13119 46278 13165
rect 46336 13119 46382 13165
rect 46440 13119 46486 13165
rect 46544 13119 46590 13165
rect 46648 13119 46694 13165
rect 46752 13119 46798 13165
rect 46856 13119 46902 13165
rect 46960 13119 47006 13165
rect 47064 13119 47110 13165
rect 47168 13119 47214 13165
rect 47272 13119 47318 13165
rect 47376 13119 47422 13165
rect 47480 13119 47526 13165
rect 47584 13119 47630 13165
rect 47688 13119 47734 13165
rect 47792 13119 47838 13165
rect 47896 13119 47942 13165
rect 48000 13119 48046 13165
rect 48104 13119 48150 13165
rect 48208 13119 48254 13165
rect 48312 13119 48358 13165
rect 48416 13119 48462 13165
rect 48520 13119 48566 13165
rect 48624 13119 48670 13165
rect 48728 13119 48774 13165
rect 48832 13119 48878 13165
rect 48936 13119 48982 13165
rect 49040 13119 49086 13165
rect 49144 13119 49190 13165
rect 49248 13119 49294 13165
rect 49352 13119 49398 13165
rect 49456 13119 49502 13165
rect 49560 13119 49606 13165
rect 49664 13119 49710 13165
rect 49768 13119 49814 13165
rect 49872 13119 49918 13165
rect 49976 13119 50022 13165
rect 50080 13119 50126 13165
rect 50184 13119 50230 13165
rect 50288 13119 50334 13165
rect 50392 13119 50438 13165
rect 50496 13119 50542 13165
rect 50600 13119 50646 13165
rect 50704 13119 50750 13165
rect 50808 13119 50854 13165
rect 50912 13119 50958 13165
rect 51016 13119 51062 13165
rect 51120 13119 51166 13165
rect 51224 13119 51270 13165
rect 51328 13119 51374 13165
rect 51432 13119 51478 13165
rect 51536 13119 51582 13165
rect 51640 13119 51686 13165
rect 51744 13119 51790 13165
rect 51848 13119 51894 13165
rect 51952 13119 51998 13165
rect 52056 13119 52102 13165
rect 52160 13119 52206 13165
rect 52264 13119 52310 13165
rect 52368 13119 52414 13165
rect 52472 13119 52518 13165
rect 52576 13119 52622 13165
rect 52680 13119 52726 13165
rect 52784 13119 52830 13165
rect 52888 13119 52934 13165
rect 52992 13119 53038 13165
rect 53096 13119 53142 13165
rect 53200 13119 53246 13165
rect 53304 13119 53350 13165
rect 53408 13119 53454 13165
rect 53512 13119 53558 13165
rect 53616 13119 53662 13165
rect 53720 13119 53766 13165
rect 53824 13119 53870 13165
rect 53928 13119 53974 13165
rect 54032 13119 54078 13165
rect 54136 13119 54182 13165
rect 54240 13119 54286 13165
rect 54344 13119 54390 13165
rect 54448 13119 54494 13165
rect 54552 13119 54598 13165
rect 54656 13119 54702 13165
rect 54760 13119 54806 13165
rect 54864 13119 54910 13165
rect 54968 13119 55014 13165
rect 55072 13119 55118 13165
rect 55176 13119 55222 13165
rect 55280 13119 55326 13165
rect 55384 13119 55430 13165
rect 55488 13119 55534 13165
rect 55592 13119 55638 13165
rect 55696 13119 55742 13165
rect 55800 13119 55846 13165
rect 55904 13119 55950 13165
rect 56008 13119 56054 13165
rect 56112 13119 56158 13165
rect 56216 13119 56262 13165
rect 56320 13119 56366 13165
rect 56424 13119 56470 13165
rect 56528 13119 56574 13165
rect 56632 13119 56678 13165
rect 56736 13119 56782 13165
rect 56840 13119 56886 13165
rect 56944 13119 56990 13165
rect 57048 13119 57094 13165
rect 57152 13119 57198 13165
rect 57256 13119 57302 13165
rect 57360 13119 57406 13165
rect 57464 13119 57510 13165
rect 57568 13119 57614 13165
rect 57672 13119 57718 13165
rect 57776 13119 57822 13165
rect 57880 13119 57926 13165
rect 57984 13119 58030 13165
rect 58088 13119 58134 13165
rect 58192 13119 58238 13165
rect 58296 13119 58342 13165
rect 58400 13119 58446 13165
rect 58504 13119 58550 13165
rect 58608 13119 58654 13165
rect 58712 13119 58758 13165
rect 58816 13119 58862 13165
rect 58920 13119 58966 13165
rect 59024 13119 59070 13165
rect 59128 13119 59174 13165
rect 59232 13119 59278 13165
rect 59336 13119 59382 13165
rect 59440 13119 59486 13165
rect 59544 13119 59590 13165
rect 59648 13119 59694 13165
rect 59752 13119 59798 13165
rect 59856 13119 59902 13165
rect 59960 13119 60006 13165
rect 60064 13119 60110 13165
rect 60168 13119 60214 13165
rect 60272 13119 60318 13165
rect 60376 13119 60422 13165
rect 60480 13119 60526 13165
rect 60584 13119 60630 13165
rect 60688 13119 60734 13165
rect 60792 13119 60838 13165
rect 60896 13119 60942 13165
rect 61000 13119 61046 13165
rect 61104 13119 61150 13165
rect 61208 13119 61254 13165
rect 61312 13119 61358 13165
rect 61416 13119 61462 13165
rect 61520 13119 61566 13165
rect 61624 13119 61670 13165
rect 61728 13119 61774 13165
rect 61832 13119 61878 13165
rect 61936 13119 61982 13165
rect 62040 13119 62086 13165
rect 62144 13119 62190 13165
rect 62248 13119 62294 13165
rect 62352 13119 62398 13165
rect 62456 13119 62502 13165
rect 62560 13119 62606 13165
rect 62664 13119 62710 13165
rect 62768 13119 62814 13165
rect 62872 13119 62918 13165
rect 62976 13119 63022 13165
rect 63080 13119 63126 13165
rect 63184 13119 63230 13165
rect 63288 13119 63334 13165
rect 63392 13119 63438 13165
rect 63496 13119 63542 13165
rect 63600 13119 63646 13165
rect 63704 13119 63750 13165
rect 63808 13119 63854 13165
rect 63912 13119 63958 13165
rect 64016 13119 64062 13165
rect 64120 13119 64166 13165
rect 64224 13119 64270 13165
rect 64328 13119 64374 13165
rect 64432 13119 64478 13165
rect 64536 13119 64582 13165
rect 64640 13119 64686 13165
rect 64744 13119 64790 13165
rect 64848 13119 64894 13165
rect 64952 13119 64998 13165
rect 65056 13119 65102 13165
rect 65160 13119 65206 13165
rect 65264 13119 65310 13165
rect 65368 13119 65414 13165
rect 65472 13119 65518 13165
rect 65576 13119 65622 13165
rect 65680 13119 65726 13165
rect 65784 13119 65830 13165
rect 65888 13119 65934 13165
rect 65992 13119 66038 13165
rect 66096 13119 66142 13165
rect 66200 13119 66246 13165
rect 66304 13119 66350 13165
rect 66408 13119 66454 13165
rect 66512 13119 66558 13165
rect 66616 13119 66662 13165
rect 66720 13119 66766 13165
rect 66824 13119 66870 13165
rect 66928 13119 66974 13165
rect 67032 13119 67078 13165
rect 67136 13119 67182 13165
rect 67240 13119 67286 13165
rect 67344 13119 67390 13165
rect 67448 13119 67494 13165
rect 67552 13119 67598 13165
rect 67656 13119 67702 13165
rect 67760 13119 67806 13165
rect 67864 13119 67910 13165
rect 67968 13119 68014 13165
rect 68072 13119 68118 13165
rect 68176 13119 68222 13165
rect 68280 13119 68326 13165
rect 68384 13119 68430 13165
rect 68488 13119 68534 13165
rect 68592 13119 68638 13165
rect 68696 13119 68742 13165
rect 68800 13119 68846 13165
rect 68904 13119 68950 13165
rect 69008 13119 69054 13165
rect 69112 13119 69158 13165
rect 69216 13119 69262 13165
rect 69320 13119 69366 13165
rect 69424 13119 69470 13165
rect 69528 13119 69574 13165
rect 69632 13119 69678 13165
rect 69736 13119 69782 13165
rect 69840 13119 69886 13165
rect 69944 13119 69990 13165
rect 70048 13119 70094 13165
rect 70152 13119 70198 13165
rect 70256 13119 70302 13165
rect 70360 13119 70406 13165
rect 70464 13119 70510 13165
rect 70568 13119 70614 13165
rect 70672 13119 70718 13165
rect 70776 13119 70822 13165
rect 70880 13119 70926 13165
<< metal1 >>
rect 13108 70975 69957 71000
rect 13108 70929 13119 70975
rect 13165 70929 13223 70975
rect 13269 70929 13377 70975
rect 13423 70929 13481 70975
rect 13527 70929 13585 70975
rect 13631 70929 13689 70975
rect 13735 70929 13793 70975
rect 13839 70929 13897 70975
rect 13943 70929 14001 70975
rect 14047 70929 14105 70975
rect 14151 70929 14209 70975
rect 14255 70929 14313 70975
rect 14359 70929 14417 70975
rect 14463 70929 14521 70975
rect 14567 70929 14625 70975
rect 14671 70929 14729 70975
rect 14775 70929 14833 70975
rect 14879 70929 14937 70975
rect 14983 70929 15041 70975
rect 15087 70929 15145 70975
rect 15191 70929 15249 70975
rect 15295 70929 15353 70975
rect 15399 70929 15457 70975
rect 15503 70929 15561 70975
rect 15607 70929 15665 70975
rect 15711 70929 15769 70975
rect 15815 70929 15873 70975
rect 15919 70929 15977 70975
rect 16023 70929 16081 70975
rect 16127 70929 16185 70975
rect 16231 70929 16289 70975
rect 16335 70929 16393 70975
rect 16439 70929 16497 70975
rect 16543 70929 16601 70975
rect 16647 70929 16705 70975
rect 16751 70929 16809 70975
rect 16855 70929 16913 70975
rect 16959 70929 17017 70975
rect 17063 70929 17121 70975
rect 17167 70929 17225 70975
rect 17271 70929 17329 70975
rect 17375 70929 17433 70975
rect 17479 70929 17537 70975
rect 17583 70929 17641 70975
rect 17687 70929 17745 70975
rect 17791 70929 17849 70975
rect 17895 70929 17953 70975
rect 17999 70929 18057 70975
rect 18103 70929 18161 70975
rect 18207 70929 18265 70975
rect 18311 70929 18369 70975
rect 18415 70929 18473 70975
rect 18519 70929 18577 70975
rect 18623 70929 18681 70975
rect 18727 70929 18785 70975
rect 18831 70929 18889 70975
rect 18935 70929 18993 70975
rect 19039 70929 19097 70975
rect 19143 70929 19201 70975
rect 19247 70929 19305 70975
rect 19351 70929 19409 70975
rect 19455 70929 19513 70975
rect 19559 70929 19617 70975
rect 19663 70929 19721 70975
rect 19767 70929 19825 70975
rect 19871 70929 19929 70975
rect 19975 70929 20033 70975
rect 20079 70929 20137 70975
rect 20183 70929 20241 70975
rect 20287 70929 20345 70975
rect 20391 70929 20449 70975
rect 20495 70929 20553 70975
rect 20599 70929 20657 70975
rect 20703 70929 20761 70975
rect 20807 70929 20865 70975
rect 20911 70929 20969 70975
rect 21015 70929 21073 70975
rect 21119 70929 21177 70975
rect 21223 70929 21281 70975
rect 21327 70929 21385 70975
rect 21431 70929 21489 70975
rect 21535 70929 21593 70975
rect 21639 70929 21697 70975
rect 21743 70929 21801 70975
rect 21847 70929 21905 70975
rect 21951 70929 22009 70975
rect 22055 70929 22113 70975
rect 22159 70929 22217 70975
rect 22263 70929 22321 70975
rect 22367 70929 22425 70975
rect 22471 70929 22529 70975
rect 22575 70929 22633 70975
rect 22679 70929 22737 70975
rect 22783 70929 22841 70975
rect 22887 70929 22945 70975
rect 22991 70929 23049 70975
rect 23095 70929 23153 70975
rect 23199 70929 23257 70975
rect 23303 70929 23361 70975
rect 23407 70929 23465 70975
rect 23511 70929 23569 70975
rect 23615 70929 23673 70975
rect 23719 70929 23777 70975
rect 23823 70929 23881 70975
rect 23927 70929 23985 70975
rect 24031 70929 24089 70975
rect 24135 70929 24193 70975
rect 24239 70929 24297 70975
rect 24343 70929 24401 70975
rect 24447 70929 24505 70975
rect 24551 70929 24609 70975
rect 24655 70929 24713 70975
rect 24759 70929 24817 70975
rect 24863 70929 24921 70975
rect 24967 70929 25025 70975
rect 25071 70929 25129 70975
rect 25175 70929 25233 70975
rect 25279 70929 25337 70975
rect 25383 70929 25441 70975
rect 25487 70929 25545 70975
rect 25591 70929 25649 70975
rect 25695 70929 25753 70975
rect 25799 70929 25857 70975
rect 25903 70929 25961 70975
rect 26007 70929 26065 70975
rect 26111 70929 26169 70975
rect 26215 70929 26273 70975
rect 26319 70929 26377 70975
rect 26423 70929 26481 70975
rect 26527 70929 26585 70975
rect 26631 70929 26689 70975
rect 26735 70929 26793 70975
rect 26839 70929 26897 70975
rect 26943 70929 27001 70975
rect 27047 70929 27105 70975
rect 27151 70929 27209 70975
rect 27255 70929 27313 70975
rect 27359 70929 27417 70975
rect 27463 70929 27521 70975
rect 27567 70929 27625 70975
rect 27671 70929 27729 70975
rect 27775 70929 27833 70975
rect 27879 70929 27937 70975
rect 27983 70929 28041 70975
rect 28087 70929 28145 70975
rect 28191 70929 28249 70975
rect 28295 70929 28353 70975
rect 28399 70929 28457 70975
rect 28503 70929 28561 70975
rect 28607 70929 28665 70975
rect 28711 70929 28769 70975
rect 28815 70929 28873 70975
rect 28919 70929 28977 70975
rect 29023 70929 29081 70975
rect 29127 70929 29185 70975
rect 29231 70929 29289 70975
rect 29335 70929 29393 70975
rect 29439 70929 29497 70975
rect 29543 70929 29601 70975
rect 29647 70929 29705 70975
rect 29751 70929 29809 70975
rect 29855 70929 29913 70975
rect 29959 70929 30017 70975
rect 30063 70929 30121 70975
rect 30167 70929 30225 70975
rect 30271 70929 30329 70975
rect 30375 70929 30433 70975
rect 30479 70929 30537 70975
rect 30583 70929 30641 70975
rect 30687 70929 30745 70975
rect 30791 70929 30849 70975
rect 30895 70929 30953 70975
rect 30999 70929 31057 70975
rect 31103 70929 31161 70975
rect 31207 70929 31265 70975
rect 31311 70929 31369 70975
rect 31415 70929 31473 70975
rect 31519 70929 31577 70975
rect 31623 70929 31681 70975
rect 31727 70929 31785 70975
rect 31831 70929 31889 70975
rect 31935 70929 31993 70975
rect 32039 70929 32097 70975
rect 32143 70929 32201 70975
rect 32247 70929 32305 70975
rect 32351 70929 32409 70975
rect 32455 70929 32513 70975
rect 32559 70929 32617 70975
rect 32663 70929 32721 70975
rect 32767 70929 32825 70975
rect 32871 70929 32929 70975
rect 32975 70929 33033 70975
rect 33079 70929 33137 70975
rect 33183 70929 33241 70975
rect 33287 70929 33345 70975
rect 33391 70929 33449 70975
rect 33495 70929 33553 70975
rect 33599 70929 33657 70975
rect 33703 70929 33761 70975
rect 33807 70929 33865 70975
rect 33911 70929 33969 70975
rect 34015 70929 34073 70975
rect 34119 70929 34177 70975
rect 34223 70929 34281 70975
rect 34327 70929 34385 70975
rect 34431 70929 34489 70975
rect 34535 70929 34593 70975
rect 34639 70929 34697 70975
rect 34743 70929 34801 70975
rect 34847 70929 34905 70975
rect 34951 70929 35009 70975
rect 35055 70929 35113 70975
rect 35159 70929 35217 70975
rect 35263 70929 35321 70975
rect 35367 70929 35425 70975
rect 35471 70929 35529 70975
rect 35575 70929 35633 70975
rect 35679 70929 35737 70975
rect 35783 70929 35841 70975
rect 35887 70929 35945 70975
rect 35991 70929 36049 70975
rect 36095 70929 36153 70975
rect 36199 70929 36257 70975
rect 36303 70929 36361 70975
rect 36407 70929 36465 70975
rect 36511 70929 36569 70975
rect 36615 70929 36673 70975
rect 36719 70929 36777 70975
rect 36823 70929 36881 70975
rect 36927 70929 36985 70975
rect 37031 70929 37089 70975
rect 37135 70929 37193 70975
rect 37239 70929 37297 70975
rect 37343 70929 37401 70975
rect 37447 70929 37505 70975
rect 37551 70929 37609 70975
rect 37655 70929 37713 70975
rect 37759 70929 37817 70975
rect 37863 70929 37921 70975
rect 37967 70929 38025 70975
rect 38071 70929 38129 70975
rect 38175 70929 38233 70975
rect 38279 70929 38337 70975
rect 38383 70929 38441 70975
rect 38487 70929 38545 70975
rect 38591 70929 38649 70975
rect 38695 70929 38753 70975
rect 38799 70929 38857 70975
rect 38903 70929 38961 70975
rect 39007 70929 39065 70975
rect 39111 70929 39169 70975
rect 39215 70929 39273 70975
rect 39319 70929 39377 70975
rect 39423 70929 39481 70975
rect 39527 70929 39585 70975
rect 39631 70929 39689 70975
rect 39735 70929 39793 70975
rect 39839 70929 39897 70975
rect 39943 70929 40001 70975
rect 40047 70929 40105 70975
rect 40151 70929 40209 70975
rect 40255 70929 40313 70975
rect 40359 70929 40417 70975
rect 40463 70929 40521 70975
rect 40567 70929 40625 70975
rect 40671 70929 40729 70975
rect 40775 70929 40833 70975
rect 40879 70929 40937 70975
rect 40983 70929 41041 70975
rect 41087 70929 41145 70975
rect 41191 70929 41249 70975
rect 41295 70929 41353 70975
rect 41399 70929 41457 70975
rect 41503 70929 41561 70975
rect 41607 70929 41665 70975
rect 41711 70929 41769 70975
rect 41815 70929 41873 70975
rect 41919 70929 41977 70975
rect 42023 70929 42081 70975
rect 42127 70929 42185 70975
rect 42231 70929 42289 70975
rect 42335 70929 42393 70975
rect 42439 70929 42497 70975
rect 42543 70929 42601 70975
rect 42647 70929 42705 70975
rect 42751 70929 42809 70975
rect 42855 70929 42913 70975
rect 42959 70929 43017 70975
rect 43063 70929 43121 70975
rect 43167 70929 43225 70975
rect 43271 70929 43329 70975
rect 43375 70929 43433 70975
rect 43479 70929 43537 70975
rect 43583 70929 43641 70975
rect 43687 70929 43745 70975
rect 43791 70929 43849 70975
rect 43895 70929 43953 70975
rect 43999 70929 44057 70975
rect 44103 70929 44161 70975
rect 44207 70929 44265 70975
rect 44311 70929 44369 70975
rect 44415 70929 44473 70975
rect 44519 70929 44577 70975
rect 44623 70929 44681 70975
rect 44727 70929 44785 70975
rect 44831 70929 44889 70975
rect 44935 70929 44993 70975
rect 45039 70929 45097 70975
rect 45143 70929 45201 70975
rect 45247 70929 45305 70975
rect 45351 70929 45409 70975
rect 45455 70929 45513 70975
rect 45559 70929 45617 70975
rect 45663 70929 45721 70975
rect 45767 70929 45825 70975
rect 45871 70929 45929 70975
rect 45975 70929 46033 70975
rect 46079 70929 46137 70975
rect 46183 70929 46241 70975
rect 46287 70929 46345 70975
rect 46391 70929 46449 70975
rect 46495 70929 46553 70975
rect 46599 70929 46657 70975
rect 46703 70929 46761 70975
rect 46807 70929 46865 70975
rect 46911 70929 46969 70975
rect 47015 70929 47073 70975
rect 47119 70929 47177 70975
rect 47223 70929 47281 70975
rect 47327 70929 47385 70975
rect 47431 70929 47489 70975
rect 47535 70929 47593 70975
rect 47639 70929 47697 70975
rect 47743 70929 47801 70975
rect 47847 70929 47905 70975
rect 47951 70929 48009 70975
rect 48055 70929 48113 70975
rect 48159 70929 48217 70975
rect 48263 70929 48321 70975
rect 48367 70929 48425 70975
rect 48471 70929 48529 70975
rect 48575 70929 48633 70975
rect 48679 70929 48737 70975
rect 48783 70929 48841 70975
rect 48887 70929 48945 70975
rect 48991 70929 49049 70975
rect 49095 70929 49153 70975
rect 49199 70929 49257 70975
rect 49303 70929 49361 70975
rect 49407 70929 49465 70975
rect 49511 70929 49569 70975
rect 49615 70929 49673 70975
rect 49719 70929 49777 70975
rect 49823 70929 49881 70975
rect 49927 70929 49985 70975
rect 50031 70929 50089 70975
rect 50135 70929 50193 70975
rect 50239 70929 50297 70975
rect 50343 70929 50401 70975
rect 50447 70929 50505 70975
rect 50551 70929 50609 70975
rect 50655 70929 50713 70975
rect 50759 70929 50817 70975
rect 50863 70929 50921 70975
rect 50967 70929 51025 70975
rect 51071 70929 51129 70975
rect 51175 70929 51233 70975
rect 51279 70929 51337 70975
rect 51383 70929 51441 70975
rect 51487 70929 51545 70975
rect 51591 70929 51649 70975
rect 51695 70929 51753 70975
rect 51799 70929 51857 70975
rect 51903 70929 51961 70975
rect 52007 70929 52065 70975
rect 52111 70929 52169 70975
rect 52215 70929 52273 70975
rect 52319 70929 52377 70975
rect 52423 70929 52481 70975
rect 52527 70929 52585 70975
rect 52631 70929 52689 70975
rect 52735 70929 52793 70975
rect 52839 70929 52897 70975
rect 52943 70929 53001 70975
rect 53047 70929 53105 70975
rect 53151 70929 53209 70975
rect 53255 70929 53313 70975
rect 53359 70929 53417 70975
rect 53463 70929 53521 70975
rect 53567 70929 53625 70975
rect 53671 70929 53729 70975
rect 53775 70929 53833 70975
rect 53879 70929 53937 70975
rect 53983 70929 54041 70975
rect 54087 70929 54145 70975
rect 54191 70929 54249 70975
rect 54295 70929 54353 70975
rect 54399 70929 54457 70975
rect 54503 70929 54561 70975
rect 54607 70929 54665 70975
rect 54711 70929 54769 70975
rect 54815 70929 54873 70975
rect 54919 70929 54977 70975
rect 55023 70929 55081 70975
rect 55127 70929 55185 70975
rect 55231 70929 55289 70975
rect 55335 70929 55393 70975
rect 55439 70929 55497 70975
rect 55543 70929 55601 70975
rect 55647 70929 55705 70975
rect 55751 70929 55809 70975
rect 55855 70929 55913 70975
rect 55959 70929 56017 70975
rect 56063 70929 56121 70975
rect 56167 70929 56225 70975
rect 56271 70929 56329 70975
rect 56375 70929 56433 70975
rect 56479 70929 56537 70975
rect 56583 70929 56641 70975
rect 56687 70929 56745 70975
rect 56791 70929 56849 70975
rect 56895 70929 56953 70975
rect 56999 70929 57057 70975
rect 57103 70929 57161 70975
rect 57207 70929 57265 70975
rect 57311 70929 57369 70975
rect 57415 70929 57473 70975
rect 57519 70929 57577 70975
rect 57623 70929 57681 70975
rect 57727 70929 57785 70975
rect 57831 70929 57889 70975
rect 57935 70929 57993 70975
rect 58039 70929 58097 70975
rect 58143 70929 58201 70975
rect 58247 70929 58305 70975
rect 58351 70929 58409 70975
rect 58455 70929 58513 70975
rect 58559 70929 58617 70975
rect 58663 70929 58721 70975
rect 58767 70929 58825 70975
rect 58871 70929 58929 70975
rect 58975 70929 59033 70975
rect 59079 70929 59137 70975
rect 59183 70929 59241 70975
rect 59287 70929 59345 70975
rect 59391 70929 59449 70975
rect 59495 70929 59553 70975
rect 59599 70929 59657 70975
rect 59703 70929 59761 70975
rect 59807 70929 59865 70975
rect 59911 70929 59969 70975
rect 60015 70929 60073 70975
rect 60119 70929 60177 70975
rect 60223 70929 60281 70975
rect 60327 70929 60385 70975
rect 60431 70929 60489 70975
rect 60535 70929 60593 70975
rect 60639 70929 60697 70975
rect 60743 70929 60801 70975
rect 60847 70929 60905 70975
rect 60951 70929 61009 70975
rect 61055 70929 61113 70975
rect 61159 70929 61217 70975
rect 61263 70929 61321 70975
rect 61367 70929 61425 70975
rect 61471 70929 61529 70975
rect 61575 70929 61633 70975
rect 61679 70929 61737 70975
rect 61783 70929 61841 70975
rect 61887 70929 61945 70975
rect 61991 70929 62049 70975
rect 62095 70929 62153 70975
rect 62199 70929 62257 70975
rect 62303 70929 62361 70975
rect 62407 70929 62465 70975
rect 62511 70929 62569 70975
rect 62615 70929 62673 70975
rect 62719 70929 62777 70975
rect 62823 70929 62881 70975
rect 62927 70929 62985 70975
rect 63031 70929 63089 70975
rect 63135 70929 63193 70975
rect 63239 70929 63297 70975
rect 63343 70929 63401 70975
rect 63447 70929 63505 70975
rect 63551 70929 63609 70975
rect 63655 70929 63713 70975
rect 63759 70929 63817 70975
rect 63863 70929 63921 70975
rect 63967 70929 64025 70975
rect 64071 70929 64129 70975
rect 64175 70929 64233 70975
rect 64279 70929 64337 70975
rect 64383 70929 64441 70975
rect 64487 70929 64545 70975
rect 64591 70929 64649 70975
rect 64695 70929 64753 70975
rect 64799 70929 64857 70975
rect 64903 70929 64961 70975
rect 65007 70929 65065 70975
rect 65111 70929 65169 70975
rect 65215 70929 65273 70975
rect 65319 70929 65377 70975
rect 65423 70929 65481 70975
rect 65527 70929 65585 70975
rect 65631 70929 65689 70975
rect 65735 70929 65793 70975
rect 65839 70929 65897 70975
rect 65943 70929 66001 70975
rect 66047 70929 66105 70975
rect 66151 70929 66209 70975
rect 66255 70929 66313 70975
rect 66359 70929 66417 70975
rect 66463 70929 66521 70975
rect 66567 70929 66625 70975
rect 66671 70929 66729 70975
rect 66775 70929 66833 70975
rect 66879 70929 66937 70975
rect 66983 70929 67041 70975
rect 67087 70929 67145 70975
rect 67191 70929 67249 70975
rect 67295 70929 67353 70975
rect 67399 70929 67457 70975
rect 67503 70929 67561 70975
rect 67607 70929 67665 70975
rect 67711 70929 67769 70975
rect 67815 70929 67873 70975
rect 67919 70929 67977 70975
rect 68023 70929 68081 70975
rect 68127 70929 68185 70975
rect 68231 70929 68289 70975
rect 68335 70929 68393 70975
rect 68439 70929 68497 70975
rect 68543 70929 68601 70975
rect 68647 70929 68705 70975
rect 68751 70929 68809 70975
rect 68855 70929 68913 70975
rect 68959 70929 69017 70975
rect 69063 70929 69121 70975
rect 69167 70929 69225 70975
rect 69271 70929 69329 70975
rect 69375 70929 69433 70975
rect 69479 70929 69537 70975
rect 69583 70929 69641 70975
rect 69687 70929 69745 70975
rect 69791 70929 69849 70975
rect 69895 70929 69957 70975
rect 13108 70871 69957 70929
rect 13108 70825 13119 70871
rect 13165 70825 13223 70871
rect 13269 70825 13377 70871
rect 13423 70825 13481 70871
rect 13527 70825 13585 70871
rect 13631 70825 13689 70871
rect 13735 70825 13793 70871
rect 13839 70825 13897 70871
rect 13943 70825 14001 70871
rect 14047 70825 14105 70871
rect 14151 70825 14209 70871
rect 14255 70825 14313 70871
rect 14359 70825 14417 70871
rect 14463 70825 14521 70871
rect 14567 70825 14625 70871
rect 14671 70825 14729 70871
rect 14775 70825 14833 70871
rect 14879 70825 14937 70871
rect 14983 70825 15041 70871
rect 15087 70825 15145 70871
rect 15191 70825 15249 70871
rect 15295 70825 15353 70871
rect 15399 70825 15457 70871
rect 15503 70825 15561 70871
rect 15607 70825 15665 70871
rect 15711 70825 15769 70871
rect 15815 70825 15873 70871
rect 15919 70825 15977 70871
rect 16023 70825 16081 70871
rect 16127 70825 16185 70871
rect 16231 70825 16289 70871
rect 16335 70825 16393 70871
rect 16439 70825 16497 70871
rect 16543 70825 16601 70871
rect 16647 70825 16705 70871
rect 16751 70825 16809 70871
rect 16855 70825 16913 70871
rect 16959 70825 17017 70871
rect 17063 70825 17121 70871
rect 17167 70825 17225 70871
rect 17271 70825 17329 70871
rect 17375 70825 17433 70871
rect 17479 70825 17537 70871
rect 17583 70825 17641 70871
rect 17687 70825 17745 70871
rect 17791 70825 17849 70871
rect 17895 70825 17953 70871
rect 17999 70825 18057 70871
rect 18103 70825 18161 70871
rect 18207 70825 18265 70871
rect 18311 70825 18369 70871
rect 18415 70825 18473 70871
rect 18519 70825 18577 70871
rect 18623 70825 18681 70871
rect 18727 70825 18785 70871
rect 18831 70825 18889 70871
rect 18935 70825 18993 70871
rect 19039 70825 19097 70871
rect 19143 70825 19201 70871
rect 19247 70825 19305 70871
rect 19351 70825 19409 70871
rect 19455 70825 19513 70871
rect 19559 70825 19617 70871
rect 19663 70825 19721 70871
rect 19767 70825 19825 70871
rect 19871 70825 19929 70871
rect 19975 70825 20033 70871
rect 20079 70825 20137 70871
rect 20183 70825 20241 70871
rect 20287 70825 20345 70871
rect 20391 70825 20449 70871
rect 20495 70825 20553 70871
rect 20599 70825 20657 70871
rect 20703 70825 20761 70871
rect 20807 70825 20865 70871
rect 20911 70825 20969 70871
rect 21015 70825 21073 70871
rect 21119 70825 21177 70871
rect 21223 70825 21281 70871
rect 21327 70825 21385 70871
rect 21431 70825 21489 70871
rect 21535 70825 21593 70871
rect 21639 70825 21697 70871
rect 21743 70825 21801 70871
rect 21847 70825 21905 70871
rect 21951 70825 22009 70871
rect 22055 70825 22113 70871
rect 22159 70825 22217 70871
rect 22263 70825 22321 70871
rect 22367 70825 22425 70871
rect 22471 70825 22529 70871
rect 22575 70825 22633 70871
rect 22679 70825 22737 70871
rect 22783 70825 22841 70871
rect 22887 70825 22945 70871
rect 22991 70825 23049 70871
rect 23095 70825 23153 70871
rect 23199 70825 23257 70871
rect 23303 70825 23361 70871
rect 23407 70825 23465 70871
rect 23511 70825 23569 70871
rect 23615 70825 23673 70871
rect 23719 70825 23777 70871
rect 23823 70825 23881 70871
rect 23927 70825 23985 70871
rect 24031 70825 24089 70871
rect 24135 70825 24193 70871
rect 24239 70825 24297 70871
rect 24343 70825 24401 70871
rect 24447 70825 24505 70871
rect 24551 70825 24609 70871
rect 24655 70825 24713 70871
rect 24759 70825 24817 70871
rect 24863 70825 24921 70871
rect 24967 70825 25025 70871
rect 25071 70825 25129 70871
rect 25175 70825 25233 70871
rect 25279 70825 25337 70871
rect 25383 70825 25441 70871
rect 25487 70825 25545 70871
rect 25591 70825 25649 70871
rect 25695 70825 25753 70871
rect 25799 70825 25857 70871
rect 25903 70825 25961 70871
rect 26007 70825 26065 70871
rect 26111 70825 26169 70871
rect 26215 70825 26273 70871
rect 26319 70825 26377 70871
rect 26423 70825 26481 70871
rect 26527 70825 26585 70871
rect 26631 70825 26689 70871
rect 26735 70825 26793 70871
rect 26839 70825 26897 70871
rect 26943 70825 27001 70871
rect 27047 70825 27105 70871
rect 27151 70825 27209 70871
rect 27255 70825 27313 70871
rect 27359 70825 27417 70871
rect 27463 70825 27521 70871
rect 27567 70825 27625 70871
rect 27671 70825 27729 70871
rect 27775 70825 27833 70871
rect 27879 70825 27937 70871
rect 27983 70825 28041 70871
rect 28087 70825 28145 70871
rect 28191 70825 28249 70871
rect 28295 70825 28353 70871
rect 28399 70825 28457 70871
rect 28503 70825 28561 70871
rect 28607 70825 28665 70871
rect 28711 70825 28769 70871
rect 28815 70825 28873 70871
rect 28919 70825 28977 70871
rect 29023 70825 29081 70871
rect 29127 70825 29185 70871
rect 29231 70825 29289 70871
rect 29335 70825 29393 70871
rect 29439 70825 29497 70871
rect 29543 70825 29601 70871
rect 29647 70825 29705 70871
rect 29751 70825 29809 70871
rect 29855 70825 29913 70871
rect 29959 70825 30017 70871
rect 30063 70825 30121 70871
rect 30167 70825 30225 70871
rect 30271 70825 30329 70871
rect 30375 70825 30433 70871
rect 30479 70825 30537 70871
rect 30583 70825 30641 70871
rect 30687 70825 30745 70871
rect 30791 70825 30849 70871
rect 30895 70825 30953 70871
rect 30999 70825 31057 70871
rect 31103 70825 31161 70871
rect 31207 70825 31265 70871
rect 31311 70825 31369 70871
rect 31415 70825 31473 70871
rect 31519 70825 31577 70871
rect 31623 70825 31681 70871
rect 31727 70825 31785 70871
rect 31831 70825 31889 70871
rect 31935 70825 31993 70871
rect 32039 70825 32097 70871
rect 32143 70825 32201 70871
rect 32247 70825 32305 70871
rect 32351 70825 32409 70871
rect 32455 70825 32513 70871
rect 32559 70825 32617 70871
rect 32663 70825 32721 70871
rect 32767 70825 32825 70871
rect 32871 70825 32929 70871
rect 32975 70825 33033 70871
rect 33079 70825 33137 70871
rect 33183 70825 33241 70871
rect 33287 70825 33345 70871
rect 33391 70825 33449 70871
rect 33495 70825 33553 70871
rect 33599 70825 33657 70871
rect 33703 70825 33761 70871
rect 33807 70825 33865 70871
rect 33911 70825 33969 70871
rect 34015 70825 34073 70871
rect 34119 70825 34177 70871
rect 34223 70825 34281 70871
rect 34327 70825 34385 70871
rect 34431 70825 34489 70871
rect 34535 70825 34593 70871
rect 34639 70825 34697 70871
rect 34743 70825 34801 70871
rect 34847 70825 34905 70871
rect 34951 70825 35009 70871
rect 35055 70825 35113 70871
rect 35159 70825 35217 70871
rect 35263 70825 35321 70871
rect 35367 70825 35425 70871
rect 35471 70825 35529 70871
rect 35575 70825 35633 70871
rect 35679 70825 35737 70871
rect 35783 70825 35841 70871
rect 35887 70825 35945 70871
rect 35991 70825 36049 70871
rect 36095 70825 36153 70871
rect 36199 70825 36257 70871
rect 36303 70825 36361 70871
rect 36407 70825 36465 70871
rect 36511 70825 36569 70871
rect 36615 70825 36673 70871
rect 36719 70825 36777 70871
rect 36823 70825 36881 70871
rect 36927 70825 36985 70871
rect 37031 70825 37089 70871
rect 37135 70825 37193 70871
rect 37239 70825 37297 70871
rect 37343 70825 37401 70871
rect 37447 70825 37505 70871
rect 37551 70825 37609 70871
rect 37655 70825 37713 70871
rect 37759 70825 37817 70871
rect 37863 70825 37921 70871
rect 37967 70825 38025 70871
rect 38071 70825 38129 70871
rect 38175 70825 38233 70871
rect 38279 70825 38337 70871
rect 38383 70825 38441 70871
rect 38487 70825 38545 70871
rect 38591 70825 38649 70871
rect 38695 70825 38753 70871
rect 38799 70825 38857 70871
rect 38903 70825 38961 70871
rect 39007 70825 39065 70871
rect 39111 70825 39169 70871
rect 39215 70825 39273 70871
rect 39319 70825 39377 70871
rect 39423 70825 39481 70871
rect 39527 70825 39585 70871
rect 39631 70825 39689 70871
rect 39735 70825 39793 70871
rect 39839 70825 39897 70871
rect 39943 70825 40001 70871
rect 40047 70825 40105 70871
rect 40151 70825 40209 70871
rect 40255 70825 40313 70871
rect 40359 70825 40417 70871
rect 40463 70825 40521 70871
rect 40567 70825 40625 70871
rect 40671 70825 40729 70871
rect 40775 70825 40833 70871
rect 40879 70825 40937 70871
rect 40983 70825 41041 70871
rect 41087 70825 41145 70871
rect 41191 70825 41249 70871
rect 41295 70825 41353 70871
rect 41399 70825 41457 70871
rect 41503 70825 41561 70871
rect 41607 70825 41665 70871
rect 41711 70825 41769 70871
rect 41815 70825 41873 70871
rect 41919 70825 41977 70871
rect 42023 70825 42081 70871
rect 42127 70825 42185 70871
rect 42231 70825 42289 70871
rect 42335 70825 42393 70871
rect 42439 70825 42497 70871
rect 42543 70825 42601 70871
rect 42647 70825 42705 70871
rect 42751 70825 42809 70871
rect 42855 70825 42913 70871
rect 42959 70825 43017 70871
rect 43063 70825 43121 70871
rect 43167 70825 43225 70871
rect 43271 70825 43329 70871
rect 43375 70825 43433 70871
rect 43479 70825 43537 70871
rect 43583 70825 43641 70871
rect 43687 70825 43745 70871
rect 43791 70825 43849 70871
rect 43895 70825 43953 70871
rect 43999 70825 44057 70871
rect 44103 70825 44161 70871
rect 44207 70825 44265 70871
rect 44311 70825 44369 70871
rect 44415 70825 44473 70871
rect 44519 70825 44577 70871
rect 44623 70825 44681 70871
rect 44727 70825 44785 70871
rect 44831 70825 44889 70871
rect 44935 70825 44993 70871
rect 45039 70825 45097 70871
rect 45143 70825 45201 70871
rect 45247 70825 45305 70871
rect 45351 70825 45409 70871
rect 45455 70825 45513 70871
rect 45559 70825 45617 70871
rect 45663 70825 45721 70871
rect 45767 70825 45825 70871
rect 45871 70825 45929 70871
rect 45975 70825 46033 70871
rect 46079 70825 46137 70871
rect 46183 70825 46241 70871
rect 46287 70825 46345 70871
rect 46391 70825 46449 70871
rect 46495 70825 46553 70871
rect 46599 70825 46657 70871
rect 46703 70825 46761 70871
rect 46807 70825 46865 70871
rect 46911 70825 46969 70871
rect 47015 70825 47073 70871
rect 47119 70825 47177 70871
rect 47223 70825 47281 70871
rect 47327 70825 47385 70871
rect 47431 70825 47489 70871
rect 47535 70825 47593 70871
rect 47639 70825 47697 70871
rect 47743 70825 47801 70871
rect 47847 70825 47905 70871
rect 47951 70825 48009 70871
rect 48055 70825 48113 70871
rect 48159 70825 48217 70871
rect 48263 70825 48321 70871
rect 48367 70825 48425 70871
rect 48471 70825 48529 70871
rect 48575 70825 48633 70871
rect 48679 70825 48737 70871
rect 48783 70825 48841 70871
rect 48887 70825 48945 70871
rect 48991 70825 49049 70871
rect 49095 70825 49153 70871
rect 49199 70825 49257 70871
rect 49303 70825 49361 70871
rect 49407 70825 49465 70871
rect 49511 70825 49569 70871
rect 49615 70825 49673 70871
rect 49719 70825 49777 70871
rect 49823 70825 49881 70871
rect 49927 70825 49985 70871
rect 50031 70825 50089 70871
rect 50135 70825 50193 70871
rect 50239 70825 50297 70871
rect 50343 70825 50401 70871
rect 50447 70825 50505 70871
rect 50551 70825 50609 70871
rect 50655 70825 50713 70871
rect 50759 70825 50817 70871
rect 50863 70825 50921 70871
rect 50967 70825 51025 70871
rect 51071 70825 51129 70871
rect 51175 70825 51233 70871
rect 51279 70825 51337 70871
rect 51383 70825 51441 70871
rect 51487 70825 51545 70871
rect 51591 70825 51649 70871
rect 51695 70825 51753 70871
rect 51799 70825 51857 70871
rect 51903 70825 51961 70871
rect 52007 70825 52065 70871
rect 52111 70825 52169 70871
rect 52215 70825 52273 70871
rect 52319 70825 52377 70871
rect 52423 70825 52481 70871
rect 52527 70825 52585 70871
rect 52631 70825 52689 70871
rect 52735 70825 52793 70871
rect 52839 70825 52897 70871
rect 52943 70825 53001 70871
rect 53047 70825 53105 70871
rect 53151 70825 53209 70871
rect 53255 70825 53313 70871
rect 53359 70825 53417 70871
rect 53463 70825 53521 70871
rect 53567 70825 53625 70871
rect 53671 70825 53729 70871
rect 53775 70825 53833 70871
rect 53879 70825 53937 70871
rect 53983 70825 54041 70871
rect 54087 70825 54145 70871
rect 54191 70825 54249 70871
rect 54295 70825 54353 70871
rect 54399 70825 54457 70871
rect 54503 70825 54561 70871
rect 54607 70825 54665 70871
rect 54711 70825 54769 70871
rect 54815 70825 54873 70871
rect 54919 70825 54977 70871
rect 55023 70825 55081 70871
rect 55127 70825 55185 70871
rect 55231 70825 55289 70871
rect 55335 70825 55393 70871
rect 55439 70825 55497 70871
rect 55543 70825 55601 70871
rect 55647 70825 55705 70871
rect 55751 70825 55809 70871
rect 55855 70825 55913 70871
rect 55959 70825 56017 70871
rect 56063 70825 56121 70871
rect 56167 70825 56225 70871
rect 56271 70825 56329 70871
rect 56375 70825 56433 70871
rect 56479 70825 56537 70871
rect 56583 70825 56641 70871
rect 56687 70825 56745 70871
rect 56791 70825 56849 70871
rect 56895 70825 56953 70871
rect 56999 70825 57057 70871
rect 57103 70825 57161 70871
rect 57207 70825 57265 70871
rect 57311 70825 57369 70871
rect 57415 70825 57473 70871
rect 57519 70825 57577 70871
rect 57623 70825 57681 70871
rect 57727 70825 57785 70871
rect 57831 70825 57889 70871
rect 57935 70825 57993 70871
rect 58039 70825 58097 70871
rect 58143 70825 58201 70871
rect 58247 70825 58305 70871
rect 58351 70825 58409 70871
rect 58455 70825 58513 70871
rect 58559 70825 58617 70871
rect 58663 70825 58721 70871
rect 58767 70825 58825 70871
rect 58871 70825 58929 70871
rect 58975 70825 59033 70871
rect 59079 70825 59137 70871
rect 59183 70825 59241 70871
rect 59287 70825 59345 70871
rect 59391 70825 59449 70871
rect 59495 70825 59553 70871
rect 59599 70825 59657 70871
rect 59703 70825 59761 70871
rect 59807 70825 59865 70871
rect 59911 70825 59969 70871
rect 60015 70825 60073 70871
rect 60119 70825 60177 70871
rect 60223 70825 60281 70871
rect 60327 70825 60385 70871
rect 60431 70825 60489 70871
rect 60535 70825 60593 70871
rect 60639 70825 60697 70871
rect 60743 70825 60801 70871
rect 60847 70825 60905 70871
rect 60951 70825 61009 70871
rect 61055 70825 61113 70871
rect 61159 70825 61217 70871
rect 61263 70825 61321 70871
rect 61367 70825 61425 70871
rect 61471 70825 61529 70871
rect 61575 70825 61633 70871
rect 61679 70825 61737 70871
rect 61783 70825 61841 70871
rect 61887 70825 61945 70871
rect 61991 70825 62049 70871
rect 62095 70825 62153 70871
rect 62199 70825 62257 70871
rect 62303 70825 62361 70871
rect 62407 70825 62465 70871
rect 62511 70825 62569 70871
rect 62615 70825 62673 70871
rect 62719 70825 62777 70871
rect 62823 70825 62881 70871
rect 62927 70825 62985 70871
rect 63031 70825 63089 70871
rect 63135 70825 63193 70871
rect 63239 70825 63297 70871
rect 63343 70825 63401 70871
rect 63447 70825 63505 70871
rect 63551 70825 63609 70871
rect 63655 70825 63713 70871
rect 63759 70825 63817 70871
rect 63863 70825 63921 70871
rect 63967 70825 64025 70871
rect 64071 70825 64129 70871
rect 64175 70825 64233 70871
rect 64279 70825 64337 70871
rect 64383 70825 64441 70871
rect 64487 70825 64545 70871
rect 64591 70825 64649 70871
rect 64695 70825 64753 70871
rect 64799 70825 64857 70871
rect 64903 70825 64961 70871
rect 65007 70825 65065 70871
rect 65111 70825 65169 70871
rect 65215 70825 65273 70871
rect 65319 70825 65377 70871
rect 65423 70825 65481 70871
rect 65527 70825 65585 70871
rect 65631 70825 65689 70871
rect 65735 70825 65793 70871
rect 65839 70825 65897 70871
rect 65943 70825 66001 70871
rect 66047 70825 66105 70871
rect 66151 70825 66209 70871
rect 66255 70825 66313 70871
rect 66359 70825 66417 70871
rect 66463 70825 66521 70871
rect 66567 70825 66625 70871
rect 66671 70825 66729 70871
rect 66775 70825 66833 70871
rect 66879 70825 66937 70871
rect 66983 70825 67041 70871
rect 67087 70825 67145 70871
rect 67191 70825 67249 70871
rect 67295 70825 67353 70871
rect 67399 70825 67457 70871
rect 67503 70825 67561 70871
rect 67607 70825 67665 70871
rect 67711 70825 67769 70871
rect 67815 70825 67873 70871
rect 67919 70825 67977 70871
rect 68023 70825 68081 70871
rect 68127 70825 68185 70871
rect 68231 70825 68289 70871
rect 68335 70825 68393 70871
rect 68439 70825 68497 70871
rect 68543 70825 68601 70871
rect 68647 70825 68705 70871
rect 68751 70825 68809 70871
rect 68855 70825 68913 70871
rect 68959 70825 69017 70871
rect 69063 70825 69121 70871
rect 69167 70825 69225 70871
rect 69271 70825 69329 70871
rect 69375 70825 69433 70871
rect 69479 70825 69537 70871
rect 69583 70825 69641 70871
rect 69687 70825 69745 70871
rect 69791 70825 69849 70871
rect 69895 70825 69957 70871
rect 13108 70814 69957 70825
rect 13108 70767 13280 70814
rect 13108 70721 13119 70767
rect 13165 70721 13223 70767
rect 13269 70721 13280 70767
rect 13108 70663 13280 70721
rect 13108 70617 13119 70663
rect 13165 70617 13223 70663
rect 13269 70617 13280 70663
rect 13108 70559 13280 70617
rect 13108 70513 13119 70559
rect 13165 70513 13223 70559
rect 13269 70513 13280 70559
rect 13108 70455 13280 70513
rect 13108 70409 13119 70455
rect 13165 70409 13223 70455
rect 13269 70409 13280 70455
rect 13108 70351 13280 70409
rect 13108 70305 13119 70351
rect 13165 70305 13223 70351
rect 13269 70305 13280 70351
rect 13108 70247 13280 70305
rect 13108 70201 13119 70247
rect 13165 70201 13223 70247
rect 13269 70201 13280 70247
rect 13108 70143 13280 70201
rect 13108 70097 13119 70143
rect 13165 70097 13223 70143
rect 13269 70097 13280 70143
rect 13108 70039 13280 70097
rect 13108 69993 13119 70039
rect 13165 69993 13223 70039
rect 13269 69993 13280 70039
rect 13108 69935 13280 69993
rect 13108 69889 13119 69935
rect 13165 69889 13223 69935
rect 13269 69889 13280 69935
rect 13108 69831 13280 69889
rect 13108 69785 13119 69831
rect 13165 69785 13223 69831
rect 13269 69785 13280 69831
rect 69785 70720 69957 70814
rect 69785 70674 69796 70720
rect 69842 70674 69900 70720
rect 69946 70674 69957 70720
rect 69785 70616 69957 70674
rect 69785 70570 69796 70616
rect 69842 70570 69900 70616
rect 69946 70570 69957 70616
rect 69785 70512 69957 70570
rect 69785 70466 69796 70512
rect 69842 70466 69900 70512
rect 69946 70466 69957 70512
rect 69785 70408 69957 70466
rect 69785 70362 69796 70408
rect 69842 70362 69900 70408
rect 69946 70362 69957 70408
rect 69785 70304 69957 70362
rect 69785 70258 69796 70304
rect 69842 70258 69900 70304
rect 69946 70258 69957 70304
rect 69785 70200 69957 70258
rect 69785 70154 69796 70200
rect 69842 70154 69900 70200
rect 69946 70154 69957 70200
rect 69785 70096 69957 70154
rect 69785 70050 69796 70096
rect 69842 70050 69900 70096
rect 69946 70050 69957 70096
rect 69785 69957 69957 70050
rect 69785 69946 71000 69957
rect 69785 69900 69796 69946
rect 69842 69900 69900 69946
rect 69946 69900 70004 69946
rect 70050 69900 70108 69946
rect 70154 69900 70212 69946
rect 70258 69900 70316 69946
rect 70362 69900 70420 69946
rect 70466 69900 70524 69946
rect 70570 69900 70628 69946
rect 70674 69908 71000 69946
rect 70674 69900 70824 69908
rect 69785 69862 70824 69900
rect 70870 69862 70928 69908
rect 70974 69862 71000 69908
rect 69785 69842 71000 69862
rect 69785 69796 69796 69842
rect 69842 69796 69900 69842
rect 69946 69796 70004 69842
rect 70050 69796 70108 69842
rect 70154 69796 70212 69842
rect 70258 69796 70316 69842
rect 70362 69796 70420 69842
rect 70466 69796 70524 69842
rect 70570 69796 70628 69842
rect 70674 69804 71000 69842
rect 70674 69796 70824 69804
rect 69785 69785 70824 69796
rect 13108 69727 13280 69785
rect 13108 69681 13119 69727
rect 13165 69681 13223 69727
rect 13269 69681 13280 69727
rect 13108 69623 13280 69681
rect 13108 69577 13119 69623
rect 13165 69577 13223 69623
rect 13269 69577 13280 69623
rect 13108 69519 13280 69577
rect 13108 69473 13119 69519
rect 13165 69473 13223 69519
rect 13269 69473 13280 69519
rect 13108 69415 13280 69473
rect 13108 69369 13119 69415
rect 13165 69369 13223 69415
rect 13269 69369 13280 69415
rect 13108 69311 13280 69369
rect 13108 69265 13119 69311
rect 13165 69265 13223 69311
rect 13269 69265 13280 69311
rect 13108 69207 13280 69265
rect 13108 69161 13119 69207
rect 13165 69161 13223 69207
rect 13269 69161 13280 69207
rect 13108 69103 13280 69161
rect 13108 69057 13119 69103
rect 13165 69057 13223 69103
rect 13269 69057 13280 69103
rect 13108 68999 13280 69057
rect 13108 68953 13119 68999
rect 13165 68953 13223 68999
rect 13269 68953 13280 68999
rect 13108 68895 13280 68953
rect 13108 68849 13119 68895
rect 13165 68849 13223 68895
rect 13269 68849 13280 68895
rect 13108 68791 13280 68849
rect 13108 68745 13119 68791
rect 13165 68745 13223 68791
rect 13269 68745 13280 68791
rect 13108 68687 13280 68745
rect 13108 68641 13119 68687
rect 13165 68641 13223 68687
rect 13269 68641 13280 68687
rect 13108 68583 13280 68641
rect 13108 68537 13119 68583
rect 13165 68537 13223 68583
rect 13269 68537 13280 68583
rect 13108 68479 13280 68537
rect 13108 68433 13119 68479
rect 13165 68433 13223 68479
rect 13269 68433 13280 68479
rect 13108 68375 13280 68433
rect 13108 68329 13119 68375
rect 13165 68329 13223 68375
rect 13269 68329 13280 68375
rect 13108 68271 13280 68329
rect 13108 68225 13119 68271
rect 13165 68225 13223 68271
rect 13269 68225 13280 68271
rect 13108 68167 13280 68225
rect 13108 68121 13119 68167
rect 13165 68121 13223 68167
rect 13269 68121 13280 68167
rect 13108 68063 13280 68121
rect 13108 68017 13119 68063
rect 13165 68017 13223 68063
rect 13269 68017 13280 68063
rect 13108 67959 13280 68017
rect 13108 67913 13119 67959
rect 13165 67913 13223 67959
rect 13269 67913 13280 67959
rect 13108 67855 13280 67913
rect 13108 67809 13119 67855
rect 13165 67809 13223 67855
rect 13269 67809 13280 67855
rect 13108 67751 13280 67809
rect 13108 67705 13119 67751
rect 13165 67705 13223 67751
rect 13269 67705 13280 67751
rect 13108 67647 13280 67705
rect 13108 67601 13119 67647
rect 13165 67601 13223 67647
rect 13269 67601 13280 67647
rect 13108 67543 13280 67601
rect 13108 67497 13119 67543
rect 13165 67497 13223 67543
rect 13269 67497 13280 67543
rect 13108 67439 13280 67497
rect 13108 67393 13119 67439
rect 13165 67393 13223 67439
rect 13269 67393 13280 67439
rect 13108 67335 13280 67393
rect 13108 67289 13119 67335
rect 13165 67289 13223 67335
rect 13269 67289 13280 67335
rect 13108 67231 13280 67289
rect 13108 67185 13119 67231
rect 13165 67185 13223 67231
rect 13269 67185 13280 67231
rect 13108 67127 13280 67185
rect 13108 67081 13119 67127
rect 13165 67081 13223 67127
rect 13269 67081 13280 67127
rect 13108 67023 13280 67081
rect 13108 66977 13119 67023
rect 13165 66977 13223 67023
rect 13269 66977 13280 67023
rect 13108 66919 13280 66977
rect 13108 66873 13119 66919
rect 13165 66873 13223 66919
rect 13269 66873 13280 66919
rect 13108 66815 13280 66873
rect 13108 66769 13119 66815
rect 13165 66769 13223 66815
rect 13269 66769 13280 66815
rect 13108 66711 13280 66769
rect 13108 66665 13119 66711
rect 13165 66665 13223 66711
rect 13269 66665 13280 66711
rect 13108 66607 13280 66665
rect 13108 66561 13119 66607
rect 13165 66561 13223 66607
rect 13269 66561 13280 66607
rect 13108 66503 13280 66561
rect 13108 66457 13119 66503
rect 13165 66457 13223 66503
rect 13269 66457 13280 66503
rect 13108 66399 13280 66457
rect 13108 66353 13119 66399
rect 13165 66353 13223 66399
rect 13269 66353 13280 66399
rect 13108 66295 13280 66353
rect 13108 66249 13119 66295
rect 13165 66249 13223 66295
rect 13269 66249 13280 66295
rect 13108 66191 13280 66249
rect 13108 66145 13119 66191
rect 13165 66145 13223 66191
rect 13269 66145 13280 66191
rect 13108 66087 13280 66145
rect 13108 66041 13119 66087
rect 13165 66041 13223 66087
rect 13269 66041 13280 66087
rect 13108 65983 13280 66041
rect 13108 65937 13119 65983
rect 13165 65937 13223 65983
rect 13269 65937 13280 65983
rect 13108 65879 13280 65937
rect 13108 65833 13119 65879
rect 13165 65833 13223 65879
rect 13269 65833 13280 65879
rect 13108 65775 13280 65833
rect 13108 65729 13119 65775
rect 13165 65729 13223 65775
rect 13269 65729 13280 65775
rect 13108 65671 13280 65729
rect 13108 65625 13119 65671
rect 13165 65625 13223 65671
rect 13269 65625 13280 65671
rect 13108 65567 13280 65625
rect 13108 65521 13119 65567
rect 13165 65521 13223 65567
rect 13269 65521 13280 65567
rect 13108 65463 13280 65521
rect 13108 65417 13119 65463
rect 13165 65417 13223 65463
rect 13269 65417 13280 65463
rect 13108 65359 13280 65417
rect 13108 65313 13119 65359
rect 13165 65313 13223 65359
rect 13269 65313 13280 65359
rect 13108 65255 13280 65313
rect 13108 65209 13119 65255
rect 13165 65209 13223 65255
rect 13269 65209 13280 65255
rect 13108 65151 13280 65209
rect 13108 65105 13119 65151
rect 13165 65105 13223 65151
rect 13269 65105 13280 65151
rect 13108 65047 13280 65105
rect 13108 65001 13119 65047
rect 13165 65001 13223 65047
rect 13269 65001 13280 65047
rect 13108 64943 13280 65001
rect 13108 64897 13119 64943
rect 13165 64897 13223 64943
rect 13269 64897 13280 64943
rect 13108 64839 13280 64897
rect 13108 64793 13119 64839
rect 13165 64793 13223 64839
rect 13269 64793 13280 64839
rect 13108 64735 13280 64793
rect 13108 64689 13119 64735
rect 13165 64689 13223 64735
rect 13269 64689 13280 64735
rect 13108 64631 13280 64689
rect 13108 64585 13119 64631
rect 13165 64585 13223 64631
rect 13269 64585 13280 64631
rect 13108 64527 13280 64585
rect 13108 64481 13119 64527
rect 13165 64481 13223 64527
rect 13269 64481 13280 64527
rect 13108 64423 13280 64481
rect 13108 64377 13119 64423
rect 13165 64377 13223 64423
rect 13269 64377 13280 64423
rect 13108 64319 13280 64377
rect 13108 64273 13119 64319
rect 13165 64273 13223 64319
rect 13269 64273 13280 64319
rect 13108 64215 13280 64273
rect 13108 64169 13119 64215
rect 13165 64169 13223 64215
rect 13269 64169 13280 64215
rect 13108 64111 13280 64169
rect 13108 64065 13119 64111
rect 13165 64065 13223 64111
rect 13269 64065 13280 64111
rect 13108 64007 13280 64065
rect 13108 63961 13119 64007
rect 13165 63961 13223 64007
rect 13269 63961 13280 64007
rect 13108 63903 13280 63961
rect 13108 63857 13119 63903
rect 13165 63857 13223 63903
rect 13269 63857 13280 63903
rect 13108 63799 13280 63857
rect 13108 63753 13119 63799
rect 13165 63753 13223 63799
rect 13269 63753 13280 63799
rect 13108 63695 13280 63753
rect 13108 63649 13119 63695
rect 13165 63649 13223 63695
rect 13269 63649 13280 63695
rect 13108 63591 13280 63649
rect 13108 63545 13119 63591
rect 13165 63545 13223 63591
rect 13269 63545 13280 63591
rect 13108 63487 13280 63545
rect 13108 63441 13119 63487
rect 13165 63441 13223 63487
rect 13269 63441 13280 63487
rect 13108 63383 13280 63441
rect 13108 63337 13119 63383
rect 13165 63337 13223 63383
rect 13269 63337 13280 63383
rect 13108 63279 13280 63337
rect 13108 63233 13119 63279
rect 13165 63233 13223 63279
rect 13269 63233 13280 63279
rect 13108 63175 13280 63233
rect 13108 63129 13119 63175
rect 13165 63129 13223 63175
rect 13269 63129 13280 63175
rect 13108 63071 13280 63129
rect 13108 63025 13119 63071
rect 13165 63025 13223 63071
rect 13269 63025 13280 63071
rect 13108 62967 13280 63025
rect 13108 62921 13119 62967
rect 13165 62921 13223 62967
rect 13269 62921 13280 62967
rect 13108 62863 13280 62921
rect 13108 62817 13119 62863
rect 13165 62817 13223 62863
rect 13269 62817 13280 62863
rect 13108 62759 13280 62817
rect 13108 62713 13119 62759
rect 13165 62713 13223 62759
rect 13269 62713 13280 62759
rect 13108 62655 13280 62713
rect 13108 62609 13119 62655
rect 13165 62609 13223 62655
rect 13269 62609 13280 62655
rect 13108 62551 13280 62609
rect 13108 62505 13119 62551
rect 13165 62505 13223 62551
rect 13269 62505 13280 62551
rect 13108 62447 13280 62505
rect 13108 62401 13119 62447
rect 13165 62401 13223 62447
rect 13269 62401 13280 62447
rect 13108 62343 13280 62401
rect 13108 62297 13119 62343
rect 13165 62297 13223 62343
rect 13269 62297 13280 62343
rect 13108 62239 13280 62297
rect 13108 62193 13119 62239
rect 13165 62193 13223 62239
rect 13269 62193 13280 62239
rect 13108 62135 13280 62193
rect 13108 62089 13119 62135
rect 13165 62089 13223 62135
rect 13269 62089 13280 62135
rect 13108 62031 13280 62089
rect 13108 61985 13119 62031
rect 13165 61985 13223 62031
rect 13269 61985 13280 62031
rect 13108 61927 13280 61985
rect 13108 61881 13119 61927
rect 13165 61881 13223 61927
rect 13269 61881 13280 61927
rect 13108 61823 13280 61881
rect 13108 61777 13119 61823
rect 13165 61777 13223 61823
rect 13269 61777 13280 61823
rect 13108 61719 13280 61777
rect 13108 61673 13119 61719
rect 13165 61673 13223 61719
rect 13269 61673 13280 61719
rect 13108 61615 13280 61673
rect 13108 61569 13119 61615
rect 13165 61569 13223 61615
rect 13269 61569 13280 61615
rect 13108 61511 13280 61569
rect 13108 61465 13119 61511
rect 13165 61465 13223 61511
rect 13269 61465 13280 61511
rect 13108 61407 13280 61465
rect 13108 61361 13119 61407
rect 13165 61361 13223 61407
rect 13269 61361 13280 61407
rect 13108 61303 13280 61361
rect 13108 61257 13119 61303
rect 13165 61257 13223 61303
rect 13269 61257 13280 61303
rect 13108 61199 13280 61257
rect 13108 61153 13119 61199
rect 13165 61153 13223 61199
rect 13269 61153 13280 61199
rect 13108 61095 13280 61153
rect 13108 61049 13119 61095
rect 13165 61049 13223 61095
rect 13269 61049 13280 61095
rect 13108 60991 13280 61049
rect 13108 60945 13119 60991
rect 13165 60945 13223 60991
rect 13269 60945 13280 60991
rect 13108 60887 13280 60945
rect 13108 60841 13119 60887
rect 13165 60841 13223 60887
rect 13269 60841 13280 60887
rect 13108 60783 13280 60841
rect 13108 60737 13119 60783
rect 13165 60737 13223 60783
rect 13269 60737 13280 60783
rect 13108 60679 13280 60737
rect 13108 60633 13119 60679
rect 13165 60633 13223 60679
rect 13269 60633 13280 60679
rect 13108 60575 13280 60633
rect 13108 60529 13119 60575
rect 13165 60529 13223 60575
rect 13269 60529 13280 60575
rect 13108 60471 13280 60529
rect 13108 60425 13119 60471
rect 13165 60425 13223 60471
rect 13269 60425 13280 60471
rect 13108 60367 13280 60425
rect 13108 60321 13119 60367
rect 13165 60321 13223 60367
rect 13269 60321 13280 60367
rect 13108 60263 13280 60321
rect 13108 60217 13119 60263
rect 13165 60217 13223 60263
rect 13269 60217 13280 60263
rect 13108 60159 13280 60217
rect 13108 60113 13119 60159
rect 13165 60113 13223 60159
rect 13269 60113 13280 60159
rect 13108 60055 13280 60113
rect 13108 60009 13119 60055
rect 13165 60009 13223 60055
rect 13269 60009 13280 60055
rect 13108 59951 13280 60009
rect 13108 59905 13119 59951
rect 13165 59905 13223 59951
rect 13269 59905 13280 59951
rect 13108 59847 13280 59905
rect 13108 59801 13119 59847
rect 13165 59801 13223 59847
rect 13269 59801 13280 59847
rect 13108 59743 13280 59801
rect 13108 59697 13119 59743
rect 13165 59697 13223 59743
rect 13269 59697 13280 59743
rect 13108 59639 13280 59697
rect 13108 59593 13119 59639
rect 13165 59593 13223 59639
rect 13269 59593 13280 59639
rect 13108 59535 13280 59593
rect 13108 59489 13119 59535
rect 13165 59489 13223 59535
rect 13269 59489 13280 59535
rect 13108 59431 13280 59489
rect 13108 59385 13119 59431
rect 13165 59385 13223 59431
rect 13269 59385 13280 59431
rect 13108 59327 13280 59385
rect 13108 59281 13119 59327
rect 13165 59281 13223 59327
rect 13269 59281 13280 59327
rect 13108 59223 13280 59281
rect 13108 59177 13119 59223
rect 13165 59177 13223 59223
rect 13269 59177 13280 59223
rect 13108 59119 13280 59177
rect 13108 59073 13119 59119
rect 13165 59073 13223 59119
rect 13269 59073 13280 59119
rect 13108 59015 13280 59073
rect 13108 58969 13119 59015
rect 13165 58969 13223 59015
rect 13269 58969 13280 59015
rect 13108 58911 13280 58969
rect 13108 58865 13119 58911
rect 13165 58865 13223 58911
rect 13269 58865 13280 58911
rect 13108 58807 13280 58865
rect 13108 58761 13119 58807
rect 13165 58761 13223 58807
rect 13269 58761 13280 58807
rect 13108 58703 13280 58761
rect 13108 58657 13119 58703
rect 13165 58657 13223 58703
rect 13269 58657 13280 58703
rect 13108 58599 13280 58657
rect 13108 58553 13119 58599
rect 13165 58553 13223 58599
rect 13269 58553 13280 58599
rect 13108 58495 13280 58553
rect 13108 58449 13119 58495
rect 13165 58449 13223 58495
rect 13269 58449 13280 58495
rect 13108 58391 13280 58449
rect 13108 58345 13119 58391
rect 13165 58345 13223 58391
rect 13269 58345 13280 58391
rect 13108 58287 13280 58345
rect 13108 58241 13119 58287
rect 13165 58241 13223 58287
rect 13269 58241 13280 58287
rect 13108 58183 13280 58241
rect 13108 58137 13119 58183
rect 13165 58137 13223 58183
rect 13269 58137 13280 58183
rect 13108 58079 13280 58137
rect 13108 58033 13119 58079
rect 13165 58033 13223 58079
rect 13269 58033 13280 58079
rect 13108 57975 13280 58033
rect 13108 57929 13119 57975
rect 13165 57929 13223 57975
rect 13269 57929 13280 57975
rect 13108 57871 13280 57929
rect 13108 57825 13119 57871
rect 13165 57825 13223 57871
rect 13269 57825 13280 57871
rect 13108 57767 13280 57825
rect 13108 57721 13119 57767
rect 13165 57721 13223 57767
rect 13269 57721 13280 57767
rect 13108 57663 13280 57721
rect 13108 57617 13119 57663
rect 13165 57617 13223 57663
rect 13269 57617 13280 57663
rect 13108 57559 13280 57617
rect 13108 57513 13119 57559
rect 13165 57513 13223 57559
rect 13269 57513 13280 57559
rect 13108 57455 13280 57513
rect 13108 57409 13119 57455
rect 13165 57409 13223 57455
rect 13269 57409 13280 57455
rect 13108 57351 13280 57409
rect 13108 57305 13119 57351
rect 13165 57305 13223 57351
rect 13269 57305 13280 57351
rect 13108 57247 13280 57305
rect 13108 57201 13119 57247
rect 13165 57201 13223 57247
rect 13269 57201 13280 57247
rect 13108 57143 13280 57201
rect 13108 57097 13119 57143
rect 13165 57097 13223 57143
rect 13269 57097 13280 57143
rect 13108 57039 13280 57097
rect 13108 56993 13119 57039
rect 13165 56993 13223 57039
rect 13269 56993 13280 57039
rect 13108 56935 13280 56993
rect 13108 56889 13119 56935
rect 13165 56889 13223 56935
rect 13269 56889 13280 56935
rect 13108 56831 13280 56889
rect 13108 56785 13119 56831
rect 13165 56785 13223 56831
rect 13269 56785 13280 56831
rect 13108 56727 13280 56785
rect 13108 56681 13119 56727
rect 13165 56681 13223 56727
rect 13269 56681 13280 56727
rect 13108 56623 13280 56681
rect 13108 56577 13119 56623
rect 13165 56577 13223 56623
rect 13269 56577 13280 56623
rect 13108 56519 13280 56577
rect 13108 56473 13119 56519
rect 13165 56473 13223 56519
rect 13269 56473 13280 56519
rect 13108 56415 13280 56473
rect 13108 56369 13119 56415
rect 13165 56369 13223 56415
rect 13269 56369 13280 56415
rect 13108 56311 13280 56369
rect 13108 56265 13119 56311
rect 13165 56265 13223 56311
rect 13269 56265 13280 56311
rect 13108 56207 13280 56265
rect 13108 56161 13119 56207
rect 13165 56161 13223 56207
rect 13269 56161 13280 56207
rect 13108 56103 13280 56161
rect 13108 56057 13119 56103
rect 13165 56057 13223 56103
rect 13269 56057 13280 56103
rect 13108 55999 13280 56057
rect 13108 55953 13119 55999
rect 13165 55953 13223 55999
rect 13269 55953 13280 55999
rect 13108 55895 13280 55953
rect 13108 55849 13119 55895
rect 13165 55849 13223 55895
rect 13269 55849 13280 55895
rect 13108 55791 13280 55849
rect 13108 55745 13119 55791
rect 13165 55745 13223 55791
rect 13269 55745 13280 55791
rect 13108 55687 13280 55745
rect 13108 55641 13119 55687
rect 13165 55641 13223 55687
rect 13269 55641 13280 55687
rect 13108 55583 13280 55641
rect 13108 55537 13119 55583
rect 13165 55537 13223 55583
rect 13269 55537 13280 55583
rect 13108 55479 13280 55537
rect 13108 55433 13119 55479
rect 13165 55433 13223 55479
rect 13269 55433 13280 55479
rect 13108 55375 13280 55433
rect 13108 55329 13119 55375
rect 13165 55329 13223 55375
rect 13269 55329 13280 55375
rect 13108 55271 13280 55329
rect 13108 55225 13119 55271
rect 13165 55225 13223 55271
rect 13269 55225 13280 55271
rect 13108 55167 13280 55225
rect 13108 55121 13119 55167
rect 13165 55121 13223 55167
rect 13269 55121 13280 55167
rect 13108 55063 13280 55121
rect 13108 55017 13119 55063
rect 13165 55017 13223 55063
rect 13269 55017 13280 55063
rect 13108 54959 13280 55017
rect 13108 54913 13119 54959
rect 13165 54913 13223 54959
rect 13269 54913 13280 54959
rect 13108 54855 13280 54913
rect 13108 54809 13119 54855
rect 13165 54809 13223 54855
rect 13269 54809 13280 54855
rect 13108 54751 13280 54809
rect 13108 54705 13119 54751
rect 13165 54705 13223 54751
rect 13269 54705 13280 54751
rect 13108 54647 13280 54705
rect 13108 54601 13119 54647
rect 13165 54601 13223 54647
rect 13269 54601 13280 54647
rect 13108 54543 13280 54601
rect 13108 54497 13119 54543
rect 13165 54497 13223 54543
rect 13269 54497 13280 54543
rect 13108 54439 13280 54497
rect 13108 54393 13119 54439
rect 13165 54393 13223 54439
rect 13269 54393 13280 54439
rect 13108 54335 13280 54393
rect 13108 54289 13119 54335
rect 13165 54289 13223 54335
rect 13269 54289 13280 54335
rect 13108 54231 13280 54289
rect 13108 54185 13119 54231
rect 13165 54185 13223 54231
rect 13269 54185 13280 54231
rect 13108 54127 13280 54185
rect 13108 54081 13119 54127
rect 13165 54081 13223 54127
rect 13269 54081 13280 54127
rect 13108 54023 13280 54081
rect 13108 53977 13119 54023
rect 13165 53977 13223 54023
rect 13269 53977 13280 54023
rect 13108 53919 13280 53977
rect 13108 53873 13119 53919
rect 13165 53873 13223 53919
rect 13269 53873 13280 53919
rect 13108 53815 13280 53873
rect 13108 53769 13119 53815
rect 13165 53769 13223 53815
rect 13269 53769 13280 53815
rect 13108 53711 13280 53769
rect 13108 53665 13119 53711
rect 13165 53665 13223 53711
rect 13269 53665 13280 53711
rect 13108 53607 13280 53665
rect 13108 53561 13119 53607
rect 13165 53561 13223 53607
rect 13269 53561 13280 53607
rect 13108 53503 13280 53561
rect 13108 53457 13119 53503
rect 13165 53457 13223 53503
rect 13269 53457 13280 53503
rect 13108 53399 13280 53457
rect 13108 53353 13119 53399
rect 13165 53353 13223 53399
rect 13269 53353 13280 53399
rect 13108 53295 13280 53353
rect 13108 53249 13119 53295
rect 13165 53249 13223 53295
rect 13269 53249 13280 53295
rect 13108 53191 13280 53249
rect 13108 53145 13119 53191
rect 13165 53145 13223 53191
rect 13269 53145 13280 53191
rect 13108 53087 13280 53145
rect 13108 53041 13119 53087
rect 13165 53041 13223 53087
rect 13269 53041 13280 53087
rect 13108 52983 13280 53041
rect 13108 52937 13119 52983
rect 13165 52937 13223 52983
rect 13269 52937 13280 52983
rect 13108 52879 13280 52937
rect 13108 52833 13119 52879
rect 13165 52833 13223 52879
rect 13269 52833 13280 52879
rect 13108 52775 13280 52833
rect 13108 52729 13119 52775
rect 13165 52729 13223 52775
rect 13269 52729 13280 52775
rect 13108 52671 13280 52729
rect 13108 52625 13119 52671
rect 13165 52625 13223 52671
rect 13269 52625 13280 52671
rect 13108 52567 13280 52625
rect 13108 52521 13119 52567
rect 13165 52521 13223 52567
rect 13269 52521 13280 52567
rect 13108 52463 13280 52521
rect 13108 52417 13119 52463
rect 13165 52417 13223 52463
rect 13269 52417 13280 52463
rect 13108 52359 13280 52417
rect 13108 52313 13119 52359
rect 13165 52313 13223 52359
rect 13269 52313 13280 52359
rect 13108 52255 13280 52313
rect 13108 52209 13119 52255
rect 13165 52209 13223 52255
rect 13269 52209 13280 52255
rect 13108 52151 13280 52209
rect 13108 52105 13119 52151
rect 13165 52105 13223 52151
rect 13269 52105 13280 52151
rect 13108 52047 13280 52105
rect 13108 52001 13119 52047
rect 13165 52001 13223 52047
rect 13269 52001 13280 52047
rect 13108 51943 13280 52001
rect 13108 51897 13119 51943
rect 13165 51897 13223 51943
rect 13269 51897 13280 51943
rect 13108 51839 13280 51897
rect 13108 51793 13119 51839
rect 13165 51793 13223 51839
rect 13269 51793 13280 51839
rect 13108 51735 13280 51793
rect 13108 51689 13119 51735
rect 13165 51689 13223 51735
rect 13269 51689 13280 51735
rect 13108 51631 13280 51689
rect 13108 51585 13119 51631
rect 13165 51585 13223 51631
rect 13269 51585 13280 51631
rect 13108 51527 13280 51585
rect 13108 51481 13119 51527
rect 13165 51481 13223 51527
rect 13269 51481 13280 51527
rect 13108 51423 13280 51481
rect 13108 51377 13119 51423
rect 13165 51377 13223 51423
rect 13269 51377 13280 51423
rect 13108 51319 13280 51377
rect 13108 51273 13119 51319
rect 13165 51273 13223 51319
rect 13269 51273 13280 51319
rect 13108 51215 13280 51273
rect 13108 51169 13119 51215
rect 13165 51169 13223 51215
rect 13269 51169 13280 51215
rect 13108 51111 13280 51169
rect 13108 51065 13119 51111
rect 13165 51065 13223 51111
rect 13269 51065 13280 51111
rect 13108 51007 13280 51065
rect 13108 50961 13119 51007
rect 13165 50961 13223 51007
rect 13269 50961 13280 51007
rect 13108 50903 13280 50961
rect 13108 50857 13119 50903
rect 13165 50857 13223 50903
rect 13269 50857 13280 50903
rect 13108 50799 13280 50857
rect 13108 50753 13119 50799
rect 13165 50753 13223 50799
rect 13269 50753 13280 50799
rect 13108 50695 13280 50753
rect 13108 50649 13119 50695
rect 13165 50649 13223 50695
rect 13269 50649 13280 50695
rect 13108 50591 13280 50649
rect 13108 50545 13119 50591
rect 13165 50545 13223 50591
rect 13269 50545 13280 50591
rect 13108 50487 13280 50545
rect 13108 50441 13119 50487
rect 13165 50441 13223 50487
rect 13269 50441 13280 50487
rect 13108 50383 13280 50441
rect 13108 50337 13119 50383
rect 13165 50337 13223 50383
rect 13269 50337 13280 50383
rect 13108 50279 13280 50337
rect 13108 50233 13119 50279
rect 13165 50233 13223 50279
rect 13269 50233 13280 50279
rect 13108 50175 13280 50233
rect 13108 50129 13119 50175
rect 13165 50129 13223 50175
rect 13269 50129 13280 50175
rect 13108 50071 13280 50129
rect 13108 50025 13119 50071
rect 13165 50025 13223 50071
rect 13269 50025 13280 50071
rect 13108 49967 13280 50025
rect 13108 49921 13119 49967
rect 13165 49921 13223 49967
rect 13269 49921 13280 49967
rect 13108 49863 13280 49921
rect 13108 49817 13119 49863
rect 13165 49817 13223 49863
rect 13269 49817 13280 49863
rect 13108 49759 13280 49817
rect 13108 49713 13119 49759
rect 13165 49713 13223 49759
rect 13269 49713 13280 49759
rect 13108 49655 13280 49713
rect 13108 49609 13119 49655
rect 13165 49609 13223 49655
rect 13269 49609 13280 49655
rect 13108 49551 13280 49609
rect 13108 49505 13119 49551
rect 13165 49505 13223 49551
rect 13269 49505 13280 49551
rect 13108 49447 13280 49505
rect 13108 49401 13119 49447
rect 13165 49401 13223 49447
rect 13269 49401 13280 49447
rect 13108 49343 13280 49401
rect 13108 49297 13119 49343
rect 13165 49297 13223 49343
rect 13269 49297 13280 49343
rect 13108 49239 13280 49297
rect 13108 49193 13119 49239
rect 13165 49193 13223 49239
rect 13269 49193 13280 49239
rect 13108 49135 13280 49193
rect 13108 49089 13119 49135
rect 13165 49089 13223 49135
rect 13269 49089 13280 49135
rect 13108 49031 13280 49089
rect 13108 48985 13119 49031
rect 13165 48985 13223 49031
rect 13269 48985 13280 49031
rect 13108 48927 13280 48985
rect 13108 48881 13119 48927
rect 13165 48881 13223 48927
rect 13269 48881 13280 48927
rect 13108 48823 13280 48881
rect 13108 48777 13119 48823
rect 13165 48777 13223 48823
rect 13269 48777 13280 48823
rect 13108 48719 13280 48777
rect 13108 48673 13119 48719
rect 13165 48673 13223 48719
rect 13269 48673 13280 48719
rect 13108 48615 13280 48673
rect 13108 48569 13119 48615
rect 13165 48569 13223 48615
rect 13269 48569 13280 48615
rect 13108 48511 13280 48569
rect 13108 48465 13119 48511
rect 13165 48465 13223 48511
rect 13269 48465 13280 48511
rect 13108 48407 13280 48465
rect 13108 48361 13119 48407
rect 13165 48361 13223 48407
rect 13269 48361 13280 48407
rect 13108 48303 13280 48361
rect 13108 48257 13119 48303
rect 13165 48257 13223 48303
rect 13269 48257 13280 48303
rect 13108 48199 13280 48257
rect 13108 48153 13119 48199
rect 13165 48153 13223 48199
rect 13269 48153 13280 48199
rect 13108 48095 13280 48153
rect 13108 48049 13119 48095
rect 13165 48049 13223 48095
rect 13269 48049 13280 48095
rect 13108 47991 13280 48049
rect 13108 47945 13119 47991
rect 13165 47945 13223 47991
rect 13269 47945 13280 47991
rect 13108 47887 13280 47945
rect 13108 47841 13119 47887
rect 13165 47841 13223 47887
rect 13269 47841 13280 47887
rect 13108 47783 13280 47841
rect 13108 47737 13119 47783
rect 13165 47737 13223 47783
rect 13269 47737 13280 47783
rect 13108 47679 13280 47737
rect 13108 47633 13119 47679
rect 13165 47633 13223 47679
rect 13269 47633 13280 47679
rect 13108 47575 13280 47633
rect 13108 47529 13119 47575
rect 13165 47529 13223 47575
rect 13269 47529 13280 47575
rect 13108 47471 13280 47529
rect 13108 47425 13119 47471
rect 13165 47425 13223 47471
rect 13269 47425 13280 47471
rect 13108 47367 13280 47425
rect 13108 47321 13119 47367
rect 13165 47321 13223 47367
rect 13269 47321 13280 47367
rect 13108 47263 13280 47321
rect 13108 47217 13119 47263
rect 13165 47217 13223 47263
rect 13269 47217 13280 47263
rect 13108 47159 13280 47217
rect 13108 47113 13119 47159
rect 13165 47113 13223 47159
rect 13269 47113 13280 47159
rect 13108 47055 13280 47113
rect 13108 47009 13119 47055
rect 13165 47009 13223 47055
rect 13269 47009 13280 47055
rect 13108 46951 13280 47009
rect 13108 46905 13119 46951
rect 13165 46905 13223 46951
rect 13269 46905 13280 46951
rect 13108 46847 13280 46905
rect 13108 46801 13119 46847
rect 13165 46801 13223 46847
rect 13269 46801 13280 46847
rect 13108 46743 13280 46801
rect 13108 46697 13119 46743
rect 13165 46697 13223 46743
rect 13269 46697 13280 46743
rect 13108 46639 13280 46697
rect 13108 46593 13119 46639
rect 13165 46593 13223 46639
rect 13269 46593 13280 46639
rect 13108 46535 13280 46593
rect 13108 46489 13119 46535
rect 13165 46489 13223 46535
rect 13269 46489 13280 46535
rect 13108 46431 13280 46489
rect 13108 46385 13119 46431
rect 13165 46385 13223 46431
rect 13269 46385 13280 46431
rect 13108 46327 13280 46385
rect 13108 46281 13119 46327
rect 13165 46281 13223 46327
rect 13269 46281 13280 46327
rect 13108 46223 13280 46281
rect 13108 46177 13119 46223
rect 13165 46177 13223 46223
rect 13269 46177 13280 46223
rect 13108 46119 13280 46177
rect 13108 46073 13119 46119
rect 13165 46073 13223 46119
rect 13269 46073 13280 46119
rect 13108 46015 13280 46073
rect 13108 45969 13119 46015
rect 13165 45969 13223 46015
rect 13269 45969 13280 46015
rect 13108 45911 13280 45969
rect 13108 45865 13119 45911
rect 13165 45865 13223 45911
rect 13269 45865 13280 45911
rect 13108 45807 13280 45865
rect 13108 45761 13119 45807
rect 13165 45761 13223 45807
rect 13269 45761 13280 45807
rect 13108 45703 13280 45761
rect 13108 45657 13119 45703
rect 13165 45657 13223 45703
rect 13269 45657 13280 45703
rect 13108 45599 13280 45657
rect 13108 45553 13119 45599
rect 13165 45553 13223 45599
rect 13269 45553 13280 45599
rect 13108 45495 13280 45553
rect 13108 45449 13119 45495
rect 13165 45449 13223 45495
rect 13269 45449 13280 45495
rect 13108 45391 13280 45449
rect 13108 45345 13119 45391
rect 13165 45345 13223 45391
rect 13269 45345 13280 45391
rect 13108 45287 13280 45345
rect 13108 45241 13119 45287
rect 13165 45241 13223 45287
rect 13269 45241 13280 45287
rect 13108 45183 13280 45241
rect 13108 45137 13119 45183
rect 13165 45137 13223 45183
rect 13269 45137 13280 45183
rect 13108 45079 13280 45137
rect 13108 45033 13119 45079
rect 13165 45033 13223 45079
rect 13269 45033 13280 45079
rect 13108 44848 13280 45033
rect 70813 69758 70824 69785
rect 70870 69758 70928 69804
rect 70974 69758 71000 69804
rect 70813 69700 71000 69758
rect 70813 69654 70824 69700
rect 70870 69654 70928 69700
rect 70974 69654 71000 69700
rect 70813 69596 71000 69654
rect 70813 69550 70824 69596
rect 70870 69550 70928 69596
rect 70974 69550 71000 69596
rect 70813 69492 71000 69550
rect 70813 69446 70824 69492
rect 70870 69446 70928 69492
rect 70974 69446 71000 69492
rect 70813 69388 71000 69446
rect 70813 69342 70824 69388
rect 70870 69342 70928 69388
rect 70974 69342 71000 69388
rect 70813 69284 71000 69342
rect 70813 69238 70824 69284
rect 70870 69238 70928 69284
rect 70974 69238 71000 69284
rect 70813 69180 71000 69238
rect 70813 69134 70824 69180
rect 70870 69134 70928 69180
rect 70974 69134 71000 69180
rect 70813 69076 71000 69134
rect 70813 69030 70824 69076
rect 70870 69030 70928 69076
rect 70974 69030 71000 69076
rect 70813 68972 71000 69030
rect 70813 68926 70824 68972
rect 70870 68926 70928 68972
rect 70974 68926 71000 68972
rect 70813 68868 71000 68926
rect 70813 68822 70824 68868
rect 70870 68822 70928 68868
rect 70974 68822 71000 68868
rect 70813 68764 71000 68822
rect 70813 68718 70824 68764
rect 70870 68718 70928 68764
rect 70974 68718 71000 68764
rect 70813 68660 71000 68718
rect 70813 68614 70824 68660
rect 70870 68614 70928 68660
rect 70974 68614 71000 68660
rect 70813 68556 71000 68614
rect 70813 68510 70824 68556
rect 70870 68510 70928 68556
rect 70974 68510 71000 68556
rect 70813 68452 71000 68510
rect 70813 68406 70824 68452
rect 70870 68406 70928 68452
rect 70974 68406 71000 68452
rect 70813 68348 71000 68406
rect 70813 68302 70824 68348
rect 70870 68302 70928 68348
rect 70974 68302 71000 68348
rect 70813 68244 71000 68302
rect 70813 68198 70824 68244
rect 70870 68198 70928 68244
rect 70974 68198 71000 68244
rect 70813 68140 71000 68198
rect 70813 68094 70824 68140
rect 70870 68094 70928 68140
rect 70974 68094 71000 68140
rect 70813 68036 71000 68094
rect 70813 67990 70824 68036
rect 70870 67990 70928 68036
rect 70974 67990 71000 68036
rect 70813 67932 71000 67990
rect 70813 67886 70824 67932
rect 70870 67886 70928 67932
rect 70974 67886 71000 67932
rect 70813 67828 71000 67886
rect 70813 67782 70824 67828
rect 70870 67782 70928 67828
rect 70974 67782 71000 67828
rect 70813 67724 71000 67782
rect 70813 67678 70824 67724
rect 70870 67678 70928 67724
rect 70974 67678 71000 67724
rect 70813 67620 71000 67678
rect 70813 67574 70824 67620
rect 70870 67574 70928 67620
rect 70974 67574 71000 67620
rect 70813 67516 71000 67574
rect 70813 67470 70824 67516
rect 70870 67470 70928 67516
rect 70974 67470 71000 67516
rect 70813 67412 71000 67470
rect 70813 67366 70824 67412
rect 70870 67366 70928 67412
rect 70974 67366 71000 67412
rect 70813 67308 71000 67366
rect 70813 67262 70824 67308
rect 70870 67262 70928 67308
rect 70974 67262 71000 67308
rect 70813 67204 71000 67262
rect 70813 67158 70824 67204
rect 70870 67158 70928 67204
rect 70974 67158 71000 67204
rect 70813 67100 71000 67158
rect 70813 67054 70824 67100
rect 70870 67054 70928 67100
rect 70974 67054 71000 67100
rect 70813 66996 71000 67054
rect 70813 66950 70824 66996
rect 70870 66950 70928 66996
rect 70974 66950 71000 66996
rect 70813 66892 71000 66950
rect 70813 66846 70824 66892
rect 70870 66846 70928 66892
rect 70974 66846 71000 66892
rect 70813 66788 71000 66846
rect 70813 66742 70824 66788
rect 70870 66742 70928 66788
rect 70974 66742 71000 66788
rect 70813 66684 71000 66742
rect 70813 66638 70824 66684
rect 70870 66638 70928 66684
rect 70974 66638 71000 66684
rect 70813 66580 71000 66638
rect 70813 66534 70824 66580
rect 70870 66534 70928 66580
rect 70974 66534 71000 66580
rect 70813 66476 71000 66534
rect 70813 66430 70824 66476
rect 70870 66430 70928 66476
rect 70974 66430 71000 66476
rect 70813 66372 71000 66430
rect 70813 66326 70824 66372
rect 70870 66326 70928 66372
rect 70974 66326 71000 66372
rect 70813 66268 71000 66326
rect 70813 66222 70824 66268
rect 70870 66222 70928 66268
rect 70974 66222 71000 66268
rect 70813 66164 71000 66222
rect 70813 66118 70824 66164
rect 70870 66118 70928 66164
rect 70974 66118 71000 66164
rect 70813 66060 71000 66118
rect 70813 66014 70824 66060
rect 70870 66014 70928 66060
rect 70974 66014 71000 66060
rect 70813 65956 71000 66014
rect 70813 65910 70824 65956
rect 70870 65910 70928 65956
rect 70974 65910 71000 65956
rect 70813 65852 71000 65910
rect 70813 65806 70824 65852
rect 70870 65806 70928 65852
rect 70974 65806 71000 65852
rect 70813 65748 71000 65806
rect 70813 65702 70824 65748
rect 70870 65702 70928 65748
rect 70974 65702 71000 65748
rect 70813 65644 71000 65702
rect 70813 65598 70824 65644
rect 70870 65598 70928 65644
rect 70974 65598 71000 65644
rect 70813 65540 71000 65598
rect 70813 65494 70824 65540
rect 70870 65494 70928 65540
rect 70974 65494 71000 65540
rect 70813 65436 71000 65494
rect 70813 65390 70824 65436
rect 70870 65390 70928 65436
rect 70974 65390 71000 65436
rect 70813 65332 71000 65390
rect 70813 65286 70824 65332
rect 70870 65286 70928 65332
rect 70974 65286 71000 65332
rect 70813 65228 71000 65286
rect 70813 65182 70824 65228
rect 70870 65182 70928 65228
rect 70974 65182 71000 65228
rect 70813 65124 71000 65182
rect 70813 65078 70824 65124
rect 70870 65078 70928 65124
rect 70974 65078 71000 65124
rect 70813 65020 71000 65078
rect 70813 64974 70824 65020
rect 70870 64974 70928 65020
rect 70974 64974 71000 65020
rect 70813 64916 71000 64974
rect 70813 64870 70824 64916
rect 70870 64870 70928 64916
rect 70974 64870 71000 64916
rect 70813 64812 71000 64870
rect 70813 64766 70824 64812
rect 70870 64766 70928 64812
rect 70974 64766 71000 64812
rect 70813 64708 71000 64766
rect 70813 64662 70824 64708
rect 70870 64662 70928 64708
rect 70974 64662 71000 64708
rect 70813 64604 71000 64662
rect 70813 64558 70824 64604
rect 70870 64558 70928 64604
rect 70974 64558 71000 64604
rect 70813 64500 71000 64558
rect 70813 64454 70824 64500
rect 70870 64454 70928 64500
rect 70974 64454 71000 64500
rect 70813 64396 71000 64454
rect 70813 64350 70824 64396
rect 70870 64350 70928 64396
rect 70974 64350 71000 64396
rect 70813 64292 71000 64350
rect 70813 64246 70824 64292
rect 70870 64246 70928 64292
rect 70974 64246 71000 64292
rect 70813 64188 71000 64246
rect 70813 64142 70824 64188
rect 70870 64142 70928 64188
rect 70974 64142 71000 64188
rect 70813 64084 71000 64142
rect 70813 64038 70824 64084
rect 70870 64038 70928 64084
rect 70974 64038 71000 64084
rect 70813 63980 71000 64038
rect 70813 63934 70824 63980
rect 70870 63934 70928 63980
rect 70974 63934 71000 63980
rect 70813 63876 71000 63934
rect 70813 63830 70824 63876
rect 70870 63830 70928 63876
rect 70974 63830 71000 63876
rect 70813 63772 71000 63830
rect 70813 63726 70824 63772
rect 70870 63726 70928 63772
rect 70974 63726 71000 63772
rect 70813 63668 71000 63726
rect 70813 63622 70824 63668
rect 70870 63622 70928 63668
rect 70974 63622 71000 63668
rect 70813 63564 71000 63622
rect 70813 63518 70824 63564
rect 70870 63518 70928 63564
rect 70974 63518 71000 63564
rect 70813 63460 71000 63518
rect 70813 63414 70824 63460
rect 70870 63414 70928 63460
rect 70974 63414 71000 63460
rect 70813 63356 71000 63414
rect 70813 63310 70824 63356
rect 70870 63310 70928 63356
rect 70974 63310 71000 63356
rect 70813 63252 71000 63310
rect 70813 63206 70824 63252
rect 70870 63206 70928 63252
rect 70974 63206 71000 63252
rect 70813 63148 71000 63206
rect 70813 63102 70824 63148
rect 70870 63102 70928 63148
rect 70974 63102 71000 63148
rect 70813 63044 71000 63102
rect 70813 62998 70824 63044
rect 70870 62998 70928 63044
rect 70974 62998 71000 63044
rect 70813 62940 71000 62998
rect 70813 62894 70824 62940
rect 70870 62894 70928 62940
rect 70974 62894 71000 62940
rect 70813 62836 71000 62894
rect 70813 62790 70824 62836
rect 70870 62790 70928 62836
rect 70974 62790 71000 62836
rect 70813 62732 71000 62790
rect 70813 62686 70824 62732
rect 70870 62686 70928 62732
rect 70974 62686 71000 62732
rect 70813 62628 71000 62686
rect 70813 62582 70824 62628
rect 70870 62582 70928 62628
rect 70974 62582 71000 62628
rect 70813 62524 71000 62582
rect 70813 62478 70824 62524
rect 70870 62478 70928 62524
rect 70974 62478 71000 62524
rect 70813 62420 71000 62478
rect 70813 62374 70824 62420
rect 70870 62374 70928 62420
rect 70974 62374 71000 62420
rect 70813 62316 71000 62374
rect 70813 62270 70824 62316
rect 70870 62270 70928 62316
rect 70974 62270 71000 62316
rect 70813 62212 71000 62270
rect 70813 62166 70824 62212
rect 70870 62166 70928 62212
rect 70974 62166 71000 62212
rect 70813 62108 71000 62166
rect 70813 62062 70824 62108
rect 70870 62062 70928 62108
rect 70974 62062 71000 62108
rect 70813 62004 71000 62062
rect 70813 61958 70824 62004
rect 70870 61958 70928 62004
rect 70974 61958 71000 62004
rect 70813 61900 71000 61958
rect 70813 61854 70824 61900
rect 70870 61854 70928 61900
rect 70974 61854 71000 61900
rect 70813 61796 71000 61854
rect 70813 61750 70824 61796
rect 70870 61750 70928 61796
rect 70974 61750 71000 61796
rect 70813 61692 71000 61750
rect 70813 61646 70824 61692
rect 70870 61646 70928 61692
rect 70974 61646 71000 61692
rect 70813 61588 71000 61646
rect 70813 61542 70824 61588
rect 70870 61542 70928 61588
rect 70974 61542 71000 61588
rect 70813 61484 71000 61542
rect 70813 61438 70824 61484
rect 70870 61438 70928 61484
rect 70974 61438 71000 61484
rect 70813 61380 71000 61438
rect 70813 61334 70824 61380
rect 70870 61334 70928 61380
rect 70974 61334 71000 61380
rect 70813 61276 71000 61334
rect 70813 61230 70824 61276
rect 70870 61230 70928 61276
rect 70974 61230 71000 61276
rect 70813 61172 71000 61230
rect 70813 61126 70824 61172
rect 70870 61126 70928 61172
rect 70974 61126 71000 61172
rect 70813 61068 71000 61126
rect 70813 61022 70824 61068
rect 70870 61022 70928 61068
rect 70974 61022 71000 61068
rect 70813 60964 71000 61022
rect 70813 60918 70824 60964
rect 70870 60918 70928 60964
rect 70974 60918 71000 60964
rect 70813 60860 71000 60918
rect 70813 60814 70824 60860
rect 70870 60814 70928 60860
rect 70974 60814 71000 60860
rect 70813 60756 71000 60814
rect 70813 60710 70824 60756
rect 70870 60710 70928 60756
rect 70974 60710 71000 60756
rect 70813 60652 71000 60710
rect 70813 60606 70824 60652
rect 70870 60606 70928 60652
rect 70974 60606 71000 60652
rect 70813 60548 71000 60606
rect 70813 60502 70824 60548
rect 70870 60502 70928 60548
rect 70974 60502 71000 60548
rect 70813 60444 71000 60502
rect 70813 60398 70824 60444
rect 70870 60398 70928 60444
rect 70974 60398 71000 60444
rect 70813 60340 71000 60398
rect 70813 60294 70824 60340
rect 70870 60294 70928 60340
rect 70974 60294 71000 60340
rect 70813 60236 71000 60294
rect 70813 60190 70824 60236
rect 70870 60190 70928 60236
rect 70974 60190 71000 60236
rect 70813 60132 71000 60190
rect 70813 60086 70824 60132
rect 70870 60086 70928 60132
rect 70974 60086 71000 60132
rect 70813 60028 71000 60086
rect 70813 59982 70824 60028
rect 70870 59982 70928 60028
rect 70974 59982 71000 60028
rect 70813 59924 71000 59982
rect 70813 59878 70824 59924
rect 70870 59878 70928 59924
rect 70974 59878 71000 59924
rect 70813 59820 71000 59878
rect 70813 59774 70824 59820
rect 70870 59774 70928 59820
rect 70974 59774 71000 59820
rect 70813 59716 71000 59774
rect 70813 59670 70824 59716
rect 70870 59670 70928 59716
rect 70974 59670 71000 59716
rect 70813 59612 71000 59670
rect 70813 59566 70824 59612
rect 70870 59566 70928 59612
rect 70974 59566 71000 59612
rect 70813 59508 71000 59566
rect 70813 59462 70824 59508
rect 70870 59462 70928 59508
rect 70974 59462 71000 59508
rect 70813 59404 71000 59462
rect 70813 59358 70824 59404
rect 70870 59358 70928 59404
rect 70974 59358 71000 59404
rect 70813 59300 71000 59358
rect 70813 59254 70824 59300
rect 70870 59254 70928 59300
rect 70974 59254 71000 59300
rect 70813 59196 71000 59254
rect 70813 59150 70824 59196
rect 70870 59150 70928 59196
rect 70974 59150 71000 59196
rect 70813 59092 71000 59150
rect 70813 59046 70824 59092
rect 70870 59046 70928 59092
rect 70974 59046 71000 59092
rect 70813 58988 71000 59046
rect 70813 58942 70824 58988
rect 70870 58942 70928 58988
rect 70974 58942 71000 58988
rect 70813 58884 71000 58942
rect 70813 58838 70824 58884
rect 70870 58838 70928 58884
rect 70974 58838 71000 58884
rect 70813 58780 71000 58838
rect 70813 58734 70824 58780
rect 70870 58734 70928 58780
rect 70974 58734 71000 58780
rect 70813 58676 71000 58734
rect 70813 58630 70824 58676
rect 70870 58630 70928 58676
rect 70974 58630 71000 58676
rect 70813 58572 71000 58630
rect 70813 58526 70824 58572
rect 70870 58526 70928 58572
rect 70974 58526 71000 58572
rect 70813 58468 71000 58526
rect 70813 58422 70824 58468
rect 70870 58422 70928 58468
rect 70974 58422 71000 58468
rect 70813 58364 71000 58422
rect 70813 58318 70824 58364
rect 70870 58318 70928 58364
rect 70974 58318 71000 58364
rect 70813 58260 71000 58318
rect 70813 58214 70824 58260
rect 70870 58214 70928 58260
rect 70974 58214 71000 58260
rect 70813 58156 71000 58214
rect 70813 58110 70824 58156
rect 70870 58110 70928 58156
rect 70974 58110 71000 58156
rect 70813 58052 71000 58110
rect 70813 58006 70824 58052
rect 70870 58006 70928 58052
rect 70974 58006 71000 58052
rect 70813 57948 71000 58006
rect 70813 57902 70824 57948
rect 70870 57902 70928 57948
rect 70974 57902 71000 57948
rect 70813 57844 71000 57902
rect 70813 57798 70824 57844
rect 70870 57798 70928 57844
rect 70974 57798 71000 57844
rect 70813 57740 71000 57798
rect 70813 57694 70824 57740
rect 70870 57694 70928 57740
rect 70974 57694 71000 57740
rect 70813 57636 71000 57694
rect 70813 57590 70824 57636
rect 70870 57590 70928 57636
rect 70974 57590 71000 57636
rect 70813 57532 71000 57590
rect 70813 57486 70824 57532
rect 70870 57486 70928 57532
rect 70974 57486 71000 57532
rect 70813 57428 71000 57486
rect 70813 57382 70824 57428
rect 70870 57382 70928 57428
rect 70974 57382 71000 57428
rect 70813 57324 71000 57382
rect 70813 57278 70824 57324
rect 70870 57278 70928 57324
rect 70974 57278 71000 57324
rect 70813 57220 71000 57278
rect 70813 57174 70824 57220
rect 70870 57174 70928 57220
rect 70974 57174 71000 57220
rect 70813 57116 71000 57174
rect 70813 57070 70824 57116
rect 70870 57070 70928 57116
rect 70974 57070 71000 57116
rect 70813 57012 71000 57070
rect 70813 56966 70824 57012
rect 70870 56966 70928 57012
rect 70974 56966 71000 57012
rect 70813 56908 71000 56966
rect 70813 56862 70824 56908
rect 70870 56862 70928 56908
rect 70974 56862 71000 56908
rect 70813 56804 71000 56862
rect 70813 56758 70824 56804
rect 70870 56758 70928 56804
rect 70974 56758 71000 56804
rect 70813 56700 71000 56758
rect 70813 56654 70824 56700
rect 70870 56654 70928 56700
rect 70974 56654 71000 56700
rect 70813 56596 71000 56654
rect 70813 56550 70824 56596
rect 70870 56550 70928 56596
rect 70974 56550 71000 56596
rect 70813 56492 71000 56550
rect 70813 56446 70824 56492
rect 70870 56446 70928 56492
rect 70974 56446 71000 56492
rect 70813 56388 71000 56446
rect 70813 56342 70824 56388
rect 70870 56342 70928 56388
rect 70974 56342 71000 56388
rect 70813 56284 71000 56342
rect 70813 56238 70824 56284
rect 70870 56238 70928 56284
rect 70974 56238 71000 56284
rect 70813 56180 71000 56238
rect 70813 56134 70824 56180
rect 70870 56134 70928 56180
rect 70974 56134 71000 56180
rect 70813 56076 71000 56134
rect 70813 56030 70824 56076
rect 70870 56030 70928 56076
rect 70974 56030 71000 56076
rect 70813 55972 71000 56030
rect 70813 55926 70824 55972
rect 70870 55926 70928 55972
rect 70974 55926 71000 55972
rect 70813 55868 71000 55926
rect 70813 55822 70824 55868
rect 70870 55822 70928 55868
rect 70974 55822 71000 55868
rect 70813 55764 71000 55822
rect 70813 55718 70824 55764
rect 70870 55718 70928 55764
rect 70974 55718 71000 55764
rect 70813 55660 71000 55718
rect 70813 55614 70824 55660
rect 70870 55614 70928 55660
rect 70974 55614 71000 55660
rect 70813 55556 71000 55614
rect 70813 55510 70824 55556
rect 70870 55510 70928 55556
rect 70974 55510 71000 55556
rect 70813 55452 71000 55510
rect 70813 55406 70824 55452
rect 70870 55406 70928 55452
rect 70974 55406 71000 55452
rect 70813 55348 71000 55406
rect 70813 55302 70824 55348
rect 70870 55302 70928 55348
rect 70974 55302 71000 55348
rect 70813 55244 71000 55302
rect 70813 55198 70824 55244
rect 70870 55198 70928 55244
rect 70974 55198 71000 55244
rect 70813 55140 71000 55198
rect 70813 55094 70824 55140
rect 70870 55094 70928 55140
rect 70974 55094 71000 55140
rect 70813 55036 71000 55094
rect 70813 54990 70824 55036
rect 70870 54990 70928 55036
rect 70974 54990 71000 55036
rect 70813 54932 71000 54990
rect 70813 54886 70824 54932
rect 70870 54886 70928 54932
rect 70974 54886 71000 54932
rect 70813 54828 71000 54886
rect 70813 54782 70824 54828
rect 70870 54782 70928 54828
rect 70974 54782 71000 54828
rect 70813 54724 71000 54782
rect 70813 54678 70824 54724
rect 70870 54678 70928 54724
rect 70974 54678 71000 54724
rect 70813 54620 71000 54678
rect 70813 54574 70824 54620
rect 70870 54574 70928 54620
rect 70974 54574 71000 54620
rect 70813 54516 71000 54574
rect 70813 54470 70824 54516
rect 70870 54470 70928 54516
rect 70974 54470 71000 54516
rect 70813 54412 71000 54470
rect 70813 54366 70824 54412
rect 70870 54366 70928 54412
rect 70974 54366 71000 54412
rect 70813 54308 71000 54366
rect 70813 54262 70824 54308
rect 70870 54262 70928 54308
rect 70974 54262 71000 54308
rect 70813 54204 71000 54262
rect 70813 54158 70824 54204
rect 70870 54158 70928 54204
rect 70974 54158 71000 54204
rect 70813 54100 71000 54158
rect 70813 54054 70824 54100
rect 70870 54054 70928 54100
rect 70974 54054 71000 54100
rect 70813 53996 71000 54054
rect 70813 53950 70824 53996
rect 70870 53950 70928 53996
rect 70974 53950 71000 53996
rect 70813 53892 71000 53950
rect 70813 53846 70824 53892
rect 70870 53846 70928 53892
rect 70974 53846 71000 53892
rect 70813 53788 71000 53846
rect 70813 53742 70824 53788
rect 70870 53742 70928 53788
rect 70974 53742 71000 53788
rect 70813 53684 71000 53742
rect 70813 53638 70824 53684
rect 70870 53638 70928 53684
rect 70974 53638 71000 53684
rect 70813 53580 71000 53638
rect 70813 53534 70824 53580
rect 70870 53534 70928 53580
rect 70974 53534 71000 53580
rect 70813 53476 71000 53534
rect 70813 53430 70824 53476
rect 70870 53430 70928 53476
rect 70974 53430 71000 53476
rect 70813 53372 71000 53430
rect 70813 53326 70824 53372
rect 70870 53326 70928 53372
rect 70974 53326 71000 53372
rect 70813 53268 71000 53326
rect 70813 53222 70824 53268
rect 70870 53222 70928 53268
rect 70974 53222 71000 53268
rect 70813 53164 71000 53222
rect 70813 53118 70824 53164
rect 70870 53118 70928 53164
rect 70974 53118 71000 53164
rect 70813 53060 71000 53118
rect 70813 53014 70824 53060
rect 70870 53014 70928 53060
rect 70974 53014 71000 53060
rect 70813 52956 71000 53014
rect 70813 52910 70824 52956
rect 70870 52910 70928 52956
rect 70974 52910 71000 52956
rect 70813 52852 71000 52910
rect 70813 52806 70824 52852
rect 70870 52806 70928 52852
rect 70974 52806 71000 52852
rect 70813 52748 71000 52806
rect 70813 52702 70824 52748
rect 70870 52702 70928 52748
rect 70974 52702 71000 52748
rect 70813 52644 71000 52702
rect 70813 52598 70824 52644
rect 70870 52598 70928 52644
rect 70974 52598 71000 52644
rect 70813 52540 71000 52598
rect 70813 52494 70824 52540
rect 70870 52494 70928 52540
rect 70974 52494 71000 52540
rect 70813 52436 71000 52494
rect 70813 52390 70824 52436
rect 70870 52390 70928 52436
rect 70974 52390 71000 52436
rect 70813 52332 71000 52390
rect 70813 52286 70824 52332
rect 70870 52286 70928 52332
rect 70974 52286 71000 52332
rect 70813 52228 71000 52286
rect 70813 52182 70824 52228
rect 70870 52182 70928 52228
rect 70974 52182 71000 52228
rect 70813 52124 71000 52182
rect 70813 52078 70824 52124
rect 70870 52078 70928 52124
rect 70974 52078 71000 52124
rect 70813 52020 71000 52078
rect 70813 51974 70824 52020
rect 70870 51974 70928 52020
rect 70974 51974 71000 52020
rect 70813 51916 71000 51974
rect 70813 51870 70824 51916
rect 70870 51870 70928 51916
rect 70974 51870 71000 51916
rect 70813 51812 71000 51870
rect 70813 51766 70824 51812
rect 70870 51766 70928 51812
rect 70974 51766 71000 51812
rect 70813 51708 71000 51766
rect 70813 51662 70824 51708
rect 70870 51662 70928 51708
rect 70974 51662 71000 51708
rect 70813 51604 71000 51662
rect 70813 51558 70824 51604
rect 70870 51558 70928 51604
rect 70974 51558 71000 51604
rect 70813 51500 71000 51558
rect 70813 51454 70824 51500
rect 70870 51454 70928 51500
rect 70974 51454 71000 51500
rect 70813 51396 71000 51454
rect 70813 51350 70824 51396
rect 70870 51350 70928 51396
rect 70974 51350 71000 51396
rect 70813 51292 71000 51350
rect 70813 51246 70824 51292
rect 70870 51246 70928 51292
rect 70974 51246 71000 51292
rect 70813 51188 71000 51246
rect 70813 51142 70824 51188
rect 70870 51142 70928 51188
rect 70974 51142 71000 51188
rect 70813 51084 71000 51142
rect 70813 51038 70824 51084
rect 70870 51038 70928 51084
rect 70974 51038 71000 51084
rect 70813 50980 71000 51038
rect 70813 50934 70824 50980
rect 70870 50934 70928 50980
rect 70974 50934 71000 50980
rect 70813 50876 71000 50934
rect 70813 50830 70824 50876
rect 70870 50830 70928 50876
rect 70974 50830 71000 50876
rect 70813 50772 71000 50830
rect 70813 50726 70824 50772
rect 70870 50726 70928 50772
rect 70974 50726 71000 50772
rect 70813 50668 71000 50726
rect 70813 50622 70824 50668
rect 70870 50622 70928 50668
rect 70974 50622 71000 50668
rect 70813 50564 71000 50622
rect 70813 50518 70824 50564
rect 70870 50518 70928 50564
rect 70974 50518 71000 50564
rect 70813 50460 71000 50518
rect 70813 50414 70824 50460
rect 70870 50414 70928 50460
rect 70974 50414 71000 50460
rect 70813 50356 71000 50414
rect 70813 50310 70824 50356
rect 70870 50310 70928 50356
rect 70974 50310 71000 50356
rect 70813 50252 71000 50310
rect 70813 50206 70824 50252
rect 70870 50206 70928 50252
rect 70974 50206 71000 50252
rect 70813 50148 71000 50206
rect 70813 50102 70824 50148
rect 70870 50102 70928 50148
rect 70974 50102 71000 50148
rect 70813 50044 71000 50102
rect 70813 49998 70824 50044
rect 70870 49998 70928 50044
rect 70974 49998 71000 50044
rect 70813 49940 71000 49998
rect 70813 49894 70824 49940
rect 70870 49894 70928 49940
rect 70974 49894 71000 49940
rect 70813 49836 71000 49894
rect 70813 49790 70824 49836
rect 70870 49790 70928 49836
rect 70974 49790 71000 49836
rect 70813 49732 71000 49790
rect 70813 49686 70824 49732
rect 70870 49686 70928 49732
rect 70974 49686 71000 49732
rect 70813 49628 71000 49686
rect 70813 49582 70824 49628
rect 70870 49582 70928 49628
rect 70974 49582 71000 49628
rect 70813 49524 71000 49582
rect 70813 49478 70824 49524
rect 70870 49478 70928 49524
rect 70974 49478 71000 49524
rect 70813 49420 71000 49478
rect 70813 49374 70824 49420
rect 70870 49374 70928 49420
rect 70974 49374 71000 49420
rect 70813 49316 71000 49374
rect 70813 49270 70824 49316
rect 70870 49270 70928 49316
rect 70974 49270 71000 49316
rect 70813 49212 71000 49270
rect 70813 49166 70824 49212
rect 70870 49166 70928 49212
rect 70974 49166 71000 49212
rect 70813 49108 71000 49166
rect 70813 49062 70824 49108
rect 70870 49062 70928 49108
rect 70974 49062 71000 49108
rect 70813 49004 71000 49062
rect 70813 48958 70824 49004
rect 70870 48958 70928 49004
rect 70974 48958 71000 49004
rect 70813 48900 71000 48958
rect 70813 48854 70824 48900
rect 70870 48854 70928 48900
rect 70974 48854 71000 48900
rect 70813 48796 71000 48854
rect 70813 48750 70824 48796
rect 70870 48750 70928 48796
rect 70974 48750 71000 48796
rect 70813 48692 71000 48750
rect 70813 48646 70824 48692
rect 70870 48646 70928 48692
rect 70974 48646 71000 48692
rect 70813 48588 71000 48646
rect 70813 48542 70824 48588
rect 70870 48542 70928 48588
rect 70974 48542 71000 48588
rect 70813 48484 71000 48542
rect 70813 48438 70824 48484
rect 70870 48438 70928 48484
rect 70974 48438 71000 48484
rect 70813 48380 71000 48438
rect 70813 48334 70824 48380
rect 70870 48334 70928 48380
rect 70974 48334 71000 48380
rect 70813 48276 71000 48334
rect 70813 48230 70824 48276
rect 70870 48230 70928 48276
rect 70974 48230 71000 48276
rect 70813 48172 71000 48230
rect 70813 48126 70824 48172
rect 70870 48126 70928 48172
rect 70974 48126 71000 48172
rect 70813 48068 71000 48126
rect 70813 48022 70824 48068
rect 70870 48022 70928 48068
rect 70974 48022 71000 48068
rect 70813 47964 71000 48022
rect 70813 47918 70824 47964
rect 70870 47918 70928 47964
rect 70974 47918 71000 47964
rect 70813 47860 71000 47918
rect 70813 47814 70824 47860
rect 70870 47814 70928 47860
rect 70974 47814 71000 47860
rect 70813 47756 71000 47814
rect 70813 47710 70824 47756
rect 70870 47710 70928 47756
rect 70974 47710 71000 47756
rect 70813 47652 71000 47710
rect 70813 47606 70824 47652
rect 70870 47606 70928 47652
rect 70974 47606 71000 47652
rect 70813 47548 71000 47606
rect 70813 47502 70824 47548
rect 70870 47502 70928 47548
rect 70974 47502 71000 47548
rect 70813 47444 71000 47502
rect 70813 47398 70824 47444
rect 70870 47398 70928 47444
rect 70974 47398 71000 47444
rect 70813 47340 71000 47398
rect 70813 47294 70824 47340
rect 70870 47294 70928 47340
rect 70974 47294 71000 47340
rect 70813 47236 71000 47294
rect 70813 47190 70824 47236
rect 70870 47190 70928 47236
rect 70974 47190 71000 47236
rect 70813 47132 71000 47190
rect 70813 47086 70824 47132
rect 70870 47086 70928 47132
rect 70974 47086 71000 47132
rect 70813 47028 71000 47086
rect 70813 46982 70824 47028
rect 70870 46982 70928 47028
rect 70974 46982 71000 47028
rect 70813 46924 71000 46982
rect 70813 46878 70824 46924
rect 70870 46878 70928 46924
rect 70974 46878 71000 46924
rect 70813 46820 71000 46878
rect 70813 46774 70824 46820
rect 70870 46774 70928 46820
rect 70974 46774 71000 46820
rect 70813 46716 71000 46774
rect 70813 46670 70824 46716
rect 70870 46670 70928 46716
rect 70974 46670 71000 46716
rect 70813 46612 71000 46670
rect 70813 46566 70824 46612
rect 70870 46566 70928 46612
rect 70974 46566 71000 46612
rect 70813 46508 71000 46566
rect 70813 46462 70824 46508
rect 70870 46462 70928 46508
rect 70974 46462 71000 46508
rect 70813 46404 71000 46462
rect 70813 46358 70824 46404
rect 70870 46358 70928 46404
rect 70974 46358 71000 46404
rect 70813 46300 71000 46358
rect 70813 46254 70824 46300
rect 70870 46254 70928 46300
rect 70974 46254 71000 46300
rect 70813 46196 71000 46254
rect 70813 46150 70824 46196
rect 70870 46150 70928 46196
rect 70974 46150 71000 46196
rect 70813 46092 71000 46150
rect 70813 46046 70824 46092
rect 70870 46046 70928 46092
rect 70974 46046 71000 46092
rect 70813 45988 71000 46046
rect 70813 45942 70824 45988
rect 70870 45942 70928 45988
rect 70974 45942 71000 45988
rect 70813 45884 71000 45942
rect 70813 45838 70824 45884
rect 70870 45838 70928 45884
rect 70974 45838 71000 45884
rect 70813 45780 71000 45838
rect 70813 45734 70824 45780
rect 70870 45734 70928 45780
rect 70974 45734 71000 45780
rect 70813 45676 71000 45734
rect 70813 45630 70824 45676
rect 70870 45630 70928 45676
rect 70974 45630 71000 45676
rect 70813 45572 71000 45630
rect 70813 45526 70824 45572
rect 70870 45526 70928 45572
rect 70974 45526 71000 45572
rect 70813 45468 71000 45526
rect 70813 45422 70824 45468
rect 70870 45422 70928 45468
rect 70974 45422 71000 45468
rect 70813 45364 71000 45422
rect 70813 45318 70824 45364
rect 70870 45318 70928 45364
rect 70974 45318 71000 45364
rect 70813 45260 71000 45318
rect 70813 45214 70824 45260
rect 70870 45214 70928 45260
rect 70974 45214 71000 45260
rect 70813 45156 71000 45214
rect 70813 45110 70824 45156
rect 70870 45110 70928 45156
rect 70974 45110 71000 45156
rect 70813 45052 71000 45110
rect 70813 45006 70824 45052
rect 70870 45006 70928 45052
rect 70974 45006 71000 45052
rect 70813 44948 71000 45006
tri 13108 44703 13253 44848 ne
rect 13253 44828 13280 44848
tri 13280 44828 13372 44920 sw
rect 70813 44902 70824 44948
rect 70870 44902 70928 44948
rect 70974 44902 71000 44948
rect 70813 44844 71000 44902
rect 13253 44824 13372 44828
rect 13253 44778 13254 44824
rect 13300 44778 13372 44824
rect 13253 44703 13372 44778
tri 13372 44703 13497 44828 sw
rect 70813 44798 70824 44844
rect 70870 44798 70928 44844
rect 70974 44798 71000 44844
rect 70813 44740 71000 44798
tri 13253 44571 13385 44703 ne
rect 13385 44692 13497 44703
rect 13385 44646 13386 44692
rect 13432 44646 13497 44692
rect 13385 44584 13497 44646
tri 13497 44584 13616 44703 sw
rect 70813 44694 70824 44740
rect 70870 44694 70928 44740
rect 70974 44694 71000 44740
rect 70813 44636 71000 44694
rect 70813 44590 70824 44636
rect 70870 44590 70928 44636
rect 70974 44590 71000 44636
rect 13385 44571 13616 44584
tri 13385 44439 13517 44571 ne
rect 13517 44560 13616 44571
rect 13517 44514 13518 44560
rect 13564 44514 13616 44560
rect 13517 44439 13616 44514
tri 13616 44439 13761 44584 sw
rect 70813 44532 71000 44590
rect 70813 44486 70824 44532
rect 70870 44486 70928 44532
rect 70974 44486 71000 44532
tri 13517 44307 13649 44439 ne
rect 13649 44428 13761 44439
rect 13649 44382 13650 44428
rect 13696 44382 13761 44428
rect 13649 44340 13761 44382
tri 13761 44340 13860 44439 sw
rect 70813 44428 71000 44486
rect 70813 44382 70824 44428
rect 70870 44382 70928 44428
rect 70974 44382 71000 44428
rect 13649 44307 13860 44340
tri 13649 44175 13781 44307 ne
rect 13781 44296 13860 44307
rect 13781 44250 13782 44296
rect 13828 44250 13860 44296
rect 13781 44175 13860 44250
tri 13860 44175 14025 44340 sw
rect 70813 44324 71000 44382
rect 70813 44278 70824 44324
rect 70870 44278 70928 44324
rect 70974 44278 71000 44324
rect 70813 44220 71000 44278
tri 13781 44043 13913 44175 ne
rect 13913 44164 14025 44175
rect 13913 44118 13914 44164
rect 13960 44118 14025 44164
rect 13913 44096 14025 44118
tri 14025 44096 14104 44175 sw
rect 70813 44174 70824 44220
rect 70870 44174 70928 44220
rect 70974 44174 71000 44220
rect 70813 44116 71000 44174
rect 13913 44043 14104 44096
tri 13913 43911 14045 44043 ne
rect 14045 44032 14104 44043
rect 14045 43986 14046 44032
rect 14092 43986 14104 44032
rect 14045 43911 14104 43986
tri 14104 43911 14289 44096 sw
rect 70813 44070 70824 44116
rect 70870 44070 70928 44116
rect 70974 44070 71000 44116
rect 70813 44012 71000 44070
rect 70813 43966 70824 44012
rect 70870 43966 70928 44012
rect 70974 43966 71000 44012
tri 14045 43779 14177 43911 ne
rect 14177 43900 14289 43911
rect 14177 43854 14178 43900
rect 14224 43854 14289 43900
rect 14177 43779 14289 43854
tri 14289 43779 14421 43911 sw
rect 70813 43908 71000 43966
rect 70813 43862 70824 43908
rect 70870 43862 70928 43908
rect 70974 43862 71000 43908
rect 70813 43804 71000 43862
tri 14177 43647 14309 43779 ne
rect 14309 43768 14421 43779
rect 14309 43722 14310 43768
rect 14356 43722 14421 43768
rect 14309 43647 14421 43722
tri 14421 43647 14553 43779 sw
rect 70813 43758 70824 43804
rect 70870 43758 70928 43804
rect 70974 43758 71000 43804
rect 70813 43700 71000 43758
rect 70813 43654 70824 43700
rect 70870 43654 70928 43700
rect 70974 43654 71000 43700
tri 14309 43515 14441 43647 ne
rect 14441 43636 14553 43647
rect 14441 43590 14442 43636
rect 14488 43590 14553 43636
rect 14441 43515 14553 43590
tri 14553 43515 14685 43647 sw
rect 70813 43596 71000 43654
rect 70813 43550 70824 43596
rect 70870 43550 70928 43596
rect 70974 43550 71000 43596
tri 14441 43383 14573 43515 ne
rect 14573 43504 14685 43515
rect 14573 43458 14574 43504
rect 14620 43458 14685 43504
rect 14573 43383 14685 43458
tri 14685 43383 14817 43515 sw
rect 70813 43492 71000 43550
rect 70813 43446 70824 43492
rect 70870 43446 70928 43492
rect 70974 43446 71000 43492
rect 70813 43388 71000 43446
tri 14573 43251 14705 43383 ne
rect 14705 43372 14817 43383
rect 14705 43326 14706 43372
rect 14752 43326 14817 43372
rect 14705 43251 14817 43326
tri 14817 43251 14949 43383 sw
rect 70813 43342 70824 43388
rect 70870 43342 70928 43388
rect 70974 43342 71000 43388
rect 70813 43284 71000 43342
tri 14705 43119 14837 43251 ne
rect 14837 43240 14949 43251
rect 14837 43194 14838 43240
rect 14884 43194 14949 43240
rect 14837 43120 14949 43194
tri 14949 43120 15080 43251 sw
rect 70813 43238 70824 43284
rect 70870 43238 70928 43284
rect 70974 43238 71000 43284
rect 70813 43180 71000 43238
rect 70813 43134 70824 43180
rect 70870 43134 70928 43180
rect 70974 43134 71000 43180
rect 14837 43119 15080 43120
tri 14837 42987 14969 43119 ne
rect 14969 43108 15080 43119
rect 14969 43062 14970 43108
rect 15016 43062 15080 43108
rect 14969 42987 15080 43062
tri 15080 42987 15213 43120 sw
rect 70813 43076 71000 43134
rect 70813 43030 70824 43076
rect 70870 43030 70928 43076
rect 70974 43030 71000 43076
tri 14969 42855 15101 42987 ne
rect 15101 42976 15213 42987
rect 15101 42930 15102 42976
rect 15148 42930 15213 42976
rect 15101 42876 15213 42930
tri 15213 42876 15324 42987 sw
rect 70813 42972 71000 43030
rect 70813 42926 70824 42972
rect 70870 42926 70928 42972
rect 70974 42926 71000 42972
rect 15101 42855 15324 42876
tri 15101 42723 15233 42855 ne
rect 15233 42844 15324 42855
rect 15233 42798 15234 42844
rect 15280 42798 15324 42844
rect 15233 42723 15324 42798
tri 15324 42723 15477 42876 sw
rect 70813 42868 71000 42926
rect 70813 42822 70824 42868
rect 70870 42822 70928 42868
rect 70974 42822 71000 42868
rect 70813 42764 71000 42822
tri 15233 42591 15365 42723 ne
rect 15365 42712 15477 42723
rect 15365 42666 15366 42712
rect 15412 42666 15477 42712
rect 15365 42632 15477 42666
tri 15477 42632 15568 42723 sw
rect 70813 42718 70824 42764
rect 70870 42718 70928 42764
rect 70974 42718 71000 42764
rect 70813 42660 71000 42718
rect 15365 42591 15568 42632
tri 15365 42459 15497 42591 ne
rect 15497 42580 15568 42591
rect 15497 42534 15498 42580
rect 15544 42534 15568 42580
rect 15497 42459 15568 42534
tri 15568 42459 15741 42632 sw
rect 70813 42614 70824 42660
rect 70870 42614 70928 42660
rect 70974 42614 71000 42660
rect 70813 42556 71000 42614
rect 70813 42510 70824 42556
rect 70870 42510 70928 42556
rect 70974 42510 71000 42556
tri 15497 42327 15629 42459 ne
rect 15629 42448 15741 42459
rect 15629 42402 15630 42448
rect 15676 42402 15741 42448
rect 15629 42327 15741 42402
tri 15741 42327 15873 42459 sw
rect 70813 42452 71000 42510
rect 70813 42406 70824 42452
rect 70870 42406 70928 42452
rect 70974 42406 71000 42452
rect 70813 42348 71000 42406
tri 15629 42195 15761 42327 ne
rect 15761 42316 15873 42327
rect 15761 42270 15762 42316
rect 15808 42270 15873 42316
rect 15761 42195 15873 42270
tri 15873 42195 16005 42327 sw
rect 70813 42302 70824 42348
rect 70870 42302 70928 42348
rect 70974 42302 71000 42348
rect 70813 42244 71000 42302
rect 70813 42198 70824 42244
rect 70870 42198 70928 42244
rect 70974 42198 71000 42244
tri 15761 42063 15893 42195 ne
rect 15893 42184 16005 42195
rect 15893 42138 15894 42184
rect 15940 42138 16005 42184
rect 15893 42063 16005 42138
tri 16005 42063 16137 42195 sw
rect 70813 42140 71000 42198
rect 70813 42094 70824 42140
rect 70870 42094 70928 42140
rect 70974 42094 71000 42140
tri 15893 41931 16025 42063 ne
rect 16025 42052 16137 42063
rect 16025 42006 16026 42052
rect 16072 42006 16137 42052
rect 16025 41931 16137 42006
tri 16137 41931 16269 42063 sw
rect 70813 42036 71000 42094
rect 70813 41990 70824 42036
rect 70870 41990 70928 42036
rect 70974 41990 71000 42036
rect 70813 41932 71000 41990
tri 16025 41799 16157 41931 ne
rect 16157 41920 16269 41931
rect 16157 41874 16158 41920
rect 16204 41874 16269 41920
rect 16157 41799 16269 41874
tri 16269 41799 16401 41931 sw
rect 70813 41886 70824 41932
rect 70870 41886 70928 41932
rect 70974 41886 71000 41932
rect 70813 41828 71000 41886
tri 16157 41667 16289 41799 ne
rect 16289 41788 16401 41799
rect 16289 41742 16290 41788
rect 16336 41742 16401 41788
rect 16289 41667 16401 41742
tri 16289 41599 16357 41667 ne
rect 16357 41656 16401 41667
tri 16401 41656 16544 41799 sw
rect 70813 41782 70824 41828
rect 70870 41782 70928 41828
rect 70974 41782 71000 41828
rect 70813 41724 71000 41782
rect 70813 41678 70824 41724
rect 70870 41678 70928 41724
rect 70974 41678 71000 41724
rect 16357 41610 16422 41656
rect 16468 41610 16544 41656
rect 16357 41599 16544 41610
tri 16357 41412 16544 41599 ne
tri 16544 41535 16665 41656 sw
rect 70813 41620 71000 41678
rect 70813 41574 70824 41620
rect 70870 41574 70928 41620
rect 70974 41574 71000 41620
rect 16544 41524 16665 41535
rect 16544 41478 16554 41524
rect 16600 41478 16665 41524
rect 16544 41412 16665 41478
tri 16665 41412 16788 41535 sw
rect 70813 41516 71000 41574
rect 70813 41470 70824 41516
rect 70870 41470 70928 41516
rect 70974 41470 71000 41516
rect 70813 41412 71000 41470
tri 16544 41271 16685 41412 ne
rect 16685 41392 16788 41412
rect 16685 41346 16686 41392
rect 16732 41346 16788 41392
rect 16685 41271 16788 41346
tri 16788 41271 16929 41412 sw
rect 70813 41366 70824 41412
rect 70870 41366 70928 41412
rect 70974 41366 71000 41412
rect 70813 41308 71000 41366
tri 16685 41139 16817 41271 ne
rect 16817 41260 16929 41271
rect 16817 41214 16818 41260
rect 16864 41214 16929 41260
rect 16817 41168 16929 41214
tri 16929 41168 17032 41271 sw
rect 70813 41262 70824 41308
rect 70870 41262 70928 41308
rect 70974 41262 71000 41308
rect 70813 41204 71000 41262
rect 16817 41139 17032 41168
tri 16817 41007 16949 41139 ne
rect 16949 41128 17032 41139
rect 16949 41082 16950 41128
rect 16996 41082 17032 41128
rect 16949 41007 17032 41082
tri 17032 41007 17193 41168 sw
rect 70813 41158 70824 41204
rect 70870 41158 70928 41204
rect 70974 41158 71000 41204
rect 70813 41100 71000 41158
rect 70813 41054 70824 41100
rect 70870 41054 70928 41100
rect 70974 41054 71000 41100
tri 16949 40875 17081 41007 ne
rect 17081 40996 17193 41007
rect 17081 40950 17082 40996
rect 17128 40950 17193 40996
rect 17081 40924 17193 40950
tri 17193 40924 17276 41007 sw
rect 70813 40996 71000 41054
rect 70813 40950 70824 40996
rect 70870 40950 70928 40996
rect 70974 40950 71000 40996
rect 17081 40875 17276 40924
tri 17081 40743 17213 40875 ne
rect 17213 40864 17276 40875
rect 17213 40818 17214 40864
rect 17260 40818 17276 40864
rect 17213 40743 17276 40818
tri 17276 40743 17457 40924 sw
rect 70813 40892 71000 40950
rect 70813 40846 70824 40892
rect 70870 40846 70928 40892
rect 70974 40846 71000 40892
rect 70813 40788 71000 40846
tri 17213 40611 17345 40743 ne
rect 17345 40732 17457 40743
rect 17345 40686 17346 40732
rect 17392 40686 17457 40732
rect 17345 40611 17457 40686
tri 17457 40611 17589 40743 sw
rect 70813 40742 70824 40788
rect 70870 40742 70928 40788
rect 70974 40742 71000 40788
rect 70813 40684 71000 40742
rect 70813 40638 70824 40684
rect 70870 40638 70928 40684
rect 70974 40638 71000 40684
tri 17345 40479 17477 40611 ne
rect 17477 40600 17589 40611
rect 17477 40554 17478 40600
rect 17524 40554 17589 40600
rect 17477 40479 17589 40554
tri 17589 40479 17721 40611 sw
rect 70813 40580 71000 40638
rect 70813 40534 70824 40580
rect 70870 40534 70928 40580
rect 70974 40534 71000 40580
tri 17477 40347 17609 40479 ne
rect 17609 40468 17721 40479
rect 17609 40422 17610 40468
rect 17656 40422 17721 40468
rect 17609 40347 17721 40422
tri 17721 40347 17853 40479 sw
rect 70813 40476 71000 40534
rect 70813 40430 70824 40476
rect 70870 40430 70928 40476
rect 70974 40430 71000 40476
rect 70813 40372 71000 40430
tri 17609 40215 17741 40347 ne
rect 17741 40336 17853 40347
rect 17741 40290 17742 40336
rect 17788 40290 17853 40336
rect 17741 40215 17853 40290
tri 17853 40215 17985 40347 sw
rect 70813 40326 70824 40372
rect 70870 40326 70928 40372
rect 70974 40326 71000 40372
rect 70813 40268 71000 40326
rect 70813 40222 70824 40268
rect 70870 40222 70928 40268
rect 70974 40222 71000 40268
tri 17741 40083 17873 40215 ne
rect 17873 40204 17985 40215
rect 17873 40158 17874 40204
rect 17920 40158 17985 40204
rect 17873 40083 17985 40158
tri 17985 40083 18117 40215 sw
rect 70813 40164 71000 40222
rect 70813 40118 70824 40164
rect 70870 40118 70928 40164
rect 70974 40118 71000 40164
tri 17873 39951 18005 40083 ne
rect 18005 40072 18117 40083
rect 18005 40026 18006 40072
rect 18052 40026 18117 40072
rect 18005 39951 18117 40026
tri 18005 39883 18073 39951 ne
rect 18073 39948 18117 39951
tri 18117 39948 18252 40083 sw
rect 70813 40060 71000 40118
rect 70813 40014 70824 40060
rect 70870 40014 70928 40060
rect 70974 40014 71000 40060
rect 70813 39956 71000 40014
rect 18073 39940 18252 39948
rect 18073 39894 18138 39940
rect 18184 39894 18252 39940
rect 18073 39883 18252 39894
tri 18073 39704 18252 39883 ne
tri 18252 39819 18381 39948 sw
rect 70813 39910 70824 39956
rect 70870 39910 70928 39956
rect 70974 39910 71000 39956
rect 70813 39852 71000 39910
rect 18252 39808 18381 39819
rect 18252 39762 18270 39808
rect 18316 39762 18381 39808
rect 18252 39704 18381 39762
tri 18381 39704 18496 39819 sw
rect 70813 39806 70824 39852
rect 70870 39806 70928 39852
rect 70974 39806 71000 39852
rect 70813 39748 71000 39806
tri 18252 39555 18401 39704 ne
rect 18401 39676 18496 39704
rect 18401 39630 18402 39676
rect 18448 39630 18496 39676
rect 18401 39555 18496 39630
tri 18496 39555 18645 39704 sw
rect 70813 39702 70824 39748
rect 70870 39702 70928 39748
rect 70974 39702 71000 39748
rect 70813 39644 71000 39702
rect 70813 39598 70824 39644
rect 70870 39598 70928 39644
rect 70974 39598 71000 39644
tri 18401 39423 18533 39555 ne
rect 18533 39544 18645 39555
rect 18533 39498 18534 39544
rect 18580 39498 18645 39544
rect 18533 39460 18645 39498
tri 18645 39460 18740 39555 sw
rect 70813 39540 71000 39598
rect 70813 39494 70824 39540
rect 70870 39494 70928 39540
rect 70974 39494 71000 39540
rect 18533 39423 18740 39460
tri 18533 39291 18665 39423 ne
rect 18665 39412 18740 39423
rect 18665 39366 18666 39412
rect 18712 39366 18740 39412
rect 18665 39291 18740 39366
tri 18740 39291 18909 39460 sw
rect 70813 39436 71000 39494
rect 70813 39390 70824 39436
rect 70870 39390 70928 39436
rect 70974 39390 71000 39436
rect 70813 39332 71000 39390
tri 18665 39159 18797 39291 ne
rect 18797 39280 18909 39291
rect 18797 39234 18798 39280
rect 18844 39234 18909 39280
rect 18797 39159 18909 39234
tri 18909 39159 19041 39291 sw
rect 70813 39286 70824 39332
rect 70870 39286 70928 39332
rect 70974 39286 71000 39332
rect 70813 39228 71000 39286
rect 70813 39182 70824 39228
rect 70870 39182 70928 39228
rect 70974 39182 71000 39228
tri 18797 39027 18929 39159 ne
rect 18929 39148 19041 39159
rect 18929 39102 18930 39148
rect 18976 39102 19041 39148
rect 18929 39027 19041 39102
tri 19041 39027 19173 39159 sw
rect 70813 39124 71000 39182
rect 70813 39078 70824 39124
rect 70870 39078 70928 39124
rect 70974 39078 71000 39124
tri 18929 38895 19061 39027 ne
rect 19061 39016 19173 39027
rect 19061 38970 19062 39016
rect 19108 38970 19173 39016
rect 19061 38895 19173 38970
tri 19173 38895 19305 39027 sw
rect 70813 39020 71000 39078
rect 70813 38974 70824 39020
rect 70870 38974 70928 39020
rect 70974 38974 71000 39020
rect 70813 38916 71000 38974
tri 19061 38763 19193 38895 ne
rect 19193 38884 19305 38895
rect 19193 38838 19194 38884
rect 19240 38838 19305 38884
rect 19193 38763 19305 38838
tri 19305 38763 19437 38895 sw
rect 70813 38870 70824 38916
rect 70870 38870 70928 38916
rect 70974 38870 71000 38916
rect 70813 38812 71000 38870
rect 70813 38766 70824 38812
rect 70870 38766 70928 38812
rect 70974 38766 71000 38812
tri 19193 38631 19325 38763 ne
rect 19325 38752 19437 38763
rect 19325 38706 19326 38752
rect 19372 38706 19437 38752
rect 19325 38631 19437 38706
tri 19437 38631 19569 38763 sw
rect 70813 38708 71000 38766
rect 70813 38662 70824 38708
rect 70870 38662 70928 38708
rect 70974 38662 71000 38708
tri 19325 38499 19457 38631 ne
rect 19457 38620 19569 38631
rect 19457 38574 19458 38620
rect 19504 38574 19569 38620
rect 19457 38499 19569 38574
tri 19569 38499 19701 38631 sw
rect 70813 38604 71000 38662
rect 70813 38558 70824 38604
rect 70870 38558 70928 38604
rect 70974 38558 71000 38604
rect 70813 38500 71000 38558
tri 19457 38367 19589 38499 ne
rect 19589 38488 19701 38499
rect 19589 38442 19590 38488
rect 19636 38442 19701 38488
rect 19589 38367 19701 38442
tri 19701 38367 19833 38499 sw
rect 70813 38454 70824 38500
rect 70870 38454 70928 38500
rect 70974 38454 71000 38500
rect 70813 38396 71000 38454
tri 19589 38235 19721 38367 ne
rect 19721 38356 19833 38367
rect 19721 38310 19722 38356
rect 19768 38310 19833 38356
rect 19721 38240 19833 38310
tri 19833 38240 19960 38367 sw
rect 70813 38350 70824 38396
rect 70870 38350 70928 38396
rect 70974 38350 71000 38396
rect 70813 38292 71000 38350
rect 70813 38246 70824 38292
rect 70870 38246 70928 38292
rect 70974 38246 71000 38292
rect 19721 38235 19960 38240
tri 19721 38103 19853 38235 ne
rect 19853 38224 19960 38235
rect 19853 38178 19854 38224
rect 19900 38178 19960 38224
rect 19853 38103 19960 38178
tri 19960 38103 20097 38240 sw
rect 70813 38188 71000 38246
rect 70813 38142 70824 38188
rect 70870 38142 70928 38188
rect 70974 38142 71000 38188
tri 19853 37971 19985 38103 ne
rect 19985 38092 20097 38103
rect 19985 38046 19986 38092
rect 20032 38046 20097 38092
rect 19985 37996 20097 38046
tri 20097 37996 20204 38103 sw
rect 70813 38084 71000 38142
rect 70813 38038 70824 38084
rect 70870 38038 70928 38084
rect 70974 38038 71000 38084
rect 19985 37971 20204 37996
tri 19985 37839 20117 37971 ne
rect 20117 37960 20204 37971
rect 20117 37914 20118 37960
rect 20164 37914 20204 37960
rect 20117 37839 20204 37914
tri 20204 37839 20361 37996 sw
rect 70813 37980 71000 38038
rect 70813 37934 70824 37980
rect 70870 37934 70928 37980
rect 70974 37934 71000 37980
rect 70813 37876 71000 37934
tri 20117 37707 20249 37839 ne
rect 20249 37828 20361 37839
rect 20249 37782 20250 37828
rect 20296 37782 20361 37828
rect 20249 37752 20361 37782
tri 20361 37752 20448 37839 sw
rect 70813 37830 70824 37876
rect 70870 37830 70928 37876
rect 70974 37830 71000 37876
rect 70813 37772 71000 37830
rect 20249 37707 20448 37752
tri 20249 37575 20381 37707 ne
rect 20381 37696 20448 37707
rect 20381 37650 20382 37696
rect 20428 37650 20448 37696
rect 20381 37575 20448 37650
tri 20448 37575 20625 37752 sw
rect 70813 37726 70824 37772
rect 70870 37726 70928 37772
rect 70974 37726 71000 37772
rect 70813 37668 71000 37726
rect 70813 37622 70824 37668
rect 70870 37622 70928 37668
rect 70974 37622 71000 37668
tri 20381 37443 20513 37575 ne
rect 20513 37564 20625 37575
rect 20513 37518 20514 37564
rect 20560 37518 20625 37564
rect 20513 37443 20625 37518
tri 20625 37443 20757 37575 sw
rect 70813 37564 71000 37622
rect 70813 37518 70824 37564
rect 70870 37518 70928 37564
rect 70974 37518 71000 37564
rect 70813 37460 71000 37518
tri 20513 37311 20645 37443 ne
rect 20645 37432 20757 37443
rect 20645 37386 20646 37432
rect 20692 37386 20757 37432
rect 20645 37311 20757 37386
tri 20757 37311 20889 37443 sw
rect 70813 37414 70824 37460
rect 70870 37414 70928 37460
rect 70974 37414 71000 37460
rect 70813 37356 71000 37414
tri 20645 37179 20777 37311 ne
rect 20777 37300 20889 37311
rect 20777 37254 20778 37300
rect 20824 37254 20889 37300
rect 20777 37179 20889 37254
tri 20889 37179 21021 37311 sw
rect 70813 37310 70824 37356
rect 70870 37310 70928 37356
rect 70974 37310 71000 37356
rect 70813 37252 71000 37310
rect 70813 37206 70824 37252
rect 70870 37206 70928 37252
rect 70974 37206 71000 37252
tri 20777 37047 20909 37179 ne
rect 20909 37168 21021 37179
rect 20909 37122 20910 37168
rect 20956 37122 21021 37168
rect 20909 37047 21021 37122
tri 21021 37047 21153 37179 sw
rect 70813 37148 71000 37206
rect 70813 37102 70824 37148
rect 70870 37102 70928 37148
rect 70974 37102 71000 37148
tri 20909 36915 21041 37047 ne
rect 21041 37036 21153 37047
rect 21041 36990 21042 37036
rect 21088 36990 21153 37036
rect 21041 36915 21153 36990
tri 21153 36915 21285 37047 sw
rect 70813 37044 71000 37102
rect 70813 36998 70824 37044
rect 70870 36998 70928 37044
rect 70974 36998 71000 37044
rect 70813 36940 71000 36998
tri 21041 36783 21173 36915 ne
rect 21173 36904 21285 36915
rect 21173 36858 21174 36904
rect 21220 36858 21285 36904
rect 21173 36783 21285 36858
tri 21173 36715 21241 36783 ne
rect 21241 36776 21285 36783
tri 21285 36776 21424 36915 sw
rect 70813 36894 70824 36940
rect 70870 36894 70928 36940
rect 70974 36894 71000 36940
rect 70813 36836 71000 36894
rect 70813 36790 70824 36836
rect 70870 36790 70928 36836
rect 70974 36790 71000 36836
rect 21241 36772 21424 36776
rect 21241 36726 21306 36772
rect 21352 36726 21424 36772
rect 21241 36715 21424 36726
tri 21241 36532 21424 36715 ne
tri 21424 36651 21549 36776 sw
rect 70813 36732 71000 36790
rect 70813 36686 70824 36732
rect 70870 36686 70928 36732
rect 70974 36686 71000 36732
rect 21424 36640 21549 36651
rect 21424 36594 21438 36640
rect 21484 36594 21549 36640
rect 21424 36532 21549 36594
tri 21549 36532 21668 36651 sw
rect 70813 36628 71000 36686
rect 70813 36582 70824 36628
rect 70870 36582 70928 36628
rect 70974 36582 71000 36628
tri 21424 36387 21569 36532 ne
rect 21569 36508 21668 36532
rect 21569 36462 21570 36508
rect 21616 36462 21668 36508
rect 21569 36387 21668 36462
tri 21668 36387 21813 36532 sw
rect 70813 36524 71000 36582
rect 70813 36478 70824 36524
rect 70870 36478 70928 36524
rect 70974 36478 71000 36524
rect 70813 36420 71000 36478
tri 21569 36255 21701 36387 ne
rect 21701 36376 21813 36387
rect 21701 36330 21702 36376
rect 21748 36330 21813 36376
rect 21701 36288 21813 36330
tri 21813 36288 21912 36387 sw
rect 70813 36374 70824 36420
rect 70870 36374 70928 36420
rect 70974 36374 71000 36420
rect 70813 36316 71000 36374
rect 21701 36255 21912 36288
tri 21701 36123 21833 36255 ne
rect 21833 36244 21912 36255
rect 21833 36198 21834 36244
rect 21880 36198 21912 36244
rect 21833 36123 21912 36198
tri 21912 36123 22077 36288 sw
rect 70813 36270 70824 36316
rect 70870 36270 70928 36316
rect 70974 36270 71000 36316
rect 70813 36212 71000 36270
rect 70813 36166 70824 36212
rect 70870 36166 70928 36212
rect 70974 36166 71000 36212
tri 21833 35991 21965 36123 ne
rect 21965 36112 22077 36123
rect 21965 36066 21966 36112
rect 22012 36066 22077 36112
rect 21965 36044 22077 36066
tri 22077 36044 22156 36123 sw
rect 70813 36108 71000 36166
rect 70813 36062 70824 36108
rect 70870 36062 70928 36108
rect 70974 36062 71000 36108
rect 21965 35991 22156 36044
tri 21965 35859 22097 35991 ne
rect 22097 35980 22156 35991
rect 22097 35934 22098 35980
rect 22144 35934 22156 35980
rect 22097 35859 22156 35934
tri 22156 35859 22341 36044 sw
rect 70813 36004 71000 36062
rect 70813 35958 70824 36004
rect 70870 35958 70928 36004
rect 70974 35958 71000 36004
rect 70813 35900 71000 35958
tri 22097 35727 22229 35859 ne
rect 22229 35848 22341 35859
rect 22229 35802 22230 35848
rect 22276 35802 22341 35848
rect 22229 35727 22341 35802
tri 22341 35727 22473 35859 sw
rect 70813 35854 70824 35900
rect 70870 35854 70928 35900
rect 70974 35854 71000 35900
rect 70813 35796 71000 35854
rect 70813 35750 70824 35796
rect 70870 35750 70928 35796
rect 70974 35750 71000 35796
tri 22229 35595 22361 35727 ne
rect 22361 35716 22473 35727
rect 22361 35670 22362 35716
rect 22408 35670 22473 35716
rect 22361 35595 22473 35670
tri 22473 35595 22605 35727 sw
rect 70813 35692 71000 35750
rect 70813 35646 70824 35692
rect 70870 35646 70928 35692
rect 70974 35646 71000 35692
tri 22361 35463 22493 35595 ne
rect 22493 35584 22605 35595
rect 22493 35538 22494 35584
rect 22540 35538 22605 35584
rect 22493 35463 22605 35538
tri 22605 35463 22737 35595 sw
rect 70813 35588 71000 35646
rect 70813 35542 70824 35588
rect 70870 35542 70928 35588
rect 70974 35542 71000 35588
rect 70813 35484 71000 35542
tri 22493 35331 22625 35463 ne
rect 22625 35452 22737 35463
rect 22625 35406 22626 35452
rect 22672 35406 22737 35452
rect 22625 35331 22737 35406
tri 22737 35331 22869 35463 sw
rect 70813 35438 70824 35484
rect 70870 35438 70928 35484
rect 70974 35438 71000 35484
rect 70813 35380 71000 35438
rect 70813 35334 70824 35380
rect 70870 35334 70928 35380
rect 70974 35334 71000 35380
tri 22625 35199 22757 35331 ne
rect 22757 35320 22869 35331
rect 22757 35274 22758 35320
rect 22804 35274 22869 35320
rect 22757 35199 22869 35274
tri 22869 35199 23001 35331 sw
rect 70813 35276 71000 35334
rect 70813 35230 70824 35276
rect 70870 35230 70928 35276
rect 70974 35230 71000 35276
tri 22757 35067 22889 35199 ne
rect 22889 35188 23001 35199
rect 22889 35142 22890 35188
rect 22936 35142 23001 35188
rect 22889 35068 23001 35142
tri 23001 35068 23132 35199 sw
rect 70813 35172 71000 35230
rect 70813 35126 70824 35172
rect 70870 35126 70928 35172
rect 70974 35126 71000 35172
rect 70813 35068 71000 35126
rect 22889 35067 23132 35068
tri 22889 34935 23021 35067 ne
rect 23021 35056 23132 35067
rect 23021 35010 23022 35056
rect 23068 35010 23132 35056
rect 23021 34935 23132 35010
tri 23132 34935 23265 35068 sw
rect 70813 35022 70824 35068
rect 70870 35022 70928 35068
rect 70974 35022 71000 35068
rect 70813 34964 71000 35022
tri 23021 34803 23153 34935 ne
rect 23153 34924 23265 34935
rect 23153 34878 23154 34924
rect 23200 34878 23265 34924
rect 23153 34824 23265 34878
tri 23265 34824 23376 34935 sw
rect 70813 34918 70824 34964
rect 70870 34918 70928 34964
rect 70974 34918 71000 34964
rect 70813 34860 71000 34918
rect 23153 34803 23376 34824
tri 23153 34671 23285 34803 ne
rect 23285 34792 23376 34803
rect 23285 34746 23286 34792
rect 23332 34746 23376 34792
rect 23285 34671 23376 34746
tri 23376 34671 23529 34824 sw
rect 70813 34814 70824 34860
rect 70870 34814 70928 34860
rect 70974 34814 71000 34860
rect 70813 34756 71000 34814
rect 70813 34710 70824 34756
rect 70870 34710 70928 34756
rect 70974 34710 71000 34756
tri 23285 34539 23417 34671 ne
rect 23417 34660 23529 34671
rect 23417 34614 23418 34660
rect 23464 34614 23529 34660
rect 23417 34580 23529 34614
tri 23529 34580 23620 34671 sw
rect 70813 34652 71000 34710
rect 70813 34606 70824 34652
rect 70870 34606 70928 34652
rect 70974 34606 71000 34652
rect 23417 34539 23620 34580
tri 23417 34407 23549 34539 ne
rect 23549 34528 23620 34539
rect 23549 34482 23550 34528
rect 23596 34482 23620 34528
rect 23549 34407 23620 34482
tri 23620 34407 23793 34580 sw
rect 70813 34548 71000 34606
rect 70813 34502 70824 34548
rect 70870 34502 70928 34548
rect 70974 34502 71000 34548
rect 70813 34444 71000 34502
tri 23549 34275 23681 34407 ne
rect 23681 34396 23793 34407
rect 23681 34350 23682 34396
rect 23728 34350 23793 34396
rect 23681 34275 23793 34350
tri 23793 34275 23925 34407 sw
rect 70813 34398 70824 34444
rect 70870 34398 70928 34444
rect 70974 34398 71000 34444
rect 70813 34340 71000 34398
rect 70813 34294 70824 34340
rect 70870 34294 70928 34340
rect 70974 34294 71000 34340
tri 23681 34143 23813 34275 ne
rect 23813 34264 23925 34275
rect 23813 34218 23814 34264
rect 23860 34218 23925 34264
rect 23813 34143 23925 34218
tri 23925 34143 24057 34275 sw
rect 70813 34236 71000 34294
rect 70813 34190 70824 34236
rect 70870 34190 70928 34236
rect 70974 34190 71000 34236
tri 23813 34011 23945 34143 ne
rect 23945 34132 24057 34143
rect 23945 34086 23946 34132
rect 23992 34086 24057 34132
rect 23945 34011 24057 34086
tri 24057 34011 24189 34143 sw
rect 70813 34132 71000 34190
rect 70813 34086 70824 34132
rect 70870 34086 70928 34132
rect 70974 34086 71000 34132
rect 70813 34028 71000 34086
tri 23945 33879 24077 34011 ne
rect 24077 34000 24189 34011
rect 24077 33954 24078 34000
rect 24124 33954 24189 34000
rect 24077 33879 24189 33954
tri 24189 33879 24321 34011 sw
rect 70813 33982 70824 34028
rect 70870 33982 70928 34028
rect 70974 33982 71000 34028
rect 70813 33924 71000 33982
tri 24077 33747 24209 33879 ne
rect 24209 33868 24321 33879
rect 24209 33822 24210 33868
rect 24256 33822 24321 33868
rect 24209 33747 24321 33822
tri 24321 33747 24453 33879 sw
rect 70813 33878 70824 33924
rect 70870 33878 70928 33924
rect 70974 33878 71000 33924
rect 70813 33820 71000 33878
rect 70813 33774 70824 33820
rect 70870 33774 70928 33820
rect 70974 33774 71000 33820
tri 24209 33615 24341 33747 ne
rect 24341 33736 24453 33747
rect 24341 33690 24342 33736
rect 24388 33690 24453 33736
rect 24341 33615 24453 33690
tri 24341 33547 24409 33615 ne
rect 24409 33604 24453 33615
tri 24453 33604 24596 33747 sw
rect 70813 33716 71000 33774
rect 70813 33670 70824 33716
rect 70870 33670 70928 33716
rect 70974 33670 71000 33716
rect 70813 33612 71000 33670
rect 24409 33558 24474 33604
rect 24520 33558 24596 33604
rect 24409 33547 24596 33558
tri 24409 33360 24596 33547 ne
tri 24596 33483 24717 33604 sw
rect 70813 33566 70824 33612
rect 70870 33566 70928 33612
rect 70974 33566 71000 33612
rect 70813 33508 71000 33566
rect 24596 33472 24717 33483
rect 24596 33426 24606 33472
rect 24652 33426 24717 33472
rect 24596 33360 24717 33426
tri 24717 33360 24840 33483 sw
rect 70813 33462 70824 33508
rect 70870 33462 70928 33508
rect 70974 33462 71000 33508
rect 70813 33404 71000 33462
tri 24596 33219 24737 33360 ne
rect 24737 33340 24840 33360
rect 24737 33294 24738 33340
rect 24784 33294 24840 33340
rect 24737 33219 24840 33294
tri 24840 33219 24981 33360 sw
rect 70813 33358 70824 33404
rect 70870 33358 70928 33404
rect 70974 33358 71000 33404
rect 70813 33300 71000 33358
rect 70813 33254 70824 33300
rect 70870 33254 70928 33300
rect 70974 33254 71000 33300
tri 24737 33087 24869 33219 ne
rect 24869 33208 24981 33219
rect 24869 33162 24870 33208
rect 24916 33162 24981 33208
rect 24869 33116 24981 33162
tri 24981 33116 25084 33219 sw
rect 70813 33196 71000 33254
rect 70813 33150 70824 33196
rect 70870 33150 70928 33196
rect 70974 33150 71000 33196
rect 24869 33087 25084 33116
tri 24869 32955 25001 33087 ne
rect 25001 33076 25084 33087
rect 25001 33030 25002 33076
rect 25048 33030 25084 33076
rect 25001 32955 25084 33030
tri 25084 32955 25245 33116 sw
rect 70813 33092 71000 33150
rect 70813 33046 70824 33092
rect 70870 33046 70928 33092
rect 70974 33046 71000 33092
rect 70813 32988 71000 33046
tri 25001 32823 25133 32955 ne
rect 25133 32944 25245 32955
rect 25133 32898 25134 32944
rect 25180 32898 25245 32944
rect 25133 32872 25245 32898
tri 25245 32872 25328 32955 sw
rect 70813 32942 70824 32988
rect 70870 32942 70928 32988
rect 70974 32942 71000 32988
rect 70813 32884 71000 32942
rect 25133 32823 25328 32872
tri 25133 32691 25265 32823 ne
rect 25265 32812 25328 32823
rect 25265 32766 25266 32812
rect 25312 32766 25328 32812
rect 25265 32691 25328 32766
tri 25328 32691 25509 32872 sw
rect 70813 32838 70824 32884
rect 70870 32838 70928 32884
rect 70974 32838 71000 32884
rect 70813 32780 71000 32838
rect 70813 32734 70824 32780
rect 70870 32734 70928 32780
rect 70974 32734 71000 32780
tri 25265 32559 25397 32691 ne
rect 25397 32680 25509 32691
rect 25397 32634 25398 32680
rect 25444 32634 25509 32680
rect 25397 32559 25509 32634
tri 25509 32559 25641 32691 sw
rect 70813 32676 71000 32734
rect 70813 32630 70824 32676
rect 70870 32630 70928 32676
rect 70974 32630 71000 32676
rect 70813 32572 71000 32630
tri 25397 32427 25529 32559 ne
rect 25529 32548 25641 32559
rect 25529 32502 25530 32548
rect 25576 32502 25641 32548
rect 25529 32427 25641 32502
tri 25641 32427 25773 32559 sw
rect 70813 32526 70824 32572
rect 70870 32526 70928 32572
rect 70974 32526 71000 32572
rect 70813 32468 71000 32526
tri 25529 32295 25661 32427 ne
rect 25661 32416 25773 32427
rect 25661 32370 25662 32416
rect 25708 32370 25773 32416
rect 25661 32295 25773 32370
tri 25773 32295 25905 32427 sw
rect 70813 32422 70824 32468
rect 70870 32422 70928 32468
rect 70974 32422 71000 32468
rect 70813 32364 71000 32422
rect 70813 32318 70824 32364
rect 70870 32318 70928 32364
rect 70974 32318 71000 32364
tri 25661 32163 25793 32295 ne
rect 25793 32284 25905 32295
rect 25793 32238 25794 32284
rect 25840 32238 25905 32284
rect 25793 32163 25905 32238
tri 25905 32163 26037 32295 sw
rect 70813 32260 71000 32318
rect 70813 32214 70824 32260
rect 70870 32214 70928 32260
rect 70974 32214 71000 32260
tri 25793 32031 25925 32163 ne
rect 25925 32152 26037 32163
rect 25925 32106 25926 32152
rect 25972 32106 26037 32152
rect 25925 32031 26037 32106
tri 26037 32031 26169 32163 sw
rect 70813 32156 71000 32214
rect 70813 32110 70824 32156
rect 70870 32110 70928 32156
rect 70974 32110 71000 32156
rect 70813 32052 71000 32110
tri 25925 31899 26057 32031 ne
rect 26057 32020 26169 32031
rect 26057 31974 26058 32020
rect 26104 31974 26169 32020
rect 26057 31899 26169 31974
tri 26057 31831 26125 31899 ne
rect 26125 31896 26169 31899
tri 26169 31896 26304 32031 sw
rect 70813 32006 70824 32052
rect 70870 32006 70928 32052
rect 70974 32006 71000 32052
rect 70813 31948 71000 32006
rect 70813 31902 70824 31948
rect 70870 31902 70928 31948
rect 70974 31902 71000 31948
rect 26125 31888 26304 31896
rect 26125 31842 26190 31888
rect 26236 31842 26304 31888
rect 26125 31831 26304 31842
tri 26125 31652 26304 31831 ne
tri 26304 31767 26433 31896 sw
rect 70813 31844 71000 31902
rect 70813 31798 70824 31844
rect 70870 31798 70928 31844
rect 70974 31798 71000 31844
rect 26304 31756 26433 31767
rect 26304 31710 26322 31756
rect 26368 31710 26433 31756
rect 26304 31652 26433 31710
tri 26433 31652 26548 31767 sw
rect 70813 31740 71000 31798
rect 70813 31694 70824 31740
rect 70870 31694 70928 31740
rect 70974 31694 71000 31740
tri 26304 31503 26453 31652 ne
rect 26453 31624 26548 31652
rect 26453 31578 26454 31624
rect 26500 31578 26548 31624
rect 26453 31503 26548 31578
tri 26548 31503 26697 31652 sw
rect 70813 31636 71000 31694
rect 70813 31590 70824 31636
rect 70870 31590 70928 31636
rect 70974 31590 71000 31636
rect 70813 31532 71000 31590
tri 26453 31371 26585 31503 ne
rect 26585 31492 26697 31503
rect 26585 31446 26586 31492
rect 26632 31446 26697 31492
rect 26585 31408 26697 31446
tri 26697 31408 26792 31503 sw
rect 70813 31486 70824 31532
rect 70870 31486 70928 31532
rect 70974 31486 71000 31532
rect 70813 31428 71000 31486
rect 26585 31371 26792 31408
tri 26585 31239 26717 31371 ne
rect 26717 31360 26792 31371
rect 26717 31314 26718 31360
rect 26764 31314 26792 31360
rect 26717 31239 26792 31314
tri 26792 31239 26961 31408 sw
rect 70813 31382 70824 31428
rect 70870 31382 70928 31428
rect 70974 31382 71000 31428
rect 70813 31324 71000 31382
rect 70813 31278 70824 31324
rect 70870 31278 70928 31324
rect 70974 31278 71000 31324
tri 26717 31107 26849 31239 ne
rect 26849 31228 26961 31239
rect 26849 31182 26850 31228
rect 26896 31182 26961 31228
rect 26849 31107 26961 31182
tri 26961 31107 27093 31239 sw
rect 70813 31220 71000 31278
rect 70813 31174 70824 31220
rect 70870 31174 70928 31220
rect 70974 31174 71000 31220
rect 70813 31116 71000 31174
tri 26849 30975 26981 31107 ne
rect 26981 31096 27093 31107
rect 26981 31050 26982 31096
rect 27028 31050 27093 31096
rect 26981 30975 27093 31050
tri 27093 30975 27225 31107 sw
rect 70813 31070 70824 31116
rect 70870 31070 70928 31116
rect 70974 31070 71000 31116
rect 70813 31012 71000 31070
tri 26981 30843 27113 30975 ne
rect 27113 30964 27225 30975
rect 27113 30918 27114 30964
rect 27160 30918 27225 30964
rect 27113 30843 27225 30918
tri 27225 30843 27357 30975 sw
rect 70813 30966 70824 31012
rect 70870 30966 70928 31012
rect 70974 30966 71000 31012
rect 70813 30908 71000 30966
rect 70813 30862 70824 30908
rect 70870 30862 70928 30908
rect 70974 30862 71000 30908
tri 27113 30711 27245 30843 ne
rect 27245 30832 27357 30843
rect 27245 30786 27246 30832
rect 27292 30786 27357 30832
rect 27245 30711 27357 30786
tri 27357 30711 27489 30843 sw
rect 70813 30804 71000 30862
rect 70813 30758 70824 30804
rect 70870 30758 70928 30804
rect 70974 30758 71000 30804
tri 27245 30579 27377 30711 ne
rect 27377 30700 27489 30711
rect 27377 30654 27378 30700
rect 27424 30654 27489 30700
rect 27377 30579 27489 30654
tri 27489 30579 27621 30711 sw
rect 70813 30700 71000 30758
rect 70813 30654 70824 30700
rect 70870 30654 70928 30700
rect 70974 30654 71000 30700
rect 70813 30596 71000 30654
tri 27377 30447 27509 30579 ne
rect 27509 30568 27621 30579
rect 27509 30522 27510 30568
rect 27556 30522 27621 30568
rect 27509 30447 27621 30522
tri 27621 30447 27753 30579 sw
rect 70813 30550 70824 30596
rect 70870 30550 70928 30596
rect 70974 30550 71000 30596
rect 70813 30492 71000 30550
tri 27509 30315 27641 30447 ne
rect 27641 30436 27753 30447
rect 27641 30390 27642 30436
rect 27688 30390 27753 30436
rect 27641 30315 27753 30390
tri 27753 30315 27885 30447 sw
rect 70813 30446 70824 30492
rect 70870 30446 70928 30492
rect 70974 30446 71000 30492
rect 70813 30388 71000 30446
rect 70813 30342 70824 30388
rect 70870 30342 70928 30388
rect 70974 30342 71000 30388
tri 27641 30183 27773 30315 ne
rect 27773 30304 27885 30315
rect 27773 30258 27774 30304
rect 27820 30258 27885 30304
rect 27773 30188 27885 30258
tri 27885 30188 28012 30315 sw
rect 70813 30284 71000 30342
rect 70813 30238 70824 30284
rect 70870 30238 70928 30284
rect 70974 30238 71000 30284
rect 27773 30183 28012 30188
tri 27773 30051 27905 30183 ne
rect 27905 30172 28012 30183
rect 27905 30126 27906 30172
rect 27952 30126 28012 30172
rect 27905 30051 28012 30126
tri 28012 30051 28149 30188 sw
rect 70813 30180 71000 30238
rect 70813 30134 70824 30180
rect 70870 30134 70928 30180
rect 70974 30134 71000 30180
rect 70813 30076 71000 30134
tri 27905 29919 28037 30051 ne
rect 28037 30040 28149 30051
rect 28037 29994 28038 30040
rect 28084 29994 28149 30040
rect 28037 29944 28149 29994
tri 28149 29944 28256 30051 sw
rect 70813 30030 70824 30076
rect 70870 30030 70928 30076
rect 70974 30030 71000 30076
rect 70813 29972 71000 30030
rect 28037 29919 28256 29944
tri 28037 29787 28169 29919 ne
rect 28169 29908 28256 29919
rect 28169 29862 28170 29908
rect 28216 29862 28256 29908
rect 28169 29787 28256 29862
tri 28256 29787 28413 29944 sw
rect 70813 29926 70824 29972
rect 70870 29926 70928 29972
rect 70974 29926 71000 29972
rect 70813 29868 71000 29926
rect 70813 29822 70824 29868
rect 70870 29822 70928 29868
rect 70974 29822 71000 29868
tri 28169 29655 28301 29787 ne
rect 28301 29776 28413 29787
rect 28301 29730 28302 29776
rect 28348 29730 28413 29776
rect 28301 29700 28413 29730
tri 28413 29700 28500 29787 sw
rect 70813 29764 71000 29822
rect 70813 29718 70824 29764
rect 70870 29718 70928 29764
rect 70974 29718 71000 29764
rect 28301 29655 28500 29700
tri 28301 29523 28433 29655 ne
rect 28433 29644 28500 29655
rect 28433 29598 28434 29644
rect 28480 29598 28500 29644
rect 28433 29523 28500 29598
tri 28500 29523 28677 29700 sw
rect 70813 29660 71000 29718
rect 70813 29614 70824 29660
rect 70870 29614 70928 29660
rect 70974 29614 71000 29660
rect 70813 29556 71000 29614
tri 28433 29391 28565 29523 ne
rect 28565 29512 28677 29523
rect 28565 29466 28566 29512
rect 28612 29466 28677 29512
rect 28565 29391 28677 29466
tri 28677 29391 28809 29523 sw
rect 70813 29510 70824 29556
rect 70870 29510 70928 29556
rect 70974 29510 71000 29556
rect 70813 29452 71000 29510
rect 70813 29406 70824 29452
rect 70870 29406 70928 29452
rect 70974 29406 71000 29452
tri 28565 29259 28697 29391 ne
rect 28697 29380 28809 29391
rect 28697 29334 28698 29380
rect 28744 29334 28809 29380
rect 28697 29259 28809 29334
tri 28809 29259 28941 29391 sw
rect 70813 29348 71000 29406
rect 70813 29302 70824 29348
rect 70870 29302 70928 29348
rect 70974 29302 71000 29348
tri 28697 29127 28829 29259 ne
rect 28829 29248 28941 29259
rect 28829 29202 28830 29248
rect 28876 29202 28941 29248
rect 28829 29127 28941 29202
tri 28941 29127 29073 29259 sw
rect 70813 29244 71000 29302
rect 70813 29198 70824 29244
rect 70870 29198 70928 29244
rect 70974 29198 71000 29244
rect 70813 29140 71000 29198
tri 28829 28995 28961 29127 ne
rect 28961 29116 29073 29127
rect 28961 29070 28962 29116
rect 29008 29070 29073 29116
rect 28961 28995 29073 29070
tri 29073 28995 29205 29127 sw
rect 70813 29094 70824 29140
rect 70870 29094 70928 29140
rect 70974 29094 71000 29140
rect 70813 29036 71000 29094
tri 28961 28863 29093 28995 ne
rect 29093 28984 29205 28995
rect 29093 28938 29094 28984
rect 29140 28938 29205 28984
rect 29093 28863 29205 28938
tri 29205 28863 29337 28995 sw
rect 70813 28990 70824 29036
rect 70870 28990 70928 29036
rect 70974 28990 71000 29036
rect 70813 28932 71000 28990
rect 70813 28886 70824 28932
rect 70870 28886 70928 28932
rect 70974 28886 71000 28932
tri 29093 28731 29225 28863 ne
rect 29225 28852 29337 28863
rect 29225 28806 29226 28852
rect 29272 28806 29337 28852
rect 29225 28731 29337 28806
tri 29225 28663 29293 28731 ne
rect 29293 28724 29337 28731
tri 29337 28724 29476 28863 sw
rect 70813 28828 71000 28886
rect 70813 28782 70824 28828
rect 70870 28782 70928 28828
rect 70974 28782 71000 28828
rect 70813 28724 71000 28782
rect 29293 28720 29476 28724
rect 29293 28674 29358 28720
rect 29404 28674 29476 28720
rect 29293 28663 29476 28674
tri 29293 28480 29476 28663 ne
tri 29476 28599 29601 28724 sw
rect 70813 28678 70824 28724
rect 70870 28678 70928 28724
rect 70974 28678 71000 28724
rect 70813 28620 71000 28678
rect 29476 28588 29601 28599
rect 29476 28542 29490 28588
rect 29536 28542 29601 28588
rect 29476 28480 29601 28542
tri 29601 28480 29720 28599 sw
rect 70813 28574 70824 28620
rect 70870 28574 70928 28620
rect 70974 28574 71000 28620
rect 70813 28516 71000 28574
tri 29476 28335 29621 28480 ne
rect 29621 28456 29720 28480
rect 29621 28410 29622 28456
rect 29668 28410 29720 28456
rect 29621 28335 29720 28410
tri 29720 28335 29865 28480 sw
rect 70813 28470 70824 28516
rect 70870 28470 70928 28516
rect 70974 28470 71000 28516
rect 70813 28412 71000 28470
rect 70813 28366 70824 28412
rect 70870 28366 70928 28412
rect 70974 28366 71000 28412
tri 29621 28203 29753 28335 ne
rect 29753 28324 29865 28335
rect 29753 28278 29754 28324
rect 29800 28278 29865 28324
rect 29753 28236 29865 28278
tri 29865 28236 29964 28335 sw
rect 70813 28308 71000 28366
rect 70813 28262 70824 28308
rect 70870 28262 70928 28308
rect 70974 28262 71000 28308
rect 29753 28203 29964 28236
tri 29753 28071 29885 28203 ne
rect 29885 28192 29964 28203
rect 29885 28146 29886 28192
rect 29932 28146 29964 28192
rect 29885 28071 29964 28146
tri 29964 28071 30129 28236 sw
rect 70813 28204 71000 28262
rect 70813 28158 70824 28204
rect 70870 28158 70928 28204
rect 70974 28158 71000 28204
rect 70813 28100 71000 28158
tri 29885 27939 30017 28071 ne
rect 30017 28060 30129 28071
rect 30017 28014 30018 28060
rect 30064 28014 30129 28060
rect 30017 27992 30129 28014
tri 30129 27992 30208 28071 sw
rect 70813 28054 70824 28100
rect 70870 28054 70928 28100
rect 70974 28054 71000 28100
rect 70813 27996 71000 28054
rect 30017 27939 30208 27992
tri 30017 27807 30149 27939 ne
rect 30149 27928 30208 27939
rect 30149 27882 30150 27928
rect 30196 27882 30208 27928
rect 30149 27807 30208 27882
tri 30208 27807 30393 27992 sw
rect 70813 27950 70824 27996
rect 70870 27950 70928 27996
rect 70974 27950 71000 27996
rect 70813 27892 71000 27950
rect 70813 27846 70824 27892
rect 70870 27846 70928 27892
rect 70974 27846 71000 27892
tri 30149 27675 30281 27807 ne
rect 30281 27796 30393 27807
rect 30281 27750 30282 27796
rect 30328 27750 30393 27796
rect 30281 27675 30393 27750
tri 30393 27675 30525 27807 sw
rect 70813 27788 71000 27846
rect 70813 27742 70824 27788
rect 70870 27742 70928 27788
rect 70974 27742 71000 27788
rect 70813 27684 71000 27742
tri 30281 27543 30413 27675 ne
rect 30413 27664 30525 27675
rect 30413 27618 30414 27664
rect 30460 27618 30525 27664
rect 30413 27543 30525 27618
tri 30525 27543 30657 27675 sw
rect 70813 27638 70824 27684
rect 70870 27638 70928 27684
rect 70974 27638 71000 27684
rect 70813 27580 71000 27638
tri 30413 27411 30545 27543 ne
rect 30545 27532 30657 27543
rect 30545 27486 30546 27532
rect 30592 27486 30657 27532
rect 30545 27411 30657 27486
tri 30657 27411 30789 27543 sw
rect 70813 27534 70824 27580
rect 70870 27534 70928 27580
rect 70974 27534 71000 27580
rect 70813 27476 71000 27534
rect 70813 27430 70824 27476
rect 70870 27430 70928 27476
rect 70974 27430 71000 27476
tri 30545 27279 30677 27411 ne
rect 30677 27400 30789 27411
rect 30677 27354 30678 27400
rect 30724 27354 30789 27400
rect 30677 27279 30789 27354
tri 30789 27279 30921 27411 sw
rect 70813 27372 71000 27430
rect 70813 27326 70824 27372
rect 70870 27326 70928 27372
rect 70974 27326 71000 27372
tri 30677 27147 30809 27279 ne
rect 30809 27268 30921 27279
rect 30809 27222 30810 27268
rect 30856 27222 30921 27268
rect 30809 27147 30921 27222
tri 30921 27147 31053 27279 sw
rect 70813 27268 71000 27326
rect 70813 27222 70824 27268
rect 70870 27222 70928 27268
rect 70974 27222 71000 27268
rect 70813 27164 71000 27222
tri 30809 27015 30941 27147 ne
rect 30941 27136 31053 27147
rect 30941 27090 30942 27136
rect 30988 27090 31053 27136
rect 30941 27016 31053 27090
tri 31053 27016 31184 27147 sw
rect 70813 27118 70824 27164
rect 70870 27118 70928 27164
rect 70974 27118 71000 27164
rect 70813 27060 71000 27118
rect 30941 27015 31184 27016
tri 30941 26883 31073 27015 ne
rect 31073 27004 31184 27015
rect 31073 26958 31074 27004
rect 31120 26958 31184 27004
rect 31073 26883 31184 26958
tri 31184 26883 31317 27016 sw
rect 70813 27014 70824 27060
rect 70870 27014 70928 27060
rect 70974 27014 71000 27060
rect 70813 26956 71000 27014
rect 70813 26910 70824 26956
rect 70870 26910 70928 26956
rect 70974 26910 71000 26956
tri 31073 26751 31205 26883 ne
rect 31205 26872 31317 26883
rect 31205 26826 31206 26872
rect 31252 26826 31317 26872
rect 31205 26772 31317 26826
tri 31317 26772 31428 26883 sw
rect 70813 26852 71000 26910
rect 70813 26806 70824 26852
rect 70870 26806 70928 26852
rect 70974 26806 71000 26852
rect 31205 26751 31428 26772
tri 31205 26619 31337 26751 ne
rect 31337 26740 31428 26751
rect 31337 26694 31338 26740
rect 31384 26694 31428 26740
rect 31337 26619 31428 26694
tri 31428 26619 31581 26772 sw
rect 70813 26748 71000 26806
rect 70813 26702 70824 26748
rect 70870 26702 70928 26748
rect 70974 26702 71000 26748
rect 70813 26644 71000 26702
tri 31337 26487 31469 26619 ne
rect 31469 26608 31581 26619
rect 31469 26562 31470 26608
rect 31516 26562 31581 26608
rect 31469 26528 31581 26562
tri 31581 26528 31672 26619 sw
rect 70813 26598 70824 26644
rect 70870 26598 70928 26644
rect 70974 26598 71000 26644
rect 70813 26540 71000 26598
rect 31469 26487 31672 26528
tri 31469 26355 31601 26487 ne
rect 31601 26476 31672 26487
rect 31601 26430 31602 26476
rect 31648 26430 31672 26476
rect 31601 26355 31672 26430
tri 31672 26355 31845 26528 sw
rect 70813 26494 70824 26540
rect 70870 26494 70928 26540
rect 70974 26494 71000 26540
rect 70813 26436 71000 26494
rect 70813 26390 70824 26436
rect 70870 26390 70928 26436
rect 70974 26390 71000 26436
tri 31601 26223 31733 26355 ne
rect 31733 26344 31845 26355
rect 31733 26298 31734 26344
rect 31780 26298 31845 26344
rect 31733 26223 31845 26298
tri 31845 26223 31977 26355 sw
rect 70813 26332 71000 26390
rect 70813 26286 70824 26332
rect 70870 26286 70928 26332
rect 70974 26286 71000 26332
rect 70813 26228 71000 26286
tri 31733 26091 31865 26223 ne
rect 31865 26212 31977 26223
rect 31865 26166 31866 26212
rect 31912 26166 31977 26212
rect 31865 26091 31977 26166
tri 31977 26091 32109 26223 sw
rect 70813 26182 70824 26228
rect 70870 26182 70928 26228
rect 70974 26182 71000 26228
rect 70813 26124 71000 26182
tri 31865 25959 31997 26091 ne
rect 31997 26080 32109 26091
rect 31997 26034 31998 26080
rect 32044 26034 32109 26080
rect 31997 25959 32109 26034
tri 32109 25959 32241 26091 sw
rect 70813 26078 70824 26124
rect 70870 26078 70928 26124
rect 70974 26078 71000 26124
rect 70813 26020 71000 26078
rect 70813 25974 70824 26020
rect 70870 25974 70928 26020
rect 70974 25974 71000 26020
tri 31997 25827 32129 25959 ne
rect 32129 25948 32241 25959
rect 32129 25902 32130 25948
rect 32176 25902 32241 25948
rect 32129 25827 32241 25902
tri 32241 25827 32373 25959 sw
rect 70813 25916 71000 25974
rect 70813 25870 70824 25916
rect 70870 25870 70928 25916
rect 70974 25870 71000 25916
tri 32129 25695 32261 25827 ne
rect 32261 25816 32373 25827
rect 32261 25770 32262 25816
rect 32308 25770 32373 25816
rect 32261 25695 32373 25770
tri 32373 25695 32505 25827 sw
rect 70813 25812 71000 25870
rect 70813 25766 70824 25812
rect 70870 25766 70928 25812
rect 70974 25766 71000 25812
rect 70813 25708 71000 25766
tri 32261 25563 32393 25695 ne
rect 32393 25684 32505 25695
rect 32393 25638 32394 25684
rect 32440 25638 32505 25684
rect 32393 25563 32505 25638
tri 32393 25495 32461 25563 ne
rect 32461 25552 32505 25563
tri 32505 25552 32648 25695 sw
rect 70813 25662 70824 25708
rect 70870 25662 70928 25708
rect 70974 25662 71000 25708
rect 70813 25604 71000 25662
rect 70813 25558 70824 25604
rect 70870 25558 70928 25604
rect 70974 25558 71000 25604
rect 32461 25506 32526 25552
rect 32572 25506 32648 25552
rect 32461 25495 32648 25506
tri 32461 25308 32648 25495 ne
tri 32648 25431 32769 25552 sw
rect 70813 25500 71000 25558
rect 70813 25454 70824 25500
rect 70870 25454 70928 25500
rect 70974 25454 71000 25500
rect 32648 25420 32769 25431
rect 32648 25374 32658 25420
rect 32704 25374 32769 25420
rect 32648 25308 32769 25374
tri 32769 25308 32892 25431 sw
rect 70813 25396 71000 25454
rect 70813 25350 70824 25396
rect 70870 25350 70928 25396
rect 70974 25350 71000 25396
tri 32648 25167 32789 25308 ne
rect 32789 25288 32892 25308
rect 32789 25242 32790 25288
rect 32836 25242 32892 25288
rect 32789 25167 32892 25242
tri 32892 25167 33033 25308 sw
rect 70813 25292 71000 25350
rect 70813 25246 70824 25292
rect 70870 25246 70928 25292
rect 70974 25246 71000 25292
rect 70813 25188 71000 25246
tri 32789 25035 32921 25167 ne
rect 32921 25156 33033 25167
rect 32921 25110 32922 25156
rect 32968 25110 33033 25156
rect 32921 25064 33033 25110
tri 33033 25064 33136 25167 sw
rect 70813 25142 70824 25188
rect 70870 25142 70928 25188
rect 70974 25142 71000 25188
rect 70813 25084 71000 25142
rect 32921 25035 33136 25064
tri 32921 24903 33053 25035 ne
rect 33053 25024 33136 25035
rect 33053 24978 33054 25024
rect 33100 24978 33136 25024
rect 33053 24903 33136 24978
tri 33136 24903 33297 25064 sw
rect 70813 25038 70824 25084
rect 70870 25038 70928 25084
rect 70974 25038 71000 25084
rect 70813 24980 71000 25038
rect 70813 24934 70824 24980
rect 70870 24934 70928 24980
rect 70974 24934 71000 24980
tri 33053 24771 33185 24903 ne
rect 33185 24892 33297 24903
rect 33185 24846 33186 24892
rect 33232 24846 33297 24892
rect 33185 24820 33297 24846
tri 33297 24820 33380 24903 sw
rect 70813 24876 71000 24934
rect 70813 24830 70824 24876
rect 70870 24830 70928 24876
rect 70974 24830 71000 24876
rect 33185 24771 33380 24820
tri 33185 24639 33317 24771 ne
rect 33317 24760 33380 24771
rect 33317 24714 33318 24760
rect 33364 24714 33380 24760
rect 33317 24639 33380 24714
tri 33380 24639 33561 24820 sw
rect 70813 24772 71000 24830
rect 70813 24726 70824 24772
rect 70870 24726 70928 24772
rect 70974 24726 71000 24772
rect 70813 24668 71000 24726
tri 33317 24507 33449 24639 ne
rect 33449 24628 33561 24639
rect 33449 24582 33450 24628
rect 33496 24582 33561 24628
rect 33449 24507 33561 24582
tri 33561 24507 33693 24639 sw
rect 70813 24622 70824 24668
rect 70870 24622 70928 24668
rect 70974 24622 71000 24668
rect 70813 24564 71000 24622
rect 70813 24518 70824 24564
rect 70870 24518 70928 24564
rect 70974 24518 71000 24564
tri 33449 24375 33581 24507 ne
rect 33581 24496 33693 24507
rect 33581 24450 33582 24496
rect 33628 24450 33693 24496
rect 33581 24375 33693 24450
tri 33693 24375 33825 24507 sw
rect 70813 24460 71000 24518
rect 70813 24414 70824 24460
rect 70870 24414 70928 24460
rect 70974 24414 71000 24460
tri 33581 24243 33713 24375 ne
rect 33713 24364 33825 24375
rect 33713 24318 33714 24364
rect 33760 24318 33825 24364
rect 33713 24243 33825 24318
tri 33825 24243 33957 24375 sw
rect 70813 24356 71000 24414
rect 70813 24310 70824 24356
rect 70870 24310 70928 24356
rect 70974 24310 71000 24356
rect 70813 24252 71000 24310
tri 33713 24111 33845 24243 ne
rect 33845 24232 33957 24243
rect 33845 24186 33846 24232
rect 33892 24186 33957 24232
rect 33845 24111 33957 24186
tri 33957 24111 34089 24243 sw
rect 70813 24206 70824 24252
rect 70870 24206 70928 24252
rect 70974 24206 71000 24252
rect 70813 24148 71000 24206
tri 33845 23979 33977 24111 ne
rect 33977 24100 34089 24111
rect 33977 24054 33978 24100
rect 34024 24054 34089 24100
rect 33977 23979 34089 24054
tri 34089 23979 34221 24111 sw
rect 70813 24102 70824 24148
rect 70870 24102 70928 24148
rect 70974 24102 71000 24148
rect 70813 24044 71000 24102
rect 70813 23998 70824 24044
rect 70870 23998 70928 24044
rect 70974 23998 71000 24044
tri 33977 23847 34109 23979 ne
rect 34109 23968 34221 23979
rect 34109 23922 34110 23968
rect 34156 23922 34221 23968
rect 34109 23847 34221 23922
tri 34109 23779 34177 23847 ne
rect 34177 23844 34221 23847
tri 34221 23844 34356 23979 sw
rect 70813 23940 71000 23998
rect 70813 23894 70824 23940
rect 70870 23894 70928 23940
rect 70974 23894 71000 23940
rect 34177 23836 34356 23844
rect 34177 23790 34242 23836
rect 34288 23790 34356 23836
rect 34177 23779 34356 23790
tri 34177 23600 34356 23779 ne
tri 34356 23715 34485 23844 sw
rect 70813 23836 71000 23894
rect 70813 23790 70824 23836
rect 70870 23790 70928 23836
rect 70974 23790 71000 23836
rect 70813 23732 71000 23790
rect 34356 23704 34485 23715
rect 34356 23658 34374 23704
rect 34420 23658 34485 23704
rect 34356 23600 34485 23658
tri 34485 23600 34600 23715 sw
rect 70813 23686 70824 23732
rect 70870 23686 70928 23732
rect 70974 23686 71000 23732
rect 70813 23628 71000 23686
tri 34356 23451 34505 23600 ne
rect 34505 23572 34600 23600
rect 34505 23526 34506 23572
rect 34552 23526 34600 23572
rect 34505 23451 34600 23526
tri 34600 23451 34749 23600 sw
rect 70813 23582 70824 23628
rect 70870 23582 70928 23628
rect 70974 23582 71000 23628
rect 70813 23524 71000 23582
rect 70813 23478 70824 23524
rect 70870 23478 70928 23524
rect 70974 23478 71000 23524
tri 34505 23319 34637 23451 ne
rect 34637 23440 34749 23451
rect 34637 23394 34638 23440
rect 34684 23394 34749 23440
rect 34637 23356 34749 23394
tri 34749 23356 34844 23451 sw
rect 70813 23420 71000 23478
rect 70813 23374 70824 23420
rect 70870 23374 70928 23420
rect 70974 23374 71000 23420
rect 34637 23319 34844 23356
tri 34637 23187 34769 23319 ne
rect 34769 23308 34844 23319
rect 34769 23262 34770 23308
rect 34816 23262 34844 23308
rect 34769 23187 34844 23262
tri 34844 23187 35013 23356 sw
rect 70813 23316 71000 23374
rect 70813 23270 70824 23316
rect 70870 23270 70928 23316
rect 70974 23270 71000 23316
rect 70813 23212 71000 23270
tri 34769 23055 34901 23187 ne
rect 34901 23176 35013 23187
rect 34901 23130 34902 23176
rect 34948 23130 35013 23176
rect 34901 23055 35013 23130
tri 35013 23055 35145 23187 sw
rect 70813 23166 70824 23212
rect 70870 23166 70928 23212
rect 70974 23166 71000 23212
rect 70813 23108 71000 23166
rect 70813 23062 70824 23108
rect 70870 23062 70928 23108
rect 70974 23062 71000 23108
tri 34901 22923 35033 23055 ne
rect 35033 23044 35145 23055
rect 35033 22998 35034 23044
rect 35080 22998 35145 23044
rect 35033 22923 35145 22998
tri 35145 22923 35277 23055 sw
rect 70813 23004 71000 23062
rect 70813 22958 70824 23004
rect 70870 22958 70928 23004
rect 70974 22958 71000 23004
tri 35033 22791 35165 22923 ne
rect 35165 22912 35277 22923
rect 35165 22866 35166 22912
rect 35212 22866 35277 22912
rect 35165 22791 35277 22866
tri 35277 22791 35409 22923 sw
rect 70813 22900 71000 22958
rect 70813 22854 70824 22900
rect 70870 22854 70928 22900
rect 70974 22854 71000 22900
rect 70813 22796 71000 22854
tri 35165 22659 35297 22791 ne
rect 35297 22780 35409 22791
rect 35297 22734 35298 22780
rect 35344 22734 35409 22780
rect 35297 22659 35409 22734
tri 35409 22659 35541 22791 sw
rect 70813 22750 70824 22796
rect 70870 22750 70928 22796
rect 70974 22750 71000 22796
rect 70813 22692 71000 22750
tri 35297 22527 35429 22659 ne
rect 35429 22648 35541 22659
rect 35429 22602 35430 22648
rect 35476 22602 35541 22648
rect 35429 22527 35541 22602
tri 35541 22527 35673 22659 sw
rect 70813 22646 70824 22692
rect 70870 22646 70928 22692
rect 70974 22646 71000 22692
rect 70813 22588 71000 22646
rect 70813 22542 70824 22588
rect 70870 22542 70928 22588
rect 70974 22542 71000 22588
tri 35429 22395 35561 22527 ne
rect 35561 22516 35673 22527
rect 35561 22470 35562 22516
rect 35608 22470 35673 22516
rect 35561 22395 35673 22470
tri 35673 22395 35805 22527 sw
rect 70813 22484 71000 22542
rect 70813 22438 70824 22484
rect 70870 22438 70928 22484
rect 70974 22438 71000 22484
tri 35561 22263 35693 22395 ne
rect 35693 22384 35805 22395
rect 35693 22338 35694 22384
rect 35740 22338 35805 22384
rect 35693 22263 35805 22338
tri 35805 22263 35937 22395 sw
rect 70813 22380 71000 22438
rect 70813 22334 70824 22380
rect 70870 22334 70928 22380
rect 70974 22334 71000 22380
rect 70813 22276 71000 22334
tri 35693 22131 35825 22263 ne
rect 35825 22252 35937 22263
rect 35825 22206 35826 22252
rect 35872 22206 35937 22252
rect 35825 22136 35937 22206
tri 35937 22136 36064 22263 sw
rect 70813 22230 70824 22276
rect 70870 22230 70928 22276
rect 70974 22230 71000 22276
rect 70813 22172 71000 22230
rect 35825 22131 36064 22136
tri 35825 21999 35957 22131 ne
rect 35957 22120 36064 22131
rect 35957 22074 35958 22120
rect 36004 22074 36064 22120
rect 35957 21999 36064 22074
tri 36064 21999 36201 22136 sw
rect 70813 22126 70824 22172
rect 70870 22126 70928 22172
rect 70974 22126 71000 22172
rect 70813 22068 71000 22126
rect 70813 22022 70824 22068
rect 70870 22022 70928 22068
rect 70974 22022 71000 22068
tri 35957 21867 36089 21999 ne
rect 36089 21988 36201 21999
rect 36089 21942 36090 21988
rect 36136 21942 36201 21988
rect 36089 21892 36201 21942
tri 36201 21892 36308 21999 sw
rect 70813 21964 71000 22022
rect 70813 21918 70824 21964
rect 70870 21918 70928 21964
rect 70974 21918 71000 21964
rect 36089 21867 36308 21892
tri 36089 21735 36221 21867 ne
rect 36221 21856 36308 21867
rect 36221 21810 36222 21856
rect 36268 21810 36308 21856
rect 36221 21735 36308 21810
tri 36308 21735 36465 21892 sw
rect 70813 21860 71000 21918
rect 70813 21814 70824 21860
rect 70870 21814 70928 21860
rect 70974 21814 71000 21860
rect 70813 21756 71000 21814
tri 36221 21603 36353 21735 ne
rect 36353 21724 36465 21735
rect 36353 21678 36354 21724
rect 36400 21678 36465 21724
rect 36353 21648 36465 21678
tri 36465 21648 36552 21735 sw
rect 70813 21710 70824 21756
rect 70870 21710 70928 21756
rect 70974 21710 71000 21756
rect 70813 21652 71000 21710
rect 36353 21603 36552 21648
tri 36353 21471 36485 21603 ne
rect 36485 21592 36552 21603
rect 36485 21546 36486 21592
rect 36532 21546 36552 21592
rect 36485 21471 36552 21546
tri 36552 21471 36729 21648 sw
rect 70813 21606 70824 21652
rect 70870 21606 70928 21652
rect 70974 21606 71000 21652
rect 70813 21548 71000 21606
rect 70813 21502 70824 21548
rect 70870 21502 70928 21548
rect 70974 21502 71000 21548
tri 36485 21339 36617 21471 ne
rect 36617 21460 36729 21471
rect 36617 21414 36618 21460
rect 36664 21414 36729 21460
rect 36617 21339 36729 21414
tri 36729 21339 36861 21471 sw
rect 70813 21444 71000 21502
rect 70813 21398 70824 21444
rect 70870 21398 70928 21444
rect 70974 21398 71000 21444
rect 70813 21340 71000 21398
tri 36617 21207 36749 21339 ne
rect 36749 21328 36861 21339
rect 36749 21282 36750 21328
rect 36796 21282 36861 21328
rect 36749 21207 36861 21282
tri 36861 21207 36993 21339 sw
rect 70813 21294 70824 21340
rect 70870 21294 70928 21340
rect 70974 21294 71000 21340
rect 70813 21236 71000 21294
tri 36749 21075 36881 21207 ne
rect 36881 21196 36993 21207
rect 36881 21150 36882 21196
rect 36928 21150 36993 21196
rect 36881 21075 36993 21150
tri 36993 21075 37125 21207 sw
rect 70813 21190 70824 21236
rect 70870 21190 70928 21236
rect 70974 21190 71000 21236
rect 70813 21132 71000 21190
rect 70813 21086 70824 21132
rect 70870 21086 70928 21132
rect 70974 21086 71000 21132
tri 36881 20943 37013 21075 ne
rect 37013 21064 37125 21075
rect 37013 21018 37014 21064
rect 37060 21018 37125 21064
rect 37013 20943 37125 21018
tri 37125 20943 37257 21075 sw
rect 70813 21028 71000 21086
rect 70813 20982 70824 21028
rect 70870 20982 70928 21028
rect 70974 20982 71000 21028
tri 37013 20811 37145 20943 ne
rect 37145 20932 37257 20943
rect 37145 20886 37146 20932
rect 37192 20886 37257 20932
rect 37145 20811 37257 20886
tri 37257 20811 37389 20943 sw
rect 70813 20924 71000 20982
rect 70813 20878 70824 20924
rect 70870 20878 70928 20924
rect 70974 20878 71000 20924
rect 70813 20820 71000 20878
tri 37145 20679 37277 20811 ne
rect 37277 20800 37389 20811
rect 37277 20754 37278 20800
rect 37324 20754 37389 20800
rect 37277 20679 37389 20754
tri 37277 20611 37345 20679 ne
rect 37345 20672 37389 20679
tri 37389 20672 37528 20811 sw
rect 70813 20774 70824 20820
rect 70870 20774 70928 20820
rect 70974 20774 71000 20820
rect 70813 20716 71000 20774
rect 37345 20668 37528 20672
rect 37345 20622 37410 20668
rect 37456 20622 37528 20668
rect 37345 20611 37528 20622
tri 37345 20428 37528 20611 ne
tri 37528 20547 37653 20672 sw
rect 70813 20670 70824 20716
rect 70870 20670 70928 20716
rect 70974 20670 71000 20716
rect 70813 20612 71000 20670
rect 70813 20566 70824 20612
rect 70870 20566 70928 20612
rect 70974 20566 71000 20612
rect 37528 20536 37653 20547
rect 37528 20490 37542 20536
rect 37588 20490 37653 20536
rect 37528 20428 37653 20490
tri 37653 20428 37772 20547 sw
rect 70813 20508 71000 20566
rect 70813 20462 70824 20508
rect 70870 20462 70928 20508
rect 70974 20462 71000 20508
tri 37528 20283 37673 20428 ne
rect 37673 20404 37772 20428
rect 37673 20358 37674 20404
rect 37720 20358 37772 20404
rect 37673 20283 37772 20358
tri 37772 20283 37917 20428 sw
rect 70813 20404 71000 20462
rect 70813 20358 70824 20404
rect 70870 20358 70928 20404
rect 70974 20358 71000 20404
rect 70813 20300 71000 20358
tri 37673 20151 37805 20283 ne
rect 37805 20272 37917 20283
rect 37805 20226 37806 20272
rect 37852 20226 37917 20272
rect 37805 20184 37917 20226
tri 37917 20184 38016 20283 sw
rect 70813 20254 70824 20300
rect 70870 20254 70928 20300
rect 70974 20254 71000 20300
rect 70813 20196 71000 20254
rect 37805 20151 38016 20184
tri 37805 20019 37937 20151 ne
rect 37937 20140 38016 20151
rect 37937 20094 37938 20140
rect 37984 20094 38016 20140
rect 37937 20019 38016 20094
tri 38016 20019 38181 20184 sw
rect 70813 20150 70824 20196
rect 70870 20150 70928 20196
rect 70974 20150 71000 20196
rect 70813 20092 71000 20150
rect 70813 20046 70824 20092
rect 70870 20046 70928 20092
rect 70974 20046 71000 20092
tri 37937 19887 38069 20019 ne
rect 38069 20008 38181 20019
rect 38069 19962 38070 20008
rect 38116 19962 38181 20008
rect 38069 19940 38181 19962
tri 38181 19940 38260 20019 sw
rect 70813 19988 71000 20046
rect 70813 19942 70824 19988
rect 70870 19942 70928 19988
rect 70974 19942 71000 19988
rect 38069 19887 38260 19940
tri 38069 19755 38201 19887 ne
rect 38201 19876 38260 19887
rect 38201 19830 38202 19876
rect 38248 19830 38260 19876
rect 38201 19755 38260 19830
tri 38260 19755 38445 19940 sw
rect 70813 19884 71000 19942
rect 70813 19838 70824 19884
rect 70870 19838 70928 19884
rect 70974 19838 71000 19884
rect 70813 19780 71000 19838
tri 38201 19623 38333 19755 ne
rect 38333 19744 38445 19755
rect 38333 19698 38334 19744
rect 38380 19698 38445 19744
rect 38333 19623 38445 19698
tri 38445 19623 38577 19755 sw
rect 70813 19734 70824 19780
rect 70870 19734 70928 19780
rect 70974 19734 71000 19780
rect 70813 19676 71000 19734
rect 70813 19630 70824 19676
rect 70870 19630 70928 19676
rect 70974 19630 71000 19676
tri 38333 19491 38465 19623 ne
rect 38465 19612 38577 19623
rect 38465 19566 38466 19612
rect 38512 19566 38577 19612
rect 38465 19491 38577 19566
tri 38577 19491 38709 19623 sw
rect 70813 19572 71000 19630
rect 70813 19526 70824 19572
rect 70870 19526 70928 19572
rect 70974 19526 71000 19572
tri 38465 19359 38597 19491 ne
rect 38597 19480 38709 19491
rect 38597 19434 38598 19480
rect 38644 19434 38709 19480
rect 38597 19359 38709 19434
tri 38709 19359 38841 19491 sw
rect 70813 19468 71000 19526
rect 70813 19422 70824 19468
rect 70870 19422 70928 19468
rect 70974 19422 71000 19468
rect 70813 19364 71000 19422
tri 38597 19227 38729 19359 ne
rect 38729 19348 38841 19359
rect 38729 19302 38730 19348
rect 38776 19302 38841 19348
rect 38729 19227 38841 19302
tri 38841 19227 38973 19359 sw
rect 70813 19318 70824 19364
rect 70870 19318 70928 19364
rect 70974 19318 71000 19364
rect 70813 19260 71000 19318
tri 38729 19095 38861 19227 ne
rect 38861 19216 38973 19227
rect 38861 19170 38862 19216
rect 38908 19170 38973 19216
rect 38861 19095 38973 19170
tri 38973 19095 39105 19227 sw
rect 70813 19214 70824 19260
rect 70870 19214 70928 19260
rect 70974 19214 71000 19260
rect 70813 19156 71000 19214
rect 70813 19110 70824 19156
rect 70870 19110 70928 19156
rect 70974 19110 71000 19156
tri 38861 18963 38993 19095 ne
rect 38993 19084 39105 19095
rect 38993 19038 38994 19084
rect 39040 19038 39105 19084
rect 38993 18964 39105 19038
tri 39105 18964 39236 19095 sw
rect 70813 19052 71000 19110
rect 70813 19006 70824 19052
rect 70870 19006 70928 19052
rect 70974 19006 71000 19052
rect 38993 18963 39236 18964
tri 38993 18831 39125 18963 ne
rect 39125 18952 39236 18963
rect 39125 18906 39126 18952
rect 39172 18906 39236 18952
rect 39125 18831 39236 18906
tri 39236 18831 39369 18964 sw
rect 70813 18948 71000 19006
rect 70813 18902 70824 18948
rect 70870 18902 70928 18948
rect 70974 18902 71000 18948
rect 70813 18844 71000 18902
tri 39125 18699 39257 18831 ne
rect 39257 18820 39369 18831
rect 39257 18774 39258 18820
rect 39304 18774 39369 18820
rect 39257 18720 39369 18774
tri 39369 18720 39480 18831 sw
rect 70813 18798 70824 18844
rect 70870 18798 70928 18844
rect 70974 18798 71000 18844
rect 70813 18740 71000 18798
rect 39257 18699 39480 18720
tri 39257 18567 39389 18699 ne
rect 39389 18688 39480 18699
rect 39389 18642 39390 18688
rect 39436 18642 39480 18688
rect 39389 18567 39480 18642
tri 39480 18567 39633 18720 sw
rect 70813 18694 70824 18740
rect 70870 18694 70928 18740
rect 70974 18694 71000 18740
rect 70813 18636 71000 18694
rect 70813 18590 70824 18636
rect 70870 18590 70928 18636
rect 70974 18590 71000 18636
tri 39389 18435 39521 18567 ne
rect 39521 18556 39633 18567
rect 39521 18510 39522 18556
rect 39568 18510 39633 18556
rect 39521 18476 39633 18510
tri 39633 18476 39724 18567 sw
rect 70813 18532 71000 18590
rect 70813 18486 70824 18532
rect 70870 18486 70928 18532
rect 70974 18486 71000 18532
rect 39521 18435 39724 18476
tri 39521 18303 39653 18435 ne
rect 39653 18424 39724 18435
rect 39653 18378 39654 18424
rect 39700 18378 39724 18424
rect 39653 18303 39724 18378
tri 39724 18303 39897 18476 sw
rect 70813 18428 71000 18486
rect 70813 18382 70824 18428
rect 70870 18382 70928 18428
rect 70974 18382 71000 18428
rect 70813 18324 71000 18382
tri 39653 18171 39785 18303 ne
rect 39785 18292 39897 18303
rect 39785 18246 39786 18292
rect 39832 18246 39897 18292
rect 39785 18171 39897 18246
tri 39897 18171 40029 18303 sw
rect 70813 18278 70824 18324
rect 70870 18278 70928 18324
rect 70974 18278 71000 18324
rect 70813 18220 71000 18278
rect 70813 18174 70824 18220
rect 70870 18174 70928 18220
rect 70974 18174 71000 18220
tri 39785 18039 39917 18171 ne
rect 39917 18160 40029 18171
rect 39917 18114 39918 18160
rect 39964 18114 40029 18160
rect 39917 18039 40029 18114
tri 40029 18039 40161 18171 sw
rect 70813 18116 71000 18174
rect 70813 18070 70824 18116
rect 70870 18070 70928 18116
rect 70974 18070 71000 18116
tri 39917 17907 40049 18039 ne
rect 40049 18028 40161 18039
rect 40049 17982 40050 18028
rect 40096 17982 40161 18028
rect 40049 17907 40161 17982
tri 40161 17907 40293 18039 sw
rect 70813 18012 71000 18070
rect 70813 17966 70824 18012
rect 70870 17966 70928 18012
rect 70974 17966 71000 18012
rect 70813 17908 71000 17966
tri 40049 17775 40181 17907 ne
rect 40181 17896 40293 17907
rect 40181 17850 40182 17896
rect 40228 17850 40293 17896
rect 40181 17775 40293 17850
tri 40293 17775 40425 17907 sw
rect 70813 17862 70824 17908
rect 70870 17862 70928 17908
rect 70974 17862 71000 17908
rect 70813 17804 71000 17862
tri 40181 17643 40313 17775 ne
rect 40313 17764 40425 17775
rect 40313 17718 40314 17764
rect 40360 17718 40425 17764
rect 40313 17643 40425 17718
tri 40425 17643 40557 17775 sw
rect 70813 17758 70824 17804
rect 70870 17758 70928 17804
rect 70974 17758 71000 17804
rect 70813 17700 71000 17758
rect 70813 17654 70824 17700
rect 70870 17654 70928 17700
rect 70974 17654 71000 17700
tri 40313 17511 40445 17643 ne
rect 40445 17632 40557 17643
rect 40445 17586 40446 17632
rect 40492 17586 40557 17632
rect 40445 17511 40557 17586
tri 40445 17443 40513 17511 ne
rect 40513 17500 40557 17511
tri 40557 17500 40700 17643 sw
rect 70813 17596 71000 17654
rect 70813 17550 70824 17596
rect 70870 17550 70928 17596
rect 70974 17550 71000 17596
rect 40513 17454 40578 17500
rect 40624 17454 40700 17500
rect 40513 17443 40700 17454
tri 40513 17256 40700 17443 ne
tri 40700 17379 40821 17500 sw
rect 70813 17492 71000 17550
rect 70813 17446 70824 17492
rect 70870 17446 70928 17492
rect 70974 17446 71000 17492
rect 70813 17388 71000 17446
rect 40700 17368 40821 17379
rect 40700 17322 40710 17368
rect 40756 17322 40821 17368
rect 40700 17256 40821 17322
tri 40821 17256 40944 17379 sw
rect 70813 17342 70824 17388
rect 70870 17342 70928 17388
rect 70974 17342 71000 17388
rect 70813 17284 71000 17342
tri 40700 17115 40841 17256 ne
rect 40841 17236 40944 17256
rect 40841 17190 40842 17236
rect 40888 17190 40944 17236
rect 40841 17115 40944 17190
tri 40944 17115 41085 17256 sw
rect 70813 17238 70824 17284
rect 70870 17238 70928 17284
rect 70974 17238 71000 17284
rect 70813 17180 71000 17238
rect 70813 17134 70824 17180
rect 70870 17134 70928 17180
rect 70974 17134 71000 17180
tri 40841 16983 40973 17115 ne
rect 40973 17104 41085 17115
rect 40973 17058 40974 17104
rect 41020 17058 41085 17104
rect 40973 17012 41085 17058
tri 41085 17012 41188 17115 sw
rect 70813 17076 71000 17134
rect 70813 17030 70824 17076
rect 70870 17030 70928 17076
rect 70974 17030 71000 17076
rect 40973 16983 41188 17012
tri 40973 16851 41105 16983 ne
rect 41105 16972 41188 16983
rect 41105 16926 41106 16972
rect 41152 16926 41188 16972
rect 41105 16851 41188 16926
tri 41188 16851 41349 17012 sw
rect 70813 16972 71000 17030
rect 70813 16926 70824 16972
rect 70870 16926 70928 16972
rect 70974 16926 71000 16972
rect 70813 16868 71000 16926
tri 41105 16719 41237 16851 ne
rect 41237 16840 41349 16851
rect 41237 16794 41238 16840
rect 41284 16794 41349 16840
rect 41237 16768 41349 16794
tri 41349 16768 41432 16851 sw
rect 70813 16822 70824 16868
rect 70870 16822 70928 16868
rect 70974 16822 71000 16868
rect 41237 16719 41432 16768
tri 41237 16587 41369 16719 ne
rect 41369 16708 41432 16719
rect 41369 16662 41370 16708
rect 41416 16662 41432 16708
rect 41369 16587 41432 16662
tri 41432 16587 41613 16768 sw
rect 70813 16764 71000 16822
rect 70813 16718 70824 16764
rect 70870 16718 70928 16764
rect 70974 16718 71000 16764
rect 70813 16660 71000 16718
rect 70813 16614 70824 16660
rect 70870 16614 70928 16660
rect 70974 16614 71000 16660
tri 41369 16455 41501 16587 ne
rect 41501 16576 41613 16587
rect 41501 16530 41502 16576
rect 41548 16530 41613 16576
rect 41501 16455 41613 16530
tri 41613 16455 41745 16587 sw
rect 70813 16556 71000 16614
rect 70813 16510 70824 16556
rect 70870 16510 70928 16556
rect 70974 16510 71000 16556
tri 41501 16323 41633 16455 ne
rect 41633 16444 41745 16455
rect 41633 16398 41634 16444
rect 41680 16398 41745 16444
rect 41633 16323 41745 16398
tri 41745 16323 41877 16455 sw
rect 70813 16452 71000 16510
rect 70813 16406 70824 16452
rect 70870 16406 70928 16452
rect 70974 16406 71000 16452
rect 70813 16348 71000 16406
tri 41633 16191 41765 16323 ne
rect 41765 16312 41877 16323
rect 41765 16266 41766 16312
rect 41812 16266 41877 16312
rect 41765 16191 41877 16266
tri 41877 16191 42009 16323 sw
rect 70813 16302 70824 16348
rect 70870 16302 70928 16348
rect 70974 16302 71000 16348
rect 70813 16244 71000 16302
rect 70813 16198 70824 16244
rect 70870 16198 70928 16244
rect 70974 16198 71000 16244
tri 41765 16059 41897 16191 ne
rect 41897 16180 42009 16191
rect 41897 16134 41898 16180
rect 41944 16134 42009 16180
rect 41897 16059 42009 16134
tri 42009 16059 42141 16191 sw
rect 70813 16140 71000 16198
rect 70813 16094 70824 16140
rect 70870 16094 70928 16140
rect 70974 16094 71000 16140
tri 41897 15927 42029 16059 ne
rect 42029 16048 42141 16059
rect 42029 16002 42030 16048
rect 42076 16002 42141 16048
rect 42029 15927 42141 16002
tri 42141 15927 42273 16059 sw
rect 70813 16036 71000 16094
rect 70813 15990 70824 16036
rect 70870 15990 70928 16036
rect 70974 15990 71000 16036
rect 70813 15932 71000 15990
tri 42029 15795 42161 15927 ne
rect 42161 15916 42273 15927
rect 42161 15870 42162 15916
rect 42208 15870 42273 15916
rect 42161 15795 42273 15870
tri 42161 15727 42229 15795 ne
rect 42229 15792 42273 15795
tri 42273 15792 42408 15927 sw
rect 70813 15886 70824 15932
rect 70870 15886 70928 15932
rect 70974 15886 71000 15932
rect 70813 15828 71000 15886
rect 42229 15784 42408 15792
rect 42229 15738 42294 15784
rect 42340 15738 42408 15784
rect 42229 15727 42408 15738
tri 42229 15548 42408 15727 ne
tri 42408 15663 42537 15792 sw
rect 70813 15782 70824 15828
rect 70870 15782 70928 15828
rect 70974 15782 71000 15828
rect 70813 15724 71000 15782
rect 70813 15678 70824 15724
rect 70870 15678 70928 15724
rect 70974 15678 71000 15724
rect 42408 15652 42537 15663
rect 42408 15606 42426 15652
rect 42472 15606 42537 15652
rect 42408 15548 42537 15606
tri 42537 15548 42652 15663 sw
rect 70813 15620 71000 15678
rect 70813 15574 70824 15620
rect 70870 15574 70928 15620
rect 70974 15574 71000 15620
tri 42408 15399 42557 15548 ne
rect 42557 15520 42652 15548
rect 42557 15474 42558 15520
rect 42604 15474 42652 15520
rect 42557 15399 42652 15474
tri 42652 15399 42801 15548 sw
rect 70813 15516 71000 15574
rect 70813 15470 70824 15516
rect 70870 15470 70928 15516
rect 70974 15470 71000 15516
rect 70813 15412 71000 15470
tri 42557 15267 42689 15399 ne
rect 42689 15388 42801 15399
rect 42689 15342 42690 15388
rect 42736 15342 42801 15388
rect 42689 15304 42801 15342
tri 42801 15304 42896 15399 sw
rect 70813 15366 70824 15412
rect 70870 15366 70928 15412
rect 70974 15366 71000 15412
rect 70813 15308 71000 15366
rect 42689 15267 42896 15304
tri 42689 15135 42821 15267 ne
rect 42821 15256 42896 15267
rect 42821 15210 42822 15256
rect 42868 15210 42896 15256
rect 42821 15135 42896 15210
tri 42896 15135 43065 15304 sw
rect 70813 15262 70824 15308
rect 70870 15262 70928 15308
rect 70974 15262 71000 15308
rect 70813 15204 71000 15262
rect 70813 15158 70824 15204
rect 70870 15158 70928 15204
rect 70974 15158 71000 15204
tri 42821 15003 42953 15135 ne
rect 42953 15124 43065 15135
rect 42953 15078 42954 15124
rect 43000 15078 43065 15124
rect 42953 15003 43065 15078
tri 43065 15003 43197 15135 sw
rect 70813 15100 71000 15158
rect 70813 15054 70824 15100
rect 70870 15054 70928 15100
rect 70974 15054 71000 15100
tri 42953 14871 43085 15003 ne
rect 43085 14992 43197 15003
rect 43085 14946 43086 14992
rect 43132 14946 43197 14992
rect 43085 14871 43197 14946
tri 43197 14871 43329 15003 sw
rect 70813 14996 71000 15054
rect 70813 14950 70824 14996
rect 70870 14950 70928 14996
rect 70974 14950 71000 14996
rect 70813 14892 71000 14950
tri 43085 14739 43217 14871 ne
rect 43217 14860 43329 14871
rect 43217 14814 43218 14860
rect 43264 14814 43329 14860
rect 43217 14739 43329 14814
tri 43329 14739 43461 14871 sw
rect 70813 14846 70824 14892
rect 70870 14846 70928 14892
rect 70974 14846 71000 14892
rect 70813 14788 71000 14846
rect 70813 14742 70824 14788
rect 70870 14742 70928 14788
rect 70974 14742 71000 14788
tri 43217 14607 43349 14739 ne
rect 43349 14728 43461 14739
rect 43349 14682 43350 14728
rect 43396 14682 43461 14728
rect 43349 14607 43461 14682
tri 43461 14607 43593 14739 sw
rect 70813 14684 71000 14742
rect 70813 14638 70824 14684
rect 70870 14638 70928 14684
rect 70974 14638 71000 14684
tri 43349 14475 43481 14607 ne
rect 43481 14596 43593 14607
rect 43481 14550 43482 14596
rect 43528 14550 43593 14596
rect 43481 14475 43593 14550
tri 43593 14475 43725 14607 sw
rect 70813 14580 71000 14638
rect 70813 14534 70824 14580
rect 70870 14534 70928 14580
rect 70974 14534 71000 14580
rect 70813 14476 71000 14534
tri 43481 14343 43613 14475 ne
rect 43613 14464 43725 14475
rect 43613 14418 43614 14464
rect 43660 14418 43725 14464
rect 43613 14343 43725 14418
tri 43725 14343 43857 14475 sw
rect 70813 14430 70824 14476
rect 70870 14430 70928 14476
rect 70974 14430 71000 14476
rect 70813 14372 71000 14430
tri 43613 14211 43745 14343 ne
rect 43745 14332 43857 14343
rect 43745 14286 43746 14332
rect 43792 14286 43857 14332
rect 43745 14211 43857 14286
tri 43857 14211 43989 14343 sw
rect 70813 14326 70824 14372
rect 70870 14326 70928 14372
rect 70974 14326 71000 14372
rect 70813 14268 71000 14326
rect 70813 14222 70824 14268
rect 70870 14222 70928 14268
rect 70974 14222 71000 14268
tri 43745 14079 43877 14211 ne
rect 43877 14200 43989 14211
rect 43877 14154 43878 14200
rect 43924 14154 43989 14200
rect 43877 14084 43989 14154
tri 43989 14084 44116 14211 sw
rect 70813 14164 71000 14222
rect 70813 14118 70824 14164
rect 70870 14118 70928 14164
rect 70974 14118 71000 14164
rect 43877 14079 44116 14084
tri 43877 13947 44009 14079 ne
rect 44009 14068 44116 14079
rect 44009 14022 44010 14068
rect 44056 14022 44116 14068
rect 44009 13947 44116 14022
tri 44116 13947 44253 14084 sw
rect 70813 14060 71000 14118
rect 70813 14014 70824 14060
rect 70870 14014 70928 14060
rect 70974 14014 71000 14060
rect 70813 13956 71000 14014
tri 44009 13815 44141 13947 ne
rect 44141 13936 44253 13947
rect 44141 13890 44142 13936
rect 44188 13890 44253 13936
rect 44141 13840 44253 13890
tri 44253 13840 44360 13947 sw
rect 70813 13910 70824 13956
rect 70870 13910 70928 13956
rect 70974 13910 71000 13956
rect 70813 13852 71000 13910
rect 44141 13815 44360 13840
tri 44141 13683 44273 13815 ne
rect 44273 13804 44360 13815
rect 44273 13758 44274 13804
rect 44320 13758 44360 13804
rect 44273 13683 44360 13758
tri 44360 13683 44517 13840 sw
rect 70813 13806 70824 13852
rect 70870 13806 70928 13852
rect 70974 13806 71000 13852
rect 70813 13748 71000 13806
rect 70813 13702 70824 13748
rect 70870 13702 70928 13748
rect 70974 13702 71000 13748
tri 44273 13551 44405 13683 ne
rect 44405 13672 44517 13683
rect 44405 13626 44406 13672
rect 44452 13626 44517 13672
rect 44405 13596 44517 13626
tri 44517 13596 44604 13683 sw
rect 70813 13644 71000 13702
rect 70813 13598 70824 13644
rect 70870 13598 70928 13644
rect 70974 13598 71000 13644
rect 44405 13551 44604 13596
tri 44405 13419 44537 13551 ne
rect 44537 13540 44604 13551
rect 44537 13494 44538 13540
rect 44584 13494 44604 13540
rect 44537 13419 44604 13494
tri 44604 13419 44781 13596 sw
rect 70813 13540 71000 13598
rect 70813 13494 70824 13540
rect 70870 13494 70928 13540
rect 70974 13494 71000 13540
rect 70813 13436 71000 13494
tri 44537 13351 44605 13419 ne
rect 44605 13408 44781 13419
rect 44605 13362 44670 13408
rect 44716 13362 44781 13408
rect 44605 13352 44781 13362
tri 44781 13352 44848 13419 sw
rect 70813 13390 70824 13436
rect 70870 13390 70928 13436
rect 70974 13390 71000 13436
rect 44605 13351 44848 13352
tri 44605 13108 44848 13351 ne
tri 44848 13280 44920 13352 sw
rect 70813 13280 71000 13390
rect 44848 13269 71000 13280
rect 44848 13256 45088 13269
rect 44848 13210 44850 13256
rect 44896 13223 45088 13256
rect 45134 13223 45192 13269
rect 45238 13223 45296 13269
rect 45342 13223 45400 13269
rect 45446 13223 45504 13269
rect 45550 13223 45608 13269
rect 45654 13223 45712 13269
rect 45758 13223 45816 13269
rect 45862 13223 45920 13269
rect 45966 13223 46024 13269
rect 46070 13223 46128 13269
rect 46174 13223 46232 13269
rect 46278 13223 46336 13269
rect 46382 13223 46440 13269
rect 46486 13223 46544 13269
rect 46590 13223 46648 13269
rect 46694 13223 46752 13269
rect 46798 13223 46856 13269
rect 46902 13223 46960 13269
rect 47006 13223 47064 13269
rect 47110 13223 47168 13269
rect 47214 13223 47272 13269
rect 47318 13223 47376 13269
rect 47422 13223 47480 13269
rect 47526 13223 47584 13269
rect 47630 13223 47688 13269
rect 47734 13223 47792 13269
rect 47838 13223 47896 13269
rect 47942 13223 48000 13269
rect 48046 13223 48104 13269
rect 48150 13223 48208 13269
rect 48254 13223 48312 13269
rect 48358 13223 48416 13269
rect 48462 13223 48520 13269
rect 48566 13223 48624 13269
rect 48670 13223 48728 13269
rect 48774 13223 48832 13269
rect 48878 13223 48936 13269
rect 48982 13223 49040 13269
rect 49086 13223 49144 13269
rect 49190 13223 49248 13269
rect 49294 13223 49352 13269
rect 49398 13223 49456 13269
rect 49502 13223 49560 13269
rect 49606 13223 49664 13269
rect 49710 13223 49768 13269
rect 49814 13223 49872 13269
rect 49918 13223 49976 13269
rect 50022 13223 50080 13269
rect 50126 13223 50184 13269
rect 50230 13223 50288 13269
rect 50334 13223 50392 13269
rect 50438 13223 50496 13269
rect 50542 13223 50600 13269
rect 50646 13223 50704 13269
rect 50750 13223 50808 13269
rect 50854 13223 50912 13269
rect 50958 13223 51016 13269
rect 51062 13223 51120 13269
rect 51166 13223 51224 13269
rect 51270 13223 51328 13269
rect 51374 13223 51432 13269
rect 51478 13223 51536 13269
rect 51582 13223 51640 13269
rect 51686 13223 51744 13269
rect 51790 13223 51848 13269
rect 51894 13223 51952 13269
rect 51998 13223 52056 13269
rect 52102 13223 52160 13269
rect 52206 13223 52264 13269
rect 52310 13223 52368 13269
rect 52414 13223 52472 13269
rect 52518 13223 52576 13269
rect 52622 13223 52680 13269
rect 52726 13223 52784 13269
rect 52830 13223 52888 13269
rect 52934 13223 52992 13269
rect 53038 13223 53096 13269
rect 53142 13223 53200 13269
rect 53246 13223 53304 13269
rect 53350 13223 53408 13269
rect 53454 13223 53512 13269
rect 53558 13223 53616 13269
rect 53662 13223 53720 13269
rect 53766 13223 53824 13269
rect 53870 13223 53928 13269
rect 53974 13223 54032 13269
rect 54078 13223 54136 13269
rect 54182 13223 54240 13269
rect 54286 13223 54344 13269
rect 54390 13223 54448 13269
rect 54494 13223 54552 13269
rect 54598 13223 54656 13269
rect 54702 13223 54760 13269
rect 54806 13223 54864 13269
rect 54910 13223 54968 13269
rect 55014 13223 55072 13269
rect 55118 13223 55176 13269
rect 55222 13223 55280 13269
rect 55326 13223 55384 13269
rect 55430 13223 55488 13269
rect 55534 13223 55592 13269
rect 55638 13223 55696 13269
rect 55742 13223 55800 13269
rect 55846 13223 55904 13269
rect 55950 13223 56008 13269
rect 56054 13223 56112 13269
rect 56158 13223 56216 13269
rect 56262 13223 56320 13269
rect 56366 13223 56424 13269
rect 56470 13223 56528 13269
rect 56574 13223 56632 13269
rect 56678 13223 56736 13269
rect 56782 13223 56840 13269
rect 56886 13223 56944 13269
rect 56990 13223 57048 13269
rect 57094 13223 57152 13269
rect 57198 13223 57256 13269
rect 57302 13223 57360 13269
rect 57406 13223 57464 13269
rect 57510 13223 57568 13269
rect 57614 13223 57672 13269
rect 57718 13223 57776 13269
rect 57822 13223 57880 13269
rect 57926 13223 57984 13269
rect 58030 13223 58088 13269
rect 58134 13223 58192 13269
rect 58238 13223 58296 13269
rect 58342 13223 58400 13269
rect 58446 13223 58504 13269
rect 58550 13223 58608 13269
rect 58654 13223 58712 13269
rect 58758 13223 58816 13269
rect 58862 13223 58920 13269
rect 58966 13223 59024 13269
rect 59070 13223 59128 13269
rect 59174 13223 59232 13269
rect 59278 13223 59336 13269
rect 59382 13223 59440 13269
rect 59486 13223 59544 13269
rect 59590 13223 59648 13269
rect 59694 13223 59752 13269
rect 59798 13223 59856 13269
rect 59902 13223 59960 13269
rect 60006 13223 60064 13269
rect 60110 13223 60168 13269
rect 60214 13223 60272 13269
rect 60318 13223 60376 13269
rect 60422 13223 60480 13269
rect 60526 13223 60584 13269
rect 60630 13223 60688 13269
rect 60734 13223 60792 13269
rect 60838 13223 60896 13269
rect 60942 13223 61000 13269
rect 61046 13223 61104 13269
rect 61150 13223 61208 13269
rect 61254 13223 61312 13269
rect 61358 13223 61416 13269
rect 61462 13223 61520 13269
rect 61566 13223 61624 13269
rect 61670 13223 61728 13269
rect 61774 13223 61832 13269
rect 61878 13223 61936 13269
rect 61982 13223 62040 13269
rect 62086 13223 62144 13269
rect 62190 13223 62248 13269
rect 62294 13223 62352 13269
rect 62398 13223 62456 13269
rect 62502 13223 62560 13269
rect 62606 13223 62664 13269
rect 62710 13223 62768 13269
rect 62814 13223 62872 13269
rect 62918 13223 62976 13269
rect 63022 13223 63080 13269
rect 63126 13223 63184 13269
rect 63230 13223 63288 13269
rect 63334 13223 63392 13269
rect 63438 13223 63496 13269
rect 63542 13223 63600 13269
rect 63646 13223 63704 13269
rect 63750 13223 63808 13269
rect 63854 13223 63912 13269
rect 63958 13223 64016 13269
rect 64062 13223 64120 13269
rect 64166 13223 64224 13269
rect 64270 13223 64328 13269
rect 64374 13223 64432 13269
rect 64478 13223 64536 13269
rect 64582 13223 64640 13269
rect 64686 13223 64744 13269
rect 64790 13223 64848 13269
rect 64894 13223 64952 13269
rect 64998 13223 65056 13269
rect 65102 13223 65160 13269
rect 65206 13223 65264 13269
rect 65310 13223 65368 13269
rect 65414 13223 65472 13269
rect 65518 13223 65576 13269
rect 65622 13223 65680 13269
rect 65726 13223 65784 13269
rect 65830 13223 65888 13269
rect 65934 13223 65992 13269
rect 66038 13223 66096 13269
rect 66142 13223 66200 13269
rect 66246 13223 66304 13269
rect 66350 13223 66408 13269
rect 66454 13223 66512 13269
rect 66558 13223 66616 13269
rect 66662 13223 66720 13269
rect 66766 13223 66824 13269
rect 66870 13223 66928 13269
rect 66974 13223 67032 13269
rect 67078 13223 67136 13269
rect 67182 13223 67240 13269
rect 67286 13223 67344 13269
rect 67390 13223 67448 13269
rect 67494 13223 67552 13269
rect 67598 13223 67656 13269
rect 67702 13223 67760 13269
rect 67806 13223 67864 13269
rect 67910 13223 67968 13269
rect 68014 13223 68072 13269
rect 68118 13223 68176 13269
rect 68222 13223 68280 13269
rect 68326 13223 68384 13269
rect 68430 13223 68488 13269
rect 68534 13223 68592 13269
rect 68638 13223 68696 13269
rect 68742 13223 68800 13269
rect 68846 13223 68904 13269
rect 68950 13223 69008 13269
rect 69054 13223 69112 13269
rect 69158 13223 69216 13269
rect 69262 13223 69320 13269
rect 69366 13223 69424 13269
rect 69470 13223 69528 13269
rect 69574 13223 69632 13269
rect 69678 13223 69736 13269
rect 69782 13223 69840 13269
rect 69886 13223 69944 13269
rect 69990 13223 70048 13269
rect 70094 13223 70152 13269
rect 70198 13223 70256 13269
rect 70302 13223 70360 13269
rect 70406 13223 70464 13269
rect 70510 13223 70568 13269
rect 70614 13223 70672 13269
rect 70718 13223 70776 13269
rect 70822 13223 70880 13269
rect 70926 13223 71000 13269
rect 44896 13210 71000 13223
rect 44848 13165 71000 13210
rect 44848 13119 45088 13165
rect 45134 13119 45192 13165
rect 45238 13119 45296 13165
rect 45342 13119 45400 13165
rect 45446 13119 45504 13165
rect 45550 13119 45608 13165
rect 45654 13119 45712 13165
rect 45758 13119 45816 13165
rect 45862 13119 45920 13165
rect 45966 13119 46024 13165
rect 46070 13119 46128 13165
rect 46174 13119 46232 13165
rect 46278 13119 46336 13165
rect 46382 13119 46440 13165
rect 46486 13119 46544 13165
rect 46590 13119 46648 13165
rect 46694 13119 46752 13165
rect 46798 13119 46856 13165
rect 46902 13119 46960 13165
rect 47006 13119 47064 13165
rect 47110 13119 47168 13165
rect 47214 13119 47272 13165
rect 47318 13119 47376 13165
rect 47422 13119 47480 13165
rect 47526 13119 47584 13165
rect 47630 13119 47688 13165
rect 47734 13119 47792 13165
rect 47838 13119 47896 13165
rect 47942 13119 48000 13165
rect 48046 13119 48104 13165
rect 48150 13119 48208 13165
rect 48254 13119 48312 13165
rect 48358 13119 48416 13165
rect 48462 13119 48520 13165
rect 48566 13119 48624 13165
rect 48670 13119 48728 13165
rect 48774 13119 48832 13165
rect 48878 13119 48936 13165
rect 48982 13119 49040 13165
rect 49086 13119 49144 13165
rect 49190 13119 49248 13165
rect 49294 13119 49352 13165
rect 49398 13119 49456 13165
rect 49502 13119 49560 13165
rect 49606 13119 49664 13165
rect 49710 13119 49768 13165
rect 49814 13119 49872 13165
rect 49918 13119 49976 13165
rect 50022 13119 50080 13165
rect 50126 13119 50184 13165
rect 50230 13119 50288 13165
rect 50334 13119 50392 13165
rect 50438 13119 50496 13165
rect 50542 13119 50600 13165
rect 50646 13119 50704 13165
rect 50750 13119 50808 13165
rect 50854 13119 50912 13165
rect 50958 13119 51016 13165
rect 51062 13119 51120 13165
rect 51166 13119 51224 13165
rect 51270 13119 51328 13165
rect 51374 13119 51432 13165
rect 51478 13119 51536 13165
rect 51582 13119 51640 13165
rect 51686 13119 51744 13165
rect 51790 13119 51848 13165
rect 51894 13119 51952 13165
rect 51998 13119 52056 13165
rect 52102 13119 52160 13165
rect 52206 13119 52264 13165
rect 52310 13119 52368 13165
rect 52414 13119 52472 13165
rect 52518 13119 52576 13165
rect 52622 13119 52680 13165
rect 52726 13119 52784 13165
rect 52830 13119 52888 13165
rect 52934 13119 52992 13165
rect 53038 13119 53096 13165
rect 53142 13119 53200 13165
rect 53246 13119 53304 13165
rect 53350 13119 53408 13165
rect 53454 13119 53512 13165
rect 53558 13119 53616 13165
rect 53662 13119 53720 13165
rect 53766 13119 53824 13165
rect 53870 13119 53928 13165
rect 53974 13119 54032 13165
rect 54078 13119 54136 13165
rect 54182 13119 54240 13165
rect 54286 13119 54344 13165
rect 54390 13119 54448 13165
rect 54494 13119 54552 13165
rect 54598 13119 54656 13165
rect 54702 13119 54760 13165
rect 54806 13119 54864 13165
rect 54910 13119 54968 13165
rect 55014 13119 55072 13165
rect 55118 13119 55176 13165
rect 55222 13119 55280 13165
rect 55326 13119 55384 13165
rect 55430 13119 55488 13165
rect 55534 13119 55592 13165
rect 55638 13119 55696 13165
rect 55742 13119 55800 13165
rect 55846 13119 55904 13165
rect 55950 13119 56008 13165
rect 56054 13119 56112 13165
rect 56158 13119 56216 13165
rect 56262 13119 56320 13165
rect 56366 13119 56424 13165
rect 56470 13119 56528 13165
rect 56574 13119 56632 13165
rect 56678 13119 56736 13165
rect 56782 13119 56840 13165
rect 56886 13119 56944 13165
rect 56990 13119 57048 13165
rect 57094 13119 57152 13165
rect 57198 13119 57256 13165
rect 57302 13119 57360 13165
rect 57406 13119 57464 13165
rect 57510 13119 57568 13165
rect 57614 13119 57672 13165
rect 57718 13119 57776 13165
rect 57822 13119 57880 13165
rect 57926 13119 57984 13165
rect 58030 13119 58088 13165
rect 58134 13119 58192 13165
rect 58238 13119 58296 13165
rect 58342 13119 58400 13165
rect 58446 13119 58504 13165
rect 58550 13119 58608 13165
rect 58654 13119 58712 13165
rect 58758 13119 58816 13165
rect 58862 13119 58920 13165
rect 58966 13119 59024 13165
rect 59070 13119 59128 13165
rect 59174 13119 59232 13165
rect 59278 13119 59336 13165
rect 59382 13119 59440 13165
rect 59486 13119 59544 13165
rect 59590 13119 59648 13165
rect 59694 13119 59752 13165
rect 59798 13119 59856 13165
rect 59902 13119 59960 13165
rect 60006 13119 60064 13165
rect 60110 13119 60168 13165
rect 60214 13119 60272 13165
rect 60318 13119 60376 13165
rect 60422 13119 60480 13165
rect 60526 13119 60584 13165
rect 60630 13119 60688 13165
rect 60734 13119 60792 13165
rect 60838 13119 60896 13165
rect 60942 13119 61000 13165
rect 61046 13119 61104 13165
rect 61150 13119 61208 13165
rect 61254 13119 61312 13165
rect 61358 13119 61416 13165
rect 61462 13119 61520 13165
rect 61566 13119 61624 13165
rect 61670 13119 61728 13165
rect 61774 13119 61832 13165
rect 61878 13119 61936 13165
rect 61982 13119 62040 13165
rect 62086 13119 62144 13165
rect 62190 13119 62248 13165
rect 62294 13119 62352 13165
rect 62398 13119 62456 13165
rect 62502 13119 62560 13165
rect 62606 13119 62664 13165
rect 62710 13119 62768 13165
rect 62814 13119 62872 13165
rect 62918 13119 62976 13165
rect 63022 13119 63080 13165
rect 63126 13119 63184 13165
rect 63230 13119 63288 13165
rect 63334 13119 63392 13165
rect 63438 13119 63496 13165
rect 63542 13119 63600 13165
rect 63646 13119 63704 13165
rect 63750 13119 63808 13165
rect 63854 13119 63912 13165
rect 63958 13119 64016 13165
rect 64062 13119 64120 13165
rect 64166 13119 64224 13165
rect 64270 13119 64328 13165
rect 64374 13119 64432 13165
rect 64478 13119 64536 13165
rect 64582 13119 64640 13165
rect 64686 13119 64744 13165
rect 64790 13119 64848 13165
rect 64894 13119 64952 13165
rect 64998 13119 65056 13165
rect 65102 13119 65160 13165
rect 65206 13119 65264 13165
rect 65310 13119 65368 13165
rect 65414 13119 65472 13165
rect 65518 13119 65576 13165
rect 65622 13119 65680 13165
rect 65726 13119 65784 13165
rect 65830 13119 65888 13165
rect 65934 13119 65992 13165
rect 66038 13119 66096 13165
rect 66142 13119 66200 13165
rect 66246 13119 66304 13165
rect 66350 13119 66408 13165
rect 66454 13119 66512 13165
rect 66558 13119 66616 13165
rect 66662 13119 66720 13165
rect 66766 13119 66824 13165
rect 66870 13119 66928 13165
rect 66974 13119 67032 13165
rect 67078 13119 67136 13165
rect 67182 13119 67240 13165
rect 67286 13119 67344 13165
rect 67390 13119 67448 13165
rect 67494 13119 67552 13165
rect 67598 13119 67656 13165
rect 67702 13119 67760 13165
rect 67806 13119 67864 13165
rect 67910 13119 67968 13165
rect 68014 13119 68072 13165
rect 68118 13119 68176 13165
rect 68222 13119 68280 13165
rect 68326 13119 68384 13165
rect 68430 13119 68488 13165
rect 68534 13119 68592 13165
rect 68638 13119 68696 13165
rect 68742 13119 68800 13165
rect 68846 13119 68904 13165
rect 68950 13119 69008 13165
rect 69054 13119 69112 13165
rect 69158 13119 69216 13165
rect 69262 13119 69320 13165
rect 69366 13119 69424 13165
rect 69470 13119 69528 13165
rect 69574 13119 69632 13165
rect 69678 13119 69736 13165
rect 69782 13119 69840 13165
rect 69886 13119 69944 13165
rect 69990 13119 70048 13165
rect 70094 13119 70152 13165
rect 70198 13119 70256 13165
rect 70302 13119 70360 13165
rect 70406 13119 70464 13165
rect 70510 13119 70568 13165
rect 70614 13119 70672 13165
rect 70718 13119 70776 13165
rect 70822 13119 70880 13165
rect 70926 13119 71000 13165
rect 44848 13108 71000 13119
<< metal2 >>
rect 70584 68116 70702 68200
rect 70584 66916 70613 68116
rect 70669 66916 70702 68116
rect 70584 60120 70702 66916
rect 70584 58920 70613 60120
rect 70669 58920 70702 60120
rect 70584 56910 70702 58920
rect 70584 55710 70613 56910
rect 70669 55710 70702 56910
rect 70584 55302 70702 55710
rect 70584 54102 70613 55302
rect 70669 54102 70702 55302
rect 70584 53722 70702 54102
rect 70584 52522 70613 53722
rect 70669 52522 70702 53722
rect 70584 45739 70702 52522
rect 70584 42875 70613 45739
rect 70669 42875 70702 45739
rect 70584 42497 70702 42875
rect 70584 41297 70613 42497
rect 70669 41297 70702 42497
rect 70584 39332 70702 41297
rect 70584 36468 70613 39332
rect 70669 36468 70702 39332
rect 70584 36132 70702 36468
rect 70584 33268 70613 36132
rect 70669 33268 70702 36132
rect 70584 32920 70702 33268
rect 70584 30056 70613 32920
rect 70669 30056 70702 32920
rect 70584 29752 70702 30056
rect 70584 26888 70613 29752
rect 70669 26888 70702 29752
rect 70584 24906 70702 26888
rect 70584 23706 70613 24906
rect 70669 23706 70702 24906
rect 70584 23599 70702 23706
<< via2 >>
rect 70613 66916 70669 68116
rect 70613 58920 70669 60120
rect 70613 55710 70669 56910
rect 70613 54102 70669 55302
rect 70613 52522 70669 53722
rect 70613 42875 70669 45739
rect 70613 41297 70669 42497
rect 70613 36468 70669 39332
rect 70613 33268 70669 36132
rect 70613 30056 70669 32920
rect 70613 26888 70669 29752
rect 70613 23706 70669 24906
<< metal3 >>
rect 14000 47020 17000 71000
rect 17200 48366 20200 71000
rect 20400 49973 23400 71000
rect 23600 50451 25000 71000
rect 25200 51120 26600 71000
rect 26800 52360 29800 71000
rect 30000 53704 33000 71000
rect 33200 55027 36200 71000
rect 36400 56664 39400 71000
rect 39600 57138 41000 71000
rect 41200 57810 42600 71000
rect 42800 59040 45800 71000
rect 46000 60708 49000 71000
rect 49200 61175 50600 71000
rect 50800 61839 52200 71000
rect 52400 62507 53800 71000
rect 54000 63320 55400 71000
rect 55600 63836 57000 71000
rect 57200 64540 58600 71000
rect 58800 65166 60200 71000
rect 60400 65831 61800 71000
rect 62000 66494 63400 71000
rect 63600 67166 65000 71000
rect 65200 67829 66600 71000
rect 66800 68493 68200 71000
rect 68400 69678 69678 71000
rect 68400 68769 71000 69678
tri 68200 68493 68400 68693 sw
tri 68400 68493 68676 68769 ne
rect 68676 68493 71000 68769
rect 66800 68400 68400 68493
tri 68400 68400 68493 68493 sw
tri 68676 68400 68769 68493 ne
rect 68769 68400 71000 68493
rect 66800 68200 68493 68400
tri 68493 68200 68693 68400 sw
rect 66800 68116 71000 68200
rect 66800 68113 70613 68116
tri 66800 68029 66884 68113 ne
rect 66884 68029 70613 68113
tri 66600 67829 66800 68029 sw
tri 66884 67829 67084 68029 ne
rect 67084 67829 70613 68029
rect 65200 67650 66800 67829
tri 66800 67650 66979 67829 sw
tri 67084 67650 67263 67829 ne
rect 67263 67650 70613 67829
rect 65200 67449 66979 67650
tri 65200 67366 65283 67449 ne
rect 65283 67366 66979 67449
tri 66979 67366 67263 67650 sw
tri 67263 67366 67547 67650 ne
rect 67547 67366 70613 67650
tri 65000 67166 65200 67366 sw
tri 65283 67166 65483 67366 ne
rect 65483 67264 67263 67366
tri 67263 67264 67365 67366 sw
tri 67547 67264 67649 67366 ne
rect 67649 67264 70613 67366
rect 65483 67166 67365 67264
rect 63600 66980 65200 67166
tri 65200 66980 65386 67166 sw
tri 65483 66980 65669 67166 ne
rect 65669 66980 67365 67166
tri 67365 66980 67649 67264 sw
tri 67649 66980 67933 67264 ne
rect 67933 66980 70613 67264
rect 63600 66906 65386 66980
tri 65386 66906 65460 66980 sw
tri 65669 66906 65743 66980 ne
rect 65743 66906 67649 66980
tri 67649 66906 67723 66980 sw
tri 67933 66906 68007 66980 ne
rect 68007 66916 70613 66980
rect 70669 66916 71000 68116
rect 68007 66906 71000 66916
rect 63600 66786 65460 66906
tri 63600 66694 63692 66786 ne
rect 63692 66694 65460 66786
tri 65460 66694 65672 66906 sw
tri 65743 66694 65955 66906 ne
rect 65955 66800 67723 66906
tri 67723 66800 67829 66906 sw
tri 68007 66800 68113 66906 ne
rect 68113 66800 71000 66906
rect 65955 66694 67829 66800
tri 67829 66694 67935 66800 sw
tri 63400 66494 63600 66694 sw
tri 63692 66494 63892 66694 ne
rect 63892 66494 65672 66694
rect 62000 66323 63600 66494
tri 63600 66323 63771 66494 sw
tri 63892 66323 64063 66494 ne
rect 64063 66411 65672 66494
tri 65672 66411 65955 66694 sw
tri 65955 66411 66238 66694 ne
rect 66238 66600 67935 66694
tri 67935 66600 68029 66694 sw
rect 66238 66411 71000 66600
rect 64063 66332 65955 66411
tri 65955 66332 66034 66411 sw
tri 66238 66332 66317 66411 ne
rect 66317 66332 71000 66411
rect 64063 66323 66034 66332
rect 62000 66114 63771 66323
tri 62000 66031 62083 66114 ne
rect 62083 66031 63771 66114
tri 63771 66031 64063 66323 sw
tri 64063 66031 64355 66323 ne
rect 64355 66049 66034 66323
tri 66034 66049 66317 66332 sw
tri 66317 66049 66600 66332 ne
rect 66600 66049 71000 66332
rect 64355 66031 66317 66049
tri 66317 66031 66335 66049 sw
tri 66600 66031 66618 66049 ne
rect 66618 66031 71000 66049
tri 61800 65831 62000 66031 sw
tri 62083 65831 62283 66031 ne
rect 62283 65831 64063 66031
rect 60400 65760 62000 65831
tri 62000 65760 62071 65831 sw
tri 62283 65760 62354 65831 ne
rect 62354 65760 64063 65831
tri 64063 65760 64334 66031 sw
tri 64355 65760 64626 66031 ne
rect 64626 65766 66335 66031
tri 66335 65766 66600 66031 sw
tri 66618 65766 66883 66031 ne
rect 66883 65766 71000 66031
rect 64626 65760 66600 65766
tri 66600 65760 66606 65766 sw
tri 66883 65760 66889 65766 ne
rect 66889 65760 71000 65766
rect 60400 65649 62071 65760
tri 62071 65649 62182 65760 sw
tri 62354 65649 62465 65760 ne
rect 62465 65672 64334 65760
tri 64334 65672 64422 65760 sw
tri 64626 65672 64714 65760 ne
rect 64714 65672 66606 65760
rect 62465 65649 64422 65672
rect 60400 65451 62182 65649
tri 60400 65366 60485 65451 ne
rect 60485 65366 62182 65451
tri 62182 65366 62465 65649 sw
tri 62465 65380 62734 65649 ne
rect 62734 65380 64422 65649
tri 64422 65380 64714 65672 sw
tri 64714 65380 65006 65672 ne
rect 65006 65663 66606 65672
tri 66606 65663 66703 65760 sw
tri 66889 65663 66986 65760 ne
rect 66986 65663 71000 65760
rect 65006 65380 66703 65663
tri 66703 65380 66986 65663 sw
tri 66986 65380 67269 65663 ne
rect 67269 65380 71000 65663
tri 62734 65366 62748 65380 ne
rect 62748 65366 64714 65380
tri 64714 65366 64728 65380 sw
tri 65006 65366 65020 65380 ne
rect 65020 65366 66986 65380
tri 66986 65366 67000 65380 sw
tri 67269 65366 67283 65380 ne
rect 67283 65366 71000 65380
tri 60200 65166 60400 65366 sw
tri 60485 65166 60685 65366 ne
rect 60685 65166 62465 65366
rect 58800 64984 60400 65166
tri 60400 64984 60582 65166 sw
tri 60685 64984 60867 65166 ne
rect 60867 65083 62465 65166
tri 62465 65083 62748 65366 sw
tri 62748 65083 63031 65366 ne
rect 63031 65292 64728 65366
tri 64728 65292 64802 65366 sw
tri 65020 65292 65094 65366 ne
rect 65094 65292 67000 65366
rect 63031 65083 64802 65292
rect 60867 64997 62748 65083
tri 62748 64997 62834 65083 sw
tri 63031 64997 63117 65083 ne
rect 63117 65000 64802 65083
tri 64802 65000 65094 65292 sw
tri 65094 65000 65386 65292 ne
rect 65386 65200 67000 65292
tri 67000 65200 67166 65366 sw
tri 67283 65200 67449 65366 ne
rect 67449 65200 71000 65366
rect 65386 65000 67166 65200
tri 67166 65000 67366 65200 sw
rect 63117 64997 65094 65000
rect 60867 64984 62834 64997
rect 58800 64786 60582 64984
tri 58800 64699 58887 64786 ne
rect 58887 64699 60582 64786
tri 60582 64699 60867 64984 sw
tri 60867 64699 61152 64984 ne
rect 61152 64714 62834 64984
tri 62834 64714 63117 64997 sw
tri 63117 64714 63400 64997 ne
rect 63400 64714 65094 64997
rect 61152 64699 63117 64714
tri 63117 64699 63132 64714 sw
tri 63400 64699 63415 64714 ne
rect 63415 64708 65094 64714
tri 65094 64708 65386 65000 sw
tri 65386 64708 65678 65000 ne
rect 65678 64708 71000 65000
rect 63415 64699 65386 64708
tri 65386 64699 65395 64708 sw
tri 65678 64699 65687 64708 ne
rect 65687 64699 71000 64708
tri 58600 64540 58759 64699 sw
tri 58887 64540 59046 64699 ne
rect 59046 64540 60867 64699
tri 60867 64540 61026 64699 sw
tri 61152 64540 61311 64699 ne
rect 61311 64540 63132 64699
tri 63132 64540 63291 64699 sw
tri 63415 64540 63574 64699 ne
rect 63574 64540 65395 64699
tri 65395 64540 65554 64699 sw
tri 65687 64540 65846 64699 ne
rect 65846 64540 71000 64699
rect 57200 64499 58759 64540
tri 58759 64499 58800 64540 sw
tri 59046 64499 59087 64540 ne
rect 59087 64499 61026 64540
rect 57200 64323 58800 64499
tri 58800 64323 58976 64499 sw
tri 59087 64323 59263 64499 ne
rect 59263 64445 61026 64499
tri 61026 64445 61121 64540 sw
tri 61311 64445 61406 64540 ne
rect 61406 64445 63291 64540
rect 59263 64323 61121 64445
rect 57200 64119 58976 64323
tri 57200 64036 57283 64119 ne
rect 57283 64036 58976 64119
tri 58976 64036 59263 64323 sw
tri 59263 64160 59426 64323 ne
rect 59426 64160 61121 64323
tri 61121 64160 61406 64445 sw
tri 61406 64160 61691 64445 ne
rect 61691 64431 63291 64445
tri 63291 64431 63400 64540 sw
tri 63574 64431 63683 64540 ne
rect 63683 64452 65554 64540
tri 65554 64452 65642 64540 sw
tri 65846 64452 65934 64540 ne
rect 65934 64452 71000 64540
rect 63683 64431 65642 64452
rect 61691 64160 63400 64431
tri 63400 64160 63671 64431 sw
tri 63683 64160 63954 64431 ne
rect 63954 64160 65642 64431
tri 65642 64160 65934 64452 sw
tri 65934 64160 66226 64452 ne
rect 66226 64160 71000 64452
tri 59426 64036 59550 64160 ne
rect 59550 64036 61406 64160
tri 61406 64036 61530 64160 sw
tri 61691 64036 61815 64160 ne
rect 61815 64036 63671 64160
tri 63671 64036 63795 64160 sw
tri 63954 64036 64078 64160 ne
rect 64078 64036 65934 64160
tri 65934 64036 66058 64160 sw
tri 66226 64036 66350 64160 ne
rect 66350 64036 71000 64160
tri 57000 63836 57200 64036 sw
tri 57283 63836 57483 64036 ne
rect 57483 63836 59263 64036
rect 55600 63656 57200 63836
tri 57200 63656 57380 63836 sw
tri 57483 63656 57663 63836 ne
rect 57663 63749 59263 63836
tri 59263 63749 59550 64036 sw
tri 59550 63749 59837 64036 ne
rect 59837 63780 61530 64036
tri 61530 63780 61786 64036 sw
tri 61815 63780 62071 64036 ne
rect 62071 63780 63795 64036
tri 63795 63780 64051 64036 sw
tri 64078 63780 64334 64036 ne
rect 64334 63780 66058 64036
tri 66058 63780 66314 64036 sw
tri 66350 63780 66606 64036 ne
rect 66606 63780 71000 64036
rect 59837 63749 61786 63780
rect 57663 63673 59550 63749
tri 59550 63673 59626 63749 sw
tri 59837 63673 59913 63749 ne
rect 59913 63673 61786 63749
rect 57663 63656 59626 63673
rect 55600 63456 57380 63656
tri 55600 63373 55683 63456 ne
rect 55683 63373 57380 63456
tri 57380 63373 57663 63656 sw
tri 57663 63373 57946 63656 ne
rect 57946 63386 59626 63656
tri 59626 63386 59913 63673 sw
tri 59913 63386 60200 63673 ne
rect 60200 63495 61786 63673
tri 61786 63495 62071 63780 sw
tri 62071 63495 62356 63780 ne
rect 62356 63683 64051 63780
tri 64051 63683 64148 63780 sw
tri 64334 63683 64431 63780 ne
rect 64431 63683 66314 63780
rect 62356 63495 64148 63683
rect 60200 63386 62071 63495
rect 57946 63373 59913 63386
tri 59913 63373 59926 63386 sw
tri 60200 63373 60213 63386 ne
rect 60213 63373 62071 63386
tri 62071 63373 62193 63495 sw
tri 62356 63373 62478 63495 ne
rect 62478 63400 64148 63495
tri 64148 63400 64431 63683 sw
tri 64431 63400 64714 63683 ne
rect 64714 63600 66314 63683
tri 66314 63600 66494 63780 sw
tri 66606 63600 66786 63780 ne
rect 66786 63600 71000 63780
rect 64714 63400 66494 63600
tri 66494 63400 66694 63600 sw
rect 62478 63373 64431 63400
tri 64431 63373 64458 63400 sw
tri 64714 63373 64741 63400 ne
rect 64741 63373 71000 63400
tri 55400 63320 55453 63373 sw
tri 55683 63320 55736 63373 ne
rect 55736 63320 57663 63373
tri 57663 63320 57716 63373 sw
tri 57946 63320 57999 63373 ne
rect 57999 63320 59926 63373
tri 59926 63320 59979 63373 sw
tri 60213 63320 60266 63373 ne
rect 60266 63320 62193 63373
tri 62193 63320 62246 63373 sw
tri 62478 63320 62531 63373 ne
rect 62531 63320 64458 63373
tri 64458 63320 64511 63373 sw
tri 64741 63320 64794 63373 ne
rect 64794 63320 71000 63373
rect 54000 63173 55453 63320
tri 55453 63173 55600 63320 sw
tri 55736 63173 55883 63320 ne
rect 55883 63223 57716 63320
tri 57716 63223 57813 63320 sw
tri 57999 63223 58096 63320 ne
rect 58096 63223 59979 63320
rect 55883 63173 57813 63223
rect 54000 62990 55600 63173
tri 55600 62990 55783 63173 sw
tri 55883 62990 56066 63173 ne
rect 56066 62990 57813 63173
rect 54000 62793 55783 62990
tri 54000 62707 54086 62793 ne
rect 54086 62707 55783 62793
tri 55783 62707 56066 62990 sw
tri 56066 62940 56116 62990 ne
rect 56116 62940 57813 62990
tri 57813 62940 58096 63223 sw
tri 58096 62940 58379 63223 ne
rect 58379 63099 59979 63223
tri 59979 63099 60200 63320 sw
tri 60266 63099 60487 63320 ne
rect 60487 63225 62246 63320
tri 62246 63225 62341 63320 sw
tri 62531 63225 62626 63320 ne
rect 62626 63225 64511 63320
rect 60487 63099 62341 63225
rect 58379 62940 60200 63099
tri 60200 62940 60359 63099 sw
tri 60487 62940 60646 63099 ne
rect 60646 62940 62341 63099
tri 62341 62940 62626 63225 sw
tri 62626 62940 62911 63225 ne
rect 62911 63117 64511 63225
tri 64511 63117 64714 63320 sw
tri 64794 63117 64997 63320 ne
rect 64997 63117 71000 63320
rect 62911 62940 64714 63117
tri 64714 62940 64891 63117 sw
tri 64997 62940 65174 63117 ne
rect 65174 62940 71000 63117
tri 56116 62707 56349 62940 ne
rect 56349 62707 58096 62940
tri 58096 62707 58329 62940 sw
tri 58379 62707 58612 62940 ne
rect 58612 62707 60359 62940
tri 60359 62707 60592 62940 sw
tri 60646 62707 60879 62940 ne
rect 60879 62707 62626 62940
tri 62626 62707 62859 62940 sw
tri 62911 62707 63144 62940 ne
rect 63144 62707 64891 62940
tri 64891 62707 65124 62940 sw
tri 65174 62707 65407 62940 ne
rect 65407 62707 71000 62940
tri 53800 62507 54000 62707 sw
tri 54086 62507 54286 62707 ne
rect 54286 62507 56066 62707
rect 52400 62325 54000 62507
tri 54000 62325 54182 62507 sw
tri 54286 62325 54468 62507 ne
rect 54468 62424 56066 62507
tri 56066 62424 56349 62707 sw
tri 56349 62424 56632 62707 ne
rect 56632 62560 58329 62707
tri 58329 62560 58476 62707 sw
tri 58612 62560 58759 62707 ne
rect 58759 62560 60592 62707
tri 60592 62560 60739 62707 sw
tri 60879 62560 61026 62707 ne
rect 61026 62560 62859 62707
tri 62859 62560 63006 62707 sw
tri 63144 62560 63291 62707 ne
rect 63291 62560 65124 62707
tri 65124 62560 65271 62707 sw
tri 65407 62560 65554 62707 ne
rect 65554 62560 71000 62707
rect 56632 62424 58476 62560
rect 54468 62339 56349 62424
tri 56349 62339 56434 62424 sw
tri 56632 62339 56717 62424 ne
rect 56717 62339 58476 62424
rect 54468 62325 56434 62339
rect 52400 62127 54182 62325
tri 52400 62039 52488 62127 ne
rect 52488 62039 54182 62127
tri 54182 62039 54468 62325 sw
tri 54468 62039 54754 62325 ne
rect 54754 62056 56434 62325
tri 56434 62056 56717 62339 sw
tri 56717 62056 57000 62339 ne
rect 57000 62277 58476 62339
tri 58476 62277 58759 62560 sw
tri 58759 62277 59042 62560 ne
rect 59042 62467 60739 62560
tri 60739 62467 60832 62560 sw
tri 61026 62467 61119 62560 ne
rect 61119 62467 63006 62560
rect 59042 62277 60832 62467
rect 57000 62056 58759 62277
rect 54754 62039 56717 62056
tri 56717 62039 56734 62056 sw
tri 57000 62039 57017 62056 ne
rect 57017 62039 58759 62056
tri 58759 62039 58997 62277 sw
tri 59042 62039 59280 62277 ne
rect 59280 62180 60832 62277
tri 60832 62180 61119 62467 sw
tri 61119 62180 61406 62467 ne
rect 61406 62465 63006 62467
tri 63006 62465 63101 62560 sw
tri 63291 62465 63386 62560 ne
rect 63386 62465 65271 62560
rect 61406 62180 63101 62465
tri 63101 62180 63386 62465 sw
tri 63386 62180 63671 62465 ne
rect 63671 62463 65271 62465
tri 65271 62463 65368 62560 sw
tri 65554 62463 65651 62560 ne
rect 65651 62463 71000 62560
rect 63671 62180 65368 62463
tri 65368 62180 65651 62463 sw
tri 65651 62180 65934 62463 ne
rect 65934 62180 71000 62463
rect 59280 62039 61119 62180
tri 61119 62039 61260 62180 sw
tri 61406 62039 61547 62180 ne
rect 61547 62039 63386 62180
tri 63386 62039 63527 62180 sw
tri 63671 62039 63812 62180 ne
rect 63812 62039 65651 62180
tri 65651 62039 65792 62180 sw
tri 65934 62039 66075 62180 ne
rect 66075 62039 71000 62180
tri 52200 61839 52400 62039 sw
tri 52488 61839 52688 62039 ne
rect 52688 62006 54468 62039
tri 54468 62006 54501 62039 sw
tri 54754 62006 54787 62039 ne
rect 54787 62006 56734 62039
rect 52688 61839 54501 62006
rect 50800 61663 52400 61839
tri 52400 61663 52576 61839 sw
tri 52688 61663 52864 61839 ne
rect 52864 61720 54501 61839
tri 54501 61720 54787 62006 sw
tri 54787 61720 55073 62006 ne
rect 55073 61773 56734 62006
tri 56734 61773 57000 62039 sw
tri 57017 61773 57283 62039 ne
rect 57283 62003 58997 62039
tri 58997 62003 59033 62039 sw
tri 59280 62003 59316 62039 ne
rect 59316 62003 61260 62039
rect 57283 61773 59033 62003
rect 55073 61720 57000 61773
tri 57000 61720 57053 61773 sw
tri 57283 61720 57336 61773 ne
rect 57336 61720 59033 61773
tri 59033 61720 59316 62003 sw
tri 59316 61720 59599 62003 ne
rect 59599 61893 61260 62003
tri 61260 61893 61406 62039 sw
tri 61547 61893 61693 62039 ne
rect 61693 61893 63527 62039
rect 59599 61720 61406 61893
tri 61406 61720 61579 61893 sw
tri 61693 61720 61866 61893 ne
rect 61866 61800 63527 61893
tri 63527 61800 63766 62039 sw
tri 63812 61800 64051 62039 ne
rect 64051 62000 65792 62039
tri 65792 62000 65831 62039 sw
tri 66075 62000 66114 62039 ne
rect 66114 62000 71000 62039
rect 64051 61800 65831 62000
tri 65831 61800 66031 62000 sw
rect 61866 61720 63766 61800
tri 63766 61720 63846 61800 sw
tri 64051 61720 64131 61800 ne
rect 64131 61720 71000 61800
rect 52864 61663 54787 61720
rect 50800 61459 52576 61663
tri 50800 61375 50884 61459 ne
rect 50884 61375 52576 61459
tri 52576 61375 52864 61663 sw
tri 52864 61375 53152 61663 ne
rect 53152 61661 54787 61663
tri 54787 61661 54846 61720 sw
tri 55073 61661 55132 61720 ne
rect 55132 61661 57053 61720
rect 53152 61375 54846 61661
tri 54846 61375 55132 61661 sw
tri 55132 61375 55418 61661 ne
rect 55418 61658 57053 61661
tri 57053 61658 57115 61720 sw
tri 57336 61658 57398 61720 ne
rect 57398 61658 59316 61720
tri 59316 61658 59378 61720 sw
tri 59599 61658 59661 61720 ne
rect 59661 61662 61579 61720
tri 61579 61662 61637 61720 sw
tri 61866 61662 61924 61720 ne
rect 61924 61662 63846 61720
rect 59661 61658 61637 61662
rect 55418 61375 57115 61658
tri 57115 61375 57398 61658 sw
tri 57398 61375 57681 61658 ne
rect 57681 61375 59378 61658
tri 59378 61375 59661 61658 sw
tri 59661 61375 59944 61658 ne
rect 59944 61375 61637 61658
tri 61637 61375 61924 61662 sw
tri 61924 61375 62211 61662 ne
rect 62211 61515 63846 61662
tri 63846 61515 64051 61720 sw
tri 64131 61515 64336 61720 ne
rect 64336 61515 71000 61720
rect 62211 61375 64051 61515
tri 64051 61375 64191 61515 sw
tri 64336 61375 64476 61515 ne
rect 64476 61375 71000 61515
tri 50600 61175 50800 61375 sw
tri 50884 61175 51084 61375 ne
rect 51084 61175 52864 61375
rect 49200 60992 50800 61175
tri 50800 60992 50983 61175 sw
tri 51084 60992 51267 61175 ne
rect 51267 61087 52864 61175
tri 52864 61087 53152 61375 sw
tri 53152 61087 53440 61375 ne
rect 53440 61340 55132 61375
tri 55132 61340 55167 61375 sw
tri 55418 61340 55453 61375 ne
rect 55453 61340 57398 61375
tri 57398 61340 57433 61375 sw
tri 57681 61340 57716 61375 ne
rect 57716 61340 59661 61375
tri 59661 61340 59696 61375 sw
tri 59944 61340 59979 61375 ne
rect 59979 61340 61924 61375
tri 61924 61340 61959 61375 sw
tri 62211 61340 62246 61375 ne
rect 62246 61340 64191 61375
tri 64191 61340 64226 61375 sw
tri 64476 61340 64511 61375 ne
rect 64511 61340 71000 61375
rect 53440 61087 55167 61340
rect 51267 61015 53152 61087
tri 53152 61015 53224 61087 sw
tri 53440 61015 53512 61087 ne
rect 53512 61054 55167 61087
tri 55167 61054 55453 61340 sw
tri 55453 61054 55739 61340 ne
rect 55739 61243 57433 61340
tri 57433 61243 57530 61340 sw
tri 57716 61243 57813 61340 ne
rect 57813 61243 59696 61340
tri 59696 61243 59793 61340 sw
tri 59979 61243 60076 61340 ne
rect 60076 61247 61959 61340
tri 61959 61247 62052 61340 sw
tri 62246 61247 62339 61340 ne
rect 62339 61247 64226 61340
rect 60076 61243 62052 61247
rect 55739 61054 57530 61243
rect 53512 61015 55453 61054
rect 51267 60992 53224 61015
rect 49200 60795 50983 60992
tri 49000 60708 49002 60710 sw
tri 49200 60708 49287 60795 ne
rect 49287 60708 50983 60795
tri 50983 60708 51267 60992 sw
tri 51267 60708 51551 60992 ne
rect 51551 60727 53224 60992
tri 53224 60727 53512 61015 sw
tri 53512 60727 53800 61015 ne
rect 53800 60994 55453 61015
tri 55453 60994 55513 61054 sw
tri 55739 60994 55799 61054 ne
rect 55799 60994 57530 61054
rect 53800 60727 55513 60994
rect 51551 60708 53512 60727
tri 53512 60708 53531 60727 sw
tri 53800 60708 53819 60727 ne
rect 53819 60708 55513 60727
tri 55513 60708 55799 60994 sw
tri 55799 60708 56085 60994 ne
rect 56085 60960 57530 60994
tri 57530 60960 57813 61243 sw
tri 57813 60960 58096 61243 ne
rect 58096 60960 59793 61243
tri 59793 60960 60076 61243 sw
tri 60076 60960 60359 61243 ne
rect 60359 60960 62052 61243
tri 62052 60960 62339 61247 sw
tri 62339 60960 62626 61247 ne
rect 62626 61245 64226 61247
tri 64226 61245 64321 61340 sw
tri 64511 61245 64606 61340 ne
rect 64606 61245 71000 61340
rect 62626 60960 64321 61245
tri 64321 60960 64606 61245 sw
tri 64606 60960 64891 61245 ne
rect 64891 60960 71000 61245
rect 56085 60708 57813 60960
tri 57813 60708 58065 60960 sw
tri 58096 60708 58348 60960 ne
rect 58348 60708 60076 60960
tri 60076 60708 60328 60960 sw
tri 60359 60708 60611 60960 ne
rect 60611 60708 62339 60960
tri 62339 60708 62591 60960 sw
tri 62626 60708 62878 60960 ne
rect 62878 60708 64606 60960
tri 64606 60708 64858 60960 sw
tri 64891 60708 65143 60960 ne
rect 65143 60708 71000 60960
rect 46000 60423 49002 60708
tri 49002 60423 49287 60708 sw
tri 49287 60508 49487 60708 ne
rect 49487 60508 51267 60708
rect 46000 60224 49287 60423
tri 49287 60224 49486 60423 sw
tri 49487 60417 49578 60508 ne
rect 49578 60500 51267 60508
tri 51267 60500 51475 60708 sw
tri 51551 60500 51759 60708 ne
rect 51759 60500 53531 60708
tri 53531 60500 53739 60708 sw
tri 53819 60500 54027 60708 ne
rect 54027 60500 55799 60708
tri 55799 60500 56007 60708 sw
tri 56085 60500 56293 60708 ne
rect 56293 60677 58065 60708
tri 58065 60677 58096 60708 sw
tri 58348 60677 58379 60708 ne
rect 58379 60677 60328 60708
rect 56293 60500 58096 60677
tri 58096 60500 58273 60677 sw
tri 58379 60500 58556 60677 ne
rect 58556 60580 60328 60677
tri 60328 60580 60456 60708 sw
tri 60611 60580 60739 60708 ne
rect 60739 60580 62591 60708
tri 62591 60580 62719 60708 sw
tri 62878 60580 63006 60708 ne
rect 63006 60580 64858 60708
tri 64858 60580 64986 60708 sw
tri 65143 60580 65271 60708 ne
rect 65271 60580 71000 60708
rect 58556 60500 60456 60580
tri 60456 60500 60536 60580 sw
tri 60739 60500 60819 60580 ne
rect 60819 60500 62719 60580
tri 62719 60500 62799 60580 sw
tri 63006 60500 63086 60580 ne
rect 63086 60500 64986 60580
tri 64986 60500 65066 60580 sw
tri 65271 60500 65351 60580 ne
rect 65351 60500 71000 60580
rect 49578 60417 51475 60500
rect 46000 60132 49486 60224
tri 49486 60132 49578 60224 sw
tri 49578 60132 49863 60417 ne
rect 49863 60414 51475 60417
tri 51475 60414 51561 60500 sw
tri 51759 60414 51845 60500 ne
rect 51845 60439 53739 60500
tri 53739 60439 53800 60500 sw
tri 54027 60439 54088 60500 ne
rect 54088 60439 56007 60500
rect 51845 60418 53800 60439
tri 53800 60418 53821 60439 sw
tri 54088 60418 54109 60439 ne
rect 54109 60418 56007 60439
rect 51845 60414 53821 60418
rect 49863 60132 51561 60414
rect 46000 59847 49578 60132
tri 49578 59847 49863 60132 sw
tri 49863 60130 49865 60132 ne
rect 49865 60130 51561 60132
tri 51561 60130 51845 60414 sw
tri 51845 60130 52129 60414 ne
rect 52129 60130 53821 60414
tri 53821 60130 54109 60418 sw
tri 54109 60130 54397 60418 ne
rect 54397 60416 56007 60418
tri 56007 60416 56091 60500 sw
tri 56293 60416 56377 60500 ne
rect 56377 60416 58273 60500
rect 54397 60130 56091 60416
tri 56091 60130 56377 60416 sw
tri 56377 60130 56663 60416 ne
rect 56663 60413 58273 60416
tri 58273 60413 58360 60500 sw
tri 58556 60413 58643 60500 ne
rect 58643 60413 60536 60500
rect 56663 60130 58360 60413
tri 58360 60130 58643 60413 sw
tri 58643 60130 58926 60413 ne
rect 58926 60297 60536 60413
tri 60536 60297 60739 60500 sw
tri 60819 60297 61022 60500 ne
rect 61022 60487 62799 60500
tri 62799 60487 62812 60500 sw
tri 63086 60487 63099 60500 ne
rect 63099 60487 65066 60500
rect 61022 60297 62812 60487
rect 58926 60130 60739 60297
tri 60739 60130 60906 60297 sw
tri 61022 60130 61189 60297 ne
rect 61189 60200 62812 60297
tri 62812 60200 63099 60487 sw
tri 63099 60200 63386 60487 ne
rect 63386 60400 65066 60487
tri 65066 60400 65166 60500 sw
tri 65351 60400 65451 60500 ne
rect 65451 60400 71000 60500
rect 63386 60200 65166 60400
tri 65166 60200 65366 60400 sw
rect 61189 60130 63099 60200
tri 63099 60130 63169 60200 sw
tri 63386 60130 63456 60200 ne
rect 63456 60130 71000 60200
rect 46000 59845 49863 59847
tri 49863 59845 49865 59847 sw
tri 49865 59845 50150 60130 ne
rect 50150 60120 51845 60130
tri 51845 60120 51855 60130 sw
tri 52129 60120 52139 60130 ne
rect 52139 60120 54109 60130
tri 54109 60120 54119 60130 sw
tri 54397 60120 54407 60130 ne
rect 54407 60120 56377 60130
tri 56377 60120 56387 60130 sw
tri 56663 60120 56673 60130 ne
rect 56673 60120 58643 60130
tri 58643 60120 58653 60130 sw
tri 58926 60120 58936 60130 ne
rect 58936 60120 60906 60130
tri 60906 60120 60916 60130 sw
tri 61189 60120 61199 60130 ne
rect 61199 60120 63169 60130
tri 63169 60120 63179 60130 sw
tri 63456 60120 63466 60130 ne
rect 63466 60120 71000 60130
rect 50150 60059 51855 60120
tri 51855 60059 51916 60120 sw
tri 52139 60059 52200 60120 ne
rect 52200 60059 54119 60120
rect 50150 59845 51916 60059
rect 46000 59561 49865 59845
tri 49865 59561 50149 59845 sw
tri 50150 59682 50313 59845 ne
rect 50313 59775 51916 59845
tri 51916 59775 52200 60059 sw
tri 52200 59775 52484 60059 ne
rect 52484 60028 54119 60059
tri 54119 60028 54211 60120 sw
tri 54407 60028 54499 60120 ne
rect 54499 60028 56387 60120
rect 52484 59775 54211 60028
rect 50313 59682 52200 59775
rect 46000 59461 50149 59561
tri 46000 59350 46111 59461 ne
rect 46111 59397 50149 59461
tri 50149 59397 50313 59561 sw
tri 50313 59461 50534 59682 ne
rect 50534 59624 52200 59682
tri 52200 59624 52351 59775 sw
tri 52484 59624 52635 59775 ne
rect 52635 59740 54211 59775
tri 54211 59740 54499 60028 sw
tri 54499 59740 54787 60028 ne
rect 54787 60026 56387 60028
tri 56387 60026 56481 60120 sw
tri 56673 60026 56767 60120 ne
rect 56767 60026 58653 60120
rect 54787 59740 56481 60026
tri 56481 59740 56767 60026 sw
tri 56767 59740 57053 60026 ne
rect 57053 60023 58653 60026
tri 58653 60023 58750 60120 sw
tri 58936 60023 59033 60120 ne
rect 59033 60023 60916 60120
tri 60916 60023 61013 60120 sw
tri 61199 60023 61296 60120 ne
rect 61296 60023 63179 60120
rect 57053 59740 58750 60023
tri 58750 59740 59033 60023 sw
tri 59033 59740 59316 60023 ne
rect 59316 59740 61013 60023
tri 61013 59740 61296 60023 sw
tri 61296 59740 61579 60023 ne
rect 61579 59913 63179 60023
tri 63179 59913 63386 60120 sw
tri 63466 59913 63673 60120 ne
rect 63673 59913 70613 60120
rect 61579 59740 63386 59913
tri 63386 59740 63559 59913 sw
tri 63673 59740 63846 59913 ne
rect 63846 59740 70613 59913
rect 52635 59624 54499 59740
rect 50534 59461 52351 59624
rect 46111 59350 50313 59397
tri 45800 59040 46110 59350 sw
tri 46111 59140 46321 59350 ne
rect 46321 59176 50313 59350
tri 50313 59176 50534 59397 sw
tri 50534 59340 50655 59461 ne
rect 50655 59340 52351 59461
tri 52351 59340 52635 59624 sw
tri 52635 59340 52919 59624 ne
rect 52919 59452 54499 59624
tri 54499 59452 54787 59740 sw
tri 54787 59452 55075 59740 ne
rect 55075 59646 56767 59740
tri 56767 59646 56861 59740 sw
tri 57053 59646 57147 59740 ne
rect 57147 59646 59033 59740
rect 55075 59452 56861 59646
rect 52919 59340 54787 59452
tri 54787 59340 54899 59452 sw
tri 55075 59340 55187 59452 ne
rect 55187 59360 56861 59452
tri 56861 59360 57147 59646 sw
tri 57147 59360 57433 59646 ne
rect 57433 59643 59033 59646
tri 59033 59643 59130 59740 sw
tri 59316 59643 59413 59740 ne
rect 59413 59643 61296 59740
tri 61296 59643 61393 59740 sw
tri 61579 59643 61676 59740 ne
rect 61676 59647 63559 59740
tri 63559 59647 63652 59740 sw
tri 63846 59647 63939 59740 ne
rect 63939 59647 70613 59740
rect 61676 59643 63652 59647
rect 57433 59360 59130 59643
tri 59130 59360 59413 59643 sw
tri 59413 59360 59696 59643 ne
rect 59696 59360 61393 59643
tri 61393 59360 61676 59643 sw
tri 61676 59360 61959 59643 ne
rect 61959 59360 63652 59643
tri 63652 59360 63939 59647 sw
tri 63939 59360 64226 59647 ne
rect 64226 59360 70613 59647
rect 55187 59340 57147 59360
tri 57147 59340 57167 59360 sw
tri 57433 59340 57453 59360 ne
rect 57453 59340 59413 59360
tri 59413 59340 59433 59360 sw
tri 59696 59340 59716 59360 ne
rect 59716 59340 61676 59360
tri 61676 59340 61696 59360 sw
tri 61959 59340 61979 59360 ne
rect 61979 59340 63939 59360
tri 63939 59340 63959 59360 sw
tri 64226 59340 64246 59360 ne
rect 64246 59340 70613 59360
rect 46321 59140 50534 59176
rect 42800 58836 46110 59040
tri 46110 58836 46314 59040 sw
tri 46321 58854 46607 59140 ne
rect 46607 59056 50534 59140
tri 50534 59056 50654 59176 sw
tri 50655 59108 50887 59340 ne
rect 50887 59194 52635 59340
tri 52635 59194 52781 59340 sw
tri 52919 59194 53065 59340 ne
rect 53065 59198 54899 59340
tri 54899 59198 55041 59340 sw
tri 55187 59198 55329 59340 ne
rect 55329 59198 57167 59340
rect 53065 59194 55041 59198
rect 50887 59108 52781 59194
rect 46607 58854 50654 59056
rect 42800 58548 46314 58836
tri 46314 58548 46602 58836 sw
tri 46607 58747 46714 58854 ne
rect 46714 58823 50654 58854
tri 50654 58823 50887 59056 sw
tri 50887 58910 51085 59108 ne
rect 51085 58910 52781 59108
tri 52781 58910 53065 59194 sw
tri 53065 58910 53349 59194 ne
rect 53349 58910 55041 59194
tri 55041 58910 55329 59198 sw
tri 55329 58910 55617 59198 ne
rect 55617 59074 57167 59198
tri 57167 59074 57433 59340 sw
tri 57453 59074 57719 59340 ne
rect 57719 59263 59433 59340
tri 59433 59263 59510 59340 sw
tri 59716 59263 59793 59340 ne
rect 59793 59263 61696 59340
tri 61696 59263 61773 59340 sw
tri 61979 59263 62056 59340 ne
rect 62056 59267 63959 59340
tri 63959 59267 64032 59340 sw
tri 64246 59267 64319 59340 ne
rect 64319 59267 70613 59340
rect 62056 59263 64032 59267
rect 57719 59074 59510 59263
rect 55617 58910 57433 59074
tri 57433 58910 57597 59074 sw
tri 57719 58910 57883 59074 ne
rect 57883 58980 59510 59074
tri 59510 58980 59793 59263 sw
tri 59793 58980 60076 59263 ne
rect 60076 58980 61773 59263
tri 61773 58980 62056 59263 sw
tri 62056 58980 62339 59263 ne
rect 62339 58980 64032 59263
tri 64032 58980 64319 59267 sw
tri 64319 58980 64606 59267 ne
rect 64606 58980 70613 59267
rect 57883 58910 59793 58980
tri 59793 58910 59863 58980 sw
tri 60076 58910 60146 58980 ne
rect 60146 58910 62056 58980
tri 62056 58910 62126 58980 sw
tri 62339 58910 62409 58980 ne
rect 62409 58910 64319 58980
tri 64319 58910 64389 58980 sw
tri 64606 58910 64676 58980 ne
rect 64676 58920 70613 58980
rect 70669 58920 71000 60120
rect 64676 58910 71000 58920
rect 46714 58747 50887 58823
rect 42800 58436 46602 58548
tri 46602 58436 46714 58548 sw
tri 46714 58436 47025 58747 ne
rect 47025 58626 50887 58747
tri 50887 58626 51084 58823 sw
tri 51085 58815 51180 58910 ne
rect 51180 58815 53065 58910
tri 51180 58747 51248 58815 ne
rect 51248 58812 53065 58815
tri 53065 58812 53163 58910 sw
tri 53349 58812 53447 58910 ne
rect 53447 58816 55329 58910
tri 55329 58816 55423 58910 sw
tri 55617 58816 55711 58910 ne
rect 55711 58816 57597 58910
rect 53447 58812 55423 58816
rect 51248 58747 53163 58812
rect 47025 58624 51084 58626
tri 51084 58624 51086 58626 sw
rect 47025 58622 51086 58624
tri 51086 58622 51088 58624 sw
rect 47025 58620 51088 58622
tri 51088 58620 51090 58622 sw
rect 47025 58618 51090 58620
tri 51090 58618 51092 58620 sw
rect 47025 58616 51092 58618
tri 51092 58616 51094 58618 sw
rect 47025 58614 51094 58616
tri 51094 58614 51096 58616 sw
rect 47025 58612 51096 58614
tri 51096 58612 51098 58614 sw
rect 47025 58610 51098 58612
tri 51098 58610 51100 58612 sw
rect 47025 58608 51100 58610
tri 51100 58608 51102 58610 sw
rect 47025 58606 51102 58608
tri 51102 58606 51104 58608 sw
rect 47025 58604 51104 58606
tri 51104 58604 51106 58606 sw
rect 47025 58602 51106 58604
tri 51106 58602 51108 58604 sw
rect 47025 58600 51108 58602
tri 51108 58600 51110 58602 sw
rect 47025 58598 51110 58600
tri 51110 58598 51112 58600 sw
rect 47025 58596 51112 58598
tri 51112 58596 51114 58598 sw
rect 47025 58594 51114 58596
tri 51114 58594 51116 58596 sw
rect 47025 58592 51116 58594
tri 51116 58592 51118 58594 sw
rect 47025 58590 51118 58592
tri 51118 58590 51120 58592 sw
rect 47025 58588 51120 58590
tri 51120 58588 51122 58590 sw
rect 47025 58586 51122 58588
tri 51122 58586 51124 58588 sw
rect 47025 58584 51124 58586
tri 51124 58584 51126 58586 sw
rect 47025 58582 51126 58584
tri 51126 58582 51128 58584 sw
rect 47025 58580 51128 58582
tri 51128 58580 51130 58582 sw
rect 47025 58578 51130 58580
tri 51130 58578 51132 58580 sw
rect 47025 58576 51132 58578
tri 51132 58576 51134 58578 sw
rect 47025 58574 51134 58576
tri 51134 58574 51136 58576 sw
rect 47025 58572 51136 58574
tri 51136 58572 51138 58574 sw
rect 47025 58570 51138 58572
tri 51138 58570 51140 58572 sw
rect 47025 58568 51140 58570
tri 51140 58568 51142 58570 sw
rect 47025 58566 51142 58568
tri 51142 58566 51144 58568 sw
rect 47025 58564 51144 58566
tri 51144 58564 51146 58566 sw
rect 47025 58562 51146 58564
tri 51146 58562 51148 58564 sw
rect 47025 58560 51148 58562
tri 51148 58560 51150 58562 sw
rect 47025 58558 51150 58560
tri 51150 58558 51152 58560 sw
rect 47025 58556 51152 58558
tri 51152 58556 51154 58558 sw
rect 47025 58554 51154 58556
tri 51154 58554 51156 58556 sw
rect 47025 58552 51156 58554
tri 51156 58552 51158 58554 sw
rect 47025 58550 51158 58552
tri 51158 58550 51160 58552 sw
rect 47025 58548 51160 58550
tri 51160 58548 51162 58550 sw
rect 47025 58546 51162 58548
tri 51162 58546 51164 58548 sw
rect 47025 58544 51164 58546
tri 51164 58544 51166 58546 sw
rect 47025 58542 51166 58544
tri 51166 58542 51168 58544 sw
rect 47025 58540 51168 58542
tri 51168 58540 51170 58542 sw
rect 47025 58538 51170 58540
tri 51170 58538 51172 58540 sw
rect 47025 58536 51172 58538
tri 51172 58536 51174 58538 sw
rect 47025 58534 51174 58536
tri 51174 58534 51176 58536 sw
rect 47025 58532 51176 58534
tri 51176 58532 51178 58534 sw
rect 47025 58530 51178 58532
tri 51178 58530 51180 58532 sw
rect 47025 58528 51180 58530
tri 51180 58528 51182 58530 sw
tri 51248 58528 51467 58747 ne
rect 51467 58528 53163 58747
tri 53163 58528 53447 58812 sw
tri 53447 58528 53731 58812 ne
rect 53731 58528 55423 58812
tri 55423 58528 55711 58816 sw
tri 55711 58528 55999 58816 ne
rect 55999 58814 57597 58816
tri 57597 58814 57693 58910 sw
tri 57883 58814 57979 58910 ne
rect 57979 58814 59863 58910
rect 55999 58528 57693 58814
tri 57693 58528 57979 58814 sw
tri 57979 58528 58265 58814 ne
rect 58265 58697 59863 58814
tri 59863 58697 60076 58910 sw
tri 60146 58697 60359 58910 ne
rect 60359 58883 62126 58910
tri 62126 58883 62153 58910 sw
tri 62409 58883 62436 58910 ne
rect 62436 58883 64389 58910
rect 60359 58697 62153 58883
rect 58265 58528 60076 58697
tri 60076 58528 60245 58697 sw
tri 60359 58528 60528 58697 ne
rect 60528 58600 62153 58697
tri 62153 58600 62436 58883 sw
tri 62436 58600 62719 58883 ne
rect 62719 58800 64389 58883
tri 64389 58800 64499 58910 sw
tri 64676 58800 64786 58910 ne
rect 64786 58800 71000 58910
rect 62719 58600 64499 58800
tri 64499 58600 64699 58800 sw
rect 60528 58528 62436 58600
tri 62436 58528 62508 58600 sw
tri 62719 58528 62791 58600 ne
rect 62791 58528 71000 58600
rect 47025 58436 51182 58528
rect 42800 58127 46714 58436
tri 46714 58127 47023 58436 sw
tri 47025 58331 47130 58436 ne
rect 47130 58331 51182 58436
rect 42800 58097 47023 58127
tri 42600 57810 42800 58010 sw
tri 42800 57810 43087 58097 ne
rect 43087 58020 47023 58097
tri 47023 58020 47130 58127 sw
tri 47130 58097 47364 58331 ne
rect 47364 58243 51182 58331
tri 51182 58243 51467 58528 sw
tri 51467 58520 51475 58528 ne
rect 51475 58520 53447 58528
rect 47364 58241 51467 58243
tri 51467 58241 51469 58243 sw
rect 47364 58239 51469 58241
tri 51469 58239 51471 58241 sw
rect 47364 58237 51471 58239
tri 51471 58237 51473 58239 sw
rect 47364 58235 51473 58237
tri 51473 58235 51475 58237 sw
tri 51475 58235 51760 58520 ne
rect 51760 58424 53447 58520
tri 53447 58424 53551 58528 sw
tri 53731 58424 53835 58528 ne
rect 53835 58520 55711 58528
tri 55711 58520 55719 58528 sw
tri 55999 58520 56007 58528 ne
rect 56007 58520 57979 58528
tri 57979 58520 57987 58528 sw
tri 58265 58520 58273 58528 ne
rect 58273 58520 60245 58528
tri 60245 58520 60253 58528 sw
tri 60528 58520 60536 58528 ne
rect 60536 58520 62508 58528
tri 62508 58520 62516 58528 sw
tri 62791 58520 62799 58528 ne
rect 62799 58520 71000 58528
rect 53835 58428 55719 58520
tri 55719 58428 55811 58520 sw
tri 56007 58428 56099 58520 ne
rect 56099 58428 57987 58520
rect 53835 58424 55811 58428
rect 51760 58235 53551 58424
rect 47364 58097 51475 58235
rect 43087 57810 47130 58020
rect 41200 57625 42800 57810
tri 42800 57625 42985 57810 sw
tri 43087 57625 43272 57810 ne
rect 43272 57793 47130 57810
tri 47130 57793 47357 58020 sw
tri 47364 58005 47456 58097 ne
rect 47456 58005 51475 58097
rect 43272 57694 47357 57793
tri 47357 57694 47456 57793 sw
tri 47456 57694 47767 58005 ne
rect 47767 57950 51475 58005
tri 51475 57950 51760 58235 sw
tri 51760 58010 51985 58235 ne
rect 51985 58140 53551 58235
tri 53551 58140 53835 58424 sw
tri 53835 58140 54119 58424 ne
rect 54119 58140 55811 58424
tri 55811 58140 56099 58428 sw
tri 56099 58140 56387 58428 ne
rect 56387 58426 57987 58428
tri 57987 58426 58081 58520 sw
tri 58273 58426 58367 58520 ne
rect 58367 58426 60253 58520
rect 56387 58140 58081 58426
tri 58081 58140 58367 58426 sw
tri 58367 58140 58653 58426 ne
rect 58653 58423 60253 58426
tri 60253 58423 60350 58520 sw
tri 60536 58423 60633 58520 ne
rect 60633 58423 62516 58520
rect 58653 58140 60350 58423
tri 60350 58140 60633 58423 sw
tri 60633 58140 60916 58423 ne
rect 60916 58317 62516 58423
tri 62516 58317 62719 58520 sw
tri 62799 58317 63002 58520 ne
rect 63002 58317 71000 58520
rect 60916 58140 62719 58317
tri 62719 58140 62896 58317 sw
tri 63002 58140 63179 58317 ne
rect 63179 58140 71000 58317
rect 51985 58010 53835 58140
rect 47767 57948 51760 57950
tri 51760 57948 51762 57950 sw
rect 47767 57946 51762 57948
tri 51762 57946 51764 57948 sw
rect 47767 57944 51764 57946
tri 51764 57944 51766 57946 sw
rect 47767 57942 51766 57944
tri 51766 57942 51768 57944 sw
rect 47767 57940 51768 57942
tri 51768 57940 51770 57942 sw
rect 47767 57938 51770 57940
tri 51770 57938 51772 57940 sw
rect 47767 57936 51772 57938
tri 51772 57936 51774 57938 sw
rect 47767 57934 51774 57936
tri 51774 57934 51776 57936 sw
rect 47767 57932 51776 57934
tri 51776 57932 51778 57934 sw
rect 47767 57930 51778 57932
tri 51778 57930 51780 57932 sw
rect 47767 57928 51780 57930
tri 51780 57928 51782 57930 sw
rect 47767 57926 51782 57928
tri 51782 57926 51784 57928 sw
rect 47767 57924 51784 57926
tri 51784 57924 51786 57926 sw
rect 47767 57922 51786 57924
tri 51786 57922 51788 57924 sw
rect 47767 57920 51788 57922
tri 51788 57920 51790 57922 sw
rect 47767 57918 51790 57920
tri 51790 57918 51792 57920 sw
rect 47767 57916 51792 57918
tri 51792 57916 51794 57918 sw
rect 47767 57914 51794 57916
tri 51794 57914 51796 57916 sw
rect 47767 57912 51796 57914
tri 51796 57912 51798 57914 sw
rect 47767 57910 51798 57912
tri 51798 57910 51800 57912 sw
rect 47767 57908 51800 57910
tri 51800 57908 51802 57910 sw
rect 47767 57906 51802 57908
tri 51802 57906 51804 57908 sw
rect 47767 57904 51804 57906
tri 51804 57904 51806 57906 sw
rect 47767 57902 51806 57904
tri 51806 57902 51808 57904 sw
rect 47767 57900 51808 57902
tri 51808 57900 51810 57902 sw
rect 47767 57898 51810 57900
tri 51810 57898 51812 57900 sw
rect 47767 57896 51812 57898
tri 51812 57896 51814 57898 sw
rect 47767 57894 51814 57896
tri 51814 57894 51816 57896 sw
rect 47767 57892 51816 57894
tri 51816 57892 51818 57894 sw
rect 47767 57890 51818 57892
tri 51818 57890 51820 57892 sw
rect 47767 57888 51820 57890
tri 51820 57888 51822 57890 sw
rect 47767 57886 51822 57888
tri 51822 57886 51824 57888 sw
rect 47767 57884 51824 57886
tri 51824 57884 51826 57886 sw
rect 47767 57882 51826 57884
tri 51826 57882 51828 57884 sw
rect 47767 57880 51828 57882
tri 51828 57880 51830 57882 sw
rect 47767 57878 51830 57880
tri 51830 57878 51832 57880 sw
rect 47767 57876 51832 57878
tri 51832 57876 51834 57878 sw
rect 47767 57874 51834 57876
tri 51834 57874 51836 57876 sw
rect 47767 57872 51836 57874
tri 51836 57872 51838 57874 sw
rect 47767 57870 51838 57872
tri 51838 57870 51840 57872 sw
rect 47767 57868 51840 57870
tri 51840 57868 51842 57870 sw
rect 47767 57866 51842 57868
tri 51842 57866 51844 57868 sw
rect 47767 57864 51844 57866
tri 51844 57864 51846 57866 sw
rect 47767 57862 51846 57864
tri 51846 57862 51848 57864 sw
rect 47767 57860 51848 57862
tri 51848 57860 51850 57862 sw
rect 47767 57858 51850 57860
tri 51850 57858 51852 57860 sw
rect 47767 57856 51852 57858
tri 51852 57856 51854 57858 sw
rect 47767 57854 51854 57856
tri 51854 57854 51856 57856 sw
rect 47767 57852 51856 57854
tri 51856 57852 51858 57854 sw
rect 47767 57850 51858 57852
tri 51858 57850 51860 57852 sw
rect 47767 57848 51860 57850
tri 51860 57848 51862 57850 sw
rect 47767 57846 51862 57848
tri 51862 57846 51864 57848 sw
rect 47767 57844 51864 57846
tri 51864 57844 51866 57846 sw
rect 47767 57842 51866 57844
tri 51866 57842 51868 57844 sw
rect 47767 57840 51868 57842
tri 51868 57840 51870 57842 sw
rect 47767 57838 51870 57840
tri 51870 57838 51872 57840 sw
rect 47767 57836 51872 57838
tri 51872 57836 51874 57838 sw
rect 47767 57834 51874 57836
tri 51874 57834 51876 57836 sw
rect 47767 57832 51876 57834
tri 51876 57832 51878 57834 sw
rect 47767 57830 51878 57832
tri 51878 57830 51880 57832 sw
rect 47767 57828 51880 57830
tri 51880 57828 51882 57830 sw
rect 47767 57826 51882 57828
tri 51882 57826 51884 57828 sw
rect 47767 57824 51884 57826
tri 51884 57824 51886 57826 sw
rect 47767 57822 51886 57824
tri 51886 57822 51888 57824 sw
rect 47767 57820 51888 57822
tri 51888 57820 51890 57822 sw
rect 47767 57818 51890 57820
tri 51890 57818 51892 57820 sw
rect 47767 57816 51892 57818
tri 51892 57816 51894 57818 sw
rect 47767 57814 51894 57816
tri 51894 57814 51896 57816 sw
rect 47767 57812 51896 57814
tri 51896 57812 51898 57814 sw
rect 47767 57810 51898 57812
tri 51898 57810 51900 57812 sw
rect 47767 57808 51900 57810
tri 51900 57808 51902 57810 sw
rect 47767 57806 51902 57808
tri 51902 57806 51904 57808 sw
rect 47767 57804 51904 57806
tri 51904 57804 51906 57806 sw
rect 47767 57802 51906 57804
tri 51906 57802 51908 57804 sw
rect 47767 57800 51908 57802
tri 51908 57800 51910 57802 sw
rect 47767 57798 51910 57800
tri 51910 57798 51912 57800 sw
rect 47767 57796 51912 57798
tri 51912 57796 51914 57798 sw
rect 47767 57794 51914 57796
tri 51914 57794 51916 57796 sw
rect 47767 57792 51916 57794
tri 51916 57792 51918 57794 sw
rect 47767 57790 51918 57792
tri 51918 57790 51920 57792 sw
rect 47767 57788 51920 57790
tri 51920 57788 51922 57790 sw
rect 47767 57786 51922 57788
tri 51922 57786 51924 57788 sw
rect 47767 57784 51924 57786
tri 51924 57784 51926 57786 sw
rect 47767 57782 51926 57784
tri 51926 57782 51928 57784 sw
rect 47767 57780 51928 57782
tri 51928 57780 51930 57782 sw
rect 47767 57778 51930 57780
tri 51930 57778 51932 57780 sw
rect 47767 57776 51932 57778
tri 51932 57776 51934 57778 sw
rect 47767 57774 51934 57776
tri 51934 57774 51936 57776 sw
rect 47767 57772 51936 57774
tri 51936 57772 51938 57774 sw
tri 51985 57772 52223 58010 ne
rect 52223 57856 53835 58010
tri 53835 57856 54119 58140 sw
tri 54119 57856 54403 58140 ne
rect 54403 58010 56099 58140
tri 56099 58010 56229 58140 sw
tri 56387 58010 56517 58140 ne
rect 56517 58010 58367 58140
tri 58367 58010 58497 58140 sw
tri 58653 58010 58783 58140 ne
rect 58783 58010 60633 58140
tri 60633 58010 60763 58140 sw
tri 60916 58010 61046 58140 ne
rect 61046 58010 62896 58140
tri 62896 58010 63026 58140 sw
tri 63179 58010 63309 58140 ne
rect 63309 58010 71000 58140
rect 54403 57856 56229 58010
rect 52223 57772 54119 57856
rect 47767 57694 51938 57772
rect 43272 57625 47456 57694
rect 41200 57430 42985 57625
tri 41200 57338 41292 57430 ne
rect 41292 57338 42985 57430
tri 42985 57338 43272 57625 sw
tri 43272 57338 43559 57625 ne
rect 43559 57388 47456 57625
tri 47456 57388 47762 57694 sw
tri 47767 57659 47802 57694 ne
rect 47802 57659 51938 57694
rect 43559 57348 47762 57388
tri 47762 57348 47802 57388 sw
tri 47802 57348 48113 57659 ne
rect 48113 57487 51938 57659
tri 51938 57487 52223 57772 sw
tri 52223 57487 52508 57772 ne
rect 52508 57770 54119 57772
tri 54119 57770 54205 57856 sw
tri 54403 57770 54489 57856 ne
rect 54489 57770 56229 57856
rect 52508 57487 54205 57770
rect 48113 57348 52223 57487
rect 43559 57338 47802 57348
tri 41000 57138 41200 57338 sw
tri 41292 57138 41492 57338 ne
rect 41492 57207 43272 57338
tri 43272 57207 43403 57338 sw
tri 43559 57207 43690 57338 ne
rect 43690 57207 47802 57338
rect 41492 57138 43403 57207
rect 39600 56920 41200 57138
tri 41200 56920 41418 57138 sw
tri 41492 56920 41710 57138 ne
rect 41710 56920 43403 57138
tri 43403 56920 43690 57207 sw
tri 43690 56920 43977 57207 ne
rect 43977 57040 47802 57207
tri 47802 57040 48110 57348 sw
tri 48113 57241 48220 57348 ne
rect 48220 57241 52223 57348
rect 43977 56930 48110 57040
tri 48110 56930 48220 57040 sw
tri 48220 56930 48531 57241 ne
rect 48531 57202 52223 57241
tri 52223 57202 52508 57487 sw
tri 52508 57207 52788 57487 ne
rect 52788 57486 54205 57487
tri 54205 57486 54489 57770 sw
tri 54489 57486 54773 57770 ne
rect 54773 57760 56229 57770
tri 56229 57760 56479 58010 sw
tri 56517 57760 56767 58010 ne
rect 56767 57760 58497 58010
tri 58497 57760 58747 58010 sw
tri 58783 57760 59033 58010 ne
rect 59033 57760 60763 58010
tri 60763 57760 61013 58010 sw
tri 61046 57760 61296 58010 ne
rect 61296 57760 63026 58010
tri 63026 57760 63276 58010 sw
tri 63309 57760 63559 58010 ne
rect 63559 57760 71000 58010
rect 54773 57486 56479 57760
tri 56479 57486 56753 57760 sw
tri 56767 57486 57041 57760 ne
rect 57041 57486 58747 57760
tri 58747 57486 59021 57760 sw
tri 59033 57486 59307 57760 ne
rect 59307 57486 61013 57760
tri 61013 57486 61287 57760 sw
tri 61296 57486 61570 57760 ne
rect 61570 57486 63276 57760
tri 63276 57486 63550 57760 sw
tri 63559 57486 63833 57760 ne
rect 63833 57486 71000 57760
rect 52788 57207 54489 57486
rect 48531 57201 52508 57202
tri 52508 57201 52509 57202 sw
rect 48531 57200 52509 57201
tri 52509 57200 52510 57201 sw
rect 48531 57199 52510 57200
tri 52510 57199 52511 57200 sw
rect 48531 57198 52511 57199
tri 52511 57198 52512 57199 sw
rect 48531 57197 52512 57198
tri 52512 57197 52513 57198 sw
rect 48531 57196 52513 57197
tri 52513 57196 52514 57197 sw
rect 48531 57195 52514 57196
tri 52514 57195 52515 57196 sw
rect 48531 57194 52515 57195
tri 52515 57194 52516 57195 sw
rect 48531 57193 52516 57194
tri 52516 57193 52517 57194 sw
rect 48531 57192 52517 57193
tri 52517 57192 52518 57193 sw
rect 48531 57191 52518 57192
tri 52518 57191 52519 57192 sw
rect 48531 57190 52519 57191
tri 52519 57190 52520 57191 sw
rect 48531 57189 52520 57190
tri 52520 57189 52521 57190 sw
rect 48531 57188 52521 57189
tri 52521 57188 52522 57189 sw
rect 48531 57187 52522 57188
tri 52522 57187 52523 57188 sw
rect 48531 57186 52523 57187
tri 52523 57186 52524 57187 sw
rect 48531 57185 52524 57186
tri 52524 57185 52525 57186 sw
rect 48531 57184 52525 57185
tri 52525 57184 52526 57185 sw
rect 48531 57183 52526 57184
tri 52526 57183 52527 57184 sw
rect 48531 57182 52527 57183
tri 52527 57182 52528 57183 sw
rect 48531 57181 52528 57182
tri 52528 57181 52529 57182 sw
rect 48531 57180 52529 57181
tri 52529 57180 52530 57181 sw
rect 48531 57179 52530 57180
tri 52530 57179 52531 57180 sw
rect 48531 57178 52531 57179
tri 52531 57178 52532 57179 sw
rect 48531 57177 52532 57178
tri 52532 57177 52533 57178 sw
rect 48531 57176 52533 57177
tri 52533 57176 52534 57177 sw
rect 48531 57175 52534 57176
tri 52534 57175 52535 57176 sw
rect 48531 57174 52535 57175
tri 52535 57174 52536 57175 sw
rect 48531 57173 52536 57174
tri 52536 57173 52537 57174 sw
rect 48531 57172 52537 57173
tri 52537 57172 52538 57173 sw
rect 48531 57171 52538 57172
tri 52538 57171 52539 57172 sw
rect 48531 57170 52539 57171
tri 52539 57170 52540 57171 sw
rect 48531 57169 52540 57170
tri 52540 57169 52541 57170 sw
rect 48531 57168 52541 57169
tri 52541 57168 52542 57169 sw
rect 48531 57167 52542 57168
tri 52542 57167 52543 57168 sw
rect 48531 57166 52543 57167
tri 52543 57166 52544 57167 sw
rect 48531 57165 52544 57166
tri 52544 57165 52545 57166 sw
rect 48531 57164 52545 57165
tri 52545 57164 52546 57165 sw
rect 48531 57163 52546 57164
tri 52546 57163 52547 57164 sw
rect 48531 57162 52547 57163
tri 52547 57162 52548 57163 sw
rect 48531 57161 52548 57162
tri 52548 57161 52549 57162 sw
rect 48531 57160 52549 57161
tri 52549 57160 52550 57161 sw
rect 48531 57159 52550 57160
tri 52550 57159 52551 57160 sw
rect 48531 57158 52551 57159
tri 52551 57158 52552 57159 sw
rect 48531 57157 52552 57158
tri 52552 57157 52553 57158 sw
rect 48531 57156 52553 57157
tri 52553 57156 52554 57157 sw
rect 48531 57155 52554 57156
tri 52554 57155 52555 57156 sw
rect 48531 57154 52555 57155
tri 52555 57154 52556 57155 sw
rect 48531 57153 52556 57154
tri 52556 57153 52557 57154 sw
rect 48531 57152 52557 57153
tri 52557 57152 52558 57153 sw
rect 48531 57151 52558 57152
tri 52558 57151 52559 57152 sw
rect 48531 57150 52559 57151
tri 52559 57150 52560 57151 sw
rect 48531 57149 52560 57150
tri 52560 57149 52561 57150 sw
rect 48531 57148 52561 57149
tri 52561 57148 52562 57149 sw
rect 48531 57147 52562 57148
tri 52562 57147 52563 57148 sw
rect 48531 57146 52563 57147
tri 52563 57146 52564 57147 sw
rect 48531 57145 52564 57146
tri 52564 57145 52565 57146 sw
rect 48531 57144 52565 57145
tri 52565 57144 52566 57145 sw
rect 48531 57143 52566 57144
tri 52566 57143 52567 57144 sw
rect 48531 57142 52567 57143
tri 52567 57142 52568 57143 sw
rect 48531 57141 52568 57142
tri 52568 57141 52569 57142 sw
rect 48531 57140 52569 57141
tri 52569 57140 52570 57141 sw
rect 48531 57139 52570 57140
tri 52570 57139 52571 57140 sw
rect 48531 57138 52571 57139
tri 52571 57138 52572 57139 sw
rect 48531 57137 52572 57138
tri 52572 57137 52573 57138 sw
rect 48531 57136 52573 57137
tri 52573 57136 52574 57137 sw
rect 48531 57135 52574 57136
tri 52574 57135 52575 57136 sw
rect 48531 57134 52575 57135
tri 52575 57134 52576 57135 sw
rect 48531 57133 52576 57134
tri 52576 57133 52577 57134 sw
rect 48531 57132 52577 57133
tri 52577 57132 52578 57133 sw
rect 48531 57131 52578 57132
tri 52578 57131 52579 57132 sw
rect 48531 57130 52579 57131
tri 52579 57130 52580 57131 sw
rect 48531 57129 52580 57130
tri 52580 57129 52581 57130 sw
rect 48531 57128 52581 57129
tri 52581 57128 52582 57129 sw
rect 48531 57127 52582 57128
tri 52582 57127 52583 57128 sw
rect 48531 57126 52583 57127
tri 52583 57126 52584 57127 sw
rect 48531 57125 52584 57126
tri 52584 57125 52585 57126 sw
rect 48531 57124 52585 57125
tri 52585 57124 52586 57125 sw
rect 48531 57123 52586 57124
tri 52586 57123 52587 57124 sw
rect 48531 57122 52587 57123
tri 52587 57122 52588 57123 sw
rect 48531 57121 52588 57122
tri 52588 57121 52589 57122 sw
rect 48531 57120 52589 57121
tri 52589 57120 52590 57121 sw
rect 48531 57119 52590 57120
tri 52590 57119 52591 57120 sw
rect 48531 57118 52591 57119
tri 52591 57118 52592 57119 sw
rect 48531 57117 52592 57118
tri 52592 57117 52593 57118 sw
rect 48531 57116 52593 57117
tri 52593 57116 52594 57117 sw
rect 48531 57115 52594 57116
tri 52594 57115 52595 57116 sw
rect 48531 57114 52595 57115
tri 52595 57114 52596 57115 sw
rect 48531 57113 52596 57114
tri 52596 57113 52597 57114 sw
rect 48531 57112 52597 57113
tri 52597 57112 52598 57113 sw
rect 48531 57110 52598 57112
tri 52598 57110 52600 57112 sw
rect 48531 57108 52600 57110
tri 52600 57108 52602 57110 sw
rect 48531 57106 52602 57108
tri 52602 57106 52604 57108 sw
rect 48531 57104 52604 57106
tri 52604 57104 52606 57106 sw
rect 48531 57102 52606 57104
tri 52606 57102 52608 57104 sw
rect 48531 57100 52608 57102
tri 52608 57100 52610 57102 sw
rect 48531 57098 52610 57100
tri 52610 57098 52612 57100 sw
rect 48531 57096 52612 57098
tri 52612 57096 52614 57098 sw
rect 48531 57094 52614 57096
tri 52614 57094 52616 57096 sw
rect 48531 57092 52616 57094
tri 52616 57092 52618 57094 sw
rect 48531 57090 52618 57092
tri 52618 57090 52620 57092 sw
rect 48531 57088 52620 57090
tri 52620 57088 52622 57090 sw
rect 48531 57086 52622 57088
tri 52622 57086 52624 57088 sw
rect 48531 57084 52624 57086
tri 52624 57084 52626 57086 sw
rect 48531 57082 52626 57084
tri 52626 57082 52628 57084 sw
rect 48531 57080 52628 57082
tri 52628 57080 52630 57082 sw
rect 48531 57078 52630 57080
tri 52630 57078 52632 57080 sw
rect 48531 57076 52632 57078
tri 52632 57076 52634 57078 sw
rect 48531 57074 52634 57076
tri 52634 57074 52636 57076 sw
rect 48531 57072 52636 57074
tri 52636 57072 52638 57074 sw
rect 48531 57070 52638 57072
tri 52638 57070 52640 57072 sw
rect 48531 57068 52640 57070
tri 52640 57068 52642 57070 sw
rect 48531 57066 52642 57068
tri 52642 57066 52644 57068 sw
rect 48531 57064 52644 57066
tri 52644 57064 52646 57066 sw
rect 48531 57062 52646 57064
tri 52646 57062 52648 57064 sw
rect 48531 57060 52648 57062
tri 52648 57060 52650 57062 sw
rect 48531 57058 52650 57060
tri 52650 57058 52652 57060 sw
rect 48531 57056 52652 57058
tri 52652 57056 52654 57058 sw
rect 48531 57054 52654 57056
tri 52654 57054 52656 57056 sw
rect 48531 57052 52656 57054
tri 52656 57052 52658 57054 sw
rect 48531 57050 52658 57052
tri 52658 57050 52660 57052 sw
rect 48531 57048 52660 57050
tri 52660 57048 52662 57050 sw
rect 48531 57046 52662 57048
tri 52662 57046 52664 57048 sw
rect 48531 57044 52664 57046
tri 52664 57044 52666 57046 sw
rect 48531 57042 52666 57044
tri 52666 57042 52668 57044 sw
rect 48531 57040 52668 57042
tri 52668 57040 52670 57042 sw
rect 48531 57038 52670 57040
tri 52670 57038 52672 57040 sw
rect 48531 57036 52672 57038
tri 52672 57036 52674 57038 sw
rect 48531 57034 52674 57036
tri 52674 57034 52676 57036 sw
rect 48531 57032 52676 57034
tri 52676 57032 52678 57034 sw
rect 48531 57030 52678 57032
tri 52678 57030 52680 57032 sw
rect 48531 57028 52680 57030
tri 52680 57028 52682 57030 sw
rect 48531 57026 52682 57028
tri 52682 57026 52684 57028 sw
rect 48531 57024 52684 57026
tri 52684 57024 52686 57026 sw
rect 48531 57022 52686 57024
tri 52686 57022 52688 57024 sw
rect 48531 57020 52688 57022
tri 52688 57020 52690 57022 sw
rect 48531 57018 52690 57020
tri 52690 57018 52692 57020 sw
rect 48531 57016 52692 57018
tri 52692 57016 52694 57018 sw
rect 48531 57014 52694 57016
tri 52694 57014 52696 57016 sw
rect 48531 57012 52696 57014
tri 52696 57012 52698 57014 sw
rect 48531 57010 52698 57012
tri 52698 57010 52700 57012 sw
rect 48531 57008 52700 57010
tri 52700 57008 52702 57010 sw
rect 48531 57006 52702 57008
tri 52702 57006 52704 57008 sw
rect 48531 57004 52704 57006
tri 52704 57004 52706 57006 sw
rect 48531 57002 52706 57004
tri 52706 57002 52708 57004 sw
rect 48531 57000 52708 57002
tri 52708 57000 52710 57002 sw
rect 48531 56998 52710 57000
tri 52710 56998 52712 57000 sw
rect 48531 56996 52712 56998
tri 52712 56996 52714 56998 sw
rect 48531 56994 52714 56996
tri 52714 56994 52716 56996 sw
rect 48531 56992 52716 56994
tri 52716 56992 52718 56994 sw
rect 48531 56990 52718 56992
tri 52718 56990 52720 56992 sw
rect 48531 56988 52720 56990
tri 52720 56988 52722 56990 sw
rect 48531 56986 52722 56988
tri 52722 56986 52724 56988 sw
rect 48531 56984 52724 56986
tri 52724 56984 52726 56986 sw
rect 48531 56982 52726 56984
tri 52726 56982 52728 56984 sw
rect 48531 56980 52728 56982
tri 52728 56980 52730 56982 sw
rect 48531 56978 52730 56980
tri 52730 56978 52732 56980 sw
rect 48531 56976 52732 56978
tri 52732 56976 52734 56978 sw
rect 48531 56974 52734 56976
tri 52734 56974 52736 56976 sw
rect 48531 56972 52736 56974
tri 52736 56972 52738 56974 sw
rect 48531 56970 52738 56972
tri 52738 56970 52740 56972 sw
rect 48531 56968 52740 56970
tri 52740 56968 52742 56970 sw
rect 48531 56966 52742 56968
tri 52742 56966 52744 56968 sw
rect 48531 56964 52744 56966
tri 52744 56964 52746 56966 sw
rect 48531 56962 52746 56964
tri 52746 56962 52748 56964 sw
rect 48531 56960 52748 56962
tri 52748 56960 52750 56962 sw
rect 48531 56958 52750 56960
tri 52750 56958 52752 56960 sw
rect 48531 56956 52752 56958
tri 52752 56956 52754 56958 sw
rect 48531 56954 52754 56956
tri 52754 56954 52756 56956 sw
rect 48531 56952 52756 56954
tri 52756 56952 52758 56954 sw
rect 48531 56950 52758 56952
tri 52758 56950 52760 56952 sw
rect 48531 56948 52760 56950
tri 52760 56948 52762 56950 sw
rect 48531 56946 52762 56948
tri 52762 56946 52764 56948 sw
rect 48531 56944 52764 56946
tri 52764 56944 52766 56946 sw
rect 48531 56942 52766 56944
tri 52766 56942 52768 56944 sw
rect 48531 56940 52768 56942
tri 52768 56940 52770 56942 sw
rect 48531 56938 52770 56940
tri 52770 56938 52772 56940 sw
rect 48531 56936 52772 56938
tri 52772 56936 52774 56938 sw
rect 48531 56934 52774 56936
tri 52774 56934 52776 56936 sw
rect 48531 56932 52776 56934
tri 52776 56932 52778 56934 sw
rect 48531 56930 52778 56932
tri 52778 56930 52780 56932 sw
rect 43977 56920 48220 56930
rect 39600 56840 41418 56920
tri 41418 56840 41498 56920 sw
tri 41710 56840 41790 56920 ne
rect 41790 56840 43690 56920
rect 39600 56758 41498 56840
tri 39400 56664 39401 56665 sw
tri 39600 56664 39694 56758 ne
rect 39694 56664 41498 56758
tri 41498 56664 41674 56840 sw
tri 41790 56664 41966 56840 ne
rect 41966 56664 43690 56840
tri 43690 56664 43946 56920 sw
tri 43977 56664 44233 56920 ne
rect 44233 56664 48220 56920
rect 36400 56371 39401 56664
tri 39401 56371 39694 56664 sw
tri 39694 56371 39987 56664 ne
rect 39987 56663 41674 56664
tri 41674 56663 41675 56664 sw
tri 41966 56663 41967 56664 ne
rect 41967 56663 43946 56664
rect 39987 56371 41675 56663
tri 41675 56371 41967 56663 sw
tri 41967 56460 42170 56663 ne
rect 42170 56460 43946 56663
tri 43946 56460 44150 56664 sw
tri 44233 56460 44437 56664 ne
rect 44437 56624 48220 56664
tri 48220 56624 48526 56930 sw
tri 48531 56664 48797 56930 ne
rect 48797 56928 52780 56930
tri 52780 56928 52782 56930 sw
rect 48797 56926 52782 56928
tri 52782 56926 52784 56928 sw
rect 48797 56924 52784 56926
tri 52784 56924 52786 56926 sw
rect 48797 56922 52786 56924
tri 52786 56922 52788 56924 sw
tri 52788 56922 53073 57207 ne
rect 53073 57204 54489 57207
tri 54489 57204 54771 57486 sw
tri 54773 57204 55055 57486 ne
rect 55055 57472 56753 57486
tri 56753 57472 56767 57486 sw
tri 57041 57472 57055 57486 ne
rect 57055 57472 59021 57486
rect 55055 57338 56767 57472
tri 56767 57338 56901 57472 sw
tri 57055 57338 57189 57472 ne
rect 57189 57380 59021 57472
tri 59021 57380 59127 57486 sw
tri 59307 57380 59413 57486 ne
rect 59413 57380 61287 57486
tri 61287 57380 61393 57486 sw
tri 61570 57380 61676 57486 ne
rect 61676 57380 63550 57486
tri 63550 57380 63656 57486 sw
tri 63833 57380 63939 57486 ne
rect 63939 57380 71000 57486
rect 57189 57338 59127 57380
tri 59127 57338 59169 57380 sw
tri 59413 57338 59455 57380 ne
rect 59455 57338 61393 57380
tri 61393 57338 61435 57380 sw
tri 61676 57338 61718 57380 ne
rect 61718 57338 63656 57380
tri 63656 57338 63698 57380 sw
tri 63939 57338 63981 57380 ne
rect 63981 57338 71000 57380
rect 55055 57208 56901 57338
tri 56901 57208 57031 57338 sw
tri 57189 57208 57319 57338 ne
rect 57319 57208 59169 57338
rect 55055 57204 57031 57208
rect 53073 56922 54771 57204
rect 48797 56664 52788 56922
rect 44437 56460 48526 56624
tri 42170 56371 42259 56460 ne
rect 42259 56371 44150 56460
tri 44150 56371 44239 56460 sw
tri 44437 56371 44526 56460 ne
rect 44526 56371 48526 56460
rect 36400 56078 39694 56371
tri 39694 56078 39987 56371 sw
tri 39987 56078 40280 56371 ne
rect 40280 56322 41967 56371
tri 41967 56322 42016 56371 sw
tri 42259 56322 42308 56371 ne
rect 42308 56322 44239 56371
rect 40280 56078 42016 56322
rect 36400 55785 39987 56078
tri 39987 55785 40280 56078 sw
tri 40280 55994 40364 56078 ne
rect 40364 56030 42016 56078
tri 42016 56030 42308 56322 sw
tri 42308 56030 42600 56322 ne
rect 42600 56084 44239 56322
tri 44239 56084 44526 56371 sw
tri 44526 56084 44813 56371 ne
rect 44813 56361 48526 56371
tri 48526 56361 48789 56624 sw
tri 48797 56371 49090 56664 ne
rect 49090 56638 52788 56664
tri 52788 56638 53072 56922 sw
tri 53073 56664 53331 56922 ne
rect 53331 56920 54771 56922
tri 54771 56920 55055 57204 sw
tri 55055 56920 55339 57204 ne
rect 55339 56920 57031 57204
tri 57031 56920 57319 57208 sw
tri 57319 56920 57607 57208 ne
rect 57607 57094 59169 57208
tri 59169 57094 59413 57338 sw
tri 59455 57094 59699 57338 ne
rect 59699 57283 61435 57338
tri 61435 57283 61490 57338 sw
tri 61718 57283 61773 57338 ne
rect 61773 57283 63698 57338
rect 59699 57094 61490 57283
rect 57607 56920 59413 57094
tri 59413 56920 59587 57094 sw
tri 59699 56920 59873 57094 ne
rect 59873 57000 61490 57094
tri 61490 57000 61773 57283 sw
tri 61773 57000 62056 57283 ne
rect 62056 57200 63698 57283
tri 63698 57200 63836 57338 sw
tri 63981 57200 64119 57338 ne
rect 64119 57200 71000 57338
rect 62056 57000 63836 57200
tri 63836 57000 64036 57200 sw
rect 59873 56920 61773 57000
tri 61773 56920 61853 57000 sw
tri 62056 56920 62136 57000 ne
rect 62136 56920 71000 57000
rect 53331 56664 55055 56920
tri 55055 56664 55311 56920 sw
tri 55339 56840 55419 56920 ne
rect 55419 56840 57319 56920
tri 57319 56840 57399 56920 sw
tri 57607 56840 57687 56920 ne
rect 57687 56840 59587 56920
tri 59587 56840 59667 56920 sw
tri 59873 56840 59953 56920 ne
rect 59953 56840 61853 56920
tri 61853 56840 61933 56920 sw
tri 62136 56840 62216 56920 ne
rect 62216 56910 71000 56920
rect 62216 56840 70613 56910
tri 55419 56664 55595 56840 ne
rect 55595 56664 57399 56840
tri 57399 56664 57575 56840 sw
tri 57687 56664 57863 56840 ne
rect 57863 56664 59667 56840
tri 59667 56664 59843 56840 sw
tri 59953 56664 60129 56840 ne
rect 60129 56717 61933 56840
tri 61933 56717 62056 56840 sw
tri 62216 56717 62339 56840 ne
rect 62339 56717 70613 56840
rect 60129 56664 62056 56717
tri 62056 56664 62109 56717 sw
tri 62339 56664 62392 56717 ne
rect 62392 56664 70613 56717
rect 49090 56379 53072 56638
tri 53072 56379 53331 56638 sw
tri 53331 56460 53535 56664 ne
rect 53535 56540 55311 56664
tri 55311 56540 55435 56664 sw
tri 55595 56540 55719 56664 ne
rect 55719 56540 57575 56664
tri 57575 56540 57699 56664 sw
tri 57863 56540 57987 56664 ne
rect 57987 56540 59843 56664
tri 59843 56540 59967 56664 sw
tri 60129 56540 60253 56664 ne
rect 60253 56540 62109 56664
tri 62109 56540 62233 56664 sw
tri 62392 56540 62516 56664 ne
rect 62516 56540 70613 56664
rect 53535 56460 55435 56540
tri 55435 56460 55515 56540 sw
tri 55719 56460 55799 56540 ne
rect 55799 56460 57699 56540
tri 57699 56460 57779 56540 sw
tri 57987 56460 58067 56540 ne
rect 58067 56460 59967 56540
tri 59967 56460 60047 56540 sw
tri 60253 56460 60333 56540 ne
rect 60333 56460 62233 56540
tri 62233 56460 62313 56540 sw
tri 62516 56460 62596 56540 ne
rect 62596 56460 70613 56540
rect 49090 56371 53331 56379
rect 44813 56084 48789 56361
rect 42600 56030 44526 56084
rect 40364 55994 42308 56030
rect 36400 55701 40280 55785
tri 40280 55701 40364 55785 sw
tri 40364 55714 40644 55994 ne
rect 40644 55738 42308 55994
tri 42308 55738 42600 56030 sw
tri 42600 55738 42892 56030 ne
rect 42892 55987 44526 56030
tri 44526 55987 44623 56084 sw
tri 44813 55987 44910 56084 ne
rect 44910 56061 48789 56084
tri 48789 56061 49089 56361 sw
tri 49090 56140 49321 56371 ne
rect 49321 56175 53331 56371
tri 53331 56175 53535 56379 sw
tri 53535 56253 53742 56460 ne
rect 53742 56371 55515 56460
tri 55515 56371 55604 56460 sw
tri 55799 56371 55888 56460 ne
rect 55888 56371 57779 56460
tri 57779 56371 57868 56460 sw
tri 58067 56371 58156 56460 ne
rect 58156 56371 60047 56460
tri 60047 56371 60136 56460 sw
tri 60333 56371 60422 56460 ne
rect 60422 56371 62313 56460
tri 62313 56371 62402 56460 sw
tri 62596 56371 62685 56460 ne
rect 62685 56371 70613 56460
rect 53742 56253 55604 56371
rect 49321 56140 53535 56175
rect 44910 55987 49089 56061
rect 42892 55738 44623 55987
rect 40644 55714 42600 55738
rect 36400 55421 40364 55701
tri 40364 55421 40644 55701 sw
tri 40644 55617 40741 55714 ne
rect 40741 55700 42600 55714
tri 42600 55700 42638 55738 sw
rect 40741 55617 42638 55700
tri 40741 55421 40937 55617 ne
rect 40937 55615 42638 55617
tri 42638 55615 42723 55700 sw
rect 40937 55538 42723 55615
tri 42723 55538 42800 55615 sw
tri 42892 55538 43092 55738 ne
rect 43092 55700 44623 55738
tri 44623 55700 44910 55987 sw
tri 44910 55700 45197 55987 ne
rect 45197 55830 49089 55987
tri 49089 55830 49320 56061 sw
tri 49321 55870 49591 56140 ne
rect 49591 55968 53535 56140
tri 53535 55968 53742 56175 sw
tri 53742 55987 54008 56253 ne
rect 54008 56160 55604 56253
tri 55604 56160 55815 56371 sw
tri 55888 56160 56099 56371 ne
rect 56099 56160 57868 56371
tri 57868 56160 58079 56371 sw
tri 58156 56160 58367 56371 ne
rect 58367 56160 60136 56371
tri 60136 56160 60347 56371 sw
tri 60422 56160 60633 56371 ne
rect 60633 56160 62402 56371
tri 62402 56160 62613 56371 sw
tri 62685 56160 62896 56371 ne
rect 62896 56160 70613 56371
rect 54008 55987 55815 56160
rect 49591 55870 53742 55968
rect 45197 55700 49320 55830
rect 43092 55559 44910 55700
tri 44910 55559 45051 55700 sw
tri 45197 55559 45338 55700 ne
rect 45338 55559 49320 55700
tri 49320 55559 49591 55830 sw
tri 49591 55644 49817 55870 ne
rect 49817 55702 53742 55870
tri 53742 55702 54008 55968 sw
tri 54008 55702 54293 55987 ne
rect 54293 55876 55815 55987
tri 55815 55876 56099 56160 sw
tri 56099 55876 56383 56160 ne
rect 56383 56068 58079 56160
tri 58079 56068 58171 56160 sw
tri 58367 56068 58459 56160 ne
rect 58459 56068 60347 56160
rect 56383 55876 58171 56068
rect 54293 55702 56099 55876
rect 49817 55644 54008 55702
tri 49817 55559 49902 55644 ne
rect 49902 55559 54008 55644
rect 43092 55538 45051 55559
rect 40937 55421 42800 55538
tri 36400 55324 36497 55421 ne
rect 36497 55324 40644 55421
tri 36200 55027 36497 55324 sw
tri 36497 55123 36698 55324 ne
rect 36698 55128 40644 55324
tri 40644 55128 40937 55421 sw
tri 40937 55154 41204 55421 ne
rect 41204 55323 42800 55421
tri 42800 55323 43015 55538 sw
tri 43092 55323 43307 55538 ne
rect 43307 55323 45051 55538
rect 41204 55312 43015 55323
tri 43015 55312 43026 55323 sw
tri 43307 55312 43318 55323 ne
rect 43318 55312 45051 55323
tri 45051 55312 45298 55559 sw
rect 41204 55154 43026 55312
rect 36698 55123 40937 55128
rect 33200 54826 36497 55027
tri 36497 54826 36698 55027 sw
tri 36698 54826 36995 55123 ne
rect 36995 54861 40937 55123
tri 40937 54861 41204 55128 sw
tri 41204 54861 41497 55154 ne
rect 41497 55152 43026 55154
tri 43026 55152 43186 55312 sw
tri 43318 55152 43478 55312 ne
rect 43478 55272 45298 55312
tri 45298 55272 45338 55312 sw
tri 45338 55272 45625 55559 ne
rect 45625 55272 49591 55559
rect 43478 55152 45338 55272
rect 41497 54861 43186 55152
rect 36995 54826 41204 54861
rect 33200 54529 36698 54826
tri 36698 54529 36995 54826 sw
tri 36995 54688 37133 54826 ne
rect 37133 54688 41204 54826
rect 33200 54391 36995 54529
tri 36995 54391 37133 54529 sw
tri 37133 54391 37430 54688 ne
rect 37430 54568 41204 54688
tri 41204 54568 41497 54861 sw
tri 41497 54860 41498 54861 ne
rect 41498 54860 43186 54861
tri 43186 54860 43478 55152 sw
tri 43478 54860 43770 55152 ne
rect 43770 55147 45338 55152
tri 45338 55147 45463 55272 sw
tri 45625 55147 45750 55272 ne
rect 45750 55251 49591 55272
tri 49591 55251 49899 55559 sw
tri 49902 55323 50138 55559 ne
rect 50138 55417 54008 55559
tri 54008 55417 54293 55702 sw
tri 54293 55610 54385 55702 ne
rect 54385 55700 56099 55702
tri 56099 55700 56275 55876 sw
tri 56383 55700 56559 55876 ne
rect 56559 55780 58171 55876
tri 58171 55780 58459 56068 sw
tri 58459 55780 58747 56068 ne
rect 58747 56066 60347 56068
tri 60347 56066 60441 56160 sw
tri 60633 56066 60727 56160 ne
rect 60727 56066 62613 56160
rect 58747 55780 60441 56066
tri 60441 55780 60727 56066 sw
tri 60727 55780 61013 56066 ne
rect 61013 56063 62613 56066
tri 62613 56063 62710 56160 sw
tri 62896 56063 62993 56160 ne
rect 62993 56063 70613 56160
rect 61013 55780 62710 56063
tri 62710 55780 62993 56063 sw
tri 62993 55780 63276 56063 ne
rect 63276 55780 70613 56063
rect 56559 55700 58459 55780
tri 58459 55700 58539 55780 sw
tri 58747 55700 58827 55780 ne
rect 58827 55700 60727 55780
tri 60727 55700 60807 55780 sw
tri 61013 55700 61093 55780 ne
rect 61093 55700 62993 55780
tri 62993 55700 63073 55780 sw
tri 63276 55700 63356 55780 ne
rect 63356 55710 70613 55780
rect 70669 55710 71000 56910
rect 63356 55700 71000 55710
rect 54385 55610 56275 55700
rect 50138 55325 54293 55417
tri 54293 55325 54385 55417 sw
tri 54385 55325 54670 55610 ne
rect 54670 55607 56275 55610
tri 56275 55607 56368 55700 sw
tri 56559 55607 56652 55700 ne
rect 56652 55607 58539 55700
rect 54670 55325 56368 55607
rect 50138 55323 54385 55325
rect 45750 55147 49899 55251
rect 43770 54860 45463 55147
tri 45463 54860 45750 55147 sw
tri 45750 54860 46037 55147 ne
rect 46037 55020 49899 55147
tri 49899 55020 50130 55251 sw
tri 50138 55181 50280 55323 ne
rect 50280 55181 54385 55323
rect 46037 54870 50130 55020
tri 50130 54870 50280 55020 sw
tri 50280 54870 50591 55181 ne
rect 50591 55040 54385 55181
tri 54385 55040 54670 55325 sw
tri 54670 55147 54848 55325 ne
rect 54848 55323 56368 55325
tri 56368 55323 56652 55607 sw
tri 56652 55323 56936 55607 ne
rect 56936 55492 58539 55607
tri 58539 55492 58747 55700 sw
tri 58827 55492 59035 55700 ne
rect 59035 55686 60807 55700
tri 60807 55686 60821 55700 sw
tri 61093 55686 61107 55700 ne
rect 61107 55686 63073 55700
rect 59035 55492 60821 55686
rect 56936 55323 58747 55492
tri 58747 55323 58916 55492 sw
tri 59035 55323 59204 55492 ne
rect 59204 55400 60821 55492
tri 60821 55400 61107 55686 sw
tri 61107 55400 61393 55686 ne
rect 61393 55600 63073 55686
tri 63073 55600 63173 55700 sw
tri 63356 55600 63456 55700 ne
rect 63456 55600 71000 55700
rect 61393 55400 63173 55600
tri 63173 55400 63373 55600 sw
rect 59204 55323 61107 55400
tri 61107 55323 61184 55400 sw
tri 61393 55323 61470 55400 ne
rect 61470 55323 71000 55400
rect 54848 55312 56652 55323
tri 56652 55312 56663 55323 sw
tri 56936 55312 56947 55323 ne
rect 56947 55312 58916 55323
tri 58916 55312 58927 55323 sw
tri 59204 55312 59215 55323 ne
rect 59215 55312 61184 55323
tri 61184 55312 61195 55323 sw
tri 61470 55312 61481 55323 ne
rect 61481 55312 71000 55323
rect 54848 55147 56663 55312
rect 50591 54870 54670 55040
rect 46037 54860 50280 54870
rect 37430 54567 41497 54568
tri 41497 54567 41498 54568 sw
tri 41498 54567 41791 54860 ne
rect 41791 54772 43478 54860
tri 43478 54772 43566 54860 sw
tri 43770 54772 43858 54860 ne
rect 43858 54772 45750 54860
rect 41791 54567 43566 54772
rect 37430 54391 41498 54567
rect 33200 54094 37133 54391
tri 37133 54094 37430 54391 sw
tri 37430 54377 37444 54391 ne
rect 37444 54377 41498 54391
rect 33200 54080 37430 54094
tri 37430 54080 37444 54094 sw
tri 37444 54092 37729 54377 ne
rect 37729 54274 41498 54377
tri 41498 54274 41791 54567 sw
tri 41791 54386 41972 54567 ne
rect 41972 54480 43566 54567
tri 43566 54480 43858 54772 sw
tri 43858 54480 44150 54772 ne
rect 44150 54767 45750 54772
tri 45750 54767 45843 54860 sw
tri 46037 54767 46130 54860 ne
rect 46130 54767 50280 54860
rect 44150 54480 45843 54767
tri 45843 54480 46130 54767 sw
tri 46130 54480 46417 54767 ne
rect 46417 54568 50280 54767
tri 50280 54568 50582 54870 sw
tri 50591 54805 50656 54870 ne
rect 50656 54862 54670 54870
tri 54670 54862 54848 55040 sw
tri 54848 54862 55133 55147 ne
rect 55133 55144 56663 55147
tri 56663 55144 56831 55312 sw
tri 56947 55144 57115 55312 ne
rect 57115 55148 58927 55312
tri 58927 55148 59091 55312 sw
tri 59215 55148 59379 55312 ne
rect 59379 55148 61195 55312
rect 57115 55144 59091 55148
rect 55133 54862 56831 55144
rect 50656 54805 54848 54862
rect 46417 54498 50582 54568
tri 50582 54498 50652 54568 sw
tri 50656 54498 50963 54805 ne
rect 50963 54578 54848 54805
tri 54848 54578 55132 54862 sw
tri 55133 54783 55212 54862 ne
rect 55212 54860 56831 54862
tri 56831 54860 57115 55144 sw
tri 57115 54860 57399 55144 ne
rect 57399 54860 59091 55144
tri 59091 54860 59379 55148 sw
tri 59379 54860 59667 55148 ne
rect 59667 55114 61195 55148
tri 61195 55114 61393 55312 sw
tri 61481 55114 61679 55312 ne
rect 61679 55302 71000 55312
rect 61679 55114 70613 55302
rect 59667 54860 61393 55114
tri 61393 54860 61647 55114 sw
tri 61679 54860 61933 55114 ne
rect 61933 54860 70613 55114
rect 55212 54844 57115 54860
tri 57115 54844 57131 54860 sw
tri 57399 54844 57415 54860 ne
rect 57415 54848 59379 54860
tri 59379 54848 59391 54860 sw
tri 59667 54848 59679 54860 ne
rect 59679 54848 61647 54860
rect 57415 54844 59391 54848
rect 55212 54783 57131 54844
rect 50963 54498 55132 54578
tri 55132 54498 55212 54578 sw
tri 55212 54560 55435 54783 ne
rect 55435 54560 57131 54783
tri 57131 54560 57415 54844 sw
tri 57415 54560 57699 54844 ne
rect 57699 54560 59391 54844
tri 59391 54560 59679 54848 sw
tri 59679 54560 59967 54848 ne
rect 59967 54846 61647 54848
tri 61647 54846 61661 54860 sw
tri 61933 54846 61947 54860 ne
rect 61947 54846 70613 54860
rect 59967 54560 61661 54846
tri 61661 54560 61947 54846 sw
tri 61947 54560 62233 54846 ne
rect 62233 54560 70613 54846
rect 46417 54480 50652 54498
rect 41972 54386 43858 54480
rect 37729 54093 41791 54274
tri 41791 54093 41972 54274 sw
tri 41972 54093 42265 54386 ne
rect 42265 54286 43858 54386
tri 43858 54286 44052 54480 sw
tri 44150 54286 44344 54480 ne
rect 44344 54286 46130 54480
tri 46130 54286 46324 54480 sw
tri 46417 54286 46611 54480 ne
rect 46611 54286 50652 54480
rect 42265 54188 44052 54286
tri 44052 54188 44150 54286 sw
tri 44344 54188 44442 54286 ne
rect 44442 54188 46324 54286
rect 42265 54093 44150 54188
rect 37729 54092 41972 54093
tri 33200 53992 33288 54080 ne
rect 33288 54079 37444 54080
tri 37444 54079 37445 54080 sw
rect 33288 54078 37445 54079
tri 37445 54078 37446 54079 sw
rect 33288 54077 37446 54078
tri 37446 54077 37447 54078 sw
rect 33288 54076 37447 54077
tri 37447 54076 37448 54077 sw
rect 33288 54075 37448 54076
tri 37448 54075 37449 54076 sw
rect 33288 54074 37449 54075
tri 37449 54074 37450 54075 sw
rect 33288 54073 37450 54074
tri 37450 54073 37451 54074 sw
rect 33288 54072 37451 54073
tri 37451 54072 37452 54073 sw
rect 33288 54071 37452 54072
tri 37452 54071 37453 54072 sw
rect 33288 54070 37453 54071
tri 37453 54070 37454 54071 sw
rect 33288 54069 37454 54070
tri 37454 54069 37455 54070 sw
rect 33288 54068 37455 54069
tri 37455 54068 37456 54069 sw
rect 33288 54067 37456 54068
tri 37456 54067 37457 54068 sw
rect 33288 54066 37457 54067
tri 37457 54066 37458 54067 sw
rect 33288 54065 37458 54066
tri 37458 54065 37459 54066 sw
rect 33288 54064 37459 54065
tri 37459 54064 37460 54065 sw
rect 33288 54063 37460 54064
tri 37460 54063 37461 54064 sw
rect 33288 54062 37461 54063
tri 37461 54062 37462 54063 sw
rect 33288 54061 37462 54062
tri 37462 54061 37463 54062 sw
rect 33288 54060 37463 54061
tri 37463 54060 37464 54061 sw
rect 33288 54059 37464 54060
tri 37464 54059 37465 54060 sw
rect 33288 54058 37465 54059
tri 37465 54058 37466 54059 sw
rect 33288 54057 37466 54058
tri 37466 54057 37467 54058 sw
rect 33288 54056 37467 54057
tri 37467 54056 37468 54057 sw
rect 33288 54055 37468 54056
tri 37468 54055 37469 54056 sw
rect 33288 54054 37469 54055
tri 37469 54054 37470 54055 sw
rect 33288 54053 37470 54054
tri 37470 54053 37471 54054 sw
rect 33288 54052 37471 54053
tri 37471 54052 37472 54053 sw
rect 33288 54051 37472 54052
tri 37472 54051 37473 54052 sw
rect 33288 54050 37473 54051
tri 37473 54050 37474 54051 sw
rect 33288 54049 37474 54050
tri 37474 54049 37475 54050 sw
rect 33288 54048 37475 54049
tri 37475 54048 37476 54049 sw
rect 33288 54047 37476 54048
tri 37476 54047 37477 54048 sw
rect 33288 54046 37477 54047
tri 37477 54046 37478 54047 sw
rect 33288 54045 37478 54046
tri 37478 54045 37479 54046 sw
rect 33288 54044 37479 54045
tri 37479 54044 37480 54045 sw
rect 33288 54043 37480 54044
tri 37480 54043 37481 54044 sw
rect 33288 54042 37481 54043
tri 37481 54042 37482 54043 sw
rect 33288 54041 37482 54042
tri 37482 54041 37483 54042 sw
rect 33288 54040 37483 54041
tri 37483 54040 37484 54041 sw
rect 33288 54039 37484 54040
tri 37484 54039 37485 54040 sw
rect 33288 54038 37485 54039
tri 37485 54038 37486 54039 sw
rect 33288 54037 37486 54038
tri 37486 54037 37487 54038 sw
rect 33288 54036 37487 54037
tri 37487 54036 37488 54037 sw
rect 33288 54035 37488 54036
tri 37488 54035 37489 54036 sw
rect 33288 54034 37489 54035
tri 37489 54034 37490 54035 sw
rect 33288 54033 37490 54034
tri 37490 54033 37491 54034 sw
rect 33288 54032 37491 54033
tri 37491 54032 37492 54033 sw
rect 33288 54031 37492 54032
tri 37492 54031 37493 54032 sw
rect 33288 54030 37493 54031
tri 37493 54030 37494 54031 sw
rect 33288 54029 37494 54030
tri 37494 54029 37495 54030 sw
rect 33288 54028 37495 54029
tri 37495 54028 37496 54029 sw
rect 33288 54027 37496 54028
tri 37496 54027 37497 54028 sw
rect 33288 54026 37497 54027
tri 37497 54026 37498 54027 sw
rect 33288 54025 37498 54026
tri 37498 54025 37499 54026 sw
rect 33288 54024 37499 54025
tri 37499 54024 37500 54025 sw
rect 33288 54023 37500 54024
tri 37500 54023 37501 54024 sw
rect 33288 54022 37501 54023
tri 37501 54022 37502 54023 sw
rect 33288 54021 37502 54022
tri 37502 54021 37503 54022 sw
rect 33288 54020 37503 54021
tri 37503 54020 37504 54021 sw
rect 33288 54019 37504 54020
tri 37504 54019 37505 54020 sw
rect 33288 54018 37505 54019
tri 37505 54018 37506 54019 sw
rect 33288 54017 37506 54018
tri 37506 54017 37507 54018 sw
rect 33288 54016 37507 54017
tri 37507 54016 37508 54017 sw
rect 33288 54015 37508 54016
tri 37508 54015 37509 54016 sw
rect 33288 54014 37509 54015
tri 37509 54014 37510 54015 sw
rect 33288 54013 37510 54014
tri 37510 54013 37511 54014 sw
rect 33288 54012 37511 54013
tri 37511 54012 37512 54013 sw
rect 33288 54011 37512 54012
tri 37512 54011 37513 54012 sw
rect 33288 54010 37513 54011
tri 37513 54010 37514 54011 sw
rect 33288 54009 37514 54010
tri 37514 54009 37515 54010 sw
rect 33288 54008 37515 54009
tri 37515 54008 37516 54009 sw
rect 33288 54007 37516 54008
tri 37516 54007 37517 54008 sw
rect 33288 54006 37517 54007
tri 37517 54006 37518 54007 sw
rect 33288 54005 37518 54006
tri 37518 54005 37519 54006 sw
rect 33288 54004 37519 54005
tri 37519 54004 37520 54005 sw
rect 33288 54003 37520 54004
tri 37520 54003 37521 54004 sw
rect 33288 54002 37521 54003
tri 37521 54002 37522 54003 sw
rect 33288 54001 37522 54002
tri 37522 54001 37523 54002 sw
rect 33288 54000 37523 54001
tri 37523 54000 37524 54001 sw
rect 33288 53999 37524 54000
tri 37524 53999 37525 54000 sw
rect 33288 53998 37525 53999
tri 37525 53998 37526 53999 sw
rect 33288 53997 37526 53998
tri 37526 53997 37527 53998 sw
rect 33288 53996 37527 53997
tri 37527 53996 37528 53997 sw
rect 33288 53995 37528 53996
tri 37528 53995 37529 53996 sw
rect 33288 53994 37529 53995
tri 37529 53994 37530 53995 sw
rect 33288 53993 37530 53994
tri 37530 53993 37531 53994 sw
rect 33288 53992 37531 53993
tri 37531 53992 37532 53993 sw
tri 33000 53704 33288 53992 sw
tri 33288 53731 33549 53992 ne
rect 33549 53991 37532 53992
tri 37532 53991 37533 53992 sw
tri 37729 53991 37830 54092 ne
rect 37830 53991 41972 54092
rect 33549 53731 37533 53991
rect 30000 53443 33288 53704
tri 33288 53443 33549 53704 sw
tri 33549 53443 33837 53731 ne
rect 33837 53694 37533 53731
tri 37533 53694 37830 53991 sw
tri 37830 53732 38089 53991 ne
rect 38089 53800 41972 53991
tri 41972 53800 42265 54093 sw
tri 42265 53991 42367 54093 ne
rect 42367 54092 44150 54093
tri 44150 54092 44246 54188 sw
tri 44442 54092 44538 54188 ne
rect 44538 54092 46324 54188
tri 46324 54092 46518 54286 sw
tri 46611 54092 46805 54286 ne
rect 46805 54187 50652 54286
tri 50652 54187 50963 54498 sw
tri 50963 54187 51274 54498 ne
rect 51274 54496 55212 54498
tri 55212 54496 55214 54498 sw
rect 51274 54494 55214 54496
tri 55214 54494 55216 54496 sw
rect 51274 54492 55216 54494
tri 55216 54492 55218 54494 sw
rect 51274 54490 55218 54492
tri 55218 54490 55220 54492 sw
rect 51274 54488 55220 54490
tri 55220 54488 55222 54490 sw
rect 51274 54486 55222 54488
tri 55222 54486 55224 54488 sw
rect 51274 54484 55224 54486
tri 55224 54484 55226 54486 sw
rect 51274 54482 55226 54484
tri 55226 54482 55228 54484 sw
rect 51274 54480 55228 54482
tri 55228 54480 55230 54482 sw
rect 51274 54478 55230 54480
tri 55230 54478 55232 54480 sw
rect 51274 54476 55232 54478
tri 55232 54476 55234 54478 sw
rect 51274 54474 55234 54476
tri 55234 54474 55236 54476 sw
rect 51274 54472 55236 54474
tri 55236 54472 55238 54474 sw
rect 51274 54470 55238 54472
tri 55238 54470 55240 54472 sw
rect 51274 54468 55240 54470
tri 55240 54468 55242 54470 sw
rect 51274 54466 55242 54468
tri 55242 54466 55244 54468 sw
rect 51274 54464 55244 54466
tri 55244 54464 55246 54466 sw
rect 51274 54462 55246 54464
tri 55246 54462 55248 54464 sw
rect 51274 54460 55248 54462
tri 55248 54460 55250 54462 sw
rect 51274 54458 55250 54460
tri 55250 54458 55252 54460 sw
rect 51274 54456 55252 54458
tri 55252 54456 55254 54458 sw
rect 51274 54454 55254 54456
tri 55254 54454 55256 54456 sw
rect 51274 54452 55256 54454
tri 55256 54452 55258 54454 sw
rect 51274 54450 55258 54452
tri 55258 54450 55260 54452 sw
rect 51274 54448 55260 54450
tri 55260 54448 55262 54450 sw
rect 51274 54446 55262 54448
tri 55262 54446 55264 54448 sw
rect 51274 54444 55264 54446
tri 55264 54444 55266 54446 sw
rect 51274 54442 55266 54444
tri 55266 54442 55268 54444 sw
rect 51274 54440 55268 54442
tri 55268 54440 55270 54442 sw
rect 51274 54438 55270 54440
tri 55270 54438 55272 54440 sw
rect 51274 54436 55272 54438
tri 55272 54436 55274 54438 sw
rect 51274 54434 55274 54436
tri 55274 54434 55276 54436 sw
rect 51274 54432 55276 54434
tri 55276 54432 55278 54434 sw
rect 51274 54430 55278 54432
tri 55278 54430 55280 54432 sw
rect 51274 54428 55280 54430
tri 55280 54428 55282 54430 sw
rect 51274 54426 55282 54428
tri 55282 54426 55284 54428 sw
rect 51274 54424 55284 54426
tri 55284 54424 55286 54426 sw
rect 51274 54422 55286 54424
tri 55286 54422 55288 54424 sw
rect 51274 54420 55288 54422
tri 55288 54420 55290 54422 sw
rect 51274 54418 55290 54420
tri 55290 54418 55292 54420 sw
rect 51274 54416 55292 54418
tri 55292 54416 55294 54418 sw
rect 51274 54414 55294 54416
tri 55294 54414 55296 54416 sw
rect 51274 54412 55296 54414
tri 55296 54412 55298 54414 sw
rect 51274 54410 55298 54412
tri 55298 54410 55300 54412 sw
rect 51274 54408 55300 54410
tri 55300 54408 55302 54410 sw
rect 51274 54406 55302 54408
tri 55302 54406 55304 54408 sw
rect 51274 54404 55304 54406
tri 55304 54404 55306 54406 sw
rect 51274 54402 55306 54404
tri 55306 54402 55308 54404 sw
rect 51274 54400 55308 54402
tri 55308 54400 55310 54402 sw
rect 51274 54398 55310 54400
tri 55310 54398 55312 54400 sw
rect 51274 54396 55312 54398
tri 55312 54396 55314 54398 sw
rect 51274 54394 55314 54396
tri 55314 54394 55316 54396 sw
rect 51274 54392 55316 54394
tri 55316 54392 55318 54394 sw
rect 51274 54390 55318 54392
tri 55318 54390 55320 54392 sw
rect 51274 54388 55320 54390
tri 55320 54388 55322 54390 sw
rect 51274 54386 55322 54388
tri 55322 54386 55324 54388 sw
rect 51274 54384 55324 54386
tri 55324 54384 55326 54386 sw
rect 51274 54382 55326 54384
tri 55326 54382 55328 54384 sw
rect 51274 54380 55328 54382
tri 55328 54380 55330 54382 sw
rect 51274 54378 55330 54380
tri 55330 54378 55332 54380 sw
rect 51274 54376 55332 54378
tri 55332 54376 55334 54378 sw
rect 51274 54374 55334 54376
tri 55334 54374 55336 54376 sw
rect 51274 54372 55336 54374
tri 55336 54372 55338 54374 sw
rect 51274 54370 55338 54372
tri 55338 54370 55340 54372 sw
rect 51274 54368 55340 54370
tri 55340 54368 55342 54370 sw
rect 51274 54366 55342 54368
tri 55342 54366 55344 54368 sw
rect 51274 54364 55344 54366
tri 55344 54364 55346 54366 sw
rect 51274 54362 55346 54364
tri 55346 54362 55348 54364 sw
rect 51274 54360 55348 54362
tri 55348 54360 55350 54362 sw
rect 51274 54358 55350 54360
tri 55350 54358 55352 54360 sw
rect 51274 54356 55352 54358
tri 55352 54356 55354 54358 sw
rect 51274 54354 55354 54356
tri 55354 54354 55356 54356 sw
rect 51274 54352 55356 54354
tri 55356 54352 55358 54354 sw
rect 51274 54351 55358 54352
tri 55358 54351 55359 54352 sw
rect 51274 54350 55359 54351
tri 55359 54350 55360 54351 sw
rect 51274 54349 55360 54350
tri 55360 54349 55361 54350 sw
rect 51274 54348 55361 54349
tri 55361 54348 55362 54349 sw
rect 51274 54347 55362 54348
tri 55362 54347 55363 54348 sw
rect 51274 54346 55363 54347
tri 55363 54346 55364 54347 sw
rect 51274 54345 55364 54346
tri 55364 54345 55365 54346 sw
rect 51274 54344 55365 54345
tri 55365 54344 55366 54345 sw
rect 51274 54343 55366 54344
tri 55366 54343 55367 54344 sw
rect 51274 54342 55367 54343
tri 55367 54342 55368 54343 sw
rect 51274 54341 55368 54342
tri 55368 54341 55369 54342 sw
rect 51274 54340 55369 54341
tri 55369 54340 55370 54341 sw
rect 51274 54339 55370 54340
tri 55370 54339 55371 54340 sw
rect 51274 54338 55371 54339
tri 55371 54338 55372 54339 sw
rect 51274 54337 55372 54338
tri 55372 54337 55373 54338 sw
rect 51274 54336 55373 54337
tri 55373 54336 55374 54337 sw
rect 51274 54335 55374 54336
tri 55374 54335 55375 54336 sw
rect 51274 54334 55375 54335
tri 55375 54334 55376 54335 sw
rect 51274 54333 55376 54334
tri 55376 54333 55377 54334 sw
rect 51274 54332 55377 54333
tri 55377 54332 55378 54333 sw
rect 51274 54331 55378 54332
tri 55378 54331 55379 54332 sw
rect 51274 54330 55379 54331
tri 55379 54330 55380 54331 sw
rect 51274 54329 55380 54330
tri 55380 54329 55381 54330 sw
rect 51274 54328 55381 54329
tri 55381 54328 55382 54329 sw
rect 51274 54327 55382 54328
tri 55382 54327 55383 54328 sw
rect 51274 54326 55383 54327
tri 55383 54326 55384 54327 sw
rect 51274 54325 55384 54326
tri 55384 54325 55385 54326 sw
rect 51274 54324 55385 54325
tri 55385 54324 55386 54325 sw
rect 51274 54323 55386 54324
tri 55386 54323 55387 54324 sw
rect 51274 54322 55387 54323
tri 55387 54322 55388 54323 sw
rect 51274 54321 55388 54322
tri 55388 54321 55389 54322 sw
rect 51274 54320 55389 54321
tri 55389 54320 55390 54321 sw
rect 51274 54319 55390 54320
tri 55390 54319 55391 54320 sw
rect 51274 54318 55391 54319
tri 55391 54318 55392 54319 sw
rect 51274 54317 55392 54318
tri 55392 54317 55393 54318 sw
rect 51274 54316 55393 54317
tri 55393 54316 55394 54317 sw
rect 51274 54315 55394 54316
tri 55394 54315 55395 54316 sw
rect 51274 54314 55395 54315
tri 55395 54314 55396 54315 sw
rect 51274 54313 55396 54314
tri 55396 54313 55397 54314 sw
rect 51274 54312 55397 54313
tri 55397 54312 55398 54313 sw
rect 51274 54311 55398 54312
tri 55398 54311 55399 54312 sw
rect 51274 54310 55399 54311
tri 55399 54310 55400 54311 sw
rect 51274 54309 55400 54310
tri 55400 54309 55401 54310 sw
rect 51274 54308 55401 54309
tri 55401 54308 55402 54309 sw
rect 51274 54307 55402 54308
tri 55402 54307 55403 54308 sw
rect 51274 54306 55403 54307
tri 55403 54306 55404 54307 sw
rect 51274 54305 55404 54306
tri 55404 54305 55405 54306 sw
rect 51274 54304 55405 54305
tri 55405 54304 55406 54305 sw
rect 51274 54303 55406 54304
tri 55406 54303 55407 54304 sw
rect 51274 54302 55407 54303
tri 55407 54302 55408 54303 sw
rect 51274 54301 55408 54302
tri 55408 54301 55409 54302 sw
rect 51274 54300 55409 54301
tri 55409 54300 55410 54301 sw
rect 51274 54299 55410 54300
tri 55410 54299 55411 54300 sw
rect 51274 54298 55411 54299
tri 55411 54298 55412 54299 sw
rect 51274 54297 55412 54298
tri 55412 54297 55413 54298 sw
rect 51274 54296 55413 54297
tri 55413 54296 55414 54297 sw
rect 51274 54295 55414 54296
tri 55414 54295 55415 54296 sw
rect 51274 54294 55415 54295
tri 55415 54294 55416 54295 sw
rect 51274 54293 55416 54294
tri 55416 54293 55417 54294 sw
rect 51274 54292 55417 54293
tri 55417 54292 55418 54293 sw
rect 51274 54291 55418 54292
tri 55418 54291 55419 54292 sw
rect 51274 54290 55419 54291
tri 55419 54290 55420 54291 sw
rect 51274 54289 55420 54290
tri 55420 54289 55421 54290 sw
rect 51274 54288 55421 54289
tri 55421 54288 55422 54289 sw
rect 51274 54287 55422 54288
tri 55422 54287 55423 54288 sw
rect 51274 54286 55423 54287
tri 55423 54286 55424 54287 sw
tri 55435 54286 55709 54560 ne
rect 55709 54286 57415 54560
tri 57415 54286 57689 54560 sw
tri 57699 54286 57973 54560 ne
rect 57973 54480 59679 54560
tri 59679 54480 59759 54560 sw
tri 59967 54480 60047 54560 ne
rect 60047 54480 61947 54560
tri 61947 54480 62027 54560 sw
tri 62233 54480 62313 54560 ne
rect 62313 54480 70613 54560
rect 57973 54286 59759 54480
tri 59759 54286 59953 54480 sw
tri 60047 54286 60241 54480 ne
rect 60241 54286 62027 54480
tri 62027 54286 62221 54480 sw
tri 62313 54286 62507 54480 ne
rect 62507 54286 70613 54480
rect 51274 54187 55424 54286
rect 46805 54092 50963 54187
rect 42367 53991 44246 54092
tri 44246 53991 44347 54092 sw
tri 44538 53991 44639 54092 ne
rect 44639 53991 46518 54092
tri 46518 53991 46619 54092 sw
tri 46805 53991 46906 54092 ne
rect 46906 53991 50963 54092
rect 38089 53732 42265 53800
rect 33837 53443 37830 53694
rect 30000 53231 33549 53443
tri 33549 53231 33761 53443 sw
tri 33837 53231 34049 53443 ne
rect 34049 53435 37830 53443
tri 37830 53435 38089 53694 sw
tri 38089 53469 38352 53732 ne
rect 38352 53698 42265 53732
tri 42265 53698 42367 53800 sw
tri 42367 53732 42626 53991 ne
rect 42626 53732 44347 53991
tri 44347 53732 44606 53991 sw
tri 44639 53732 44898 53991 ne
rect 44898 53732 46619 53991
tri 46619 53732 46878 53991 sw
tri 46906 53732 47165 53991 ne
rect 47165 53881 50963 53991
tri 50963 53881 51269 54187 sw
tri 51274 53991 51470 54187 ne
rect 51470 54001 55424 54187
tri 55424 54001 55709 54286 sw
tri 55709 54092 55903 54286 ne
rect 55903 54092 57689 54286
tri 57689 54092 57883 54286 sw
tri 57973 54092 58167 54286 ne
rect 58167 54180 59953 54286
tri 59953 54180 60059 54286 sw
tri 60241 54180 60347 54286 ne
rect 60347 54180 62221 54286
tri 62221 54180 62327 54286 sw
tri 62507 54180 62613 54286 ne
rect 62613 54180 70613 54286
rect 58167 54092 60059 54180
tri 60059 54092 60147 54180 sw
tri 60347 54092 60435 54180 ne
rect 60435 54092 62327 54180
tri 62327 54092 62415 54180 sw
tri 62613 54092 62701 54180 ne
rect 62701 54102 70613 54180
rect 70669 54102 71000 55302
rect 62701 54092 71000 54102
rect 51470 53991 55709 54001
rect 47165 53732 51269 53881
rect 38352 53469 42367 53698
rect 34049 53231 38089 53435
rect 30000 52943 33761 53231
tri 33761 52943 34049 53231 sw
tri 34049 52943 34337 53231 ne
rect 34337 53172 38089 53231
tri 38089 53172 38352 53435 sw
tri 38352 53172 38649 53469 ne
rect 38649 53465 42367 53469
tri 42367 53465 42600 53698 sw
tri 42626 53465 42893 53732 ne
rect 42893 53465 44606 53732
rect 38649 53172 42600 53465
tri 42600 53172 42893 53465 sw
tri 42893 53376 42982 53465 ne
rect 42982 53463 44606 53465
tri 44606 53463 44875 53732 sw
tri 44898 53463 45167 53732 ne
rect 45167 53463 46878 53732
rect 42982 53376 44875 53463
rect 34337 52943 38352 53172
rect 30000 52748 34049 52943
tri 30000 52654 30094 52748 ne
rect 30094 52655 34049 52748
tri 34049 52655 34337 52943 sw
tri 34337 52942 34338 52943 ne
rect 34338 52942 38352 52943
tri 34338 52748 34532 52942 ne
rect 34532 52875 38352 52942
tri 38352 52875 38649 53172 sw
tri 38649 52951 38870 53172 ne
rect 38870 53171 42893 53172
tri 42893 53171 42894 53172 sw
tri 42982 53171 43187 53376 ne
rect 43187 53171 44875 53376
tri 44875 53171 45167 53463 sw
tri 45167 53171 45459 53463 ne
rect 45459 53458 46878 53463
tri 46878 53458 47152 53732 sw
tri 47165 53458 47439 53732 ne
rect 47439 53682 51269 53732
tri 51269 53682 51468 53881 sw
tri 51470 53732 51729 53991 ne
rect 51729 53808 55709 53991
tri 55709 53808 55902 54001 sw
tri 55903 53991 56004 54092 ne
rect 56004 53991 57883 54092
rect 51729 53806 55902 53808
tri 55902 53806 55904 53808 sw
rect 51729 53804 55904 53806
tri 55904 53804 55906 53806 sw
rect 51729 53802 55906 53804
tri 55906 53802 55908 53804 sw
rect 51729 53800 55908 53802
tri 55908 53800 55910 53802 sw
rect 51729 53798 55910 53800
tri 55910 53798 55912 53800 sw
rect 51729 53796 55912 53798
tri 55912 53796 55914 53798 sw
rect 51729 53794 55914 53796
tri 55914 53794 55916 53796 sw
rect 51729 53792 55916 53794
tri 55916 53792 55918 53794 sw
rect 51729 53790 55918 53792
tri 55918 53790 55920 53792 sw
rect 51729 53788 55920 53790
tri 55920 53788 55922 53790 sw
rect 51729 53786 55922 53788
tri 55922 53786 55924 53788 sw
rect 51729 53784 55924 53786
tri 55924 53784 55926 53786 sw
rect 51729 53782 55926 53784
tri 55926 53782 55928 53784 sw
rect 51729 53780 55928 53782
tri 55928 53780 55930 53782 sw
rect 51729 53778 55930 53780
tri 55930 53778 55932 53780 sw
rect 51729 53776 55932 53778
tri 55932 53776 55934 53778 sw
rect 51729 53774 55934 53776
tri 55934 53774 55936 53776 sw
rect 51729 53772 55936 53774
tri 55936 53772 55938 53774 sw
rect 51729 53770 55938 53772
tri 55938 53770 55940 53772 sw
rect 51729 53768 55940 53770
tri 55940 53768 55942 53770 sw
rect 51729 53766 55942 53768
tri 55942 53766 55944 53768 sw
rect 51729 53764 55944 53766
tri 55944 53764 55946 53766 sw
rect 51729 53762 55946 53764
tri 55946 53762 55948 53764 sw
rect 51729 53760 55948 53762
tri 55948 53760 55950 53762 sw
rect 51729 53758 55950 53760
tri 55950 53758 55952 53760 sw
rect 51729 53756 55952 53758
tri 55952 53756 55954 53758 sw
rect 51729 53754 55954 53756
tri 55954 53754 55956 53756 sw
rect 51729 53752 55956 53754
tri 55956 53752 55958 53754 sw
rect 51729 53750 55958 53752
tri 55958 53750 55960 53752 sw
rect 51729 53748 55960 53750
tri 55960 53748 55962 53750 sw
rect 51729 53746 55962 53748
tri 55962 53746 55964 53748 sw
rect 51729 53744 55964 53746
tri 55964 53744 55966 53746 sw
rect 51729 53742 55966 53744
tri 55966 53742 55968 53744 sw
rect 51729 53740 55968 53742
tri 55968 53740 55970 53742 sw
rect 51729 53738 55970 53740
tri 55970 53738 55972 53740 sw
rect 51729 53736 55972 53738
tri 55972 53736 55974 53738 sw
rect 51729 53734 55974 53736
tri 55974 53734 55976 53736 sw
rect 51729 53732 55976 53734
tri 55976 53732 55978 53734 sw
tri 56004 53732 56263 53991 ne
rect 56263 53896 57883 53991
tri 57883 53896 58079 54092 sw
tri 58167 53896 58363 54092 ne
rect 58363 53991 60147 54092
tri 60147 53991 60248 54092 sw
tri 60435 53991 60536 54092 ne
rect 60536 54000 62415 54092
tri 62415 54000 62507 54092 sw
tri 62701 54000 62793 54092 ne
rect 62793 54000 71000 54092
rect 60536 53991 62507 54000
tri 62507 53991 62516 54000 sw
rect 58363 53896 60248 53991
rect 56263 53732 58079 53896
tri 58079 53732 58243 53896 sw
tri 58363 53732 58527 53896 ne
rect 58527 53800 60248 53896
tri 60248 53800 60439 53991 sw
tri 60536 53800 60727 53991 ne
rect 60727 53800 62516 53991
tri 62516 53800 62707 53991 sw
rect 58527 53732 60439 53800
tri 60439 53732 60507 53800 sw
tri 60727 53732 60795 53800 ne
rect 60795 53732 71000 53800
rect 47439 53458 51468 53682
rect 45459 53171 47152 53458
tri 47152 53171 47439 53458 sw
tri 47439 53171 47726 53458 ne
rect 47726 53423 51468 53458
tri 51468 53423 51727 53682 sw
tri 51729 53563 51898 53732 ne
rect 51898 53563 55978 53732
rect 47726 53252 51727 53423
tri 51727 53252 51898 53423 sw
tri 51898 53252 52209 53563 ne
rect 52209 53447 55978 53563
tri 55978 53447 56263 53732 sw
tri 56263 53529 56466 53732 ne
rect 56466 53529 58243 53732
rect 52209 53252 56263 53447
rect 47726 53171 51898 53252
rect 38870 52951 42894 53171
rect 34532 52748 38649 52875
rect 30094 52654 34337 52655
tri 29800 52360 30094 52654 sw
tri 30094 52453 30295 52654 ne
rect 30295 52460 34337 52654
tri 34337 52460 34532 52655 sw
tri 34532 52511 34769 52748 ne
rect 34769 52654 38649 52748
tri 38649 52654 38870 52875 sw
tri 38870 52654 39167 52951 ne
rect 39167 52878 42894 52951
tri 42894 52878 43187 53171 sw
tri 43187 52880 43478 53171 ne
rect 43478 52880 45167 53171
tri 45167 52880 45458 53171 sw
tri 45459 52880 45750 53171 ne
rect 45750 53167 47439 53171
tri 47439 53167 47443 53171 sw
tri 47726 53167 47730 53171 ne
rect 47730 53167 51898 53171
rect 45750 52880 47443 53167
tri 47443 52880 47730 53167 sw
tri 47730 52880 48017 53167 ne
rect 48017 52945 51898 53167
tri 51898 52945 52205 53252 sw
tri 52209 53171 52290 53252 ne
rect 52290 53244 56263 53252
tri 56263 53244 56466 53447 sw
tri 56466 53244 56751 53529 ne
rect 56751 53527 58243 53529
tri 58243 53527 58448 53732 sw
tri 58527 53527 58732 53732 ne
rect 58732 53527 60507 53732
rect 56751 53244 58448 53527
rect 52290 53171 56466 53244
rect 48017 52880 52205 52945
rect 39167 52654 43187 52878
rect 34769 52511 38870 52654
rect 30295 52453 34532 52460
rect 26800 52159 30094 52360
tri 30094 52159 30295 52360 sw
tri 30295 52159 30589 52453 ne
rect 30589 52223 34532 52453
tri 34532 52223 34769 52460 sw
tri 34769 52223 35057 52511 ne
rect 35057 52357 38870 52511
tri 38870 52357 39167 52654 sw
tri 39167 52426 39395 52654 ne
rect 39395 52587 43187 52654
tri 43187 52587 43478 52878 sw
tri 43478 52653 43705 52880 ne
rect 43705 52653 45458 52880
tri 45458 52653 45685 52880 sw
tri 45750 52653 45977 52880 ne
rect 45977 52653 47730 52880
tri 47730 52653 47957 52880 sw
tri 48017 52653 48244 52880 ne
rect 48244 52860 52205 52880
tri 52205 52860 52290 52945 sw
tri 52290 52880 52581 53171 ne
rect 52581 52960 56466 53171
tri 56466 52960 56750 53244 sw
tri 56751 53167 56828 53244 ne
rect 56828 53243 58448 53244
tri 58448 53243 58732 53527 sw
tri 58732 53243 59016 53527 ne
rect 59016 53512 60507 53527
tri 60507 53512 60727 53732 sw
tri 60795 53512 61015 53732 ne
rect 61015 53722 71000 53732
rect 61015 53512 70613 53722
rect 59016 53243 60727 53512
tri 60727 53243 60996 53512 sw
tri 61015 53243 61284 53512 ne
rect 61284 53243 70613 53512
rect 56828 53167 58732 53243
rect 52581 52958 56750 52960
tri 56750 52958 56752 52960 sw
rect 52581 52956 56752 52958
tri 56752 52956 56754 52958 sw
rect 52581 52954 56754 52956
tri 56754 52954 56756 52956 sw
rect 52581 52952 56756 52954
tri 56756 52952 56758 52954 sw
rect 52581 52950 56758 52952
tri 56758 52950 56760 52952 sw
rect 52581 52948 56760 52950
tri 56760 52948 56762 52950 sw
rect 52581 52946 56762 52948
tri 56762 52946 56764 52948 sw
rect 52581 52944 56764 52946
tri 56764 52944 56766 52946 sw
rect 52581 52942 56766 52944
tri 56766 52942 56768 52944 sw
rect 52581 52940 56768 52942
tri 56768 52940 56770 52942 sw
rect 52581 52938 56770 52940
tri 56770 52938 56772 52940 sw
rect 52581 52936 56772 52938
tri 56772 52936 56774 52938 sw
rect 52581 52934 56774 52936
tri 56774 52934 56776 52936 sw
rect 52581 52932 56776 52934
tri 56776 52932 56778 52934 sw
rect 52581 52930 56778 52932
tri 56778 52930 56780 52932 sw
rect 52581 52928 56780 52930
tri 56780 52928 56782 52930 sw
rect 52581 52926 56782 52928
tri 56782 52926 56784 52928 sw
rect 52581 52924 56784 52926
tri 56784 52924 56786 52926 sw
rect 52581 52922 56786 52924
tri 56786 52922 56788 52924 sw
rect 52581 52920 56788 52922
tri 56788 52920 56790 52922 sw
rect 52581 52918 56790 52920
tri 56790 52918 56792 52920 sw
rect 52581 52916 56792 52918
tri 56792 52916 56794 52918 sw
rect 52581 52914 56794 52916
tri 56794 52914 56796 52916 sw
rect 52581 52912 56796 52914
tri 56796 52912 56798 52914 sw
rect 52581 52910 56798 52912
tri 56798 52910 56800 52912 sw
rect 52581 52908 56800 52910
tri 56800 52908 56802 52910 sw
rect 52581 52906 56802 52908
tri 56802 52906 56804 52908 sw
rect 52581 52904 56804 52906
tri 56804 52904 56806 52906 sw
rect 52581 52902 56806 52904
tri 56806 52902 56808 52904 sw
rect 52581 52900 56808 52902
tri 56808 52900 56810 52902 sw
rect 52581 52898 56810 52900
tri 56810 52898 56812 52900 sw
rect 52581 52896 56812 52898
tri 56812 52896 56814 52898 sw
rect 52581 52894 56814 52896
tri 56814 52894 56816 52896 sw
rect 52581 52892 56816 52894
tri 56816 52892 56818 52894 sw
rect 52581 52890 56818 52892
tri 56818 52890 56820 52892 sw
rect 52581 52888 56820 52890
tri 56820 52888 56822 52890 sw
rect 52581 52886 56822 52888
tri 56822 52886 56824 52888 sw
rect 52581 52884 56824 52886
tri 56824 52884 56826 52886 sw
rect 52581 52882 56826 52884
tri 56826 52882 56828 52884 sw
tri 56828 52882 57113 53167 ne
rect 57113 53164 58732 53167
tri 58732 53164 58811 53243 sw
tri 59016 53164 59095 53243 ne
rect 59095 53171 60996 53243
tri 60996 53171 61068 53243 sw
tri 61284 53171 61356 53243 ne
rect 61356 53171 70613 53243
rect 59095 53168 61068 53171
tri 61068 53168 61071 53171 sw
tri 61356 53168 61359 53171 ne
rect 61359 53168 70613 53171
rect 59095 53164 61071 53168
rect 57113 52882 58811 53164
rect 52581 52880 56828 52882
rect 48244 52653 52290 52860
rect 39395 52426 43478 52587
rect 35057 52223 39167 52357
rect 30589 52222 34769 52223
tri 34769 52222 34770 52223 sw
tri 35057 52222 35058 52223 ne
rect 35058 52222 39167 52223
rect 30589 52159 34770 52222
rect 26800 51865 30295 52159
tri 30295 51865 30589 52159 sw
tri 30589 51910 30838 52159 ne
rect 30838 51934 34770 52159
tri 34770 51934 35058 52222 sw
tri 35058 51934 35346 52222 ne
rect 35346 52129 39167 52222
tri 39167 52129 39395 52357 sw
tri 39395 52129 39692 52426 ne
rect 39692 52360 43478 52426
tri 43478 52360 43705 52587 sw
tri 43705 52422 43936 52653 ne
rect 43936 52500 45685 52653
tri 45685 52500 45838 52653 sw
tri 45977 52500 46130 52653 ne
rect 46130 52500 47957 52653
rect 43936 52422 45838 52500
rect 39692 52129 43705 52360
tri 43705 52129 43936 52360 sw
tri 43936 52129 44229 52422 ne
rect 44229 52208 45838 52422
tri 45838 52208 46130 52500 sw
tri 46130 52208 46422 52500 ne
rect 46422 52415 47957 52500
tri 47957 52415 48195 52653 sw
tri 48244 52415 48482 52653 ne
rect 48482 52570 52290 52653
tri 52290 52570 52580 52860 sw
tri 52581 52653 52808 52880 ne
rect 52808 52653 56828 52880
rect 48482 52415 52580 52570
rect 46422 52208 48195 52415
rect 44229 52129 46130 52208
rect 35346 51934 39395 52129
rect 30838 51910 35058 51934
rect 26800 51616 30589 51865
tri 30589 51616 30838 51865 sw
tri 30838 51704 31044 51910 ne
rect 31044 51704 35058 51910
rect 26800 51410 30838 51616
tri 30838 51410 31044 51616 sw
tri 31044 51615 31133 51704 ne
rect 31133 51646 35058 51704
tri 35058 51646 35346 51934 sw
tri 35346 51898 35382 51934 ne
rect 35382 51898 39395 51934
rect 31133 51615 35346 51646
tri 31133 51410 31338 51615 ne
rect 31338 51610 35346 51615
tri 35346 51610 35382 51646 sw
tri 35382 51610 35670 51898 ne
rect 35670 51832 39395 51898
tri 39395 51832 39692 52129 sw
tri 39692 52128 39693 52129 ne
rect 39693 52128 43936 52129
rect 35670 51831 39692 51832
tri 39692 51831 39693 51832 sw
tri 39693 51831 39990 52128 ne
rect 39990 51836 43936 52128
tri 43936 51836 44229 52129 sw
tri 44229 52128 44230 52129 ne
rect 44230 52128 46130 52129
tri 46130 52128 46210 52208 sw
tri 46422 52128 46502 52208 ne
rect 46502 52128 48195 52208
tri 48195 52128 48482 52415 sw
tri 48482 52128 48769 52415 ne
rect 48769 52350 52580 52415
tri 52580 52350 52800 52570 sw
tri 52808 52449 53012 52653 ne
rect 53012 52598 56828 52653
tri 56828 52598 57112 52882 sw
tri 57113 52653 57342 52882 ne
rect 57342 52880 58811 52882
tri 58811 52880 59095 53164 sw
tri 59095 52880 59379 53164 ne
rect 59379 52880 61071 53164
tri 61071 52880 61359 53168 sw
tri 61359 52880 61647 53168 ne
rect 61647 52880 70613 53168
rect 57342 52653 59095 52880
tri 59095 52653 59322 52880 sw
tri 59379 52653 59606 52880 ne
rect 59606 52653 61359 52880
tri 61359 52653 61586 52880 sw
tri 61647 52653 61874 52880 ne
rect 61874 52653 70613 52880
rect 53012 52449 57112 52598
rect 48769 52138 52800 52350
tri 52800 52138 53012 52350 sw
tri 53012 52138 53323 52449 ne
rect 53323 52369 57112 52449
tri 57112 52369 57341 52598 sw
tri 57342 52500 57495 52653 ne
rect 57495 52500 59322 52653
rect 53323 52367 57341 52369
tri 57341 52367 57343 52369 sw
rect 53323 52365 57343 52367
tri 57343 52365 57345 52367 sw
rect 53323 52363 57345 52365
tri 57345 52363 57347 52365 sw
rect 53323 52361 57347 52363
tri 57347 52361 57349 52363 sw
rect 53323 52359 57349 52361
tri 57349 52359 57351 52361 sw
rect 53323 52357 57351 52359
tri 57351 52357 57353 52359 sw
rect 53323 52355 57353 52357
tri 57353 52355 57355 52357 sw
rect 53323 52353 57355 52355
tri 57355 52353 57357 52355 sw
rect 53323 52351 57357 52353
tri 57357 52351 57359 52353 sw
rect 53323 52349 57359 52351
tri 57359 52349 57361 52351 sw
rect 53323 52347 57361 52349
tri 57361 52347 57363 52349 sw
rect 53323 52345 57363 52347
tri 57363 52345 57365 52347 sw
rect 53323 52343 57365 52345
tri 57365 52343 57367 52345 sw
rect 53323 52341 57367 52343
tri 57367 52341 57369 52343 sw
rect 53323 52339 57369 52341
tri 57369 52339 57371 52341 sw
rect 53323 52337 57371 52339
tri 57371 52337 57373 52339 sw
rect 53323 52335 57373 52337
tri 57373 52335 57375 52337 sw
rect 53323 52333 57375 52335
tri 57375 52333 57377 52335 sw
rect 53323 52331 57377 52333
tri 57377 52331 57379 52333 sw
rect 53323 52329 57379 52331
tri 57379 52329 57381 52331 sw
rect 53323 52327 57381 52329
tri 57381 52327 57383 52329 sw
rect 53323 52325 57383 52327
tri 57383 52325 57385 52327 sw
rect 53323 52323 57385 52325
tri 57385 52323 57387 52325 sw
rect 53323 52321 57387 52323
tri 57387 52321 57389 52323 sw
rect 53323 52319 57389 52321
tri 57389 52319 57391 52321 sw
rect 53323 52317 57391 52319
tri 57391 52317 57393 52319 sw
rect 53323 52315 57393 52317
tri 57393 52315 57395 52317 sw
rect 53323 52313 57395 52315
tri 57395 52313 57397 52315 sw
rect 53323 52311 57397 52313
tri 57397 52311 57399 52313 sw
rect 53323 52309 57399 52311
tri 57399 52309 57401 52311 sw
rect 53323 52307 57401 52309
tri 57401 52307 57403 52309 sw
rect 53323 52305 57403 52307
tri 57403 52305 57405 52307 sw
rect 53323 52303 57405 52305
tri 57405 52303 57407 52305 sw
rect 53323 52301 57407 52303
tri 57407 52301 57409 52303 sw
rect 53323 52299 57409 52301
tri 57409 52299 57411 52301 sw
rect 53323 52297 57411 52299
tri 57411 52297 57413 52299 sw
rect 53323 52295 57413 52297
tri 57413 52295 57415 52297 sw
rect 53323 52293 57415 52295
tri 57415 52293 57417 52295 sw
tri 57495 52293 57702 52500 ne
rect 57702 52484 59322 52500
tri 59322 52484 59491 52653 sw
tri 59606 52580 59679 52653 ne
rect 59679 52580 61586 52653
tri 61586 52580 61659 52653 sw
tri 61874 52580 61947 52653 ne
rect 61947 52580 70613 52653
tri 59679 52512 59747 52580 ne
rect 59747 52512 61659 52580
tri 61659 52512 61727 52580 sw
tri 61947 52512 62015 52580 ne
rect 62015 52522 70613 52580
rect 70669 52522 71000 53722
rect 62015 52512 71000 52522
tri 59747 52500 59759 52512 ne
rect 59759 52500 61727 52512
tri 61727 52500 61739 52512 sw
tri 62015 52500 62027 52512 ne
rect 62027 52500 71000 52512
tri 59759 52484 59775 52500 ne
rect 59775 52484 61739 52500
rect 57702 52293 59491 52484
rect 53323 52138 57417 52293
rect 48769 52128 53012 52138
rect 39990 51835 44229 51836
tri 44229 51835 44230 51836 sw
tri 44230 51835 44523 52128 ne
rect 44523 51836 46210 52128
tri 46210 51836 46502 52128 sw
tri 46502 51836 46794 52128 ne
rect 46794 51841 48482 52128
tri 48482 51841 48769 52128 sw
tri 48769 51841 49056 52128 ne
rect 49056 51841 53012 52128
rect 46794 51836 48769 51841
rect 44523 51835 46502 51836
rect 39990 51831 44230 51835
rect 35670 51610 39693 51831
rect 31338 51410 35382 51610
tri 26600 51120 26800 51320 sw
tri 26800 51120 27090 51410 ne
rect 27090 51120 31044 51410
rect 25200 50941 26800 51120
tri 26800 50941 26979 51120 sw
tri 27090 50941 27269 51120 ne
rect 27269 51116 31044 51120
tri 31044 51116 31338 51410 sw
tri 31338 51220 31528 51410 ne
rect 31528 51322 35382 51410
tri 35382 51322 35670 51610 sw
tri 35670 51508 35772 51610 ne
rect 35772 51534 39693 51610
tri 39693 51534 39990 51831 sw
tri 39990 51618 40203 51831 ne
rect 40203 51618 44230 51831
rect 35772 51508 39990 51534
rect 31528 51220 35670 51322
tri 35670 51220 35772 51322 sw
tri 35772 51320 35960 51508 ne
rect 35960 51321 39990 51508
tri 39990 51321 40203 51534 sw
tri 40203 51321 40500 51618 ne
rect 40500 51542 44230 51618
tri 44230 51542 44523 51835 sw
tri 44523 51614 44744 51835 ne
rect 44744 51614 46502 51835
rect 40500 51321 44523 51542
tri 44523 51321 44744 51542 sw
tri 44744 51321 45037 51614 ne
rect 45037 51612 46502 51614
tri 46502 51612 46726 51836 sw
tri 46794 51612 47018 51836 ne
rect 47018 51612 48769 51836
rect 45037 51321 46726 51612
rect 35960 51320 40203 51321
rect 27269 50941 31338 51116
rect 25200 50740 26979 50941
tri 25200 50651 25289 50740 ne
rect 25289 50651 26979 50740
tri 26979 50651 27269 50941 sw
tri 27269 50651 27559 50941 ne
rect 27559 50926 31338 50941
tri 31338 50926 31528 51116 sw
tri 31528 50926 31822 51220 ne
rect 31822 51219 35772 51220
tri 35772 51219 35773 51220 sw
rect 31822 51218 35773 51219
tri 35773 51218 35774 51219 sw
rect 31822 51217 35774 51218
tri 35774 51217 35775 51218 sw
rect 31822 51216 35775 51217
tri 35775 51216 35776 51217 sw
rect 31822 51215 35776 51216
tri 35776 51215 35777 51216 sw
rect 31822 51214 35777 51215
tri 35777 51214 35778 51215 sw
rect 31822 51213 35778 51214
tri 35778 51213 35779 51214 sw
rect 31822 51212 35779 51213
tri 35779 51212 35780 51213 sw
rect 31822 51211 35780 51212
tri 35780 51211 35781 51212 sw
rect 31822 51210 35781 51211
tri 35781 51210 35782 51211 sw
rect 31822 51209 35782 51210
tri 35782 51209 35783 51210 sw
rect 31822 51208 35783 51209
tri 35783 51208 35784 51209 sw
rect 31822 51207 35784 51208
tri 35784 51207 35785 51208 sw
rect 31822 51206 35785 51207
tri 35785 51206 35786 51207 sw
rect 31822 51205 35786 51206
tri 35786 51205 35787 51206 sw
rect 31822 51204 35787 51205
tri 35787 51204 35788 51205 sw
rect 31822 51203 35788 51204
tri 35788 51203 35789 51204 sw
rect 31822 51202 35789 51203
tri 35789 51202 35790 51203 sw
rect 31822 51201 35790 51202
tri 35790 51201 35791 51202 sw
rect 31822 51200 35791 51201
tri 35791 51200 35792 51201 sw
rect 31822 51199 35792 51200
tri 35792 51199 35793 51200 sw
rect 31822 51198 35793 51199
tri 35793 51198 35794 51199 sw
rect 31822 51197 35794 51198
tri 35794 51197 35795 51198 sw
rect 31822 51196 35795 51197
tri 35795 51196 35796 51197 sw
rect 31822 51195 35796 51196
tri 35796 51195 35797 51196 sw
rect 31822 51194 35797 51195
tri 35797 51194 35798 51195 sw
rect 31822 51193 35798 51194
tri 35798 51193 35799 51194 sw
rect 31822 51192 35799 51193
tri 35799 51192 35800 51193 sw
rect 31822 51191 35800 51192
tri 35800 51191 35801 51192 sw
rect 31822 51190 35801 51191
tri 35801 51190 35802 51191 sw
rect 31822 51189 35802 51190
tri 35802 51189 35803 51190 sw
rect 31822 51188 35803 51189
tri 35803 51188 35804 51189 sw
rect 31822 51187 35804 51188
tri 35804 51187 35805 51188 sw
rect 31822 51186 35805 51187
tri 35805 51186 35806 51187 sw
rect 31822 51185 35806 51186
tri 35806 51185 35807 51186 sw
rect 31822 51184 35807 51185
tri 35807 51184 35808 51185 sw
rect 31822 51183 35808 51184
tri 35808 51183 35809 51184 sw
rect 31822 51182 35809 51183
tri 35809 51182 35810 51183 sw
rect 31822 51181 35810 51182
tri 35810 51181 35811 51182 sw
rect 31822 51180 35811 51181
tri 35811 51180 35812 51181 sw
rect 31822 51179 35812 51180
tri 35812 51179 35813 51180 sw
rect 31822 51178 35813 51179
tri 35813 51178 35814 51179 sw
rect 31822 51177 35814 51178
tri 35814 51177 35815 51178 sw
rect 31822 51176 35815 51177
tri 35815 51176 35816 51177 sw
rect 31822 51175 35816 51176
tri 35816 51175 35817 51176 sw
rect 31822 51174 35817 51175
tri 35817 51174 35818 51175 sw
rect 31822 51173 35818 51174
tri 35818 51173 35819 51174 sw
rect 31822 51172 35819 51173
tri 35819 51172 35820 51173 sw
rect 31822 51171 35820 51172
tri 35820 51171 35821 51172 sw
rect 31822 51170 35821 51171
tri 35821 51170 35822 51171 sw
rect 31822 51169 35822 51170
tri 35822 51169 35823 51170 sw
rect 31822 51168 35823 51169
tri 35823 51168 35824 51169 sw
rect 31822 51167 35824 51168
tri 35824 51167 35825 51168 sw
rect 31822 51166 35825 51167
tri 35825 51166 35826 51167 sw
rect 31822 51165 35826 51166
tri 35826 51165 35827 51166 sw
rect 31822 51164 35827 51165
tri 35827 51164 35828 51165 sw
rect 31822 51163 35828 51164
tri 35828 51163 35829 51164 sw
rect 31822 51162 35829 51163
tri 35829 51162 35830 51163 sw
rect 31822 51161 35830 51162
tri 35830 51161 35831 51162 sw
rect 31822 51160 35831 51161
tri 35831 51160 35832 51161 sw
rect 31822 51159 35832 51160
tri 35832 51159 35833 51160 sw
rect 31822 51158 35833 51159
tri 35833 51158 35834 51159 sw
rect 31822 51157 35834 51158
tri 35834 51157 35835 51158 sw
rect 31822 51156 35835 51157
tri 35835 51156 35836 51157 sw
rect 31822 51155 35836 51156
tri 35836 51155 35837 51156 sw
rect 31822 51154 35837 51155
tri 35837 51154 35838 51155 sw
rect 31822 51153 35838 51154
tri 35838 51153 35839 51154 sw
rect 31822 51152 35839 51153
tri 35839 51152 35840 51153 sw
rect 31822 51151 35840 51152
tri 35840 51151 35841 51152 sw
rect 31822 51150 35841 51151
tri 35841 51150 35842 51151 sw
rect 31822 51149 35842 51150
tri 35842 51149 35843 51150 sw
rect 31822 51148 35843 51149
tri 35843 51148 35844 51149 sw
rect 31822 51147 35844 51148
tri 35844 51147 35845 51148 sw
rect 31822 51146 35845 51147
tri 35845 51146 35846 51147 sw
rect 31822 51145 35846 51146
tri 35846 51145 35847 51146 sw
rect 31822 51144 35847 51145
tri 35847 51144 35848 51145 sw
rect 31822 51143 35848 51144
tri 35848 51143 35849 51144 sw
rect 31822 51142 35849 51143
tri 35849 51142 35850 51143 sw
rect 31822 51141 35850 51142
tri 35850 51141 35851 51142 sw
rect 31822 51140 35851 51141
tri 35851 51140 35852 51141 sw
rect 31822 51139 35852 51140
tri 35852 51139 35853 51140 sw
rect 31822 51138 35853 51139
tri 35853 51138 35854 51139 sw
rect 31822 51137 35854 51138
tri 35854 51137 35855 51138 sw
rect 31822 51136 35855 51137
tri 35855 51136 35856 51137 sw
rect 31822 51135 35856 51136
tri 35856 51135 35857 51136 sw
rect 31822 51134 35857 51135
tri 35857 51134 35858 51135 sw
rect 31822 51133 35858 51134
tri 35858 51133 35859 51134 sw
rect 31822 51132 35859 51133
tri 35859 51132 35860 51133 sw
rect 31822 51131 35860 51132
tri 35860 51131 35861 51132 sw
rect 31822 51130 35861 51131
tri 35861 51130 35862 51131 sw
rect 31822 51129 35862 51130
tri 35862 51129 35863 51130 sw
rect 31822 51128 35863 51129
tri 35863 51128 35864 51129 sw
rect 31822 51127 35864 51128
tri 35864 51127 35865 51128 sw
rect 31822 51126 35865 51127
tri 35865 51126 35866 51127 sw
rect 31822 51125 35866 51126
tri 35866 51125 35867 51126 sw
rect 31822 51124 35867 51125
tri 35867 51124 35868 51125 sw
rect 31822 51123 35868 51124
tri 35868 51123 35869 51124 sw
rect 31822 51122 35869 51123
tri 35869 51122 35870 51123 sw
rect 31822 51121 35870 51122
tri 35870 51121 35871 51122 sw
rect 31822 51120 35871 51121
tri 35871 51120 35872 51121 sw
rect 31822 51119 35872 51120
tri 35872 51119 35873 51120 sw
rect 31822 51118 35873 51119
tri 35873 51118 35874 51119 sw
rect 31822 51117 35874 51118
tri 35874 51117 35875 51118 sw
rect 31822 51116 35875 51117
tri 35875 51116 35876 51117 sw
rect 31822 51115 35876 51116
tri 35876 51115 35877 51116 sw
rect 31822 51114 35877 51115
tri 35877 51114 35878 51115 sw
rect 31822 51113 35878 51114
tri 35878 51113 35879 51114 sw
rect 31822 51112 35879 51113
tri 35879 51112 35880 51113 sw
rect 31822 51111 35880 51112
tri 35880 51111 35881 51112 sw
rect 31822 51110 35881 51111
tri 35881 51110 35882 51111 sw
rect 31822 51109 35882 51110
tri 35882 51109 35883 51110 sw
rect 31822 51108 35883 51109
tri 35883 51108 35884 51109 sw
rect 31822 51107 35884 51108
tri 35884 51107 35885 51108 sw
rect 31822 51106 35885 51107
tri 35885 51106 35886 51107 sw
rect 31822 51105 35886 51106
tri 35886 51105 35887 51106 sw
rect 31822 51104 35887 51105
tri 35887 51104 35888 51105 sw
rect 31822 51103 35888 51104
tri 35888 51103 35889 51104 sw
rect 31822 51102 35889 51103
tri 35889 51102 35890 51103 sw
rect 31822 51101 35890 51102
tri 35890 51101 35891 51102 sw
rect 31822 51100 35891 51101
tri 35891 51100 35892 51101 sw
rect 31822 51099 35892 51100
tri 35892 51099 35893 51100 sw
rect 31822 51098 35893 51099
tri 35893 51098 35894 51099 sw
rect 31822 51097 35894 51098
tri 35894 51097 35895 51098 sw
rect 31822 51096 35895 51097
tri 35895 51096 35896 51097 sw
rect 31822 51095 35896 51096
tri 35896 51095 35897 51096 sw
rect 31822 51094 35897 51095
tri 35897 51094 35898 51095 sw
rect 31822 51093 35898 51094
tri 35898 51093 35899 51094 sw
rect 31822 51092 35899 51093
tri 35899 51092 35900 51093 sw
rect 31822 51091 35900 51092
tri 35900 51091 35901 51092 sw
rect 31822 51090 35901 51091
tri 35901 51090 35902 51091 sw
rect 31822 51089 35902 51090
tri 35902 51089 35903 51090 sw
rect 31822 51088 35903 51089
tri 35903 51088 35904 51089 sw
rect 31822 51087 35904 51088
tri 35904 51087 35905 51088 sw
rect 31822 51086 35905 51087
tri 35905 51086 35906 51087 sw
rect 31822 51085 35906 51086
tri 35906 51085 35907 51086 sw
rect 31822 51084 35907 51085
tri 35907 51084 35908 51085 sw
rect 31822 51083 35908 51084
tri 35908 51083 35909 51084 sw
rect 31822 51082 35909 51083
tri 35909 51082 35910 51083 sw
rect 31822 51081 35910 51082
tri 35910 51081 35911 51082 sw
tri 35960 51081 36199 51320 ne
rect 36199 51081 40203 51320
rect 31822 50926 35911 51081
rect 27559 50651 31528 50926
tri 25000 50451 25200 50651 sw
tri 25289 50451 25489 50651 ne
rect 25489 50650 27269 50651
tri 27269 50650 27270 50651 sw
tri 27559 50650 27560 50651 ne
rect 27560 50650 31528 50651
rect 25489 50451 27270 50650
rect 23600 50262 25200 50451
tri 25200 50262 25389 50451 sw
tri 25489 50262 25678 50451 ne
rect 25678 50360 27270 50451
tri 27270 50360 27560 50650 sw
tri 27560 50360 27850 50650 ne
rect 27850 50632 31528 50650
tri 31528 50632 31822 50926 sw
tri 31822 50651 32097 50926 ne
rect 32097 50793 35911 50926
tri 35911 50793 36199 51081 sw
tri 36199 51014 36266 51081 ne
rect 36266 51024 40203 51081
tri 40203 51024 40500 51321 sw
tri 40500 51312 40509 51321 ne
rect 40509 51320 44744 51321
tri 44744 51320 44745 51321 sw
tri 45037 51320 45038 51321 ne
rect 45038 51320 46726 51321
tri 46726 51320 47018 51612 sw
tri 47018 51320 47310 51612 ne
rect 47310 51607 48769 51612
tri 48769 51607 49003 51841 sw
tri 49056 51607 49290 51841 ne
rect 49290 51833 53012 51841
tri 53012 51833 53317 52138 sw
tri 53323 52124 53337 52138 ne
rect 53337 52124 57417 52138
rect 49290 51813 53317 51833
tri 53317 51813 53337 51833 sw
tri 53337 51813 53648 52124 ne
rect 53648 52008 57417 52124
tri 57417 52008 57702 52293 sw
tri 57702 52128 57867 52293 ne
rect 57867 52200 59491 52293
tri 59491 52200 59775 52484 sw
tri 59775 52200 60059 52484 ne
rect 60059 52400 61739 52484
tri 61739 52400 61839 52500 sw
tri 62027 52400 62127 52500 ne
rect 62127 52400 71000 52500
rect 60059 52200 61839 52400
tri 61839 52200 62039 52400 sw
rect 57867 52128 59775 52200
tri 59775 52128 59847 52200 sw
tri 60059 52128 60131 52200 ne
rect 60131 52128 71000 52200
rect 53648 51843 57702 52008
tri 57702 51843 57867 52008 sw
tri 57867 51843 58152 52128 ne
rect 58152 51916 59847 52128
tri 59847 51916 60059 52128 sw
tri 60131 51916 60343 52128 ne
rect 60343 51916 71000 52128
rect 58152 51843 60059 51916
rect 53648 51813 57867 51843
rect 49290 51607 53337 51813
rect 47310 51320 49003 51607
tri 49003 51320 49290 51607 sw
tri 49290 51320 49577 51607 ne
rect 49577 51511 53337 51607
tri 53337 51511 53639 51813 sw
tri 53648 51617 53844 51813 ne
rect 53844 51617 57867 51813
rect 49577 51320 53639 51511
rect 40509 51312 44745 51320
rect 36266 51015 40500 51024
tri 40500 51015 40509 51024 sw
tri 40509 51015 40806 51312 ne
rect 40806 51027 44745 51312
tri 44745 51027 45038 51320 sw
tri 45038 51306 45052 51320 ne
rect 45052 51306 47018 51320
tri 47018 51306 47032 51320 sw
tri 47310 51306 47324 51320 ne
rect 47324 51306 49290 51320
rect 40806 51015 45038 51027
rect 36266 51014 40509 51015
rect 32097 50726 36199 50793
tri 36199 50726 36266 50793 sw
tri 36266 50791 36489 51014 ne
rect 36489 50791 40509 51014
rect 32097 50651 36266 50726
rect 27850 50360 31822 50632
rect 25678 50263 27560 50360
tri 27560 50263 27657 50360 sw
tri 27850 50263 27947 50360 ne
rect 27947 50357 31822 50360
tri 31822 50357 32097 50632 sw
tri 32097 50360 32388 50651 ne
rect 32388 50503 36266 50651
tri 36266 50503 36489 50726 sw
tri 36489 50649 36631 50791 ne
rect 36631 50718 40509 50791
tri 40509 50718 40806 51015 sw
tri 40806 50949 40872 51015 ne
rect 40872 51013 45038 51015
tri 45038 51013 45052 51027 sw
tri 45052 51014 45344 51306 ne
rect 45344 51014 47032 51306
tri 47032 51014 47324 51306 sw
tri 47324 51014 47616 51306 ne
rect 47616 51302 49290 51306
tri 49290 51302 49308 51320 sw
tri 49577 51302 49595 51320 ne
rect 49595 51306 53639 51320
tri 53639 51306 53844 51511 sw
tri 53844 51320 54141 51617 ne
rect 54141 51558 57867 51617
tri 57867 51558 58152 51843 sw
tri 58152 51607 58388 51843 ne
rect 58388 51632 60059 51843
tri 60059 51632 60343 51916 sw
tri 60343 51632 60627 51916 ne
rect 60627 51632 71000 51916
rect 58388 51607 60343 51632
rect 54141 51322 58152 51558
tri 58152 51322 58388 51558 sw
tri 58388 51322 58673 51607 ne
rect 58673 51604 60343 51607
tri 60343 51604 60371 51632 sw
tri 60627 51604 60655 51632 ne
rect 60655 51604 71000 51632
rect 58673 51322 60371 51604
rect 54141 51320 58388 51322
rect 49595 51302 53844 51306
rect 47616 51019 49308 51302
tri 49308 51019 49591 51302 sw
tri 49595 51019 49878 51302 ne
rect 49878 51296 53844 51302
tri 53844 51296 53854 51306 sw
rect 49878 51286 53854 51296
tri 53854 51286 53864 51296 sw
rect 49878 51276 53864 51286
tri 53864 51276 53874 51286 sw
rect 49878 51266 53874 51276
tri 53874 51266 53884 51276 sw
rect 49878 51256 53884 51266
tri 53884 51256 53894 51266 sw
rect 49878 51246 53894 51256
tri 53894 51246 53904 51256 sw
rect 49878 51236 53904 51246
tri 53904 51236 53914 51246 sw
rect 49878 51226 53914 51236
tri 53914 51226 53924 51236 sw
rect 49878 51216 53924 51226
tri 53924 51216 53934 51226 sw
rect 49878 51206 53934 51216
tri 53934 51206 53944 51216 sw
rect 49878 51196 53944 51206
tri 53944 51196 53954 51206 sw
rect 49878 51186 53954 51196
tri 53954 51186 53964 51196 sw
rect 49878 51176 53964 51186
tri 53964 51176 53974 51186 sw
rect 49878 51166 53974 51176
tri 53974 51166 53984 51176 sw
rect 49878 51156 53984 51166
tri 53984 51156 53994 51166 sw
rect 49878 51154 53994 51156
tri 53994 51154 53996 51156 sw
rect 49878 51144 53996 51154
tri 53996 51144 54006 51154 sw
rect 49878 51134 54006 51144
tri 54006 51134 54016 51144 sw
rect 49878 51124 54016 51134
tri 54016 51124 54026 51134 sw
rect 49878 51114 54026 51124
tri 54026 51114 54036 51124 sw
rect 49878 51104 54036 51114
tri 54036 51104 54046 51114 sw
rect 49878 51094 54046 51104
tri 54046 51094 54056 51104 sw
rect 49878 51084 54056 51094
tri 54056 51084 54066 51094 sw
rect 49878 51074 54066 51084
tri 54066 51074 54076 51084 sw
rect 49878 51064 54076 51074
tri 54076 51064 54086 51074 sw
rect 49878 51054 54086 51064
tri 54086 51054 54096 51064 sw
rect 49878 51044 54096 51054
tri 54096 51044 54106 51054 sw
rect 49878 51034 54106 51044
tri 54106 51034 54116 51044 sw
rect 49878 51024 54116 51034
tri 54116 51024 54126 51034 sw
rect 49878 51019 54126 51024
rect 47616 51014 49591 51019
rect 40872 50949 45052 51013
rect 36631 50652 40806 50718
tri 40806 50652 40872 50718 sw
tri 40872 50652 41169 50949 ne
rect 41169 50721 45052 50949
tri 45052 50721 45344 51013 sw
tri 45344 50900 45458 51014 ne
rect 45458 50900 47324 51014
tri 47324 50900 47438 51014 sw
tri 47616 50900 47730 51014 ne
rect 47730 50900 49591 51014
tri 49591 50900 49710 51019 sw
tri 49878 50900 49997 51019 ne
rect 49997 51014 54126 51019
tri 54126 51014 54136 51024 sw
tri 54141 51014 54447 51320 ne
rect 54447 51038 58388 51320
tri 58388 51038 58672 51322 sw
tri 58673 51301 58694 51322 ne
rect 58694 51320 60371 51322
tri 60371 51320 60655 51604 sw
tri 60655 51320 60939 51604 ne
rect 60939 51320 71000 51604
rect 58694 51301 60655 51320
rect 54447 51016 58672 51038
tri 58672 51016 58694 51038 sw
tri 58694 51016 58979 51301 ne
rect 58979 51298 60655 51301
tri 60655 51298 60677 51320 sw
tri 60939 51298 60961 51320 ne
rect 60961 51298 71000 51320
rect 58979 51016 60677 51298
rect 54447 51014 58694 51016
rect 49997 50900 54136 51014
rect 41169 50652 45344 50721
rect 36631 50649 40872 50652
rect 32388 50361 36489 50503
tri 36489 50361 36631 50503 sw
tri 36631 50361 36919 50649 ne
rect 36919 50361 40872 50649
rect 32388 50360 36631 50361
rect 27947 50263 32097 50357
rect 25678 50262 27657 50263
rect 23600 50071 25389 50262
tri 23400 49973 23401 49974 sw
tri 23600 49973 23698 50071 ne
rect 23698 49973 25389 50071
tri 25389 49973 25678 50262 sw
tri 25678 49973 25967 50262 ne
rect 25967 49973 27657 50262
tri 27657 49973 27947 50263 sw
tri 27947 49973 28237 50263 ne
rect 28237 50066 32097 50263
tri 32097 50066 32388 50357 sw
tri 32388 50268 32480 50360 ne
rect 32480 50268 36631 50360
rect 28237 49974 32388 50066
tri 32388 49974 32480 50066 sw
tri 32480 49974 32774 50268 ne
rect 32774 50073 36631 50268
tri 36631 50073 36919 50361 sw
tri 36919 50176 37104 50361 ne
rect 37104 50355 40872 50361
tri 40872 50355 41169 50652 sw
tri 41169 50360 41461 50652 ne
rect 41461 50607 45344 50652
tri 45344 50607 45458 50721 sw
tri 45458 50651 45707 50900 ne
rect 45707 50651 47438 50900
tri 47438 50651 47687 50900 sw
tri 47730 50651 47979 50900 ne
rect 47979 50651 49710 50900
tri 49710 50651 49959 50900 sw
tri 49997 50651 50246 50900 ne
rect 50246 50711 54136 50900
tri 54136 50711 54439 51014 sw
tri 54447 50900 54561 51014 ne
rect 54561 50900 58694 51014
rect 50246 50651 54439 50711
rect 41461 50360 45458 50607
rect 37104 50176 41169 50355
rect 32774 49974 36919 50073
rect 28237 49973 32480 49974
rect 20400 49676 23401 49973
tri 23401 49676 23698 49973 sw
tri 23698 49773 23898 49973 ne
rect 23898 49773 25678 49973
rect 20400 49476 23698 49676
tri 23698 49476 23898 49676 sw
tri 23898 49476 24195 49773 ne
rect 24195 49684 25678 49773
tri 25678 49684 25967 49973 sw
tri 25967 49684 26256 49973 ne
rect 26256 49684 27947 49973
rect 24195 49629 25967 49684
tri 25967 49629 26022 49684 sw
tri 26256 49629 26311 49684 ne
rect 26311 49683 27947 49684
tri 27947 49683 28237 49973 sw
tri 28237 49683 28527 49973 ne
rect 28527 49683 32480 49973
rect 26311 49629 28237 49683
rect 24195 49476 26022 49629
rect 20400 49179 23898 49476
tri 23898 49179 24195 49476 sw
tri 24195 49452 24219 49476 ne
rect 24219 49452 26022 49476
rect 20400 49155 24195 49179
tri 24195 49155 24219 49179 sw
tri 24219 49155 24516 49452 ne
rect 24516 49340 26022 49452
tri 26022 49340 26311 49629 sw
tri 26311 49340 26600 49629 ne
rect 26600 49437 28237 49629
tri 28237 49437 28483 49683 sw
tri 28527 49437 28773 49683 ne
rect 28773 49680 32480 49683
tri 32480 49680 32774 49974 sw
tri 32774 49748 33000 49974 ne
rect 33000 49888 36919 49974
tri 36919 49888 37104 50073 sw
tri 37104 49888 37392 50176 ne
rect 37392 50063 41169 50176
tri 41169 50063 41461 50355 sw
tri 41461 50271 41550 50360 ne
rect 41550 50358 45458 50360
tri 45458 50358 45707 50607 sw
tri 45707 50360 45998 50651 ne
rect 45998 50520 47687 50651
tri 47687 50520 47818 50651 sw
tri 47979 50520 48110 50651 ne
rect 48110 50520 49959 50651
tri 49959 50520 50090 50651 sw
tri 50246 50520 50377 50651 ne
rect 50377 50591 54439 50651
tri 54439 50591 54559 50711 sw
tri 54561 50651 54810 50900 ne
rect 54810 50731 58694 50900
tri 58694 50731 58979 51016 sw
tri 58979 50900 59095 51016 ne
rect 59095 51014 60677 51016
tri 60677 51014 60961 51298 sw
tri 60961 51014 61245 51298 ne
rect 61245 51014 71000 51298
rect 59095 50900 60961 51014
tri 60961 50900 61075 51014 sw
tri 61245 50900 61359 51014 ne
rect 61359 50900 71000 51014
rect 54810 50651 58979 50731
rect 50377 50520 54559 50591
rect 45998 50360 47818 50520
tri 47818 50360 47978 50520 sw
tri 48110 50360 48270 50520 ne
rect 48270 50360 50090 50520
rect 41550 50271 45707 50358
tri 41550 50176 41645 50271 ne
rect 41645 50176 45707 50271
rect 37392 49888 41461 50063
rect 33000 49748 37104 49888
rect 28773 49454 32774 49680
tri 32774 49454 33000 49680 sw
tri 33000 49454 33294 49748 ne
rect 33294 49600 37104 49748
tri 37104 49600 37392 49888 sw
tri 37392 49682 37598 49888 ne
rect 37598 49879 41461 49888
tri 41461 49879 41645 50063 sw
tri 41645 49971 41850 50176 ne
rect 41850 50067 45707 50176
tri 45707 50067 45998 50358 sw
tri 45998 50267 46091 50360 ne
rect 46091 50267 47978 50360
rect 41850 49974 45998 50067
tri 45998 49974 46091 50067 sw
tri 46091 49974 46384 50267 ne
rect 46384 50228 47978 50267
tri 47978 50228 48110 50360 sw
tri 48270 50228 48402 50360 ne
rect 48402 50330 50090 50360
tri 50090 50330 50280 50520 sw
tri 50377 50330 50567 50520 ne
rect 50567 50340 54559 50520
tri 54559 50340 54810 50591 sw
tri 54810 50360 55101 50651 ne
rect 55101 50616 58979 50651
tri 58979 50616 59094 50731 sw
tri 59095 50651 59344 50900 ne
rect 59344 50800 61075 50900
tri 61075 50800 61175 50900 sw
tri 61359 50800 61459 50900 ne
rect 61459 50800 71000 50900
rect 59344 50651 61175 50800
tri 61175 50651 61324 50800 sw
rect 55101 50366 59094 50616
tri 59094 50366 59344 50616 sw
tri 59344 50520 59475 50651 ne
rect 59475 50600 61324 50651
tri 61324 50600 61375 50651 sw
rect 59475 50520 71000 50600
rect 55101 50360 59344 50366
rect 50567 50330 54810 50340
rect 48402 50228 50280 50330
rect 46384 50043 48110 50228
tri 48110 50043 48295 50228 sw
tri 48402 50043 48587 50228 ne
rect 48587 50043 50280 50228
tri 50280 50043 50567 50330 sw
tri 50567 50043 50854 50330 ne
rect 50854 50049 54810 50330
tri 54810 50049 55101 50340 sw
tri 55101 50049 55412 50360 ne
rect 55412 50235 59344 50360
tri 59344 50235 59475 50366 sw
tri 59475 50360 59635 50520 ne
rect 59635 50360 71000 50520
tri 59635 50313 59682 50360 ne
rect 59682 50313 71000 50360
rect 55412 50233 59475 50235
tri 59475 50233 59477 50235 sw
rect 55412 50231 59477 50233
tri 59477 50231 59479 50233 sw
rect 55412 50229 59479 50231
tri 59479 50229 59481 50231 sw
rect 55412 50227 59481 50229
tri 59481 50227 59483 50229 sw
rect 55412 50225 59483 50227
tri 59483 50225 59485 50227 sw
rect 55412 50223 59485 50225
tri 59485 50223 59487 50225 sw
rect 55412 50221 59487 50223
tri 59487 50221 59489 50223 sw
rect 55412 50219 59489 50221
tri 59489 50219 59491 50221 sw
rect 55412 50217 59491 50219
tri 59491 50217 59493 50219 sw
rect 55412 50215 59493 50217
tri 59493 50215 59495 50217 sw
rect 55412 50213 59495 50215
tri 59495 50213 59497 50215 sw
rect 55412 50211 59497 50213
tri 59497 50211 59499 50213 sw
rect 55412 50209 59499 50211
tri 59499 50209 59501 50211 sw
rect 55412 50207 59501 50209
tri 59501 50207 59503 50209 sw
rect 55412 50205 59503 50207
tri 59503 50205 59505 50207 sw
rect 55412 50203 59505 50205
tri 59505 50203 59507 50205 sw
rect 55412 50201 59507 50203
tri 59507 50201 59509 50203 sw
rect 55412 50199 59509 50201
tri 59509 50199 59511 50201 sw
rect 55412 50197 59511 50199
tri 59511 50197 59513 50199 sw
rect 55412 50195 59513 50197
tri 59513 50195 59515 50197 sw
rect 55412 50193 59515 50195
tri 59515 50193 59517 50195 sw
rect 55412 50191 59517 50193
tri 59517 50191 59519 50193 sw
rect 55412 50189 59519 50191
tri 59519 50189 59521 50191 sw
rect 55412 50187 59521 50189
tri 59521 50187 59523 50189 sw
rect 55412 50185 59523 50187
tri 59523 50185 59525 50187 sw
rect 55412 50183 59525 50185
tri 59525 50183 59527 50185 sw
rect 55412 50181 59527 50183
tri 59527 50181 59529 50183 sw
rect 55412 50179 59529 50181
tri 59529 50179 59531 50181 sw
rect 55412 50177 59531 50179
tri 59531 50177 59533 50179 sw
rect 55412 50175 59533 50177
tri 59533 50175 59535 50177 sw
rect 55412 50173 59535 50175
tri 59535 50173 59537 50175 sw
rect 55412 50171 59537 50173
tri 59537 50171 59539 50173 sw
rect 55412 50169 59539 50171
tri 59539 50169 59541 50171 sw
rect 55412 50167 59541 50169
tri 59541 50167 59543 50169 sw
rect 55412 50165 59543 50167
tri 59543 50165 59545 50167 sw
rect 55412 50163 59545 50165
tri 59545 50163 59547 50165 sw
rect 55412 50161 59547 50163
tri 59547 50161 59549 50163 sw
rect 55412 50159 59549 50161
tri 59549 50159 59551 50161 sw
rect 55412 50157 59551 50159
tri 59551 50157 59553 50159 sw
rect 55412 50155 59553 50157
tri 59553 50155 59555 50157 sw
rect 55412 50153 59555 50155
tri 59555 50153 59557 50155 sw
rect 55412 50151 59557 50153
tri 59557 50151 59559 50153 sw
rect 55412 50149 59559 50151
tri 59559 50149 59561 50151 sw
rect 55412 50147 59561 50149
tri 59561 50147 59563 50149 sw
rect 55412 50145 59563 50147
tri 59563 50145 59565 50147 sw
rect 55412 50143 59565 50145
tri 59565 50143 59567 50145 sw
rect 55412 50141 59567 50143
tri 59567 50141 59569 50143 sw
rect 55412 50139 59569 50141
tri 59569 50139 59571 50141 sw
rect 55412 50137 59571 50139
tri 59571 50137 59573 50139 sw
rect 55412 50135 59573 50137
tri 59573 50135 59575 50137 sw
rect 55412 50133 59575 50135
tri 59575 50133 59577 50135 sw
rect 55412 50131 59577 50133
tri 59577 50131 59579 50133 sw
rect 55412 50129 59579 50131
tri 59579 50129 59581 50131 sw
rect 55412 50127 59581 50129
tri 59581 50127 59583 50129 sw
rect 55412 50125 59583 50127
tri 59583 50125 59585 50127 sw
rect 55412 50123 59585 50125
tri 59585 50123 59587 50125 sw
rect 55412 50121 59587 50123
tri 59587 50121 59589 50123 sw
rect 55412 50119 59589 50121
tri 59589 50119 59591 50121 sw
rect 55412 50117 59591 50119
tri 59591 50117 59593 50119 sw
rect 55412 50115 59593 50117
tri 59593 50115 59595 50117 sw
rect 55412 50113 59595 50115
tri 59595 50113 59597 50115 sw
rect 55412 50111 59597 50113
tri 59597 50111 59599 50113 sw
rect 55412 50110 59599 50111
tri 59599 50110 59600 50111 sw
rect 55412 50109 59600 50110
tri 59600 50109 59601 50110 sw
rect 55412 50108 59601 50109
tri 59601 50108 59602 50109 sw
rect 55412 50107 59602 50108
tri 59602 50107 59603 50108 sw
rect 55412 50106 59603 50107
tri 59603 50106 59604 50107 sw
rect 55412 50105 59604 50106
tri 59604 50105 59605 50106 sw
rect 55412 50104 59605 50105
tri 59605 50104 59606 50105 sw
rect 55412 50103 59606 50104
tri 59606 50103 59607 50104 sw
rect 55412 50102 59607 50103
tri 59607 50102 59608 50103 sw
rect 55412 50101 59608 50102
tri 59608 50101 59609 50102 sw
rect 55412 50100 59609 50101
tri 59609 50100 59610 50101 sw
rect 55412 50099 59610 50100
tri 59610 50099 59611 50100 sw
rect 55412 50098 59611 50099
tri 59611 50098 59612 50099 sw
rect 55412 50097 59612 50098
tri 59612 50097 59613 50098 sw
rect 55412 50096 59613 50097
tri 59613 50096 59614 50097 sw
rect 55412 50095 59614 50096
tri 59614 50095 59615 50096 sw
rect 55412 50094 59615 50095
tri 59615 50094 59616 50095 sw
rect 55412 50093 59616 50094
tri 59616 50093 59617 50094 sw
rect 55412 50092 59617 50093
tri 59617 50092 59618 50093 sw
rect 55412 50091 59618 50092
tri 59618 50091 59619 50092 sw
rect 55412 50090 59619 50091
tri 59619 50090 59620 50091 sw
rect 55412 50089 59620 50090
tri 59620 50089 59621 50090 sw
rect 55412 50088 59621 50089
tri 59621 50088 59622 50089 sw
rect 55412 50087 59622 50088
tri 59622 50087 59623 50088 sw
rect 55412 50086 59623 50087
tri 59623 50086 59624 50087 sw
rect 55412 50085 59624 50086
tri 59624 50085 59625 50086 sw
rect 55412 50084 59625 50085
tri 59625 50084 59626 50085 sw
rect 55412 50083 59626 50084
tri 59626 50083 59627 50084 sw
rect 55412 50082 59627 50083
tri 59627 50082 59628 50083 sw
rect 55412 50081 59628 50082
tri 59628 50081 59629 50082 sw
rect 55412 50080 59629 50081
tri 59629 50080 59630 50081 sw
rect 55412 50079 59630 50080
tri 59630 50079 59631 50080 sw
rect 55412 50078 59631 50079
tri 59631 50078 59632 50079 sw
rect 55412 50077 59632 50078
tri 59632 50077 59633 50078 sw
rect 55412 50076 59633 50077
tri 59633 50076 59634 50077 sw
rect 55412 50075 59634 50076
tri 59634 50075 59635 50076 sw
rect 55412 50074 59635 50075
tri 59635 50074 59636 50075 sw
rect 55412 50073 59636 50074
tri 59636 50073 59637 50074 sw
rect 55412 50072 59637 50073
tri 59637 50072 59638 50073 sw
rect 55412 50071 59638 50072
tri 59638 50071 59639 50072 sw
rect 55412 50070 59639 50071
tri 59639 50070 59640 50071 sw
rect 55412 50069 59640 50070
tri 59640 50069 59641 50070 sw
rect 55412 50068 59641 50069
tri 59641 50068 59642 50069 sw
rect 55412 50067 59642 50068
tri 59642 50067 59643 50068 sw
rect 55412 50066 59643 50067
tri 59643 50066 59644 50067 sw
rect 55412 50065 59644 50066
tri 59644 50065 59645 50066 sw
rect 55412 50064 59645 50065
tri 59645 50064 59646 50065 sw
rect 55412 50063 59646 50064
tri 59646 50063 59647 50064 sw
rect 55412 50062 59647 50063
tri 59647 50062 59648 50063 sw
rect 55412 50061 59648 50062
tri 59648 50061 59649 50062 sw
rect 55412 50060 59649 50061
tri 59649 50060 59650 50061 sw
rect 55412 50059 59650 50060
tri 59650 50059 59651 50060 sw
rect 55412 50058 59651 50059
tri 59651 50058 59652 50059 sw
rect 55412 50057 59652 50058
tri 59652 50057 59653 50058 sw
rect 55412 50056 59653 50057
tri 59653 50056 59654 50057 sw
rect 55412 50055 59654 50056
tri 59654 50055 59655 50056 sw
rect 55412 50054 59655 50055
tri 59655 50054 59656 50055 sw
rect 55412 50053 59656 50054
tri 59656 50053 59657 50054 sw
rect 55412 50052 59657 50053
tri 59657 50052 59658 50053 sw
rect 55412 50051 59658 50052
tri 59658 50051 59659 50052 sw
rect 55412 50050 59659 50051
tri 59659 50050 59660 50051 sw
rect 55412 50049 59660 50050
tri 59660 50049 59661 50050 sw
rect 50854 50043 55101 50049
rect 46384 49974 48295 50043
rect 41850 49971 46091 49974
rect 37598 49682 41645 49879
rect 33294 49506 37392 49600
tri 37392 49506 37486 49600 sw
tri 37598 49506 37774 49682 ne
rect 37774 49674 41645 49682
tri 41645 49674 41850 49879 sw
tri 41850 49674 42147 49971 ne
rect 42147 49681 46091 49971
tri 46091 49681 46384 49974 sw
tri 46384 49971 46387 49974 ne
rect 46387 49973 48295 49974
tri 48295 49973 48365 50043 sw
tri 48587 49973 48657 50043 ne
rect 48657 49973 50567 50043
rect 46387 49971 48365 49973
tri 48365 49971 48367 49973 sw
tri 48657 49971 48659 49973 ne
rect 48659 49971 50567 49973
tri 50567 49971 50639 50043 sw
tri 50854 49971 50926 50043 ne
rect 50926 49971 55101 50043
rect 42147 49678 46384 49681
tri 46384 49678 46387 49681 sw
tri 46387 49678 46680 49971 ne
rect 46680 49679 48367 49971
tri 48367 49679 48659 49971 sw
tri 48659 49679 48951 49971 ne
rect 48951 49755 50639 49971
tri 50639 49755 50855 49971 sw
tri 50926 49755 51142 49971 ne
rect 51142 49755 55101 49971
rect 48951 49679 50855 49755
rect 46680 49678 48659 49679
rect 42147 49674 46387 49678
rect 37774 49524 41850 49674
tri 41850 49524 42000 49674 sw
tri 42147 49524 42297 49674 ne
rect 42297 49524 46387 49674
rect 37774 49506 42000 49524
rect 33294 49454 37486 49506
rect 28773 49437 33000 49454
rect 26600 49340 28483 49437
rect 24516 49155 26311 49340
rect 20400 48858 24219 49155
tri 24219 48858 24516 49155 sw
tri 24516 49027 24644 49155 ne
rect 24644 49051 26311 49155
tri 26311 49051 26600 49340 sw
tri 26600 49051 26889 49340 ne
rect 26889 49147 28483 49340
tri 28483 49147 28773 49437 sw
tri 28773 49147 29063 49437 ne
rect 29063 49160 33000 49437
tri 33000 49160 33294 49454 sw
tri 33294 49453 33295 49454 ne
rect 33295 49453 37486 49454
rect 29063 49159 33294 49160
tri 33294 49159 33295 49160 sw
tri 33295 49159 33589 49453 ne
rect 33589 49218 37486 49453
tri 37486 49218 37774 49506 sw
tri 37774 49218 38062 49506 ne
rect 38062 49227 42000 49506
tri 42000 49227 42297 49524 sw
tri 42297 49227 42594 49524 ne
rect 42594 49385 46387 49524
tri 46387 49385 46680 49678 sw
tri 46680 49425 46933 49678 ne
rect 46933 49512 48659 49678
tri 48659 49512 48826 49679 sw
tri 48951 49512 49118 49679 ne
rect 49118 49512 50855 49679
rect 46933 49425 48826 49512
rect 42594 49227 46680 49385
rect 38062 49218 42297 49227
rect 33589 49159 37774 49218
rect 29063 49147 33295 49159
rect 26889 49051 28773 49147
rect 24644 49027 26600 49051
rect 20400 48730 24516 48858
tri 24516 48730 24644 48858 sw
tri 24644 48760 24911 49027 ne
rect 24911 48857 26600 49027
tri 26600 48857 26794 49051 sw
rect 24911 48851 26794 48857
tri 26794 48851 26800 48857 sw
tri 26889 48851 27089 49051 ne
rect 27089 48857 28773 49051
tri 28773 48857 29063 49147 sw
tri 29063 48857 29353 49147 ne
rect 29353 48865 33295 49147
tri 33295 48865 33589 49159 sw
tri 33589 49151 33597 49159 ne
rect 33597 49151 37774 49159
rect 29353 48857 33589 48865
tri 33589 48857 33597 48865 sw
tri 33597 48857 33891 49151 ne
rect 33891 48930 37774 49151
tri 37774 48930 38062 49218 sw
tri 38062 49217 38063 49218 ne
rect 38063 49217 42297 49218
rect 33891 48929 38062 48930
tri 38062 48929 38063 48930 sw
tri 38063 48929 38351 49217 ne
rect 38351 48930 42297 49217
tri 42297 48930 42594 49227 sw
tri 42594 49132 42689 49227 ne
rect 42689 49132 46680 49227
tri 46680 49132 46933 49385 sw
tri 46933 49222 47136 49425 ne
rect 47136 49222 48826 49425
tri 47136 49132 47226 49222 ne
rect 47226 49220 48826 49222
tri 48826 49220 49118 49512 sw
tri 49118 49220 49410 49512 ne
rect 49410 49468 50855 49512
tri 50855 49468 51142 49755 sw
tri 51142 49468 51429 49755 ne
rect 51429 49746 55101 49755
tri 55101 49746 55404 50049 sw
tri 55412 49928 55533 50049 ne
rect 55533 50048 59661 50049
tri 59661 50048 59662 50049 sw
rect 55533 50047 59662 50048
tri 59662 50047 59663 50048 sw
rect 55533 50046 59663 50047
tri 59663 50046 59664 50047 sw
rect 55533 50045 59664 50046
tri 59664 50045 59665 50046 sw
rect 55533 50044 59665 50045
tri 59665 50044 59666 50045 sw
rect 55533 50043 59666 50044
tri 59666 50043 59667 50044 sw
tri 59682 50043 59952 50313 ne
rect 59952 50043 71000 50313
rect 55533 49928 59667 50043
rect 51429 49626 55404 49746
tri 55404 49626 55524 49746 sw
tri 55533 49646 55815 49928 ne
rect 55815 49758 59667 49928
tri 59667 49758 59952 50043 sw
tri 59952 49971 60024 50043 ne
rect 60024 49971 71000 50043
rect 55815 49686 59952 49758
tri 59952 49686 60024 49758 sw
tri 60024 49686 60309 49971 ne
rect 60309 49686 71000 49971
rect 55815 49646 60024 49686
rect 51429 49468 55524 49626
rect 49410 49220 51142 49468
rect 47226 49132 49118 49220
rect 38351 48929 42594 48930
rect 33891 48857 38063 48929
rect 27089 48851 29063 48857
rect 24911 48760 26800 48851
tri 20400 48648 20482 48730 ne
rect 20482 48729 24644 48730
tri 24644 48729 24645 48730 sw
rect 20482 48728 24645 48729
tri 24645 48728 24646 48729 sw
rect 20482 48727 24646 48728
tri 24646 48727 24647 48728 sw
rect 20482 48726 24647 48727
tri 24647 48726 24648 48727 sw
rect 20482 48725 24648 48726
tri 24648 48725 24649 48726 sw
rect 20482 48724 24649 48725
tri 24649 48724 24650 48725 sw
rect 20482 48723 24650 48724
tri 24650 48723 24651 48724 sw
rect 20482 48722 24651 48723
tri 24651 48722 24652 48723 sw
rect 20482 48721 24652 48722
tri 24652 48721 24653 48722 sw
rect 20482 48720 24653 48721
tri 24653 48720 24654 48721 sw
rect 20482 48719 24654 48720
tri 24654 48719 24655 48720 sw
rect 20482 48718 24655 48719
tri 24655 48718 24656 48719 sw
rect 20482 48717 24656 48718
tri 24656 48717 24657 48718 sw
rect 20482 48716 24657 48717
tri 24657 48716 24658 48717 sw
rect 20482 48715 24658 48716
tri 24658 48715 24659 48716 sw
rect 20482 48714 24659 48715
tri 24659 48714 24660 48715 sw
rect 20482 48713 24660 48714
tri 24660 48713 24661 48714 sw
rect 20482 48712 24661 48713
tri 24661 48712 24662 48713 sw
rect 20482 48711 24662 48712
tri 24662 48711 24663 48712 sw
rect 20482 48710 24663 48711
tri 24663 48710 24664 48711 sw
rect 20482 48709 24664 48710
tri 24664 48709 24665 48710 sw
rect 20482 48708 24665 48709
tri 24665 48708 24666 48709 sw
rect 20482 48707 24666 48708
tri 24666 48707 24667 48708 sw
rect 20482 48706 24667 48707
tri 24667 48706 24668 48707 sw
rect 20482 48705 24668 48706
tri 24668 48705 24669 48706 sw
rect 20482 48704 24669 48705
tri 24669 48704 24670 48705 sw
rect 20482 48703 24670 48704
tri 24670 48703 24671 48704 sw
rect 20482 48702 24671 48703
tri 24671 48702 24672 48703 sw
rect 20482 48701 24672 48702
tri 24672 48701 24673 48702 sw
rect 20482 48700 24673 48701
tri 24673 48700 24674 48701 sw
rect 20482 48699 24674 48700
tri 24674 48699 24675 48700 sw
rect 20482 48698 24675 48699
tri 24675 48698 24676 48699 sw
rect 20482 48697 24676 48698
tri 24676 48697 24677 48698 sw
rect 20482 48696 24677 48697
tri 24677 48696 24678 48697 sw
rect 20482 48695 24678 48696
tri 24678 48695 24679 48696 sw
rect 20482 48694 24679 48695
tri 24679 48694 24680 48695 sw
rect 20482 48693 24680 48694
tri 24680 48693 24681 48694 sw
rect 20482 48692 24681 48693
tri 24681 48692 24682 48693 sw
rect 20482 48691 24682 48692
tri 24682 48691 24683 48692 sw
rect 20482 48690 24683 48691
tri 24683 48690 24684 48691 sw
rect 20482 48689 24684 48690
tri 24684 48689 24685 48690 sw
rect 20482 48688 24685 48689
tri 24685 48688 24686 48689 sw
rect 20482 48687 24686 48688
tri 24686 48687 24687 48688 sw
rect 20482 48686 24687 48687
tri 24687 48686 24688 48687 sw
rect 20482 48685 24688 48686
tri 24688 48685 24689 48686 sw
rect 20482 48684 24689 48685
tri 24689 48684 24690 48685 sw
rect 20482 48683 24690 48684
tri 24690 48683 24691 48684 sw
rect 20482 48682 24691 48683
tri 24691 48682 24692 48683 sw
rect 20482 48681 24692 48682
tri 24692 48681 24693 48682 sw
rect 20482 48680 24693 48681
tri 24693 48680 24694 48681 sw
rect 20482 48679 24694 48680
tri 24694 48679 24695 48680 sw
rect 20482 48678 24695 48679
tri 24695 48678 24696 48679 sw
rect 20482 48677 24696 48678
tri 24696 48677 24697 48678 sw
rect 20482 48676 24697 48677
tri 24697 48676 24698 48677 sw
rect 20482 48675 24698 48676
tri 24698 48675 24699 48676 sw
rect 20482 48674 24699 48675
tri 24699 48674 24700 48675 sw
rect 20482 48673 24700 48674
tri 24700 48673 24701 48674 sw
rect 20482 48672 24701 48673
tri 24701 48672 24702 48673 sw
rect 20482 48671 24702 48672
tri 24702 48671 24703 48672 sw
rect 20482 48670 24703 48671
tri 24703 48670 24704 48671 sw
rect 20482 48669 24704 48670
tri 24704 48669 24705 48670 sw
rect 20482 48668 24705 48669
tri 24705 48668 24706 48669 sw
rect 20482 48667 24706 48668
tri 24706 48667 24707 48668 sw
rect 20482 48666 24707 48667
tri 24707 48666 24708 48667 sw
rect 20482 48665 24708 48666
tri 24708 48665 24709 48666 sw
rect 20482 48664 24709 48665
tri 24709 48664 24710 48665 sw
rect 20482 48663 24710 48664
tri 24710 48663 24711 48664 sw
rect 20482 48662 24711 48663
tri 24711 48662 24712 48663 sw
rect 20482 48661 24712 48662
tri 24712 48661 24713 48662 sw
rect 20482 48660 24713 48661
tri 24713 48660 24714 48661 sw
rect 20482 48659 24714 48660
tri 24714 48659 24715 48660 sw
rect 20482 48658 24715 48659
tri 24715 48658 24716 48659 sw
rect 20482 48657 24716 48658
tri 24716 48657 24717 48658 sw
rect 20482 48656 24717 48657
tri 24717 48656 24718 48657 sw
rect 20482 48655 24718 48656
tri 24718 48655 24719 48656 sw
rect 20482 48654 24719 48655
tri 24719 48654 24720 48655 sw
rect 20482 48653 24720 48654
tri 24720 48653 24721 48654 sw
rect 20482 48652 24721 48653
tri 24721 48652 24722 48653 sw
rect 20482 48651 24722 48652
tri 24722 48651 24723 48652 sw
rect 20482 48650 24723 48651
tri 24723 48650 24724 48651 sw
rect 20482 48649 24724 48650
tri 24724 48649 24725 48650 sw
rect 20482 48648 24725 48649
tri 24725 48648 24726 48649 sw
tri 20200 48366 20482 48648 sw
tri 20482 48447 20683 48648 ne
rect 20683 48647 24726 48648
tri 24726 48647 24727 48648 sw
tri 24911 48647 25024 48760 ne
rect 25024 48647 26800 48760
tri 26800 48647 27004 48851 sw
tri 27089 48647 27293 48851 ne
rect 27293 48647 29063 48851
tri 29063 48647 29273 48857 sw
tri 29353 48647 29563 48857 ne
rect 29563 48647 33597 48857
rect 20683 48447 24727 48647
rect 17200 48165 20482 48366
tri 20482 48165 20683 48366 sw
tri 20683 48165 20965 48447 ne
rect 20965 48350 24727 48447
tri 24727 48350 25024 48647 sw
tri 25024 48373 25298 48647 ne
rect 25298 48380 27004 48647
tri 27004 48380 27271 48647 sw
tri 27293 48380 27560 48647 ne
rect 27560 48380 29273 48647
tri 29273 48380 29540 48647 sw
tri 29563 48380 29830 48647 ne
rect 29830 48563 33597 48647
tri 33597 48563 33891 48857 sw
tri 33891 48647 34101 48857 ne
rect 34101 48647 38063 48857
rect 29830 48380 33891 48563
rect 25298 48373 27271 48380
rect 20965 48165 25024 48350
rect 17200 47883 20683 48165
tri 20683 47883 20965 48165 sw
tri 20965 48164 20966 48165 ne
rect 20966 48164 25024 48165
rect 17200 47882 20965 47883
tri 20965 47882 20966 47883 sw
tri 20966 47882 21248 48164 ne
rect 21248 48076 25024 48164
tri 25024 48076 25298 48350 sw
tri 25298 48076 25595 48373 ne
rect 25595 48091 27271 48373
tri 27271 48091 27560 48380 sw
tri 27560 48091 27849 48380 ne
rect 27849 48120 29540 48380
tri 29540 48120 29800 48380 sw
tri 29830 48120 30090 48380 ne
rect 30090 48353 33891 48380
tri 33891 48353 34101 48563 sw
tri 34101 48379 34369 48647 ne
rect 34369 48641 38063 48647
tri 38063 48641 38351 48929 sw
tri 38351 48928 38352 48929 ne
rect 38352 48928 42594 48929
rect 34369 48640 38351 48641
tri 38351 48640 38352 48641 sw
tri 38352 48640 38640 48928 ne
rect 38640 48835 42594 48928
tri 42594 48835 42689 48930 sw
tri 42689 48835 42986 49132 ne
rect 42986 49131 46933 49132
tri 46933 49131 46934 49132 sw
rect 42986 49130 46934 49131
tri 46934 49130 46935 49131 sw
rect 42986 49129 46935 49130
tri 46935 49129 46936 49130 sw
rect 42986 49128 46936 49129
tri 46936 49128 46937 49129 sw
rect 42986 49127 46937 49128
tri 46937 49127 46938 49128 sw
rect 42986 49126 46938 49127
tri 46938 49126 46939 49127 sw
rect 42986 49125 46939 49126
tri 46939 49125 46940 49126 sw
rect 42986 49124 46940 49125
tri 46940 49124 46941 49125 sw
rect 42986 49123 46941 49124
tri 46941 49123 46942 49124 sw
rect 42986 49122 46942 49123
tri 46942 49122 46943 49123 sw
rect 42986 49121 46943 49122
tri 46943 49121 46944 49122 sw
rect 42986 49120 46944 49121
tri 46944 49120 46945 49121 sw
rect 42986 49119 46945 49120
tri 46945 49119 46946 49120 sw
rect 42986 49118 46946 49119
tri 46946 49118 46947 49119 sw
rect 42986 49117 46947 49118
tri 46947 49117 46948 49118 sw
rect 42986 49116 46948 49117
tri 46948 49116 46949 49117 sw
rect 42986 49115 46949 49116
tri 46949 49115 46950 49116 sw
rect 42986 49114 46950 49115
tri 46950 49114 46951 49115 sw
rect 42986 49113 46951 49114
tri 46951 49113 46952 49114 sw
rect 42986 49112 46952 49113
tri 46952 49112 46953 49113 sw
rect 42986 49111 46953 49112
tri 46953 49111 46954 49112 sw
rect 42986 49110 46954 49111
tri 46954 49110 46955 49111 sw
rect 42986 49109 46955 49110
tri 46955 49109 46956 49110 sw
rect 42986 49108 46956 49109
tri 46956 49108 46957 49109 sw
rect 42986 49107 46957 49108
tri 46957 49107 46958 49108 sw
rect 42986 49106 46958 49107
tri 46958 49106 46959 49107 sw
rect 42986 49105 46959 49106
tri 46959 49105 46960 49106 sw
rect 42986 49104 46960 49105
tri 46960 49104 46961 49105 sw
rect 42986 49103 46961 49104
tri 46961 49103 46962 49104 sw
rect 42986 49102 46962 49103
tri 46962 49102 46963 49103 sw
rect 42986 49101 46963 49102
tri 46963 49101 46964 49102 sw
rect 42986 49100 46964 49101
tri 46964 49100 46965 49101 sw
rect 42986 49099 46965 49100
tri 46965 49099 46966 49100 sw
rect 42986 49098 46966 49099
tri 46966 49098 46967 49099 sw
rect 42986 49097 46967 49098
tri 46967 49097 46968 49098 sw
rect 42986 49096 46968 49097
tri 46968 49096 46969 49097 sw
rect 42986 49095 46969 49096
tri 46969 49095 46970 49096 sw
rect 42986 49094 46970 49095
tri 46970 49094 46971 49095 sw
rect 42986 49093 46971 49094
tri 46971 49093 46972 49094 sw
rect 42986 49092 46972 49093
tri 46972 49092 46973 49093 sw
rect 42986 49091 46973 49092
tri 46973 49091 46974 49092 sw
rect 42986 49090 46974 49091
tri 46974 49090 46975 49091 sw
rect 42986 49089 46975 49090
tri 46975 49089 46976 49090 sw
rect 42986 49088 46976 49089
tri 46976 49088 46977 49089 sw
rect 42986 49087 46977 49088
tri 46977 49087 46978 49088 sw
rect 42986 49086 46978 49087
tri 46978 49086 46979 49087 sw
rect 42986 49085 46979 49086
tri 46979 49085 46980 49086 sw
rect 42986 49084 46980 49085
tri 46980 49084 46981 49085 sw
rect 42986 49083 46981 49084
tri 46981 49083 46982 49084 sw
rect 42986 49082 46982 49083
tri 46982 49082 46983 49083 sw
rect 42986 49081 46983 49082
tri 46983 49081 46984 49082 sw
rect 42986 49080 46984 49081
tri 46984 49080 46985 49081 sw
rect 42986 49079 46985 49080
tri 46985 49079 46986 49080 sw
rect 42986 49078 46986 49079
tri 46986 49078 46987 49079 sw
rect 42986 49077 46987 49078
tri 46987 49077 46988 49078 sw
rect 42986 49076 46988 49077
tri 46988 49076 46989 49077 sw
rect 42986 49075 46989 49076
tri 46989 49075 46990 49076 sw
rect 42986 49074 46990 49075
tri 46990 49074 46991 49075 sw
rect 42986 49073 46991 49074
tri 46991 49073 46992 49074 sw
rect 42986 49072 46992 49073
tri 46992 49072 46993 49073 sw
rect 42986 49071 46993 49072
tri 46993 49071 46994 49072 sw
rect 42986 49070 46994 49071
tri 46994 49070 46995 49071 sw
rect 42986 49069 46995 49070
tri 46995 49069 46996 49070 sw
rect 42986 49068 46996 49069
tri 46996 49068 46997 49069 sw
rect 42986 49067 46997 49068
tri 46997 49067 46998 49068 sw
rect 42986 49066 46998 49067
tri 46998 49066 46999 49067 sw
rect 42986 49065 46999 49066
tri 46999 49065 47000 49066 sw
rect 42986 49064 47000 49065
tri 47000 49064 47001 49065 sw
rect 42986 49063 47001 49064
tri 47001 49063 47002 49064 sw
rect 42986 49062 47002 49063
tri 47002 49062 47003 49063 sw
rect 42986 49061 47003 49062
tri 47003 49061 47004 49062 sw
rect 42986 49060 47004 49061
tri 47004 49060 47005 49061 sw
rect 42986 49059 47005 49060
tri 47005 49059 47006 49060 sw
rect 42986 49058 47006 49059
tri 47006 49058 47007 49059 sw
rect 42986 49057 47007 49058
tri 47007 49057 47008 49058 sw
rect 42986 49056 47008 49057
tri 47008 49056 47009 49057 sw
rect 42986 49055 47009 49056
tri 47009 49055 47010 49056 sw
rect 42986 49054 47010 49055
tri 47010 49054 47011 49055 sw
rect 42986 49053 47011 49054
tri 47011 49053 47012 49054 sw
rect 42986 49052 47012 49053
tri 47012 49052 47013 49053 sw
rect 42986 49051 47013 49052
tri 47013 49051 47014 49052 sw
rect 42986 49050 47014 49051
tri 47014 49050 47015 49051 sw
rect 42986 49049 47015 49050
tri 47015 49049 47016 49050 sw
rect 42986 49048 47016 49049
tri 47016 49048 47017 49049 sw
rect 42986 49047 47017 49048
tri 47017 49047 47018 49048 sw
rect 42986 49046 47018 49047
tri 47018 49046 47019 49047 sw
rect 42986 49045 47019 49046
tri 47019 49045 47020 49046 sw
rect 42986 49044 47020 49045
tri 47020 49044 47021 49045 sw
rect 42986 49043 47021 49044
tri 47021 49043 47022 49044 sw
rect 42986 49042 47022 49043
tri 47022 49042 47023 49043 sw
rect 42986 49041 47023 49042
tri 47023 49041 47024 49042 sw
rect 42986 49040 47024 49041
tri 47024 49040 47025 49041 sw
rect 42986 49039 47025 49040
tri 47025 49039 47026 49040 sw
rect 42986 49038 47026 49039
tri 47026 49038 47027 49039 sw
rect 42986 49037 47027 49038
tri 47027 49037 47028 49038 sw
rect 42986 49036 47028 49037
tri 47028 49036 47029 49037 sw
rect 42986 49035 47029 49036
tri 47029 49035 47030 49036 sw
rect 42986 49034 47030 49035
tri 47030 49034 47031 49035 sw
rect 42986 49033 47031 49034
tri 47031 49033 47032 49034 sw
rect 42986 49032 47032 49033
tri 47032 49032 47033 49033 sw
rect 42986 49031 47033 49032
tri 47033 49031 47034 49032 sw
rect 42986 49030 47034 49031
tri 47034 49030 47035 49031 sw
rect 42986 49029 47035 49030
tri 47035 49029 47036 49030 sw
rect 42986 49028 47036 49029
tri 47036 49028 47037 49029 sw
rect 42986 49027 47037 49028
tri 47037 49027 47038 49028 sw
rect 42986 49026 47038 49027
tri 47038 49026 47039 49027 sw
rect 42986 49025 47039 49026
tri 47039 49025 47040 49026 sw
rect 42986 49024 47040 49025
tri 47040 49024 47041 49025 sw
rect 42986 49023 47041 49024
tri 47041 49023 47042 49024 sw
rect 42986 49022 47042 49023
tri 47042 49022 47043 49023 sw
rect 42986 49021 47043 49022
tri 47043 49021 47044 49022 sw
rect 42986 49020 47044 49021
tri 47044 49020 47045 49021 sw
rect 42986 49019 47045 49020
tri 47045 49019 47046 49020 sw
rect 42986 49018 47046 49019
tri 47046 49018 47047 49019 sw
rect 42986 49017 47047 49018
tri 47047 49017 47048 49018 sw
rect 42986 49016 47048 49017
tri 47048 49016 47049 49017 sw
rect 42986 49015 47049 49016
tri 47049 49015 47050 49016 sw
rect 42986 49014 47050 49015
tri 47050 49014 47051 49015 sw
rect 42986 49013 47051 49014
tri 47051 49013 47052 49014 sw
rect 42986 49012 47052 49013
tri 47052 49012 47053 49013 sw
rect 42986 49011 47053 49012
tri 47053 49011 47054 49012 sw
rect 42986 49010 47054 49011
tri 47054 49010 47055 49011 sw
rect 42986 49009 47055 49010
tri 47055 49009 47056 49010 sw
rect 42986 49008 47056 49009
tri 47056 49008 47057 49009 sw
rect 42986 49007 47057 49008
tri 47057 49007 47058 49008 sw
rect 42986 49006 47058 49007
tri 47058 49006 47059 49007 sw
rect 42986 49005 47059 49006
tri 47059 49005 47060 49006 sw
rect 42986 49004 47060 49005
tri 47060 49004 47061 49005 sw
rect 42986 49003 47061 49004
tri 47061 49003 47062 49004 sw
rect 42986 49002 47062 49003
tri 47062 49002 47063 49003 sw
rect 42986 49001 47063 49002
tri 47063 49001 47064 49002 sw
rect 42986 49000 47064 49001
tri 47064 49000 47065 49001 sw
rect 42986 48999 47065 49000
tri 47065 48999 47066 49000 sw
rect 42986 48998 47066 48999
tri 47066 48998 47067 48999 sw
rect 42986 48997 47067 48998
tri 47067 48997 47068 48998 sw
rect 42986 48996 47068 48997
tri 47068 48996 47069 48997 sw
rect 42986 48995 47069 48996
tri 47069 48995 47070 48996 sw
rect 42986 48994 47070 48995
tri 47070 48994 47071 48995 sw
rect 42986 48993 47071 48994
tri 47071 48993 47072 48994 sw
rect 42986 48992 47072 48993
tri 47072 48992 47073 48993 sw
rect 42986 48991 47073 48992
tri 47073 48991 47074 48992 sw
rect 42986 48990 47074 48991
tri 47074 48990 47075 48991 sw
rect 42986 48989 47075 48990
tri 47075 48989 47076 48990 sw
rect 42986 48988 47076 48989
tri 47076 48988 47077 48989 sw
rect 42986 48987 47077 48988
tri 47077 48987 47078 48988 sw
rect 42986 48986 47078 48987
tri 47078 48986 47079 48987 sw
rect 42986 48985 47079 48986
tri 47079 48985 47080 48986 sw
rect 42986 48984 47080 48985
tri 47080 48984 47081 48985 sw
rect 42986 48983 47081 48984
tri 47081 48983 47082 48984 sw
rect 42986 48982 47082 48983
tri 47082 48982 47083 48983 sw
rect 42986 48981 47083 48982
tri 47083 48981 47084 48982 sw
rect 42986 48980 47084 48981
tri 47084 48980 47085 48981 sw
rect 42986 48979 47085 48980
tri 47085 48979 47086 48980 sw
rect 42986 48978 47086 48979
tri 47086 48978 47087 48979 sw
rect 42986 48977 47087 48978
tri 47087 48977 47088 48978 sw
rect 42986 48976 47088 48977
tri 47088 48976 47089 48977 sw
rect 42986 48975 47089 48976
tri 47089 48975 47090 48976 sw
rect 42986 48974 47090 48975
tri 47090 48974 47091 48975 sw
rect 42986 48973 47091 48974
tri 47091 48973 47092 48974 sw
rect 42986 48972 47092 48973
tri 47092 48972 47093 48973 sw
rect 42986 48971 47093 48972
tri 47093 48971 47094 48972 sw
rect 42986 48970 47094 48971
tri 47094 48970 47095 48971 sw
rect 42986 48969 47095 48970
tri 47095 48969 47096 48970 sw
rect 42986 48968 47096 48969
tri 47096 48968 47097 48969 sw
rect 42986 48967 47097 48968
tri 47097 48967 47098 48968 sw
rect 42986 48966 47098 48967
tri 47098 48966 47099 48967 sw
rect 42986 48965 47099 48966
tri 47099 48965 47100 48966 sw
rect 42986 48964 47100 48965
tri 47100 48964 47101 48965 sw
rect 42986 48963 47101 48964
tri 47101 48963 47102 48964 sw
rect 42986 48962 47102 48963
tri 47102 48962 47103 48963 sw
rect 42986 48961 47103 48962
tri 47103 48961 47104 48962 sw
rect 42986 48960 47104 48961
tri 47104 48960 47105 48961 sw
rect 42986 48959 47105 48960
tri 47105 48959 47106 48960 sw
rect 42986 48958 47106 48959
tri 47106 48958 47107 48959 sw
rect 42986 48957 47107 48958
tri 47107 48957 47108 48958 sw
rect 42986 48956 47108 48957
tri 47108 48956 47109 48957 sw
rect 42986 48955 47109 48956
tri 47109 48955 47110 48956 sw
rect 42986 48954 47110 48955
tri 47110 48954 47111 48955 sw
rect 42986 48953 47111 48954
tri 47111 48953 47112 48954 sw
rect 42986 48952 47112 48953
tri 47112 48952 47113 48953 sw
rect 42986 48951 47113 48952
tri 47113 48951 47114 48952 sw
rect 42986 48950 47114 48951
tri 47114 48950 47115 48951 sw
rect 42986 48949 47115 48950
tri 47115 48949 47116 48950 sw
rect 42986 48948 47116 48949
tri 47116 48948 47117 48949 sw
rect 42986 48947 47117 48948
tri 47117 48947 47118 48948 sw
rect 42986 48946 47118 48947
tri 47118 48946 47119 48947 sw
rect 42986 48945 47119 48946
tri 47119 48945 47120 48946 sw
rect 42986 48944 47120 48945
tri 47120 48944 47121 48945 sw
rect 42986 48943 47121 48944
tri 47121 48943 47122 48944 sw
rect 42986 48942 47122 48943
tri 47122 48942 47123 48943 sw
rect 42986 48941 47123 48942
tri 47123 48941 47124 48942 sw
rect 42986 48940 47124 48941
tri 47124 48940 47125 48941 sw
rect 42986 48939 47125 48940
tri 47125 48939 47126 48940 sw
rect 42986 48938 47126 48939
tri 47126 48938 47127 48939 sw
rect 42986 48937 47127 48938
tri 47127 48937 47128 48938 sw
rect 42986 48936 47128 48937
tri 47128 48936 47129 48937 sw
rect 42986 48935 47129 48936
tri 47129 48935 47130 48936 sw
rect 42986 48934 47130 48935
tri 47130 48934 47131 48935 sw
rect 42986 48933 47131 48934
tri 47131 48933 47132 48934 sw
rect 42986 48932 47132 48933
tri 47132 48932 47133 48933 sw
rect 42986 48931 47133 48932
tri 47133 48931 47134 48932 sw
rect 42986 48930 47134 48931
tri 47134 48930 47135 48931 sw
rect 42986 48929 47135 48930
tri 47135 48929 47136 48930 sw
rect 42986 48928 47136 48929
tri 47136 48928 47137 48929 sw
tri 47226 48928 47430 49132 ne
rect 47430 48928 49118 49132
tri 49118 48928 49410 49220 sw
tri 49410 48928 49702 49220 ne
rect 49702 49215 51142 49220
tri 51142 49215 51395 49468 sw
tri 51429 49215 51682 49468 ne
rect 51682 49335 55524 49468
tri 55524 49335 55815 49626 sw
tri 55815 49335 56126 49646 ne
rect 56126 49401 60024 49646
tri 60024 49401 60309 49686 sw
tri 60309 49487 60508 49686 ne
rect 60508 49487 71000 49686
rect 56126 49335 60309 49401
rect 51682 49215 55815 49335
rect 49702 48928 51395 49215
tri 51395 48928 51682 49215 sw
tri 51682 48928 51969 49215 ne
rect 51969 49030 55815 49215
tri 55815 49030 56120 49335 sw
tri 56126 49321 56140 49335 ne
rect 56140 49321 60309 49335
rect 51969 49010 56120 49030
tri 56120 49010 56140 49030 sw
tri 56140 49010 56451 49321 ne
rect 56451 49202 60309 49321
tri 60309 49202 60508 49401 sw
tri 60508 49285 60710 49487 ne
rect 60710 49285 71000 49487
rect 56451 49010 60508 49202
rect 51969 48928 56140 49010
rect 42986 48835 47137 48928
rect 38640 48640 42689 48835
rect 34369 48379 38352 48640
rect 30090 48120 34101 48353
rect 27849 48091 29800 48120
rect 25595 48076 27560 48091
rect 21248 47882 25298 48076
rect 17200 47877 20966 47882
tri 20966 47877 20971 47882 sw
tri 21248 47877 21253 47882 ne
rect 21253 47877 25298 47882
rect 17200 47595 20971 47877
tri 20971 47595 21253 47877 sw
tri 21253 47595 21535 47877 ne
rect 21535 47779 25298 47877
tri 25298 47779 25595 48076 sw
tri 25595 47907 25764 48076 ne
rect 25764 47907 27560 48076
rect 21535 47610 25595 47779
tri 25595 47610 25764 47779 sw
tri 25764 47610 26061 47907 ne
rect 26061 47802 27560 47907
tri 27560 47802 27849 48091 sw
tri 27849 47802 28138 48091 ne
rect 28138 48020 29800 48091
tri 29800 48020 29900 48120 sw
tri 30090 48020 30190 48120 ne
rect 30190 48085 34101 48120
tri 34101 48085 34369 48353 sw
tri 34369 48085 34663 48379 ne
rect 34663 48352 38352 48379
tri 38352 48352 38640 48640 sw
tri 38640 48379 38901 48640 ne
rect 38901 48538 42689 48640
tri 42689 48538 42986 48835 sw
tri 42986 48647 43174 48835 ne
rect 43174 48647 47137 48835
rect 38901 48379 42986 48538
rect 34663 48091 38640 48352
tri 38640 48091 38901 48352 sw
tri 38901 48091 39189 48379 ne
rect 39189 48350 42986 48379
tri 42986 48350 43174 48538 sw
tri 43174 48380 43441 48647 ne
rect 43441 48635 47137 48647
tri 47137 48635 47430 48928 sw
tri 47430 48647 47711 48928 ne
rect 47711 48647 49410 48928
tri 49410 48647 49691 48928 sw
tri 49702 48647 49983 48928 ne
rect 49983 48647 51682 48928
tri 51682 48647 51963 48928 sw
tri 51969 48647 52250 48928 ne
rect 52250 48702 56140 48928
tri 56140 48702 56448 49010 sw
tri 56451 48760 56701 49010 ne
rect 56701 49000 60508 49010
tri 60508 49000 60710 49202 sw
tri 60710 49200 60795 49285 ne
rect 60795 49200 71000 49285
rect 56701 48760 71000 49000
rect 52250 48647 56448 48702
rect 43441 48380 47430 48635
rect 39189 48183 43174 48350
tri 43174 48183 43341 48350 sw
tri 43441 48183 43638 48380 ne
rect 43638 48354 47430 48380
tri 47430 48354 47711 48635 sw
tri 47711 48380 47978 48647 ne
rect 47978 48380 49691 48647
tri 49691 48380 49958 48647 sw
tri 49983 48380 50250 48647 ne
rect 50250 48380 51963 48647
tri 51963 48380 52230 48647 sw
tri 52250 48380 52517 48647 ne
rect 52517 48450 56448 48647
tri 56448 48450 56700 48702 sw
tri 56701 48540 56921 48760 ne
rect 56921 48540 71000 48760
rect 52517 48380 56700 48450
rect 43638 48183 47711 48354
rect 39189 48091 43341 48183
rect 34663 48085 38901 48091
rect 30190 48020 34369 48085
rect 28138 47829 29900 48020
tri 29900 47829 30091 48020 sw
tri 30190 48019 30191 48020 ne
rect 30191 48019 34369 48020
tri 30191 48018 30192 48019 ne
rect 30192 48018 34369 48019
tri 30192 48017 30193 48018 ne
rect 30193 48017 34369 48018
tri 30193 48016 30194 48017 ne
rect 30194 48016 34369 48017
tri 30194 48015 30195 48016 ne
rect 30195 48015 34369 48016
tri 30195 48014 30196 48015 ne
rect 30196 48014 34369 48015
tri 30196 48013 30197 48014 ne
rect 30197 48013 34369 48014
tri 30197 48012 30198 48013 ne
rect 30198 48012 34369 48013
tri 30198 48011 30199 48012 ne
rect 30199 48011 34369 48012
tri 30199 48010 30200 48011 ne
rect 30200 48010 34369 48011
tri 30200 48009 30201 48010 ne
rect 30201 48009 34369 48010
tri 30201 48008 30202 48009 ne
rect 30202 48008 34369 48009
tri 30202 48007 30203 48008 ne
rect 30203 48007 34369 48008
tri 30203 48006 30204 48007 ne
rect 30204 48006 34369 48007
tri 30204 48005 30205 48006 ne
rect 30205 48005 34369 48006
tri 30205 48004 30206 48005 ne
rect 30206 48004 34369 48005
tri 30206 48003 30207 48004 ne
rect 30207 48003 34369 48004
tri 30207 48002 30208 48003 ne
rect 30208 48002 34369 48003
tri 30208 48001 30209 48002 ne
rect 30209 48001 34369 48002
tri 30209 48000 30210 48001 ne
rect 30210 48000 34369 48001
tri 30210 47999 30211 48000 ne
rect 30211 47999 34369 48000
tri 30211 47998 30212 47999 ne
rect 30212 47998 34369 47999
tri 30212 47997 30213 47998 ne
rect 30213 47997 34369 47998
tri 30213 47996 30214 47997 ne
rect 30214 47996 34369 47997
tri 30214 47995 30215 47996 ne
rect 30215 47995 34369 47996
tri 30215 47994 30216 47995 ne
rect 30216 47994 34369 47995
tri 30216 47993 30217 47994 ne
rect 30217 47993 34369 47994
tri 30217 47992 30218 47993 ne
rect 30218 47992 34369 47993
tri 30218 47991 30219 47992 ne
rect 30219 47991 34369 47992
tri 30219 47990 30220 47991 ne
rect 30220 47990 34369 47991
tri 30220 47989 30221 47990 ne
rect 30221 47989 34369 47990
tri 30221 47988 30222 47989 ne
rect 30222 47988 34369 47989
tri 30222 47987 30223 47988 ne
rect 30223 47987 34369 47988
tri 30223 47986 30224 47987 ne
rect 30224 47986 34369 47987
tri 30224 47985 30225 47986 ne
rect 30225 47985 34369 47986
tri 30225 47984 30226 47985 ne
rect 30226 47984 34369 47985
tri 30226 47983 30227 47984 ne
rect 30227 47983 34369 47984
tri 30227 47982 30228 47983 ne
rect 30228 47982 34369 47983
tri 30228 47981 30229 47982 ne
rect 30229 47981 34369 47982
tri 30229 47980 30230 47981 ne
rect 30230 47980 34369 47981
tri 30230 47979 30231 47980 ne
rect 30231 47979 34369 47980
tri 30231 47978 30232 47979 ne
rect 30232 47978 34369 47979
tri 30232 47977 30233 47978 ne
rect 30233 47977 34369 47978
tri 30233 47976 30234 47977 ne
rect 30234 47976 34369 47977
tri 30234 47975 30235 47976 ne
rect 30235 47975 34369 47976
tri 30235 47974 30236 47975 ne
rect 30236 47974 34369 47975
tri 30236 47973 30237 47974 ne
rect 30237 47973 34369 47974
tri 30237 47972 30238 47973 ne
rect 30238 47972 34369 47973
tri 30238 47971 30239 47972 ne
rect 30239 47971 34369 47972
tri 30239 47970 30240 47971 ne
rect 30240 47970 34369 47971
tri 30240 47969 30241 47970 ne
rect 30241 47969 34369 47970
tri 30241 47968 30242 47969 ne
rect 30242 47968 34369 47969
tri 30242 47967 30243 47968 ne
rect 30243 47967 34369 47968
tri 30243 47966 30244 47967 ne
rect 30244 47966 34369 47967
tri 30244 47965 30245 47966 ne
rect 30245 47965 34369 47966
tri 30245 47964 30246 47965 ne
rect 30246 47964 34369 47965
tri 30246 47963 30247 47964 ne
rect 30247 47963 34369 47964
tri 30247 47962 30248 47963 ne
rect 30248 47962 34369 47963
tri 30248 47961 30249 47962 ne
rect 30249 47961 34369 47962
tri 30249 47960 30250 47961 ne
rect 30250 47960 34369 47961
tri 30250 47959 30251 47960 ne
rect 30251 47959 34369 47960
tri 30251 47958 30252 47959 ne
rect 30252 47958 34369 47959
tri 30252 47957 30253 47958 ne
rect 30253 47957 34369 47958
tri 30253 47956 30254 47957 ne
rect 30254 47956 34369 47957
tri 30254 47955 30255 47956 ne
rect 30255 47955 34369 47956
tri 30255 47954 30256 47955 ne
rect 30256 47954 34369 47955
tri 30256 47953 30257 47954 ne
rect 30257 47953 34369 47954
tri 30257 47952 30258 47953 ne
rect 30258 47952 34369 47953
tri 30258 47951 30259 47952 ne
rect 30259 47951 34369 47952
tri 30259 47950 30260 47951 ne
rect 30260 47950 34369 47951
tri 30260 47949 30261 47950 ne
rect 30261 47949 34369 47950
tri 30261 47948 30262 47949 ne
rect 30262 47948 34369 47949
tri 30262 47947 30263 47948 ne
rect 30263 47947 34369 47948
tri 30263 47946 30264 47947 ne
rect 30264 47946 34369 47947
tri 30264 47945 30265 47946 ne
rect 30265 47945 34369 47946
tri 30265 47944 30266 47945 ne
rect 30266 47944 34369 47945
tri 30266 47943 30267 47944 ne
rect 30267 47943 34369 47944
tri 30267 47942 30268 47943 ne
rect 30268 47942 34369 47943
tri 30268 47941 30269 47942 ne
rect 30269 47941 34369 47942
tri 30269 47940 30270 47941 ne
rect 30270 47940 34369 47941
tri 30270 47939 30271 47940 ne
rect 30271 47939 34369 47940
tri 30271 47938 30272 47939 ne
rect 30272 47938 34369 47939
tri 30272 47937 30273 47938 ne
rect 30273 47937 34369 47938
tri 30273 47936 30274 47937 ne
rect 30274 47936 34369 47937
tri 30274 47935 30275 47936 ne
rect 30275 47935 34369 47936
tri 30275 47934 30276 47935 ne
rect 30276 47934 34369 47935
tri 30276 47933 30277 47934 ne
rect 30277 47933 34369 47934
tri 30277 47932 30278 47933 ne
rect 30278 47932 34369 47933
tri 30278 47931 30279 47932 ne
rect 30279 47931 34369 47932
tri 30279 47930 30280 47931 ne
rect 30280 47930 34369 47931
tri 30280 47929 30281 47930 ne
rect 30281 47929 34369 47930
tri 30281 47928 30282 47929 ne
rect 30282 47928 34369 47929
tri 30282 47927 30283 47928 ne
rect 30283 47927 34369 47928
tri 30283 47926 30284 47927 ne
rect 30284 47926 34369 47927
tri 30284 47925 30285 47926 ne
rect 30285 47925 34369 47926
tri 30285 47924 30286 47925 ne
rect 30286 47924 34369 47925
tri 30286 47923 30287 47924 ne
rect 30287 47923 34369 47924
tri 30287 47922 30288 47923 ne
rect 30288 47922 34369 47923
tri 30288 47921 30289 47922 ne
rect 30289 47921 34369 47922
tri 30289 47920 30290 47921 ne
rect 30290 47920 34369 47921
tri 30290 47919 30291 47920 ne
rect 30291 47919 34369 47920
tri 30291 47918 30292 47919 ne
rect 30292 47918 34369 47919
tri 30292 47917 30293 47918 ne
rect 30293 47917 34369 47918
tri 30293 47916 30294 47917 ne
rect 30294 47916 34369 47917
tri 30294 47915 30295 47916 ne
rect 30295 47915 34369 47916
tri 30295 47914 30296 47915 ne
rect 30296 47914 34369 47915
tri 30296 47913 30297 47914 ne
rect 30297 47913 34369 47914
tri 30297 47912 30298 47913 ne
rect 30298 47912 34369 47913
tri 30298 47911 30299 47912 ne
rect 30299 47911 34369 47912
tri 30299 47910 30300 47911 ne
rect 30300 47910 34369 47911
tri 30300 47909 30301 47910 ne
rect 30301 47909 34369 47910
tri 30301 47908 30302 47909 ne
rect 30302 47908 34369 47909
tri 30302 47907 30303 47908 ne
rect 30303 47907 34369 47908
tri 30303 47906 30304 47907 ne
rect 30304 47906 34369 47907
tri 30304 47905 30305 47906 ne
rect 30305 47905 34369 47906
tri 30305 47904 30306 47905 ne
rect 30306 47904 34369 47905
tri 30306 47903 30307 47904 ne
rect 30307 47903 34369 47904
tri 30307 47902 30308 47903 ne
rect 30308 47902 34369 47903
tri 30308 47901 30309 47902 ne
rect 30309 47901 34369 47902
tri 34369 47901 34553 48085 sw
tri 34663 47901 34847 48085 ne
rect 34847 47901 38901 48085
rect 28138 47802 30091 47829
rect 26061 47610 27849 47802
rect 21535 47595 25764 47610
rect 17200 47404 21253 47595
tri 17200 47312 17292 47404 ne
rect 17292 47313 21253 47404
tri 21253 47313 21535 47595 sw
tri 21535 47594 21536 47595 ne
rect 21536 47594 25764 47595
tri 21536 47404 21726 47594 ne
rect 21726 47404 25764 47594
rect 17292 47312 21535 47313
tri 17000 47020 17292 47312 sw
tri 17292 47111 17493 47312 ne
rect 17493 47122 21535 47312
tri 21535 47122 21726 47313 sw
tri 21726 47190 21940 47404 ne
rect 21940 47313 25764 47404
tri 25764 47313 26061 47610 sw
tri 26061 47609 26062 47610 ne
rect 26062 47609 27849 47610
rect 21940 47312 26061 47313
tri 26061 47312 26062 47313 sw
tri 26062 47312 26359 47609 ne
rect 26359 47600 27849 47609
tri 27849 47600 28051 47802 sw
tri 28138 47600 28340 47802 ne
rect 28340 47730 30091 47802
tri 30091 47730 30190 47829 sw
tri 30309 47730 30480 47901 ne
rect 30480 47730 34553 47901
rect 28340 47601 30190 47730
tri 30190 47601 30319 47730 sw
tri 30480 47601 30609 47730 ne
rect 30609 47607 34553 47730
tri 34553 47607 34847 47901 sw
tri 34847 47607 35141 47901 ne
rect 35141 47889 38901 47901
tri 38901 47889 39103 48091 sw
tri 39189 47889 39391 48091 ne
rect 39391 47889 43341 48091
rect 35141 47607 39103 47889
rect 30609 47601 34847 47607
rect 28340 47600 30319 47601
rect 26359 47312 28051 47600
rect 21940 47190 26062 47312
rect 17493 47111 21726 47122
rect 14000 46908 17292 47020
tri 17292 46908 17404 47020 sw
tri 17493 46908 17696 47111 ne
rect 17696 46908 21726 47111
tri 21726 46908 21940 47122 sw
tri 21940 46982 22148 47190 ne
rect 22148 47015 26062 47190
tri 26062 47015 26359 47312 sw
tri 26359 47078 26593 47312 ne
rect 26593 47311 28051 47312
tri 28051 47311 28340 47600 sw
tri 28340 47311 28629 47600 ne
rect 28629 47311 30319 47600
tri 30319 47311 30609 47601 sw
tri 30609 47311 30899 47601 ne
rect 30899 47313 34847 47601
tri 34847 47313 35141 47607 sw
tri 35141 47606 35142 47607 ne
rect 35142 47606 39103 47607
rect 30899 47312 35141 47313
tri 35141 47312 35142 47313 sw
tri 35142 47312 35436 47606 ne
rect 35436 47601 39103 47606
tri 39103 47601 39391 47889 sw
tri 39391 47601 39679 47889 ne
rect 39679 47886 43341 47889
tri 43341 47886 43638 48183 sw
tri 43638 47886 43935 48183 ne
rect 43935 48087 47711 48183
tri 47711 48087 47978 48354 sw
tri 47978 48179 48179 48380 ne
rect 48179 48179 49958 48380
rect 43935 47886 47978 48087
tri 47978 47886 48179 48087 sw
tri 48179 47886 48472 48179 ne
rect 48472 48178 49958 48179
tri 49958 48178 50160 48380 sw
tri 50250 48178 50452 48380 ne
rect 50452 48178 52230 48380
rect 48472 47886 50160 48178
tri 50160 47886 50452 48178 sw
tri 50452 47886 50744 48178 ne
rect 50744 48173 52230 48178
tri 52230 48173 52437 48380 sw
tri 52517 48173 52724 48380 ne
rect 52724 48229 56700 48380
tri 56700 48229 56921 48450 sw
tri 56921 48380 57081 48540 ne
rect 57081 48380 71000 48540
rect 52724 48173 56921 48229
rect 50744 47886 52437 48173
tri 52437 47886 52724 48173 sw
tri 52724 47886 53011 48173 ne
rect 53011 48071 56921 48173
tri 56921 48071 57079 48229 sw
tri 57081 48206 57255 48380 ne
rect 57255 48206 71000 48380
rect 53011 47895 57079 48071
tri 57079 47895 57255 48071 sw
tri 57255 47895 57566 48206 ne
rect 57566 47895 71000 48206
rect 53011 47886 57255 47895
rect 39679 47601 43638 47886
rect 35436 47313 39391 47601
tri 39391 47313 39679 47601 sw
tri 39679 47600 39680 47601 ne
rect 39680 47600 43638 47601
rect 35436 47312 39679 47313
tri 39679 47312 39680 47313 sw
tri 39680 47312 39968 47600 ne
rect 39968 47589 43638 47600
tri 43638 47589 43935 47886 sw
tri 43935 47885 43936 47886 ne
rect 43936 47885 48179 47886
rect 39968 47588 43935 47589
tri 43935 47588 43936 47589 sw
tri 43936 47588 44233 47885 ne
rect 44233 47593 48179 47885
tri 48179 47593 48472 47886 sw
tri 48472 47605 48753 47886 ne
rect 48753 47605 50452 47886
rect 44233 47588 48472 47593
rect 39968 47312 43936 47588
rect 30899 47311 35142 47312
rect 26593 47078 28340 47311
rect 22148 46982 26359 47015
rect 14000 46616 17404 46908
tri 17404 46616 17696 46908 sw
tri 17696 46616 17988 46908 ne
rect 17988 46700 21940 46908
tri 21940 46700 22148 46908 sw
tri 22148 46700 22430 46982 ne
rect 22430 46781 26359 46982
tri 26359 46781 26593 47015 sw
tri 26593 46781 26890 47078 ne
rect 26890 47069 28340 47078
tri 28340 47069 28582 47311 sw
tri 28629 47069 28871 47311 ne
rect 28871 47070 30609 47311
tri 30609 47070 30850 47311 sw
tri 30899 47070 31140 47311 ne
rect 31140 47070 35142 47311
rect 28871 47069 30850 47070
rect 26890 46781 28582 47069
rect 22430 46700 26593 46781
rect 17988 46616 22148 46700
rect 14000 46324 17696 46616
tri 17696 46324 17988 46616 sw
tri 17988 46335 18269 46616 ne
rect 18269 46418 22148 46616
tri 22148 46418 22430 46700 sw
tri 22430 46699 22431 46700 ne
rect 22431 46699 26593 46700
rect 18269 46417 22430 46418
tri 22430 46417 22431 46418 sw
tri 22431 46417 22713 46699 ne
rect 22713 46484 26593 46699
tri 26593 46484 26890 46781 sw
tri 26890 46700 26971 46781 ne
rect 26971 46780 28582 46781
tri 28582 46780 28871 47069 sw
tri 28871 46780 29160 47069 ne
rect 29160 46780 30850 47069
tri 30850 46780 31140 47070 sw
tri 31140 46780 31430 47070 ne
rect 31430 47018 35142 47070
tri 35142 47018 35436 47312 sw
tri 35436 47075 35673 47312 ne
rect 35673 47075 39680 47312
rect 31430 46781 35436 47018
tri 35436 46781 35673 47018 sw
tri 35673 46781 35967 47075 ne
rect 35967 47024 39680 47075
tri 39680 47024 39968 47312 sw
tri 39968 47069 40211 47312 ne
rect 40211 47291 43936 47312
tri 43936 47291 44233 47588 sw
tri 44233 47311 44510 47588 ne
rect 44510 47312 48472 47588
tri 48472 47312 48753 47593 sw
tri 48753 47312 49046 47605 ne
rect 49046 47603 50452 47605
tri 50452 47603 50735 47886 sw
tri 50744 47603 51027 47886 ne
rect 51027 47603 52724 47886
rect 49046 47312 50735 47603
rect 44510 47311 48753 47312
rect 40211 47069 44233 47291
rect 35967 46781 39968 47024
tri 39968 46781 40211 47024 sw
tri 40211 46976 40304 47069 ne
rect 40304 47014 44233 47069
tri 44233 47014 44510 47291 sw
tri 44510 47078 44743 47311 ne
rect 44743 47078 48753 47311
rect 40304 46976 44510 47014
rect 31430 46780 35673 46781
rect 26971 46700 28871 46780
tri 28871 46700 28951 46780 sw
tri 29160 46700 29240 46780 ne
rect 29240 46700 31140 46780
tri 31140 46700 31220 46780 sw
tri 31430 46700 31510 46780 ne
rect 31510 46700 35673 46780
rect 22713 46417 26890 46484
rect 18269 46335 22431 46417
rect 14000 46068 17988 46324
tri 14000 42080 17988 46068 ne
tri 17988 46043 18269 46324 sw
tri 18269 46068 18536 46335 ne
rect 18536 46135 22431 46335
tri 22431 46135 22713 46417 sw
tri 22713 46315 22815 46417 ne
rect 22815 46403 26890 46417
tri 26890 46403 26971 46484 sw
tri 26971 46482 27189 46700 ne
rect 27189 46689 28951 46700
tri 28951 46689 28962 46700 sw
tri 29240 46689 29251 46700 ne
rect 29251 46689 31220 46700
rect 27189 46482 28962 46689
rect 22815 46315 26971 46403
rect 18536 46068 22713 46135
rect 17988 45776 18269 46043
tri 18269 45776 18536 46043 sw
tri 18536 46042 18562 46068 ne
rect 18562 46042 22713 46068
rect 17988 45750 18536 45776
tri 18536 45750 18562 45776 sw
tri 18562 45750 18854 46042 ne
rect 18854 46033 22713 46042
tri 22713 46033 22815 46135 sw
tri 22815 46033 23097 46315 ne
rect 23097 46185 26971 46315
tri 26971 46185 27189 46403 sw
tri 27189 46185 27486 46482 ne
rect 27486 46400 28962 46482
tri 28962 46400 29251 46689 sw
tri 29251 46400 29540 46689 ne
rect 29540 46481 31220 46689
tri 31220 46481 31439 46700 sw
tri 31510 46481 31729 46700 ne
rect 31729 46487 35673 46700
tri 35673 46487 35967 46781 sw
tri 35967 46681 36067 46781 ne
rect 36067 46688 40211 46781
tri 40211 46688 40304 46781 sw
tri 40304 46689 40591 46976 ne
rect 40591 46781 44510 46976
tri 44510 46781 44743 47014 sw
tri 44743 46781 45040 47078 ne
rect 45040 47019 48753 47078
tri 48753 47019 49046 47312 sw
tri 49046 47234 49124 47312 ne
rect 49124 47311 50735 47312
tri 50735 47311 51027 47603 sw
tri 51027 47311 51319 47603 ne
rect 51319 47599 52724 47603
tri 52724 47599 53011 47886 sw
tri 53011 47599 53298 47886 ne
rect 53298 47599 57255 47886
rect 51319 47598 53011 47599
tri 53011 47598 53012 47599 sw
tri 53298 47598 53299 47599 ne
rect 53299 47598 57255 47599
rect 51319 47311 53012 47598
tri 53012 47311 53299 47598 sw
tri 53299 47311 53586 47598 ne
rect 53586 47587 57255 47598
tri 57255 47587 57563 47895 sw
tri 57566 47632 57829 47895 ne
rect 57829 47632 71000 47895
rect 53586 47321 57563 47587
tri 57563 47321 57829 47587 sw
tri 57829 47364 58097 47632 ne
rect 58097 47364 71000 47632
rect 53586 47311 57829 47321
rect 49124 47234 51027 47311
rect 45040 46941 49046 47019
tri 49046 46941 49124 47019 sw
tri 49124 46941 49417 47234 ne
rect 49417 47053 51027 47234
tri 51027 47053 51285 47311 sw
tri 51319 47053 51577 47311 ne
rect 51577 47053 53299 47311
tri 53299 47053 53557 47311 sw
tri 53586 47053 53844 47311 ne
rect 53844 47053 57829 47311
tri 57829 47053 58097 47321 sw
tri 58097 47261 58200 47364 ne
rect 58200 47261 71000 47364
tri 58200 47053 58408 47261 ne
rect 58408 47053 71000 47261
rect 49417 46941 51285 47053
rect 45040 46781 49124 46941
rect 40591 46689 44743 46781
rect 36067 46681 40304 46688
rect 31729 46481 35967 46487
rect 29540 46400 31439 46481
rect 27486 46185 29251 46400
rect 23097 46033 27189 46185
rect 18854 45751 22815 46033
tri 22815 45751 23097 46033 sw
tri 23097 46032 23098 46033 ne
rect 23098 46032 27189 46033
rect 18854 45750 23097 45751
tri 23097 45750 23098 45751 sw
tri 23098 45750 23380 46032 ne
rect 23380 45888 27189 46032
tri 27189 45888 27486 46185 sw
tri 27486 46047 27624 46185 ne
rect 27624 46111 29251 46185
tri 29251 46111 29540 46400 sw
tri 29540 46111 29829 46400 ne
rect 29829 46399 31439 46400
tri 31439 46399 31521 46481 sw
tri 31729 46399 31811 46481 ne
rect 31811 46399 35967 46481
rect 29829 46111 31521 46399
rect 27624 46047 29540 46111
rect 23380 45750 27486 45888
tri 27486 45750 27624 45888 sw
tri 27624 45864 27807 46047 ne
rect 27807 46038 29540 46047
tri 29540 46038 29613 46111 sw
tri 29829 46038 29902 46111 ne
rect 29902 46109 31521 46111
tri 31521 46109 31811 46399 sw
tri 31811 46109 32101 46399 ne
rect 32101 46387 35967 46399
tri 35967 46387 36067 46487 sw
tri 36067 46399 36349 46681 ne
rect 36349 46401 40304 46681
tri 40304 46401 40591 46688 sw
tri 40591 46401 40879 46689 ne
rect 40879 46484 44743 46689
tri 44743 46484 45040 46781 sw
tri 45040 46698 45123 46781 ne
rect 45123 46698 49124 46781
rect 40879 46401 45040 46484
tri 45040 46401 45123 46484 sw
tri 45123 46401 45420 46698 ne
rect 45420 46648 49124 46698
tri 49124 46648 49417 46941 sw
tri 49417 46700 49658 46941 ne
rect 49658 46940 51285 46941
tri 51285 46940 51398 47053 sw
tri 51577 46940 51690 47053 ne
rect 51690 46940 53557 47053
tri 53557 46940 53670 47053 sw
rect 49658 46780 51398 46940
tri 51398 46780 51558 46940 sw
tri 51690 46780 51850 46940 ne
rect 51850 46780 53670 46940
tri 53670 46780 53830 46940 sw
rect 49658 46771 51558 46780
tri 51558 46771 51567 46780 sw
tri 51850 46771 51859 46780 ne
rect 51859 46771 53830 46780
tri 53830 46771 53839 46780 sw
rect 49658 46700 51567 46771
tri 51567 46700 51638 46771 sw
tri 51859 46700 51930 46771 ne
rect 51930 46766 53839 46771
tri 53839 46766 53844 46771 sw
tri 53844 46766 54131 47053 ne
rect 54131 46766 58097 47053
rect 51930 46700 53844 46766
rect 45420 46407 49417 46648
tri 49417 46407 49658 46648 sw
tri 49658 46646 49712 46700 ne
rect 49712 46646 51638 46700
rect 45420 46401 49658 46407
rect 36349 46399 40591 46401
rect 32101 46109 36067 46387
rect 29902 46039 31811 46109
tri 31811 46039 31881 46109 sw
tri 32101 46039 32171 46109 ne
rect 32171 46105 36067 46109
tri 36067 46105 36349 46387 sw
tri 36349 46105 36643 46399 ne
rect 36643 46113 40591 46399
tri 40591 46113 40879 46401 sw
tri 40879 46399 40881 46401 ne
rect 40881 46399 45123 46401
rect 36643 46111 40879 46113
tri 40879 46111 40881 46113 sw
tri 40881 46111 41169 46399 ne
rect 41169 46111 45123 46399
rect 36643 46105 40881 46111
rect 32171 46039 36349 46105
rect 29902 46038 31881 46039
rect 27807 45864 29613 46038
rect 17988 45656 18562 45750
tri 18562 45656 18656 45750 sw
tri 18854 45656 18948 45750 ne
rect 18948 45656 23098 45750
rect 17988 45364 18656 45656
tri 18656 45364 18948 45656 sw
tri 18948 45364 19240 45656 ne
rect 19240 45582 23098 45656
tri 23098 45582 23266 45750 sw
tri 23380 45582 23548 45750 ne
rect 23548 45749 27624 45750
tri 27624 45749 27625 45750 sw
tri 27807 45749 27922 45864 ne
rect 27922 45749 29613 45864
tri 29613 45749 29902 46038 sw
tri 29902 45749 30191 46038 ne
rect 30191 45749 31881 46038
tri 31881 45749 32171 46039 sw
tri 32171 45749 32461 46039 ne
rect 32461 45811 36349 46039
tri 36349 45811 36643 46105 sw
tri 36643 46044 36704 46105 ne
rect 36704 46044 40881 46105
rect 32461 45750 36643 45811
tri 36643 45750 36704 45811 sw
tri 36704 45750 36998 46044 ne
rect 36998 45823 40881 46044
tri 40881 45823 41169 46111 sw
tri 41169 45932 41348 46111 ne
rect 41348 46104 45123 46111
tri 45123 46104 45420 46401 sw
tri 45420 46229 45592 46401 ne
rect 45592 46353 49658 46401
tri 49658 46353 49712 46407 sw
tri 49712 46400 49958 46646 ne
rect 49958 46560 51638 46646
tri 51638 46560 51778 46700 sw
tri 51930 46560 52070 46700 ne
rect 52070 46560 53844 46700
tri 53844 46560 54050 46766 sw
tri 54131 46560 54337 46766 ne
rect 54337 46751 58097 46766
tri 58097 46751 58399 47053 sw
tri 58408 46940 58521 47053 ne
rect 58521 46940 71000 47053
rect 54337 46630 58399 46751
tri 58399 46630 58520 46751 sw
tri 58521 46700 58761 46940 ne
rect 58761 46700 71000 46940
rect 54337 46560 58520 46630
rect 49958 46400 51778 46560
tri 51778 46400 51938 46560 sw
tri 52070 46400 52230 46560 ne
rect 52230 46400 54050 46560
rect 45592 46229 49712 46353
rect 41348 45932 45420 46104
tri 45420 45932 45592 46104 sw
tri 45592 46047 45774 46229 ne
rect 45774 46107 49712 46229
tri 49712 46107 49958 46353 sw
tri 49958 46107 50251 46400 ne
rect 50251 46268 51938 46400
tri 51938 46268 52070 46400 sw
tri 52230 46268 52362 46400 ne
rect 52362 46399 54050 46400
tri 54050 46399 54211 46560 sw
tri 54337 46399 54498 46560 ne
rect 54498 46399 58520 46560
rect 52362 46268 54211 46399
rect 50251 46107 52070 46268
rect 45774 46047 49958 46107
tri 45774 45932 45889 46047 ne
rect 45889 45932 49958 46047
rect 36998 45750 41169 45823
rect 32461 45749 36704 45750
rect 23548 45582 27625 45749
rect 19240 45364 23266 45582
rect 17988 45072 18948 45364
tri 18948 45072 19240 45364 sw
tri 19240 45363 19241 45364 ne
rect 19241 45363 23266 45364
rect 17988 45071 19240 45072
tri 19240 45071 19241 45072 sw
tri 19241 45071 19533 45363 ne
rect 19533 45300 23266 45363
tri 23266 45300 23548 45582 sw
tri 23548 45374 23756 45582 ne
rect 23756 45452 27625 45582
tri 27625 45452 27922 45749 sw
tri 27922 45657 28014 45749 ne
rect 28014 45657 29902 45749
rect 23756 45451 27922 45452
tri 27922 45451 27923 45452 sw
rect 23756 45450 27923 45451
tri 27923 45450 27924 45451 sw
rect 23756 45449 27924 45450
tri 27924 45449 27925 45450 sw
rect 23756 45448 27925 45449
tri 27925 45448 27926 45449 sw
rect 23756 45447 27926 45448
tri 27926 45447 27927 45448 sw
rect 23756 45446 27927 45447
tri 27927 45446 27928 45447 sw
rect 23756 45445 27928 45446
tri 27928 45445 27929 45446 sw
rect 23756 45444 27929 45445
tri 27929 45444 27930 45445 sw
rect 23756 45443 27930 45444
tri 27930 45443 27931 45444 sw
rect 23756 45442 27931 45443
tri 27931 45442 27932 45443 sw
rect 23756 45441 27932 45442
tri 27932 45441 27933 45442 sw
rect 23756 45440 27933 45441
tri 27933 45440 27934 45441 sw
rect 23756 45439 27934 45440
tri 27934 45439 27935 45440 sw
rect 23756 45438 27935 45439
tri 27935 45438 27936 45439 sw
rect 23756 45437 27936 45438
tri 27936 45437 27937 45438 sw
rect 23756 45436 27937 45437
tri 27937 45436 27938 45437 sw
rect 23756 45435 27938 45436
tri 27938 45435 27939 45436 sw
rect 23756 45434 27939 45435
tri 27939 45434 27940 45435 sw
rect 23756 45433 27940 45434
tri 27940 45433 27941 45434 sw
rect 23756 45432 27941 45433
tri 27941 45432 27942 45433 sw
rect 23756 45431 27942 45432
tri 27942 45431 27943 45432 sw
rect 23756 45430 27943 45431
tri 27943 45430 27944 45431 sw
rect 23756 45429 27944 45430
tri 27944 45429 27945 45430 sw
rect 23756 45428 27945 45429
tri 27945 45428 27946 45429 sw
rect 23756 45427 27946 45428
tri 27946 45427 27947 45428 sw
rect 23756 45426 27947 45427
tri 27947 45426 27948 45427 sw
rect 23756 45425 27948 45426
tri 27948 45425 27949 45426 sw
rect 23756 45424 27949 45425
tri 27949 45424 27950 45425 sw
rect 23756 45423 27950 45424
tri 27950 45423 27951 45424 sw
rect 23756 45422 27951 45423
tri 27951 45422 27952 45423 sw
rect 23756 45421 27952 45422
tri 27952 45421 27953 45422 sw
rect 23756 45420 27953 45421
tri 27953 45420 27954 45421 sw
rect 23756 45419 27954 45420
tri 27954 45419 27955 45420 sw
rect 23756 45418 27955 45419
tri 27955 45418 27956 45419 sw
rect 23756 45417 27956 45418
tri 27956 45417 27957 45418 sw
rect 23756 45416 27957 45417
tri 27957 45416 27958 45417 sw
rect 23756 45415 27958 45416
tri 27958 45415 27959 45416 sw
rect 23756 45414 27959 45415
tri 27959 45414 27960 45415 sw
rect 23756 45413 27960 45414
tri 27960 45413 27961 45414 sw
rect 23756 45412 27961 45413
tri 27961 45412 27962 45413 sw
rect 23756 45411 27962 45412
tri 27962 45411 27963 45412 sw
rect 23756 45410 27963 45411
tri 27963 45410 27964 45411 sw
rect 23756 45409 27964 45410
tri 27964 45409 27965 45410 sw
rect 23756 45408 27965 45409
tri 27965 45408 27966 45409 sw
rect 23756 45407 27966 45408
tri 27966 45407 27967 45408 sw
rect 23756 45406 27967 45407
tri 27967 45406 27968 45407 sw
rect 23756 45405 27968 45406
tri 27968 45405 27969 45406 sw
rect 23756 45404 27969 45405
tri 27969 45404 27970 45405 sw
rect 23756 45403 27970 45404
tri 27970 45403 27971 45404 sw
rect 23756 45402 27971 45403
tri 27971 45402 27972 45403 sw
rect 23756 45401 27972 45402
tri 27972 45401 27973 45402 sw
rect 23756 45400 27973 45401
tri 27973 45400 27974 45401 sw
rect 23756 45399 27974 45400
tri 27974 45399 27975 45400 sw
rect 23756 45398 27975 45399
tri 27975 45398 27976 45399 sw
rect 23756 45397 27976 45398
tri 27976 45397 27977 45398 sw
rect 23756 45396 27977 45397
tri 27977 45396 27978 45397 sw
rect 23756 45395 27978 45396
tri 27978 45395 27979 45396 sw
rect 23756 45394 27979 45395
tri 27979 45394 27980 45395 sw
rect 23756 45393 27980 45394
tri 27980 45393 27981 45394 sw
rect 23756 45392 27981 45393
tri 27981 45392 27982 45393 sw
rect 23756 45391 27982 45392
tri 27982 45391 27983 45392 sw
rect 23756 45390 27983 45391
tri 27983 45390 27984 45391 sw
rect 23756 45389 27984 45390
tri 27984 45389 27985 45390 sw
rect 23756 45388 27985 45389
tri 27985 45388 27986 45389 sw
rect 23756 45387 27986 45388
tri 27986 45387 27987 45388 sw
rect 23756 45386 27987 45387
tri 27987 45386 27988 45387 sw
rect 23756 45385 27988 45386
tri 27988 45385 27989 45386 sw
rect 23756 45384 27989 45385
tri 27989 45384 27990 45385 sw
rect 23756 45383 27990 45384
tri 27990 45383 27991 45384 sw
rect 23756 45382 27991 45383
tri 27991 45382 27992 45383 sw
rect 23756 45381 27992 45382
tri 27992 45381 27993 45382 sw
rect 23756 45380 27993 45381
tri 27993 45380 27994 45381 sw
rect 23756 45379 27994 45380
tri 27994 45379 27995 45380 sw
rect 23756 45378 27995 45379
tri 27995 45378 27996 45379 sw
rect 23756 45377 27996 45378
tri 27996 45377 27997 45378 sw
rect 23756 45376 27997 45377
tri 27997 45376 27998 45377 sw
rect 23756 45375 27998 45376
tri 27998 45375 27999 45376 sw
rect 23756 45374 27999 45375
tri 27999 45374 28000 45375 sw
rect 19533 45092 23548 45300
tri 23548 45092 23756 45300 sw
tri 23756 45180 23950 45374 ne
rect 23950 45373 28000 45374
tri 28000 45373 28001 45374 sw
rect 23950 45372 28001 45373
tri 28001 45372 28002 45373 sw
rect 23950 45371 28002 45372
tri 28002 45371 28003 45372 sw
rect 23950 45370 28003 45371
tri 28003 45370 28004 45371 sw
rect 23950 45369 28004 45370
tri 28004 45369 28005 45370 sw
rect 23950 45368 28005 45369
tri 28005 45368 28006 45369 sw
rect 23950 45367 28006 45368
tri 28006 45367 28007 45368 sw
rect 23950 45366 28007 45367
tri 28007 45366 28008 45367 sw
rect 23950 45365 28008 45366
tri 28008 45365 28009 45366 sw
rect 23950 45364 28009 45365
tri 28009 45364 28010 45365 sw
rect 23950 45363 28010 45364
tri 28010 45363 28011 45364 sw
rect 23950 45362 28011 45363
tri 28011 45362 28012 45363 sw
rect 23950 45361 28012 45362
tri 28012 45361 28013 45362 sw
rect 23950 45360 28013 45361
tri 28013 45360 28014 45361 sw
tri 28014 45360 28311 45657 ne
rect 28311 45461 29902 45657
tri 29902 45461 30190 45749 sw
tri 30191 45657 30283 45749 ne
rect 30283 45657 32171 45749
rect 28311 45368 30190 45461
tri 30190 45368 30283 45461 sw
tri 30283 45368 30572 45657 ne
rect 30572 45656 32171 45657
tri 32171 45656 32264 45749 sw
tri 32461 45656 32554 45749 ne
rect 32554 45656 36704 45749
rect 30572 45368 32264 45656
rect 28311 45360 30283 45368
rect 23950 45180 28014 45360
rect 19533 45071 23756 45092
rect 17988 44779 19241 45071
tri 19241 44779 19533 45071 sw
tri 19533 44990 19614 45071 ne
rect 19614 44990 23756 45071
rect 17988 44698 19533 44779
tri 19533 44698 19614 44779 sw
tri 19614 44698 19906 44990 ne
rect 19906 44898 23756 44990
tri 23756 44898 23950 45092 sw
tri 23950 44898 24232 45180 ne
rect 24232 45063 28014 45180
tri 28014 45063 28311 45360 sw
tri 28311 45098 28573 45360 ne
rect 28573 45098 30283 45360
rect 24232 44898 28311 45063
rect 19906 44698 23950 44898
rect 17988 44697 19614 44698
tri 19614 44697 19615 44698 sw
tri 19906 44697 19907 44698 ne
rect 19907 44697 23950 44698
rect 17988 44405 19615 44697
tri 19615 44405 19907 44697 sw
tri 19907 44405 20199 44697 ne
rect 20199 44616 23950 44697
tri 23950 44616 24232 44898 sw
tri 24232 44897 24233 44898 ne
rect 24233 44897 28311 44898
rect 20199 44615 24232 44616
tri 24232 44615 24233 44616 sw
tri 24233 44615 24515 44897 ne
rect 24515 44801 28311 44897
tri 28311 44801 28573 45063 sw
tri 28573 44801 28870 45098 ne
rect 28870 45089 30283 45098
tri 30283 45089 30562 45368 sw
tri 30572 45089 30851 45368 ne
rect 30851 45366 32264 45368
tri 32264 45366 32554 45656 sw
tri 32554 45366 32844 45656 ne
rect 32844 45456 36704 45656
tri 36704 45456 36998 45750 sw
tri 36998 45657 37091 45750 ne
rect 37091 45657 41169 45750
rect 32844 45366 36998 45456
rect 30851 45090 32554 45366
tri 32554 45090 32830 45366 sw
tri 32844 45090 33120 45366 ne
rect 33120 45363 36998 45366
tri 36998 45363 37091 45456 sw
tri 37091 45433 37315 45657 ne
rect 37315 45644 41169 45657
tri 41169 45644 41348 45823 sw
tri 41348 45644 41636 45932 ne
rect 41636 45656 45592 45932
tri 45592 45656 45868 45932 sw
tri 45889 45656 46165 45932 ne
rect 46165 45814 49958 45932
tri 49958 45814 50251 46107 sw
tri 50251 46043 50315 46107 ne
rect 50315 46043 52070 46107
rect 46165 45750 50251 45814
tri 50251 45750 50315 45814 sw
tri 50315 45750 50608 46043 ne
rect 50608 46041 52070 46043
tri 52070 46041 52297 46268 sw
tri 52362 46041 52589 46268 ne
rect 52589 46112 54211 46268
tri 54211 46112 54498 46399 sw
tri 54498 46112 54785 46399 ne
rect 54785 46390 58520 46399
tri 58520 46390 58760 46630 sw
tri 58761 46400 59061 46700 ne
rect 59061 46400 71000 46700
rect 54785 46112 58760 46390
rect 52589 46087 54498 46112
tri 54498 46087 54523 46112 sw
tri 54785 46087 54810 46112 ne
rect 54810 46090 58760 46112
tri 58760 46090 59060 46390 sw
tri 59061 46110 59351 46400 ne
rect 59351 46110 71000 46400
rect 54810 46087 59060 46090
rect 52589 46041 54523 46087
rect 50608 45800 52297 46041
tri 52297 45800 52538 46041 sw
tri 52589 45800 52830 46041 ne
rect 52830 45800 54523 46041
tri 54523 45800 54810 46087 sw
tri 54810 45800 55097 46087 ne
rect 55097 45800 59060 46087
tri 59060 45800 59350 46090 sw
tri 59351 46000 59461 46110 ne
rect 59461 46000 71000 46110
rect 50608 45750 52538 45800
rect 46165 45656 50315 45750
rect 41636 45644 45868 45656
rect 37315 45433 41348 45644
rect 33120 45139 37091 45363
tri 37091 45139 37315 45363 sw
tri 37315 45139 37609 45433 ne
rect 37609 45356 41348 45433
tri 41348 45356 41636 45644 sw
tri 41636 45368 41912 45644 ne
rect 41912 45368 45868 45644
rect 37609 45139 41636 45356
rect 33120 45090 37315 45139
rect 30851 45089 32830 45090
rect 28870 44801 30562 45089
rect 24515 44615 28573 44801
rect 20199 44405 24233 44615
rect 17988 44113 19907 44405
tri 19907 44113 20199 44405 sw
tri 20199 44404 20200 44405 ne
rect 20200 44404 24233 44405
rect 17988 44112 20199 44113
tri 20199 44112 20200 44113 sw
tri 20200 44112 20492 44404 ne
rect 20492 44333 24233 44404
tri 24233 44333 24515 44615 sw
tri 24515 44613 24517 44615 ne
rect 24517 44613 28573 44615
rect 20492 44331 24515 44333
tri 24515 44331 24517 44333 sw
tri 24517 44331 24799 44613 ne
rect 24799 44504 28573 44613
tri 28573 44504 28870 44801 sw
tri 28870 44614 29057 44801 ne
rect 29057 44800 30562 44801
tri 30562 44800 30851 45089 sw
tri 30851 44800 31140 45089 ne
rect 31140 44800 32830 45089
tri 32830 44800 33120 45090 sw
tri 33120 44800 33410 45090 ne
rect 33410 44845 37315 45090
tri 37315 44845 37609 45139 sw
tri 37609 45095 37653 45139 ne
rect 37653 45095 41636 45139
rect 33410 44801 37609 44845
tri 37609 44801 37653 44845 sw
tri 37653 44801 37947 45095 ne
rect 37947 45080 41636 45095
tri 41636 45080 41912 45356 sw
tri 41912 45089 42191 45368 ne
rect 42191 45359 45868 45368
tri 45868 45359 46165 45656 sw
tri 46165 45359 46462 45656 ne
rect 46462 45457 50315 45656
tri 50315 45457 50608 45750 sw
tri 50608 45657 50701 45750 ne
rect 50701 45749 52538 45750
tri 52538 45749 52589 45800 sw
tri 52830 45749 52881 45800 ne
rect 52881 45749 54810 45800
rect 50701 45728 52589 45749
tri 52589 45728 52610 45749 sw
tri 52881 45728 52902 45749 ne
rect 52902 45728 54810 45749
rect 50701 45657 52610 45728
tri 52610 45657 52681 45728 sw
tri 52902 45657 52973 45728 ne
rect 52973 45657 54810 45728
tri 54810 45657 54953 45800 sw
tri 55097 45657 55240 45800 ne
rect 55240 45739 71000 45800
rect 55240 45657 70613 45739
rect 46462 45364 50608 45457
tri 50608 45364 50701 45457 sw
tri 50701 45364 50994 45657 ne
rect 50994 45365 52681 45657
tri 52681 45365 52973 45657 sw
tri 52973 45365 53265 45657 ne
rect 53265 45512 54953 45657
tri 54953 45512 55098 45657 sw
tri 55240 45512 55385 45657 ne
rect 55385 45512 70613 45657
rect 53265 45365 55098 45512
rect 50994 45364 52973 45365
rect 46462 45359 50701 45364
rect 42191 45089 46165 45359
rect 37947 44801 41912 45080
tri 41912 44801 42191 45080 sw
tri 42191 44801 42479 45089 ne
rect 42479 45062 46165 45089
tri 46165 45062 46462 45359 sw
tri 46462 45098 46723 45359 ne
rect 46723 45098 50701 45359
rect 42479 44801 46462 45062
tri 46462 44801 46723 45062 sw
tri 46723 44801 47020 45098 ne
rect 47020 45071 50701 45098
tri 50701 45071 50994 45364 sw
tri 50994 45181 51177 45364 ne
rect 51177 45252 52973 45364
tri 52973 45252 53086 45365 sw
tri 53265 45252 53378 45365 ne
rect 53378 45252 55098 45365
rect 51177 45181 53086 45252
rect 47020 44888 50994 45071
tri 50994 44888 51177 45071 sw
tri 51177 44960 51398 45181 ne
rect 51398 44960 53086 45181
tri 53086 44960 53378 45252 sw
tri 53378 44960 53670 45252 ne
rect 53670 45247 55098 45252
tri 55098 45247 55363 45512 sw
tri 55385 45247 55650 45512 ne
rect 55650 45247 70613 45512
rect 53670 44960 55363 45247
tri 55363 44960 55650 45247 sw
tri 55650 44960 55937 45247 ne
rect 55937 44960 70613 45247
rect 47020 44887 51177 44888
tri 51177 44887 51178 44888 sw
rect 47020 44886 51178 44887
tri 51178 44886 51179 44887 sw
rect 47020 44885 51179 44886
tri 51179 44885 51180 44886 sw
rect 47020 44884 51180 44885
tri 51180 44884 51181 44885 sw
rect 47020 44883 51181 44884
tri 51181 44883 51182 44884 sw
rect 47020 44882 51182 44883
tri 51182 44882 51183 44883 sw
rect 47020 44881 51183 44882
tri 51183 44881 51184 44882 sw
rect 47020 44880 51184 44881
tri 51184 44880 51185 44881 sw
rect 47020 44879 51185 44880
tri 51185 44879 51186 44880 sw
rect 47020 44878 51186 44879
tri 51186 44878 51187 44879 sw
rect 47020 44877 51187 44878
tri 51187 44877 51188 44878 sw
rect 47020 44876 51188 44877
tri 51188 44876 51189 44877 sw
rect 47020 44875 51189 44876
tri 51189 44875 51190 44876 sw
rect 47020 44874 51190 44875
tri 51190 44874 51191 44875 sw
rect 47020 44873 51191 44874
tri 51191 44873 51192 44874 sw
rect 47020 44872 51192 44873
tri 51192 44872 51193 44873 sw
rect 47020 44871 51193 44872
tri 51193 44871 51194 44872 sw
rect 47020 44870 51194 44871
tri 51194 44870 51195 44871 sw
rect 47020 44869 51195 44870
tri 51195 44869 51196 44870 sw
rect 47020 44868 51196 44869
tri 51196 44868 51197 44869 sw
rect 47020 44867 51197 44868
tri 51197 44867 51198 44868 sw
rect 47020 44866 51198 44867
tri 51198 44866 51199 44867 sw
rect 47020 44865 51199 44866
tri 51199 44865 51200 44866 sw
rect 47020 44864 51200 44865
tri 51200 44864 51201 44865 sw
rect 47020 44863 51201 44864
tri 51201 44863 51202 44864 sw
rect 47020 44862 51202 44863
tri 51202 44862 51203 44863 sw
rect 47020 44861 51203 44862
tri 51203 44861 51204 44862 sw
rect 47020 44860 51204 44861
tri 51204 44860 51205 44861 sw
rect 47020 44859 51205 44860
tri 51205 44859 51206 44860 sw
rect 47020 44858 51206 44859
tri 51206 44858 51207 44859 sw
rect 47020 44857 51207 44858
tri 51207 44857 51208 44858 sw
rect 47020 44856 51208 44857
tri 51208 44856 51209 44857 sw
rect 47020 44855 51209 44856
tri 51209 44855 51210 44856 sw
rect 47020 44854 51210 44855
tri 51210 44854 51211 44855 sw
rect 47020 44853 51211 44854
tri 51211 44853 51212 44854 sw
rect 47020 44852 51212 44853
tri 51212 44852 51213 44853 sw
rect 47020 44851 51213 44852
tri 51213 44851 51214 44852 sw
rect 47020 44850 51214 44851
tri 51214 44850 51215 44851 sw
rect 47020 44849 51215 44850
tri 51215 44849 51216 44850 sw
rect 47020 44848 51216 44849
tri 51216 44848 51217 44849 sw
rect 47020 44847 51217 44848
tri 51217 44847 51218 44848 sw
rect 47020 44846 51218 44847
tri 51218 44846 51219 44847 sw
rect 47020 44845 51219 44846
tri 51219 44845 51220 44846 sw
rect 47020 44844 51220 44845
tri 51220 44844 51221 44845 sw
rect 47020 44843 51221 44844
tri 51221 44843 51222 44844 sw
rect 47020 44842 51222 44843
tri 51222 44842 51223 44843 sw
rect 47020 44841 51223 44842
tri 51223 44841 51224 44842 sw
rect 47020 44840 51224 44841
tri 51224 44840 51225 44841 sw
rect 47020 44839 51225 44840
tri 51225 44839 51226 44840 sw
rect 47020 44838 51226 44839
tri 51226 44838 51227 44839 sw
rect 47020 44837 51227 44838
tri 51227 44837 51228 44838 sw
rect 47020 44836 51228 44837
tri 51228 44836 51229 44837 sw
rect 47020 44835 51229 44836
tri 51229 44835 51230 44836 sw
rect 47020 44834 51230 44835
tri 51230 44834 51231 44835 sw
rect 47020 44833 51231 44834
tri 51231 44833 51232 44834 sw
rect 47020 44832 51232 44833
tri 51232 44832 51233 44833 sw
rect 47020 44831 51233 44832
tri 51233 44831 51234 44832 sw
rect 47020 44830 51234 44831
tri 51234 44830 51235 44831 sw
rect 47020 44829 51235 44830
tri 51235 44829 51236 44830 sw
rect 47020 44828 51236 44829
tri 51236 44828 51237 44829 sw
rect 47020 44827 51237 44828
tri 51237 44827 51238 44828 sw
rect 47020 44826 51238 44827
tri 51238 44826 51239 44827 sw
rect 47020 44825 51239 44826
tri 51239 44825 51240 44826 sw
rect 47020 44824 51240 44825
tri 51240 44824 51241 44825 sw
rect 47020 44823 51241 44824
tri 51241 44823 51242 44824 sw
rect 47020 44822 51242 44823
tri 51242 44822 51243 44823 sw
rect 47020 44821 51243 44822
tri 51243 44821 51244 44822 sw
rect 47020 44820 51244 44821
tri 51244 44820 51245 44821 sw
rect 47020 44819 51245 44820
tri 51245 44819 51246 44820 sw
rect 47020 44818 51246 44819
tri 51246 44818 51247 44819 sw
rect 47020 44817 51247 44818
tri 51247 44817 51248 44818 sw
rect 47020 44816 51248 44817
tri 51248 44816 51249 44817 sw
rect 47020 44815 51249 44816
tri 51249 44815 51250 44816 sw
rect 47020 44814 51250 44815
tri 51250 44814 51251 44815 sw
rect 47020 44813 51251 44814
tri 51251 44813 51252 44814 sw
rect 47020 44812 51252 44813
tri 51252 44812 51253 44813 sw
rect 47020 44811 51253 44812
tri 51253 44811 51254 44812 sw
rect 47020 44810 51254 44811
tri 51254 44810 51255 44811 sw
rect 47020 44809 51255 44810
tri 51255 44809 51256 44810 sw
rect 47020 44808 51256 44809
tri 51256 44808 51257 44809 sw
rect 47020 44807 51257 44808
tri 51257 44807 51258 44808 sw
rect 47020 44806 51258 44807
tri 51258 44806 51259 44807 sw
rect 47020 44805 51259 44806
tri 51259 44805 51260 44806 sw
rect 47020 44804 51260 44805
tri 51260 44804 51261 44805 sw
rect 47020 44803 51261 44804
tri 51261 44803 51262 44804 sw
rect 47020 44802 51262 44803
tri 51262 44802 51263 44803 sw
rect 47020 44801 51263 44802
tri 51263 44801 51264 44802 sw
rect 33410 44800 37653 44801
rect 29057 44614 30851 44800
tri 30851 44614 31037 44800 sw
tri 31140 44614 31326 44800 ne
rect 31326 44614 33120 44800
tri 33120 44614 33306 44800 sw
tri 33410 44614 33596 44800 ne
rect 33596 44614 37653 44800
rect 24799 44331 28870 44504
rect 20492 44330 24517 44331
tri 24517 44330 24518 44331 sw
tri 24799 44330 24800 44331 ne
rect 24800 44330 28870 44331
rect 20492 44112 24518 44330
rect 17988 43820 20200 44112
tri 20200 43820 20492 44112 sw
tri 20492 44000 20604 44112 ne
rect 20604 44048 24518 44112
tri 24518 44048 24800 44330 sw
tri 24800 44048 25082 44330 ne
rect 25082 44317 28870 44330
tri 28870 44317 29057 44504 sw
tri 29057 44502 29169 44614 ne
rect 29169 44502 31037 44614
rect 25082 44205 29057 44317
tri 29057 44205 29169 44317 sw
tri 29169 44205 29466 44502 ne
rect 29466 44420 31037 44502
tri 31037 44420 31231 44614 sw
tri 31326 44420 31520 44614 ne
rect 31520 44420 33306 44614
rect 29466 44205 31231 44420
rect 25082 44204 29169 44205
tri 29169 44204 29170 44205 sw
rect 25082 44203 29170 44204
tri 29170 44203 29171 44204 sw
rect 25082 44202 29171 44203
tri 29171 44202 29172 44203 sw
rect 25082 44201 29172 44202
tri 29172 44201 29173 44202 sw
rect 25082 44200 29173 44201
tri 29173 44200 29174 44201 sw
rect 25082 44199 29174 44200
tri 29174 44199 29175 44200 sw
rect 25082 44198 29175 44199
tri 29175 44198 29176 44199 sw
rect 25082 44197 29176 44198
tri 29176 44197 29177 44198 sw
rect 25082 44196 29177 44197
tri 29177 44196 29178 44197 sw
rect 25082 44195 29178 44196
tri 29178 44195 29179 44196 sw
rect 25082 44194 29179 44195
tri 29179 44194 29180 44195 sw
rect 25082 44193 29180 44194
tri 29180 44193 29181 44194 sw
rect 25082 44192 29181 44193
tri 29181 44192 29182 44193 sw
rect 25082 44191 29182 44192
tri 29182 44191 29183 44192 sw
rect 25082 44190 29183 44191
tri 29183 44190 29184 44191 sw
rect 25082 44189 29184 44190
tri 29184 44189 29185 44190 sw
rect 25082 44188 29185 44189
tri 29185 44188 29186 44189 sw
rect 25082 44187 29186 44188
tri 29186 44187 29187 44188 sw
rect 25082 44186 29187 44187
tri 29187 44186 29188 44187 sw
rect 25082 44185 29188 44186
tri 29188 44185 29189 44186 sw
rect 25082 44184 29189 44185
tri 29189 44184 29190 44185 sw
rect 25082 44183 29190 44184
tri 29190 44183 29191 44184 sw
rect 25082 44182 29191 44183
tri 29191 44182 29192 44183 sw
rect 25082 44181 29192 44182
tri 29192 44181 29193 44182 sw
rect 25082 44180 29193 44181
tri 29193 44180 29194 44181 sw
rect 25082 44179 29194 44180
tri 29194 44179 29195 44180 sw
rect 25082 44178 29195 44179
tri 29195 44178 29196 44179 sw
rect 25082 44177 29196 44178
tri 29196 44177 29197 44178 sw
rect 25082 44176 29197 44177
tri 29197 44176 29198 44177 sw
rect 25082 44175 29198 44176
tri 29198 44175 29199 44176 sw
rect 25082 44174 29199 44175
tri 29199 44174 29200 44175 sw
rect 25082 44173 29200 44174
tri 29200 44173 29201 44174 sw
rect 25082 44172 29201 44173
tri 29201 44172 29202 44173 sw
rect 25082 44171 29202 44172
tri 29202 44171 29203 44172 sw
rect 25082 44170 29203 44171
tri 29203 44170 29204 44171 sw
rect 25082 44169 29204 44170
tri 29204 44169 29205 44170 sw
rect 25082 44168 29205 44169
tri 29205 44168 29206 44169 sw
rect 25082 44167 29206 44168
tri 29206 44167 29207 44168 sw
rect 25082 44166 29207 44167
tri 29207 44166 29208 44167 sw
rect 25082 44165 29208 44166
tri 29208 44165 29209 44166 sw
rect 25082 44164 29209 44165
tri 29209 44164 29210 44165 sw
rect 25082 44163 29210 44164
tri 29210 44163 29211 44164 sw
rect 25082 44162 29211 44163
tri 29211 44162 29212 44163 sw
rect 25082 44161 29212 44162
tri 29212 44161 29213 44162 sw
rect 25082 44160 29213 44161
tri 29213 44160 29214 44161 sw
rect 25082 44159 29214 44160
tri 29214 44159 29215 44160 sw
rect 25082 44158 29215 44159
tri 29215 44158 29216 44159 sw
rect 25082 44157 29216 44158
tri 29216 44157 29217 44158 sw
rect 25082 44156 29217 44157
tri 29217 44156 29218 44157 sw
rect 25082 44155 29218 44156
tri 29218 44155 29219 44156 sw
rect 25082 44154 29219 44155
tri 29219 44154 29220 44155 sw
rect 25082 44153 29220 44154
tri 29220 44153 29221 44154 sw
rect 25082 44152 29221 44153
tri 29221 44152 29222 44153 sw
rect 25082 44151 29222 44152
tri 29222 44151 29223 44152 sw
rect 25082 44150 29223 44151
tri 29223 44150 29224 44151 sw
rect 25082 44149 29224 44150
tri 29224 44149 29225 44150 sw
rect 25082 44148 29225 44149
tri 29225 44148 29226 44149 sw
rect 25082 44147 29226 44148
tri 29226 44147 29227 44148 sw
rect 25082 44146 29227 44147
tri 29227 44146 29228 44147 sw
rect 25082 44145 29228 44146
tri 29228 44145 29229 44146 sw
rect 25082 44144 29229 44145
tri 29229 44144 29230 44145 sw
rect 25082 44143 29230 44144
tri 29230 44143 29231 44144 sw
rect 25082 44142 29231 44143
tri 29231 44142 29232 44143 sw
rect 25082 44141 29232 44142
tri 29232 44141 29233 44142 sw
rect 25082 44140 29233 44141
tri 29233 44140 29234 44141 sw
rect 25082 44139 29234 44140
tri 29234 44139 29235 44140 sw
rect 25082 44138 29235 44139
tri 29235 44138 29236 44139 sw
rect 25082 44137 29236 44138
tri 29236 44137 29237 44138 sw
rect 25082 44136 29237 44137
tri 29237 44136 29238 44137 sw
rect 25082 44135 29238 44136
tri 29238 44135 29239 44136 sw
rect 25082 44134 29239 44135
tri 29239 44134 29240 44135 sw
rect 25082 44133 29240 44134
tri 29240 44133 29241 44134 sw
rect 25082 44132 29241 44133
tri 29241 44132 29242 44133 sw
rect 25082 44131 29242 44132
tri 29242 44131 29243 44132 sw
rect 25082 44130 29243 44131
tri 29243 44130 29244 44131 sw
rect 25082 44129 29244 44130
tri 29244 44129 29245 44130 sw
rect 25082 44128 29245 44129
tri 29245 44128 29246 44129 sw
rect 25082 44127 29246 44128
tri 29246 44127 29247 44128 sw
rect 25082 44126 29247 44127
tri 29247 44126 29248 44127 sw
rect 25082 44125 29248 44126
tri 29248 44125 29249 44126 sw
rect 25082 44124 29249 44125
tri 29249 44124 29250 44125 sw
rect 25082 44123 29250 44124
tri 29250 44123 29251 44124 sw
rect 25082 44122 29251 44123
tri 29251 44122 29252 44123 sw
rect 25082 44121 29252 44122
tri 29252 44121 29253 44122 sw
rect 25082 44120 29253 44121
tri 29253 44120 29254 44121 sw
rect 25082 44119 29254 44120
tri 29254 44119 29255 44120 sw
rect 25082 44118 29255 44119
tri 29255 44118 29256 44119 sw
rect 25082 44117 29256 44118
tri 29256 44117 29257 44118 sw
rect 25082 44116 29257 44117
tri 29257 44116 29258 44117 sw
rect 25082 44115 29258 44116
tri 29258 44115 29259 44116 sw
rect 25082 44114 29259 44115
tri 29259 44114 29260 44115 sw
rect 25082 44113 29260 44114
tri 29260 44113 29261 44114 sw
rect 25082 44112 29261 44113
tri 29261 44112 29262 44113 sw
rect 25082 44111 29262 44112
tri 29262 44111 29263 44112 sw
rect 25082 44110 29263 44111
tri 29263 44110 29264 44111 sw
rect 25082 44109 29264 44110
tri 29264 44109 29265 44110 sw
rect 25082 44108 29265 44109
tri 29265 44108 29266 44109 sw
rect 25082 44107 29266 44108
tri 29266 44107 29267 44108 sw
rect 25082 44106 29267 44107
tri 29267 44106 29268 44107 sw
rect 25082 44105 29268 44106
tri 29268 44105 29269 44106 sw
rect 25082 44104 29269 44105
tri 29269 44104 29270 44105 sw
rect 25082 44103 29270 44104
tri 29270 44103 29271 44104 sw
rect 25082 44102 29271 44103
tri 29271 44102 29272 44103 sw
rect 25082 44101 29272 44102
tri 29272 44101 29273 44102 sw
rect 25082 44100 29273 44101
tri 29273 44100 29274 44101 sw
rect 25082 44099 29274 44100
tri 29274 44099 29275 44100 sw
rect 25082 44098 29275 44099
tri 29275 44098 29276 44099 sw
rect 25082 44097 29276 44098
tri 29276 44097 29277 44098 sw
rect 25082 44096 29277 44097
tri 29277 44096 29278 44097 sw
rect 25082 44095 29278 44096
tri 29278 44095 29279 44096 sw
rect 25082 44094 29279 44095
tri 29279 44094 29280 44095 sw
rect 25082 44093 29280 44094
tri 29280 44093 29281 44094 sw
rect 25082 44092 29281 44093
tri 29281 44092 29282 44093 sw
rect 25082 44091 29282 44092
tri 29282 44091 29283 44092 sw
rect 25082 44090 29283 44091
tri 29283 44090 29284 44091 sw
rect 25082 44089 29284 44090
tri 29284 44089 29285 44090 sw
rect 25082 44088 29285 44089
tri 29285 44088 29286 44089 sw
rect 25082 44087 29286 44088
tri 29286 44087 29287 44088 sw
rect 25082 44086 29287 44087
tri 29287 44086 29288 44087 sw
rect 25082 44085 29288 44086
tri 29288 44085 29289 44086 sw
rect 25082 44084 29289 44085
tri 29289 44084 29290 44085 sw
rect 25082 44083 29290 44084
tri 29290 44083 29291 44084 sw
rect 25082 44082 29291 44083
tri 29291 44082 29292 44083 sw
rect 25082 44081 29292 44082
tri 29292 44081 29293 44082 sw
rect 25082 44080 29293 44081
tri 29293 44080 29294 44081 sw
rect 25082 44079 29294 44080
tri 29294 44079 29295 44080 sw
rect 25082 44078 29295 44079
tri 29295 44078 29296 44079 sw
rect 25082 44077 29296 44078
tri 29296 44077 29297 44078 sw
rect 25082 44076 29297 44077
tri 29297 44076 29298 44077 sw
rect 25082 44075 29298 44076
tri 29298 44075 29299 44076 sw
rect 25082 44074 29299 44075
tri 29299 44074 29300 44075 sw
rect 25082 44073 29300 44074
tri 29300 44073 29301 44074 sw
rect 25082 44072 29301 44073
tri 29301 44072 29302 44073 sw
rect 25082 44071 29302 44072
tri 29302 44071 29303 44072 sw
rect 25082 44070 29303 44071
tri 29303 44070 29304 44071 sw
rect 25082 44069 29304 44070
tri 29304 44069 29305 44070 sw
rect 25082 44068 29305 44069
tri 29305 44068 29306 44069 sw
rect 25082 44067 29306 44068
tri 29306 44067 29307 44068 sw
rect 25082 44066 29307 44067
tri 29307 44066 29308 44067 sw
rect 25082 44065 29308 44066
tri 29308 44065 29309 44066 sw
rect 25082 44064 29309 44065
tri 29309 44064 29310 44065 sw
rect 25082 44063 29310 44064
tri 29310 44063 29311 44064 sw
rect 25082 44062 29311 44063
tri 29311 44062 29312 44063 sw
rect 25082 44061 29312 44062
tri 29312 44061 29313 44062 sw
rect 25082 44060 29313 44061
tri 29313 44060 29314 44061 sw
rect 25082 44059 29314 44060
tri 29314 44059 29315 44060 sw
rect 25082 44058 29315 44059
tri 29315 44058 29316 44059 sw
rect 25082 44057 29316 44058
tri 29316 44057 29317 44058 sw
rect 25082 44056 29317 44057
tri 29317 44056 29318 44057 sw
rect 25082 44055 29318 44056
tri 29318 44055 29319 44056 sw
rect 25082 44054 29319 44055
tri 29319 44054 29320 44055 sw
rect 25082 44053 29320 44054
tri 29320 44053 29321 44054 sw
rect 25082 44052 29321 44053
tri 29321 44052 29322 44053 sw
rect 25082 44051 29322 44052
tri 29322 44051 29323 44052 sw
rect 25082 44050 29323 44051
tri 29323 44050 29324 44051 sw
rect 25082 44049 29324 44050
tri 29324 44049 29325 44050 sw
rect 25082 44048 29325 44049
tri 29325 44048 29326 44049 sw
rect 20604 44000 24800 44048
rect 17988 43708 20492 43820
tri 20492 43708 20604 43820 sw
tri 20604 43818 20786 44000 ne
rect 20786 43818 24800 44000
tri 20786 43708 20896 43818 ne
rect 20896 43766 24800 43818
tri 24800 43766 25082 44048 sw
tri 25082 44047 25083 44048 ne
rect 25083 44047 29326 44048
tri 29326 44047 29327 44048 sw
rect 20896 43765 25082 43766
tri 25082 43765 25083 43766 sw
tri 25083 43765 25365 44047 ne
rect 25365 44046 29327 44047
tri 29327 44046 29328 44047 sw
rect 25365 44045 29328 44046
tri 29328 44045 29329 44046 sw
rect 25365 44044 29329 44045
tri 29329 44044 29330 44045 sw
rect 25365 44043 29330 44044
tri 29330 44043 29331 44044 sw
rect 25365 44042 29331 44043
tri 29331 44042 29332 44043 sw
rect 25365 44041 29332 44042
tri 29332 44041 29333 44042 sw
rect 25365 44040 29333 44041
tri 29333 44040 29334 44041 sw
rect 25365 44039 29334 44040
tri 29334 44039 29335 44040 sw
rect 25365 44038 29335 44039
tri 29335 44038 29336 44039 sw
rect 25365 44037 29336 44038
tri 29336 44037 29337 44038 sw
rect 25365 44036 29337 44037
tri 29337 44036 29338 44037 sw
rect 25365 44035 29338 44036
tri 29338 44035 29339 44036 sw
rect 25365 44034 29339 44035
tri 29339 44034 29340 44035 sw
rect 25365 44033 29340 44034
tri 29340 44033 29341 44034 sw
rect 25365 44032 29341 44033
tri 29341 44032 29342 44033 sw
rect 25365 44031 29342 44032
tri 29342 44031 29343 44032 sw
rect 25365 44030 29343 44031
tri 29343 44030 29344 44031 sw
rect 25365 44029 29344 44030
tri 29344 44029 29345 44030 sw
rect 25365 44028 29345 44029
tri 29345 44028 29346 44029 sw
rect 25365 44027 29346 44028
tri 29346 44027 29347 44028 sw
rect 25365 44026 29347 44027
tri 29347 44026 29348 44027 sw
rect 25365 44025 29348 44026
tri 29348 44025 29349 44026 sw
rect 25365 44024 29349 44025
tri 29349 44024 29350 44025 sw
rect 25365 44023 29350 44024
tri 29350 44023 29351 44024 sw
rect 25365 44022 29351 44023
tri 29351 44022 29352 44023 sw
rect 25365 44021 29352 44022
tri 29352 44021 29353 44022 sw
rect 25365 44020 29353 44021
tri 29353 44020 29354 44021 sw
rect 25365 44019 29354 44020
tri 29354 44019 29355 44020 sw
rect 25365 44018 29355 44019
tri 29355 44018 29356 44019 sw
rect 25365 44017 29356 44018
tri 29356 44017 29357 44018 sw
rect 25365 44016 29357 44017
tri 29357 44016 29358 44017 sw
rect 25365 44015 29358 44016
tri 29358 44015 29359 44016 sw
rect 25365 44014 29359 44015
tri 29359 44014 29360 44015 sw
rect 25365 44013 29360 44014
tri 29360 44013 29361 44014 sw
rect 25365 44012 29361 44013
tri 29361 44012 29362 44013 sw
rect 25365 44011 29362 44012
tri 29362 44011 29363 44012 sw
rect 25365 44010 29363 44011
tri 29363 44010 29364 44011 sw
rect 25365 44009 29364 44010
tri 29364 44009 29365 44010 sw
rect 25365 44008 29365 44009
tri 29365 44008 29366 44009 sw
rect 25365 44007 29366 44008
tri 29366 44007 29367 44008 sw
rect 25365 44006 29367 44007
tri 29367 44006 29368 44007 sw
rect 25365 44005 29368 44006
tri 29368 44005 29369 44006 sw
rect 25365 44004 29369 44005
tri 29369 44004 29370 44005 sw
rect 25365 44003 29370 44004
tri 29370 44003 29371 44004 sw
rect 25365 44002 29371 44003
tri 29371 44002 29372 44003 sw
rect 25365 44001 29372 44002
tri 29372 44001 29373 44002 sw
rect 25365 44000 29373 44001
tri 29373 44000 29374 44001 sw
rect 25365 43999 29374 44000
tri 29374 43999 29375 44000 sw
rect 25365 43998 29375 43999
tri 29375 43998 29376 43999 sw
rect 25365 43997 29376 43998
tri 29376 43997 29377 43998 sw
rect 25365 43996 29377 43997
tri 29377 43996 29378 43997 sw
rect 25365 43995 29378 43996
tri 29378 43995 29379 43996 sw
rect 25365 43994 29379 43995
tri 29379 43994 29380 43995 sw
rect 25365 43993 29380 43994
tri 29380 43993 29381 43994 sw
rect 25365 43992 29381 43993
tri 29381 43992 29382 43993 sw
rect 25365 43991 29382 43992
tri 29382 43991 29383 43992 sw
rect 25365 43990 29383 43991
tri 29383 43990 29384 43991 sw
rect 25365 43989 29384 43990
tri 29384 43989 29385 43990 sw
rect 25365 43988 29385 43989
tri 29385 43988 29386 43989 sw
rect 25365 43987 29386 43988
tri 29386 43987 29387 43988 sw
rect 25365 43986 29387 43987
tri 29387 43986 29388 43987 sw
rect 25365 43985 29388 43986
tri 29388 43985 29389 43986 sw
rect 25365 43984 29389 43985
tri 29389 43984 29390 43985 sw
rect 25365 43983 29390 43984
tri 29390 43983 29391 43984 sw
rect 25365 43982 29391 43983
tri 29391 43982 29392 43983 sw
rect 25365 43981 29392 43982
tri 29392 43981 29393 43982 sw
rect 25365 43980 29393 43981
tri 29393 43980 29394 43981 sw
rect 25365 43979 29394 43980
tri 29394 43979 29395 43980 sw
rect 25365 43978 29395 43979
tri 29395 43978 29396 43979 sw
rect 25365 43977 29396 43978
tri 29396 43977 29397 43978 sw
rect 25365 43976 29397 43977
tri 29397 43976 29398 43977 sw
rect 25365 43975 29398 43976
tri 29398 43975 29399 43976 sw
rect 25365 43974 29399 43975
tri 29399 43974 29400 43975 sw
rect 25365 43973 29400 43974
tri 29400 43973 29401 43974 sw
rect 25365 43972 29401 43973
tri 29401 43972 29402 43973 sw
rect 25365 43971 29402 43972
tri 29402 43971 29403 43972 sw
rect 25365 43970 29403 43971
tri 29403 43970 29404 43971 sw
rect 25365 43969 29404 43970
tri 29404 43969 29405 43970 sw
rect 25365 43968 29405 43969
tri 29405 43968 29406 43969 sw
rect 25365 43967 29406 43968
tri 29406 43967 29407 43968 sw
rect 25365 43966 29407 43967
tri 29407 43966 29408 43967 sw
rect 25365 43965 29408 43966
tri 29408 43965 29409 43966 sw
rect 25365 43964 29409 43965
tri 29409 43964 29410 43965 sw
rect 25365 43963 29410 43964
tri 29410 43963 29411 43964 sw
rect 25365 43962 29411 43963
tri 29411 43962 29412 43963 sw
rect 25365 43961 29412 43962
tri 29412 43961 29413 43962 sw
rect 25365 43960 29413 43961
tri 29413 43960 29414 43961 sw
rect 25365 43959 29414 43960
tri 29414 43959 29415 43960 sw
rect 25365 43958 29415 43959
tri 29415 43958 29416 43959 sw
rect 25365 43957 29416 43958
tri 29416 43957 29417 43958 sw
rect 25365 43956 29417 43957
tri 29417 43956 29418 43957 sw
rect 25365 43955 29418 43956
tri 29418 43955 29419 43956 sw
rect 25365 43954 29419 43955
tri 29419 43954 29420 43955 sw
rect 25365 43953 29420 43954
tri 29420 43953 29421 43954 sw
rect 25365 43952 29421 43953
tri 29421 43952 29422 43953 sw
rect 25365 43951 29422 43952
tri 29422 43951 29423 43952 sw
rect 25365 43950 29423 43951
tri 29423 43950 29424 43951 sw
rect 25365 43949 29424 43950
tri 29424 43949 29425 43950 sw
rect 25365 43948 29425 43949
tri 29425 43948 29426 43949 sw
rect 25365 43947 29426 43948
tri 29426 43947 29427 43948 sw
rect 25365 43946 29427 43947
tri 29427 43946 29428 43947 sw
rect 25365 43945 29428 43946
tri 29428 43945 29429 43946 sw
rect 25365 43944 29429 43945
tri 29429 43944 29430 43945 sw
rect 25365 43943 29430 43944
tri 29430 43943 29431 43944 sw
rect 25365 43942 29431 43943
tri 29431 43942 29432 43943 sw
rect 25365 43941 29432 43942
tri 29432 43941 29433 43942 sw
rect 25365 43940 29433 43941
tri 29433 43940 29434 43941 sw
rect 25365 43939 29434 43940
tri 29434 43939 29435 43940 sw
rect 25365 43938 29435 43939
tri 29435 43938 29436 43939 sw
rect 25365 43937 29436 43938
tri 29436 43937 29437 43938 sw
rect 25365 43936 29437 43937
tri 29437 43936 29438 43937 sw
rect 25365 43935 29438 43936
tri 29438 43935 29439 43936 sw
rect 25365 43934 29439 43935
tri 29439 43934 29440 43935 sw
rect 25365 43933 29440 43934
tri 29440 43933 29441 43934 sw
rect 25365 43932 29441 43933
tri 29441 43932 29442 43933 sw
rect 25365 43931 29442 43932
tri 29442 43931 29443 43932 sw
rect 25365 43930 29443 43931
tri 29443 43930 29444 43931 sw
rect 25365 43929 29444 43930
tri 29444 43929 29445 43930 sw
rect 25365 43928 29445 43929
tri 29445 43928 29446 43929 sw
rect 25365 43927 29446 43928
tri 29446 43927 29447 43928 sw
rect 25365 43926 29447 43927
tri 29447 43926 29448 43927 sw
rect 25365 43925 29448 43926
tri 29448 43925 29449 43926 sw
rect 25365 43924 29449 43925
tri 29449 43924 29450 43925 sw
rect 25365 43923 29450 43924
tri 29450 43923 29451 43924 sw
rect 25365 43922 29451 43923
tri 29451 43922 29452 43923 sw
rect 25365 43921 29452 43922
tri 29452 43921 29453 43922 sw
rect 25365 43920 29453 43921
tri 29453 43920 29454 43921 sw
rect 25365 43919 29454 43920
tri 29454 43919 29455 43920 sw
rect 25365 43918 29455 43919
tri 29455 43918 29456 43919 sw
rect 25365 43917 29456 43918
tri 29456 43917 29457 43918 sw
rect 25365 43916 29457 43917
tri 29457 43916 29458 43917 sw
rect 25365 43915 29458 43916
tri 29458 43915 29459 43916 sw
rect 25365 43914 29459 43915
tri 29459 43914 29460 43915 sw
rect 25365 43913 29460 43914
tri 29460 43913 29461 43914 sw
rect 25365 43912 29461 43913
tri 29461 43912 29462 43913 sw
rect 25365 43911 29462 43912
tri 29462 43911 29463 43912 sw
rect 25365 43910 29463 43911
tri 29463 43910 29464 43911 sw
rect 25365 43909 29464 43910
tri 29464 43909 29465 43910 sw
rect 25365 43908 29465 43909
tri 29465 43908 29466 43909 sw
tri 29466 43908 29763 44205 ne
rect 29763 44131 31231 44205
tri 31231 44131 31520 44420 sw
tri 31520 44131 31809 44420 ne
rect 31809 44419 33306 44420
tri 33306 44419 33501 44614 sw
tri 33596 44419 33791 44614 ne
rect 33791 44507 37653 44614
tri 37653 44507 37947 44801 sw
tri 37947 44614 38134 44801 ne
rect 38134 44614 42191 44801
rect 33791 44419 37947 44507
rect 31809 44131 33501 44419
rect 29763 43908 31520 44131
rect 25365 43765 29466 43908
rect 20896 43708 25083 43765
rect 17988 43416 20604 43708
tri 20604 43416 20896 43708 sw
tri 20896 43451 21153 43708 ne
rect 21153 43483 25083 43708
tri 25083 43483 25365 43765 sw
tri 25365 43714 25416 43765 ne
rect 25416 43714 29466 43765
rect 21153 43451 25365 43483
rect 17988 43159 20896 43416
tri 20896 43159 21153 43416 sw
tri 21153 43159 21445 43451 ne
rect 21445 43432 25365 43451
tri 25365 43432 25416 43483 sw
tri 25416 43432 25698 43714 ne
rect 25698 43611 29466 43714
tri 29466 43611 29763 43908 sw
tri 29763 43758 29913 43908 ne
rect 29913 43842 31520 43908
tri 31520 43842 31809 44131 sw
tri 31809 43842 32098 44131 ne
rect 32098 44129 33501 44131
tri 33501 44129 33791 44419 sw
tri 33791 44129 34081 44419 ne
rect 34081 44320 37947 44419
tri 37947 44320 38134 44507 sw
tri 38134 44419 38329 44614 ne
rect 38329 44513 42191 44614
tri 42191 44513 42479 44801 sw
tri 42479 44614 42666 44801 ne
rect 42666 44614 46723 44801
rect 38329 44419 42479 44513
rect 34081 44129 38134 44320
rect 32098 43842 33791 44129
rect 29913 43758 31809 43842
rect 25698 43461 29763 43611
tri 29763 43461 29913 43611 sw
tri 29913 43461 30210 43758 ne
rect 30210 43553 31809 43758
tri 31809 43553 32098 43842 sw
tri 32098 43553 32387 43842 ne
rect 32387 43839 33791 43842
tri 33791 43839 34081 44129 sw
tri 34081 43839 34371 44129 ne
rect 34371 44125 38134 44129
tri 38134 44125 38329 44320 sw
tri 38329 44125 38623 44419 ne
rect 38623 44326 42479 44419
tri 42479 44326 42666 44513 sw
tri 42666 44396 42884 44614 ne
rect 42884 44504 46723 44614
tri 46723 44504 47020 44801 sw
tri 47020 44590 47231 44801 ne
rect 47231 44800 51264 44801
tri 51264 44800 51265 44801 sw
rect 47231 44799 51265 44800
tri 51265 44799 51266 44800 sw
rect 47231 44798 51266 44799
tri 51266 44798 51267 44799 sw
rect 47231 44797 51267 44798
tri 51267 44797 51268 44798 sw
rect 47231 44796 51268 44797
tri 51268 44796 51269 44797 sw
rect 47231 44795 51269 44796
tri 51269 44795 51270 44796 sw
rect 47231 44794 51270 44795
tri 51270 44794 51271 44795 sw
rect 47231 44793 51271 44794
tri 51271 44793 51272 44794 sw
rect 47231 44792 51272 44793
tri 51272 44792 51273 44793 sw
rect 47231 44791 51273 44792
tri 51273 44791 51274 44792 sw
rect 47231 44790 51274 44791
tri 51274 44790 51275 44791 sw
rect 47231 44789 51275 44790
tri 51275 44789 51276 44790 sw
rect 47231 44788 51276 44789
tri 51276 44788 51277 44789 sw
rect 47231 44787 51277 44788
tri 51277 44787 51278 44788 sw
rect 47231 44786 51278 44787
tri 51278 44786 51279 44787 sw
rect 47231 44785 51279 44786
tri 51279 44785 51280 44786 sw
rect 47231 44784 51280 44785
tri 51280 44784 51281 44785 sw
rect 47231 44783 51281 44784
tri 51281 44783 51282 44784 sw
rect 47231 44782 51282 44783
tri 51282 44782 51283 44783 sw
rect 47231 44781 51283 44782
tri 51283 44781 51284 44782 sw
rect 47231 44780 51284 44781
tri 51284 44780 51285 44781 sw
rect 47231 44779 51285 44780
tri 51285 44779 51286 44780 sw
rect 47231 44778 51286 44779
tri 51286 44778 51287 44779 sw
rect 47231 44777 51287 44778
tri 51287 44777 51288 44778 sw
rect 47231 44776 51288 44777
tri 51288 44776 51289 44777 sw
rect 47231 44775 51289 44776
tri 51289 44775 51290 44776 sw
rect 47231 44774 51290 44775
tri 51290 44774 51291 44775 sw
rect 47231 44773 51291 44774
tri 51291 44773 51292 44774 sw
rect 47231 44772 51292 44773
tri 51292 44772 51293 44773 sw
rect 47231 44771 51293 44772
tri 51293 44771 51294 44772 sw
rect 47231 44770 51294 44771
tri 51294 44770 51295 44771 sw
rect 47231 44769 51295 44770
tri 51295 44769 51296 44770 sw
rect 47231 44768 51296 44769
tri 51296 44768 51297 44769 sw
rect 47231 44767 51297 44768
tri 51297 44767 51298 44768 sw
rect 47231 44766 51298 44767
tri 51298 44766 51299 44767 sw
rect 47231 44765 51299 44766
tri 51299 44765 51300 44766 sw
rect 47231 44764 51300 44765
tri 51300 44764 51301 44765 sw
rect 47231 44763 51301 44764
tri 51301 44763 51302 44764 sw
rect 47231 44762 51302 44763
tri 51302 44762 51303 44763 sw
rect 47231 44761 51303 44762
tri 51303 44761 51304 44762 sw
rect 47231 44760 51304 44761
tri 51304 44760 51305 44761 sw
rect 47231 44759 51305 44760
tri 51305 44759 51306 44760 sw
rect 47231 44758 51306 44759
tri 51306 44758 51307 44759 sw
rect 47231 44757 51307 44758
tri 51307 44757 51308 44758 sw
rect 47231 44756 51308 44757
tri 51308 44756 51309 44757 sw
rect 47231 44755 51309 44756
tri 51309 44755 51310 44756 sw
rect 47231 44754 51310 44755
tri 51310 44754 51311 44755 sw
rect 47231 44753 51311 44754
tri 51311 44753 51312 44754 sw
rect 47231 44752 51312 44753
tri 51312 44752 51313 44753 sw
rect 47231 44751 51313 44752
tri 51313 44751 51314 44752 sw
rect 47231 44750 51314 44751
tri 51314 44750 51315 44751 sw
rect 47231 44749 51315 44750
tri 51315 44749 51316 44750 sw
rect 47231 44748 51316 44749
tri 51316 44748 51317 44749 sw
rect 47231 44747 51317 44748
tri 51317 44747 51318 44748 sw
rect 47231 44746 51318 44747
tri 51318 44746 51319 44747 sw
rect 47231 44745 51319 44746
tri 51319 44745 51320 44746 sw
rect 47231 44744 51320 44745
tri 51320 44744 51321 44745 sw
rect 47231 44743 51321 44744
tri 51321 44743 51322 44744 sw
rect 47231 44742 51322 44743
tri 51322 44742 51323 44743 sw
rect 47231 44741 51323 44742
tri 51323 44741 51324 44742 sw
rect 47231 44740 51324 44741
tri 51324 44740 51325 44741 sw
rect 47231 44739 51325 44740
tri 51325 44739 51326 44740 sw
rect 47231 44738 51326 44739
tri 51326 44738 51327 44739 sw
rect 47231 44737 51327 44738
tri 51327 44737 51328 44738 sw
rect 47231 44736 51328 44737
tri 51328 44736 51329 44737 sw
rect 47231 44735 51329 44736
tri 51329 44735 51330 44736 sw
rect 47231 44734 51330 44735
tri 51330 44734 51331 44735 sw
rect 47231 44733 51331 44734
tri 51331 44733 51332 44734 sw
rect 47231 44732 51332 44733
tri 51332 44732 51333 44733 sw
rect 47231 44731 51333 44732
tri 51333 44731 51334 44732 sw
rect 47231 44730 51334 44731
tri 51334 44730 51335 44731 sw
rect 47231 44729 51335 44730
tri 51335 44729 51336 44730 sw
rect 47231 44728 51336 44729
tri 51336 44728 51337 44729 sw
rect 47231 44727 51337 44728
tri 51337 44727 51338 44728 sw
rect 47231 44726 51338 44727
tri 51338 44726 51339 44727 sw
rect 47231 44725 51339 44726
tri 51339 44725 51340 44726 sw
rect 47231 44724 51340 44725
tri 51340 44724 51341 44725 sw
rect 47231 44723 51341 44724
tri 51341 44723 51342 44724 sw
rect 47231 44722 51342 44723
tri 51342 44722 51343 44723 sw
rect 47231 44721 51343 44722
tri 51343 44721 51344 44722 sw
rect 47231 44720 51344 44721
tri 51344 44720 51345 44721 sw
rect 47231 44719 51345 44720
tri 51345 44719 51346 44720 sw
rect 47231 44718 51346 44719
tri 51346 44718 51347 44719 sw
rect 47231 44717 51347 44718
tri 51347 44717 51348 44718 sw
rect 47231 44716 51348 44717
tri 51348 44716 51349 44717 sw
rect 47231 44715 51349 44716
tri 51349 44715 51350 44716 sw
rect 47231 44714 51350 44715
tri 51350 44714 51351 44715 sw
rect 47231 44713 51351 44714
tri 51351 44713 51352 44714 sw
rect 47231 44712 51352 44713
tri 51352 44712 51353 44713 sw
rect 47231 44711 51353 44712
tri 51353 44711 51354 44712 sw
rect 47231 44710 51354 44711
tri 51354 44710 51355 44711 sw
rect 47231 44709 51355 44710
tri 51355 44709 51356 44710 sw
rect 47231 44708 51356 44709
tri 51356 44708 51357 44709 sw
rect 47231 44707 51357 44708
tri 51357 44707 51358 44708 sw
rect 47231 44706 51358 44707
tri 51358 44706 51359 44707 sw
rect 47231 44705 51359 44706
tri 51359 44705 51360 44706 sw
rect 47231 44704 51360 44705
tri 51360 44704 51361 44705 sw
rect 47231 44703 51361 44704
tri 51361 44703 51362 44704 sw
rect 47231 44702 51362 44703
tri 51362 44702 51363 44703 sw
rect 47231 44701 51363 44702
tri 51363 44701 51364 44702 sw
rect 47231 44700 51364 44701
tri 51364 44700 51365 44701 sw
rect 47231 44699 51365 44700
tri 51365 44699 51366 44700 sw
rect 47231 44698 51366 44699
tri 51366 44698 51367 44699 sw
rect 47231 44697 51367 44698
tri 51367 44697 51368 44698 sw
rect 47231 44696 51368 44697
tri 51368 44696 51369 44697 sw
rect 47231 44695 51369 44696
tri 51369 44695 51370 44696 sw
rect 47231 44694 51370 44695
tri 51370 44694 51371 44695 sw
rect 47231 44693 51371 44694
tri 51371 44693 51372 44694 sw
rect 47231 44692 51372 44693
tri 51372 44692 51373 44693 sw
rect 47231 44691 51373 44692
tri 51373 44691 51374 44692 sw
rect 47231 44690 51374 44691
tri 51374 44690 51375 44691 sw
rect 47231 44689 51375 44690
tri 51375 44689 51376 44690 sw
rect 47231 44688 51376 44689
tri 51376 44688 51377 44689 sw
rect 47231 44687 51377 44688
tri 51377 44687 51378 44688 sw
rect 47231 44686 51378 44687
tri 51378 44686 51379 44687 sw
tri 51398 44686 51672 44960 ne
rect 51672 44686 53378 44960
tri 53378 44686 53652 44960 sw
tri 53670 44686 53944 44960 ne
rect 53944 44686 55650 44960
tri 55650 44686 55924 44960 sw
tri 55937 44686 56211 44960 ne
rect 56211 44686 70613 44960
rect 47231 44590 51379 44686
rect 42884 44396 47020 44504
rect 38623 44125 42666 44326
rect 34371 44124 38329 44125
tri 38329 44124 38330 44125 sw
tri 38623 44124 38624 44125 ne
rect 38624 44124 42666 44125
rect 34371 43839 38330 44124
rect 32387 43737 34081 43839
tri 34081 43737 34183 43839 sw
tri 34371 43737 34473 43839 ne
rect 34473 43830 38330 43839
tri 38330 43830 38624 44124 sw
tri 38624 43830 38918 44124 ne
rect 38918 44108 42666 44124
tri 42666 44108 42884 44326 sw
tri 42884 44108 43172 44396 ne
rect 43172 44293 47020 44396
tri 47020 44293 47231 44504 sw
tri 47231 44419 47402 44590 ne
rect 47402 44419 51379 44590
rect 43172 44122 47231 44293
tri 47231 44122 47402 44293 sw
tri 47402 44122 47699 44419 ne
rect 47699 44393 51379 44419
tri 51379 44393 51672 44686 sw
tri 51672 44420 51938 44686 ne
rect 51938 44420 53652 44686
tri 53652 44420 53918 44686 sw
tri 53944 44420 54210 44686 ne
rect 54210 44420 55924 44686
rect 47699 44127 51672 44393
tri 51672 44127 51938 44393 sw
tri 51938 44127 52231 44420 ne
rect 52231 44288 53918 44420
tri 53918 44288 54050 44420 sw
tri 54210 44288 54342 44420 ne
rect 54342 44419 55924 44420
tri 55924 44419 56191 44686 sw
tri 56211 44419 56478 44686 ne
rect 56478 44419 70613 44686
rect 54342 44288 56191 44419
rect 52231 44127 54050 44288
rect 47699 44122 51938 44127
rect 43172 44108 47402 44122
rect 38918 43830 42884 44108
rect 34473 43737 38624 43830
rect 32387 43553 34183 43737
rect 30210 43461 32098 43553
rect 25698 43432 29913 43461
rect 21445 43159 25416 43432
rect 17988 42867 21153 43159
tri 21153 42867 21445 43159 sw
tri 21445 43158 21446 43159 ne
rect 21446 43158 25416 43159
rect 17988 42866 21445 42867
tri 21445 42866 21446 42867 sw
tri 21446 42866 21738 43158 ne
rect 21738 43150 25416 43158
tri 25416 43150 25698 43432 sw
tri 25698 43431 25699 43432 ne
rect 25699 43431 29913 43432
rect 21738 43149 25698 43150
tri 25698 43149 25699 43150 sw
tri 25699 43149 25981 43431 ne
rect 25981 43164 29913 43431
tri 29913 43164 30210 43461 sw
tri 30210 43460 30211 43461 ne
rect 30211 43460 32098 43461
rect 25981 43163 30210 43164
tri 30210 43163 30211 43164 sw
tri 30211 43163 30508 43460 ne
rect 30508 43443 32098 43460
tri 32098 43443 32208 43553 sw
tri 32387 43443 32497 43553 ne
rect 32497 43486 34183 43553
tri 34183 43486 34434 43737 sw
tri 34473 43486 34724 43737 ne
rect 34724 43536 38624 43737
tri 38624 43536 38918 43830 sw
tri 38918 43750 38998 43830 ne
rect 38998 43820 42884 43830
tri 42884 43820 43172 44108 sw
tri 43172 44107 43173 44108 ne
rect 43173 44107 47402 44108
rect 38998 43819 43172 43820
tri 43172 43819 43173 43820 sw
tri 43173 43819 43461 44107 ne
rect 43461 43825 47402 44107
tri 47402 43825 47699 44122 sw
tri 47699 43940 47881 44122 ne
rect 47881 43940 51938 44122
rect 43461 43819 47699 43825
rect 38998 43750 43173 43819
rect 34724 43486 38918 43536
rect 32497 43446 34434 43486
tri 34434 43446 34474 43486 sw
tri 34724 43446 34764 43486 ne
rect 34764 43456 38918 43486
tri 38918 43456 38998 43536 sw
tri 38998 43456 39292 43750 ne
rect 39292 43531 43173 43750
tri 43173 43531 43461 43819 sw
tri 43461 43732 43548 43819 ne
rect 43548 43732 47699 43819
rect 39292 43456 43461 43531
rect 34764 43446 38998 43456
rect 32497 43443 34474 43446
rect 30508 43163 32208 43443
rect 25981 43149 30211 43163
rect 21738 42867 25699 43149
tri 25699 42867 25981 43149 sw
tri 25981 42946 26184 43149 ne
rect 26184 42946 30211 43149
rect 21738 42866 25981 42867
rect 17988 42574 21446 42866
tri 21446 42574 21738 42866 sw
tri 21738 42664 21940 42866 ne
rect 21940 42664 25981 42866
tri 25981 42664 26184 42867 sw
tri 26184 42790 26340 42946 ne
rect 26340 42866 30211 42946
tri 30211 42866 30508 43163 sw
tri 30508 42866 30805 43163 ne
rect 30805 43154 32208 43163
tri 32208 43154 32497 43443 sw
tri 32497 43154 32786 43443 ne
rect 32786 43156 34474 43443
tri 34474 43156 34764 43446 sw
tri 34764 43156 35054 43446 ne
rect 35054 43162 38998 43446
tri 38998 43162 39292 43456 sw
tri 39292 43455 39293 43456 ne
rect 39293 43455 43461 43456
rect 35054 43161 39292 43162
tri 39292 43161 39293 43162 sw
tri 39293 43161 39587 43455 ne
rect 39587 43444 43461 43455
tri 43461 43444 43548 43531 sw
tri 43548 43444 43836 43732 ne
rect 43836 43643 47699 43732
tri 47699 43643 47881 43825 sw
tri 47881 43643 48178 43940 ne
rect 48178 43834 51938 43940
tri 51938 43834 52231 44127 sw
tri 52231 43936 52422 44127 ne
rect 52422 43996 54050 44127
tri 54050 43996 54342 44288 sw
tri 54342 43996 54634 44288 ne
rect 54634 44132 56191 44288
tri 56191 44132 56478 44419 sw
tri 56478 44132 56765 44419 ne
rect 56765 44132 70613 44419
rect 54634 43996 56478 44132
rect 52422 43936 54342 43996
rect 48178 43643 52231 43834
tri 52231 43643 52422 43834 sw
tri 52422 43643 52715 43936 ne
rect 52715 43935 54342 43936
tri 54342 43935 54403 43996 sw
tri 54634 43935 54695 43996 ne
rect 54695 43935 56478 43996
rect 52715 43643 54403 43935
tri 54403 43643 54695 43935 sw
tri 54695 43643 54987 43935 ne
rect 54987 43930 56478 43935
tri 56478 43930 56680 44132 sw
tri 56765 43930 56967 44132 ne
rect 56967 43930 70613 44132
rect 54987 43643 56680 43930
tri 56680 43643 56967 43930 sw
tri 56967 43643 57254 43930 ne
rect 57254 43643 70613 43930
rect 43836 43642 47881 43643
tri 47881 43642 47882 43643 sw
tri 48178 43642 48179 43643 ne
rect 48179 43642 52422 43643
rect 43836 43444 47882 43642
rect 39587 43161 43548 43444
rect 35054 43156 39293 43161
rect 32786 43155 34764 43156
tri 34764 43155 34765 43156 sw
tri 35054 43155 35055 43156 ne
rect 35055 43155 39293 43156
rect 32786 43154 34765 43155
rect 30805 42866 32497 43154
rect 26340 42790 30508 42866
tri 26340 42664 26466 42790 ne
rect 26466 42664 30508 42790
rect 17988 42372 21738 42574
tri 21738 42372 21940 42574 sw
tri 21940 42372 22232 42664 ne
rect 22232 42456 26184 42664
tri 26184 42456 26392 42664 sw
tri 26466 42456 26674 42664 ne
rect 26674 42569 30508 42664
tri 30508 42569 30805 42866 sw
tri 30805 42820 30851 42866 ne
rect 30851 42865 32497 42866
tri 32497 42865 32786 43154 sw
tri 32786 42865 33075 43154 ne
rect 33075 42865 34765 43154
tri 34765 42865 35055 43155 sw
tri 35055 42865 35345 43155 ne
rect 35345 42867 39293 43155
tri 39293 42867 39587 43161 sw
tri 39587 43160 39588 43161 ne
rect 39588 43160 43548 43161
rect 35345 42866 39587 42867
tri 39587 42866 39588 42867 sw
tri 39588 42866 39882 43160 ne
rect 39882 43156 43548 43160
tri 43548 43156 43836 43444 sw
tri 43836 43443 43837 43444 ne
rect 43837 43443 47882 43444
rect 39882 43155 43836 43156
tri 43836 43155 43837 43156 sw
tri 43837 43155 44125 43443 ne
rect 44125 43345 47882 43443
tri 47882 43345 48179 43642 sw
tri 48179 43345 48476 43642 ne
rect 48476 43350 52422 43642
tri 52422 43350 52715 43643 sw
tri 52715 43350 53008 43643 ne
rect 53008 43351 54695 43643
tri 54695 43351 54987 43643 sw
tri 54987 43351 55279 43643 ne
rect 55279 43642 56967 43643
tri 56967 43642 56968 43643 sw
tri 57254 43642 57255 43643 ne
rect 57255 43642 70613 43643
rect 55279 43355 56968 43642
tri 56968 43355 57255 43642 sw
tri 57255 43355 57542 43642 ne
rect 57542 43355 70613 43642
rect 55279 43351 57255 43355
rect 53008 43350 54987 43351
rect 48476 43345 52715 43350
rect 44125 43155 48179 43345
rect 39882 42867 43837 43155
tri 43837 42867 44125 43155 sw
tri 44125 43020 44260 43155 ne
rect 44260 43048 48179 43155
tri 48179 43048 48476 43345 sw
tri 48476 43163 48658 43345 ne
rect 48658 43163 52715 43345
rect 44260 43020 48476 43048
rect 39882 42866 44125 42867
rect 35345 42865 39588 42866
rect 30851 42820 32786 42865
tri 32786 42820 32831 42865 sw
tri 33075 42820 33120 42865 ne
rect 33120 42820 35055 42865
rect 26674 42523 30805 42569
tri 30805 42523 30851 42569 sw
tri 30851 42523 31148 42820 ne
rect 31148 42796 32831 42820
tri 32831 42796 32855 42820 sw
tri 33120 42796 33144 42820 ne
rect 33144 42818 35055 42820
tri 35055 42818 35102 42865 sw
tri 35345 42818 35392 42865 ne
rect 35392 42818 39588 42865
rect 33144 42796 35102 42818
rect 31148 42528 32855 42796
tri 32855 42528 33123 42796 sw
tri 33144 42528 33412 42796 ne
rect 33412 42528 35102 42796
tri 35102 42528 35392 42818 sw
tri 35392 42528 35682 42818 ne
rect 35682 42572 39588 42818
tri 39588 42572 39882 42866 sw
tri 39882 42732 40016 42866 ne
rect 40016 42732 44125 42866
tri 44125 42732 44260 42867 sw
tri 44260 42817 44463 43020 ne
rect 44463 42866 48476 43020
tri 48476 42866 48658 43048 sw
tri 48658 42866 48955 43163 ne
rect 48955 43057 52715 43163
tri 52715 43057 53008 43350 sw
tri 53008 43274 53084 43350 ne
rect 53084 43274 54987 43350
rect 48955 42981 53008 43057
tri 53008 42981 53084 43057 sw
tri 53084 42981 53377 43274 ne
rect 53377 43240 54987 43274
tri 54987 43240 55098 43351 sw
tri 55279 43240 55390 43351 ne
rect 55390 43267 57255 43351
tri 57255 43267 57343 43355 sw
tri 57542 43267 57630 43355 ne
rect 57630 43267 70613 43355
rect 55390 43240 57343 43267
rect 53377 42981 55098 43240
rect 48955 42866 53084 42981
rect 44463 42817 48658 42866
tri 44463 42732 44548 42817 ne
rect 44548 42732 48658 42817
rect 35682 42528 39882 42572
rect 31148 42523 33123 42528
rect 26674 42456 30851 42523
rect 22232 42372 26392 42456
rect 17988 42080 21940 42372
tri 21940 42080 22232 42372 sw
tri 22232 42164 22440 42372 ne
rect 22440 42174 26392 42372
tri 26392 42174 26674 42456 sw
tri 26674 42174 26956 42456 ne
rect 26956 42226 30851 42456
tri 30851 42226 31148 42523 sw
tri 31148 42457 31214 42523 ne
rect 31214 42507 33123 42523
tri 33123 42507 33144 42528 sw
tri 33412 42507 33433 42528 ne
rect 33433 42507 35392 42528
rect 31214 42457 33144 42507
tri 33144 42457 33194 42507 sw
tri 33433 42457 33483 42507 ne
rect 33483 42457 35392 42507
rect 26956 42174 31148 42226
rect 22440 42164 26674 42174
tri 17988 37836 22232 42080 ne
tri 22232 41872 22440 42080 sw
tri 22440 42000 22604 42164 ne
rect 22604 42000 26674 42164
rect 22232 41708 22440 41872
tri 22440 41708 22604 41872 sw
tri 22604 41708 22896 42000 ne
rect 22896 41892 26674 42000
tri 26674 41892 26956 42174 sw
tri 26956 41980 27150 42174 ne
rect 27150 42160 31148 42174
tri 31148 42160 31214 42226 sw
tri 31214 42160 31511 42457 ne
rect 31511 42440 33194 42457
tri 33194 42440 33211 42457 sw
tri 33483 42440 33500 42457 ne
rect 33500 42440 35392 42457
rect 31511 42160 33211 42440
rect 27150 41980 31214 42160
rect 22896 41708 26956 41892
rect 22232 41416 22604 41708
tri 22604 41416 22896 41708 sw
tri 22896 41707 22897 41708 ne
rect 22897 41707 26956 41708
rect 22232 41415 22896 41416
tri 22896 41415 22897 41416 sw
tri 22897 41415 23189 41707 ne
rect 23189 41698 26956 41707
tri 26956 41698 27150 41892 sw
tri 27150 41698 27432 41980 ne
rect 27432 41863 31214 41980
tri 31214 41863 31511 42160 sw
tri 31511 41917 31754 42160 ne
rect 31754 42151 33211 42160
tri 33211 42151 33500 42440 sw
tri 33500 42151 33789 42440 ne
rect 33789 42238 35392 42440
tri 35392 42238 35682 42528 sw
tri 35682 42238 35972 42528 ne
rect 35972 42438 39882 42528
tri 39882 42438 40016 42572 sw
tri 40016 42438 40310 42732 ne
rect 40310 42444 44260 42732
tri 44260 42444 44548 42732 sw
tri 44548 42528 44752 42732 ne
rect 44752 42569 48658 42732
tri 48658 42569 48955 42866 sw
tri 48955 42820 49001 42866 ne
rect 49001 42820 53084 42866
rect 44752 42528 48955 42569
rect 40310 42438 44548 42444
rect 35972 42238 40016 42438
rect 33789 42237 35682 42238
tri 35682 42237 35683 42238 sw
tri 35972 42237 35973 42238 ne
rect 35973 42237 40016 42238
rect 33789 42151 35683 42237
rect 31754 41917 33500 42151
rect 27432 41698 31511 41863
rect 23189 41416 27150 41698
tri 27150 41416 27432 41698 sw
tri 27432 41697 27433 41698 ne
rect 27433 41697 31511 41698
rect 23189 41415 27432 41416
tri 27432 41415 27433 41416 sw
tri 27433 41415 27715 41697 ne
rect 27715 41620 31511 41697
tri 31511 41620 31754 41863 sw
tri 31754 41712 31959 41917 ne
rect 31959 41862 33500 41917
tri 33500 41862 33789 42151 sw
tri 33789 41862 34078 42151 ne
rect 34078 41947 35683 42151
tri 35683 41947 35973 42237 sw
tri 35973 41947 36263 42237 ne
rect 36263 42144 40016 42237
tri 40016 42144 40310 42438 sw
tri 40310 42145 40603 42438 ne
rect 40603 42240 44548 42438
tri 44548 42240 44752 42444 sw
tri 44752 42439 44841 42528 ne
rect 44841 42523 48955 42528
tri 48955 42523 49001 42569 sw
tri 49001 42528 49293 42820 ne
rect 49293 42688 53084 42820
tri 53084 42688 53377 42981 sw
tri 53377 42820 53538 42981 ne
rect 53538 42980 55098 42981
tri 55098 42980 55358 43240 sw
tri 55390 42980 55650 43240 ne
rect 55650 42980 57343 43240
tri 57343 42980 57630 43267 sw
tri 57630 42980 57917 43267 ne
rect 57917 42980 70613 43267
rect 53538 42820 55358 42980
rect 49293 42687 53377 42688
tri 53377 42687 53378 42688 sw
rect 49293 42686 53378 42687
tri 53378 42686 53379 42687 sw
tri 53538 42686 53672 42820 ne
rect 53672 42800 55358 42820
tri 55358 42800 55538 42980 sw
tri 55650 42800 55830 42980 ne
rect 55830 42800 57630 42980
tri 57630 42800 57810 42980 sw
tri 57917 42800 58097 42980 ne
rect 58097 42875 70613 42980
rect 70669 42875 71000 45739
rect 58097 42800 71000 42875
rect 53672 42686 55538 42800
rect 49293 42528 53379 42686
rect 44841 42439 49001 42523
rect 40603 42151 44752 42240
tri 44752 42151 44841 42240 sw
tri 44841 42151 45129 42439 ne
rect 45129 42231 49001 42439
tri 49001 42231 49293 42523 sw
tri 49293 42439 49382 42528 ne
rect 49382 42439 53379 42528
rect 45129 42151 49293 42231
rect 40603 42145 44841 42151
rect 36263 41947 40310 42144
rect 34078 41862 35973 41947
rect 31959 41712 33789 41862
tri 31959 41620 32051 41712 ne
rect 32051 41703 33789 41712
tri 33789 41703 33948 41862 sw
tri 34078 41703 34237 41862 ne
rect 34237 41704 35973 41862
tri 35973 41704 36216 41947 sw
tri 36263 41704 36506 41947 ne
rect 36506 41851 40310 41947
tri 40310 41851 40603 42144 sw
tri 40603 42075 40673 42145 ne
rect 40673 42075 44841 42145
rect 36506 41781 40603 41851
tri 40603 41781 40673 41851 sw
tri 40673 41781 40967 42075 ne
rect 40967 41863 44841 42075
tri 44841 41863 45129 42151 sw
tri 45129 42063 45217 42151 ne
rect 45217 42142 49293 42151
tri 49293 42142 49382 42231 sw
tri 49382 42142 49679 42439 ne
rect 49679 42393 53379 42439
tri 53379 42393 53672 42686 sw
tri 53672 42440 53918 42686 ne
rect 53918 42528 55538 42686
tri 55538 42528 55810 42800 sw
tri 55830 42528 56102 42800 ne
rect 56102 42600 57810 42800
tri 57810 42600 58010 42800 sw
rect 56102 42528 71000 42600
rect 53918 42507 55810 42528
tri 55810 42507 55831 42528 sw
tri 56102 42507 56123 42528 ne
rect 56123 42507 71000 42528
rect 53918 42457 55831 42507
tri 55831 42457 55881 42507 sw
tri 56123 42457 56173 42507 ne
rect 56173 42497 71000 42507
rect 56173 42457 70613 42497
rect 53918 42440 55881 42457
tri 55881 42440 55898 42457 sw
tri 56173 42440 56190 42457 ne
rect 56190 42440 70613 42457
rect 49679 42147 53672 42393
tri 53672 42147 53918 42393 sw
tri 53918 42147 54211 42440 ne
rect 54211 42308 55898 42440
tri 55898 42308 56030 42440 sw
tri 56190 42308 56322 42440 ne
rect 56322 42308 70613 42440
rect 54211 42147 56030 42308
rect 49679 42142 53918 42147
rect 45217 42063 49382 42142
rect 40967 41781 45129 41863
rect 36506 41780 40673 41781
tri 40673 41780 40674 41781 sw
tri 40967 41780 40968 41781 ne
rect 40968 41780 45129 41781
rect 36506 41704 40674 41780
rect 34237 41703 36216 41704
rect 32051 41620 33948 41703
rect 27715 41619 31754 41620
tri 31754 41619 31755 41620 sw
rect 27715 41618 31755 41619
tri 31755 41618 31756 41619 sw
rect 27715 41617 31756 41618
tri 31756 41617 31757 41618 sw
rect 27715 41616 31757 41617
tri 31757 41616 31758 41617 sw
rect 27715 41615 31758 41616
tri 31758 41615 31759 41616 sw
rect 27715 41614 31759 41615
tri 31759 41614 31760 41615 sw
rect 27715 41613 31760 41614
tri 31760 41613 31761 41614 sw
rect 27715 41612 31761 41613
tri 31761 41612 31762 41613 sw
rect 27715 41611 31762 41612
tri 31762 41611 31763 41612 sw
rect 27715 41610 31763 41611
tri 31763 41610 31764 41611 sw
rect 27715 41609 31764 41610
tri 31764 41609 31765 41610 sw
rect 27715 41608 31765 41609
tri 31765 41608 31766 41609 sw
rect 27715 41607 31766 41608
tri 31766 41607 31767 41608 sw
rect 27715 41606 31767 41607
tri 31767 41606 31768 41607 sw
rect 27715 41605 31768 41606
tri 31768 41605 31769 41606 sw
rect 27715 41604 31769 41605
tri 31769 41604 31770 41605 sw
rect 27715 41603 31770 41604
tri 31770 41603 31771 41604 sw
rect 27715 41602 31771 41603
tri 31771 41602 31772 41603 sw
rect 27715 41601 31772 41602
tri 31772 41601 31773 41602 sw
rect 27715 41600 31773 41601
tri 31773 41600 31774 41601 sw
rect 27715 41599 31774 41600
tri 31774 41599 31775 41600 sw
rect 27715 41598 31775 41599
tri 31775 41598 31776 41599 sw
rect 27715 41597 31776 41598
tri 31776 41597 31777 41598 sw
rect 27715 41596 31777 41597
tri 31777 41596 31778 41597 sw
rect 27715 41595 31778 41596
tri 31778 41595 31779 41596 sw
rect 27715 41594 31779 41595
tri 31779 41594 31780 41595 sw
rect 27715 41593 31780 41594
tri 31780 41593 31781 41594 sw
rect 27715 41592 31781 41593
tri 31781 41592 31782 41593 sw
rect 27715 41591 31782 41592
tri 31782 41591 31783 41592 sw
rect 27715 41590 31783 41591
tri 31783 41590 31784 41591 sw
rect 27715 41589 31784 41590
tri 31784 41589 31785 41590 sw
rect 27715 41588 31785 41589
tri 31785 41588 31786 41589 sw
rect 27715 41587 31786 41588
tri 31786 41587 31787 41588 sw
rect 27715 41586 31787 41587
tri 31787 41586 31788 41587 sw
rect 27715 41585 31788 41586
tri 31788 41585 31789 41586 sw
rect 27715 41584 31789 41585
tri 31789 41584 31790 41585 sw
rect 27715 41583 31790 41584
tri 31790 41583 31791 41584 sw
rect 27715 41582 31791 41583
tri 31791 41582 31792 41583 sw
rect 27715 41581 31792 41582
tri 31792 41581 31793 41582 sw
rect 27715 41580 31793 41581
tri 31793 41580 31794 41581 sw
rect 27715 41579 31794 41580
tri 31794 41579 31795 41580 sw
rect 27715 41578 31795 41579
tri 31795 41578 31796 41579 sw
rect 27715 41577 31796 41578
tri 31796 41577 31797 41578 sw
rect 27715 41576 31797 41577
tri 31797 41576 31798 41577 sw
rect 27715 41575 31798 41576
tri 31798 41575 31799 41576 sw
rect 27715 41574 31799 41575
tri 31799 41574 31800 41575 sw
rect 27715 41573 31800 41574
tri 31800 41573 31801 41574 sw
rect 27715 41572 31801 41573
tri 31801 41572 31802 41573 sw
rect 27715 41571 31802 41572
tri 31802 41571 31803 41572 sw
rect 27715 41570 31803 41571
tri 31803 41570 31804 41571 sw
rect 27715 41569 31804 41570
tri 31804 41569 31805 41570 sw
rect 27715 41568 31805 41569
tri 31805 41568 31806 41569 sw
rect 27715 41567 31806 41568
tri 31806 41567 31807 41568 sw
rect 27715 41566 31807 41567
tri 31807 41566 31808 41567 sw
rect 27715 41565 31808 41566
tri 31808 41565 31809 41566 sw
rect 27715 41564 31809 41565
tri 31809 41564 31810 41565 sw
rect 27715 41563 31810 41564
tri 31810 41563 31811 41564 sw
rect 27715 41562 31811 41563
tri 31811 41562 31812 41563 sw
rect 27715 41561 31812 41562
tri 31812 41561 31813 41562 sw
rect 27715 41560 31813 41561
tri 31813 41560 31814 41561 sw
rect 27715 41559 31814 41560
tri 31814 41559 31815 41560 sw
rect 27715 41558 31815 41559
tri 31815 41558 31816 41559 sw
rect 27715 41557 31816 41558
tri 31816 41557 31817 41558 sw
rect 27715 41556 31817 41557
tri 31817 41556 31818 41557 sw
rect 27715 41555 31818 41556
tri 31818 41555 31819 41556 sw
rect 27715 41554 31819 41555
tri 31819 41554 31820 41555 sw
rect 27715 41553 31820 41554
tri 31820 41553 31821 41554 sw
rect 27715 41552 31821 41553
tri 31821 41552 31822 41553 sw
rect 27715 41551 31822 41552
tri 31822 41551 31823 41552 sw
rect 27715 41550 31823 41551
tri 31823 41550 31824 41551 sw
rect 27715 41549 31824 41550
tri 31824 41549 31825 41550 sw
rect 27715 41548 31825 41549
tri 31825 41548 31826 41549 sw
rect 27715 41547 31826 41548
tri 31826 41547 31827 41548 sw
rect 27715 41546 31827 41547
tri 31827 41546 31828 41547 sw
rect 27715 41545 31828 41546
tri 31828 41545 31829 41546 sw
rect 27715 41544 31829 41545
tri 31829 41544 31830 41545 sw
rect 27715 41543 31830 41544
tri 31830 41543 31831 41544 sw
rect 27715 41542 31831 41543
tri 31831 41542 31832 41543 sw
rect 27715 41541 31832 41542
tri 31832 41541 31833 41542 sw
rect 27715 41540 31833 41541
tri 31833 41540 31834 41541 sw
rect 27715 41539 31834 41540
tri 31834 41539 31835 41540 sw
rect 27715 41538 31835 41539
tri 31835 41538 31836 41539 sw
rect 27715 41537 31836 41538
tri 31836 41537 31837 41538 sw
rect 27715 41536 31837 41537
tri 31837 41536 31838 41537 sw
rect 27715 41535 31838 41536
tri 31838 41535 31839 41536 sw
rect 27715 41534 31839 41535
tri 31839 41534 31840 41535 sw
rect 27715 41533 31840 41534
tri 31840 41533 31841 41534 sw
rect 27715 41532 31841 41533
tri 31841 41532 31842 41533 sw
rect 27715 41531 31842 41532
tri 31842 41531 31843 41532 sw
rect 27715 41530 31843 41531
tri 31843 41530 31844 41531 sw
rect 27715 41529 31844 41530
tri 31844 41529 31845 41530 sw
rect 27715 41528 31845 41529
tri 31845 41528 31846 41529 sw
rect 27715 41527 31846 41528
tri 31846 41527 31847 41528 sw
rect 27715 41526 31847 41527
tri 31847 41526 31848 41527 sw
rect 27715 41525 31848 41526
tri 31848 41525 31849 41526 sw
rect 27715 41524 31849 41525
tri 31849 41524 31850 41525 sw
rect 27715 41523 31850 41524
tri 31850 41523 31851 41524 sw
rect 27715 41522 31851 41523
tri 31851 41522 31852 41523 sw
rect 27715 41521 31852 41522
tri 31852 41521 31853 41522 sw
rect 27715 41520 31853 41521
tri 31853 41520 31854 41521 sw
rect 27715 41519 31854 41520
tri 31854 41519 31855 41520 sw
rect 27715 41518 31855 41519
tri 31855 41518 31856 41519 sw
rect 27715 41517 31856 41518
tri 31856 41517 31857 41518 sw
rect 27715 41516 31857 41517
tri 31857 41516 31858 41517 sw
rect 27715 41515 31858 41516
tri 31858 41515 31859 41516 sw
rect 27715 41514 31859 41515
tri 31859 41514 31860 41515 sw
rect 27715 41513 31860 41514
tri 31860 41513 31861 41514 sw
rect 27715 41512 31861 41513
tri 31861 41512 31862 41513 sw
rect 27715 41511 31862 41512
tri 31862 41511 31863 41512 sw
rect 27715 41510 31863 41511
tri 31863 41510 31864 41511 sw
rect 27715 41509 31864 41510
tri 31864 41509 31865 41510 sw
rect 27715 41508 31865 41509
tri 31865 41508 31866 41509 sw
rect 27715 41507 31866 41508
tri 31866 41507 31867 41508 sw
rect 27715 41506 31867 41507
tri 31867 41506 31868 41507 sw
rect 27715 41505 31868 41506
tri 31868 41505 31869 41506 sw
rect 27715 41504 31869 41505
tri 31869 41504 31870 41505 sw
rect 27715 41503 31870 41504
tri 31870 41503 31871 41504 sw
rect 27715 41502 31871 41503
tri 31871 41502 31872 41503 sw
rect 27715 41501 31872 41502
tri 31872 41501 31873 41502 sw
rect 27715 41500 31873 41501
tri 31873 41500 31874 41501 sw
rect 27715 41499 31874 41500
tri 31874 41499 31875 41500 sw
rect 27715 41498 31875 41499
tri 31875 41498 31876 41499 sw
rect 27715 41497 31876 41498
tri 31876 41497 31877 41498 sw
rect 27715 41496 31877 41497
tri 31877 41496 31878 41497 sw
rect 27715 41495 31878 41496
tri 31878 41495 31879 41496 sw
rect 27715 41494 31879 41495
tri 31879 41494 31880 41495 sw
rect 27715 41493 31880 41494
tri 31880 41493 31881 41494 sw
rect 27715 41492 31881 41493
tri 31881 41492 31882 41493 sw
rect 27715 41491 31882 41492
tri 31882 41491 31883 41492 sw
rect 27715 41490 31883 41491
tri 31883 41490 31884 41491 sw
rect 27715 41489 31884 41490
tri 31884 41489 31885 41490 sw
rect 27715 41488 31885 41489
tri 31885 41488 31886 41489 sw
rect 27715 41487 31886 41488
tri 31886 41487 31887 41488 sw
rect 27715 41486 31887 41487
tri 31887 41486 31888 41487 sw
rect 27715 41485 31888 41486
tri 31888 41485 31889 41486 sw
rect 27715 41484 31889 41485
tri 31889 41484 31890 41485 sw
rect 27715 41483 31890 41484
tri 31890 41483 31891 41484 sw
rect 27715 41482 31891 41483
tri 31891 41482 31892 41483 sw
rect 27715 41481 31892 41482
tri 31892 41481 31893 41482 sw
rect 27715 41480 31893 41481
tri 31893 41480 31894 41481 sw
rect 27715 41479 31894 41480
tri 31894 41479 31895 41480 sw
rect 27715 41478 31895 41479
tri 31895 41478 31896 41479 sw
rect 27715 41477 31896 41478
tri 31896 41477 31897 41478 sw
rect 27715 41476 31897 41477
tri 31897 41476 31898 41477 sw
rect 27715 41475 31898 41476
tri 31898 41475 31899 41476 sw
rect 27715 41474 31899 41475
tri 31899 41474 31900 41475 sw
rect 27715 41473 31900 41474
tri 31900 41473 31901 41474 sw
rect 27715 41472 31901 41473
tri 31901 41472 31902 41473 sw
rect 27715 41471 31902 41472
tri 31902 41471 31903 41472 sw
rect 27715 41470 31903 41471
tri 31903 41470 31904 41471 sw
rect 27715 41469 31904 41470
tri 31904 41469 31905 41470 sw
rect 27715 41468 31905 41469
tri 31905 41468 31906 41469 sw
rect 27715 41467 31906 41468
tri 31906 41467 31907 41468 sw
rect 27715 41466 31907 41467
tri 31907 41466 31908 41467 sw
rect 27715 41465 31908 41466
tri 31908 41465 31909 41466 sw
rect 27715 41464 31909 41465
tri 31909 41464 31910 41465 sw
rect 27715 41463 31910 41464
tri 31910 41463 31911 41464 sw
rect 27715 41462 31911 41463
tri 31911 41462 31912 41463 sw
rect 27715 41461 31912 41462
tri 31912 41461 31913 41462 sw
rect 27715 41460 31913 41461
tri 31913 41460 31914 41461 sw
rect 27715 41459 31914 41460
tri 31914 41459 31915 41460 sw
rect 27715 41458 31915 41459
tri 31915 41458 31916 41459 sw
rect 27715 41457 31916 41458
tri 31916 41457 31917 41458 sw
rect 27715 41456 31917 41457
tri 31917 41456 31918 41457 sw
rect 27715 41455 31918 41456
tri 31918 41455 31919 41456 sw
rect 27715 41454 31919 41455
tri 31919 41454 31920 41455 sw
rect 27715 41453 31920 41454
tri 31920 41453 31921 41454 sw
rect 27715 41452 31921 41453
tri 31921 41452 31922 41453 sw
rect 27715 41451 31922 41452
tri 31922 41451 31923 41452 sw
rect 27715 41450 31923 41451
tri 31923 41450 31924 41451 sw
rect 27715 41449 31924 41450
tri 31924 41449 31925 41450 sw
rect 27715 41448 31925 41449
tri 31925 41448 31926 41449 sw
rect 27715 41447 31926 41448
tri 31926 41447 31927 41448 sw
rect 27715 41446 31927 41447
tri 31927 41446 31928 41447 sw
rect 27715 41445 31928 41446
tri 31928 41445 31929 41446 sw
rect 27715 41444 31929 41445
tri 31929 41444 31930 41445 sw
rect 27715 41443 31930 41444
tri 31930 41443 31931 41444 sw
rect 27715 41442 31931 41443
tri 31931 41442 31932 41443 sw
rect 27715 41441 31932 41442
tri 31932 41441 31933 41442 sw
rect 27715 41440 31933 41441
tri 31933 41440 31934 41441 sw
rect 27715 41439 31934 41440
tri 31934 41439 31935 41440 sw
rect 27715 41438 31935 41439
tri 31935 41438 31936 41439 sw
rect 27715 41437 31936 41438
tri 31936 41437 31937 41438 sw
rect 27715 41436 31937 41437
tri 31937 41436 31938 41437 sw
rect 27715 41435 31938 41436
tri 31938 41435 31939 41436 sw
rect 27715 41434 31939 41435
tri 31939 41434 31940 41435 sw
rect 27715 41433 31940 41434
tri 31940 41433 31941 41434 sw
rect 27715 41432 31941 41433
tri 31941 41432 31942 41433 sw
rect 27715 41431 31942 41432
tri 31942 41431 31943 41432 sw
rect 27715 41430 31943 41431
tri 31943 41430 31944 41431 sw
rect 27715 41429 31944 41430
tri 31944 41429 31945 41430 sw
rect 27715 41428 31945 41429
tri 31945 41428 31946 41429 sw
rect 27715 41427 31946 41428
tri 31946 41427 31947 41428 sw
rect 27715 41426 31947 41427
tri 31947 41426 31948 41427 sw
rect 27715 41425 31948 41426
tri 31948 41425 31949 41426 sw
rect 27715 41424 31949 41425
tri 31949 41424 31950 41425 sw
rect 27715 41423 31950 41424
tri 31950 41423 31951 41424 sw
rect 27715 41422 31951 41423
tri 31951 41422 31952 41423 sw
rect 27715 41421 31952 41422
tri 31952 41421 31953 41422 sw
rect 27715 41420 31953 41421
tri 31953 41420 31954 41421 sw
rect 27715 41419 31954 41420
tri 31954 41419 31955 41420 sw
rect 27715 41418 31955 41419
tri 31955 41418 31956 41419 sw
rect 27715 41417 31956 41418
tri 31956 41417 31957 41418 sw
rect 27715 41416 31957 41417
tri 31957 41416 31958 41417 sw
rect 27715 41415 31958 41416
tri 31958 41415 31959 41416 sw
rect 22232 41123 22897 41415
tri 22897 41123 23189 41415 sw
tri 23189 41287 23317 41415 ne
rect 23317 41287 27433 41415
rect 22232 41120 23189 41123
tri 23189 41120 23192 41123 sw
tri 23317 41120 23484 41287 ne
rect 23484 41133 27433 41287
tri 27433 41133 27715 41415 sw
tri 27715 41286 27844 41415 ne
rect 27844 41414 31959 41415
tri 31959 41414 31960 41415 sw
tri 32051 41414 32257 41620 ne
rect 32257 41414 33948 41620
tri 33948 41414 34237 41703 sw
tri 34237 41414 34526 41703 ne
rect 34526 41414 36216 41703
tri 36216 41414 36506 41704 sw
tri 36506 41414 36796 41704 ne
rect 36796 41486 40674 41704
tri 40674 41486 40968 41780 sw
tri 40968 41486 41262 41780 ne
rect 41262 41775 45129 41780
tri 45129 41775 45217 41863 sw
tri 45217 41775 45505 42063 ne
rect 45505 41845 49382 42063
tri 49382 41845 49679 42142 sw
tri 49679 41985 49836 42142 ne
rect 49836 41985 53918 42142
rect 45505 41775 49679 41845
rect 41262 41688 45217 41775
tri 45217 41688 45304 41775 sw
tri 45505 41688 45592 41775 ne
rect 45592 41688 49679 41775
tri 49679 41688 49836 41845 sw
tri 49836 41783 50038 41985 ne
rect 50038 41854 53918 41985
tri 53918 41854 54211 42147 sw
tri 54211 42073 54285 42147 ne
rect 54285 42073 56030 42147
rect 50038 41783 54211 41854
rect 41262 41486 45304 41688
rect 36796 41414 40968 41486
rect 27844 41286 31960 41414
rect 23484 41120 27715 41133
rect 22232 40828 23192 41120
tri 23192 40828 23484 41120 sw
tri 23484 40828 23776 41120 ne
rect 23776 41004 27715 41120
tri 27715 41004 27844 41133 sw
tri 27844 41004 28126 41286 ne
rect 28126 41117 31960 41286
tri 31960 41117 32257 41414 sw
tri 32257 41138 32533 41414 ne
rect 32533 41138 34237 41414
rect 28126 41116 32257 41117
tri 32257 41116 32258 41117 sw
rect 28126 41115 32258 41116
tri 32258 41115 32259 41116 sw
rect 28126 41114 32259 41115
tri 32259 41114 32260 41115 sw
rect 28126 41113 32260 41114
tri 32260 41113 32261 41114 sw
rect 28126 41112 32261 41113
tri 32261 41112 32262 41113 sw
rect 28126 41111 32262 41112
tri 32262 41111 32263 41112 sw
rect 28126 41110 32263 41111
tri 32263 41110 32264 41111 sw
rect 28126 41109 32264 41110
tri 32264 41109 32265 41110 sw
rect 28126 41108 32265 41109
tri 32265 41108 32266 41109 sw
rect 28126 41107 32266 41108
tri 32266 41107 32267 41108 sw
rect 28126 41106 32267 41107
tri 32267 41106 32268 41107 sw
rect 28126 41105 32268 41106
tri 32268 41105 32269 41106 sw
rect 28126 41104 32269 41105
tri 32269 41104 32270 41105 sw
rect 28126 41103 32270 41104
tri 32270 41103 32271 41104 sw
rect 28126 41102 32271 41103
tri 32271 41102 32272 41103 sw
rect 28126 41101 32272 41102
tri 32272 41101 32273 41102 sw
rect 28126 41100 32273 41101
tri 32273 41100 32274 41101 sw
rect 28126 41099 32274 41100
tri 32274 41099 32275 41100 sw
rect 28126 41098 32275 41099
tri 32275 41098 32276 41099 sw
rect 28126 41097 32276 41098
tri 32276 41097 32277 41098 sw
rect 28126 41096 32277 41097
tri 32277 41096 32278 41097 sw
rect 28126 41095 32278 41096
tri 32278 41095 32279 41096 sw
rect 28126 41094 32279 41095
tri 32279 41094 32280 41095 sw
rect 28126 41093 32280 41094
tri 32280 41093 32281 41094 sw
rect 28126 41092 32281 41093
tri 32281 41092 32282 41093 sw
rect 28126 41091 32282 41092
tri 32282 41091 32283 41092 sw
rect 28126 41090 32283 41091
tri 32283 41090 32284 41091 sw
rect 28126 41089 32284 41090
tri 32284 41089 32285 41090 sw
rect 28126 41088 32285 41089
tri 32285 41088 32286 41089 sw
rect 28126 41087 32286 41088
tri 32286 41087 32287 41088 sw
rect 28126 41086 32287 41087
tri 32287 41086 32288 41087 sw
rect 28126 41085 32288 41086
tri 32288 41085 32289 41086 sw
rect 28126 41084 32289 41085
tri 32289 41084 32290 41085 sw
rect 28126 41083 32290 41084
tri 32290 41083 32291 41084 sw
rect 28126 41082 32291 41083
tri 32291 41082 32292 41083 sw
rect 28126 41081 32292 41082
tri 32292 41081 32293 41082 sw
rect 28126 41080 32293 41081
tri 32293 41080 32294 41081 sw
rect 28126 41079 32294 41080
tri 32294 41079 32295 41080 sw
rect 28126 41078 32295 41079
tri 32295 41078 32296 41079 sw
rect 28126 41077 32296 41078
tri 32296 41077 32297 41078 sw
rect 28126 41076 32297 41077
tri 32297 41076 32298 41077 sw
rect 28126 41075 32298 41076
tri 32298 41075 32299 41076 sw
rect 28126 41074 32299 41075
tri 32299 41074 32300 41075 sw
rect 28126 41073 32300 41074
tri 32300 41073 32301 41074 sw
rect 28126 41072 32301 41073
tri 32301 41072 32302 41073 sw
rect 28126 41071 32302 41072
tri 32302 41071 32303 41072 sw
rect 28126 41070 32303 41071
tri 32303 41070 32304 41071 sw
rect 28126 41069 32304 41070
tri 32304 41069 32305 41070 sw
rect 28126 41068 32305 41069
tri 32305 41068 32306 41069 sw
rect 28126 41067 32306 41068
tri 32306 41067 32307 41068 sw
rect 28126 41066 32307 41067
tri 32307 41066 32308 41067 sw
rect 28126 41065 32308 41066
tri 32308 41065 32309 41066 sw
rect 28126 41064 32309 41065
tri 32309 41064 32310 41065 sw
rect 28126 41063 32310 41064
tri 32310 41063 32311 41064 sw
rect 28126 41062 32311 41063
tri 32311 41062 32312 41063 sw
rect 28126 41061 32312 41062
tri 32312 41061 32313 41062 sw
rect 28126 41060 32313 41061
tri 32313 41060 32314 41061 sw
rect 28126 41059 32314 41060
tri 32314 41059 32315 41060 sw
rect 28126 41058 32315 41059
tri 32315 41058 32316 41059 sw
rect 28126 41057 32316 41058
tri 32316 41057 32317 41058 sw
rect 28126 41056 32317 41057
tri 32317 41056 32318 41057 sw
rect 28126 41055 32318 41056
tri 32318 41055 32319 41056 sw
rect 28126 41054 32319 41055
tri 32319 41054 32320 41055 sw
rect 28126 41053 32320 41054
tri 32320 41053 32321 41054 sw
rect 28126 41052 32321 41053
tri 32321 41052 32322 41053 sw
rect 28126 41051 32322 41052
tri 32322 41051 32323 41052 sw
rect 28126 41050 32323 41051
tri 32323 41050 32324 41051 sw
rect 28126 41049 32324 41050
tri 32324 41049 32325 41050 sw
rect 28126 41048 32325 41049
tri 32325 41048 32326 41049 sw
rect 28126 41047 32326 41048
tri 32326 41047 32327 41048 sw
rect 28126 41046 32327 41047
tri 32327 41046 32328 41047 sw
rect 28126 41045 32328 41046
tri 32328 41045 32329 41046 sw
rect 28126 41044 32329 41045
tri 32329 41044 32330 41045 sw
rect 28126 41043 32330 41044
tri 32330 41043 32331 41044 sw
rect 28126 41042 32331 41043
tri 32331 41042 32332 41043 sw
rect 28126 41041 32332 41042
tri 32332 41041 32333 41042 sw
rect 28126 41040 32333 41041
tri 32333 41040 32334 41041 sw
rect 28126 41039 32334 41040
tri 32334 41039 32335 41040 sw
rect 28126 41038 32335 41039
tri 32335 41038 32336 41039 sw
rect 28126 41037 32336 41038
tri 32336 41037 32337 41038 sw
rect 28126 41036 32337 41037
tri 32337 41036 32338 41037 sw
rect 28126 41035 32338 41036
tri 32338 41035 32339 41036 sw
rect 28126 41034 32339 41035
tri 32339 41034 32340 41035 sw
rect 28126 41033 32340 41034
tri 32340 41033 32341 41034 sw
rect 28126 41032 32341 41033
tri 32341 41032 32342 41033 sw
rect 28126 41031 32342 41032
tri 32342 41031 32343 41032 sw
rect 28126 41030 32343 41031
tri 32343 41030 32344 41031 sw
rect 28126 41029 32344 41030
tri 32344 41029 32345 41030 sw
rect 28126 41028 32345 41029
tri 32345 41028 32346 41029 sw
rect 28126 41027 32346 41028
tri 32346 41027 32347 41028 sw
rect 28126 41026 32347 41027
tri 32347 41026 32348 41027 sw
rect 28126 41025 32348 41026
tri 32348 41025 32349 41026 sw
rect 28126 41024 32349 41025
tri 32349 41024 32350 41025 sw
rect 28126 41023 32350 41024
tri 32350 41023 32351 41024 sw
rect 28126 41022 32351 41023
tri 32351 41022 32352 41023 sw
rect 28126 41021 32352 41022
tri 32352 41021 32353 41022 sw
rect 28126 41020 32353 41021
tri 32353 41020 32354 41021 sw
rect 28126 41019 32354 41020
tri 32354 41019 32355 41020 sw
rect 28126 41018 32355 41019
tri 32355 41018 32356 41019 sw
rect 28126 41017 32356 41018
tri 32356 41017 32357 41018 sw
rect 28126 41016 32357 41017
tri 32357 41016 32358 41017 sw
rect 28126 41015 32358 41016
tri 32358 41015 32359 41016 sw
rect 28126 41014 32359 41015
tri 32359 41014 32360 41015 sw
rect 28126 41013 32360 41014
tri 32360 41013 32361 41014 sw
rect 28126 41012 32361 41013
tri 32361 41012 32362 41013 sw
rect 28126 41011 32362 41012
tri 32362 41011 32363 41012 sw
rect 28126 41010 32363 41011
tri 32363 41010 32364 41011 sw
rect 28126 41009 32364 41010
tri 32364 41009 32365 41010 sw
rect 28126 41008 32365 41009
tri 32365 41008 32366 41009 sw
rect 28126 41007 32366 41008
tri 32366 41007 32367 41008 sw
rect 28126 41006 32367 41007
tri 32367 41006 32368 41007 sw
rect 28126 41005 32368 41006
tri 32368 41005 32369 41006 sw
rect 28126 41004 32369 41005
tri 32369 41004 32370 41005 sw
rect 23776 40828 27844 41004
rect 22232 40536 23484 40828
tri 23484 40536 23776 40828 sw
tri 23776 40827 23777 40828 ne
rect 23777 40827 27844 40828
rect 22232 40535 23776 40536
tri 23776 40535 23777 40536 sw
tri 23777 40535 24069 40827 ne
rect 24069 40722 27844 40827
tri 27844 40722 28126 41004 sw
tri 28126 40937 28193 41004 ne
rect 28193 41003 32370 41004
tri 32370 41003 32371 41004 sw
rect 28193 41002 32371 41003
tri 32371 41002 32372 41003 sw
rect 28193 41001 32372 41002
tri 32372 41001 32373 41002 sw
rect 28193 41000 32373 41001
tri 32373 41000 32374 41001 sw
rect 28193 40999 32374 41000
tri 32374 40999 32375 41000 sw
rect 28193 40998 32375 40999
tri 32375 40998 32376 40999 sw
rect 28193 40997 32376 40998
tri 32376 40997 32377 40998 sw
rect 28193 40996 32377 40997
tri 32377 40996 32378 40997 sw
rect 28193 40995 32378 40996
tri 32378 40995 32379 40996 sw
rect 28193 40994 32379 40995
tri 32379 40994 32380 40995 sw
rect 28193 40993 32380 40994
tri 32380 40993 32381 40994 sw
rect 28193 40992 32381 40993
tri 32381 40992 32382 40993 sw
rect 28193 40991 32382 40992
tri 32382 40991 32383 40992 sw
rect 28193 40990 32383 40991
tri 32383 40990 32384 40991 sw
rect 28193 40989 32384 40990
tri 32384 40989 32385 40990 sw
rect 28193 40988 32385 40989
tri 32385 40988 32386 40989 sw
rect 28193 40987 32386 40988
tri 32386 40987 32387 40988 sw
rect 28193 40986 32387 40987
tri 32387 40986 32388 40987 sw
rect 28193 40985 32388 40986
tri 32388 40985 32389 40986 sw
rect 28193 40984 32389 40985
tri 32389 40984 32390 40985 sw
rect 28193 40983 32390 40984
tri 32390 40983 32391 40984 sw
rect 28193 40982 32391 40983
tri 32391 40982 32392 40983 sw
rect 28193 40981 32392 40982
tri 32392 40981 32393 40982 sw
rect 28193 40980 32393 40981
tri 32393 40980 32394 40981 sw
rect 28193 40979 32394 40980
tri 32394 40979 32395 40980 sw
rect 28193 40978 32395 40979
tri 32395 40978 32396 40979 sw
rect 28193 40977 32396 40978
tri 32396 40977 32397 40978 sw
rect 28193 40976 32397 40977
tri 32397 40976 32398 40977 sw
rect 28193 40975 32398 40976
tri 32398 40975 32399 40976 sw
rect 28193 40974 32399 40975
tri 32399 40974 32400 40975 sw
rect 28193 40973 32400 40974
tri 32400 40973 32401 40974 sw
rect 28193 40972 32401 40973
tri 32401 40972 32402 40973 sw
rect 28193 40971 32402 40972
tri 32402 40971 32403 40972 sw
rect 28193 40970 32403 40971
tri 32403 40970 32404 40971 sw
rect 28193 40969 32404 40970
tri 32404 40969 32405 40970 sw
rect 28193 40968 32405 40969
tri 32405 40968 32406 40969 sw
rect 28193 40967 32406 40968
tri 32406 40967 32407 40968 sw
rect 28193 40966 32407 40967
tri 32407 40966 32408 40967 sw
rect 28193 40965 32408 40966
tri 32408 40965 32409 40966 sw
rect 28193 40964 32409 40965
tri 32409 40964 32410 40965 sw
rect 28193 40963 32410 40964
tri 32410 40963 32411 40964 sw
rect 28193 40962 32411 40963
tri 32411 40962 32412 40963 sw
rect 28193 40961 32412 40962
tri 32412 40961 32413 40962 sw
rect 28193 40960 32413 40961
tri 32413 40960 32414 40961 sw
rect 28193 40959 32414 40960
tri 32414 40959 32415 40960 sw
rect 28193 40958 32415 40959
tri 32415 40958 32416 40959 sw
rect 28193 40957 32416 40958
tri 32416 40957 32417 40958 sw
rect 28193 40956 32417 40957
tri 32417 40956 32418 40957 sw
rect 28193 40955 32418 40956
tri 32418 40955 32419 40956 sw
rect 28193 40954 32419 40955
tri 32419 40954 32420 40955 sw
rect 28193 40953 32420 40954
tri 32420 40953 32421 40954 sw
rect 28193 40952 32421 40953
tri 32421 40952 32422 40953 sw
rect 28193 40951 32422 40952
tri 32422 40951 32423 40952 sw
rect 28193 40950 32423 40951
tri 32423 40950 32424 40951 sw
rect 28193 40949 32424 40950
tri 32424 40949 32425 40950 sw
rect 28193 40948 32425 40949
tri 32425 40948 32426 40949 sw
rect 28193 40947 32426 40948
tri 32426 40947 32427 40948 sw
rect 28193 40946 32427 40947
tri 32427 40946 32428 40947 sw
rect 28193 40945 32428 40946
tri 32428 40945 32429 40946 sw
rect 28193 40944 32429 40945
tri 32429 40944 32430 40945 sw
rect 28193 40943 32430 40944
tri 32430 40943 32431 40944 sw
rect 28193 40942 32431 40943
tri 32431 40942 32432 40943 sw
rect 28193 40941 32432 40942
tri 32432 40941 32433 40942 sw
rect 28193 40940 32433 40941
tri 32433 40940 32434 40941 sw
rect 28193 40939 32434 40940
tri 32434 40939 32435 40940 sw
rect 28193 40938 32435 40939
tri 32435 40938 32436 40939 sw
rect 28193 40937 32436 40938
tri 32436 40937 32437 40938 sw
rect 24069 40655 28126 40722
tri 28126 40655 28193 40722 sw
tri 28193 40655 28475 40937 ne
rect 28475 40936 32437 40937
tri 32437 40936 32438 40937 sw
rect 28475 40935 32438 40936
tri 32438 40935 32439 40936 sw
rect 28475 40934 32439 40935
tri 32439 40934 32440 40935 sw
rect 28475 40933 32440 40934
tri 32440 40933 32441 40934 sw
rect 28475 40932 32441 40933
tri 32441 40932 32442 40933 sw
rect 28475 40931 32442 40932
tri 32442 40931 32443 40932 sw
rect 28475 40930 32443 40931
tri 32443 40930 32444 40931 sw
rect 28475 40929 32444 40930
tri 32444 40929 32445 40930 sw
rect 28475 40928 32445 40929
tri 32445 40928 32446 40929 sw
rect 28475 40927 32446 40928
tri 32446 40927 32447 40928 sw
rect 28475 40926 32447 40927
tri 32447 40926 32448 40927 sw
rect 28475 40925 32448 40926
tri 32448 40925 32449 40926 sw
rect 28475 40924 32449 40925
tri 32449 40924 32450 40925 sw
rect 28475 40923 32450 40924
tri 32450 40923 32451 40924 sw
rect 28475 40922 32451 40923
tri 32451 40922 32452 40923 sw
rect 28475 40921 32452 40922
tri 32452 40921 32453 40922 sw
rect 28475 40920 32453 40921
tri 32453 40920 32454 40921 sw
rect 28475 40919 32454 40920
tri 32454 40919 32455 40920 sw
rect 28475 40918 32455 40919
tri 32455 40918 32456 40919 sw
rect 28475 40917 32456 40918
tri 32456 40917 32457 40918 sw
rect 28475 40916 32457 40917
tri 32457 40916 32458 40917 sw
rect 28475 40915 32458 40916
tri 32458 40915 32459 40916 sw
rect 28475 40914 32459 40915
tri 32459 40914 32460 40915 sw
rect 28475 40913 32460 40914
tri 32460 40913 32461 40914 sw
rect 28475 40912 32461 40913
tri 32461 40912 32462 40913 sw
rect 28475 40911 32462 40912
tri 32462 40911 32463 40912 sw
rect 28475 40910 32463 40911
tri 32463 40910 32464 40911 sw
rect 28475 40909 32464 40910
tri 32464 40909 32465 40910 sw
rect 28475 40908 32465 40909
tri 32465 40908 32466 40909 sw
rect 28475 40907 32466 40908
tri 32466 40907 32467 40908 sw
rect 28475 40906 32467 40907
tri 32467 40906 32468 40907 sw
rect 28475 40905 32468 40906
tri 32468 40905 32469 40906 sw
rect 28475 40904 32469 40905
tri 32469 40904 32470 40905 sw
rect 28475 40903 32470 40904
tri 32470 40903 32471 40904 sw
rect 28475 40902 32471 40903
tri 32471 40902 32472 40903 sw
rect 28475 40901 32472 40902
tri 32472 40901 32473 40902 sw
rect 28475 40900 32473 40901
tri 32473 40900 32474 40901 sw
rect 28475 40899 32474 40900
tri 32474 40899 32475 40900 sw
rect 28475 40898 32475 40899
tri 32475 40898 32476 40899 sw
rect 28475 40897 32476 40898
tri 32476 40897 32477 40898 sw
rect 28475 40896 32477 40897
tri 32477 40896 32478 40897 sw
rect 28475 40895 32478 40896
tri 32478 40895 32479 40896 sw
rect 28475 40894 32479 40895
tri 32479 40894 32480 40895 sw
rect 28475 40893 32480 40894
tri 32480 40893 32481 40894 sw
rect 28475 40892 32481 40893
tri 32481 40892 32482 40893 sw
rect 28475 40891 32482 40892
tri 32482 40891 32483 40892 sw
rect 28475 40890 32483 40891
tri 32483 40890 32484 40891 sw
rect 28475 40889 32484 40890
tri 32484 40889 32485 40890 sw
rect 28475 40888 32485 40889
tri 32485 40888 32486 40889 sw
rect 28475 40887 32486 40888
tri 32486 40887 32487 40888 sw
rect 28475 40886 32487 40887
tri 32487 40886 32488 40887 sw
rect 28475 40885 32488 40886
tri 32488 40885 32489 40886 sw
rect 28475 40884 32489 40885
tri 32489 40884 32490 40885 sw
rect 28475 40883 32490 40884
tri 32490 40883 32491 40884 sw
rect 28475 40882 32491 40883
tri 32491 40882 32492 40883 sw
rect 28475 40881 32492 40882
tri 32492 40881 32493 40882 sw
rect 28475 40880 32493 40881
tri 32493 40880 32494 40881 sw
rect 28475 40879 32494 40880
tri 32494 40879 32495 40880 sw
rect 28475 40878 32495 40879
tri 32495 40878 32496 40879 sw
rect 28475 40877 32496 40878
tri 32496 40877 32497 40878 sw
rect 28475 40876 32497 40877
tri 32497 40876 32498 40877 sw
rect 28475 40875 32498 40876
tri 32498 40875 32499 40876 sw
rect 28475 40874 32499 40875
tri 32499 40874 32500 40875 sw
rect 28475 40873 32500 40874
tri 32500 40873 32501 40874 sw
rect 28475 40872 32501 40873
tri 32501 40872 32502 40873 sw
rect 28475 40871 32502 40872
tri 32502 40871 32503 40872 sw
rect 28475 40870 32503 40871
tri 32503 40870 32504 40871 sw
rect 28475 40869 32504 40870
tri 32504 40869 32505 40870 sw
rect 28475 40868 32505 40869
tri 32505 40868 32506 40869 sw
rect 28475 40867 32506 40868
tri 32506 40867 32507 40868 sw
rect 28475 40866 32507 40867
tri 32507 40866 32508 40867 sw
rect 28475 40865 32508 40866
tri 32508 40865 32509 40866 sw
rect 28475 40864 32509 40865
tri 32509 40864 32510 40865 sw
rect 28475 40863 32510 40864
tri 32510 40863 32511 40864 sw
rect 28475 40862 32511 40863
tri 32511 40862 32512 40863 sw
rect 28475 40861 32512 40862
tri 32512 40861 32513 40862 sw
rect 28475 40860 32513 40861
tri 32513 40860 32514 40861 sw
rect 28475 40859 32514 40860
tri 32514 40859 32515 40860 sw
rect 28475 40858 32515 40859
tri 32515 40858 32516 40859 sw
rect 28475 40857 32516 40858
tri 32516 40857 32517 40858 sw
rect 28475 40856 32517 40857
tri 32517 40856 32518 40857 sw
rect 28475 40855 32518 40856
tri 32518 40855 32519 40856 sw
rect 28475 40854 32519 40855
tri 32519 40854 32520 40855 sw
rect 28475 40853 32520 40854
tri 32520 40853 32521 40854 sw
rect 28475 40852 32521 40853
tri 32521 40852 32522 40853 sw
rect 28475 40851 32522 40852
tri 32522 40851 32523 40852 sw
rect 28475 40850 32523 40851
tri 32523 40850 32524 40851 sw
rect 28475 40849 32524 40850
tri 32524 40849 32525 40850 sw
rect 28475 40848 32525 40849
tri 32525 40848 32526 40849 sw
rect 28475 40847 32526 40848
tri 32526 40847 32527 40848 sw
rect 28475 40846 32527 40847
tri 32527 40846 32528 40847 sw
rect 28475 40845 32528 40846
tri 32528 40845 32529 40846 sw
rect 28475 40844 32529 40845
tri 32529 40844 32530 40845 sw
rect 28475 40843 32530 40844
tri 32530 40843 32531 40844 sw
rect 28475 40842 32531 40843
tri 32531 40842 32532 40843 sw
rect 28475 40841 32532 40842
tri 32532 40841 32533 40842 sw
tri 32533 40841 32830 41138 ne
rect 32830 41129 34237 41138
tri 34237 41129 34522 41414 sw
tri 34526 41129 34811 41414 ne
rect 34811 41130 36506 41414
tri 36506 41130 36790 41414 sw
tri 36796 41130 37080 41414 ne
rect 37080 41192 40968 41414
tri 40968 41192 41262 41486 sw
tri 41262 41287 41461 41486 ne
rect 41461 41400 45304 41486
tri 45304 41400 45592 41688 sw
tri 45592 41400 45880 41688 ne
rect 45880 41486 49836 41688
tri 49836 41486 50038 41688 sw
tri 50038 41486 50335 41783 ne
rect 50335 41780 54211 41783
tri 54211 41780 54285 41854 sw
tri 54285 41780 54578 42073 ne
rect 54578 42016 56030 42073
tri 56030 42016 56322 42308 sw
tri 56322 42016 56614 42308 ne
rect 56614 42016 70613 42308
rect 54578 41780 56322 42016
rect 50335 41487 54285 41780
tri 54285 41487 54578 41780 sw
tri 54578 41779 54579 41780 ne
rect 54579 41779 56322 41780
rect 50335 41486 54578 41487
tri 54578 41486 54579 41487 sw
tri 54579 41486 54872 41779 ne
rect 54872 41778 56322 41779
tri 56322 41778 56560 42016 sw
tri 56614 41778 56852 42016 ne
rect 56852 41778 70613 42016
rect 54872 41486 56560 41778
tri 56560 41486 56852 41778 sw
tri 56852 41486 57144 41778 ne
rect 57144 41486 70613 41778
rect 45880 41400 50038 41486
rect 41461 41287 45592 41400
rect 37080 41130 41262 41192
rect 34811 41129 36790 41130
rect 32830 40841 34522 41129
rect 28475 40655 32533 40841
rect 24069 40535 28193 40655
rect 22232 40243 23777 40535
tri 23777 40243 24069 40535 sw
tri 24069 40534 24070 40535 ne
rect 24070 40534 28193 40535
rect 22232 40242 24069 40243
tri 24069 40242 24070 40243 sw
tri 24070 40242 24362 40534 ne
rect 24362 40373 28193 40534
tri 28193 40373 28475 40655 sw
tri 28475 40654 28476 40655 ne
rect 28476 40654 32533 40655
rect 24362 40372 28475 40373
tri 28475 40372 28476 40373 sw
tri 28476 40372 28758 40654 ne
rect 28758 40544 32533 40654
tri 32533 40544 32830 40841 sw
tri 32830 40840 32831 40841 ne
rect 32831 40840 34522 40841
tri 34522 40840 34811 41129 sw
tri 34811 40840 35100 41129 ne
rect 35100 40840 36790 41129
tri 36790 40840 37080 41130 sw
tri 37080 40840 37370 41130 ne
rect 37370 40993 41262 41130
tri 41262 40993 41461 41192 sw
tri 41461 41135 41613 41287 ne
rect 41613 41135 45592 41287
rect 37370 40841 41461 40993
tri 41461 40841 41613 40993 sw
tri 41613 40841 41907 41135 ne
rect 41907 41112 45592 41135
tri 45592 41112 45880 41400 sw
tri 45880 41129 46151 41400 ne
rect 46151 41189 50038 41400
tri 50038 41189 50335 41486 sw
tri 50335 41287 50534 41486 ne
rect 50534 41287 54579 41486
rect 46151 41129 50335 41189
rect 41907 40841 45880 41112
tri 45880 40841 46151 41112 sw
tri 46151 40841 46439 41129 ne
rect 46439 40990 50335 41129
tri 50335 40990 50534 41189 sw
tri 50534 41138 50683 41287 ne
rect 50683 41193 54579 41287
tri 54579 41193 54872 41486 sw
tri 54872 41287 55071 41486 ne
rect 55071 41414 56852 41486
tri 56852 41414 56924 41486 sw
tri 57144 41414 57216 41486 ne
rect 57216 41414 70613 41486
rect 55071 41287 56924 41414
tri 56924 41287 57051 41414 sw
tri 57216 41287 57343 41414 ne
rect 57343 41297 70613 41414
rect 70669 41297 71000 42497
rect 57343 41287 71000 41297
rect 50683 41138 54872 41193
rect 46439 40841 50534 40990
tri 50534 40841 50683 40990 sw
tri 50683 40841 50980 41138 ne
rect 50980 40994 54872 41138
tri 54872 40994 55071 41193 sw
tri 55071 41000 55358 41287 ne
rect 55358 41200 57051 41287
tri 57051 41200 57138 41287 sw
tri 57343 41200 57430 41287 ne
rect 57430 41200 71000 41287
rect 55358 41000 57138 41200
tri 57138 41000 57338 41200 sw
rect 50980 40841 55071 40994
rect 37370 40840 41613 40841
rect 28758 40543 32830 40544
tri 32830 40543 32831 40544 sw
tri 32831 40543 33128 40840 ne
rect 33128 40749 34811 40840
tri 34811 40749 34902 40840 sw
tri 35100 40749 35191 40840 ne
rect 35191 40750 37080 40840
tri 37080 40750 37170 40840 sw
tri 37370 40750 37460 40840 ne
rect 37460 40750 41613 40840
rect 35191 40749 37170 40750
rect 33128 40543 34902 40749
rect 28758 40372 32831 40543
rect 24362 40242 28476 40372
rect 22232 39950 24070 40242
tri 24070 39950 24362 40242 sw
tri 24362 40221 24383 40242 ne
rect 24383 40221 28476 40242
rect 22232 39929 24362 39950
tri 24362 39929 24383 39950 sw
tri 24383 39929 24675 40221 ne
rect 24675 40090 28476 40221
tri 28476 40090 28758 40372 sw
tri 28758 40371 28759 40372 ne
rect 28759 40371 32831 40372
rect 24675 40089 28758 40090
tri 28758 40089 28759 40090 sw
tri 28759 40089 29041 40371 ne
rect 29041 40246 32831 40371
tri 32831 40246 33128 40543 sw
tri 33128 40371 33300 40543 ne
rect 33300 40460 34902 40543
tri 34902 40460 35191 40749 sw
tri 35191 40460 35480 40749 ne
rect 35480 40460 37170 40749
tri 37170 40460 37460 40750 sw
tri 37460 40460 37750 40750 ne
rect 37750 40547 41613 40750
tri 41613 40547 41907 40841 sw
tri 41907 40755 41993 40841 ne
rect 41993 40755 46151 40841
rect 37750 40461 41907 40547
tri 41907 40461 41993 40547 sw
tri 41993 40461 42287 40755 ne
rect 42287 40553 46151 40755
tri 46151 40553 46439 40841 sw
tri 46439 40749 46531 40841 ne
rect 46531 40749 50683 40841
rect 42287 40461 46439 40553
tri 46439 40461 46531 40553 sw
tri 46531 40461 46819 40749 ne
rect 46819 40544 50683 40749
tri 50683 40544 50980 40841 sw
tri 50980 40644 51177 40841 ne
rect 51177 40707 55071 40841
tri 55071 40707 55358 40994 sw
tri 55358 40840 55518 41000 ne
rect 55518 40840 71000 41000
rect 51177 40644 55358 40707
rect 46819 40461 50980 40544
rect 37750 40460 41993 40461
rect 33300 40371 35191 40460
rect 29041 40089 33128 40246
rect 24675 39929 28759 40089
rect 22232 39637 24383 39929
tri 24383 39637 24675 39929 sw
tri 24675 39756 24848 39929 ne
rect 24848 39807 28759 39929
tri 28759 39807 29041 40089 sw
tri 29041 40087 29043 40089 ne
rect 29043 40087 33128 40089
rect 24848 39805 29041 39807
tri 29041 39805 29043 39807 sw
tri 29043 39805 29325 40087 ne
rect 29325 40074 33128 40087
tri 33128 40074 33300 40246 sw
tri 33300 40074 33597 40371 ne
rect 33597 40171 35191 40371
tri 35191 40171 35480 40460 sw
tri 35480 40171 35769 40460 ne
rect 35769 40371 37460 40460
tri 37460 40371 37549 40460 sw
tri 37750 40371 37839 40460 ne
rect 37839 40371 41993 40460
rect 35769 40171 37549 40371
rect 33597 40074 35480 40171
rect 29325 39805 33300 40074
rect 24848 39756 29043 39805
rect 22232 39464 24675 39637
tri 24675 39464 24848 39637 sw
tri 24848 39635 24969 39756 ne
rect 24969 39635 29043 39756
tri 24969 39464 25140 39635 ne
rect 25140 39523 29043 39635
tri 29043 39523 29325 39805 sw
tri 29325 39625 29505 39805 ne
rect 29505 39777 33300 39805
tri 33300 39777 33597 40074 sw
tri 33597 39937 33734 40074 ne
rect 33734 39937 35480 40074
rect 29505 39640 33597 39777
tri 33597 39640 33734 39777 sw
tri 33734 39640 34031 39937 ne
rect 34031 39882 35480 39937
tri 35480 39882 35769 40171 sw
tri 35769 39882 36058 40171 ne
rect 36058 40081 37549 40171
tri 37549 40081 37839 40371 sw
tri 37839 40081 38129 40371 ne
rect 38129 40167 41993 40371
tri 41993 40167 42287 40461 sw
tri 42287 40371 42377 40461 ne
rect 42377 40371 46531 40461
rect 38129 40081 42287 40167
rect 36058 39923 37839 40081
tri 37839 39923 37997 40081 sw
tri 38129 39923 38287 40081 ne
rect 38287 40077 42287 40081
tri 42287 40077 42377 40167 sw
tri 42377 40077 42671 40371 ne
rect 42671 40173 46531 40371
tri 46531 40173 46819 40461 sw
tri 46819 40371 46909 40461 ne
rect 46909 40371 50980 40461
rect 42671 40083 46819 40173
tri 46819 40083 46909 40173 sw
tri 46909 40153 47127 40371 ne
rect 47127 40347 50980 40371
tri 50980 40347 51177 40544 sw
tri 51177 40347 51474 40644 ne
rect 51474 40547 55358 40644
tri 55358 40547 55518 40707 sw
tri 55518 40706 55652 40840 ne
rect 55652 40706 71000 40840
rect 51474 40546 55518 40547
tri 55518 40546 55519 40547 sw
rect 51474 40545 55519 40546
tri 55519 40545 55520 40546 sw
rect 51474 40544 55520 40545
tri 55520 40544 55521 40545 sw
rect 51474 40543 55521 40544
tri 55521 40543 55522 40544 sw
rect 51474 40542 55522 40543
tri 55522 40542 55523 40543 sw
rect 51474 40541 55523 40542
tri 55523 40541 55524 40542 sw
rect 51474 40540 55524 40541
tri 55524 40540 55525 40541 sw
rect 51474 40539 55525 40540
tri 55525 40539 55526 40540 sw
rect 51474 40538 55526 40539
tri 55526 40538 55527 40539 sw
rect 51474 40537 55527 40538
tri 55527 40537 55528 40538 sw
rect 51474 40536 55528 40537
tri 55528 40536 55529 40537 sw
rect 51474 40535 55529 40536
tri 55529 40535 55530 40536 sw
rect 51474 40534 55530 40535
tri 55530 40534 55531 40535 sw
rect 51474 40533 55531 40534
tri 55531 40533 55532 40534 sw
rect 51474 40532 55532 40533
tri 55532 40532 55533 40533 sw
rect 51474 40531 55533 40532
tri 55533 40531 55534 40532 sw
rect 51474 40530 55534 40531
tri 55534 40530 55535 40531 sw
rect 51474 40529 55535 40530
tri 55535 40529 55536 40530 sw
rect 51474 40528 55536 40529
tri 55536 40528 55537 40529 sw
rect 51474 40527 55537 40528
tri 55537 40527 55538 40528 sw
rect 51474 40526 55538 40527
tri 55538 40526 55539 40527 sw
rect 51474 40525 55539 40526
tri 55539 40525 55540 40526 sw
rect 51474 40524 55540 40525
tri 55540 40524 55541 40525 sw
rect 51474 40523 55541 40524
tri 55541 40523 55542 40524 sw
rect 51474 40522 55542 40523
tri 55542 40522 55543 40523 sw
rect 51474 40521 55543 40522
tri 55543 40521 55544 40522 sw
rect 51474 40520 55544 40521
tri 55544 40520 55545 40521 sw
rect 51474 40519 55545 40520
tri 55545 40519 55546 40520 sw
rect 51474 40518 55546 40519
tri 55546 40518 55547 40519 sw
rect 51474 40517 55547 40518
tri 55547 40517 55548 40518 sw
rect 51474 40516 55548 40517
tri 55548 40516 55549 40517 sw
rect 51474 40515 55549 40516
tri 55549 40515 55550 40516 sw
rect 51474 40514 55550 40515
tri 55550 40514 55551 40515 sw
rect 51474 40513 55551 40514
tri 55551 40513 55552 40514 sw
rect 51474 40512 55552 40513
tri 55552 40512 55553 40513 sw
rect 51474 40511 55553 40512
tri 55553 40511 55554 40512 sw
rect 51474 40510 55554 40511
tri 55554 40510 55555 40511 sw
rect 51474 40509 55555 40510
tri 55555 40509 55556 40510 sw
rect 51474 40508 55556 40509
tri 55556 40508 55557 40509 sw
rect 51474 40507 55557 40508
tri 55557 40507 55558 40508 sw
rect 51474 40506 55558 40507
tri 55558 40506 55559 40507 sw
rect 51474 40505 55559 40506
tri 55559 40505 55560 40506 sw
rect 51474 40504 55560 40505
tri 55560 40504 55561 40505 sw
rect 51474 40503 55561 40504
tri 55561 40503 55562 40504 sw
rect 51474 40502 55562 40503
tri 55562 40502 55563 40503 sw
rect 51474 40501 55563 40502
tri 55563 40501 55564 40502 sw
rect 51474 40500 55564 40501
tri 55564 40500 55565 40501 sw
rect 51474 40499 55565 40500
tri 55565 40499 55566 40500 sw
rect 51474 40498 55566 40499
tri 55566 40498 55567 40499 sw
rect 51474 40497 55567 40498
tri 55567 40497 55568 40498 sw
rect 51474 40496 55568 40497
tri 55568 40496 55569 40497 sw
rect 51474 40495 55569 40496
tri 55569 40495 55570 40496 sw
rect 51474 40494 55570 40495
tri 55570 40494 55571 40495 sw
rect 51474 40493 55571 40494
tri 55571 40493 55572 40494 sw
rect 51474 40492 55572 40493
tri 55572 40492 55573 40493 sw
rect 51474 40491 55573 40492
tri 55573 40491 55574 40492 sw
rect 51474 40490 55574 40491
tri 55574 40490 55575 40491 sw
rect 51474 40489 55575 40490
tri 55575 40489 55576 40490 sw
rect 51474 40488 55576 40489
tri 55576 40488 55577 40489 sw
rect 51474 40487 55577 40488
tri 55577 40487 55578 40488 sw
rect 51474 40486 55578 40487
tri 55578 40486 55579 40487 sw
rect 51474 40485 55579 40486
tri 55579 40485 55580 40486 sw
rect 51474 40484 55580 40485
tri 55580 40484 55581 40485 sw
rect 51474 40483 55581 40484
tri 55581 40483 55582 40484 sw
rect 51474 40482 55582 40483
tri 55582 40482 55583 40483 sw
rect 51474 40481 55583 40482
tri 55583 40481 55584 40482 sw
rect 51474 40480 55584 40481
tri 55584 40480 55585 40481 sw
rect 51474 40479 55585 40480
tri 55585 40479 55586 40480 sw
rect 51474 40478 55586 40479
tri 55586 40478 55587 40479 sw
rect 51474 40477 55587 40478
tri 55587 40477 55588 40478 sw
rect 51474 40476 55588 40477
tri 55588 40476 55589 40477 sw
rect 51474 40475 55589 40476
tri 55589 40475 55590 40476 sw
rect 51474 40474 55590 40475
tri 55590 40474 55591 40475 sw
rect 51474 40473 55591 40474
tri 55591 40473 55592 40474 sw
rect 51474 40472 55592 40473
tri 55592 40472 55593 40473 sw
rect 51474 40471 55593 40472
tri 55593 40471 55594 40472 sw
rect 51474 40470 55594 40471
tri 55594 40470 55595 40471 sw
rect 51474 40469 55595 40470
tri 55595 40469 55596 40470 sw
rect 51474 40468 55596 40469
tri 55596 40468 55597 40469 sw
rect 51474 40467 55597 40468
tri 55597 40467 55598 40468 sw
rect 51474 40466 55598 40467
tri 55598 40466 55599 40467 sw
rect 51474 40465 55599 40466
tri 55599 40465 55600 40466 sw
rect 51474 40464 55600 40465
tri 55600 40464 55601 40465 sw
rect 51474 40463 55601 40464
tri 55601 40463 55602 40464 sw
rect 51474 40462 55602 40463
tri 55602 40462 55603 40463 sw
rect 51474 40461 55603 40462
tri 55603 40461 55604 40462 sw
rect 51474 40460 55604 40461
tri 55604 40460 55605 40461 sw
rect 51474 40459 55605 40460
tri 55605 40459 55606 40460 sw
rect 51474 40458 55606 40459
tri 55606 40458 55607 40459 sw
rect 51474 40457 55607 40458
tri 55607 40457 55608 40458 sw
rect 51474 40456 55608 40457
tri 55608 40456 55609 40457 sw
rect 51474 40455 55609 40456
tri 55609 40455 55610 40456 sw
rect 51474 40454 55610 40455
tri 55610 40454 55611 40455 sw
rect 51474 40453 55611 40454
tri 55611 40453 55612 40454 sw
rect 51474 40452 55612 40453
tri 55612 40452 55613 40453 sw
rect 51474 40451 55613 40452
tri 55613 40451 55614 40452 sw
rect 51474 40450 55614 40451
tri 55614 40450 55615 40451 sw
rect 51474 40449 55615 40450
tri 55615 40449 55616 40450 sw
rect 51474 40448 55616 40449
tri 55616 40448 55617 40449 sw
rect 51474 40447 55617 40448
tri 55617 40447 55618 40448 sw
rect 51474 40446 55618 40447
tri 55618 40446 55619 40447 sw
rect 51474 40445 55619 40446
tri 55619 40445 55620 40446 sw
rect 51474 40444 55620 40445
tri 55620 40444 55621 40445 sw
rect 51474 40443 55621 40444
tri 55621 40443 55622 40444 sw
tri 55652 40443 55915 40706 ne
rect 55915 40443 71000 40706
rect 51474 40347 55622 40443
rect 47127 40153 51177 40347
rect 42671 40077 46909 40083
rect 38287 39923 42377 40077
rect 36058 39882 37997 39923
rect 34031 39640 35769 39882
rect 29505 39639 33734 39640
tri 33734 39639 33735 39640 sw
rect 29505 39638 33735 39639
tri 33735 39638 33736 39639 sw
rect 29505 39637 33736 39638
tri 33736 39637 33737 39638 sw
rect 29505 39636 33737 39637
tri 33737 39636 33738 39637 sw
rect 29505 39635 33738 39636
tri 33738 39635 33739 39636 sw
rect 29505 39634 33739 39635
tri 33739 39634 33740 39635 sw
rect 29505 39633 33740 39634
tri 33740 39633 33741 39634 sw
rect 29505 39632 33741 39633
tri 33741 39632 33742 39633 sw
rect 29505 39631 33742 39632
tri 33742 39631 33743 39632 sw
rect 29505 39630 33743 39631
tri 33743 39630 33744 39631 sw
rect 29505 39629 33744 39630
tri 33744 39629 33745 39630 sw
rect 29505 39628 33745 39629
tri 33745 39628 33746 39629 sw
rect 29505 39627 33746 39628
tri 33746 39627 33747 39628 sw
rect 29505 39626 33747 39627
tri 33747 39626 33748 39627 sw
rect 29505 39625 33748 39626
tri 33748 39625 33749 39626 sw
rect 25140 39464 29325 39523
rect 22232 39172 24848 39464
tri 24848 39172 25140 39464 sw
tri 25140 39341 25263 39464 ne
rect 25263 39343 29325 39464
tri 29325 39343 29505 39523 sw
tri 29505 39343 29787 39625 ne
rect 29787 39624 33749 39625
tri 33749 39624 33750 39625 sw
rect 29787 39623 33750 39624
tri 33750 39623 33751 39624 sw
rect 29787 39622 33751 39623
tri 33751 39622 33752 39623 sw
rect 29787 39621 33752 39622
tri 33752 39621 33753 39622 sw
rect 29787 39620 33753 39621
tri 33753 39620 33754 39621 sw
rect 29787 39619 33754 39620
tri 33754 39619 33755 39620 sw
rect 29787 39618 33755 39619
tri 33755 39618 33756 39619 sw
rect 29787 39617 33756 39618
tri 33756 39617 33757 39618 sw
rect 29787 39616 33757 39617
tri 33757 39616 33758 39617 sw
rect 29787 39615 33758 39616
tri 33758 39615 33759 39616 sw
rect 29787 39614 33759 39615
tri 33759 39614 33760 39615 sw
rect 29787 39613 33760 39614
tri 33760 39613 33761 39614 sw
rect 29787 39612 33761 39613
tri 33761 39612 33762 39613 sw
rect 29787 39611 33762 39612
tri 33762 39611 33763 39612 sw
rect 29787 39610 33763 39611
tri 33763 39610 33764 39611 sw
rect 29787 39609 33764 39610
tri 33764 39609 33765 39610 sw
rect 29787 39608 33765 39609
tri 33765 39608 33766 39609 sw
rect 29787 39607 33766 39608
tri 33766 39607 33767 39608 sw
rect 29787 39606 33767 39607
tri 33767 39606 33768 39607 sw
rect 29787 39605 33768 39606
tri 33768 39605 33769 39606 sw
rect 29787 39604 33769 39605
tri 33769 39604 33770 39605 sw
rect 29787 39603 33770 39604
tri 33770 39603 33771 39604 sw
rect 29787 39602 33771 39603
tri 33771 39602 33772 39603 sw
rect 29787 39601 33772 39602
tri 33772 39601 33773 39602 sw
rect 29787 39600 33773 39601
tri 33773 39600 33774 39601 sw
rect 29787 39599 33774 39600
tri 33774 39599 33775 39600 sw
rect 29787 39598 33775 39599
tri 33775 39598 33776 39599 sw
rect 29787 39597 33776 39598
tri 33776 39597 33777 39598 sw
rect 29787 39596 33777 39597
tri 33777 39596 33778 39597 sw
rect 29787 39595 33778 39596
tri 33778 39595 33779 39596 sw
rect 29787 39594 33779 39595
tri 33779 39594 33780 39595 sw
rect 29787 39593 33780 39594
tri 33780 39593 33781 39594 sw
rect 29787 39592 33781 39593
tri 33781 39592 33782 39593 sw
rect 29787 39591 33782 39592
tri 33782 39591 33783 39592 sw
rect 29787 39590 33783 39591
tri 33783 39590 33784 39591 sw
rect 29787 39589 33784 39590
tri 33784 39589 33785 39590 sw
rect 29787 39588 33785 39589
tri 33785 39588 33786 39589 sw
rect 29787 39587 33786 39588
tri 33786 39587 33787 39588 sw
rect 29787 39586 33787 39587
tri 33787 39586 33788 39587 sw
rect 29787 39585 33788 39586
tri 33788 39585 33789 39586 sw
rect 29787 39584 33789 39585
tri 33789 39584 33790 39585 sw
rect 29787 39583 33790 39584
tri 33790 39583 33791 39584 sw
rect 29787 39582 33791 39583
tri 33791 39582 33792 39583 sw
rect 29787 39581 33792 39582
tri 33792 39581 33793 39582 sw
rect 29787 39580 33793 39581
tri 33793 39580 33794 39581 sw
rect 29787 39579 33794 39580
tri 33794 39579 33795 39580 sw
rect 29787 39578 33795 39579
tri 33795 39578 33796 39579 sw
rect 29787 39577 33796 39578
tri 33796 39577 33797 39578 sw
rect 29787 39576 33797 39577
tri 33797 39576 33798 39577 sw
rect 29787 39575 33798 39576
tri 33798 39575 33799 39576 sw
rect 29787 39574 33799 39575
tri 33799 39574 33800 39575 sw
rect 29787 39573 33800 39574
tri 33800 39573 33801 39574 sw
rect 29787 39572 33801 39573
tri 33801 39572 33802 39573 sw
rect 29787 39571 33802 39572
tri 33802 39571 33803 39572 sw
rect 29787 39570 33803 39571
tri 33803 39570 33804 39571 sw
rect 29787 39569 33804 39570
tri 33804 39569 33805 39570 sw
rect 29787 39568 33805 39569
tri 33805 39568 33806 39569 sw
rect 29787 39567 33806 39568
tri 33806 39567 33807 39568 sw
rect 29787 39566 33807 39567
tri 33807 39566 33808 39567 sw
rect 29787 39565 33808 39566
tri 33808 39565 33809 39566 sw
rect 29787 39564 33809 39565
tri 33809 39564 33810 39565 sw
rect 29787 39563 33810 39564
tri 33810 39563 33811 39564 sw
rect 29787 39562 33811 39563
tri 33811 39562 33812 39563 sw
rect 29787 39561 33812 39562
tri 33812 39561 33813 39562 sw
rect 29787 39560 33813 39561
tri 33813 39560 33814 39561 sw
rect 29787 39559 33814 39560
tri 33814 39559 33815 39560 sw
rect 29787 39558 33815 39559
tri 33815 39558 33816 39559 sw
rect 29787 39557 33816 39558
tri 33816 39557 33817 39558 sw
rect 29787 39556 33817 39557
tri 33817 39556 33818 39557 sw
rect 29787 39555 33818 39556
tri 33818 39555 33819 39556 sw
rect 29787 39554 33819 39555
tri 33819 39554 33820 39555 sw
rect 29787 39553 33820 39554
tri 33820 39553 33821 39554 sw
rect 29787 39552 33821 39553
tri 33821 39552 33822 39553 sw
rect 29787 39551 33822 39552
tri 33822 39551 33823 39552 sw
rect 29787 39550 33823 39551
tri 33823 39550 33824 39551 sw
rect 29787 39549 33824 39550
tri 33824 39549 33825 39550 sw
rect 29787 39548 33825 39549
tri 33825 39548 33826 39549 sw
rect 29787 39547 33826 39548
tri 33826 39547 33827 39548 sw
rect 29787 39546 33827 39547
tri 33827 39546 33828 39547 sw
rect 29787 39545 33828 39546
tri 33828 39545 33829 39546 sw
rect 29787 39544 33829 39545
tri 33829 39544 33830 39545 sw
rect 29787 39543 33830 39544
tri 33830 39543 33831 39544 sw
rect 29787 39542 33831 39543
tri 33831 39542 33832 39543 sw
rect 29787 39541 33832 39542
tri 33832 39541 33833 39542 sw
rect 29787 39540 33833 39541
tri 33833 39540 33834 39541 sw
rect 29787 39539 33834 39540
tri 33834 39539 33835 39540 sw
rect 29787 39538 33835 39539
tri 33835 39538 33836 39539 sw
rect 29787 39537 33836 39538
tri 33836 39537 33837 39538 sw
rect 29787 39536 33837 39537
tri 33837 39536 33838 39537 sw
rect 29787 39535 33838 39536
tri 33838 39535 33839 39536 sw
rect 29787 39534 33839 39535
tri 33839 39534 33840 39535 sw
rect 29787 39533 33840 39534
tri 33840 39533 33841 39534 sw
rect 29787 39532 33841 39533
tri 33841 39532 33842 39533 sw
rect 29787 39531 33842 39532
tri 33842 39531 33843 39532 sw
rect 29787 39530 33843 39531
tri 33843 39530 33844 39531 sw
rect 29787 39529 33844 39530
tri 33844 39529 33845 39530 sw
rect 29787 39528 33845 39529
tri 33845 39528 33846 39529 sw
rect 29787 39527 33846 39528
tri 33846 39527 33847 39528 sw
rect 29787 39526 33847 39527
tri 33847 39526 33848 39527 sw
rect 29787 39525 33848 39526
tri 33848 39525 33849 39526 sw
rect 29787 39524 33849 39525
tri 33849 39524 33850 39525 sw
rect 29787 39523 33850 39524
tri 33850 39523 33851 39524 sw
rect 29787 39522 33851 39523
tri 33851 39522 33852 39523 sw
rect 29787 39521 33852 39522
tri 33852 39521 33853 39522 sw
rect 29787 39520 33853 39521
tri 33853 39520 33854 39521 sw
rect 29787 39519 33854 39520
tri 33854 39519 33855 39520 sw
rect 29787 39518 33855 39519
tri 33855 39518 33856 39519 sw
rect 29787 39517 33856 39518
tri 33856 39517 33857 39518 sw
rect 29787 39516 33857 39517
tri 33857 39516 33858 39517 sw
rect 29787 39515 33858 39516
tri 33858 39515 33859 39516 sw
rect 29787 39514 33859 39515
tri 33859 39514 33860 39515 sw
rect 29787 39513 33860 39514
tri 33860 39513 33861 39514 sw
rect 29787 39512 33861 39513
tri 33861 39512 33862 39513 sw
rect 29787 39511 33862 39512
tri 33862 39511 33863 39512 sw
rect 29787 39510 33863 39511
tri 33863 39510 33864 39511 sw
rect 29787 39509 33864 39510
tri 33864 39509 33865 39510 sw
rect 29787 39508 33865 39509
tri 33865 39508 33866 39509 sw
rect 29787 39507 33866 39508
tri 33866 39507 33867 39508 sw
rect 29787 39506 33867 39507
tri 33867 39506 33868 39507 sw
rect 29787 39505 33868 39506
tri 33868 39505 33869 39506 sw
rect 29787 39504 33869 39505
tri 33869 39504 33870 39505 sw
rect 29787 39503 33870 39504
tri 33870 39503 33871 39504 sw
rect 29787 39502 33871 39503
tri 33871 39502 33872 39503 sw
rect 29787 39501 33872 39502
tri 33872 39501 33873 39502 sw
rect 29787 39500 33873 39501
tri 33873 39500 33874 39501 sw
rect 29787 39499 33874 39500
tri 33874 39499 33875 39500 sw
rect 29787 39498 33875 39499
tri 33875 39498 33876 39499 sw
rect 29787 39497 33876 39498
tri 33876 39497 33877 39498 sw
rect 29787 39496 33877 39497
tri 33877 39496 33878 39497 sw
rect 29787 39495 33878 39496
tri 33878 39495 33879 39496 sw
rect 29787 39494 33879 39495
tri 33879 39494 33880 39495 sw
rect 29787 39493 33880 39494
tri 33880 39493 33881 39494 sw
rect 29787 39492 33881 39493
tri 33881 39492 33882 39493 sw
rect 29787 39491 33882 39492
tri 33882 39491 33883 39492 sw
rect 29787 39490 33883 39491
tri 33883 39490 33884 39491 sw
rect 29787 39489 33884 39490
tri 33884 39489 33885 39490 sw
rect 29787 39488 33885 39489
tri 33885 39488 33886 39489 sw
rect 29787 39487 33886 39488
tri 33886 39487 33887 39488 sw
rect 29787 39486 33887 39487
tri 33887 39486 33888 39487 sw
rect 29787 39485 33888 39486
tri 33888 39485 33889 39486 sw
rect 29787 39484 33889 39485
tri 33889 39484 33890 39485 sw
rect 29787 39483 33890 39484
tri 33890 39483 33891 39484 sw
rect 29787 39482 33891 39483
tri 33891 39482 33892 39483 sw
rect 29787 39481 33892 39482
tri 33892 39481 33893 39482 sw
rect 29787 39480 33893 39481
tri 33893 39480 33894 39481 sw
rect 29787 39479 33894 39480
tri 33894 39479 33895 39480 sw
rect 29787 39478 33895 39479
tri 33895 39478 33896 39479 sw
rect 29787 39477 33896 39478
tri 33896 39477 33897 39478 sw
rect 29787 39476 33897 39477
tri 33897 39476 33898 39477 sw
rect 29787 39475 33898 39476
tri 33898 39475 33899 39476 sw
rect 29787 39474 33899 39475
tri 33899 39474 33900 39475 sw
rect 29787 39473 33900 39474
tri 33900 39473 33901 39474 sw
rect 29787 39472 33901 39473
tri 33901 39472 33902 39473 sw
rect 29787 39471 33902 39472
tri 33902 39471 33903 39472 sw
rect 29787 39470 33903 39471
tri 33903 39470 33904 39471 sw
rect 29787 39469 33904 39470
tri 33904 39469 33905 39470 sw
rect 29787 39468 33905 39469
tri 33905 39468 33906 39469 sw
rect 29787 39467 33906 39468
tri 33906 39467 33907 39468 sw
rect 29787 39466 33907 39467
tri 33907 39466 33908 39467 sw
rect 29787 39465 33908 39466
tri 33908 39465 33909 39466 sw
rect 29787 39464 33909 39465
tri 33909 39464 33910 39465 sw
rect 29787 39463 33910 39464
tri 33910 39463 33911 39464 sw
rect 29787 39462 33911 39463
tri 33911 39462 33912 39463 sw
rect 29787 39461 33912 39462
tri 33912 39461 33913 39462 sw
rect 29787 39460 33913 39461
tri 33913 39460 33914 39461 sw
rect 29787 39459 33914 39460
tri 33914 39459 33915 39460 sw
rect 29787 39458 33915 39459
tri 33915 39458 33916 39459 sw
rect 29787 39457 33916 39458
tri 33916 39457 33917 39458 sw
rect 29787 39456 33917 39457
tri 33917 39456 33918 39457 sw
rect 29787 39455 33918 39456
tri 33918 39455 33919 39456 sw
rect 29787 39454 33919 39455
tri 33919 39454 33920 39455 sw
rect 29787 39453 33920 39454
tri 33920 39453 33921 39454 sw
rect 29787 39452 33921 39453
tri 33921 39452 33922 39453 sw
rect 29787 39451 33922 39452
tri 33922 39451 33923 39452 sw
rect 29787 39450 33923 39451
tri 33923 39450 33924 39451 sw
rect 29787 39449 33924 39450
tri 33924 39449 33925 39450 sw
rect 29787 39448 33925 39449
tri 33925 39448 33926 39449 sw
rect 29787 39447 33926 39448
tri 33926 39447 33927 39448 sw
rect 29787 39446 33927 39447
tri 33927 39446 33928 39447 sw
rect 29787 39445 33928 39446
tri 33928 39445 33929 39446 sw
rect 29787 39444 33929 39445
tri 33929 39444 33930 39445 sw
rect 29787 39443 33930 39444
tri 33930 39443 33931 39444 sw
rect 29787 39442 33931 39443
tri 33931 39442 33932 39443 sw
rect 29787 39441 33932 39442
tri 33932 39441 33933 39442 sw
rect 29787 39440 33933 39441
tri 33933 39440 33934 39441 sw
rect 29787 39439 33934 39440
tri 33934 39439 33935 39440 sw
rect 29787 39438 33935 39439
tri 33935 39438 33936 39439 sw
rect 29787 39437 33936 39438
tri 33936 39437 33937 39438 sw
rect 29787 39436 33937 39437
tri 33937 39436 33938 39437 sw
rect 29787 39435 33938 39436
tri 33938 39435 33939 39436 sw
rect 29787 39434 33939 39435
tri 33939 39434 33940 39435 sw
rect 29787 39433 33940 39434
tri 33940 39433 33941 39434 sw
rect 29787 39432 33941 39433
tri 33941 39432 33942 39433 sw
rect 29787 39431 33942 39432
tri 33942 39431 33943 39432 sw
rect 29787 39430 33943 39431
tri 33943 39430 33944 39431 sw
rect 29787 39429 33944 39430
tri 33944 39429 33945 39430 sw
rect 29787 39428 33945 39429
tri 33945 39428 33946 39429 sw
rect 29787 39427 33946 39428
tri 33946 39427 33947 39428 sw
rect 29787 39426 33947 39427
tri 33947 39426 33948 39427 sw
rect 29787 39425 33948 39426
tri 33948 39425 33949 39426 sw
rect 29787 39424 33949 39425
tri 33949 39424 33950 39425 sw
rect 29787 39423 33950 39424
tri 33950 39423 33951 39424 sw
rect 29787 39422 33951 39423
tri 33951 39422 33952 39423 sw
rect 29787 39421 33952 39422
tri 33952 39421 33953 39422 sw
rect 29787 39420 33953 39421
tri 33953 39420 33954 39421 sw
rect 29787 39419 33954 39420
tri 33954 39419 33955 39420 sw
rect 29787 39418 33955 39419
tri 33955 39418 33956 39419 sw
rect 29787 39417 33956 39418
tri 33956 39417 33957 39418 sw
rect 29787 39416 33957 39417
tri 33957 39416 33958 39417 sw
rect 29787 39415 33958 39416
tri 33958 39415 33959 39416 sw
rect 29787 39414 33959 39415
tri 33959 39414 33960 39415 sw
rect 29787 39413 33960 39414
tri 33960 39413 33961 39414 sw
rect 29787 39412 33961 39413
tri 33961 39412 33962 39413 sw
rect 29787 39411 33962 39412
tri 33962 39411 33963 39412 sw
rect 29787 39410 33963 39411
tri 33963 39410 33964 39411 sw
rect 29787 39409 33964 39410
tri 33964 39409 33965 39410 sw
rect 29787 39408 33965 39409
tri 33965 39408 33966 39409 sw
rect 29787 39407 33966 39408
tri 33966 39407 33967 39408 sw
rect 29787 39406 33967 39407
tri 33967 39406 33968 39407 sw
rect 29787 39405 33968 39406
tri 33968 39405 33969 39406 sw
rect 29787 39404 33969 39405
tri 33969 39404 33970 39405 sw
rect 29787 39403 33970 39404
tri 33970 39403 33971 39404 sw
rect 29787 39402 33971 39403
tri 33971 39402 33972 39403 sw
rect 29787 39401 33972 39402
tri 33972 39401 33973 39402 sw
rect 29787 39400 33973 39401
tri 33973 39400 33974 39401 sw
rect 29787 39399 33974 39400
tri 33974 39399 33975 39400 sw
rect 29787 39398 33975 39399
tri 33975 39398 33976 39399 sw
rect 29787 39397 33976 39398
tri 33976 39397 33977 39398 sw
rect 29787 39396 33977 39397
tri 33977 39396 33978 39397 sw
rect 29787 39395 33978 39396
tri 33978 39395 33979 39396 sw
rect 29787 39394 33979 39395
tri 33979 39394 33980 39395 sw
rect 29787 39393 33980 39394
tri 33980 39393 33981 39394 sw
rect 29787 39392 33981 39393
tri 33981 39392 33982 39393 sw
rect 29787 39391 33982 39392
tri 33982 39391 33983 39392 sw
rect 29787 39390 33983 39391
tri 33983 39390 33984 39391 sw
rect 29787 39389 33984 39390
tri 33984 39389 33985 39390 sw
rect 29787 39388 33985 39389
tri 33985 39388 33986 39389 sw
rect 29787 39387 33986 39388
tri 33986 39387 33987 39388 sw
rect 29787 39386 33987 39387
tri 33987 39386 33988 39387 sw
rect 29787 39385 33988 39386
tri 33988 39385 33989 39386 sw
rect 29787 39384 33989 39385
tri 33989 39384 33990 39385 sw
rect 29787 39383 33990 39384
tri 33990 39383 33991 39384 sw
rect 29787 39382 33991 39383
tri 33991 39382 33992 39383 sw
rect 29787 39381 33992 39382
tri 33992 39381 33993 39382 sw
rect 29787 39380 33993 39381
tri 33993 39380 33994 39381 sw
rect 29787 39379 33994 39380
tri 33994 39379 33995 39380 sw
rect 29787 39378 33995 39379
tri 33995 39378 33996 39379 sw
rect 29787 39377 33996 39378
tri 33996 39377 33997 39378 sw
rect 29787 39376 33997 39377
tri 33997 39376 33998 39377 sw
rect 29787 39375 33998 39376
tri 33998 39375 33999 39376 sw
rect 29787 39374 33999 39375
tri 33999 39374 34000 39375 sw
rect 29787 39373 34000 39374
tri 34000 39373 34001 39374 sw
rect 29787 39372 34001 39373
tri 34001 39372 34002 39373 sw
rect 29787 39371 34002 39372
tri 34002 39371 34003 39372 sw
rect 29787 39370 34003 39371
tri 34003 39370 34004 39371 sw
rect 29787 39369 34004 39370
tri 34004 39369 34005 39370 sw
rect 29787 39368 34005 39369
tri 34005 39368 34006 39369 sw
rect 29787 39367 34006 39368
tri 34006 39367 34007 39368 sw
rect 29787 39366 34007 39367
tri 34007 39366 34008 39367 sw
rect 29787 39365 34008 39366
tri 34008 39365 34009 39366 sw
rect 29787 39364 34009 39365
tri 34009 39364 34010 39365 sw
rect 29787 39363 34010 39364
tri 34010 39363 34011 39364 sw
rect 29787 39362 34011 39363
tri 34011 39362 34012 39363 sw
rect 29787 39361 34012 39362
tri 34012 39361 34013 39362 sw
rect 29787 39360 34013 39361
tri 34013 39360 34014 39361 sw
rect 29787 39359 34014 39360
tri 34014 39359 34015 39360 sw
rect 29787 39358 34015 39359
tri 34015 39358 34016 39359 sw
rect 29787 39357 34016 39358
tri 34016 39357 34017 39358 sw
rect 29787 39356 34017 39357
tri 34017 39356 34018 39357 sw
rect 29787 39355 34018 39356
tri 34018 39355 34019 39356 sw
rect 29787 39354 34019 39355
tri 34019 39354 34020 39355 sw
rect 29787 39353 34020 39354
tri 34020 39353 34021 39354 sw
rect 29787 39352 34021 39353
tri 34021 39352 34022 39353 sw
rect 29787 39351 34022 39352
tri 34022 39351 34023 39352 sw
rect 29787 39350 34023 39351
tri 34023 39350 34024 39351 sw
rect 29787 39349 34024 39350
tri 34024 39349 34025 39350 sw
rect 29787 39348 34025 39349
tri 34025 39348 34026 39349 sw
rect 29787 39347 34026 39348
tri 34026 39347 34027 39348 sw
rect 29787 39346 34027 39347
tri 34027 39346 34028 39347 sw
rect 29787 39345 34028 39346
tri 34028 39345 34029 39346 sw
rect 29787 39344 34029 39345
tri 34029 39344 34030 39345 sw
rect 29787 39343 34030 39344
tri 34030 39343 34031 39344 sw
tri 34031 39343 34328 39640 ne
rect 34328 39631 35769 39640
tri 35769 39631 36020 39882 sw
tri 36058 39631 36309 39882 ne
rect 36309 39633 37997 39882
tri 37997 39633 38287 39923 sw
tri 38287 39633 38577 39923 ne
rect 38577 39783 42377 39923
tri 42377 39783 42671 40077 sw
tri 42671 39826 42922 40077 ne
rect 42922 39865 46909 40077
tri 46909 39865 47127 40083 sw
tri 47127 39865 47415 40153 ne
rect 47415 40050 51177 40153
tri 51177 40050 51474 40347 sw
tri 51474 40073 51748 40347 ne
rect 51748 40150 55622 40347
tri 55622 40150 55915 40443 sw
tri 55915 40371 55987 40443 ne
rect 55987 40371 71000 40443
rect 51748 40078 55915 40150
tri 55915 40078 55987 40150 sw
tri 55987 40078 56280 40371 ne
rect 56280 40078 71000 40371
rect 51748 40073 55987 40078
rect 47415 39865 51474 40050
rect 42922 39826 47127 39865
rect 38577 39633 42671 39783
rect 36309 39631 38287 39633
rect 34328 39343 36020 39631
rect 25263 39341 29505 39343
rect 22232 39049 25140 39172
tri 25140 39049 25263 39172 sw
tri 25263 39049 25555 39341 ne
rect 25555 39061 29505 39341
tri 29505 39061 29787 39343 sw
tri 29787 39341 29789 39343 ne
rect 29789 39341 34031 39343
rect 25555 39059 29787 39061
tri 29787 39059 29789 39061 sw
tri 29789 39059 30071 39341 ne
rect 30071 39059 34031 39341
rect 25555 39049 29789 39059
rect 22232 38757 25263 39049
tri 25263 38757 25555 39049 sw
tri 25555 38800 25804 39049 ne
rect 25804 38800 29789 39049
rect 22232 38508 25555 38757
tri 25555 38508 25804 38757 sw
tri 25804 38508 26096 38800 ne
rect 26096 38777 29789 38800
tri 29789 38777 30071 39059 sw
tri 30071 38780 30350 39059 ne
rect 30350 39046 34031 39059
tri 34031 39046 34328 39343 sw
tri 34328 39158 34513 39343 ne
rect 34513 39342 36020 39343
tri 36020 39342 36309 39631 sw
tri 36309 39342 36598 39631 ne
rect 36598 39532 38287 39631
tri 38287 39532 38388 39633 sw
tri 38577 39532 38678 39633 ne
rect 38678 39532 42671 39633
tri 42671 39532 42922 39783 sw
tri 42922 39637 43111 39826 ne
rect 43111 39637 47127 39826
tri 43111 39532 43216 39637 ne
rect 43216 39577 47127 39637
tri 47127 39577 47415 39865 sw
tri 47415 39631 47649 39865 ne
rect 47649 39776 51474 39865
tri 51474 39776 51748 40050 sw
tri 51748 39996 51825 40073 ne
rect 51825 39996 55987 40073
rect 47649 39699 51748 39776
tri 51748 39699 51825 39776 sw
tri 51825 39699 52122 39996 ne
rect 52122 39785 55987 39996
tri 55987 39785 56280 40078 sw
tri 56280 39894 56464 40078 ne
rect 56464 39894 71000 40078
rect 52122 39699 56280 39785
rect 47649 39631 51825 39699
rect 43216 39532 47415 39577
rect 36598 39342 38388 39532
tri 38388 39342 38578 39532 sw
rect 34513 39158 36309 39342
rect 30350 38861 34328 39046
tri 34328 38861 34513 39046 sw
tri 34513 38861 34810 39158 ne
rect 34810 39149 36309 39158
tri 36309 39149 36502 39342 sw
tri 36598 39149 36791 39342 ne
rect 36791 39242 38578 39342
tri 38578 39242 38678 39342 sw
tri 38678 39242 38968 39532 ne
rect 38968 39242 42922 39532
rect 36791 39150 38678 39242
tri 38678 39150 38770 39242 sw
tri 38968 39150 39060 39242 ne
rect 39060 39238 42922 39242
tri 42922 39238 43216 39532 sw
tri 43216 39342 43406 39532 ne
rect 43406 39343 47415 39532
tri 47415 39343 47649 39577 sw
tri 47649 39343 47937 39631 ne
rect 47937 39402 51825 39631
tri 51825 39402 52122 39699 sw
tri 52122 39698 52123 39699 ne
rect 52123 39698 56280 39699
rect 47937 39401 52122 39402
tri 52122 39401 52123 39402 sw
tri 52123 39401 52420 39698 ne
rect 52420 39601 56280 39698
tri 56280 39601 56464 39785 sw
tri 56464 39693 56665 39894 ne
rect 56665 39693 71000 39894
rect 52420 39401 56464 39601
rect 47937 39343 52123 39401
rect 43406 39342 47649 39343
rect 39060 39150 43216 39238
rect 36791 39149 38770 39150
rect 34810 38861 36502 39149
rect 30350 38780 34513 38861
rect 26096 38508 30071 38777
rect 22232 38216 25804 38508
tri 25804 38216 26096 38508 sw
tri 26096 38507 26097 38508 ne
rect 26097 38507 30071 38508
rect 22232 38215 26096 38216
tri 26096 38215 26097 38216 sw
tri 26097 38215 26389 38507 ne
rect 26389 38498 30071 38507
tri 30071 38498 30350 38777 sw
tri 30350 38702 30428 38780 ne
rect 30428 38702 34513 38780
rect 26389 38420 30350 38498
tri 30350 38420 30428 38498 sw
tri 30428 38497 30633 38702 ne
rect 30633 38564 34513 38702
tri 34513 38564 34810 38861 sw
tri 34810 38860 34811 38861 ne
rect 34811 38860 36502 38861
tri 36502 38860 36791 39149 sw
tri 36791 38860 37080 39149 ne
rect 37080 38860 38770 39149
tri 38770 38860 39060 39150 sw
tri 39060 38860 39350 39150 ne
rect 39350 39048 43216 39150
tri 43216 39048 43406 39238 sw
tri 43406 39155 43593 39342 ne
rect 43593 39155 47649 39342
rect 39350 38861 43406 39048
tri 43406 38861 43593 39048 sw
tri 43593 38861 43887 39155 ne
rect 43887 39055 47649 39155
tri 47649 39055 47937 39343 sw
tri 47937 39149 48131 39343 ne
rect 48131 39149 52123 39343
rect 43887 38861 47937 39055
tri 47937 38861 48131 39055 sw
tri 48131 38861 48419 39149 ne
rect 48419 39104 52123 39149
tri 52123 39104 52420 39401 sw
tri 52420 39342 52479 39401 ne
rect 52479 39400 56464 39401
tri 56464 39400 56665 39601 sw
tri 56665 39600 56758 39693 ne
rect 56758 39600 71000 39693
rect 52479 39342 71000 39400
rect 48419 39045 52420 39104
tri 52420 39045 52479 39104 sw
tri 52479 39102 52719 39342 ne
rect 52719 39332 71000 39342
rect 52719 39102 70613 39332
rect 48419 38861 52479 39045
rect 39350 38860 43593 38861
rect 30633 38563 34810 38564
tri 34810 38563 34811 38564 sw
tri 34811 38563 35108 38860 ne
rect 35108 38769 36791 38860
tri 36791 38769 36882 38860 sw
tri 37080 38769 37171 38860 ne
rect 37171 38770 39060 38860
tri 39060 38770 39150 38860 sw
tri 39350 38770 39440 38860 ne
rect 39440 38770 43593 38860
rect 37171 38769 39150 38770
rect 35108 38563 36882 38769
rect 30633 38497 34811 38563
tri 30633 38420 30710 38497 ne
rect 30710 38420 34811 38497
rect 26389 38215 30428 38420
rect 22232 37923 26097 38215
tri 26097 37923 26389 38215 sw
tri 26389 38127 26477 38215 ne
rect 26477 38138 30428 38215
tri 30428 38138 30710 38420 sw
tri 30710 38213 30917 38420 ne
rect 30917 38266 34811 38420
tri 34811 38266 35108 38563 sw
tri 35108 38512 35159 38563 ne
rect 35159 38512 36882 38563
rect 30917 38215 35108 38266
tri 35108 38215 35159 38266 sw
tri 35159 38215 35456 38512 ne
rect 35456 38480 36882 38512
tri 36882 38480 37171 38769 sw
tri 37171 38480 37460 38769 ne
rect 37460 38480 39150 38769
tri 39150 38480 39440 38770 sw
tri 39440 38480 39730 38770 ne
rect 39730 38567 43593 38770
tri 43593 38567 43887 38861 sw
tri 43887 38775 43973 38861 ne
rect 43973 38775 48131 38861
rect 39730 38481 43887 38567
tri 43887 38481 43973 38567 sw
tri 43973 38481 44267 38775 ne
rect 44267 38573 48131 38775
tri 48131 38573 48419 38861 sw
tri 48419 38769 48511 38861 ne
rect 48511 38805 52479 38861
tri 52479 38805 52719 39045 sw
tri 52719 38860 52961 39102 ne
rect 52961 38860 70613 39102
rect 48511 38769 52719 38805
rect 44267 38481 48419 38573
tri 48419 38481 48511 38573 sw
tri 48511 38488 48792 38769 ne
rect 48792 38563 52719 38769
tri 52719 38563 52961 38805 sw
tri 52961 38778 53043 38860 ne
rect 53043 38778 70613 38860
rect 48792 38488 52961 38563
rect 39730 38480 43973 38481
rect 35456 38286 37171 38480
tri 37171 38286 37365 38480 sw
tri 37460 38286 37654 38480 ne
rect 37654 38286 39440 38480
rect 35456 38215 37365 38286
rect 30917 38213 35159 38215
rect 26477 38127 30710 38138
rect 22232 37921 26389 37923
tri 26389 37921 26391 37923 sw
tri 26477 37921 26683 38127 ne
rect 26683 37931 30710 38127
tri 30710 37931 30917 38138 sw
tri 30917 37931 31199 38213 ne
rect 31199 37931 35159 38213
rect 26683 37921 30917 37931
rect 22232 37836 26391 37921
tri 22232 33971 26097 37836 ne
rect 26097 37629 26391 37836
tri 26391 37629 26683 37921 sw
tri 26683 37757 26847 37921 ne
rect 26847 37757 30917 37921
rect 26097 37465 26683 37629
tri 26683 37465 26847 37629 sw
tri 26847 37465 27139 37757 ne
rect 27139 37649 30917 37757
tri 30917 37649 31199 37931 sw
tri 31199 37737 31393 37931 ne
rect 31393 37918 35159 37931
tri 35159 37918 35456 38215 sw
tri 35456 38214 35457 38215 ne
rect 35457 38214 37365 38215
tri 37365 38214 37437 38286 sw
tri 37654 38214 37726 38286 ne
rect 37726 38214 39440 38286
tri 39440 38214 39706 38480 sw
tri 39730 38214 39996 38480 ne
rect 39996 38214 43973 38480
rect 31393 37917 35456 37918
tri 35456 37917 35457 37918 sw
tri 35457 37917 35754 38214 ne
rect 35754 38191 37437 38214
tri 37437 38191 37460 38214 sw
tri 37726 38191 37749 38214 ne
rect 37749 38191 39706 38214
rect 35754 37917 37460 38191
rect 31393 37737 35457 37917
rect 27139 37465 31199 37649
rect 26097 37173 26847 37465
tri 26847 37173 27139 37465 sw
tri 27139 37464 27140 37465 ne
rect 27140 37464 31199 37465
rect 26097 37172 27139 37173
tri 27139 37172 27140 37173 sw
tri 27140 37172 27432 37464 ne
rect 27432 37455 31199 37464
tri 31199 37455 31393 37649 sw
tri 31393 37455 31675 37737 ne
rect 31675 37620 35457 37737
tri 35457 37620 35754 37917 sw
tri 35754 37673 35998 37917 ne
rect 35998 37902 37460 37917
tri 37460 37902 37749 38191 sw
tri 37749 37902 38038 38191 ne
rect 38038 37994 39706 38191
tri 39706 37994 39926 38214 sw
tri 39996 37994 40216 38214 ne
rect 40216 38187 43973 38214
tri 43973 38187 44267 38481 sw
tri 44267 38193 44555 38481 ne
rect 44555 38200 48511 38481
tri 48511 38200 48792 38481 sw
tri 48792 38213 49067 38488 ne
rect 49067 38481 52961 38488
tri 52961 38481 53043 38563 sw
tri 53043 38481 53340 38778 ne
rect 53340 38481 70613 38778
rect 49067 38213 53043 38481
rect 44555 38193 48792 38200
rect 40216 37994 44267 38187
rect 38038 37902 39926 37994
rect 35998 37749 37749 37902
tri 37749 37749 37902 37902 sw
tri 38038 37749 38191 37902 ne
rect 38191 37749 39926 37902
rect 35998 37673 37902 37749
rect 31675 37455 35754 37620
rect 27432 37173 31393 37455
tri 31393 37173 31675 37455 sw
tri 31675 37454 31676 37455 ne
rect 31676 37454 35754 37455
rect 27432 37172 31675 37173
tri 31675 37172 31676 37173 sw
tri 31676 37172 31958 37454 ne
rect 31958 37376 35754 37454
tri 35754 37376 35998 37620 sw
tri 35998 37469 36202 37673 ne
rect 36202 37469 37902 37673
tri 36202 37376 36295 37469 ne
rect 36295 37460 37902 37469
tri 37902 37460 38191 37749 sw
tri 38191 37460 38480 37749 ne
rect 38480 37704 39926 37749
tri 39926 37704 40216 37994 sw
tri 40216 37704 40506 37994 ne
rect 40506 37899 44267 37994
tri 44267 37899 44555 38187 sw
tri 44555 37919 44829 38193 ne
rect 44829 37925 48792 38193
tri 48792 37925 49067 38200 sw
tri 49067 37925 49355 38213 ne
rect 49355 38184 53043 38213
tri 53043 38184 53340 38481 sw
tri 53340 38213 53608 38481 ne
rect 53608 38213 70613 38481
rect 49355 37925 53340 38184
rect 44829 37919 49067 37925
rect 40506 37704 44555 37899
rect 38480 37461 40216 37704
tri 40216 37461 40459 37704 sw
tri 40506 37461 40749 37704 ne
rect 40749 37625 44555 37704
tri 44555 37625 44829 37899 sw
tri 44829 37833 44915 37919 ne
rect 44915 37833 49067 37919
rect 40749 37539 44829 37625
tri 44829 37539 44915 37625 sw
tri 44915 37539 45209 37833 ne
rect 45209 37637 49067 37833
tri 49067 37637 49355 37925 sw
tri 49355 37821 49459 37925 ne
rect 49459 37916 53340 37925
tri 53340 37916 53608 38184 sw
tri 53608 37916 53905 38213 ne
rect 53905 37916 70613 38213
rect 49459 37821 53608 37916
rect 45209 37539 49355 37637
rect 40749 37461 44915 37539
rect 38480 37460 40459 37461
rect 36295 37376 38191 37460
rect 31958 37375 35998 37376
tri 35998 37375 35999 37376 sw
rect 31958 37374 35999 37375
tri 35999 37374 36000 37375 sw
rect 31958 37373 36000 37374
tri 36000 37373 36001 37374 sw
rect 31958 37372 36001 37373
tri 36001 37372 36002 37373 sw
rect 31958 37371 36002 37372
tri 36002 37371 36003 37372 sw
rect 31958 37370 36003 37371
tri 36003 37370 36004 37371 sw
rect 31958 37369 36004 37370
tri 36004 37369 36005 37370 sw
rect 31958 37368 36005 37369
tri 36005 37368 36006 37369 sw
rect 31958 37367 36006 37368
tri 36006 37367 36007 37368 sw
rect 31958 37366 36007 37367
tri 36007 37366 36008 37367 sw
rect 31958 37365 36008 37366
tri 36008 37365 36009 37366 sw
rect 31958 37364 36009 37365
tri 36009 37364 36010 37365 sw
rect 31958 37363 36010 37364
tri 36010 37363 36011 37364 sw
rect 31958 37362 36011 37363
tri 36011 37362 36012 37363 sw
rect 31958 37361 36012 37362
tri 36012 37361 36013 37362 sw
rect 31958 37360 36013 37361
tri 36013 37360 36014 37361 sw
rect 31958 37359 36014 37360
tri 36014 37359 36015 37360 sw
rect 31958 37358 36015 37359
tri 36015 37358 36016 37359 sw
rect 31958 37357 36016 37358
tri 36016 37357 36017 37358 sw
rect 31958 37356 36017 37357
tri 36017 37356 36018 37357 sw
rect 31958 37355 36018 37356
tri 36018 37355 36019 37356 sw
rect 31958 37354 36019 37355
tri 36019 37354 36020 37355 sw
rect 31958 37353 36020 37354
tri 36020 37353 36021 37354 sw
rect 31958 37352 36021 37353
tri 36021 37352 36022 37353 sw
rect 31958 37351 36022 37352
tri 36022 37351 36023 37352 sw
rect 31958 37350 36023 37351
tri 36023 37350 36024 37351 sw
rect 31958 37349 36024 37350
tri 36024 37349 36025 37350 sw
rect 31958 37348 36025 37349
tri 36025 37348 36026 37349 sw
rect 31958 37347 36026 37348
tri 36026 37347 36027 37348 sw
rect 31958 37346 36027 37347
tri 36027 37346 36028 37347 sw
rect 31958 37345 36028 37346
tri 36028 37345 36029 37346 sw
rect 31958 37344 36029 37345
tri 36029 37344 36030 37345 sw
rect 31958 37343 36030 37344
tri 36030 37343 36031 37344 sw
rect 31958 37342 36031 37343
tri 36031 37342 36032 37343 sw
rect 31958 37341 36032 37342
tri 36032 37341 36033 37342 sw
rect 31958 37340 36033 37341
tri 36033 37340 36034 37341 sw
rect 31958 37339 36034 37340
tri 36034 37339 36035 37340 sw
rect 31958 37338 36035 37339
tri 36035 37338 36036 37339 sw
rect 31958 37337 36036 37338
tri 36036 37337 36037 37338 sw
rect 31958 37336 36037 37337
tri 36037 37336 36038 37337 sw
rect 31958 37335 36038 37336
tri 36038 37335 36039 37336 sw
rect 31958 37334 36039 37335
tri 36039 37334 36040 37335 sw
rect 31958 37333 36040 37334
tri 36040 37333 36041 37334 sw
rect 31958 37332 36041 37333
tri 36041 37332 36042 37333 sw
rect 31958 37331 36042 37332
tri 36042 37331 36043 37332 sw
rect 31958 37330 36043 37331
tri 36043 37330 36044 37331 sw
rect 31958 37329 36044 37330
tri 36044 37329 36045 37330 sw
rect 31958 37328 36045 37329
tri 36045 37328 36046 37329 sw
rect 31958 37327 36046 37328
tri 36046 37327 36047 37328 sw
rect 31958 37326 36047 37327
tri 36047 37326 36048 37327 sw
rect 31958 37325 36048 37326
tri 36048 37325 36049 37326 sw
rect 31958 37324 36049 37325
tri 36049 37324 36050 37325 sw
rect 31958 37323 36050 37324
tri 36050 37323 36051 37324 sw
rect 31958 37322 36051 37323
tri 36051 37322 36052 37323 sw
rect 31958 37321 36052 37322
tri 36052 37321 36053 37322 sw
rect 31958 37320 36053 37321
tri 36053 37320 36054 37321 sw
rect 31958 37319 36054 37320
tri 36054 37319 36055 37320 sw
rect 31958 37318 36055 37319
tri 36055 37318 36056 37319 sw
rect 31958 37317 36056 37318
tri 36056 37317 36057 37318 sw
rect 31958 37316 36057 37317
tri 36057 37316 36058 37317 sw
rect 31958 37315 36058 37316
tri 36058 37315 36059 37316 sw
rect 31958 37314 36059 37315
tri 36059 37314 36060 37315 sw
rect 31958 37313 36060 37314
tri 36060 37313 36061 37314 sw
rect 31958 37312 36061 37313
tri 36061 37312 36062 37313 sw
rect 31958 37311 36062 37312
tri 36062 37311 36063 37312 sw
rect 31958 37310 36063 37311
tri 36063 37310 36064 37311 sw
rect 31958 37309 36064 37310
tri 36064 37309 36065 37310 sw
rect 31958 37308 36065 37309
tri 36065 37308 36066 37309 sw
rect 31958 37307 36066 37308
tri 36066 37307 36067 37308 sw
rect 31958 37306 36067 37307
tri 36067 37306 36068 37307 sw
rect 31958 37305 36068 37306
tri 36068 37305 36069 37306 sw
rect 31958 37304 36069 37305
tri 36069 37304 36070 37305 sw
rect 31958 37303 36070 37304
tri 36070 37303 36071 37304 sw
rect 31958 37302 36071 37303
tri 36071 37302 36072 37303 sw
rect 31958 37301 36072 37302
tri 36072 37301 36073 37302 sw
rect 31958 37300 36073 37301
tri 36073 37300 36074 37301 sw
rect 31958 37299 36074 37300
tri 36074 37299 36075 37300 sw
rect 31958 37298 36075 37299
tri 36075 37298 36076 37299 sw
rect 31958 37297 36076 37298
tri 36076 37297 36077 37298 sw
rect 31958 37296 36077 37297
tri 36077 37296 36078 37297 sw
rect 31958 37295 36078 37296
tri 36078 37295 36079 37296 sw
rect 31958 37294 36079 37295
tri 36079 37294 36080 37295 sw
rect 31958 37293 36080 37294
tri 36080 37293 36081 37294 sw
rect 31958 37292 36081 37293
tri 36081 37292 36082 37293 sw
rect 31958 37291 36082 37292
tri 36082 37291 36083 37292 sw
rect 31958 37290 36083 37291
tri 36083 37290 36084 37291 sw
rect 31958 37289 36084 37290
tri 36084 37289 36085 37290 sw
rect 31958 37288 36085 37289
tri 36085 37288 36086 37289 sw
rect 31958 37287 36086 37288
tri 36086 37287 36087 37288 sw
rect 31958 37286 36087 37287
tri 36087 37286 36088 37287 sw
rect 31958 37285 36088 37286
tri 36088 37285 36089 37286 sw
rect 31958 37284 36089 37285
tri 36089 37284 36090 37285 sw
rect 31958 37283 36090 37284
tri 36090 37283 36091 37284 sw
rect 31958 37282 36091 37283
tri 36091 37282 36092 37283 sw
rect 31958 37281 36092 37282
tri 36092 37281 36093 37282 sw
rect 31958 37280 36093 37281
tri 36093 37280 36094 37281 sw
rect 31958 37279 36094 37280
tri 36094 37279 36095 37280 sw
rect 31958 37278 36095 37279
tri 36095 37278 36096 37279 sw
rect 31958 37277 36096 37278
tri 36096 37277 36097 37278 sw
rect 31958 37276 36097 37277
tri 36097 37276 36098 37277 sw
rect 31958 37275 36098 37276
tri 36098 37275 36099 37276 sw
rect 31958 37274 36099 37275
tri 36099 37274 36100 37275 sw
rect 31958 37273 36100 37274
tri 36100 37273 36101 37274 sw
rect 31958 37272 36101 37273
tri 36101 37272 36102 37273 sw
rect 31958 37271 36102 37272
tri 36102 37271 36103 37272 sw
rect 31958 37270 36103 37271
tri 36103 37270 36104 37271 sw
rect 31958 37269 36104 37270
tri 36104 37269 36105 37270 sw
rect 31958 37268 36105 37269
tri 36105 37268 36106 37269 sw
rect 31958 37267 36106 37268
tri 36106 37267 36107 37268 sw
rect 31958 37266 36107 37267
tri 36107 37266 36108 37267 sw
rect 31958 37265 36108 37266
tri 36108 37265 36109 37266 sw
rect 31958 37264 36109 37265
tri 36109 37264 36110 37265 sw
rect 31958 37263 36110 37264
tri 36110 37263 36111 37264 sw
rect 31958 37262 36111 37263
tri 36111 37262 36112 37263 sw
rect 31958 37261 36112 37262
tri 36112 37261 36113 37262 sw
rect 31958 37260 36113 37261
tri 36113 37260 36114 37261 sw
rect 31958 37259 36114 37260
tri 36114 37259 36115 37260 sw
rect 31958 37258 36115 37259
tri 36115 37258 36116 37259 sw
rect 31958 37257 36116 37258
tri 36116 37257 36117 37258 sw
rect 31958 37256 36117 37257
tri 36117 37256 36118 37257 sw
rect 31958 37255 36118 37256
tri 36118 37255 36119 37256 sw
rect 31958 37254 36119 37255
tri 36119 37254 36120 37255 sw
rect 31958 37253 36120 37254
tri 36120 37253 36121 37254 sw
rect 31958 37252 36121 37253
tri 36121 37252 36122 37253 sw
rect 31958 37251 36122 37252
tri 36122 37251 36123 37252 sw
rect 31958 37250 36123 37251
tri 36123 37250 36124 37251 sw
rect 31958 37249 36124 37250
tri 36124 37249 36125 37250 sw
rect 31958 37248 36125 37249
tri 36125 37248 36126 37249 sw
rect 31958 37247 36126 37248
tri 36126 37247 36127 37248 sw
rect 31958 37246 36127 37247
tri 36127 37246 36128 37247 sw
rect 31958 37245 36128 37246
tri 36128 37245 36129 37246 sw
rect 31958 37244 36129 37245
tri 36129 37244 36130 37245 sw
rect 31958 37243 36130 37244
tri 36130 37243 36131 37244 sw
rect 31958 37242 36131 37243
tri 36131 37242 36132 37243 sw
rect 31958 37241 36132 37242
tri 36132 37241 36133 37242 sw
rect 31958 37240 36133 37241
tri 36133 37240 36134 37241 sw
rect 31958 37239 36134 37240
tri 36134 37239 36135 37240 sw
rect 31958 37238 36135 37239
tri 36135 37238 36136 37239 sw
rect 31958 37237 36136 37238
tri 36136 37237 36137 37238 sw
rect 31958 37236 36137 37237
tri 36137 37236 36138 37237 sw
rect 31958 37235 36138 37236
tri 36138 37235 36139 37236 sw
rect 31958 37234 36139 37235
tri 36139 37234 36140 37235 sw
rect 31958 37233 36140 37234
tri 36140 37233 36141 37234 sw
rect 31958 37232 36141 37233
tri 36141 37232 36142 37233 sw
rect 31958 37231 36142 37232
tri 36142 37231 36143 37232 sw
rect 31958 37230 36143 37231
tri 36143 37230 36144 37231 sw
rect 31958 37229 36144 37230
tri 36144 37229 36145 37230 sw
rect 31958 37228 36145 37229
tri 36145 37228 36146 37229 sw
rect 31958 37227 36146 37228
tri 36146 37227 36147 37228 sw
rect 31958 37226 36147 37227
tri 36147 37226 36148 37227 sw
rect 31958 37225 36148 37226
tri 36148 37225 36149 37226 sw
rect 31958 37224 36149 37225
tri 36149 37224 36150 37225 sw
rect 31958 37223 36150 37224
tri 36150 37223 36151 37224 sw
rect 31958 37222 36151 37223
tri 36151 37222 36152 37223 sw
rect 31958 37221 36152 37222
tri 36152 37221 36153 37222 sw
rect 31958 37220 36153 37221
tri 36153 37220 36154 37221 sw
rect 31958 37219 36154 37220
tri 36154 37219 36155 37220 sw
rect 31958 37218 36155 37219
tri 36155 37218 36156 37219 sw
rect 31958 37217 36156 37218
tri 36156 37217 36157 37218 sw
rect 31958 37216 36157 37217
tri 36157 37216 36158 37217 sw
rect 31958 37215 36158 37216
tri 36158 37215 36159 37216 sw
rect 31958 37214 36159 37215
tri 36159 37214 36160 37215 sw
rect 31958 37213 36160 37214
tri 36160 37213 36161 37214 sw
rect 31958 37212 36161 37213
tri 36161 37212 36162 37213 sw
rect 31958 37211 36162 37212
tri 36162 37211 36163 37212 sw
rect 31958 37210 36163 37211
tri 36163 37210 36164 37211 sw
rect 31958 37209 36164 37210
tri 36164 37209 36165 37210 sw
rect 31958 37208 36165 37209
tri 36165 37208 36166 37209 sw
rect 31958 37207 36166 37208
tri 36166 37207 36167 37208 sw
rect 31958 37206 36167 37207
tri 36167 37206 36168 37207 sw
rect 31958 37205 36168 37206
tri 36168 37205 36169 37206 sw
rect 31958 37204 36169 37205
tri 36169 37204 36170 37205 sw
rect 31958 37203 36170 37204
tri 36170 37203 36171 37204 sw
rect 31958 37202 36171 37203
tri 36171 37202 36172 37203 sw
rect 31958 37201 36172 37202
tri 36172 37201 36173 37202 sw
rect 31958 37200 36173 37201
tri 36173 37200 36174 37201 sw
rect 31958 37199 36174 37200
tri 36174 37199 36175 37200 sw
rect 31958 37198 36175 37199
tri 36175 37198 36176 37199 sw
rect 31958 37197 36176 37198
tri 36176 37197 36177 37198 sw
rect 31958 37196 36177 37197
tri 36177 37196 36178 37197 sw
rect 31958 37195 36178 37196
tri 36178 37195 36179 37196 sw
rect 31958 37194 36179 37195
tri 36179 37194 36180 37195 sw
rect 31958 37193 36180 37194
tri 36180 37193 36181 37194 sw
rect 31958 37192 36181 37193
tri 36181 37192 36182 37193 sw
rect 31958 37191 36182 37192
tri 36182 37191 36183 37192 sw
rect 31958 37190 36183 37191
tri 36183 37190 36184 37191 sw
rect 31958 37189 36184 37190
tri 36184 37189 36185 37190 sw
rect 31958 37188 36185 37189
tri 36185 37188 36186 37189 sw
rect 31958 37187 36186 37188
tri 36186 37187 36187 37188 sw
rect 31958 37186 36187 37187
tri 36187 37186 36188 37187 sw
rect 31958 37185 36188 37186
tri 36188 37185 36189 37186 sw
rect 31958 37184 36189 37185
tri 36189 37184 36190 37185 sw
rect 31958 37183 36190 37184
tri 36190 37183 36191 37184 sw
rect 31958 37182 36191 37183
tri 36191 37182 36192 37183 sw
rect 31958 37181 36192 37182
tri 36192 37181 36193 37182 sw
rect 31958 37180 36193 37181
tri 36193 37180 36194 37181 sw
rect 31958 37179 36194 37180
tri 36194 37179 36195 37180 sw
rect 31958 37178 36195 37179
tri 36195 37178 36196 37179 sw
rect 31958 37177 36196 37178
tri 36196 37177 36197 37178 sw
rect 31958 37176 36197 37177
tri 36197 37176 36198 37177 sw
rect 31958 37175 36198 37176
tri 36198 37175 36199 37176 sw
rect 31958 37174 36199 37175
tri 36199 37174 36200 37175 sw
rect 31958 37173 36200 37174
tri 36200 37173 36201 37174 sw
rect 31958 37172 36201 37173
tri 36201 37172 36202 37173 sw
rect 26097 36880 27140 37172
tri 27140 36880 27432 37172 sw
tri 27432 37171 27433 37172 ne
rect 27433 37171 31676 37172
rect 26097 36879 27432 36880
tri 27432 36879 27433 36880 sw
tri 27433 36879 27725 37171 ne
rect 27725 36890 31676 37171
tri 31676 36890 31958 37172 sw
tri 31958 37171 31959 37172 ne
rect 31959 37171 36202 37172
tri 36202 37171 36203 37172 sw
tri 36295 37171 36500 37376 ne
rect 36500 37171 38191 37376
tri 38191 37171 38480 37460 sw
tri 38480 37171 38769 37460 ne
rect 38769 37171 40459 37460
tri 40459 37171 40749 37461 sw
tri 40749 37171 41039 37461 ne
rect 41039 37245 44915 37461
tri 44915 37245 45209 37539 sw
tri 45209 37537 45211 37539 ne
rect 45211 37537 49355 37539
rect 41039 37243 45209 37245
tri 45209 37243 45211 37245 sw
tri 45211 37243 45505 37537 ne
rect 45505 37533 49355 37537
tri 49355 37533 49459 37637 sw
tri 49459 37533 49747 37821 ne
rect 49747 37619 53608 37821
tri 53608 37619 53905 37916 sw
tri 53905 37741 54080 37916 ne
rect 54080 37741 70613 37916
rect 49747 37533 53905 37619
rect 45505 37245 49459 37533
tri 49459 37245 49747 37533 sw
tri 49747 37444 49836 37533 ne
rect 49836 37444 53905 37533
tri 53905 37444 54080 37619 sw
tri 54080 37540 54281 37741 ne
rect 54281 37540 70613 37741
rect 45505 37243 49747 37245
rect 41039 37171 45211 37243
rect 27725 36889 31958 36890
tri 31958 36889 31959 36890 sw
tri 31959 36889 32241 37171 ne
rect 32241 36889 36203 37171
rect 27725 36879 31959 36889
rect 26097 36587 27433 36879
tri 27433 36587 27725 36879 sw
tri 27725 36751 27853 36879 ne
rect 27853 36751 31959 36879
rect 26097 36459 27725 36587
tri 27725 36459 27853 36587 sw
tri 27853 36459 28145 36751 ne
rect 28145 36607 31959 36751
tri 31959 36607 32241 36889 sw
tri 32241 36741 32389 36889 ne
rect 32389 36874 36203 36889
tri 36203 36874 36500 37171 sw
tri 36500 36880 36791 37171 ne
rect 36791 37169 38480 37171
tri 38480 37169 38482 37171 sw
tri 38769 37169 38771 37171 ne
rect 38771 37170 40749 37171
tri 40749 37170 40750 37171 sw
tri 41039 37170 41040 37171 ne
rect 41040 37170 45211 37171
rect 38771 37169 40750 37170
rect 36791 36880 38482 37169
tri 38482 36880 38771 37169 sw
tri 38771 36880 39060 37169 ne
rect 39060 36880 40750 37169
tri 40750 36880 41040 37170 sw
tri 41040 36880 41330 37170 ne
rect 41330 36949 45211 37170
tri 45211 36949 45505 37243 sw
tri 45505 37171 45577 37243 ne
rect 45577 37171 49747 37243
rect 41330 36880 45505 36949
rect 32389 36741 36500 36874
rect 28145 36459 32241 36607
tri 32241 36459 32389 36607 sw
tri 32389 36459 32671 36741 ne
rect 32671 36583 36500 36741
tri 36500 36583 36791 36874 sw
tri 36791 36583 37088 36880 ne
rect 37088 36789 38771 36880
tri 38771 36789 38862 36880 sw
tri 39060 36789 39151 36880 ne
rect 39151 36790 41040 36880
tri 41040 36790 41130 36880 sw
tri 41330 36790 41420 36880 ne
rect 41420 36877 45505 36880
tri 45505 36877 45577 36949 sw
tri 45577 36880 45868 37171 ne
rect 45868 37156 49747 37171
tri 49747 37156 49836 37245 sw
tri 49836 37156 50124 37444 ne
rect 50124 37443 54080 37444
tri 54080 37443 54081 37444 sw
rect 50124 37442 54081 37443
tri 54081 37442 54082 37443 sw
rect 50124 37441 54082 37442
tri 54082 37441 54083 37442 sw
rect 50124 37440 54083 37441
tri 54083 37440 54084 37441 sw
rect 50124 37439 54084 37440
tri 54084 37439 54085 37440 sw
rect 50124 37438 54085 37439
tri 54085 37438 54086 37439 sw
rect 50124 37437 54086 37438
tri 54086 37437 54087 37438 sw
rect 50124 37436 54087 37437
tri 54087 37436 54088 37437 sw
rect 50124 37435 54088 37436
tri 54088 37435 54089 37436 sw
rect 50124 37434 54089 37435
tri 54089 37434 54090 37435 sw
rect 50124 37433 54090 37434
tri 54090 37433 54091 37434 sw
rect 50124 37432 54091 37433
tri 54091 37432 54092 37433 sw
rect 50124 37431 54092 37432
tri 54092 37431 54093 37432 sw
rect 50124 37430 54093 37431
tri 54093 37430 54094 37431 sw
rect 50124 37429 54094 37430
tri 54094 37429 54095 37430 sw
rect 50124 37428 54095 37429
tri 54095 37428 54096 37429 sw
rect 50124 37427 54096 37428
tri 54096 37427 54097 37428 sw
rect 50124 37426 54097 37427
tri 54097 37426 54098 37427 sw
rect 50124 37425 54098 37426
tri 54098 37425 54099 37426 sw
rect 50124 37424 54099 37425
tri 54099 37424 54100 37425 sw
rect 50124 37423 54100 37424
tri 54100 37423 54101 37424 sw
rect 50124 37422 54101 37423
tri 54101 37422 54102 37423 sw
rect 50124 37421 54102 37422
tri 54102 37421 54103 37422 sw
rect 50124 37420 54103 37421
tri 54103 37420 54104 37421 sw
rect 50124 37419 54104 37420
tri 54104 37419 54105 37420 sw
rect 50124 37418 54105 37419
tri 54105 37418 54106 37419 sw
rect 50124 37417 54106 37418
tri 54106 37417 54107 37418 sw
rect 50124 37416 54107 37417
tri 54107 37416 54108 37417 sw
rect 50124 37415 54108 37416
tri 54108 37415 54109 37416 sw
rect 50124 37414 54109 37415
tri 54109 37414 54110 37415 sw
rect 50124 37413 54110 37414
tri 54110 37413 54111 37414 sw
rect 50124 37412 54111 37413
tri 54111 37412 54112 37413 sw
rect 50124 37411 54112 37412
tri 54112 37411 54113 37412 sw
rect 50124 37410 54113 37411
tri 54113 37410 54114 37411 sw
rect 50124 37409 54114 37410
tri 54114 37409 54115 37410 sw
rect 50124 37408 54115 37409
tri 54115 37408 54116 37409 sw
rect 50124 37407 54116 37408
tri 54116 37407 54117 37408 sw
rect 50124 37406 54117 37407
tri 54117 37406 54118 37407 sw
rect 50124 37405 54118 37406
tri 54118 37405 54119 37406 sw
rect 50124 37404 54119 37405
tri 54119 37404 54120 37405 sw
rect 50124 37403 54120 37404
tri 54120 37403 54121 37404 sw
rect 50124 37402 54121 37403
tri 54121 37402 54122 37403 sw
rect 50124 37401 54122 37402
tri 54122 37401 54123 37402 sw
rect 50124 37400 54123 37401
tri 54123 37400 54124 37401 sw
rect 50124 37399 54124 37400
tri 54124 37399 54125 37400 sw
rect 50124 37398 54125 37399
tri 54125 37398 54126 37399 sw
rect 50124 37397 54126 37398
tri 54126 37397 54127 37398 sw
rect 50124 37396 54127 37397
tri 54127 37396 54128 37397 sw
rect 50124 37395 54128 37396
tri 54128 37395 54129 37396 sw
rect 50124 37394 54129 37395
tri 54129 37394 54130 37395 sw
rect 50124 37393 54130 37394
tri 54130 37393 54131 37394 sw
rect 50124 37392 54131 37393
tri 54131 37392 54132 37393 sw
rect 50124 37391 54132 37392
tri 54132 37391 54133 37392 sw
rect 50124 37390 54133 37391
tri 54133 37390 54134 37391 sw
rect 50124 37389 54134 37390
tri 54134 37389 54135 37390 sw
rect 50124 37388 54135 37389
tri 54135 37388 54136 37389 sw
rect 50124 37387 54136 37388
tri 54136 37387 54137 37388 sw
rect 50124 37386 54137 37387
tri 54137 37386 54138 37387 sw
rect 50124 37385 54138 37386
tri 54138 37385 54139 37386 sw
rect 50124 37384 54139 37385
tri 54139 37384 54140 37385 sw
rect 50124 37383 54140 37384
tri 54140 37383 54141 37384 sw
rect 50124 37382 54141 37383
tri 54141 37382 54142 37383 sw
rect 50124 37381 54142 37382
tri 54142 37381 54143 37382 sw
rect 50124 37380 54143 37381
tri 54143 37380 54144 37381 sw
rect 50124 37379 54144 37380
tri 54144 37379 54145 37380 sw
rect 50124 37378 54145 37379
tri 54145 37378 54146 37379 sw
rect 50124 37377 54146 37378
tri 54146 37377 54147 37378 sw
rect 50124 37376 54147 37377
tri 54147 37376 54148 37377 sw
rect 50124 37375 54148 37376
tri 54148 37375 54149 37376 sw
rect 50124 37374 54149 37375
tri 54149 37374 54150 37375 sw
rect 50124 37373 54150 37374
tri 54150 37373 54151 37374 sw
rect 50124 37372 54151 37373
tri 54151 37372 54152 37373 sw
rect 50124 37371 54152 37372
tri 54152 37371 54153 37372 sw
rect 50124 37370 54153 37371
tri 54153 37370 54154 37371 sw
rect 50124 37369 54154 37370
tri 54154 37369 54155 37370 sw
rect 50124 37368 54155 37369
tri 54155 37368 54156 37369 sw
rect 50124 37367 54156 37368
tri 54156 37367 54157 37368 sw
rect 50124 37366 54157 37367
tri 54157 37366 54158 37367 sw
rect 50124 37365 54158 37366
tri 54158 37365 54159 37366 sw
rect 50124 37364 54159 37365
tri 54159 37364 54160 37365 sw
rect 50124 37363 54160 37364
tri 54160 37363 54161 37364 sw
rect 50124 37362 54161 37363
tri 54161 37362 54162 37363 sw
rect 50124 37361 54162 37362
tri 54162 37361 54163 37362 sw
rect 50124 37360 54163 37361
tri 54163 37360 54164 37361 sw
rect 50124 37359 54164 37360
tri 54164 37359 54165 37360 sw
rect 50124 37358 54165 37359
tri 54165 37358 54166 37359 sw
rect 50124 37357 54166 37358
tri 54166 37357 54167 37358 sw
rect 50124 37356 54167 37357
tri 54167 37356 54168 37357 sw
rect 50124 37355 54168 37356
tri 54168 37355 54169 37356 sw
rect 50124 37354 54169 37355
tri 54169 37354 54170 37355 sw
rect 50124 37353 54170 37354
tri 54170 37353 54171 37354 sw
rect 50124 37352 54171 37353
tri 54171 37352 54172 37353 sw
rect 50124 37351 54172 37352
tri 54172 37351 54173 37352 sw
rect 50124 37350 54173 37351
tri 54173 37350 54174 37351 sw
rect 50124 37349 54174 37350
tri 54174 37349 54175 37350 sw
rect 50124 37348 54175 37349
tri 54175 37348 54176 37349 sw
rect 50124 37347 54176 37348
tri 54176 37347 54177 37348 sw
rect 50124 37346 54177 37347
tri 54177 37346 54178 37347 sw
rect 50124 37345 54178 37346
tri 54178 37345 54179 37346 sw
rect 50124 37344 54179 37345
tri 54179 37344 54180 37345 sw
rect 50124 37343 54180 37344
tri 54180 37343 54181 37344 sw
rect 50124 37342 54181 37343
tri 54181 37342 54182 37343 sw
rect 50124 37341 54182 37342
tri 54182 37341 54183 37342 sw
rect 50124 37340 54183 37341
tri 54183 37340 54184 37341 sw
rect 50124 37339 54184 37340
tri 54184 37339 54185 37340 sw
rect 50124 37338 54185 37339
tri 54185 37338 54186 37339 sw
rect 50124 37337 54186 37338
tri 54186 37337 54187 37338 sw
rect 50124 37336 54187 37337
tri 54187 37336 54188 37337 sw
rect 50124 37335 54188 37336
tri 54188 37335 54189 37336 sw
rect 50124 37334 54189 37335
tri 54189 37334 54190 37335 sw
rect 50124 37333 54190 37334
tri 54190 37333 54191 37334 sw
rect 50124 37332 54191 37333
tri 54191 37332 54192 37333 sw
rect 50124 37331 54192 37332
tri 54192 37331 54193 37332 sw
rect 50124 37330 54193 37331
tri 54193 37330 54194 37331 sw
rect 50124 37329 54194 37330
tri 54194 37329 54195 37330 sw
rect 50124 37328 54195 37329
tri 54195 37328 54196 37329 sw
rect 50124 37327 54196 37328
tri 54196 37327 54197 37328 sw
rect 50124 37326 54197 37327
tri 54197 37326 54198 37327 sw
rect 50124 37325 54198 37326
tri 54198 37325 54199 37326 sw
rect 50124 37324 54199 37325
tri 54199 37324 54200 37325 sw
rect 50124 37323 54200 37324
tri 54200 37323 54201 37324 sw
rect 50124 37322 54201 37323
tri 54201 37322 54202 37323 sw
rect 50124 37321 54202 37322
tri 54202 37321 54203 37322 sw
rect 50124 37320 54203 37321
tri 54203 37320 54204 37321 sw
rect 50124 37319 54204 37320
tri 54204 37319 54205 37320 sw
rect 50124 37318 54205 37319
tri 54205 37318 54206 37319 sw
rect 50124 37317 54206 37318
tri 54206 37317 54207 37318 sw
rect 50124 37316 54207 37317
tri 54207 37316 54208 37317 sw
rect 50124 37315 54208 37316
tri 54208 37315 54209 37316 sw
rect 50124 37314 54209 37315
tri 54209 37314 54210 37315 sw
rect 50124 37313 54210 37314
tri 54210 37313 54211 37314 sw
rect 50124 37312 54211 37313
tri 54211 37312 54212 37313 sw
rect 50124 37311 54212 37312
tri 54212 37311 54213 37312 sw
rect 50124 37310 54213 37311
tri 54213 37310 54214 37311 sw
rect 50124 37309 54214 37310
tri 54214 37309 54215 37310 sw
rect 50124 37308 54215 37309
tri 54215 37308 54216 37309 sw
rect 50124 37307 54216 37308
tri 54216 37307 54217 37308 sw
rect 50124 37306 54217 37307
tri 54217 37306 54218 37307 sw
rect 50124 37305 54218 37306
tri 54218 37305 54219 37306 sw
rect 50124 37304 54219 37305
tri 54219 37304 54220 37305 sw
rect 50124 37303 54220 37304
tri 54220 37303 54221 37304 sw
rect 50124 37302 54221 37303
tri 54221 37302 54222 37303 sw
rect 50124 37301 54222 37302
tri 54222 37301 54223 37302 sw
rect 50124 37300 54223 37301
tri 54223 37300 54224 37301 sw
rect 50124 37299 54224 37300
tri 54224 37299 54225 37300 sw
rect 50124 37298 54225 37299
tri 54225 37298 54226 37299 sw
rect 50124 37297 54226 37298
tri 54226 37297 54227 37298 sw
rect 50124 37296 54227 37297
tri 54227 37296 54228 37297 sw
rect 50124 37295 54228 37296
tri 54228 37295 54229 37296 sw
rect 50124 37294 54229 37295
tri 54229 37294 54230 37295 sw
rect 50124 37293 54230 37294
tri 54230 37293 54231 37294 sw
rect 50124 37292 54231 37293
tri 54231 37292 54232 37293 sw
rect 50124 37291 54232 37292
tri 54232 37291 54233 37292 sw
rect 50124 37290 54233 37291
tri 54233 37290 54234 37291 sw
rect 50124 37289 54234 37290
tri 54234 37289 54235 37290 sw
rect 50124 37288 54235 37289
tri 54235 37288 54236 37289 sw
rect 50124 37287 54236 37288
tri 54236 37287 54237 37288 sw
rect 50124 37286 54237 37287
tri 54237 37286 54238 37287 sw
rect 50124 37285 54238 37286
tri 54238 37285 54239 37286 sw
rect 50124 37284 54239 37285
tri 54239 37284 54240 37285 sw
rect 50124 37283 54240 37284
tri 54240 37283 54241 37284 sw
rect 50124 37282 54241 37283
tri 54241 37282 54242 37283 sw
rect 50124 37281 54242 37282
tri 54242 37281 54243 37282 sw
rect 50124 37280 54243 37281
tri 54243 37280 54244 37281 sw
rect 50124 37279 54244 37280
tri 54244 37279 54245 37280 sw
rect 50124 37278 54245 37279
tri 54245 37278 54246 37279 sw
rect 50124 37277 54246 37278
tri 54246 37277 54247 37278 sw
rect 50124 37276 54247 37277
tri 54247 37276 54248 37277 sw
rect 50124 37275 54248 37276
tri 54248 37275 54249 37276 sw
rect 50124 37274 54249 37275
tri 54249 37274 54250 37275 sw
rect 50124 37273 54250 37274
tri 54250 37273 54251 37274 sw
rect 50124 37272 54251 37273
tri 54251 37272 54252 37273 sw
rect 50124 37271 54252 37272
tri 54252 37271 54253 37272 sw
rect 50124 37270 54253 37271
tri 54253 37270 54254 37271 sw
rect 50124 37269 54254 37270
tri 54254 37269 54255 37270 sw
rect 50124 37268 54255 37269
tri 54255 37268 54256 37269 sw
rect 50124 37267 54256 37268
tri 54256 37267 54257 37268 sw
rect 50124 37266 54257 37267
tri 54257 37266 54258 37267 sw
rect 50124 37265 54258 37266
tri 54258 37265 54259 37266 sw
rect 50124 37264 54259 37265
tri 54259 37264 54260 37265 sw
rect 50124 37263 54260 37264
tri 54260 37263 54261 37264 sw
rect 50124 37262 54261 37263
tri 54261 37262 54262 37263 sw
rect 50124 37261 54262 37262
tri 54262 37261 54263 37262 sw
rect 50124 37260 54263 37261
tri 54263 37260 54264 37261 sw
rect 50124 37259 54264 37260
tri 54264 37259 54265 37260 sw
rect 50124 37258 54265 37259
tri 54265 37258 54266 37259 sw
rect 50124 37257 54266 37258
tri 54266 37257 54267 37258 sw
rect 50124 37256 54267 37257
tri 54267 37256 54268 37257 sw
rect 50124 37255 54268 37256
tri 54268 37255 54269 37256 sw
rect 50124 37254 54269 37255
tri 54269 37254 54270 37255 sw
rect 50124 37253 54270 37254
tri 54270 37253 54271 37254 sw
rect 50124 37252 54271 37253
tri 54271 37252 54272 37253 sw
rect 50124 37251 54272 37252
tri 54272 37251 54273 37252 sw
rect 50124 37250 54273 37251
tri 54273 37250 54274 37251 sw
rect 50124 37249 54274 37250
tri 54274 37249 54275 37250 sw
rect 50124 37248 54275 37249
tri 54275 37248 54276 37249 sw
rect 50124 37247 54276 37248
tri 54276 37247 54277 37248 sw
rect 50124 37246 54277 37247
tri 54277 37246 54278 37247 sw
rect 50124 37245 54278 37246
tri 54278 37245 54279 37246 sw
rect 50124 37244 54279 37245
tri 54279 37244 54280 37245 sw
rect 50124 37243 54280 37244
tri 54280 37243 54281 37244 sw
tri 54281 37243 54578 37540 ne
rect 54578 37243 70613 37540
rect 50124 37156 54281 37243
rect 45868 36880 49836 37156
rect 41420 36790 45577 36877
rect 39151 36789 41130 36790
rect 37088 36583 38862 36789
rect 32671 36459 36791 36583
rect 26097 36167 27853 36459
tri 27853 36167 28145 36459 sw
tri 28145 36435 28169 36459 ne
rect 28169 36435 32389 36459
rect 26097 36143 28145 36167
tri 28145 36143 28169 36167 sw
tri 28169 36143 28461 36435 ne
rect 28461 36177 32389 36435
tri 32389 36177 32671 36459 sw
tri 32671 36425 32705 36459 ne
rect 32705 36425 36791 36459
rect 28461 36143 32671 36177
tri 32671 36143 32705 36177 sw
tri 32705 36143 32987 36425 ne
rect 32987 36286 36791 36425
tri 36791 36286 37088 36583 sw
tri 37088 36440 37231 36583 ne
rect 37231 36500 38862 36583
tri 38862 36500 39151 36789 sw
tri 39151 36500 39440 36789 ne
rect 39440 36500 41130 36789
tri 41130 36500 41420 36790 sw
tri 41420 36500 41710 36790 ne
rect 41710 36586 45577 36790
tri 45577 36586 45868 36877 sw
tri 45868 36795 45953 36880 ne
rect 45953 36868 49836 36880
tri 49836 36868 50124 37156 sw
tri 50124 36880 50400 37156 ne
rect 50400 36946 54281 37156
tri 54281 36946 54578 37243 sw
tri 54578 37171 54650 37243 ne
rect 54650 37171 70613 37243
rect 50400 36880 54578 36946
rect 45953 36795 50124 36868
rect 41710 36501 45868 36586
tri 45868 36501 45953 36586 sw
tri 45953 36501 46247 36795 ne
rect 46247 36592 50124 36795
tri 50124 36592 50400 36868 sw
tri 50400 36789 50491 36880 ne
rect 50491 36874 54578 36880
tri 54578 36874 54650 36946 sw
tri 54650 36880 54941 37171 ne
rect 54941 36880 70613 37171
rect 50491 36789 54650 36874
rect 46247 36501 50400 36592
tri 50400 36501 50491 36592 sw
tri 50491 36501 50779 36789 ne
rect 50779 36583 54650 36789
tri 54650 36583 54941 36874 sw
tri 54941 36798 55023 36880 ne
rect 55023 36798 70613 36880
rect 50779 36501 54941 36583
tri 54941 36501 55023 36583 sw
tri 55023 36501 55320 36798 ne
rect 55320 36501 70613 36798
rect 41710 36500 45953 36501
rect 37231 36440 39151 36500
rect 32987 36143 37088 36286
tri 37088 36143 37231 36286 sw
tri 37231 36143 37528 36440 ne
rect 37528 36211 39151 36440
tri 39151 36211 39440 36500 sw
tri 39440 36211 39729 36500 ne
rect 39729 36432 41420 36500
tri 41420 36432 41488 36500 sw
tri 41710 36432 41778 36500 ne
rect 41778 36432 45953 36500
rect 39729 36211 41488 36432
rect 37528 36143 39440 36211
rect 26097 35851 28169 36143
tri 28169 35851 28461 36143 sw
tri 28461 36141 28463 36143 ne
rect 28463 36141 32705 36143
rect 26097 35849 28461 35851
tri 28461 35849 28463 35851 sw
tri 28463 35849 28755 36141 ne
rect 28755 35861 32705 36141
tri 32705 35861 32987 36143 sw
tri 32987 36128 33002 36143 ne
rect 33002 36128 37231 36143
rect 28755 35849 32987 35861
rect 26097 35848 28463 35849
tri 28463 35848 28464 35849 sw
tri 28755 35848 28756 35849 ne
rect 28756 35848 32987 35849
rect 26097 35556 28464 35848
tri 28464 35556 28756 35848 sw
tri 28756 35556 29048 35848 ne
rect 29048 35846 32987 35848
tri 32987 35846 33002 35861 sw
tri 33002 35846 33284 36128 ne
rect 33284 35846 37231 36128
tri 37231 35846 37528 36143 sw
tri 37528 36128 37543 36143 ne
rect 37543 36128 39440 36143
tri 39440 36128 39523 36211 sw
tri 39729 36128 39812 36211 ne
rect 39812 36142 41488 36211
tri 41488 36142 41778 36432 sw
tri 41778 36142 42068 36432 ne
rect 42068 36207 45953 36432
tri 45953 36207 46247 36501 sw
tri 46247 36437 46311 36501 ne
rect 46311 36437 50491 36501
rect 42068 36143 46247 36207
tri 46247 36143 46311 36207 sw
tri 46311 36143 46605 36437 ne
rect 46605 36213 50491 36437
tri 50491 36213 50779 36501 sw
tri 50779 36458 50822 36501 ne
rect 50822 36458 55023 36501
rect 46605 36170 50779 36213
tri 50779 36170 50822 36213 sw
tri 50822 36200 51080 36458 ne
rect 51080 36204 55023 36458
tri 55023 36204 55320 36501 sw
tri 55320 36400 55421 36501 ne
rect 55421 36468 70613 36501
rect 70669 36468 71000 39332
rect 55421 36400 71000 36468
rect 51080 36200 55320 36204
tri 55320 36200 55324 36204 sw
rect 46605 36143 50822 36170
rect 42068 36142 46311 36143
rect 39812 36128 41778 36142
tri 41778 36128 41792 36142 sw
tri 42068 36128 42082 36142 ne
rect 42082 36128 46311 36142
rect 29048 35564 33002 35846
tri 33002 35564 33284 35846 sw
tri 33284 35845 33285 35846 ne
rect 33285 35845 37528 35846
rect 29048 35563 33284 35564
tri 33284 35563 33285 35564 sw
tri 33285 35563 33567 35845 ne
rect 33567 35831 37528 35845
tri 37528 35831 37543 35846 sw
tri 37543 35831 37840 36128 ne
rect 37840 35839 39523 36128
tri 39523 35839 39812 36128 sw
tri 39812 35839 40101 36128 ne
rect 40101 35839 41792 36128
rect 37840 35831 39812 35839
rect 33567 35563 37543 35831
rect 29048 35556 33285 35563
rect 26097 35264 28756 35556
tri 28756 35264 29048 35556 sw
tri 29048 35512 29092 35556 ne
rect 29092 35512 33285 35556
rect 26097 35220 29048 35264
tri 29048 35220 29092 35264 sw
tri 29092 35262 29342 35512 ne
rect 29342 35281 33285 35512
tri 33285 35281 33567 35563 sw
tri 33567 35561 33569 35563 ne
rect 33569 35561 37543 35563
rect 29342 35279 33567 35281
tri 33567 35279 33569 35281 sw
tri 33569 35279 33851 35561 ne
rect 33851 35534 37543 35561
tri 37543 35534 37840 35831 sw
tri 37840 35534 38137 35831 ne
rect 38137 35550 39812 35831
tri 39812 35550 40101 35839 sw
tri 40101 35550 40390 35839 ne
rect 40390 35838 41792 35839
tri 41792 35838 42082 36128 sw
tri 42082 35838 42372 36128 ne
rect 42372 35849 46311 36128
tri 46311 35849 46605 36143 sw
tri 46605 36128 46620 36143 ne
rect 46620 36128 50822 36143
rect 42372 35838 46605 35849
rect 40390 35837 42082 35838
tri 42082 35837 42083 35838 sw
tri 42372 35837 42373 35838 ne
rect 42373 35837 46605 35838
rect 40390 35550 42083 35837
rect 38137 35534 40101 35550
rect 33851 35279 37840 35534
rect 29342 35278 33569 35279
tri 33569 35278 33570 35279 sw
tri 33851 35278 33852 35279 ne
rect 33852 35278 37840 35279
rect 29342 35262 33570 35278
rect 26097 35219 29092 35220
tri 29092 35219 29093 35220 sw
rect 26097 35218 29093 35219
tri 29093 35218 29094 35219 sw
rect 26097 35217 29094 35218
tri 29094 35217 29095 35218 sw
rect 26097 35216 29095 35217
tri 29095 35216 29096 35217 sw
rect 26097 35215 29096 35216
tri 29096 35215 29097 35216 sw
rect 26097 35214 29097 35215
tri 29097 35214 29098 35215 sw
rect 26097 35213 29098 35214
tri 29098 35213 29099 35214 sw
rect 26097 35212 29099 35213
tri 29099 35212 29100 35213 sw
rect 26097 35211 29100 35212
tri 29100 35211 29101 35212 sw
rect 26097 35210 29101 35211
tri 29101 35210 29102 35211 sw
rect 26097 35209 29102 35210
tri 29102 35209 29103 35210 sw
rect 26097 35208 29103 35209
tri 29103 35208 29104 35209 sw
rect 26097 35207 29104 35208
tri 29104 35207 29105 35208 sw
rect 26097 35206 29105 35207
tri 29105 35206 29106 35207 sw
rect 26097 35205 29106 35206
tri 29106 35205 29107 35206 sw
rect 26097 35204 29107 35205
tri 29107 35204 29108 35205 sw
rect 26097 35203 29108 35204
tri 29108 35203 29109 35204 sw
rect 26097 35202 29109 35203
tri 29109 35202 29110 35203 sw
rect 26097 35201 29110 35202
tri 29110 35201 29111 35202 sw
rect 26097 35200 29111 35201
tri 29111 35200 29112 35201 sw
rect 26097 35199 29112 35200
tri 29112 35199 29113 35200 sw
rect 26097 35198 29113 35199
tri 29113 35198 29114 35199 sw
rect 26097 35197 29114 35198
tri 29114 35197 29115 35198 sw
rect 26097 35196 29115 35197
tri 29115 35196 29116 35197 sw
rect 26097 35195 29116 35196
tri 29116 35195 29117 35196 sw
rect 26097 35194 29117 35195
tri 29117 35194 29118 35195 sw
rect 26097 35193 29118 35194
tri 29118 35193 29119 35194 sw
rect 26097 35192 29119 35193
tri 29119 35192 29120 35193 sw
rect 26097 35191 29120 35192
tri 29120 35191 29121 35192 sw
rect 26097 35190 29121 35191
tri 29121 35190 29122 35191 sw
rect 26097 35189 29122 35190
tri 29122 35189 29123 35190 sw
rect 26097 35188 29123 35189
tri 29123 35188 29124 35189 sw
rect 26097 35187 29124 35188
tri 29124 35187 29125 35188 sw
rect 26097 35186 29125 35187
tri 29125 35186 29126 35187 sw
rect 26097 35185 29126 35186
tri 29126 35185 29127 35186 sw
rect 26097 35184 29127 35185
tri 29127 35184 29128 35185 sw
rect 26097 35183 29128 35184
tri 29128 35183 29129 35184 sw
rect 26097 35182 29129 35183
tri 29129 35182 29130 35183 sw
rect 26097 35181 29130 35182
tri 29130 35181 29131 35182 sw
rect 26097 35180 29131 35181
tri 29131 35180 29132 35181 sw
rect 26097 35179 29132 35180
tri 29132 35179 29133 35180 sw
rect 26097 35178 29133 35179
tri 29133 35178 29134 35179 sw
rect 26097 35177 29134 35178
tri 29134 35177 29135 35178 sw
rect 26097 35176 29135 35177
tri 29135 35176 29136 35177 sw
rect 26097 35175 29136 35176
tri 29136 35175 29137 35176 sw
rect 26097 35174 29137 35175
tri 29137 35174 29138 35175 sw
rect 26097 35173 29138 35174
tri 29138 35173 29139 35174 sw
rect 26097 35172 29139 35173
tri 29139 35172 29140 35173 sw
rect 26097 35171 29140 35172
tri 29140 35171 29141 35172 sw
rect 26097 35170 29141 35171
tri 29141 35170 29142 35171 sw
rect 26097 35169 29142 35170
tri 29142 35169 29143 35170 sw
rect 26097 35168 29143 35169
tri 29143 35168 29144 35169 sw
rect 26097 35167 29144 35168
tri 29144 35167 29145 35168 sw
rect 26097 35166 29145 35167
tri 29145 35166 29146 35167 sw
rect 26097 35165 29146 35166
tri 29146 35165 29147 35166 sw
rect 26097 35164 29147 35165
tri 29147 35164 29148 35165 sw
rect 26097 35163 29148 35164
tri 29148 35163 29149 35164 sw
rect 26097 35162 29149 35163
tri 29149 35162 29150 35163 sw
rect 26097 35161 29150 35162
tri 29150 35161 29151 35162 sw
rect 26097 35160 29151 35161
tri 29151 35160 29152 35161 sw
rect 26097 35159 29152 35160
tri 29152 35159 29153 35160 sw
rect 26097 35158 29153 35159
tri 29153 35158 29154 35159 sw
rect 26097 35157 29154 35158
tri 29154 35157 29155 35158 sw
rect 26097 35156 29155 35157
tri 29155 35156 29156 35157 sw
rect 26097 35155 29156 35156
tri 29156 35155 29157 35156 sw
rect 26097 35154 29157 35155
tri 29157 35154 29158 35155 sw
rect 26097 35153 29158 35154
tri 29158 35153 29159 35154 sw
rect 26097 35152 29159 35153
tri 29159 35152 29160 35153 sw
rect 26097 35151 29160 35152
tri 29160 35151 29161 35152 sw
rect 26097 35150 29161 35151
tri 29161 35150 29162 35151 sw
rect 26097 35149 29162 35150
tri 29162 35149 29163 35150 sw
rect 26097 35148 29163 35149
tri 29163 35148 29164 35149 sw
rect 26097 35147 29164 35148
tri 29164 35147 29165 35148 sw
rect 26097 35146 29165 35147
tri 29165 35146 29166 35147 sw
rect 26097 35145 29166 35146
tri 29166 35145 29167 35146 sw
rect 26097 35144 29167 35145
tri 29167 35144 29168 35145 sw
rect 26097 35143 29168 35144
tri 29168 35143 29169 35144 sw
tri 29342 35143 29461 35262 ne
rect 29461 35143 33570 35262
rect 26097 34851 29169 35143
tri 29169 34851 29461 35143 sw
tri 29461 34851 29753 35143 ne
rect 29753 34996 33570 35143
tri 33570 34996 33852 35278 sw
tri 33852 34996 34134 35278 ne
rect 34134 35237 37840 35278
tri 37840 35237 38137 35534 sw
tri 38137 35495 38176 35534 ne
rect 38176 35495 40101 35534
rect 34134 35198 38137 35237
tri 38137 35198 38176 35237 sw
tri 38176 35198 38473 35495 ne
rect 38473 35288 40101 35495
tri 40101 35288 40363 35550 sw
tri 40390 35288 40652 35550 ne
rect 40652 35547 42083 35550
tri 42083 35547 42373 35837 sw
tri 42373 35547 42663 35837 ne
rect 42663 35834 46605 35837
tri 46605 35834 46620 35849 sw
tri 46620 35834 46914 36128 ne
rect 46914 35912 50822 36128
tri 50822 35912 51080 36170 sw
tri 51080 36128 51152 36200 ne
rect 51152 36132 71000 36200
rect 51152 36128 70613 36132
rect 46914 35910 51080 35912
tri 51080 35910 51082 35912 sw
tri 51152 35910 51370 36128 ne
rect 51370 35910 70613 36128
rect 46914 35834 51082 35910
rect 42663 35547 46620 35834
rect 40652 35288 42373 35547
tri 42373 35288 42632 35547 sw
tri 42663 35288 42922 35547 ne
rect 42922 35540 46620 35547
tri 46620 35540 46914 35834 sw
tri 46914 35582 47166 35834 ne
rect 47166 35622 51082 35834
tri 51082 35622 51370 35910 sw
tri 51370 35622 51658 35910 ne
rect 51658 35622 70613 35910
rect 47166 35582 51370 35622
rect 42922 35288 46914 35540
tri 46914 35288 47166 35540 sw
tri 47166 35490 47258 35582 ne
rect 47258 35490 51370 35582
tri 47258 35288 47460 35490 ne
rect 47460 35334 51370 35490
tri 51370 35334 51658 35622 sw
tri 51658 35478 51802 35622 ne
rect 51802 35478 70613 35622
rect 47460 35288 51658 35334
rect 38473 35198 40363 35288
rect 34134 34996 38176 35198
rect 29753 34851 33852 34996
rect 26097 34850 29461 34851
tri 29461 34850 29462 34851 sw
tri 29753 34850 29754 34851 ne
rect 29754 34850 33852 34851
rect 26097 34558 29462 34850
tri 29462 34558 29754 34850 sw
tri 29754 34558 30046 34850 ne
rect 30046 34820 33852 34850
tri 33852 34820 34028 34996 sw
tri 34134 34820 34310 34996 ne
rect 34310 34901 38176 34996
tri 38176 34901 38473 35198 sw
tri 38473 34901 38770 35198 ne
rect 38770 35189 40363 35198
tri 40363 35189 40462 35288 sw
tri 40652 35189 40751 35288 ne
rect 40751 35191 42632 35288
tri 42632 35191 42729 35288 sw
rect 40751 35189 42729 35191
rect 38770 34901 40462 35189
rect 34310 34820 38473 34901
rect 30046 34558 34028 34820
rect 26097 34266 29754 34558
tri 29754 34266 30046 34558 sw
tri 30046 34557 30047 34558 ne
rect 30047 34557 34028 34558
rect 26097 34265 30046 34266
tri 30046 34265 30047 34266 sw
tri 30047 34265 30339 34557 ne
rect 30339 34538 34028 34557
tri 34028 34538 34310 34820 sw
tri 34310 34538 34592 34820 ne
rect 34592 34604 38473 34820
tri 38473 34604 38770 34901 sw
tri 38770 34900 38771 34901 ne
rect 38771 34900 40462 34901
tri 40462 34900 40751 35189 sw
tri 40751 34900 41040 35189 ne
rect 41040 34998 42729 35189
tri 42729 34998 42922 35191 sw
tri 42922 34998 43212 35288 ne
rect 43212 34998 47166 35288
rect 41040 34900 42922 34998
rect 34592 34603 38770 34604
tri 38770 34603 38771 34604 sw
tri 38771 34603 39068 34900 ne
rect 39068 34809 40751 34900
tri 40751 34809 40842 34900 sw
tri 41040 34809 41131 34900 ne
rect 41131 34810 42922 34900
tri 42922 34810 43110 34998 sw
tri 43212 34810 43400 34998 ne
rect 43400 34994 47166 34998
tri 47166 34994 47460 35288 sw
tri 47460 35195 47553 35288 ne
rect 47553 35195 51658 35288
rect 43400 34901 47460 34994
tri 47460 34901 47553 34994 sw
tri 47553 34901 47847 35195 ne
rect 47847 35190 51658 35195
tri 51658 35190 51802 35334 sw
tri 51802 35190 52090 35478 ne
rect 52090 35190 70613 35478
rect 47847 34902 51802 35190
tri 51802 34902 52090 35190 sw
tri 52090 35189 52091 35190 ne
rect 52091 35189 70613 35190
rect 47847 34901 52090 34902
tri 52090 34901 52091 34902 sw
tri 52091 34901 52379 35189 ne
rect 52379 34901 70613 35189
rect 43400 34810 47553 34901
rect 41131 34809 43110 34810
rect 39068 34603 40842 34809
rect 34592 34538 38771 34603
rect 30339 34265 34310 34538
rect 26097 33973 30047 34265
tri 30047 33973 30339 34265 sw
tri 30339 34264 30340 34265 ne
rect 30340 34264 34310 34265
rect 26097 33972 30339 33973
tri 30339 33972 30340 33973 sw
tri 30340 33972 30632 34264 ne
rect 30632 34256 34310 34264
tri 34310 34256 34592 34538 sw
tri 34592 34458 34672 34538 ne
rect 34672 34458 38771 34538
rect 30632 34176 34592 34256
tri 34592 34176 34672 34256 sw
tri 34672 34254 34876 34458 ne
rect 34876 34306 38771 34458
tri 38771 34306 39068 34603 sw
tri 39068 34602 39069 34603 ne
rect 39069 34602 40842 34603
rect 34876 34305 39068 34306
tri 39068 34305 39069 34306 sw
tri 39069 34305 39366 34602 ne
rect 39366 34520 40842 34602
tri 40842 34520 41131 34809 sw
tri 41131 34520 41420 34809 ne
rect 41420 34520 43110 34809
tri 43110 34520 43400 34810 sw
tri 43400 34520 43690 34810 ne
rect 43690 34607 47553 34810
tri 47553 34607 47847 34901 sw
tri 47847 34815 47933 34901 ne
rect 47933 34815 52091 34901
rect 43690 34521 47847 34607
tri 47847 34521 47933 34607 sw
tri 47933 34521 48227 34815 ne
rect 48227 34613 52091 34815
tri 52091 34613 52379 34901 sw
tri 52379 34809 52471 34901 ne
rect 52471 34809 70613 34901
rect 48227 34521 52379 34613
tri 52379 34521 52471 34613 sw
tri 52471 34532 52748 34809 ne
rect 52748 34532 70613 34809
rect 43690 34520 47933 34521
rect 39366 34305 41131 34520
rect 34876 34254 39069 34305
tri 34876 34176 34954 34254 ne
rect 34954 34176 39069 34254
rect 30632 33972 34672 34176
rect 26097 33971 30340 33972
tri 26097 29728 30340 33971 ne
tri 30340 33680 30632 33972 sw
tri 30632 33971 30633 33972 ne
rect 30633 33971 34672 33972
rect 30340 33679 30632 33680
tri 30632 33679 30633 33680 sw
tri 30633 33679 30925 33971 ne
rect 30925 33894 34672 33971
tri 34672 33894 34954 34176 sw
tri 34954 33971 35159 34176 ne
rect 35159 34008 39069 34176
tri 39069 34008 39366 34305 sw
tri 39366 34269 39402 34305 ne
rect 39402 34269 41131 34305
rect 35159 33972 39366 34008
tri 39366 33972 39402 34008 sw
tri 39402 33972 39699 34269 ne
rect 39699 34231 41131 34269
tri 41131 34231 41420 34520 sw
tri 41420 34231 41709 34520 ne
rect 41709 34333 43400 34520
tri 43400 34333 43587 34520 sw
tri 43690 34333 43877 34520 ne
rect 43877 34333 47933 34520
rect 41709 34231 43587 34333
rect 39699 34043 41420 34231
tri 41420 34043 41608 34231 sw
tri 41709 34043 41897 34231 ne
rect 41897 34043 43587 34231
tri 43587 34043 43877 34333 sw
tri 43877 34043 44167 34333 ne
rect 44167 34227 47933 34333
tri 47933 34227 48227 34521 sw
tri 48227 34244 48504 34521 ne
rect 48504 34244 52471 34521
tri 52471 34244 52748 34521 sw
tri 52748 34331 52949 34532 ne
rect 52949 34331 70613 34532
rect 44167 34043 48227 34227
rect 39699 33972 41608 34043
rect 35159 33971 39402 33972
rect 30925 33689 34954 33894
tri 34954 33689 35159 33894 sw
tri 35159 33689 35441 33971 ne
rect 35441 33689 39402 33971
rect 30925 33679 35159 33689
rect 30340 33387 30633 33679
tri 30633 33387 30925 33679 sw
tri 30925 33551 31053 33679 ne
rect 31053 33551 35159 33679
rect 30340 33259 30925 33387
tri 30925 33259 31053 33387 sw
tri 31053 33259 31345 33551 ne
rect 31345 33407 35159 33551
tri 35159 33407 35441 33689 sw
tri 35441 33541 35589 33689 ne
rect 35589 33675 39402 33689
tri 39402 33675 39699 33972 sw
tri 39699 33971 39700 33972 ne
rect 39700 33971 41608 33972
tri 41608 33971 41680 34043 sw
tri 41897 33971 41969 34043 ne
rect 41969 33971 43877 34043
tri 43877 33971 43949 34043 sw
tri 44167 33971 44239 34043 ne
rect 44239 33971 48227 34043
rect 35589 33674 39699 33675
tri 39699 33674 39700 33675 sw
tri 39700 33674 39997 33971 ne
rect 39997 33682 41680 33971
tri 41680 33682 41969 33971 sw
tri 41969 33682 42258 33971 ne
rect 42258 33752 43949 33971
tri 43949 33752 44168 33971 sw
tri 44239 33752 44458 33971 ne
rect 44458 33950 48227 33971
tri 48227 33950 48504 34227 sw
tri 48504 33950 48798 34244 ne
rect 48798 34243 52748 34244
tri 52748 34243 52749 34244 sw
rect 48798 34242 52749 34243
tri 52749 34242 52750 34243 sw
rect 48798 34241 52750 34242
tri 52750 34241 52751 34242 sw
rect 48798 34240 52751 34241
tri 52751 34240 52752 34241 sw
rect 48798 34239 52752 34240
tri 52752 34239 52753 34240 sw
rect 48798 34238 52753 34239
tri 52753 34238 52754 34239 sw
rect 48798 34237 52754 34238
tri 52754 34237 52755 34238 sw
rect 48798 34236 52755 34237
tri 52755 34236 52756 34237 sw
rect 48798 34235 52756 34236
tri 52756 34235 52757 34236 sw
rect 48798 34234 52757 34235
tri 52757 34234 52758 34235 sw
rect 48798 34233 52758 34234
tri 52758 34233 52759 34234 sw
rect 48798 34232 52759 34233
tri 52759 34232 52760 34233 sw
rect 48798 34231 52760 34232
tri 52760 34231 52761 34232 sw
rect 48798 34230 52761 34231
tri 52761 34230 52762 34231 sw
rect 48798 34229 52762 34230
tri 52762 34229 52763 34230 sw
rect 48798 34228 52763 34229
tri 52763 34228 52764 34229 sw
rect 48798 34227 52764 34228
tri 52764 34227 52765 34228 sw
rect 48798 34226 52765 34227
tri 52765 34226 52766 34227 sw
rect 48798 34225 52766 34226
tri 52766 34225 52767 34226 sw
rect 48798 34224 52767 34225
tri 52767 34224 52768 34225 sw
rect 48798 34223 52768 34224
tri 52768 34223 52769 34224 sw
rect 48798 34222 52769 34223
tri 52769 34222 52770 34223 sw
rect 48798 34221 52770 34222
tri 52770 34221 52771 34222 sw
rect 48798 34220 52771 34221
tri 52771 34220 52772 34221 sw
rect 48798 34219 52772 34220
tri 52772 34219 52773 34220 sw
rect 48798 34218 52773 34219
tri 52773 34218 52774 34219 sw
rect 48798 34217 52774 34218
tri 52774 34217 52775 34218 sw
rect 48798 34216 52775 34217
tri 52775 34216 52776 34217 sw
rect 48798 34215 52776 34216
tri 52776 34215 52777 34216 sw
rect 48798 34214 52777 34215
tri 52777 34214 52778 34215 sw
rect 48798 34213 52778 34214
tri 52778 34213 52779 34214 sw
rect 48798 34212 52779 34213
tri 52779 34212 52780 34213 sw
rect 48798 34211 52780 34212
tri 52780 34211 52781 34212 sw
rect 48798 34210 52781 34211
tri 52781 34210 52782 34211 sw
rect 48798 34209 52782 34210
tri 52782 34209 52783 34210 sw
rect 48798 34208 52783 34209
tri 52783 34208 52784 34209 sw
rect 48798 34207 52784 34208
tri 52784 34207 52785 34208 sw
rect 48798 34206 52785 34207
tri 52785 34206 52786 34207 sw
rect 48798 34205 52786 34206
tri 52786 34205 52787 34206 sw
rect 48798 34204 52787 34205
tri 52787 34204 52788 34205 sw
rect 48798 34203 52788 34204
tri 52788 34203 52789 34204 sw
rect 48798 34202 52789 34203
tri 52789 34202 52790 34203 sw
rect 48798 34201 52790 34202
tri 52790 34201 52791 34202 sw
rect 48798 34200 52791 34201
tri 52791 34200 52792 34201 sw
rect 48798 34199 52792 34200
tri 52792 34199 52793 34200 sw
rect 48798 34198 52793 34199
tri 52793 34198 52794 34199 sw
rect 48798 34197 52794 34198
tri 52794 34197 52795 34198 sw
rect 48798 34196 52795 34197
tri 52795 34196 52796 34197 sw
rect 48798 34195 52796 34196
tri 52796 34195 52797 34196 sw
rect 48798 34194 52797 34195
tri 52797 34194 52798 34195 sw
rect 48798 34193 52798 34194
tri 52798 34193 52799 34194 sw
rect 48798 34192 52799 34193
tri 52799 34192 52800 34193 sw
rect 48798 34191 52800 34192
tri 52800 34191 52801 34192 sw
rect 48798 34190 52801 34191
tri 52801 34190 52802 34191 sw
rect 48798 34189 52802 34190
tri 52802 34189 52803 34190 sw
rect 48798 34188 52803 34189
tri 52803 34188 52804 34189 sw
rect 48798 34187 52804 34188
tri 52804 34187 52805 34188 sw
rect 48798 34186 52805 34187
tri 52805 34186 52806 34187 sw
rect 48798 34185 52806 34186
tri 52806 34185 52807 34186 sw
rect 48798 34184 52807 34185
tri 52807 34184 52808 34185 sw
rect 48798 34183 52808 34184
tri 52808 34183 52809 34184 sw
rect 48798 34182 52809 34183
tri 52809 34182 52810 34183 sw
rect 48798 34181 52810 34182
tri 52810 34181 52811 34182 sw
rect 48798 34180 52811 34181
tri 52811 34180 52812 34181 sw
rect 48798 34179 52812 34180
tri 52812 34179 52813 34180 sw
rect 48798 34178 52813 34179
tri 52813 34178 52814 34179 sw
rect 48798 34177 52814 34178
tri 52814 34177 52815 34178 sw
rect 48798 34176 52815 34177
tri 52815 34176 52816 34177 sw
rect 48798 34175 52816 34176
tri 52816 34175 52817 34176 sw
rect 48798 34174 52817 34175
tri 52817 34174 52818 34175 sw
rect 48798 34173 52818 34174
tri 52818 34173 52819 34174 sw
rect 48798 34172 52819 34173
tri 52819 34172 52820 34173 sw
rect 48798 34171 52820 34172
tri 52820 34171 52821 34172 sw
rect 48798 34170 52821 34171
tri 52821 34170 52822 34171 sw
rect 48798 34169 52822 34170
tri 52822 34169 52823 34170 sw
rect 48798 34168 52823 34169
tri 52823 34168 52824 34169 sw
rect 48798 34167 52824 34168
tri 52824 34167 52825 34168 sw
rect 48798 34166 52825 34167
tri 52825 34166 52826 34167 sw
rect 48798 34165 52826 34166
tri 52826 34165 52827 34166 sw
rect 48798 34164 52827 34165
tri 52827 34164 52828 34165 sw
rect 48798 34163 52828 34164
tri 52828 34163 52829 34164 sw
rect 48798 34162 52829 34163
tri 52829 34162 52830 34163 sw
rect 48798 34161 52830 34162
tri 52830 34161 52831 34162 sw
rect 48798 34160 52831 34161
tri 52831 34160 52832 34161 sw
rect 48798 34159 52832 34160
tri 52832 34159 52833 34160 sw
rect 48798 34158 52833 34159
tri 52833 34158 52834 34159 sw
rect 48798 34157 52834 34158
tri 52834 34157 52835 34158 sw
rect 48798 34156 52835 34157
tri 52835 34156 52836 34157 sw
rect 48798 34155 52836 34156
tri 52836 34155 52837 34156 sw
rect 48798 34154 52837 34155
tri 52837 34154 52838 34155 sw
rect 48798 34153 52838 34154
tri 52838 34153 52839 34154 sw
rect 48798 34152 52839 34153
tri 52839 34152 52840 34153 sw
rect 48798 34151 52840 34152
tri 52840 34151 52841 34152 sw
rect 48798 34150 52841 34151
tri 52841 34150 52842 34151 sw
rect 48798 34149 52842 34150
tri 52842 34149 52843 34150 sw
rect 48798 34148 52843 34149
tri 52843 34148 52844 34149 sw
rect 48798 34147 52844 34148
tri 52844 34147 52845 34148 sw
rect 48798 34146 52845 34147
tri 52845 34146 52846 34147 sw
rect 48798 34145 52846 34146
tri 52846 34145 52847 34146 sw
rect 48798 34144 52847 34145
tri 52847 34144 52848 34145 sw
rect 48798 34143 52848 34144
tri 52848 34143 52849 34144 sw
rect 48798 34142 52849 34143
tri 52849 34142 52850 34143 sw
rect 48798 34141 52850 34142
tri 52850 34141 52851 34142 sw
rect 48798 34140 52851 34141
tri 52851 34140 52852 34141 sw
rect 48798 34139 52852 34140
tri 52852 34139 52853 34140 sw
rect 48798 34138 52853 34139
tri 52853 34138 52854 34139 sw
rect 48798 34137 52854 34138
tri 52854 34137 52855 34138 sw
rect 48798 34136 52855 34137
tri 52855 34136 52856 34137 sw
rect 48798 34135 52856 34136
tri 52856 34135 52857 34136 sw
rect 48798 34134 52857 34135
tri 52857 34134 52858 34135 sw
rect 48798 34133 52858 34134
tri 52858 34133 52859 34134 sw
rect 48798 34132 52859 34133
tri 52859 34132 52860 34133 sw
rect 48798 34131 52860 34132
tri 52860 34131 52861 34132 sw
rect 48798 34130 52861 34131
tri 52861 34130 52862 34131 sw
rect 48798 34129 52862 34130
tri 52862 34129 52863 34130 sw
rect 48798 34128 52863 34129
tri 52863 34128 52864 34129 sw
rect 48798 34127 52864 34128
tri 52864 34127 52865 34128 sw
rect 48798 34126 52865 34127
tri 52865 34126 52866 34127 sw
rect 48798 34125 52866 34126
tri 52866 34125 52867 34126 sw
rect 48798 34124 52867 34125
tri 52867 34124 52868 34125 sw
rect 48798 34123 52868 34124
tri 52868 34123 52869 34124 sw
rect 48798 34122 52869 34123
tri 52869 34122 52870 34123 sw
rect 48798 34121 52870 34122
tri 52870 34121 52871 34122 sw
rect 48798 34120 52871 34121
tri 52871 34120 52872 34121 sw
rect 48798 34119 52872 34120
tri 52872 34119 52873 34120 sw
rect 48798 34118 52873 34119
tri 52873 34118 52874 34119 sw
rect 48798 34117 52874 34118
tri 52874 34117 52875 34118 sw
rect 48798 34116 52875 34117
tri 52875 34116 52876 34117 sw
rect 48798 34115 52876 34116
tri 52876 34115 52877 34116 sw
rect 48798 34114 52877 34115
tri 52877 34114 52878 34115 sw
rect 48798 34113 52878 34114
tri 52878 34113 52879 34114 sw
rect 48798 34112 52879 34113
tri 52879 34112 52880 34113 sw
rect 48798 34111 52880 34112
tri 52880 34111 52881 34112 sw
rect 48798 34110 52881 34111
tri 52881 34110 52882 34111 sw
rect 48798 34109 52882 34110
tri 52882 34109 52883 34110 sw
rect 48798 34108 52883 34109
tri 52883 34108 52884 34109 sw
rect 48798 34107 52884 34108
tri 52884 34107 52885 34108 sw
rect 48798 34106 52885 34107
tri 52885 34106 52886 34107 sw
rect 48798 34105 52886 34106
tri 52886 34105 52887 34106 sw
rect 48798 34104 52887 34105
tri 52887 34104 52888 34105 sw
rect 48798 34103 52888 34104
tri 52888 34103 52889 34104 sw
rect 48798 34102 52889 34103
tri 52889 34102 52890 34103 sw
rect 48798 34101 52890 34102
tri 52890 34101 52891 34102 sw
rect 48798 34100 52891 34101
tri 52891 34100 52892 34101 sw
rect 48798 34099 52892 34100
tri 52892 34099 52893 34100 sw
rect 48798 34098 52893 34099
tri 52893 34098 52894 34099 sw
rect 48798 34097 52894 34098
tri 52894 34097 52895 34098 sw
rect 48798 34096 52895 34097
tri 52895 34096 52896 34097 sw
rect 48798 34095 52896 34096
tri 52896 34095 52897 34096 sw
rect 48798 34094 52897 34095
tri 52897 34094 52898 34095 sw
rect 48798 34093 52898 34094
tri 52898 34093 52899 34094 sw
rect 48798 34092 52899 34093
tri 52899 34092 52900 34093 sw
rect 48798 34091 52900 34092
tri 52900 34091 52901 34092 sw
rect 48798 34090 52901 34091
tri 52901 34090 52902 34091 sw
rect 48798 34089 52902 34090
tri 52902 34089 52903 34090 sw
rect 48798 34088 52903 34089
tri 52903 34088 52904 34089 sw
rect 48798 34087 52904 34088
tri 52904 34087 52905 34088 sw
rect 48798 34086 52905 34087
tri 52905 34086 52906 34087 sw
rect 48798 34085 52906 34086
tri 52906 34085 52907 34086 sw
rect 48798 34084 52907 34085
tri 52907 34084 52908 34085 sw
rect 48798 34083 52908 34084
tri 52908 34083 52909 34084 sw
rect 48798 34082 52909 34083
tri 52909 34082 52910 34083 sw
rect 48798 34081 52910 34082
tri 52910 34081 52911 34082 sw
rect 48798 34080 52911 34081
tri 52911 34080 52912 34081 sw
rect 48798 34079 52912 34080
tri 52912 34079 52913 34080 sw
rect 48798 34078 52913 34079
tri 52913 34078 52914 34079 sw
rect 48798 34077 52914 34078
tri 52914 34077 52915 34078 sw
rect 48798 34076 52915 34077
tri 52915 34076 52916 34077 sw
rect 48798 34075 52916 34076
tri 52916 34075 52917 34076 sw
rect 48798 34074 52917 34075
tri 52917 34074 52918 34075 sw
rect 48798 34073 52918 34074
tri 52918 34073 52919 34074 sw
rect 48798 34072 52919 34073
tri 52919 34072 52920 34073 sw
rect 48798 34071 52920 34072
tri 52920 34071 52921 34072 sw
rect 48798 34070 52921 34071
tri 52921 34070 52922 34071 sw
rect 48798 34069 52922 34070
tri 52922 34069 52923 34070 sw
rect 48798 34068 52923 34069
tri 52923 34068 52924 34069 sw
rect 48798 34067 52924 34068
tri 52924 34067 52925 34068 sw
rect 48798 34066 52925 34067
tri 52925 34066 52926 34067 sw
rect 48798 34065 52926 34066
tri 52926 34065 52927 34066 sw
rect 48798 34064 52927 34065
tri 52927 34064 52928 34065 sw
rect 48798 34063 52928 34064
tri 52928 34063 52929 34064 sw
rect 48798 34062 52929 34063
tri 52929 34062 52930 34063 sw
rect 48798 34061 52930 34062
tri 52930 34061 52931 34062 sw
rect 48798 34060 52931 34061
tri 52931 34060 52932 34061 sw
rect 48798 34059 52932 34060
tri 52932 34059 52933 34060 sw
rect 48798 34058 52933 34059
tri 52933 34058 52934 34059 sw
rect 48798 34057 52934 34058
tri 52934 34057 52935 34058 sw
rect 48798 34056 52935 34057
tri 52935 34056 52936 34057 sw
rect 48798 34055 52936 34056
tri 52936 34055 52937 34056 sw
rect 48798 34054 52937 34055
tri 52937 34054 52938 34055 sw
rect 48798 34053 52938 34054
tri 52938 34053 52939 34054 sw
rect 48798 34052 52939 34053
tri 52939 34052 52940 34053 sw
rect 48798 34051 52940 34052
tri 52940 34051 52941 34052 sw
rect 48798 34050 52941 34051
tri 52941 34050 52942 34051 sw
rect 48798 34049 52942 34050
tri 52942 34049 52943 34050 sw
rect 48798 34048 52943 34049
tri 52943 34048 52944 34049 sw
rect 48798 34047 52944 34048
tri 52944 34047 52945 34048 sw
rect 48798 34046 52945 34047
tri 52945 34046 52946 34047 sw
rect 48798 34045 52946 34046
tri 52946 34045 52947 34046 sw
rect 48798 34044 52947 34045
tri 52947 34044 52948 34045 sw
rect 48798 34043 52948 34044
tri 52948 34043 52949 34044 sw
tri 52949 34043 53237 34331 ne
rect 53237 34043 70613 34331
rect 48798 33950 52949 34043
rect 44458 33752 48504 33950
rect 42258 33682 44168 33752
rect 39997 33674 41969 33682
rect 35589 33541 39700 33674
rect 31345 33259 35441 33407
tri 35441 33259 35589 33407 sw
tri 35589 33259 35871 33541 ne
rect 35871 33377 39700 33541
tri 39700 33377 39997 33674 sw
tri 39997 33429 40242 33674 ne
rect 40242 33547 41969 33674
tri 41969 33547 42104 33682 sw
tri 42258 33547 42393 33682 ne
rect 42393 33548 44168 33682
tri 44168 33548 44372 33752 sw
tri 44458 33548 44662 33752 ne
rect 44662 33656 48504 33752
tri 48504 33656 48798 33950 sw
tri 48798 33676 49072 33950 ne
rect 49072 33755 52949 33950
tri 52949 33755 53237 34043 sw
tri 53237 33971 53309 34043 ne
rect 53309 33971 70613 34043
rect 49072 33683 53237 33755
tri 53237 33683 53309 33755 sw
tri 53309 33683 53597 33971 ne
rect 53597 33683 70613 33971
rect 49072 33676 53309 33683
rect 44662 33548 48798 33656
rect 42393 33547 44372 33548
rect 40242 33429 42104 33547
rect 35871 33259 39997 33377
rect 30340 32967 31053 33259
tri 31053 32967 31345 33259 sw
tri 31345 33223 31381 33259 ne
rect 31381 33223 35589 33259
rect 30340 32931 31345 32967
tri 31345 32931 31381 32967 sw
tri 31381 32931 31673 33223 ne
rect 31673 32977 35589 33223
tri 35589 32977 35871 33259 sw
tri 35871 33132 35998 33259 ne
rect 35998 33132 39997 33259
tri 39997 33132 40242 33377 sw
tri 40242 33228 40443 33429 ne
rect 40443 33258 42104 33429
tri 42104 33258 42393 33547 sw
tri 42393 33258 42682 33547 ne
rect 42682 33258 44372 33547
tri 44372 33258 44662 33548 sw
tri 44662 33258 44952 33548 ne
rect 44952 33382 48798 33548
tri 48798 33382 49072 33656 sw
tri 49072 33553 49195 33676 ne
rect 49195 33553 53309 33676
rect 44952 33259 49072 33382
tri 49072 33259 49195 33382 sw
tri 49195 33259 49489 33553 ne
rect 49489 33395 53309 33553
tri 53309 33395 53597 33683 sw
tri 53597 33547 53733 33683 ne
rect 53733 33547 70613 33683
rect 49489 33259 53597 33395
tri 53597 33259 53733 33395 sw
tri 53733 33288 53992 33547 ne
rect 53992 33288 70613 33547
rect 44952 33258 49195 33259
rect 40443 33228 42393 33258
tri 40443 33132 40539 33228 ne
rect 40539 33219 42393 33228
tri 42393 33219 42432 33258 sw
tri 42682 33219 42721 33258 ne
rect 42721 33220 44662 33258
tri 44662 33220 44700 33258 sw
tri 44952 33220 44990 33258 ne
rect 44990 33220 49195 33258
rect 42721 33219 44700 33220
rect 40539 33132 42432 33219
rect 31673 32931 35871 32977
rect 30340 32639 31381 32931
tri 31381 32639 31673 32931 sw
tri 31673 32928 31676 32931 ne
rect 31676 32928 35871 32931
rect 30340 32636 31673 32639
tri 31673 32636 31676 32639 sw
tri 31676 32636 31968 32928 ne
rect 31968 32850 35871 32928
tri 35871 32850 35998 32977 sw
tri 35998 32928 36202 33132 ne
rect 36202 33131 40242 33132
tri 40242 33131 40243 33132 sw
rect 36202 33130 40243 33131
tri 40243 33130 40244 33131 sw
rect 36202 33129 40244 33130
tri 40244 33129 40245 33130 sw
rect 36202 33128 40245 33129
tri 40245 33128 40246 33129 sw
rect 36202 33127 40246 33128
tri 40246 33127 40247 33128 sw
rect 36202 33126 40247 33127
tri 40247 33126 40248 33127 sw
rect 36202 33125 40248 33126
tri 40248 33125 40249 33126 sw
rect 36202 33124 40249 33125
tri 40249 33124 40250 33125 sw
rect 36202 33123 40250 33124
tri 40250 33123 40251 33124 sw
rect 36202 33122 40251 33123
tri 40251 33122 40252 33123 sw
rect 36202 33121 40252 33122
tri 40252 33121 40253 33122 sw
rect 36202 33120 40253 33121
tri 40253 33120 40254 33121 sw
rect 36202 33119 40254 33120
tri 40254 33119 40255 33120 sw
rect 36202 33118 40255 33119
tri 40255 33118 40256 33119 sw
rect 36202 33117 40256 33118
tri 40256 33117 40257 33118 sw
rect 36202 33116 40257 33117
tri 40257 33116 40258 33117 sw
rect 36202 33115 40258 33116
tri 40258 33115 40259 33116 sw
rect 36202 33114 40259 33115
tri 40259 33114 40260 33115 sw
rect 36202 33113 40260 33114
tri 40260 33113 40261 33114 sw
rect 36202 33112 40261 33113
tri 40261 33112 40262 33113 sw
rect 36202 33111 40262 33112
tri 40262 33111 40263 33112 sw
rect 36202 33110 40263 33111
tri 40263 33110 40264 33111 sw
rect 36202 33109 40264 33110
tri 40264 33109 40265 33110 sw
rect 36202 33108 40265 33109
tri 40265 33108 40266 33109 sw
rect 36202 33107 40266 33108
tri 40266 33107 40267 33108 sw
rect 36202 33106 40267 33107
tri 40267 33106 40268 33107 sw
rect 36202 33105 40268 33106
tri 40268 33105 40269 33106 sw
rect 36202 33104 40269 33105
tri 40269 33104 40270 33105 sw
rect 36202 33103 40270 33104
tri 40270 33103 40271 33104 sw
rect 36202 33102 40271 33103
tri 40271 33102 40272 33103 sw
rect 36202 33101 40272 33102
tri 40272 33101 40273 33102 sw
rect 36202 33100 40273 33101
tri 40273 33100 40274 33101 sw
rect 36202 33099 40274 33100
tri 40274 33099 40275 33100 sw
rect 36202 33098 40275 33099
tri 40275 33098 40276 33099 sw
rect 36202 33097 40276 33098
tri 40276 33097 40277 33098 sw
rect 36202 33096 40277 33097
tri 40277 33096 40278 33097 sw
rect 36202 33095 40278 33096
tri 40278 33095 40279 33096 sw
rect 36202 33094 40279 33095
tri 40279 33094 40280 33095 sw
rect 36202 33093 40280 33094
tri 40280 33093 40281 33094 sw
rect 36202 33092 40281 33093
tri 40281 33092 40282 33093 sw
rect 36202 33091 40282 33092
tri 40282 33091 40283 33092 sw
rect 36202 33090 40283 33091
tri 40283 33090 40284 33091 sw
rect 36202 33089 40284 33090
tri 40284 33089 40285 33090 sw
rect 36202 33088 40285 33089
tri 40285 33088 40286 33089 sw
rect 36202 33087 40286 33088
tri 40286 33087 40287 33088 sw
rect 36202 33086 40287 33087
tri 40287 33086 40288 33087 sw
rect 36202 33085 40288 33086
tri 40288 33085 40289 33086 sw
rect 36202 33084 40289 33085
tri 40289 33084 40290 33085 sw
rect 36202 33083 40290 33084
tri 40290 33083 40291 33084 sw
rect 36202 33082 40291 33083
tri 40291 33082 40292 33083 sw
rect 36202 33081 40292 33082
tri 40292 33081 40293 33082 sw
rect 36202 33080 40293 33081
tri 40293 33080 40294 33081 sw
rect 36202 33079 40294 33080
tri 40294 33079 40295 33080 sw
rect 36202 33078 40295 33079
tri 40295 33078 40296 33079 sw
rect 36202 33077 40296 33078
tri 40296 33077 40297 33078 sw
rect 36202 33076 40297 33077
tri 40297 33076 40298 33077 sw
rect 36202 33075 40298 33076
tri 40298 33075 40299 33076 sw
rect 36202 33074 40299 33075
tri 40299 33074 40300 33075 sw
rect 36202 33073 40300 33074
tri 40300 33073 40301 33074 sw
rect 36202 33072 40301 33073
tri 40301 33072 40302 33073 sw
rect 36202 33071 40302 33072
tri 40302 33071 40303 33072 sw
rect 36202 33070 40303 33071
tri 40303 33070 40304 33071 sw
rect 36202 33069 40304 33070
tri 40304 33069 40305 33070 sw
rect 36202 33068 40305 33069
tri 40305 33068 40306 33069 sw
rect 36202 33067 40306 33068
tri 40306 33067 40307 33068 sw
rect 36202 33066 40307 33067
tri 40307 33066 40308 33067 sw
rect 36202 33065 40308 33066
tri 40308 33065 40309 33066 sw
rect 36202 33064 40309 33065
tri 40309 33064 40310 33065 sw
rect 36202 33063 40310 33064
tri 40310 33063 40311 33064 sw
rect 36202 33062 40311 33063
tri 40311 33062 40312 33063 sw
rect 36202 33061 40312 33062
tri 40312 33061 40313 33062 sw
rect 36202 33060 40313 33061
tri 40313 33060 40314 33061 sw
rect 36202 33059 40314 33060
tri 40314 33059 40315 33060 sw
rect 36202 33058 40315 33059
tri 40315 33058 40316 33059 sw
rect 36202 33057 40316 33058
tri 40316 33057 40317 33058 sw
rect 36202 33056 40317 33057
tri 40317 33056 40318 33057 sw
rect 36202 33055 40318 33056
tri 40318 33055 40319 33056 sw
rect 36202 33054 40319 33055
tri 40319 33054 40320 33055 sw
rect 36202 33053 40320 33054
tri 40320 33053 40321 33054 sw
rect 36202 33052 40321 33053
tri 40321 33052 40322 33053 sw
rect 36202 33051 40322 33052
tri 40322 33051 40323 33052 sw
rect 36202 33050 40323 33051
tri 40323 33050 40324 33051 sw
rect 36202 33049 40324 33050
tri 40324 33049 40325 33050 sw
rect 36202 33048 40325 33049
tri 40325 33048 40326 33049 sw
rect 36202 33047 40326 33048
tri 40326 33047 40327 33048 sw
rect 36202 33046 40327 33047
tri 40327 33046 40328 33047 sw
rect 36202 33045 40328 33046
tri 40328 33045 40329 33046 sw
rect 36202 33044 40329 33045
tri 40329 33044 40330 33045 sw
rect 36202 33043 40330 33044
tri 40330 33043 40331 33044 sw
rect 36202 33042 40331 33043
tri 40331 33042 40332 33043 sw
rect 36202 33041 40332 33042
tri 40332 33041 40333 33042 sw
rect 36202 33040 40333 33041
tri 40333 33040 40334 33041 sw
rect 36202 33039 40334 33040
tri 40334 33039 40335 33040 sw
rect 36202 33038 40335 33039
tri 40335 33038 40336 33039 sw
rect 36202 33037 40336 33038
tri 40336 33037 40337 33038 sw
rect 36202 33036 40337 33037
tri 40337 33036 40338 33037 sw
rect 36202 33035 40338 33036
tri 40338 33035 40339 33036 sw
rect 36202 33034 40339 33035
tri 40339 33034 40340 33035 sw
rect 36202 33033 40340 33034
tri 40340 33033 40341 33034 sw
rect 36202 33032 40341 33033
tri 40341 33032 40342 33033 sw
rect 36202 33031 40342 33032
tri 40342 33031 40343 33032 sw
rect 36202 33030 40343 33031
tri 40343 33030 40344 33031 sw
rect 36202 33029 40344 33030
tri 40344 33029 40345 33030 sw
rect 36202 33028 40345 33029
tri 40345 33028 40346 33029 sw
rect 36202 33027 40346 33028
tri 40346 33027 40347 33028 sw
rect 36202 33026 40347 33027
tri 40347 33026 40348 33027 sw
rect 36202 33025 40348 33026
tri 40348 33025 40349 33026 sw
rect 36202 33024 40349 33025
tri 40349 33024 40350 33025 sw
rect 36202 33023 40350 33024
tri 40350 33023 40351 33024 sw
rect 36202 33022 40351 33023
tri 40351 33022 40352 33023 sw
rect 36202 33021 40352 33022
tri 40352 33021 40353 33022 sw
rect 36202 33020 40353 33021
tri 40353 33020 40354 33021 sw
rect 36202 33019 40354 33020
tri 40354 33019 40355 33020 sw
rect 36202 33018 40355 33019
tri 40355 33018 40356 33019 sw
rect 36202 33017 40356 33018
tri 40356 33017 40357 33018 sw
rect 36202 33016 40357 33017
tri 40357 33016 40358 33017 sw
rect 36202 33015 40358 33016
tri 40358 33015 40359 33016 sw
rect 36202 33014 40359 33015
tri 40359 33014 40360 33015 sw
rect 36202 33013 40360 33014
tri 40360 33013 40361 33014 sw
rect 36202 33012 40361 33013
tri 40361 33012 40362 33013 sw
rect 36202 33011 40362 33012
tri 40362 33011 40363 33012 sw
rect 36202 33010 40363 33011
tri 40363 33010 40364 33011 sw
rect 36202 33009 40364 33010
tri 40364 33009 40365 33010 sw
rect 36202 33008 40365 33009
tri 40365 33008 40366 33009 sw
rect 36202 33007 40366 33008
tri 40366 33007 40367 33008 sw
rect 36202 33006 40367 33007
tri 40367 33006 40368 33007 sw
rect 36202 33005 40368 33006
tri 40368 33005 40369 33006 sw
rect 36202 33004 40369 33005
tri 40369 33004 40370 33005 sw
rect 36202 33003 40370 33004
tri 40370 33003 40371 33004 sw
rect 36202 33002 40371 33003
tri 40371 33002 40372 33003 sw
rect 36202 33001 40372 33002
tri 40372 33001 40373 33002 sw
rect 36202 33000 40373 33001
tri 40373 33000 40374 33001 sw
rect 36202 32999 40374 33000
tri 40374 32999 40375 33000 sw
rect 36202 32998 40375 32999
tri 40375 32998 40376 32999 sw
rect 36202 32997 40376 32998
tri 40376 32997 40377 32998 sw
rect 36202 32996 40377 32997
tri 40377 32996 40378 32997 sw
rect 36202 32995 40378 32996
tri 40378 32995 40379 32996 sw
rect 36202 32994 40379 32995
tri 40379 32994 40380 32995 sw
rect 36202 32993 40380 32994
tri 40380 32993 40381 32994 sw
rect 36202 32992 40381 32993
tri 40381 32992 40382 32993 sw
rect 36202 32991 40382 32992
tri 40382 32991 40383 32992 sw
rect 36202 32990 40383 32991
tri 40383 32990 40384 32991 sw
rect 36202 32989 40384 32990
tri 40384 32989 40385 32990 sw
rect 36202 32988 40385 32989
tri 40385 32988 40386 32989 sw
rect 36202 32987 40386 32988
tri 40386 32987 40387 32988 sw
rect 36202 32986 40387 32987
tri 40387 32986 40388 32987 sw
rect 36202 32985 40388 32986
tri 40388 32985 40389 32986 sw
rect 36202 32984 40389 32985
tri 40389 32984 40390 32985 sw
rect 36202 32983 40390 32984
tri 40390 32983 40391 32984 sw
rect 36202 32982 40391 32983
tri 40391 32982 40392 32983 sw
rect 36202 32981 40392 32982
tri 40392 32981 40393 32982 sw
rect 36202 32980 40393 32981
tri 40393 32980 40394 32981 sw
rect 36202 32979 40394 32980
tri 40394 32979 40395 32980 sw
rect 36202 32978 40395 32979
tri 40395 32978 40396 32979 sw
rect 36202 32977 40396 32978
tri 40396 32977 40397 32978 sw
rect 36202 32976 40397 32977
tri 40397 32976 40398 32977 sw
rect 36202 32975 40398 32976
tri 40398 32975 40399 32976 sw
rect 36202 32974 40399 32975
tri 40399 32974 40400 32975 sw
rect 36202 32973 40400 32974
tri 40400 32973 40401 32974 sw
rect 36202 32972 40401 32973
tri 40401 32972 40402 32973 sw
rect 36202 32971 40402 32972
tri 40402 32971 40403 32972 sw
rect 36202 32970 40403 32971
tri 40403 32970 40404 32971 sw
rect 36202 32969 40404 32970
tri 40404 32969 40405 32970 sw
rect 36202 32968 40405 32969
tri 40405 32968 40406 32969 sw
rect 36202 32967 40406 32968
tri 40406 32967 40407 32968 sw
rect 36202 32966 40407 32967
tri 40407 32966 40408 32967 sw
rect 36202 32965 40408 32966
tri 40408 32965 40409 32966 sw
rect 36202 32964 40409 32965
tri 40409 32964 40410 32965 sw
rect 36202 32963 40410 32964
tri 40410 32963 40411 32964 sw
rect 36202 32962 40411 32963
tri 40411 32962 40412 32963 sw
rect 36202 32961 40412 32962
tri 40412 32961 40413 32962 sw
rect 36202 32960 40413 32961
tri 40413 32960 40414 32961 sw
rect 36202 32959 40414 32960
tri 40414 32959 40415 32960 sw
rect 36202 32958 40415 32959
tri 40415 32958 40416 32959 sw
rect 36202 32957 40416 32958
tri 40416 32957 40417 32958 sw
rect 36202 32956 40417 32957
tri 40417 32956 40418 32957 sw
rect 36202 32955 40418 32956
tri 40418 32955 40419 32956 sw
rect 36202 32954 40419 32955
tri 40419 32954 40420 32955 sw
rect 36202 32953 40420 32954
tri 40420 32953 40421 32954 sw
rect 36202 32952 40421 32953
tri 40421 32952 40422 32953 sw
rect 36202 32951 40422 32952
tri 40422 32951 40423 32952 sw
rect 36202 32950 40423 32951
tri 40423 32950 40424 32951 sw
rect 36202 32949 40424 32950
tri 40424 32949 40425 32950 sw
rect 36202 32948 40425 32949
tri 40425 32948 40426 32949 sw
rect 36202 32947 40426 32948
tri 40426 32947 40427 32948 sw
rect 36202 32946 40427 32947
tri 40427 32946 40428 32947 sw
rect 36202 32945 40428 32946
tri 40428 32945 40429 32946 sw
rect 36202 32944 40429 32945
tri 40429 32944 40430 32945 sw
rect 36202 32943 40430 32944
tri 40430 32943 40431 32944 sw
rect 36202 32942 40431 32943
tri 40431 32942 40432 32943 sw
rect 36202 32941 40432 32942
tri 40432 32941 40433 32942 sw
rect 36202 32940 40433 32941
tri 40433 32940 40434 32941 sw
rect 36202 32939 40434 32940
tri 40434 32939 40435 32940 sw
rect 36202 32938 40435 32939
tri 40435 32938 40436 32939 sw
rect 36202 32937 40436 32938
tri 40436 32937 40437 32938 sw
rect 36202 32936 40437 32937
tri 40437 32936 40438 32937 sw
rect 36202 32935 40438 32936
tri 40438 32935 40439 32936 sw
rect 36202 32934 40439 32935
tri 40439 32934 40440 32935 sw
rect 36202 32933 40440 32934
tri 40440 32933 40441 32934 sw
rect 36202 32932 40441 32933
tri 40441 32932 40442 32933 sw
rect 36202 32931 40442 32932
tri 40442 32931 40443 32932 sw
rect 36202 32930 40443 32931
tri 40443 32930 40444 32931 sw
tri 40539 32930 40741 33132 ne
rect 40741 32930 42432 33132
tri 42432 32930 42721 33219 sw
tri 42721 32930 43010 33219 ne
rect 43010 32930 44700 33219
tri 44700 32930 44990 33220 sw
tri 44990 32930 45280 33220 ne
rect 45280 32965 49195 33220
tri 49195 32965 49489 33259 sw
tri 49489 33000 49748 33259 ne
rect 49748 33000 53733 33259
tri 53733 33000 53992 33259 sw
tri 53992 33200 54080 33288 ne
rect 54080 33268 70613 33288
rect 70669 33268 71000 36132
rect 54080 33200 71000 33268
rect 45280 32930 49489 32965
rect 36202 32928 40444 32930
rect 31968 32646 35998 32850
tri 35998 32646 36202 32850 sw
tri 36202 32646 36484 32928 ne
rect 36484 32646 40444 32928
rect 31968 32636 36202 32646
rect 30340 32344 31676 32636
tri 31676 32344 31968 32636 sw
tri 31968 32635 31969 32636 ne
rect 31969 32635 36202 32636
rect 30340 32343 31968 32344
tri 31968 32343 31969 32344 sw
tri 31969 32343 32261 32635 ne
rect 32261 32364 36202 32635
tri 36202 32364 36484 32646 sw
tri 36484 32451 36679 32646 ne
rect 36679 32633 40444 32646
tri 40444 32633 40741 32930 sw
tri 40741 32920 40751 32930 ne
rect 40751 32920 42721 32930
rect 36679 32632 40741 32633
tri 40741 32632 40742 32633 sw
rect 36679 32631 40742 32632
tri 40742 32631 40743 32632 sw
rect 36679 32630 40743 32631
tri 40743 32630 40744 32631 sw
rect 36679 32629 40744 32630
tri 40744 32629 40745 32630 sw
rect 36679 32628 40745 32629
tri 40745 32628 40746 32629 sw
rect 36679 32627 40746 32628
tri 40746 32627 40747 32628 sw
rect 36679 32626 40747 32627
tri 40747 32626 40748 32627 sw
rect 36679 32625 40748 32626
tri 40748 32625 40749 32626 sw
rect 36679 32624 40749 32625
tri 40749 32624 40750 32625 sw
rect 36679 32623 40750 32624
tri 40750 32623 40751 32624 sw
tri 40751 32623 41048 32920 ne
rect 41048 32829 42721 32920
tri 42721 32829 42822 32930 sw
tri 43010 32829 43111 32930 ne
rect 43111 32830 44990 32930
tri 44990 32830 45090 32930 sw
tri 45280 32830 45380 32930 ne
rect 45380 32830 49489 32930
rect 43111 32829 45090 32830
rect 41048 32623 42822 32829
rect 36679 32451 40751 32623
rect 32261 32343 36484 32364
rect 30340 32051 31969 32343
tri 31969 32051 32261 32343 sw
tri 32261 32341 32263 32343 ne
rect 32263 32341 36484 32343
rect 30340 32049 32261 32051
tri 32261 32049 32263 32051 sw
tri 32263 32049 32555 32341 ne
rect 32555 32169 36484 32341
tri 36484 32169 36679 32364 sw
tri 36679 32169 36961 32451 ne
rect 36961 32326 40751 32451
tri 40751 32326 41048 32623 sw
tri 41048 32622 41049 32623 ne
rect 41049 32622 42822 32623
rect 36961 32325 41048 32326
tri 41048 32325 41049 32326 sw
tri 41049 32325 41346 32622 ne
rect 41346 32540 42822 32622
tri 42822 32540 43111 32829 sw
tri 43111 32540 43400 32829 ne
rect 43400 32540 45090 32829
tri 45090 32540 45380 32830 sw
tri 45380 32540 45670 32830 ne
rect 45670 32706 49489 32830
tri 49489 32706 49748 32965 sw
tri 49748 32920 49828 33000 ne
rect 49828 32920 71000 33000
rect 45670 32626 49748 32706
tri 49748 32626 49828 32706 sw
tri 49828 32705 50043 32920 ne
rect 50043 32705 70613 32920
rect 45670 32540 49828 32626
rect 41346 32325 43111 32540
rect 36961 32169 41049 32325
rect 32555 32168 36679 32169
tri 36679 32168 36680 32169 sw
tri 36961 32168 36962 32169 ne
rect 36962 32168 41049 32169
rect 32555 32049 36680 32168
rect 30340 32048 32263 32049
tri 32263 32048 32264 32049 sw
tri 32555 32048 32556 32049 ne
rect 32556 32048 36680 32049
rect 30340 31756 32264 32048
tri 32264 31756 32556 32048 sw
tri 32556 31756 32848 32048 ne
rect 32848 31886 36680 32048
tri 36680 31886 36962 32168 sw
tri 36962 31886 37244 32168 ne
rect 37244 32028 41049 32168
tri 41049 32028 41346 32325 sw
tri 41346 32183 41488 32325 ne
rect 41488 32251 43111 32325
tri 43111 32251 43400 32540 sw
tri 43400 32251 43689 32540 ne
rect 43689 32539 45380 32540
tri 45380 32539 45381 32540 sw
tri 45670 32539 45671 32540 ne
rect 45671 32539 49828 32540
rect 43689 32251 45381 32539
rect 41488 32183 43400 32251
rect 37244 31886 41346 32028
tri 41346 31886 41488 32028 sw
tri 41488 31886 41785 32183 ne
rect 41785 32175 43400 32183
tri 43400 32175 43476 32251 sw
tri 43689 32175 43765 32251 ne
rect 43765 32249 45381 32251
tri 45381 32249 45671 32539 sw
tri 45671 32249 45961 32539 ne
rect 45961 32411 49828 32539
tri 49828 32411 50043 32626 sw
tri 50043 32539 50209 32705 ne
rect 50209 32539 70613 32705
rect 45961 32249 50043 32411
rect 43765 32176 45671 32249
tri 45671 32176 45744 32249 sw
tri 45961 32176 46034 32249 ne
rect 46034 32245 50043 32249
tri 50043 32245 50209 32411 sw
tri 50209 32245 50503 32539 ne
rect 50503 32245 70613 32539
rect 46034 32180 50209 32245
tri 50209 32180 50274 32245 sw
tri 50503 32180 50568 32245 ne
rect 50568 32180 70613 32245
rect 46034 32176 50274 32180
rect 43765 32175 45744 32176
rect 41785 31886 43476 32175
tri 43476 31886 43765 32175 sw
tri 43765 31886 44054 32175 ne
rect 44054 31886 45744 32175
tri 45744 31886 46034 32176 sw
tri 46034 31886 46324 32176 ne
rect 46324 31886 50274 32176
tri 50274 31886 50568 32180 sw
tri 50568 31886 50862 32180 ne
rect 50862 31886 70613 32180
rect 32848 31756 36962 31886
rect 30340 31464 32556 31756
tri 32556 31464 32848 31756 sw
tri 32848 31755 32849 31756 ne
rect 32849 31755 36962 31756
rect 30340 31463 32848 31464
tri 32848 31463 32849 31464 sw
tri 32849 31463 33141 31755 ne
rect 33141 31604 36962 31755
tri 36962 31604 37244 31886 sw
tri 37244 31885 37245 31886 ne
rect 37245 31885 41488 31886
rect 33141 31603 37244 31604
tri 37244 31603 37245 31604 sw
tri 37245 31603 37527 31885 ne
rect 37527 31603 41488 31885
rect 33141 31463 37245 31603
rect 30340 31218 32849 31463
tri 32849 31218 33094 31463 sw
tri 33141 31218 33386 31463 ne
rect 33386 31321 37245 31463
tri 37245 31321 37527 31603 sw
tri 37527 31602 37528 31603 ne
rect 37528 31602 41488 31603
rect 33386 31320 37527 31321
tri 37527 31320 37528 31321 sw
tri 37528 31320 37810 31602 ne
rect 37810 31589 41488 31602
tri 41488 31589 41785 31886 sw
tri 41785 31589 42082 31886 ne
rect 42082 31597 43765 31886
tri 43765 31597 44054 31886 sw
tri 44054 31597 44343 31886 ne
rect 44343 31885 46034 31886
tri 46034 31885 46035 31886 sw
tri 46324 31885 46325 31886 ne
rect 46325 31885 50568 31886
rect 44343 31597 46035 31885
rect 42082 31589 44054 31597
rect 37810 31320 41785 31589
rect 33386 31218 37528 31320
rect 30340 30926 33094 31218
tri 33094 30926 33386 31218 sw
tri 33386 30926 33678 31218 ne
rect 33678 31038 37528 31218
tri 37528 31038 37810 31320 sw
tri 37810 31319 37811 31320 ne
rect 37811 31319 41785 31320
rect 33678 31037 37810 31038
tri 37810 31037 37811 31038 sw
tri 37811 31037 38093 31319 ne
rect 38093 31292 41785 31319
tri 41785 31292 42082 31589 sw
tri 42082 31535 42136 31589 ne
rect 42136 31535 44054 31589
rect 38093 31238 42082 31292
tri 42082 31238 42136 31292 sw
tri 42136 31238 42433 31535 ne
rect 42433 31483 44054 31535
tri 44054 31483 44168 31597 sw
tri 44343 31483 44457 31597 ne
rect 44457 31595 46035 31597
tri 46035 31595 46325 31885 sw
tri 46325 31595 46615 31885 ne
rect 46615 31595 50568 31885
rect 44457 31521 46325 31595
tri 46325 31521 46399 31595 sw
tri 46615 31521 46689 31595 ne
rect 46689 31592 50568 31595
tri 50568 31592 50862 31886 sw
tri 50862 31885 50863 31886 ne
rect 50863 31885 70613 31886
rect 46689 31591 50862 31592
tri 50862 31591 50863 31592 sw
tri 50863 31591 51157 31885 ne
rect 51157 31591 70613 31885
rect 46689 31521 50863 31591
rect 44457 31483 46399 31521
rect 42433 31238 44168 31483
rect 38093 31037 42136 31238
rect 33678 30926 37811 31037
rect 30340 30634 33386 30926
tri 33386 30634 33678 30926 sw
tri 33678 30925 33679 30926 ne
rect 33679 30925 37811 30926
rect 30340 30633 33678 30634
tri 33678 30633 33679 30634 sw
tri 33679 30633 33971 30925 ne
rect 33971 30755 37811 30925
tri 37811 30755 38093 31037 sw
tri 38093 30895 38235 31037 ne
rect 38235 30941 42136 31037
tri 42136 30941 42433 31238 sw
tri 42433 30941 42730 31238 ne
rect 42730 31229 44168 31238
tri 44168 31229 44422 31483 sw
tri 44457 31229 44711 31483 ne
rect 44711 31231 46399 31483
tri 46399 31231 46689 31521 sw
tri 46689 31231 46979 31521 ne
rect 46979 31297 50863 31521
tri 50863 31297 51157 31591 sw
tri 51157 31338 51410 31591 ne
rect 51410 31338 70613 31591
rect 46979 31231 51157 31297
rect 44711 31229 46689 31231
rect 42730 30941 44422 31229
rect 38235 30940 42433 30941
tri 42433 30940 42434 30941 sw
tri 42730 30940 42731 30941 ne
rect 42731 30940 44422 30941
tri 44422 30940 44711 31229 sw
tri 44711 30940 45000 31229 ne
rect 45000 31044 46689 31229
tri 46689 31044 46876 31231 sw
tri 46979 31044 47166 31231 ne
rect 47166 31044 51157 31231
tri 51157 31044 51410 31297 sw
tri 51410 31235 51513 31338 ne
rect 51513 31235 70613 31338
tri 51513 31044 51704 31235 ne
rect 51704 31044 70613 31235
rect 45000 30940 46876 31044
tri 46876 30940 46980 31044 sw
rect 38235 30895 42434 30940
rect 33971 30633 38093 30755
rect 30340 30341 33679 30633
tri 33679 30341 33971 30633 sw
tri 33971 30632 33972 30633 ne
rect 33972 30632 38093 30633
rect 30340 30340 33971 30341
tri 33971 30340 33972 30341 sw
tri 33972 30340 34264 30632 ne
rect 34264 30613 38093 30632
tri 38093 30613 38235 30755 sw
tri 38235 30613 38517 30895 ne
rect 38517 30643 42434 30895
tri 42434 30643 42731 30940 sw
tri 42731 30643 43028 30940 ne
rect 43028 30849 44711 30940
tri 44711 30849 44802 30940 sw
tri 45000 30849 45091 30940 ne
rect 45091 30851 46980 30940
tri 46980 30851 47069 30940 sw
rect 45091 30849 47069 30851
rect 43028 30643 44802 30849
rect 38517 30613 42731 30643
rect 34264 30340 38235 30613
rect 30340 30048 33972 30340
tri 33972 30048 34264 30340 sw
tri 34264 30339 34265 30340 ne
rect 34265 30339 38235 30340
rect 30340 30047 34264 30048
tri 34264 30047 34265 30048 sw
tri 34265 30047 34557 30339 ne
rect 34557 30331 38235 30339
tri 38235 30331 38517 30613 sw
tri 38517 30612 38518 30613 ne
rect 38518 30612 42731 30613
rect 34557 30330 38517 30331
tri 38517 30330 38518 30331 sw
tri 38518 30330 38800 30612 ne
rect 38800 30346 42731 30612
tri 42731 30346 43028 30643 sw
tri 43028 30642 43029 30643 ne
rect 43029 30642 44802 30643
rect 38800 30345 43028 30346
tri 43028 30345 43029 30346 sw
tri 43029 30345 43326 30642 ne
rect 43326 30560 44802 30642
tri 44802 30560 45091 30849 sw
tri 45091 30560 45380 30849 ne
rect 45380 30754 47069 30849
tri 47069 30754 47166 30851 sw
tri 47166 30754 47456 31044 ne
rect 47456 30754 51410 31044
rect 45380 30560 47166 30754
tri 47166 30560 47360 30754 sw
tri 47456 30560 47650 30754 ne
rect 47650 30750 51410 30754
tri 51410 30750 51704 31044 sw
tri 51704 30855 51893 31044 ne
rect 51893 30855 70613 31044
rect 47650 30561 51704 30750
tri 51704 30561 51893 30750 sw
tri 51893 30561 52187 30855 ne
rect 52187 30561 70613 30855
rect 47650 30560 51893 30561
rect 43326 30345 45091 30560
rect 38800 30330 43029 30345
rect 34557 30048 38518 30330
tri 38518 30048 38800 30330 sw
tri 38800 30214 38916 30330 ne
rect 38916 30214 43029 30330
rect 34557 30047 38800 30048
rect 30340 29755 34265 30047
tri 34265 29755 34557 30047 sw
tri 34557 29762 34842 30047 ne
rect 34842 29932 38800 30047
tri 38800 29932 38916 30048 sw
tri 38916 30045 39085 30214 ne
rect 39085 30048 43029 30214
tri 43029 30048 43326 30345 sw
tri 43326 30344 43327 30345 ne
rect 43327 30344 45091 30345
rect 39085 30047 43326 30048
tri 43326 30047 43327 30048 sw
tri 43327 30047 43624 30344 ne
rect 43624 30271 45091 30344
tri 45091 30271 45380 30560 sw
tri 45380 30271 45669 30560 ne
rect 45669 30336 47360 30560
tri 47360 30336 47584 30560 sw
tri 47650 30336 47874 30560 ne
rect 47874 30336 51893 30560
rect 45669 30271 47584 30336
rect 43624 30047 45380 30271
rect 39085 30045 43327 30047
tri 39085 29932 39198 30045 ne
rect 39198 29932 43327 30045
rect 34842 29762 38916 29932
rect 30340 29728 34557 29755
tri 30340 25511 34557 29728 ne
tri 34557 29470 34842 29755 sw
tri 34842 29728 34876 29762 ne
rect 34876 29728 38916 29762
rect 34557 29436 34842 29470
tri 34842 29436 34876 29470 sw
tri 34876 29436 35168 29728 ne
rect 35168 29650 38916 29728
tri 38916 29650 39198 29932 sw
tri 39198 29728 39402 29932 ne
rect 39402 29750 43327 29932
tri 43327 29750 43624 30047 sw
tri 43624 29762 43909 30047 ne
rect 43909 30046 45380 30047
tri 45380 30046 45605 30271 sw
tri 45669 30046 45894 30271 ne
rect 45894 30046 47584 30271
tri 47584 30046 47874 30336 sw
tri 47874 30046 48164 30336 ne
rect 48164 30267 51893 30336
tri 51893 30267 52187 30561 sw
tri 52187 30341 52407 30561 ne
rect 52407 30341 70613 30561
rect 48164 30047 52187 30267
tri 52187 30047 52407 30267 sw
tri 52407 30094 52654 30341 ne
rect 52654 30094 70613 30341
rect 48164 30046 52407 30047
rect 43909 29800 45605 30046
tri 45605 29800 45851 30046 sw
tri 45894 29800 46140 30046 ne
rect 46140 29800 47874 30046
rect 43909 29762 45851 29800
tri 45851 29762 45889 29800 sw
tri 46140 29762 46178 29800 ne
rect 46178 29762 47874 29800
tri 47874 29762 48158 30046 sw
tri 48164 29762 48448 30046 ne
rect 48448 29800 52407 30046
tri 52407 29800 52654 30047 sw
tri 52654 30000 52748 30094 ne
rect 52748 30056 70613 30094
rect 70669 30056 71000 32920
rect 52748 30000 71000 30056
rect 48448 29762 71000 29800
rect 39402 29728 43624 29750
rect 35168 29446 39198 29650
tri 39198 29446 39402 29650 sw
tri 39402 29446 39684 29728 ne
rect 39684 29465 43624 29728
tri 43624 29465 43909 29750 sw
tri 43909 29728 43943 29762 ne
rect 43943 29728 45889 29762
tri 45889 29728 45923 29762 sw
tri 46178 29728 46212 29762 ne
rect 46212 29728 48158 29762
rect 39684 29446 43909 29465
rect 35168 29436 39402 29446
rect 34557 29144 34876 29436
tri 34876 29144 35168 29436 sw
tri 35168 29271 35333 29436 ne
rect 35333 29271 39402 29436
rect 34557 28979 35168 29144
tri 35168 28979 35333 29144 sw
tri 35333 28979 35625 29271 ne
rect 35625 29164 39402 29271
tri 39402 29164 39684 29446 sw
tri 39684 29251 39879 29446 ne
rect 39879 29431 43909 29446
tri 43909 29431 43943 29465 sw
tri 43943 29431 44240 29728 ne
rect 44240 29439 45923 29728
tri 45923 29439 46212 29728 sw
tri 46212 29439 46501 29728 ne
rect 46501 29509 48158 29728
tri 48158 29509 48411 29762 sw
tri 48448 29509 48701 29762 ne
rect 48701 29752 71000 29762
rect 48701 29509 70613 29752
rect 46501 29439 48411 29509
rect 44240 29431 46212 29439
rect 39879 29251 43943 29431
rect 35625 28979 39684 29164
rect 34557 28978 35333 28979
tri 35333 28978 35334 28979 sw
tri 35625 28978 35626 28979 ne
rect 35626 28978 39684 28979
rect 34557 28686 35334 28978
tri 35334 28686 35626 28978 sw
tri 35626 28686 35918 28978 ne
rect 35918 28969 39684 28978
tri 39684 28969 39879 29164 sw
tri 39879 28969 40161 29251 ne
rect 40161 29134 43943 29251
tri 43943 29134 44240 29431 sw
tri 44240 29185 44486 29431 ne
rect 44486 29249 46212 29431
tri 46212 29249 46402 29439 sw
tri 46501 29249 46691 29439 ne
rect 46691 29250 48411 29439
tri 48411 29250 48670 29509 sw
tri 48701 29250 48960 29509 ne
rect 48960 29250 70613 29509
rect 46691 29249 48670 29250
rect 44486 29185 46402 29249
rect 40161 28969 44240 29134
rect 35918 28888 39879 28969
tri 39879 28888 39960 28969 sw
tri 40161 28888 40242 28969 ne
rect 40242 28888 44240 28969
tri 44240 28888 44486 29134 sw
tri 44486 28960 44711 29185 ne
rect 44711 28960 46402 29185
tri 46402 28960 46691 29249 sw
tri 46691 28960 46980 29249 ne
rect 46980 28960 48670 29249
tri 48670 28960 48960 29250 sw
tri 48960 28960 49250 29250 ne
rect 49250 28960 70613 29250
rect 35918 28686 39960 28888
rect 34557 28394 35626 28686
tri 35626 28394 35918 28686 sw
tri 35918 28685 35919 28686 ne
rect 35919 28685 39960 28686
rect 34557 28393 35918 28394
tri 35918 28393 35919 28394 sw
tri 35919 28393 36211 28685 ne
rect 36211 28606 39960 28685
tri 39960 28606 40242 28888 sw
tri 40242 28606 40524 28888 ne
rect 40524 28887 44486 28888
tri 44486 28887 44487 28888 sw
rect 40524 28886 44487 28887
tri 44487 28886 44488 28887 sw
rect 40524 28885 44488 28886
tri 44488 28885 44489 28886 sw
rect 40524 28884 44489 28885
tri 44489 28884 44490 28885 sw
rect 40524 28883 44490 28884
tri 44490 28883 44491 28884 sw
rect 40524 28882 44491 28883
tri 44491 28882 44492 28883 sw
rect 40524 28881 44492 28882
tri 44492 28881 44493 28882 sw
rect 40524 28880 44493 28881
tri 44493 28880 44494 28881 sw
rect 40524 28879 44494 28880
tri 44494 28879 44495 28880 sw
rect 40524 28878 44495 28879
tri 44495 28878 44496 28879 sw
rect 40524 28877 44496 28878
tri 44496 28877 44497 28878 sw
rect 40524 28876 44497 28877
tri 44497 28876 44498 28877 sw
rect 40524 28875 44498 28876
tri 44498 28875 44499 28876 sw
rect 40524 28874 44499 28875
tri 44499 28874 44500 28875 sw
rect 40524 28873 44500 28874
tri 44500 28873 44501 28874 sw
rect 40524 28872 44501 28873
tri 44501 28872 44502 28873 sw
rect 40524 28871 44502 28872
tri 44502 28871 44503 28872 sw
rect 40524 28870 44503 28871
tri 44503 28870 44504 28871 sw
rect 40524 28869 44504 28870
tri 44504 28869 44505 28870 sw
rect 40524 28868 44505 28869
tri 44505 28868 44506 28869 sw
rect 40524 28867 44506 28868
tri 44506 28867 44507 28868 sw
rect 40524 28866 44507 28867
tri 44507 28866 44508 28867 sw
rect 40524 28865 44508 28866
tri 44508 28865 44509 28866 sw
rect 40524 28864 44509 28865
tri 44509 28864 44510 28865 sw
rect 40524 28863 44510 28864
tri 44510 28863 44511 28864 sw
rect 40524 28862 44511 28863
tri 44511 28862 44512 28863 sw
rect 40524 28861 44512 28862
tri 44512 28861 44513 28862 sw
rect 40524 28860 44513 28861
tri 44513 28860 44514 28861 sw
rect 40524 28859 44514 28860
tri 44514 28859 44515 28860 sw
rect 40524 28858 44515 28859
tri 44515 28858 44516 28859 sw
rect 40524 28857 44516 28858
tri 44516 28857 44517 28858 sw
rect 40524 28856 44517 28857
tri 44517 28856 44518 28857 sw
rect 40524 28855 44518 28856
tri 44518 28855 44519 28856 sw
rect 40524 28854 44519 28855
tri 44519 28854 44520 28855 sw
rect 40524 28853 44520 28854
tri 44520 28853 44521 28854 sw
rect 40524 28852 44521 28853
tri 44521 28852 44522 28853 sw
rect 40524 28851 44522 28852
tri 44522 28851 44523 28852 sw
rect 40524 28850 44523 28851
tri 44523 28850 44524 28851 sw
rect 40524 28849 44524 28850
tri 44524 28849 44525 28850 sw
rect 40524 28848 44525 28849
tri 44525 28848 44526 28849 sw
rect 40524 28847 44526 28848
tri 44526 28847 44527 28848 sw
rect 40524 28846 44527 28847
tri 44527 28846 44528 28847 sw
rect 40524 28845 44528 28846
tri 44528 28845 44529 28846 sw
rect 40524 28844 44529 28845
tri 44529 28844 44530 28845 sw
rect 40524 28843 44530 28844
tri 44530 28843 44531 28844 sw
rect 40524 28842 44531 28843
tri 44531 28842 44532 28843 sw
rect 40524 28841 44532 28842
tri 44532 28841 44533 28842 sw
rect 40524 28840 44533 28841
tri 44533 28840 44534 28841 sw
rect 40524 28839 44534 28840
tri 44534 28839 44535 28840 sw
rect 40524 28838 44535 28839
tri 44535 28838 44536 28839 sw
rect 40524 28837 44536 28838
tri 44536 28837 44537 28838 sw
rect 40524 28836 44537 28837
tri 44537 28836 44538 28837 sw
rect 40524 28835 44538 28836
tri 44538 28835 44539 28836 sw
rect 40524 28834 44539 28835
tri 44539 28834 44540 28835 sw
rect 40524 28833 44540 28834
tri 44540 28833 44541 28834 sw
rect 40524 28832 44541 28833
tri 44541 28832 44542 28833 sw
rect 40524 28831 44542 28832
tri 44542 28831 44543 28832 sw
rect 40524 28830 44543 28831
tri 44543 28830 44544 28831 sw
rect 40524 28829 44544 28830
tri 44544 28829 44545 28830 sw
rect 40524 28828 44545 28829
tri 44545 28828 44546 28829 sw
rect 40524 28827 44546 28828
tri 44546 28827 44547 28828 sw
rect 40524 28826 44547 28827
tri 44547 28826 44548 28827 sw
rect 40524 28825 44548 28826
tri 44548 28825 44549 28826 sw
rect 40524 28824 44549 28825
tri 44549 28824 44550 28825 sw
rect 40524 28823 44550 28824
tri 44550 28823 44551 28824 sw
rect 40524 28822 44551 28823
tri 44551 28822 44552 28823 sw
rect 40524 28821 44552 28822
tri 44552 28821 44553 28822 sw
rect 40524 28820 44553 28821
tri 44553 28820 44554 28821 sw
rect 40524 28819 44554 28820
tri 44554 28819 44555 28820 sw
rect 40524 28818 44555 28819
tri 44555 28818 44556 28819 sw
rect 40524 28817 44556 28818
tri 44556 28817 44557 28818 sw
rect 40524 28816 44557 28817
tri 44557 28816 44558 28817 sw
rect 40524 28815 44558 28816
tri 44558 28815 44559 28816 sw
rect 40524 28814 44559 28815
tri 44559 28814 44560 28815 sw
rect 40524 28813 44560 28814
tri 44560 28813 44561 28814 sw
rect 40524 28812 44561 28813
tri 44561 28812 44562 28813 sw
rect 40524 28811 44562 28812
tri 44562 28811 44563 28812 sw
rect 40524 28810 44563 28811
tri 44563 28810 44564 28811 sw
rect 40524 28809 44564 28810
tri 44564 28809 44565 28810 sw
rect 40524 28808 44565 28809
tri 44565 28808 44566 28809 sw
rect 40524 28807 44566 28808
tri 44566 28807 44567 28808 sw
rect 40524 28806 44567 28807
tri 44567 28806 44568 28807 sw
rect 40524 28805 44568 28806
tri 44568 28805 44569 28806 sw
rect 40524 28804 44569 28805
tri 44569 28804 44570 28805 sw
rect 40524 28803 44570 28804
tri 44570 28803 44571 28804 sw
rect 40524 28802 44571 28803
tri 44571 28802 44572 28803 sw
rect 40524 28801 44572 28802
tri 44572 28801 44573 28802 sw
rect 40524 28800 44573 28801
tri 44573 28800 44574 28801 sw
rect 40524 28799 44574 28800
tri 44574 28799 44575 28800 sw
rect 40524 28798 44575 28799
tri 44575 28798 44576 28799 sw
rect 40524 28797 44576 28798
tri 44576 28797 44577 28798 sw
rect 40524 28796 44577 28797
tri 44577 28796 44578 28797 sw
rect 40524 28795 44578 28796
tri 44578 28795 44579 28796 sw
rect 40524 28794 44579 28795
tri 44579 28794 44580 28795 sw
rect 40524 28793 44580 28794
tri 44580 28793 44581 28794 sw
rect 40524 28792 44581 28793
tri 44581 28792 44582 28793 sw
rect 40524 28791 44582 28792
tri 44582 28791 44583 28792 sw
rect 40524 28790 44583 28791
tri 44583 28790 44584 28791 sw
rect 40524 28789 44584 28790
tri 44584 28789 44585 28790 sw
rect 40524 28788 44585 28789
tri 44585 28788 44586 28789 sw
rect 40524 28787 44586 28788
tri 44586 28787 44587 28788 sw
rect 40524 28786 44587 28787
tri 44587 28786 44588 28787 sw
rect 40524 28785 44588 28786
tri 44588 28785 44589 28786 sw
rect 40524 28784 44589 28785
tri 44589 28784 44590 28785 sw
rect 40524 28783 44590 28784
tri 44590 28783 44591 28784 sw
rect 40524 28782 44591 28783
tri 44591 28782 44592 28783 sw
rect 40524 28781 44592 28782
tri 44592 28781 44593 28782 sw
rect 40524 28780 44593 28781
tri 44593 28780 44594 28781 sw
rect 40524 28779 44594 28780
tri 44594 28779 44595 28780 sw
rect 40524 28778 44595 28779
tri 44595 28778 44596 28779 sw
rect 40524 28777 44596 28778
tri 44596 28777 44597 28778 sw
rect 40524 28776 44597 28777
tri 44597 28776 44598 28777 sw
rect 40524 28775 44598 28776
tri 44598 28775 44599 28776 sw
rect 40524 28774 44599 28775
tri 44599 28774 44600 28775 sw
rect 40524 28773 44600 28774
tri 44600 28773 44601 28774 sw
rect 40524 28772 44601 28773
tri 44601 28772 44602 28773 sw
rect 40524 28771 44602 28772
tri 44602 28771 44603 28772 sw
rect 40524 28770 44603 28771
tri 44603 28770 44604 28771 sw
rect 40524 28769 44604 28770
tri 44604 28769 44605 28770 sw
rect 40524 28768 44605 28769
tri 44605 28768 44606 28769 sw
rect 40524 28767 44606 28768
tri 44606 28767 44607 28768 sw
rect 40524 28766 44607 28767
tri 44607 28766 44608 28767 sw
rect 40524 28765 44608 28766
tri 44608 28765 44609 28766 sw
rect 40524 28764 44609 28765
tri 44609 28764 44610 28765 sw
rect 40524 28763 44610 28764
tri 44610 28763 44611 28764 sw
rect 40524 28762 44611 28763
tri 44611 28762 44612 28763 sw
rect 40524 28761 44612 28762
tri 44612 28761 44613 28762 sw
rect 40524 28760 44613 28761
tri 44613 28760 44614 28761 sw
rect 40524 28759 44614 28760
tri 44614 28759 44615 28760 sw
rect 40524 28758 44615 28759
tri 44615 28758 44616 28759 sw
rect 40524 28757 44616 28758
tri 44616 28757 44617 28758 sw
rect 40524 28756 44617 28757
tri 44617 28756 44618 28757 sw
rect 40524 28755 44618 28756
tri 44618 28755 44619 28756 sw
rect 40524 28754 44619 28755
tri 44619 28754 44620 28755 sw
rect 40524 28753 44620 28754
tri 44620 28753 44621 28754 sw
rect 40524 28752 44621 28753
tri 44621 28752 44622 28753 sw
rect 40524 28751 44622 28752
tri 44622 28751 44623 28752 sw
rect 40524 28750 44623 28751
tri 44623 28750 44624 28751 sw
rect 40524 28749 44624 28750
tri 44624 28749 44625 28750 sw
rect 40524 28748 44625 28749
tri 44625 28748 44626 28749 sw
rect 40524 28747 44626 28748
tri 44626 28747 44627 28748 sw
rect 40524 28746 44627 28747
tri 44627 28746 44628 28747 sw
rect 40524 28745 44628 28746
tri 44628 28745 44629 28746 sw
rect 40524 28744 44629 28745
tri 44629 28744 44630 28745 sw
rect 40524 28743 44630 28744
tri 44630 28743 44631 28744 sw
rect 40524 28742 44631 28743
tri 44631 28742 44632 28743 sw
rect 40524 28741 44632 28742
tri 44632 28741 44633 28742 sw
rect 40524 28740 44633 28741
tri 44633 28740 44634 28741 sw
rect 40524 28739 44634 28740
tri 44634 28739 44635 28740 sw
rect 40524 28738 44635 28739
tri 44635 28738 44636 28739 sw
rect 40524 28737 44636 28738
tri 44636 28737 44637 28738 sw
rect 40524 28736 44637 28737
tri 44637 28736 44638 28737 sw
rect 40524 28735 44638 28736
tri 44638 28735 44639 28736 sw
rect 40524 28734 44639 28735
tri 44639 28734 44640 28735 sw
rect 40524 28733 44640 28734
tri 44640 28733 44641 28734 sw
rect 40524 28732 44641 28733
tri 44641 28732 44642 28733 sw
rect 40524 28731 44642 28732
tri 44642 28731 44643 28732 sw
rect 40524 28730 44643 28731
tri 44643 28730 44644 28731 sw
rect 40524 28729 44644 28730
tri 44644 28729 44645 28730 sw
rect 40524 28728 44645 28729
tri 44645 28728 44646 28729 sw
rect 40524 28727 44646 28728
tri 44646 28727 44647 28728 sw
rect 40524 28726 44647 28727
tri 44647 28726 44648 28727 sw
rect 40524 28725 44648 28726
tri 44648 28725 44649 28726 sw
rect 40524 28724 44649 28725
tri 44649 28724 44650 28725 sw
rect 40524 28723 44650 28724
tri 44650 28723 44651 28724 sw
rect 40524 28722 44651 28723
tri 44651 28722 44652 28723 sw
rect 40524 28721 44652 28722
tri 44652 28721 44653 28722 sw
rect 40524 28720 44653 28721
tri 44653 28720 44654 28721 sw
rect 40524 28719 44654 28720
tri 44654 28719 44655 28720 sw
rect 40524 28718 44655 28719
tri 44655 28718 44656 28719 sw
rect 40524 28717 44656 28718
tri 44656 28717 44657 28718 sw
rect 40524 28716 44657 28717
tri 44657 28716 44658 28717 sw
rect 40524 28715 44658 28716
tri 44658 28715 44659 28716 sw
rect 40524 28714 44659 28715
tri 44659 28714 44660 28715 sw
rect 40524 28713 44660 28714
tri 44660 28713 44661 28714 sw
rect 40524 28712 44661 28713
tri 44661 28712 44662 28713 sw
rect 40524 28711 44662 28712
tri 44662 28711 44663 28712 sw
rect 40524 28710 44663 28711
tri 44663 28710 44664 28711 sw
rect 40524 28709 44664 28710
tri 44664 28709 44665 28710 sw
rect 40524 28708 44665 28709
tri 44665 28708 44666 28709 sw
rect 40524 28707 44666 28708
tri 44666 28707 44667 28708 sw
rect 40524 28706 44667 28707
tri 44667 28706 44668 28707 sw
rect 40524 28705 44668 28706
tri 44668 28705 44669 28706 sw
rect 40524 28704 44669 28705
tri 44669 28704 44670 28705 sw
rect 40524 28703 44670 28704
tri 44670 28703 44671 28704 sw
rect 40524 28702 44671 28703
tri 44671 28702 44672 28703 sw
rect 40524 28701 44672 28702
tri 44672 28701 44673 28702 sw
rect 40524 28700 44673 28701
tri 44673 28700 44674 28701 sw
rect 40524 28699 44674 28700
tri 44674 28699 44675 28700 sw
rect 40524 28698 44675 28699
tri 44675 28698 44676 28699 sw
rect 40524 28697 44676 28698
tri 44676 28697 44677 28698 sw
rect 40524 28696 44677 28697
tri 44677 28696 44678 28697 sw
rect 40524 28695 44678 28696
tri 44678 28695 44679 28696 sw
rect 40524 28694 44679 28695
tri 44679 28694 44680 28695 sw
rect 40524 28693 44680 28694
tri 44680 28693 44681 28694 sw
rect 40524 28692 44681 28693
tri 44681 28692 44682 28693 sw
rect 40524 28691 44682 28692
tri 44682 28691 44683 28692 sw
rect 40524 28690 44683 28691
tri 44683 28690 44684 28691 sw
rect 40524 28689 44684 28690
tri 44684 28689 44685 28690 sw
rect 40524 28688 44685 28689
tri 44685 28688 44686 28689 sw
rect 40524 28687 44686 28688
tri 44686 28687 44687 28688 sw
rect 40524 28686 44687 28687
tri 44687 28686 44688 28687 sw
tri 44711 28686 44985 28960 ne
rect 44985 28686 46691 28960
tri 46691 28686 46965 28960 sw
tri 46980 28686 47254 28960 ne
rect 47254 28686 48960 28960
tri 48960 28686 49234 28960 sw
tri 49250 28686 49524 28960 ne
rect 49524 28686 70613 28960
rect 40524 28606 44688 28686
rect 36211 28393 40242 28606
rect 34557 28101 35919 28393
tri 35919 28101 36211 28393 sw
tri 36211 28392 36212 28393 ne
rect 36212 28392 40242 28393
rect 34557 28100 36211 28101
tri 36211 28100 36212 28101 sw
tri 36212 28100 36504 28392 ne
rect 36504 28324 40242 28392
tri 40242 28324 40524 28606 sw
tri 40524 28402 40728 28606 ne
rect 40728 28402 44688 28606
rect 36504 28120 40524 28324
tri 40524 28120 40728 28324 sw
tri 40728 28209 40921 28402 ne
rect 40921 28389 44688 28402
tri 44688 28389 44985 28686 sw
tri 44985 28662 45009 28686 ne
rect 45009 28662 46965 28686
rect 40921 28365 44985 28389
tri 44985 28365 45009 28389 sw
tri 45009 28365 45306 28662 ne
rect 45306 28485 46965 28662
tri 46965 28485 47166 28686 sw
tri 47254 28580 47360 28686 ne
rect 47360 28580 49234 28686
rect 45306 28365 47166 28485
rect 40921 28209 45009 28365
rect 36504 28100 40728 28120
rect 34557 27808 36212 28100
tri 36212 27808 36504 28100 sw
tri 36504 28099 36505 28100 ne
rect 36505 28099 40728 28100
rect 34557 27807 36504 27808
tri 36504 27807 36505 27808 sw
tri 36505 27807 36797 28099 ne
rect 36797 27927 40728 28099
tri 40728 27927 40921 28120 sw
tri 40921 27927 41203 28209 ne
rect 41203 28068 45009 28209
tri 45009 28068 45306 28365 sw
tri 45306 28238 45433 28365 ne
rect 45433 28291 47166 28365
tri 47166 28291 47360 28485 sw
tri 47360 28291 47649 28580 ne
rect 47649 28579 49234 28580
tri 49234 28579 49341 28686 sw
tri 49524 28579 49631 28686 ne
rect 49631 28579 70613 28686
rect 47649 28291 49341 28579
rect 45433 28238 47360 28291
rect 41203 27941 45306 28068
tri 45306 27941 45433 28068 sw
tri 45433 27941 45730 28238 ne
rect 45730 28002 47360 28238
tri 47360 28002 47649 28291 sw
tri 47649 28002 47938 28291 ne
rect 47938 28289 49341 28291
tri 49341 28289 49631 28579 sw
tri 49631 28289 49921 28579 ne
rect 49921 28289 70613 28579
rect 47938 28223 49631 28289
tri 49631 28223 49697 28289 sw
tri 49921 28223 49987 28289 ne
rect 49987 28223 70613 28289
rect 47938 28002 49697 28223
rect 45730 27941 47649 28002
rect 41203 27927 45433 27941
rect 36797 27807 40921 27927
rect 34557 27515 36505 27807
tri 36505 27515 36797 27807 sw
tri 36797 27757 36847 27807 ne
rect 36847 27757 40921 27807
rect 34557 27465 36797 27515
tri 36797 27465 36847 27515 sw
tri 36847 27465 37139 27757 ne
rect 37139 27645 40921 27757
tri 40921 27645 41203 27927 sw
tri 41203 27925 41205 27927 ne
rect 41205 27925 45433 27927
rect 37139 27643 41203 27645
tri 41203 27643 41205 27645 sw
tri 41205 27643 41487 27925 ne
rect 41487 27644 45433 27925
tri 45433 27644 45730 27941 sw
tri 45730 27940 45731 27941 ne
rect 45731 27940 47649 27941
rect 41487 27643 45730 27644
tri 45730 27643 45731 27644 sw
tri 45731 27643 46028 27940 ne
rect 46028 27932 47649 27940
tri 47649 27932 47719 28002 sw
tri 47938 27932 48008 28002 ne
rect 48008 27933 49697 28002
tri 49697 27933 49987 28223 sw
tri 49987 27933 50277 28223 ne
rect 50277 27933 70613 28223
rect 48008 27932 49987 27933
rect 46028 27643 47719 27932
tri 47719 27643 48008 27932 sw
tri 48008 27643 48297 27932 ne
rect 48297 27643 49987 27932
tri 49987 27643 50277 27933 sw
tri 50277 27643 50567 27933 ne
rect 50567 27643 70613 27933
rect 37139 27642 41205 27643
tri 41205 27642 41206 27643 sw
tri 41487 27642 41488 27643 ne
rect 41488 27642 45731 27643
rect 37139 27465 41206 27642
rect 34557 27173 36847 27465
tri 36847 27173 37139 27465 sw
tri 37139 27464 37140 27465 ne
rect 37140 27464 41206 27465
rect 34557 27172 37139 27173
tri 37139 27172 37140 27173 sw
tri 37140 27172 37432 27464 ne
rect 37432 27360 41206 27464
tri 41206 27360 41488 27642 sw
tri 41488 27360 41770 27642 ne
rect 41770 27360 45731 27642
rect 37432 27172 41488 27360
rect 34557 26880 37140 27172
tri 37140 26880 37432 27172 sw
tri 37432 27024 37580 27172 ne
rect 37580 27078 41488 27172
tri 41488 27078 41770 27360 sw
tri 41770 27161 41969 27360 ne
rect 41969 27346 45731 27360
tri 45731 27346 46028 27643 sw
tri 46028 27346 46325 27643 ne
rect 46325 27354 48008 27643
tri 48008 27354 48297 27643 sw
tri 48297 27354 48586 27643 ne
rect 48586 27642 50277 27643
tri 50277 27642 50278 27643 sw
tri 50567 27642 50568 27643 ne
rect 50568 27642 70613 27643
rect 48586 27354 50278 27642
rect 46325 27346 48297 27354
rect 41969 27161 46028 27346
rect 37580 27024 41770 27078
rect 34557 26732 37432 26880
tri 37432 26732 37580 26880 sw
tri 37580 26877 37727 27024 ne
rect 37727 26879 41770 27024
tri 41770 26879 41969 27078 sw
tri 41969 26879 42251 27161 ne
rect 42251 27049 46028 27161
tri 46028 27049 46325 27346 sw
tri 46325 27278 46393 27346 ne
rect 46393 27278 48297 27346
rect 42251 26981 46325 27049
tri 46325 26981 46393 27049 sw
tri 46393 26981 46690 27278 ne
rect 46690 27240 48297 27278
tri 48297 27240 48411 27354 sw
tri 48586 27240 48700 27354 ne
rect 48700 27352 50278 27354
tri 50278 27352 50568 27642 sw
tri 50568 27352 50858 27642 ne
rect 50858 27352 70613 27642
rect 48700 27270 50568 27352
tri 50568 27270 50650 27352 sw
tri 50858 27270 50940 27352 ne
rect 50940 27270 70613 27352
rect 48700 27240 50650 27270
rect 46690 26981 48411 27240
rect 42251 26879 46393 26981
rect 37727 26877 41969 26879
rect 34557 26731 37580 26732
tri 37580 26731 37581 26732 sw
rect 34557 26730 37581 26731
tri 37581 26730 37582 26731 sw
rect 34557 26729 37582 26730
tri 37582 26729 37583 26730 sw
rect 34557 26728 37583 26729
tri 37583 26728 37584 26729 sw
rect 34557 26727 37584 26728
tri 37584 26727 37585 26728 sw
rect 34557 26726 37585 26727
tri 37585 26726 37586 26727 sw
rect 34557 26725 37586 26726
tri 37586 26725 37587 26726 sw
rect 34557 26724 37587 26725
tri 37587 26724 37588 26725 sw
rect 34557 26723 37588 26724
tri 37588 26723 37589 26724 sw
rect 34557 26722 37589 26723
tri 37589 26722 37590 26723 sw
rect 34557 26721 37590 26722
tri 37590 26721 37591 26722 sw
rect 34557 26720 37591 26721
tri 37591 26720 37592 26721 sw
rect 34557 26719 37592 26720
tri 37592 26719 37593 26720 sw
rect 34557 26718 37593 26719
tri 37593 26718 37594 26719 sw
rect 34557 26717 37594 26718
tri 37594 26717 37595 26718 sw
rect 34557 26716 37595 26717
tri 37595 26716 37596 26717 sw
rect 34557 26715 37596 26716
tri 37596 26715 37597 26716 sw
rect 34557 26714 37597 26715
tri 37597 26714 37598 26715 sw
rect 34557 26713 37598 26714
tri 37598 26713 37599 26714 sw
rect 34557 26712 37599 26713
tri 37599 26712 37600 26713 sw
rect 34557 26711 37600 26712
tri 37600 26711 37601 26712 sw
rect 34557 26710 37601 26711
tri 37601 26710 37602 26711 sw
rect 34557 26709 37602 26710
tri 37602 26709 37603 26710 sw
rect 34557 26708 37603 26709
tri 37603 26708 37604 26709 sw
rect 34557 26707 37604 26708
tri 37604 26707 37605 26708 sw
rect 34557 26706 37605 26707
tri 37605 26706 37606 26707 sw
rect 34557 26705 37606 26706
tri 37606 26705 37607 26706 sw
rect 34557 26704 37607 26705
tri 37607 26704 37608 26705 sw
rect 34557 26703 37608 26704
tri 37608 26703 37609 26704 sw
rect 34557 26702 37609 26703
tri 37609 26702 37610 26703 sw
rect 34557 26701 37610 26702
tri 37610 26701 37611 26702 sw
rect 34557 26700 37611 26701
tri 37611 26700 37612 26701 sw
rect 34557 26699 37612 26700
tri 37612 26699 37613 26700 sw
rect 34557 26698 37613 26699
tri 37613 26698 37614 26699 sw
rect 34557 26697 37614 26698
tri 37614 26697 37615 26698 sw
rect 34557 26696 37615 26697
tri 37615 26696 37616 26697 sw
rect 34557 26695 37616 26696
tri 37616 26695 37617 26696 sw
rect 34557 26694 37617 26695
tri 37617 26694 37618 26695 sw
rect 34557 26693 37618 26694
tri 37618 26693 37619 26694 sw
rect 34557 26692 37619 26693
tri 37619 26692 37620 26693 sw
rect 34557 26691 37620 26692
tri 37620 26691 37621 26692 sw
rect 34557 26690 37621 26691
tri 37621 26690 37622 26691 sw
rect 34557 26689 37622 26690
tri 37622 26689 37623 26690 sw
rect 34557 26688 37623 26689
tri 37623 26688 37624 26689 sw
rect 34557 26687 37624 26688
tri 37624 26687 37625 26688 sw
rect 34557 26686 37625 26687
tri 37625 26686 37626 26687 sw
rect 34557 26685 37626 26686
tri 37626 26685 37627 26686 sw
rect 34557 26684 37627 26685
tri 37627 26684 37628 26685 sw
rect 34557 26683 37628 26684
tri 37628 26683 37629 26684 sw
rect 34557 26682 37629 26683
tri 37629 26682 37630 26683 sw
rect 34557 26681 37630 26682
tri 37630 26681 37631 26682 sw
rect 34557 26680 37631 26681
tri 37631 26680 37632 26681 sw
rect 34557 26679 37632 26680
tri 37632 26679 37633 26680 sw
rect 34557 26678 37633 26679
tri 37633 26678 37634 26679 sw
rect 34557 26677 37634 26678
tri 37634 26677 37635 26678 sw
rect 34557 26676 37635 26677
tri 37635 26676 37636 26677 sw
rect 34557 26675 37636 26676
tri 37636 26675 37637 26676 sw
rect 34557 26674 37637 26675
tri 37637 26674 37638 26675 sw
rect 34557 26673 37638 26674
tri 37638 26673 37639 26674 sw
rect 34557 26672 37639 26673
tri 37639 26672 37640 26673 sw
rect 34557 26671 37640 26672
tri 37640 26671 37641 26672 sw
rect 34557 26670 37641 26671
tri 37641 26670 37642 26671 sw
rect 34557 26669 37642 26670
tri 37642 26669 37643 26670 sw
rect 34557 26668 37643 26669
tri 37643 26668 37644 26669 sw
rect 34557 26667 37644 26668
tri 37644 26667 37645 26668 sw
rect 34557 26666 37645 26667
tri 37645 26666 37646 26667 sw
rect 34557 26665 37646 26666
tri 37646 26665 37647 26666 sw
rect 34557 26664 37647 26665
tri 37647 26664 37648 26665 sw
rect 34557 26663 37648 26664
tri 37648 26663 37649 26664 sw
rect 34557 26662 37649 26663
tri 37649 26662 37650 26663 sw
rect 34557 26661 37650 26662
tri 37650 26661 37651 26662 sw
rect 34557 26660 37651 26661
tri 37651 26660 37652 26661 sw
rect 34557 26659 37652 26660
tri 37652 26659 37653 26660 sw
rect 34557 26658 37653 26659
tri 37653 26658 37654 26659 sw
rect 34557 26657 37654 26658
tri 37654 26657 37655 26658 sw
rect 34557 26656 37655 26657
tri 37655 26656 37656 26657 sw
rect 34557 26655 37656 26656
tri 37656 26655 37657 26656 sw
rect 34557 26654 37657 26655
tri 37657 26654 37658 26655 sw
rect 34557 26653 37658 26654
tri 37658 26653 37659 26654 sw
rect 34557 26652 37659 26653
tri 37659 26652 37660 26653 sw
rect 34557 26651 37660 26652
tri 37660 26651 37661 26652 sw
rect 34557 26650 37661 26651
tri 37661 26650 37662 26651 sw
rect 34557 26649 37662 26650
tri 37662 26649 37663 26650 sw
rect 34557 26648 37663 26649
tri 37663 26648 37664 26649 sw
rect 34557 26647 37664 26648
tri 37664 26647 37665 26648 sw
rect 34557 26646 37665 26647
tri 37665 26646 37666 26647 sw
rect 34557 26645 37666 26646
tri 37666 26645 37667 26646 sw
rect 34557 26644 37667 26645
tri 37667 26644 37668 26645 sw
rect 34557 26643 37668 26644
tri 37668 26643 37669 26644 sw
rect 34557 26642 37669 26643
tri 37669 26642 37670 26643 sw
rect 34557 26641 37670 26642
tri 37670 26641 37671 26642 sw
rect 34557 26640 37671 26641
tri 37671 26640 37672 26641 sw
rect 34557 26639 37672 26640
tri 37672 26639 37673 26640 sw
rect 34557 26638 37673 26639
tri 37673 26638 37674 26639 sw
rect 34557 26637 37674 26638
tri 37674 26637 37675 26638 sw
rect 34557 26636 37675 26637
tri 37675 26636 37676 26637 sw
rect 34557 26635 37676 26636
tri 37676 26635 37677 26636 sw
rect 34557 26634 37677 26635
tri 37677 26634 37678 26635 sw
rect 34557 26633 37678 26634
tri 37678 26633 37679 26634 sw
rect 34557 26632 37679 26633
tri 37679 26632 37680 26633 sw
rect 34557 26631 37680 26632
tri 37680 26631 37681 26632 sw
rect 34557 26630 37681 26631
tri 37681 26630 37682 26631 sw
rect 34557 26629 37682 26630
tri 37682 26629 37683 26630 sw
rect 34557 26628 37683 26629
tri 37683 26628 37684 26629 sw
rect 34557 26627 37684 26628
tri 37684 26627 37685 26628 sw
rect 34557 26626 37685 26627
tri 37685 26626 37686 26627 sw
rect 34557 26625 37686 26626
tri 37686 26625 37687 26626 sw
rect 34557 26624 37687 26625
tri 37687 26624 37688 26625 sw
rect 34557 26623 37688 26624
tri 37688 26623 37689 26624 sw
rect 34557 26622 37689 26623
tri 37689 26622 37690 26623 sw
rect 34557 26621 37690 26622
tri 37690 26621 37691 26622 sw
rect 34557 26620 37691 26621
tri 37691 26620 37692 26621 sw
rect 34557 26619 37692 26620
tri 37692 26619 37693 26620 sw
rect 34557 26618 37693 26619
tri 37693 26618 37694 26619 sw
rect 34557 26617 37694 26618
tri 37694 26617 37695 26618 sw
rect 34557 26616 37695 26617
tri 37695 26616 37696 26617 sw
rect 34557 26615 37696 26616
tri 37696 26615 37697 26616 sw
rect 34557 26614 37697 26615
tri 37697 26614 37698 26615 sw
rect 34557 26613 37698 26614
tri 37698 26613 37699 26614 sw
rect 34557 26612 37699 26613
tri 37699 26612 37700 26613 sw
rect 34557 26611 37700 26612
tri 37700 26611 37701 26612 sw
rect 34557 26610 37701 26611
tri 37701 26610 37702 26611 sw
rect 34557 26609 37702 26610
tri 37702 26609 37703 26610 sw
rect 34557 26608 37703 26609
tri 37703 26608 37704 26609 sw
rect 34557 26607 37704 26608
tri 37704 26607 37705 26608 sw
rect 34557 26606 37705 26607
tri 37705 26606 37706 26607 sw
rect 34557 26605 37706 26606
tri 37706 26605 37707 26606 sw
rect 34557 26604 37707 26605
tri 37707 26604 37708 26605 sw
rect 34557 26603 37708 26604
tri 37708 26603 37709 26604 sw
rect 34557 26602 37709 26603
tri 37709 26602 37710 26603 sw
rect 34557 26601 37710 26602
tri 37710 26601 37711 26602 sw
rect 34557 26600 37711 26601
tri 37711 26600 37712 26601 sw
rect 34557 26599 37712 26600
tri 37712 26599 37713 26600 sw
rect 34557 26598 37713 26599
tri 37713 26598 37714 26599 sw
rect 34557 26597 37714 26598
tri 37714 26597 37715 26598 sw
rect 34557 26596 37715 26597
tri 37715 26596 37716 26597 sw
rect 34557 26595 37716 26596
tri 37716 26595 37717 26596 sw
rect 34557 26594 37717 26595
tri 37717 26594 37718 26595 sw
rect 34557 26593 37718 26594
tri 37718 26593 37719 26594 sw
rect 34557 26592 37719 26593
tri 37719 26592 37720 26593 sw
rect 34557 26591 37720 26592
tri 37720 26591 37721 26592 sw
rect 34557 26590 37721 26591
tri 37721 26590 37722 26591 sw
rect 34557 26589 37722 26590
tri 37722 26589 37723 26590 sw
rect 34557 26588 37723 26589
tri 37723 26588 37724 26589 sw
rect 34557 26587 37724 26588
tri 37724 26587 37725 26588 sw
rect 34557 26586 37725 26587
tri 37725 26586 37726 26587 sw
rect 34557 26585 37726 26586
tri 37726 26585 37727 26586 sw
tri 37727 26585 38019 26877 ne
rect 38019 26597 41969 26877
tri 41969 26597 42251 26879 sw
tri 42251 26877 42253 26879 ne
rect 42253 26877 46393 26879
rect 38019 26595 42251 26597
tri 42251 26595 42253 26597 sw
tri 42253 26595 42535 26877 ne
rect 42535 26684 46393 26877
tri 46393 26684 46690 26981 sw
tri 46690 26878 46793 26981 ne
rect 46793 26980 48411 26981
tri 48411 26980 48671 27240 sw
tri 48700 26980 48960 27240 ne
rect 48960 26980 50650 27240
tri 50650 26980 50940 27270 sw
tri 50940 26980 51230 27270 ne
rect 51230 26980 70613 27270
rect 46793 26878 48671 26980
rect 42535 26683 46690 26684
tri 46690 26683 46691 26684 sw
rect 42535 26682 46691 26683
tri 46691 26682 46692 26683 sw
tri 46793 26682 46989 26878 ne
rect 46989 26800 48671 26878
tri 48671 26800 48851 26980 sw
tri 48960 26800 49140 26980 ne
rect 49140 26800 50940 26980
tri 50940 26800 51120 26980 sw
tri 51230 26800 51410 26980 ne
rect 51410 26888 70613 26980
rect 70669 26888 71000 29752
rect 51410 26800 71000 26888
rect 46989 26682 48851 26800
rect 42535 26595 46692 26682
rect 38019 26594 42253 26595
tri 42253 26594 42254 26595 sw
tri 42535 26594 42536 26595 ne
rect 42536 26594 46692 26595
rect 38019 26585 42254 26594
rect 34557 26584 37727 26585
tri 37727 26584 37728 26585 sw
tri 38019 26584 38020 26585 ne
rect 38020 26584 42254 26585
rect 34557 26292 37728 26584
tri 37728 26292 38020 26584 sw
tri 38020 26292 38312 26584 ne
rect 38312 26312 42254 26584
tri 42254 26312 42536 26594 sw
tri 42536 26312 42818 26594 ne
rect 42818 26385 46692 26594
tri 46692 26385 46989 26682 sw
tri 46989 26385 47286 26682 ne
rect 47286 26600 48851 26682
tri 48851 26600 49051 26800 sw
tri 49140 26600 49340 26800 ne
rect 49340 26600 51120 26800
tri 51120 26600 51320 26800 sw
rect 47286 26385 49051 26600
rect 42818 26312 46989 26385
rect 38312 26292 42536 26312
rect 34557 26000 38020 26292
tri 38020 26000 38312 26292 sw
tri 38312 26071 38533 26292 ne
rect 38533 26071 42536 26292
rect 34557 25779 38312 26000
tri 38312 25779 38533 26000 sw
tri 38533 25779 38825 26071 ne
rect 38825 26030 42536 26071
tri 42536 26030 42818 26312 sw
tri 42818 26051 43079 26312 ne
rect 43079 26088 46989 26312
tri 46989 26088 47286 26385 sw
tri 47286 26088 47583 26385 ne
rect 47583 26311 49051 26385
tri 49051 26311 49340 26600 sw
tri 49340 26311 49629 26600 ne
rect 49629 26311 71000 26600
rect 47583 26088 49340 26311
rect 43079 26051 47286 26088
rect 38825 25779 42818 26030
rect 34557 25688 38533 25779
tri 38533 25688 38624 25779 sw
tri 38825 25688 38916 25779 ne
rect 38916 25769 42818 25779
tri 42818 25769 43079 26030 sw
tri 43079 25769 43361 26051 ne
rect 43361 25791 47286 26051
tri 47286 25791 47583 26088 sw
tri 47583 26081 47590 26088 ne
rect 47590 26081 49340 26088
rect 43361 25784 47583 25791
tri 47583 25784 47590 25791 sw
tri 47590 25784 47887 26081 ne
rect 47887 26022 49340 26081
tri 49340 26022 49629 26311 sw
tri 49629 26022 49918 26311 ne
rect 49918 26022 71000 26311
rect 47887 25784 49629 26022
rect 43361 25769 47590 25784
rect 38916 25688 43079 25769
tri 43079 25688 43160 25769 sw
tri 43361 25768 43362 25769 ne
rect 43362 25768 47590 25769
rect 34557 25511 38624 25688
tri 34557 21444 38624 25511 ne
tri 38624 25396 38916 25688 sw
tri 38916 25396 39208 25688 ne
rect 39208 25486 43160 25688
tri 43160 25486 43362 25688 sw
tri 43362 25486 43644 25768 ne
rect 43644 25487 47590 25768
tri 47590 25487 47887 25784 sw
tri 47887 25783 47888 25784 ne
rect 47888 25783 49629 25784
rect 43644 25486 47887 25487
tri 47887 25486 47888 25487 sw
tri 47888 25486 48185 25783 ne
rect 48185 25775 49629 25783
tri 49629 25775 49876 26022 sw
tri 49918 25775 50165 26022 ne
rect 50165 25775 71000 26022
rect 48185 25486 49876 25775
tri 49876 25486 50165 25775 sw
tri 50165 25486 50454 25775 ne
rect 50454 25486 71000 25775
rect 39208 25396 43362 25486
rect 38624 25104 38916 25396
tri 38916 25104 39208 25396 sw
tri 39208 25209 39395 25396 ne
rect 39395 25209 43362 25396
rect 38624 24917 39208 25104
tri 39208 24917 39395 25104 sw
tri 39395 24917 39687 25209 ne
rect 39687 25204 43362 25209
tri 43362 25204 43644 25486 sw
tri 43644 25485 43645 25486 ne
rect 43645 25485 47888 25486
rect 39687 25203 43644 25204
tri 43644 25203 43645 25204 sw
tri 43645 25203 43927 25485 ne
rect 43927 25203 47888 25485
rect 39687 24921 43645 25203
tri 43645 24921 43927 25203 sw
tri 43927 25199 43931 25203 ne
rect 43931 25199 47888 25203
rect 39687 24917 43927 24921
tri 43927 24917 43931 24921 sw
tri 43931 24917 44213 25199 ne
rect 44213 25189 47888 25199
tri 47888 25189 48185 25486 sw
tri 48185 25298 48373 25486 ne
rect 48373 25298 50165 25486
rect 44213 25001 48185 25189
tri 48185 25001 48373 25189 sw
tri 48373 25001 48670 25298 ne
rect 48670 25200 50165 25298
tri 50165 25200 50451 25486 sw
tri 50454 25200 50740 25486 ne
rect 50740 25200 71000 25486
rect 48670 25001 50451 25200
rect 44213 24917 48373 25001
rect 38624 24625 39395 24917
tri 39395 24625 39687 24917 sw
tri 39687 24735 39869 24917 ne
rect 39869 24735 43931 24917
rect 38624 24443 39687 24625
tri 39687 24443 39869 24625 sw
tri 39869 24443 40161 24735 ne
rect 40161 24635 43931 24735
tri 43931 24635 44213 24917 sw
tri 44213 24644 44486 24917 ne
rect 44486 24704 48373 24917
tri 48373 24704 48670 25001 sw
tri 48670 24916 48755 25001 ne
rect 48755 25000 50451 25001
tri 50451 25000 50651 25200 sw
rect 48755 24916 71000 25000
rect 44486 24644 48670 24704
rect 40161 24443 44213 24635
rect 38624 24442 39869 24443
tri 39869 24442 39870 24443 sw
tri 40161 24442 40162 24443 ne
rect 40162 24442 44213 24443
rect 38624 24150 39870 24442
tri 39870 24150 40162 24442 sw
tri 40162 24150 40454 24442 ne
rect 40454 24362 44213 24442
tri 44213 24362 44486 24635 sw
tri 44486 24362 44768 24644 ne
rect 44768 24619 48670 24644
tri 48670 24619 48755 24704 sw
tri 48755 24702 48969 24916 ne
rect 48969 24906 71000 24916
rect 48969 24702 70613 24906
rect 44768 24618 48755 24619
tri 48755 24618 48756 24619 sw
rect 44768 24617 48756 24618
tri 48756 24617 48757 24618 sw
rect 44768 24616 48757 24617
tri 48757 24616 48758 24617 sw
rect 44768 24615 48758 24616
tri 48758 24615 48759 24616 sw
rect 44768 24614 48759 24615
tri 48759 24614 48760 24615 sw
rect 44768 24613 48760 24614
tri 48760 24613 48761 24614 sw
rect 44768 24612 48761 24613
tri 48761 24612 48762 24613 sw
rect 44768 24611 48762 24612
tri 48762 24611 48763 24612 sw
rect 44768 24610 48763 24611
tri 48763 24610 48764 24611 sw
rect 44768 24609 48764 24610
tri 48764 24609 48765 24610 sw
rect 44768 24608 48765 24609
tri 48765 24608 48766 24609 sw
rect 44768 24607 48766 24608
tri 48766 24607 48767 24608 sw
rect 44768 24606 48767 24607
tri 48767 24606 48768 24607 sw
rect 44768 24605 48768 24606
tri 48768 24605 48769 24606 sw
rect 44768 24604 48769 24605
tri 48769 24604 48770 24605 sw
rect 44768 24603 48770 24604
tri 48770 24603 48771 24604 sw
rect 44768 24602 48771 24603
tri 48771 24602 48772 24603 sw
rect 44768 24601 48772 24602
tri 48772 24601 48773 24602 sw
rect 44768 24600 48773 24601
tri 48773 24600 48774 24601 sw
rect 44768 24599 48774 24600
tri 48774 24599 48775 24600 sw
rect 44768 24598 48775 24599
tri 48775 24598 48776 24599 sw
rect 44768 24597 48776 24598
tri 48776 24597 48777 24598 sw
rect 44768 24596 48777 24597
tri 48777 24596 48778 24597 sw
rect 44768 24595 48778 24596
tri 48778 24595 48779 24596 sw
rect 44768 24594 48779 24595
tri 48779 24594 48780 24595 sw
rect 44768 24593 48780 24594
tri 48780 24593 48781 24594 sw
rect 44768 24592 48781 24593
tri 48781 24592 48782 24593 sw
rect 44768 24591 48782 24592
tri 48782 24591 48783 24592 sw
rect 44768 24590 48783 24591
tri 48783 24590 48784 24591 sw
rect 44768 24589 48784 24590
tri 48784 24589 48785 24590 sw
rect 44768 24588 48785 24589
tri 48785 24588 48786 24589 sw
rect 44768 24587 48786 24588
tri 48786 24587 48787 24588 sw
rect 44768 24586 48787 24587
tri 48787 24586 48788 24587 sw
rect 44768 24585 48788 24586
tri 48788 24585 48789 24586 sw
rect 44768 24584 48789 24585
tri 48789 24584 48790 24585 sw
rect 44768 24583 48790 24584
tri 48790 24583 48791 24584 sw
rect 44768 24582 48791 24583
tri 48791 24582 48792 24583 sw
rect 44768 24581 48792 24582
tri 48792 24581 48793 24582 sw
rect 44768 24580 48793 24581
tri 48793 24580 48794 24581 sw
rect 44768 24579 48794 24580
tri 48794 24579 48795 24580 sw
rect 44768 24578 48795 24579
tri 48795 24578 48796 24579 sw
rect 44768 24577 48796 24578
tri 48796 24577 48797 24578 sw
rect 44768 24576 48797 24577
tri 48797 24576 48798 24577 sw
rect 44768 24575 48798 24576
tri 48798 24575 48799 24576 sw
rect 44768 24574 48799 24575
tri 48799 24574 48800 24575 sw
rect 44768 24573 48800 24574
tri 48800 24573 48801 24574 sw
rect 44768 24572 48801 24573
tri 48801 24572 48802 24573 sw
rect 44768 24571 48802 24572
tri 48802 24571 48803 24572 sw
rect 44768 24570 48803 24571
tri 48803 24570 48804 24571 sw
rect 44768 24569 48804 24570
tri 48804 24569 48805 24570 sw
rect 44768 24568 48805 24569
tri 48805 24568 48806 24569 sw
rect 44768 24567 48806 24568
tri 48806 24567 48807 24568 sw
rect 44768 24566 48807 24567
tri 48807 24566 48808 24567 sw
rect 44768 24565 48808 24566
tri 48808 24565 48809 24566 sw
rect 44768 24564 48809 24565
tri 48809 24564 48810 24565 sw
rect 44768 24563 48810 24564
tri 48810 24563 48811 24564 sw
rect 44768 24562 48811 24563
tri 48811 24562 48812 24563 sw
rect 44768 24561 48812 24562
tri 48812 24561 48813 24562 sw
rect 44768 24560 48813 24561
tri 48813 24560 48814 24561 sw
rect 44768 24559 48814 24560
tri 48814 24559 48815 24560 sw
rect 44768 24558 48815 24559
tri 48815 24558 48816 24559 sw
rect 44768 24557 48816 24558
tri 48816 24557 48817 24558 sw
rect 44768 24556 48817 24557
tri 48817 24556 48818 24557 sw
rect 44768 24555 48818 24556
tri 48818 24555 48819 24556 sw
rect 44768 24554 48819 24555
tri 48819 24554 48820 24555 sw
rect 44768 24553 48820 24554
tri 48820 24553 48821 24554 sw
rect 44768 24552 48821 24553
tri 48821 24552 48822 24553 sw
rect 44768 24551 48822 24552
tri 48822 24551 48823 24552 sw
rect 44768 24550 48823 24551
tri 48823 24550 48824 24551 sw
rect 44768 24549 48824 24550
tri 48824 24549 48825 24550 sw
rect 44768 24548 48825 24549
tri 48825 24548 48826 24549 sw
rect 44768 24547 48826 24548
tri 48826 24547 48827 24548 sw
rect 44768 24546 48827 24547
tri 48827 24546 48828 24547 sw
rect 44768 24545 48828 24546
tri 48828 24545 48829 24546 sw
rect 44768 24544 48829 24545
tri 48829 24544 48830 24545 sw
rect 44768 24543 48830 24544
tri 48830 24543 48831 24544 sw
rect 44768 24542 48831 24543
tri 48831 24542 48832 24543 sw
rect 44768 24541 48832 24542
tri 48832 24541 48833 24542 sw
rect 44768 24540 48833 24541
tri 48833 24540 48834 24541 sw
rect 44768 24539 48834 24540
tri 48834 24539 48835 24540 sw
rect 44768 24538 48835 24539
tri 48835 24538 48836 24539 sw
rect 44768 24537 48836 24538
tri 48836 24537 48837 24538 sw
rect 44768 24536 48837 24537
tri 48837 24536 48838 24537 sw
rect 44768 24535 48838 24536
tri 48838 24535 48839 24536 sw
rect 44768 24534 48839 24535
tri 48839 24534 48840 24535 sw
rect 44768 24533 48840 24534
tri 48840 24533 48841 24534 sw
rect 44768 24532 48841 24533
tri 48841 24532 48842 24533 sw
rect 44768 24531 48842 24532
tri 48842 24531 48843 24532 sw
rect 44768 24530 48843 24531
tri 48843 24530 48844 24531 sw
rect 44768 24529 48844 24530
tri 48844 24529 48845 24530 sw
rect 44768 24528 48845 24529
tri 48845 24528 48846 24529 sw
rect 44768 24527 48846 24528
tri 48846 24527 48847 24528 sw
rect 44768 24526 48847 24527
tri 48847 24526 48848 24527 sw
rect 44768 24525 48848 24526
tri 48848 24525 48849 24526 sw
rect 44768 24524 48849 24525
tri 48849 24524 48850 24525 sw
rect 44768 24523 48850 24524
tri 48850 24523 48851 24524 sw
rect 44768 24522 48851 24523
tri 48851 24522 48852 24523 sw
rect 44768 24521 48852 24522
tri 48852 24521 48853 24522 sw
rect 44768 24520 48853 24521
tri 48853 24520 48854 24521 sw
rect 44768 24519 48854 24520
tri 48854 24519 48855 24520 sw
rect 44768 24518 48855 24519
tri 48855 24518 48856 24519 sw
rect 44768 24517 48856 24518
tri 48856 24517 48857 24518 sw
rect 44768 24516 48857 24517
tri 48857 24516 48858 24517 sw
rect 44768 24515 48858 24516
tri 48858 24515 48859 24516 sw
rect 44768 24514 48859 24515
tri 48859 24514 48860 24515 sw
rect 44768 24513 48860 24514
tri 48860 24513 48861 24514 sw
rect 44768 24512 48861 24513
tri 48861 24512 48862 24513 sw
rect 44768 24511 48862 24512
tri 48862 24511 48863 24512 sw
rect 44768 24510 48863 24511
tri 48863 24510 48864 24511 sw
rect 44768 24509 48864 24510
tri 48864 24509 48865 24510 sw
rect 44768 24508 48865 24509
tri 48865 24508 48866 24509 sw
rect 44768 24507 48866 24508
tri 48866 24507 48867 24508 sw
rect 44768 24506 48867 24507
tri 48867 24506 48868 24507 sw
rect 44768 24505 48868 24506
tri 48868 24505 48869 24506 sw
rect 44768 24504 48869 24505
tri 48869 24504 48870 24505 sw
rect 44768 24503 48870 24504
tri 48870 24503 48871 24504 sw
rect 44768 24502 48871 24503
tri 48871 24502 48872 24503 sw
rect 44768 24501 48872 24502
tri 48872 24501 48873 24502 sw
rect 44768 24500 48873 24501
tri 48873 24500 48874 24501 sw
rect 44768 24499 48874 24500
tri 48874 24499 48875 24500 sw
rect 44768 24498 48875 24499
tri 48875 24498 48876 24499 sw
rect 44768 24497 48876 24498
tri 48876 24497 48877 24498 sw
rect 44768 24496 48877 24497
tri 48877 24496 48878 24497 sw
rect 44768 24495 48878 24496
tri 48878 24495 48879 24496 sw
rect 44768 24494 48879 24495
tri 48879 24494 48880 24495 sw
rect 44768 24493 48880 24494
tri 48880 24493 48881 24494 sw
rect 44768 24492 48881 24493
tri 48881 24492 48882 24493 sw
rect 44768 24491 48882 24492
tri 48882 24491 48883 24492 sw
rect 44768 24490 48883 24491
tri 48883 24490 48884 24491 sw
rect 44768 24489 48884 24490
tri 48884 24489 48885 24490 sw
rect 44768 24488 48885 24489
tri 48885 24488 48886 24489 sw
rect 44768 24487 48886 24488
tri 48886 24487 48887 24488 sw
rect 44768 24486 48887 24487
tri 48887 24486 48888 24487 sw
rect 44768 24485 48888 24486
tri 48888 24485 48889 24486 sw
rect 44768 24484 48889 24485
tri 48889 24484 48890 24485 sw
rect 44768 24483 48890 24484
tri 48890 24483 48891 24484 sw
rect 44768 24482 48891 24483
tri 48891 24482 48892 24483 sw
rect 44768 24481 48892 24482
tri 48892 24481 48893 24482 sw
rect 44768 24480 48893 24481
tri 48893 24480 48894 24481 sw
rect 44768 24479 48894 24480
tri 48894 24479 48895 24480 sw
rect 44768 24478 48895 24479
tri 48895 24478 48896 24479 sw
rect 44768 24477 48896 24478
tri 48896 24477 48897 24478 sw
rect 44768 24476 48897 24477
tri 48897 24476 48898 24477 sw
rect 44768 24475 48898 24476
tri 48898 24475 48899 24476 sw
rect 44768 24474 48899 24475
tri 48899 24474 48900 24475 sw
rect 44768 24473 48900 24474
tri 48900 24473 48901 24474 sw
rect 44768 24472 48901 24473
tri 48901 24472 48902 24473 sw
rect 44768 24471 48902 24472
tri 48902 24471 48903 24472 sw
rect 44768 24470 48903 24471
tri 48903 24470 48904 24471 sw
rect 44768 24469 48904 24470
tri 48904 24469 48905 24470 sw
rect 44768 24468 48905 24469
tri 48905 24468 48906 24469 sw
rect 44768 24467 48906 24468
tri 48906 24467 48907 24468 sw
rect 44768 24466 48907 24467
tri 48907 24466 48908 24467 sw
rect 44768 24465 48908 24466
tri 48908 24465 48909 24466 sw
rect 44768 24464 48909 24465
tri 48909 24464 48910 24465 sw
rect 44768 24463 48910 24464
tri 48910 24463 48911 24464 sw
rect 44768 24462 48911 24463
tri 48911 24462 48912 24463 sw
rect 44768 24461 48912 24462
tri 48912 24461 48913 24462 sw
rect 44768 24460 48913 24461
tri 48913 24460 48914 24461 sw
rect 44768 24459 48914 24460
tri 48914 24459 48915 24460 sw
rect 44768 24458 48915 24459
tri 48915 24458 48916 24459 sw
rect 44768 24457 48916 24458
tri 48916 24457 48917 24458 sw
rect 44768 24456 48917 24457
tri 48917 24456 48918 24457 sw
rect 44768 24455 48918 24456
tri 48918 24455 48919 24456 sw
rect 44768 24454 48919 24455
tri 48919 24454 48920 24455 sw
rect 44768 24453 48920 24454
tri 48920 24453 48921 24454 sw
rect 44768 24452 48921 24453
tri 48921 24452 48922 24453 sw
rect 44768 24451 48922 24452
tri 48922 24451 48923 24452 sw
rect 44768 24450 48923 24451
tri 48923 24450 48924 24451 sw
rect 44768 24449 48924 24450
tri 48924 24449 48925 24450 sw
rect 44768 24448 48925 24449
tri 48925 24448 48926 24449 sw
rect 44768 24447 48926 24448
tri 48926 24447 48927 24448 sw
rect 44768 24446 48927 24447
tri 48927 24446 48928 24447 sw
rect 44768 24445 48928 24446
tri 48928 24445 48929 24446 sw
rect 44768 24444 48929 24445
tri 48929 24444 48930 24445 sw
rect 44768 24443 48930 24444
tri 48930 24443 48931 24444 sw
tri 48969 24443 49228 24702 ne
rect 49228 24443 70613 24702
rect 44768 24362 48931 24443
rect 40454 24150 44486 24362
rect 38624 23858 40162 24150
tri 40162 23858 40454 24150 sw
tri 40454 23989 40615 24150 ne
rect 40615 24080 44486 24150
tri 44486 24080 44768 24362 sw
tri 44768 24160 44970 24362 ne
rect 44970 24160 48931 24362
rect 40615 23989 44768 24080
rect 38624 23697 40454 23858
tri 40454 23697 40615 23858 sw
tri 40615 23697 40907 23989 ne
rect 40907 23878 44768 23989
tri 44768 23878 44970 24080 sw
tri 44970 23979 45151 24160 ne
rect 45151 24146 48931 24160
tri 48931 24146 49228 24443 sw
tri 49228 24146 49525 24443 ne
rect 49525 24146 70613 24443
rect 45151 23979 49228 24146
rect 40907 23697 44970 23878
tri 44970 23697 45151 23878 sw
tri 45151 23697 45433 23979 ne
rect 45433 23849 49228 23979
tri 49228 23849 49525 24146 sw
tri 49525 23994 49677 24146 ne
rect 49677 23994 70613 24146
rect 45433 23697 49525 23849
tri 49525 23697 49677 23849 sw
tri 49677 23697 49974 23994 ne
rect 49974 23706 70613 23994
rect 70669 23706 71000 24906
rect 49974 23697 71000 23706
rect 38624 23405 40615 23697
tri 40615 23405 40907 23697 sw
tri 40907 23695 40909 23697 ne
rect 40909 23695 45151 23697
rect 38624 23403 40907 23405
tri 40907 23403 40909 23405 sw
tri 40909 23403 41201 23695 ne
rect 41201 23415 45151 23695
tri 45151 23415 45433 23697 sw
tri 45433 23683 45447 23697 ne
rect 45447 23683 49677 23697
rect 41201 23403 45433 23415
rect 38624 23402 40909 23403
tri 40909 23402 40910 23403 sw
tri 41201 23402 41202 23403 ne
rect 41202 23402 45433 23403
rect 38624 23110 40910 23402
tri 40910 23110 41202 23402 sw
tri 41202 23110 41494 23402 ne
rect 41494 23401 45433 23402
tri 45433 23401 45447 23415 sw
tri 45447 23401 45729 23683 ne
rect 45729 23401 49677 23683
rect 41494 23119 45447 23401
tri 45447 23119 45729 23401 sw
tri 45729 23399 45731 23401 ne
rect 45731 23400 49677 23401
tri 49677 23400 49974 23697 sw
tri 49974 23600 50071 23697 ne
rect 50071 23600 71000 23697
rect 45731 23399 71000 23400
rect 41494 23117 45729 23119
tri 45729 23117 45731 23119 sw
tri 45731 23117 46013 23399 ne
rect 46013 23117 71000 23399
rect 41494 23116 45731 23117
tri 45731 23116 45732 23117 sw
tri 46013 23116 46014 23117 ne
rect 46014 23116 71000 23117
rect 41494 23110 45732 23116
rect 38624 22818 41202 23110
tri 41202 22818 41494 23110 sw
tri 41494 23109 41495 23110 ne
rect 41495 23109 45732 23110
rect 38624 22817 41494 22818
tri 41494 22817 41495 22818 sw
tri 41495 22817 41787 23109 ne
rect 41787 22834 45732 23109
tri 45732 22834 46014 23116 sw
tri 46014 22834 46296 23116 ne
rect 46296 22834 71000 23116
rect 41787 22817 46014 22834
rect 38624 22525 41495 22817
tri 41495 22525 41787 22817 sw
tri 41787 22780 41824 22817 ne
rect 41824 22780 46014 22817
rect 38624 22488 41787 22525
tri 41787 22488 41824 22525 sw
tri 41824 22523 42081 22780 ne
rect 42081 22552 46014 22780
tri 46014 22552 46296 22834 sw
tri 46296 22833 46297 22834 ne
rect 46297 22833 71000 22834
rect 42081 22551 46296 22552
tri 46296 22551 46297 22552 sw
tri 46297 22551 46579 22833 ne
rect 46579 22551 71000 22833
rect 42081 22523 46297 22551
rect 38624 22487 41824 22488
tri 41824 22487 41825 22488 sw
rect 38624 22486 41825 22487
tri 41825 22486 41826 22487 sw
rect 38624 22485 41826 22486
tri 41826 22485 41827 22486 sw
rect 38624 22484 41827 22485
tri 41827 22484 41828 22485 sw
rect 38624 22483 41828 22484
tri 41828 22483 41829 22484 sw
rect 38624 22482 41829 22483
tri 41829 22482 41830 22483 sw
rect 38624 22481 41830 22482
tri 41830 22481 41831 22482 sw
rect 38624 22480 41831 22481
tri 41831 22480 41832 22481 sw
rect 38624 22479 41832 22480
tri 41832 22479 41833 22480 sw
rect 38624 22478 41833 22479
tri 41833 22478 41834 22479 sw
rect 38624 22477 41834 22478
tri 41834 22477 41835 22478 sw
rect 38624 22476 41835 22477
tri 41835 22476 41836 22477 sw
rect 38624 22475 41836 22476
tri 41836 22475 41837 22476 sw
rect 38624 22474 41837 22475
tri 41837 22474 41838 22475 sw
rect 38624 22473 41838 22474
tri 41838 22473 41839 22474 sw
rect 38624 22472 41839 22473
tri 41839 22472 41840 22473 sw
rect 38624 22471 41840 22472
tri 41840 22471 41841 22472 sw
rect 38624 22470 41841 22471
tri 41841 22470 41842 22471 sw
rect 38624 22469 41842 22470
tri 41842 22469 41843 22470 sw
rect 38624 22468 41843 22469
tri 41843 22468 41844 22469 sw
rect 38624 22467 41844 22468
tri 41844 22467 41845 22468 sw
rect 38624 22466 41845 22467
tri 41845 22466 41846 22467 sw
rect 38624 22465 41846 22466
tri 41846 22465 41847 22466 sw
rect 38624 22464 41847 22465
tri 41847 22464 41848 22465 sw
rect 38624 22463 41848 22464
tri 41848 22463 41849 22464 sw
rect 38624 22462 41849 22463
tri 41849 22462 41850 22463 sw
rect 38624 22461 41850 22462
tri 41850 22461 41851 22462 sw
rect 38624 22460 41851 22461
tri 41851 22460 41852 22461 sw
rect 38624 22459 41852 22460
tri 41852 22459 41853 22460 sw
rect 38624 22458 41853 22459
tri 41853 22458 41854 22459 sw
rect 38624 22457 41854 22458
tri 41854 22457 41855 22458 sw
rect 38624 22456 41855 22457
tri 41855 22456 41856 22457 sw
rect 38624 22455 41856 22456
tri 41856 22455 41857 22456 sw
rect 38624 22454 41857 22455
tri 41857 22454 41858 22455 sw
rect 38624 22453 41858 22454
tri 41858 22453 41859 22454 sw
rect 38624 22452 41859 22453
tri 41859 22452 41860 22453 sw
rect 38624 22451 41860 22452
tri 41860 22451 41861 22452 sw
rect 38624 22450 41861 22451
tri 41861 22450 41862 22451 sw
rect 38624 22449 41862 22450
tri 41862 22449 41863 22450 sw
rect 38624 22448 41863 22449
tri 41863 22448 41864 22449 sw
rect 38624 22447 41864 22448
tri 41864 22447 41865 22448 sw
rect 38624 22446 41865 22447
tri 41865 22446 41866 22447 sw
rect 38624 22445 41866 22446
tri 41866 22445 41867 22446 sw
rect 38624 22444 41867 22445
tri 41867 22444 41868 22445 sw
rect 38624 22443 41868 22444
tri 41868 22443 41869 22444 sw
rect 38624 22442 41869 22443
tri 41869 22442 41870 22443 sw
rect 38624 22441 41870 22442
tri 41870 22441 41871 22442 sw
rect 38624 22440 41871 22441
tri 41871 22440 41872 22441 sw
rect 38624 22439 41872 22440
tri 41872 22439 41873 22440 sw
rect 38624 22438 41873 22439
tri 41873 22438 41874 22439 sw
rect 38624 22437 41874 22438
tri 41874 22437 41875 22438 sw
rect 38624 22436 41875 22437
tri 41875 22436 41876 22437 sw
rect 38624 22435 41876 22436
tri 41876 22435 41877 22436 sw
rect 38624 22434 41877 22435
tri 41877 22434 41878 22435 sw
rect 38624 22433 41878 22434
tri 41878 22433 41879 22434 sw
rect 38624 22432 41879 22433
tri 41879 22432 41880 22433 sw
rect 38624 22431 41880 22432
tri 41880 22431 41881 22432 sw
rect 38624 22430 41881 22431
tri 41881 22430 41882 22431 sw
rect 38624 22429 41882 22430
tri 41882 22429 41883 22430 sw
rect 38624 22428 41883 22429
tri 41883 22428 41884 22429 sw
rect 38624 22427 41884 22428
tri 41884 22427 41885 22428 sw
rect 38624 22426 41885 22427
tri 41885 22426 41886 22427 sw
rect 38624 22425 41886 22426
tri 41886 22425 41887 22426 sw
rect 38624 22424 41887 22425
tri 41887 22424 41888 22425 sw
rect 38624 22423 41888 22424
tri 41888 22423 41889 22424 sw
rect 38624 22422 41889 22423
tri 41889 22422 41890 22423 sw
rect 38624 22421 41890 22422
tri 41890 22421 41891 22422 sw
rect 38624 22420 41891 22421
tri 41891 22420 41892 22421 sw
rect 38624 22419 41892 22420
tri 41892 22419 41893 22420 sw
rect 38624 22418 41893 22419
tri 41893 22418 41894 22419 sw
rect 38624 22417 41894 22418
tri 41894 22417 41895 22418 sw
rect 38624 22416 41895 22417
tri 41895 22416 41896 22417 sw
rect 38624 22415 41896 22416
tri 41896 22415 41897 22416 sw
tri 42081 22415 42189 22523 ne
rect 42189 22415 46297 22523
rect 38624 22123 41897 22415
tri 41897 22123 42189 22415 sw
tri 42189 22123 42481 22415 ne
rect 42481 22269 46297 22415
tri 46297 22269 46579 22551 sw
tri 46579 22550 46580 22551 ne
rect 46580 22550 71000 22551
rect 42481 22268 46579 22269
tri 46579 22268 46580 22269 sw
tri 46580 22268 46862 22550 ne
rect 46862 22268 71000 22550
rect 42481 22123 46580 22268
rect 38624 21831 42189 22123
tri 42189 21831 42481 22123 sw
tri 42481 22122 42482 22123 ne
rect 42482 22122 46580 22123
rect 38624 21830 42481 21831
tri 42481 21830 42482 21831 sw
tri 42482 21830 42774 22122 ne
rect 42774 21986 46580 22122
tri 46580 21986 46862 22268 sw
tri 46862 22092 47038 22268 ne
rect 47038 22092 71000 22268
rect 42774 21830 46862 21986
rect 38624 21538 42482 21830
tri 42482 21538 42774 21830 sw
tri 42774 21829 42775 21830 ne
rect 42775 21829 46862 21830
rect 38624 21537 42774 21538
tri 42774 21537 42775 21538 sw
tri 42775 21537 43067 21829 ne
rect 43067 21810 46862 21829
tri 46862 21810 47038 21986 sw
tri 47038 21810 47320 22092 ne
rect 47320 21810 71000 22092
rect 43067 21537 47038 21810
rect 38624 21444 42775 21537
tri 38624 17293 42775 21444 ne
tri 42775 21245 43067 21537 sw
tri 43067 21444 43160 21537 ne
rect 43160 21528 47038 21537
tri 47038 21528 47320 21810 sw
tri 47320 21726 47404 21810 ne
rect 47404 21726 71000 21810
rect 43160 21444 47320 21528
tri 47320 21444 47404 21528 sw
tri 47404 21525 47605 21726 ne
rect 47605 21525 71000 21726
rect 42775 21152 43067 21245
tri 43067 21152 43160 21245 sw
tri 43160 21152 43452 21444 ne
rect 43452 21443 47404 21444
tri 47404 21443 47405 21444 sw
rect 43452 21442 47405 21443
tri 47405 21442 47406 21443 sw
rect 43452 21441 47406 21442
tri 47406 21441 47407 21442 sw
rect 43452 21440 47407 21441
tri 47407 21440 47408 21441 sw
rect 43452 21439 47408 21440
tri 47408 21439 47409 21440 sw
rect 43452 21438 47409 21439
tri 47409 21438 47410 21439 sw
rect 43452 21437 47410 21438
tri 47410 21437 47411 21438 sw
rect 43452 21436 47411 21437
tri 47411 21436 47412 21437 sw
rect 43452 21435 47412 21436
tri 47412 21435 47413 21436 sw
rect 43452 21434 47413 21435
tri 47413 21434 47414 21435 sw
rect 43452 21433 47414 21434
tri 47414 21433 47415 21434 sw
rect 43452 21432 47415 21433
tri 47415 21432 47416 21433 sw
rect 43452 21431 47416 21432
tri 47416 21431 47417 21432 sw
rect 43452 21430 47417 21431
tri 47417 21430 47418 21431 sw
rect 43452 21429 47418 21430
tri 47418 21429 47419 21430 sw
rect 43452 21428 47419 21429
tri 47419 21428 47420 21429 sw
rect 43452 21427 47420 21428
tri 47420 21427 47421 21428 sw
rect 43452 21426 47421 21427
tri 47421 21426 47422 21427 sw
rect 43452 21425 47422 21426
tri 47422 21425 47423 21426 sw
rect 43452 21424 47423 21425
tri 47423 21424 47424 21425 sw
rect 43452 21423 47424 21424
tri 47424 21423 47425 21424 sw
rect 43452 21422 47425 21423
tri 47425 21422 47426 21423 sw
rect 43452 21421 47426 21422
tri 47426 21421 47427 21422 sw
rect 43452 21420 47427 21421
tri 47427 21420 47428 21421 sw
rect 43452 21419 47428 21420
tri 47428 21419 47429 21420 sw
rect 43452 21418 47429 21419
tri 47429 21418 47430 21419 sw
rect 43452 21417 47430 21418
tri 47430 21417 47431 21418 sw
rect 43452 21416 47431 21417
tri 47431 21416 47432 21417 sw
rect 43452 21415 47432 21416
tri 47432 21415 47433 21416 sw
rect 43452 21414 47433 21415
tri 47433 21414 47434 21415 sw
rect 43452 21413 47434 21414
tri 47434 21413 47435 21414 sw
rect 43452 21412 47435 21413
tri 47435 21412 47436 21413 sw
rect 43452 21411 47436 21412
tri 47436 21411 47437 21412 sw
rect 43452 21410 47437 21411
tri 47437 21410 47438 21411 sw
rect 43452 21409 47438 21410
tri 47438 21409 47439 21410 sw
rect 43452 21408 47439 21409
tri 47439 21408 47440 21409 sw
rect 43452 21407 47440 21408
tri 47440 21407 47441 21408 sw
rect 43452 21406 47441 21407
tri 47441 21406 47442 21407 sw
rect 43452 21405 47442 21406
tri 47442 21405 47443 21406 sw
rect 43452 21404 47443 21405
tri 47443 21404 47444 21405 sw
rect 43452 21403 47444 21404
tri 47444 21403 47445 21404 sw
rect 43452 21402 47445 21403
tri 47445 21402 47446 21403 sw
rect 43452 21401 47446 21402
tri 47446 21401 47447 21402 sw
rect 43452 21400 47447 21401
tri 47447 21400 47448 21401 sw
rect 43452 21399 47448 21400
tri 47448 21399 47449 21400 sw
rect 43452 21398 47449 21399
tri 47449 21398 47450 21399 sw
rect 43452 21397 47450 21398
tri 47450 21397 47451 21398 sw
rect 43452 21396 47451 21397
tri 47451 21396 47452 21397 sw
rect 43452 21395 47452 21396
tri 47452 21395 47453 21396 sw
rect 43452 21394 47453 21395
tri 47453 21394 47454 21395 sw
rect 43452 21393 47454 21394
tri 47454 21393 47455 21394 sw
rect 43452 21392 47455 21393
tri 47455 21392 47456 21393 sw
rect 43452 21391 47456 21392
tri 47456 21391 47457 21392 sw
rect 43452 21390 47457 21391
tri 47457 21390 47458 21391 sw
rect 43452 21389 47458 21390
tri 47458 21389 47459 21390 sw
rect 43452 21388 47459 21389
tri 47459 21388 47460 21389 sw
rect 43452 21387 47460 21388
tri 47460 21387 47461 21388 sw
rect 43452 21386 47461 21387
tri 47461 21386 47462 21387 sw
rect 43452 21385 47462 21386
tri 47462 21385 47463 21386 sw
rect 43452 21384 47463 21385
tri 47463 21384 47464 21385 sw
rect 43452 21383 47464 21384
tri 47464 21383 47465 21384 sw
rect 43452 21382 47465 21383
tri 47465 21382 47466 21383 sw
rect 43452 21381 47466 21382
tri 47466 21381 47467 21382 sw
rect 43452 21380 47467 21381
tri 47467 21380 47468 21381 sw
rect 43452 21379 47468 21380
tri 47468 21379 47469 21380 sw
rect 43452 21378 47469 21379
tri 47469 21378 47470 21379 sw
rect 43452 21377 47470 21378
tri 47470 21377 47471 21378 sw
rect 43452 21376 47471 21377
tri 47471 21376 47472 21377 sw
rect 43452 21375 47472 21376
tri 47472 21375 47473 21376 sw
rect 43452 21374 47473 21375
tri 47473 21374 47474 21375 sw
rect 43452 21373 47474 21374
tri 47474 21373 47475 21374 sw
rect 43452 21372 47475 21373
tri 47475 21372 47476 21373 sw
rect 43452 21371 47476 21372
tri 47476 21371 47477 21372 sw
rect 43452 21370 47477 21371
tri 47477 21370 47478 21371 sw
rect 43452 21369 47478 21370
tri 47478 21369 47479 21370 sw
rect 43452 21368 47479 21369
tri 47479 21368 47480 21369 sw
rect 43452 21367 47480 21368
tri 47480 21367 47481 21368 sw
rect 43452 21366 47481 21367
tri 47481 21366 47482 21367 sw
rect 43452 21365 47482 21366
tri 47482 21365 47483 21366 sw
rect 43452 21364 47483 21365
tri 47483 21364 47484 21365 sw
rect 43452 21363 47484 21364
tri 47484 21363 47485 21364 sw
rect 43452 21362 47485 21363
tri 47485 21362 47486 21363 sw
rect 43452 21361 47486 21362
tri 47486 21361 47487 21362 sw
rect 43452 21360 47487 21361
tri 47487 21360 47488 21361 sw
rect 43452 21359 47488 21360
tri 47488 21359 47489 21360 sw
rect 43452 21358 47489 21359
tri 47489 21358 47490 21359 sw
rect 43452 21357 47490 21358
tri 47490 21357 47491 21358 sw
rect 43452 21356 47491 21357
tri 47491 21356 47492 21357 sw
rect 43452 21355 47492 21356
tri 47492 21355 47493 21356 sw
rect 43452 21354 47493 21355
tri 47493 21354 47494 21355 sw
rect 43452 21353 47494 21354
tri 47494 21353 47495 21354 sw
rect 43452 21352 47495 21353
tri 47495 21352 47496 21353 sw
rect 43452 21351 47496 21352
tri 47496 21351 47497 21352 sw
rect 43452 21350 47497 21351
tri 47497 21350 47498 21351 sw
rect 43452 21349 47498 21350
tri 47498 21349 47499 21350 sw
rect 43452 21348 47499 21349
tri 47499 21348 47500 21349 sw
rect 43452 21347 47500 21348
tri 47500 21347 47501 21348 sw
rect 43452 21346 47501 21347
tri 47501 21346 47502 21347 sw
rect 43452 21345 47502 21346
tri 47502 21345 47503 21346 sw
rect 43452 21344 47503 21345
tri 47503 21344 47504 21345 sw
rect 43452 21343 47504 21344
tri 47504 21343 47505 21344 sw
rect 43452 21342 47505 21343
tri 47505 21342 47506 21343 sw
rect 43452 21341 47506 21342
tri 47506 21341 47507 21342 sw
rect 43452 21340 47507 21341
tri 47507 21340 47508 21341 sw
rect 43452 21339 47508 21340
tri 47508 21339 47509 21340 sw
rect 43452 21338 47509 21339
tri 47509 21338 47510 21339 sw
rect 43452 21337 47510 21338
tri 47510 21337 47511 21338 sw
rect 43452 21336 47511 21337
tri 47511 21336 47512 21337 sw
rect 43452 21335 47512 21336
tri 47512 21335 47513 21336 sw
rect 43452 21334 47513 21335
tri 47513 21334 47514 21335 sw
rect 43452 21333 47514 21334
tri 47514 21333 47515 21334 sw
rect 43452 21332 47515 21333
tri 47515 21332 47516 21333 sw
rect 43452 21331 47516 21332
tri 47516 21331 47517 21332 sw
rect 43452 21330 47517 21331
tri 47517 21330 47518 21331 sw
rect 43452 21329 47518 21330
tri 47518 21329 47519 21330 sw
rect 43452 21328 47519 21329
tri 47519 21328 47520 21329 sw
rect 43452 21327 47520 21328
tri 47520 21327 47521 21328 sw
rect 43452 21326 47521 21327
tri 47521 21326 47522 21327 sw
rect 43452 21325 47522 21326
tri 47522 21325 47523 21326 sw
rect 43452 21324 47523 21325
tri 47523 21324 47524 21325 sw
rect 43452 21323 47524 21324
tri 47524 21323 47525 21324 sw
rect 43452 21322 47525 21323
tri 47525 21322 47526 21323 sw
rect 43452 21321 47526 21322
tri 47526 21321 47527 21322 sw
rect 43452 21320 47527 21321
tri 47527 21320 47528 21321 sw
rect 43452 21319 47528 21320
tri 47528 21319 47529 21320 sw
rect 43452 21318 47529 21319
tri 47529 21318 47530 21319 sw
rect 43452 21317 47530 21318
tri 47530 21317 47531 21318 sw
rect 43452 21316 47531 21317
tri 47531 21316 47532 21317 sw
rect 43452 21315 47532 21316
tri 47532 21315 47533 21316 sw
rect 43452 21314 47533 21315
tri 47533 21314 47534 21315 sw
rect 43452 21313 47534 21314
tri 47534 21313 47535 21314 sw
rect 43452 21312 47535 21313
tri 47535 21312 47536 21313 sw
rect 43452 21311 47536 21312
tri 47536 21311 47537 21312 sw
rect 43452 21310 47537 21311
tri 47537 21310 47538 21311 sw
rect 43452 21309 47538 21310
tri 47538 21309 47539 21310 sw
rect 43452 21308 47539 21309
tri 47539 21308 47540 21309 sw
rect 43452 21307 47540 21308
tri 47540 21307 47541 21308 sw
rect 43452 21306 47541 21307
tri 47541 21306 47542 21307 sw
rect 43452 21305 47542 21306
tri 47542 21305 47543 21306 sw
rect 43452 21304 47543 21305
tri 47543 21304 47544 21305 sw
rect 43452 21303 47544 21304
tri 47544 21303 47545 21304 sw
rect 43452 21302 47545 21303
tri 47545 21302 47546 21303 sw
rect 43452 21301 47546 21302
tri 47546 21301 47547 21302 sw
rect 43452 21300 47547 21301
tri 47547 21300 47548 21301 sw
rect 43452 21299 47548 21300
tri 47548 21299 47549 21300 sw
rect 43452 21298 47549 21299
tri 47549 21298 47550 21299 sw
rect 43452 21297 47550 21298
tri 47550 21297 47551 21298 sw
rect 43452 21296 47551 21297
tri 47551 21296 47552 21297 sw
rect 43452 21295 47552 21296
tri 47552 21295 47553 21296 sw
rect 43452 21294 47553 21295
tri 47553 21294 47554 21295 sw
rect 43452 21293 47554 21294
tri 47554 21293 47555 21294 sw
rect 43452 21292 47555 21293
tri 47555 21292 47556 21293 sw
rect 43452 21291 47556 21292
tri 47556 21291 47557 21292 sw
rect 43452 21290 47557 21291
tri 47557 21290 47558 21291 sw
rect 43452 21289 47558 21290
tri 47558 21289 47559 21290 sw
rect 43452 21288 47559 21289
tri 47559 21288 47560 21289 sw
rect 43452 21287 47560 21288
tri 47560 21287 47561 21288 sw
rect 43452 21286 47561 21287
tri 47561 21286 47562 21287 sw
rect 43452 21285 47562 21286
tri 47562 21285 47563 21286 sw
rect 43452 21284 47563 21285
tri 47563 21284 47564 21285 sw
rect 43452 21283 47564 21284
tri 47564 21283 47565 21284 sw
rect 43452 21282 47565 21283
tri 47565 21282 47566 21283 sw
rect 43452 21281 47566 21282
tri 47566 21281 47567 21282 sw
rect 43452 21280 47567 21281
tri 47567 21280 47568 21281 sw
rect 43452 21279 47568 21280
tri 47568 21279 47569 21280 sw
rect 43452 21278 47569 21279
tri 47569 21278 47570 21279 sw
rect 43452 21277 47570 21278
tri 47570 21277 47571 21278 sw
rect 43452 21276 47571 21277
tri 47571 21276 47572 21277 sw
rect 43452 21275 47572 21276
tri 47572 21275 47573 21276 sw
rect 43452 21274 47573 21275
tri 47573 21274 47574 21275 sw
rect 43452 21273 47574 21274
tri 47574 21273 47575 21274 sw
rect 43452 21272 47575 21273
tri 47575 21272 47576 21273 sw
rect 43452 21271 47576 21272
tri 47576 21271 47577 21272 sw
rect 43452 21270 47577 21271
tri 47577 21270 47578 21271 sw
rect 43452 21269 47578 21270
tri 47578 21269 47579 21270 sw
rect 43452 21268 47579 21269
tri 47579 21268 47580 21269 sw
rect 43452 21267 47580 21268
tri 47580 21267 47581 21268 sw
rect 43452 21266 47581 21267
tri 47581 21266 47582 21267 sw
rect 43452 21265 47582 21266
tri 47582 21265 47583 21266 sw
rect 43452 21264 47583 21265
tri 47583 21264 47584 21265 sw
rect 43452 21263 47584 21264
tri 47584 21263 47585 21264 sw
rect 43452 21262 47585 21263
tri 47585 21262 47586 21263 sw
rect 43452 21261 47586 21262
tri 47586 21261 47587 21262 sw
rect 43452 21260 47587 21261
tri 47587 21260 47588 21261 sw
rect 43452 21259 47588 21260
tri 47588 21259 47589 21260 sw
rect 43452 21258 47589 21259
tri 47589 21258 47590 21259 sw
rect 43452 21257 47590 21258
tri 47590 21257 47591 21258 sw
rect 43452 21256 47591 21257
tri 47591 21256 47592 21257 sw
rect 43452 21255 47592 21256
tri 47592 21255 47593 21256 sw
rect 43452 21254 47593 21255
tri 47593 21254 47594 21255 sw
rect 43452 21253 47594 21254
tri 47594 21253 47595 21254 sw
rect 43452 21252 47595 21253
tri 47595 21252 47596 21253 sw
rect 43452 21251 47596 21252
tri 47596 21251 47597 21252 sw
rect 43452 21250 47597 21251
tri 47597 21250 47598 21251 sw
rect 43452 21249 47598 21250
tri 47598 21249 47599 21250 sw
rect 43452 21248 47599 21249
tri 47599 21248 47600 21249 sw
rect 43452 21247 47600 21248
tri 47600 21247 47601 21248 sw
rect 43452 21246 47601 21247
tri 47601 21246 47602 21247 sw
rect 43452 21245 47602 21246
tri 47602 21245 47603 21246 sw
rect 43452 21244 47603 21245
tri 47603 21244 47604 21245 sw
rect 43452 21243 47604 21244
tri 47604 21243 47605 21244 sw
tri 47605 21243 47887 21525 ne
rect 47887 21243 71000 21525
rect 43452 21242 47605 21243
tri 47605 21242 47606 21243 sw
tri 47887 21242 47888 21243 ne
rect 47888 21242 71000 21243
rect 43452 21152 47606 21242
rect 42775 20860 43160 21152
tri 43160 20860 43452 21152 sw
tri 43452 20950 43654 21152 ne
rect 43654 20960 47606 21152
tri 47606 20960 47888 21242 sw
tri 47888 20960 48170 21242 ne
rect 48170 20960 71000 21242
rect 43654 20950 47888 20960
rect 42775 20658 43452 20860
tri 43452 20658 43654 20860 sw
tri 43654 20786 43818 20950 ne
rect 43818 20786 47888 20950
rect 42775 20494 43654 20658
tri 43654 20494 43818 20658 sw
tri 43818 20494 44110 20786 ne
rect 44110 20678 47888 20786
tri 47888 20678 48170 20960 sw
tri 48170 20683 48447 20960 ne
rect 48447 20683 71000 20960
rect 44110 20494 48170 20678
rect 42775 20202 43818 20494
tri 43818 20202 44110 20494 sw
tri 44110 20493 44111 20494 ne
rect 44111 20493 48170 20494
rect 42775 20201 44110 20202
tri 44110 20201 44111 20202 sw
tri 44111 20201 44403 20493 ne
rect 44403 20401 48170 20493
tri 48170 20401 48447 20678 sw
tri 48447 20482 48648 20683 ne
rect 48648 20482 71000 20683
rect 44403 20201 48447 20401
rect 42775 19909 44111 20201
tri 44111 19909 44403 20201 sw
tri 44403 20199 44405 20201 ne
rect 44405 20200 48447 20201
tri 48447 20200 48648 20401 sw
tri 48648 20400 48730 20482 ne
rect 48730 20400 71000 20482
rect 44405 20199 71000 20200
rect 42775 19907 44403 19909
tri 44403 19907 44405 19909 sw
tri 44405 19907 44697 20199 ne
rect 44697 19907 71000 20199
rect 42775 19906 44405 19907
tri 44405 19906 44406 19907 sw
tri 44697 19906 44698 19907 ne
rect 44698 19906 71000 19907
rect 42775 19614 44406 19906
tri 44406 19614 44698 19906 sw
tri 44698 19614 44990 19906 ne
rect 44990 19614 71000 19906
rect 42775 19322 44698 19614
tri 44698 19322 44990 19614 sw
tri 44990 19613 44991 19614 ne
rect 44991 19613 71000 19614
rect 42775 19321 44990 19322
tri 44990 19321 44991 19322 sw
tri 44991 19321 45283 19613 ne
rect 45283 19321 71000 19613
rect 42775 19029 44991 19321
tri 44991 19029 45283 19321 sw
tri 45283 19320 45284 19321 ne
rect 45284 19320 71000 19321
rect 42775 19028 45283 19029
tri 45283 19028 45284 19029 sw
tri 45284 19028 45576 19320 ne
rect 45576 19028 71000 19320
rect 42775 18736 45284 19028
tri 45284 18736 45576 19028 sw
tri 45576 19027 45577 19028 ne
rect 45577 19027 71000 19028
rect 42775 18735 45576 18736
tri 45576 18735 45577 18736 sw
tri 45577 18735 45869 19027 ne
rect 45869 18735 71000 19027
rect 42775 18443 45577 18735
tri 45577 18443 45869 18735 sw
tri 45869 18536 46068 18735 ne
rect 46068 18536 71000 18735
rect 42775 18244 45869 18443
tri 45869 18244 46068 18443 sw
tri 46068 18372 46232 18536 ne
rect 46232 18372 71000 18536
rect 42775 18080 46068 18244
tri 46068 18080 46232 18244 sw
tri 46232 18080 46524 18372 ne
rect 46524 18080 71000 18372
rect 42775 17788 46232 18080
tri 46232 17788 46524 18080 sw
tri 46524 18079 46525 18080 ne
rect 46525 18079 71000 18080
rect 42775 17787 46524 17788
tri 46524 17787 46525 17788 sw
tri 46525 17787 46817 18079 ne
rect 46817 17787 71000 18079
rect 42775 17495 46525 17787
tri 46525 17495 46817 17787 sw
tri 46817 17786 46818 17787 ne
rect 46818 17786 71000 17787
rect 42775 17494 46817 17495
tri 46817 17494 46818 17495 sw
tri 46818 17494 47110 17786 ne
rect 47110 17494 71000 17786
rect 42775 17293 46818 17494
tri 42775 14000 46068 17293 ne
rect 46068 17202 46818 17293
tri 46818 17202 47110 17494 sw
tri 47110 17292 47312 17494 ne
rect 47312 17292 71000 17494
rect 46068 17000 47110 17202
tri 47110 17000 47312 17202 sw
tri 47312 17200 47404 17292 ne
rect 47404 17200 71000 17292
rect 46068 14000 71000 17000
use M1_PSUB_CDNS_40661954729127  M1_PSUB_CDNS_40661954729127_0
timestamp 1698431365
transform -1 0 58007 0 -1 13194
box 0 0 1 1
use M1_PSUB_CDNS_40661954729128  M1_PSUB_CDNS_40661954729128_0
timestamp 1698431365
transform 0 -1 69871 1 0 70385
box 0 0 1 1
use M1_PSUB_CDNS_40661954729129  M1_PSUB_CDNS_40661954729129_0
timestamp 1698431365
transform 1 0 70235 0 1 69871
box 0 0 1 1
use M1_PSUB_CDNS_40661954729130  M1_PSUB_CDNS_40661954729130_0
timestamp 1698431365
transform 0 -1 70899 1 0 41649
box 0 0 1 1
use M1_PSUB_CDNS_40661954729130  M1_PSUB_CDNS_40661954729130_1
timestamp 1698431365
transform 1 0 41636 0 1 70900
box 0 0 1 1
use M1_PSUB_CDNS_40661954729131  M1_PSUB_CDNS_40661954729131_0
timestamp 1698431365
transform 0 -1 13194 1 0 58004
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_0
timestamp 1698431365
transform 1 0 42317 0 1 15761
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_1
timestamp 1698431365
transform 1 0 42185 0 1 15893
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_2
timestamp 1698431365
transform 1 0 42977 0 1 15101
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_3
timestamp 1698431365
transform 1 0 44873 0 1 13233
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_4
timestamp 1698431365
transform 1 0 44693 0 1 13385
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_5
timestamp 1698431365
transform 1 0 44561 0 1 13517
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_6
timestamp 1698431365
transform 1 0 44429 0 1 13649
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_7
timestamp 1698431365
transform 1 0 44297 0 1 13781
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_8
timestamp 1698431365
transform 1 0 44165 0 1 13913
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_9
timestamp 1698431365
transform 1 0 44033 0 1 14045
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_10
timestamp 1698431365
transform 1 0 43901 0 1 14177
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_11
timestamp 1698431365
transform 1 0 43769 0 1 14309
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_12
timestamp 1698431365
transform 1 0 43637 0 1 14441
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_13
timestamp 1698431365
transform 1 0 43505 0 1 14573
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_14
timestamp 1698431365
transform 1 0 43373 0 1 14705
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_15
timestamp 1698431365
transform 1 0 43241 0 1 14837
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_16
timestamp 1698431365
transform 1 0 43109 0 1 14969
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_17
timestamp 1698431365
transform 1 0 42845 0 1 15233
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_18
timestamp 1698431365
transform 1 0 42713 0 1 15365
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_19
timestamp 1698431365
transform 1 0 42581 0 1 15497
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_20
timestamp 1698431365
transform 1 0 42449 0 1 15629
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_21
timestamp 1698431365
transform 1 0 33605 0 1 24473
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_22
timestamp 1698431365
transform 1 0 39017 0 1 19061
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_23
timestamp 1698431365
transform 1 0 38885 0 1 19193
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_24
timestamp 1698431365
transform 1 0 38753 0 1 19325
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_25
timestamp 1698431365
transform 1 0 38621 0 1 19457
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_26
timestamp 1698431365
transform 1 0 38489 0 1 19589
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_27
timestamp 1698431365
transform 1 0 38357 0 1 19721
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_28
timestamp 1698431365
transform 1 0 33737 0 1 24341
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_29
timestamp 1698431365
transform 1 0 33869 0 1 24209
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_30
timestamp 1698431365
transform 1 0 34001 0 1 24077
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_31
timestamp 1698431365
transform 1 0 34133 0 1 23945
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_32
timestamp 1698431365
transform 1 0 34265 0 1 23813
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_33
timestamp 1698431365
transform 1 0 34397 0 1 23681
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_34
timestamp 1698431365
transform 1 0 34529 0 1 23549
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_35
timestamp 1698431365
transform 1 0 34661 0 1 23417
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_36
timestamp 1698431365
transform 1 0 34793 0 1 23285
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_37
timestamp 1698431365
transform 1 0 33209 0 1 24869
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_38
timestamp 1698431365
transform 1 0 39413 0 1 18665
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_39
timestamp 1698431365
transform 1 0 41261 0 1 16817
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_40
timestamp 1698431365
transform 1 0 36245 0 1 21833
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_41
timestamp 1698431365
transform 1 0 37301 0 1 20777
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_42
timestamp 1698431365
transform 1 0 37169 0 1 20909
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_43
timestamp 1698431365
transform 1 0 37037 0 1 21041
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_44
timestamp 1698431365
transform 1 0 36905 0 1 21173
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_45
timestamp 1698431365
transform 1 0 36773 0 1 21305
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_46
timestamp 1698431365
transform 1 0 36641 0 1 21437
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_47
timestamp 1698431365
transform 1 0 36509 0 1 21569
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_48
timestamp 1698431365
transform 1 0 36377 0 1 21701
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_49
timestamp 1698431365
transform 1 0 32945 0 1 25133
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_50
timestamp 1698431365
transform 1 0 32813 0 1 25265
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_51
timestamp 1698431365
transform 1 0 32681 0 1 25397
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_52
timestamp 1698431365
transform 1 0 32549 0 1 25529
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_53
timestamp 1698431365
transform 1 0 32417 0 1 25661
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_54
timestamp 1698431365
transform 1 0 32285 0 1 25793
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_55
timestamp 1698431365
transform 1 0 32153 0 1 25925
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_56
timestamp 1698431365
transform 1 0 32021 0 1 26057
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_57
timestamp 1698431365
transform 1 0 31889 0 1 26189
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_58
timestamp 1698431365
transform 1 0 31757 0 1 26321
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_59
timestamp 1698431365
transform 1 0 31625 0 1 26453
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_60
timestamp 1698431365
transform 1 0 31493 0 1 26585
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_61
timestamp 1698431365
transform 1 0 31361 0 1 26717
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_62
timestamp 1698431365
transform 1 0 31229 0 1 26849
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_63
timestamp 1698431365
transform 1 0 33077 0 1 25001
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_64
timestamp 1698431365
transform 1 0 30965 0 1 27113
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_65
timestamp 1698431365
transform 1 0 30833 0 1 27245
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_66
timestamp 1698431365
transform 1 0 30701 0 1 27377
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_67
timestamp 1698431365
transform 1 0 31097 0 1 26981
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_68
timestamp 1698431365
transform 1 0 36113 0 1 21965
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_69
timestamp 1698431365
transform 1 0 35981 0 1 22097
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_70
timestamp 1698431365
transform 1 0 35849 0 1 22229
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_71
timestamp 1698431365
transform 1 0 35717 0 1 22361
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_72
timestamp 1698431365
transform 1 0 35585 0 1 22493
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_73
timestamp 1698431365
transform 1 0 35453 0 1 22625
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_74
timestamp 1698431365
transform 1 0 35321 0 1 22757
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_75
timestamp 1698431365
transform 1 0 35189 0 1 22889
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_76
timestamp 1698431365
transform 1 0 34925 0 1 23153
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_77
timestamp 1698431365
transform 1 0 41921 0 1 16157
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_78
timestamp 1698431365
transform 1 0 41789 0 1 16289
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_79
timestamp 1698431365
transform 1 0 41657 0 1 16421
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_80
timestamp 1698431365
transform 1 0 41525 0 1 16553
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_81
timestamp 1698431365
transform 1 0 41393 0 1 16685
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_82
timestamp 1698431365
transform 1 0 39281 0 1 18797
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_83
timestamp 1698431365
transform 1 0 41129 0 1 16949
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_84
timestamp 1698431365
transform 1 0 40997 0 1 17081
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_85
timestamp 1698431365
transform 1 0 40865 0 1 17213
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_86
timestamp 1698431365
transform 1 0 40733 0 1 17345
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_87
timestamp 1698431365
transform 1 0 40601 0 1 17477
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_88
timestamp 1698431365
transform 1 0 40469 0 1 17609
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_89
timestamp 1698431365
transform 1 0 40337 0 1 17741
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_90
timestamp 1698431365
transform 1 0 40205 0 1 17873
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_91
timestamp 1698431365
transform 1 0 40073 0 1 18005
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_92
timestamp 1698431365
transform 1 0 39941 0 1 18137
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_93
timestamp 1698431365
transform 1 0 39809 0 1 18269
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_94
timestamp 1698431365
transform 1 0 39677 0 1 18401
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_95
timestamp 1698431365
transform 1 0 38225 0 1 19853
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_96
timestamp 1698431365
transform 1 0 38093 0 1 19985
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_97
timestamp 1698431365
transform 1 0 37961 0 1 20117
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_98
timestamp 1698431365
transform 1 0 37829 0 1 20249
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_99
timestamp 1698431365
transform 1 0 37697 0 1 20381
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_100
timestamp 1698431365
transform 1 0 37565 0 1 20513
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_101
timestamp 1698431365
transform 1 0 37433 0 1 20645
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_102
timestamp 1698431365
transform 1 0 39545 0 1 18533
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_103
timestamp 1698431365
transform 1 0 35057 0 1 23021
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_104
timestamp 1698431365
transform 1 0 39149 0 1 18929
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_105
timestamp 1698431365
transform 1 0 33341 0 1 24737
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_106
timestamp 1698431365
transform 1 0 33473 0 1 24605
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_107
timestamp 1698431365
transform 1 0 18689 0 1 39389
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_108
timestamp 1698431365
transform 1 0 23969 0 1 34109
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_109
timestamp 1698431365
transform 1 0 23045 0 1 35033
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_110
timestamp 1698431365
transform 1 0 23309 0 1 34769
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_111
timestamp 1698431365
transform 1 0 23441 0 1 34637
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_112
timestamp 1698431365
transform 1 0 23573 0 1 34505
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_113
timestamp 1698431365
transform 1 0 23705 0 1 34373
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_114
timestamp 1698431365
transform 1 0 23837 0 1 34241
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_115
timestamp 1698431365
transform 1 0 24101 0 1 33977
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_116
timestamp 1698431365
transform 1 0 24233 0 1 33845
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_117
timestamp 1698431365
transform 1 0 24365 0 1 33713
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_118
timestamp 1698431365
transform 1 0 24497 0 1 33581
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_119
timestamp 1698431365
transform 1 0 24629 0 1 33449
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_120
timestamp 1698431365
transform 1 0 24761 0 1 33317
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_121
timestamp 1698431365
transform 1 0 25025 0 1 33053
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_122
timestamp 1698431365
transform 1 0 23177 0 1 34901
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_123
timestamp 1698431365
transform 1 0 22913 0 1 35165
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_124
timestamp 1698431365
transform 1 0 22781 0 1 35297
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_125
timestamp 1698431365
transform 1 0 22649 0 1 35429
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_126
timestamp 1698431365
transform 1 0 22517 0 1 35561
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_127
timestamp 1698431365
transform 1 0 22385 0 1 35693
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_128
timestamp 1698431365
transform 1 0 22253 0 1 35825
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_129
timestamp 1698431365
transform 1 0 22121 0 1 35957
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_130
timestamp 1698431365
transform 1 0 21989 0 1 36089
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_131
timestamp 1698431365
transform 1 0 21857 0 1 36221
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_132
timestamp 1698431365
transform 1 0 21725 0 1 36353
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_133
timestamp 1698431365
transform 1 0 21593 0 1 36485
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_134
timestamp 1698431365
transform 1 0 21461 0 1 36617
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_135
timestamp 1698431365
transform 1 0 21329 0 1 36749
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_136
timestamp 1698431365
transform 1 0 21065 0 1 37013
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_137
timestamp 1698431365
transform 1 0 24893 0 1 33185
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_138
timestamp 1698431365
transform 1 0 18557 0 1 39521
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_139
timestamp 1698431365
transform 1 0 18425 0 1 39653
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_140
timestamp 1698431365
transform 1 0 18293 0 1 39785
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_141
timestamp 1698431365
transform 1 0 18161 0 1 39917
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_142
timestamp 1698431365
transform 1 0 16973 0 1 41105
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_143
timestamp 1698431365
transform 1 0 18029 0 1 40049
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_144
timestamp 1698431365
transform 1 0 17897 0 1 40181
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_145
timestamp 1698431365
transform 1 0 17765 0 1 40313
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_146
timestamp 1698431365
transform 1 0 17633 0 1 40445
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_147
timestamp 1698431365
transform 1 0 17501 0 1 40577
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_148
timestamp 1698431365
transform 1 0 17369 0 1 40709
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_149
timestamp 1698431365
transform 1 0 27401 0 1 30677
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_150
timestamp 1698431365
transform 1 0 27269 0 1 30809
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_151
timestamp 1698431365
transform 1 0 27137 0 1 30941
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_152
timestamp 1698431365
transform 1 0 21197 0 1 36881
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_153
timestamp 1698431365
transform 1 0 26873 0 1 31205
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_154
timestamp 1698431365
transform 1 0 26741 0 1 31337
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_155
timestamp 1698431365
transform 1 0 26609 0 1 31469
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_156
timestamp 1698431365
transform 1 0 26477 0 1 31601
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_157
timestamp 1698431365
transform 1 0 26345 0 1 31733
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_158
timestamp 1698431365
transform 1 0 26213 0 1 31865
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_159
timestamp 1698431365
transform 1 0 26081 0 1 31997
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_160
timestamp 1698431365
transform 1 0 25949 0 1 32129
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_161
timestamp 1698431365
transform 1 0 25817 0 1 32261
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_162
timestamp 1698431365
transform 1 0 25685 0 1 32393
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_163
timestamp 1698431365
transform 1 0 25553 0 1 32525
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_164
timestamp 1698431365
transform 1 0 25421 0 1 32657
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_165
timestamp 1698431365
transform 1 0 25289 0 1 32789
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_166
timestamp 1698431365
transform 1 0 25157 0 1 32921
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_167
timestamp 1698431365
transform 1 0 27005 0 1 31073
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_168
timestamp 1698431365
transform 1 0 17105 0 1 40973
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_169
timestamp 1698431365
transform 1 0 16841 0 1 41237
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_170
timestamp 1698431365
transform 1 0 16709 0 1 41369
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_171
timestamp 1698431365
transform 1 0 16577 0 1 41501
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_172
timestamp 1698431365
transform 1 0 16445 0 1 41633
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_173
timestamp 1698431365
transform 1 0 16313 0 1 41765
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_174
timestamp 1698431365
transform 1 0 16181 0 1 41897
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_175
timestamp 1698431365
transform 1 0 19085 0 1 38993
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_176
timestamp 1698431365
transform 1 0 20933 0 1 37145
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_177
timestamp 1698431365
transform 1 0 20801 0 1 37277
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_178
timestamp 1698431365
transform 1 0 20669 0 1 37409
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_179
timestamp 1698431365
transform 1 0 20537 0 1 37541
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_180
timestamp 1698431365
transform 1 0 20405 0 1 37673
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_181
timestamp 1698431365
transform 1 0 20273 0 1 37805
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_182
timestamp 1698431365
transform 1 0 20141 0 1 37937
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_183
timestamp 1698431365
transform 1 0 20009 0 1 38069
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_184
timestamp 1698431365
transform 1 0 19877 0 1 38201
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_185
timestamp 1698431365
transform 1 0 19745 0 1 38333
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_186
timestamp 1698431365
transform 1 0 19613 0 1 38465
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_187
timestamp 1698431365
transform 1 0 19481 0 1 38597
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_188
timestamp 1698431365
transform 1 0 19349 0 1 38729
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_189
timestamp 1698431365
transform 1 0 19217 0 1 38861
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_190
timestamp 1698431365
transform 1 0 17237 0 1 40841
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_191
timestamp 1698431365
transform 1 0 18953 0 1 39125
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_192
timestamp 1698431365
transform 1 0 18821 0 1 39257
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_193
timestamp 1698431365
transform 1 0 29117 0 1 28961
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_194
timestamp 1698431365
transform 1 0 28985 0 1 29093
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_195
timestamp 1698431365
transform 1 0 28721 0 1 29357
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_196
timestamp 1698431365
transform 1 0 28589 0 1 29489
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_197
timestamp 1698431365
transform 1 0 28457 0 1 29621
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_198
timestamp 1698431365
transform 1 0 28325 0 1 29753
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_199
timestamp 1698431365
transform 1 0 28193 0 1 29885
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_200
timestamp 1698431365
transform 1 0 28061 0 1 30017
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_201
timestamp 1698431365
transform 1 0 27929 0 1 30149
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_202
timestamp 1698431365
transform 1 0 27797 0 1 30281
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_203
timestamp 1698431365
transform 1 0 27665 0 1 30413
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_204
timestamp 1698431365
transform 1 0 29249 0 1 28829
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_205
timestamp 1698431365
transform 1 0 28853 0 1 29225
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_206
timestamp 1698431365
transform 1 0 29513 0 1 28565
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_207
timestamp 1698431365
transform 1 0 30437 0 1 27641
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_208
timestamp 1698431365
transform 1 0 30305 0 1 27773
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_209
timestamp 1698431365
transform 1 0 30173 0 1 27905
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_210
timestamp 1698431365
transform 1 0 30041 0 1 28037
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_211
timestamp 1698431365
transform 1 0 29909 0 1 28169
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_212
timestamp 1698431365
transform 1 0 29777 0 1 28301
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_213
timestamp 1698431365
transform 1 0 29645 0 1 28433
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_214
timestamp 1698431365
transform 1 0 29381 0 1 28697
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_215
timestamp 1698431365
transform 1 0 27533 0 1 30545
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_216
timestamp 1698431365
transform 1 0 30569 0 1 27509
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_217
timestamp 1698431365
transform 1 0 13937 0 1 44141
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_218
timestamp 1698431365
transform 1 0 13805 0 1 44273
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_219
timestamp 1698431365
transform 1 0 13673 0 1 44405
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_220
timestamp 1698431365
transform 1 0 13541 0 1 44537
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_221
timestamp 1698431365
transform 1 0 13409 0 1 44669
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_222
timestamp 1698431365
transform 1 0 13277 0 1 44801
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_223
timestamp 1698431365
transform 1 0 15125 0 1 42953
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_224
timestamp 1698431365
transform 1 0 15917 0 1 42161
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_225
timestamp 1698431365
transform 1 0 15785 0 1 42293
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_226
timestamp 1698431365
transform 1 0 15653 0 1 42425
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_227
timestamp 1698431365
transform 1 0 15521 0 1 42557
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_228
timestamp 1698431365
transform 1 0 15389 0 1 42689
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_229
timestamp 1698431365
transform 1 0 15257 0 1 42821
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_230
timestamp 1698431365
transform 1 0 14993 0 1 43085
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_231
timestamp 1698431365
transform 1 0 14861 0 1 43217
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_232
timestamp 1698431365
transform 1 0 14729 0 1 43349
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_233
timestamp 1698431365
transform 1 0 14597 0 1 43481
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_234
timestamp 1698431365
transform 1 0 14465 0 1 43613
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_235
timestamp 1698431365
transform 1 0 14333 0 1 43745
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_236
timestamp 1698431365
transform 1 0 14201 0 1 43877
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_237
timestamp 1698431365
transform 1 0 14069 0 1 44009
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_238
timestamp 1698431365
transform 1 0 16049 0 1 42029
box 0 0 1 1
use M1_PSUB_CDNS_40661954729132  M1_PSUB_CDNS_40661954729132_239
timestamp 1698431365
transform 1 0 42053 0 1 16025
box 0 0 1 1
use M3_M2_CDNS_40661954729133  M3_M2_CDNS_40661954729133_0
timestamp 1698431365
transform 1 0 70641 0 1 24306
box 0 0 1 1
use M3_M2_CDNS_40661954729133  M3_M2_CDNS_40661954729133_1
timestamp 1698431365
transform 1 0 70641 0 1 67516
box 0 0 1 1
use M3_M2_CDNS_40661954729133  M3_M2_CDNS_40661954729133_2
timestamp 1698431365
transform 1 0 70641 0 1 59520
box 0 0 1 1
use M3_M2_CDNS_40661954729133  M3_M2_CDNS_40661954729133_3
timestamp 1698431365
transform 1 0 70641 0 1 54702
box 0 0 1 1
use M3_M2_CDNS_40661954729133  M3_M2_CDNS_40661954729133_4
timestamp 1698431365
transform 1 0 70641 0 1 53122
box 0 0 1 1
use M3_M2_CDNS_40661954729133  M3_M2_CDNS_40661954729133_5
timestamp 1698431365
transform 1 0 70641 0 1 56310
box 0 0 1 1
use M3_M2_CDNS_40661954729133  M3_M2_CDNS_40661954729133_6
timestamp 1698431365
transform 1 0 70641 0 1 41897
box 0 0 1 1
use M3_M2_CDNS_40661954729134  M3_M2_CDNS_40661954729134_0
timestamp 1698431365
transform 1 0 70641 0 1 28320
box 0 0 1 1
use M3_M2_CDNS_40661954729134  M3_M2_CDNS_40661954729134_1
timestamp 1698431365
transform 1 0 70641 0 1 31488
box 0 0 1 1
use M3_M2_CDNS_40661954729134  M3_M2_CDNS_40661954729134_2
timestamp 1698431365
transform 1 0 70641 0 1 34700
box 0 0 1 1
use M3_M2_CDNS_40661954729134  M3_M2_CDNS_40661954729134_3
timestamp 1698431365
transform 1 0 70641 0 1 37900
box 0 0 1 1
use M3_M2_CDNS_40661954729134  M3_M2_CDNS_40661954729134_4
timestamp 1698431365
transform 1 0 70641 0 1 44307
box 0 0 1 1
<< labels >>
rlabel metal3 s 70454 64211 70454 64211 4 VSS
port 1 nsew
rlabel metal3 s 70454 62776 70454 62776 4 VDD
port 2 nsew
rlabel metal3 s 70454 61011 70454 61011 4 DVSS
port 3 nsew
rlabel metal3 s 70454 65976 70454 65976 4 DVSS
port 3 nsew
rlabel metal3 s 70454 69002 70454 69002 4 DVSS
port 3 nsew
rlabel metal3 s 70454 67411 70454 67411 4 DVDD
port 4 nsew
rlabel metal3 s 70454 59576 70454 59576 4 DVDD
port 4 nsew
rlabel metal3 s 70454 57811 70454 57811 4 DVSS
port 3 nsew
rlabel metal3 s 70454 56376 70454 56376 4 DVDD
port 4 nsew
rlabel metal3 s 70454 54611 70454 54611 4 DVDD
port 4 nsew
rlabel metal3 s 70454 53176 70454 53176 4 DVDD
port 4 nsew
rlabel metal3 s 70559 51411 70559 51411 4 VDD
port 2 nsew
rlabel metal3 s 70559 49976 70559 49976 4 VSS
port 1 nsew
rlabel metal3 s 70454 47548 70454 47548 4 DVSS
port 3 nsew
rlabel metal3 s 70454 44321 70454 44321 4 DVDD
port 4 nsew
rlabel metal3 s 70454 40295 70454 40295 4 DVSS
port 3 nsew
rlabel metal3 s 70454 41930 70454 41930 4 DVDD
port 4 nsew
rlabel metal3 s 70454 37912 70454 37912 4 DVDD
port 4 nsew
rlabel metal3 s 70454 34676 70454 34676 4 DVDD
port 4 nsew
rlabel metal3 s 70454 31562 70454 31562 4 DVDD
port 4 nsew
rlabel metal3 s 70454 28347 70454 28347 4 DVDD
port 4 nsew
rlabel metal3 s 70454 26053 70454 26053 4 DVSS
port 3 nsew
rlabel metal3 s 70454 24237 70454 24237 4 DVDD
port 4 nsew
rlabel metal3 s 70454 21860 70454 21860 4 DVSS
port 3 nsew
rlabel metal3 s 70385 18874 70385 18874 4 DVSS
port 3 nsew
rlabel metal3 s 70432 15703 70432 15703 4 DVSS
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 71000 71000
string GDS_END 11911992
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 11893050
string path 1687.500 1775.000 1687.500 1710.075 1710.075 1687.500 1775.000 1687.500 
<< end >>
