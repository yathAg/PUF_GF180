magic
tech gf180mcuD
magscale 1 10
timestamp 1698431365
<< deepnwell >>
rect -680 -680 788 3880
<< pbase >>
rect -180 -180 288 3380
<< ndiff >>
rect 0 3127 108 3200
rect 0 73 31 3127
rect 77 73 108 3127
rect 0 0 108 73
<< ndiffc >>
rect 31 73 77 3127
<< psubdiff >>
rect -1264 4445 1372 4464
rect -1264 4399 -1097 4445
rect 1205 4399 1372 4445
rect -1264 4380 1372 4399
rect -1264 4302 -1180 4380
rect -1264 -1102 -1245 4302
rect -1199 -1102 -1180 4302
rect 1288 4302 1372 4380
rect -148 3329 256 3348
rect -148 3283 -109 3329
rect 219 3283 256 3329
rect -148 3264 256 3283
rect -148 3220 -64 3264
rect -148 -22 -129 3220
rect -83 -22 -64 3220
rect 172 3220 256 3264
rect -148 -64 -64 -22
rect 172 -22 191 3220
rect 237 -22 256 3220
rect 172 -64 256 -22
rect -148 -148 256 -64
rect -1264 -1180 -1180 -1102
rect 1288 -1102 1307 4302
rect 1353 -1102 1372 4302
rect 1288 -1180 1372 -1102
rect -1264 -1199 1372 -1180
rect -1264 -1245 -1097 -1199
rect -769 -1245 877 -1199
rect 1205 -1245 1372 -1199
rect -1264 -1264 1372 -1245
<< nsubdiff >>
rect -296 3477 404 3496
rect -296 3431 -251 3477
rect 359 3431 404 3477
rect -296 3412 404 3431
rect -296 3361 -212 3412
rect -296 -163 -277 3361
rect -231 -163 -212 3361
rect 320 3361 404 3412
rect -296 -212 -212 -163
rect 320 -163 339 3361
rect 385 -163 404 3361
rect 320 -212 404 -163
rect -296 -296 404 -212
<< psubdiffcont >>
rect -1097 4399 1205 4445
rect -1245 -1102 -1199 4302
rect -109 3283 219 3329
rect -129 -22 -83 3220
rect 191 -22 237 3220
rect 1307 -1102 1353 4302
rect -1097 -1245 -769 -1199
rect 877 -1245 1205 -1199
<< nsubdiffcont >>
rect -251 3431 359 3477
rect -277 -163 -231 3361
rect 339 -163 385 3361
<< metal1 >>
rect -1264 4445 1372 4464
rect -1264 4399 -1097 4445
rect 1205 4399 1372 4445
rect -1264 4380 1372 4399
rect -1264 4302 -1180 4380
rect -1264 -1102 -1245 4302
rect -1199 -1102 -1180 4302
rect 1288 4302 1372 4380
rect -296 3477 404 3496
rect -296 3431 -251 3477
rect 359 3431 404 3477
rect -296 3412 404 3431
rect -296 3361 -212 3412
rect -296 -163 -277 3361
rect -231 -163 -212 3361
rect 320 3361 404 3412
rect -148 3329 256 3348
rect -148 3283 -109 3329
rect 219 3283 256 3329
rect -148 3264 256 3283
rect -148 3220 -64 3264
rect -148 -22 -129 3220
rect -83 -22 -64 3220
rect 172 3220 256 3264
rect 0 3127 108 3200
rect 0 73 31 3127
rect 77 73 108 3127
rect 0 0 108 73
rect -148 -148 -64 -22
rect 172 -22 191 3220
rect 237 -22 256 3220
rect 172 -148 256 -22
rect -296 -296 -212 -163
rect 320 -163 339 3361
rect 385 -163 404 3361
rect 320 -296 404 -163
rect -1264 -1180 -1180 -1102
rect 1288 -1102 1307 4302
rect 1353 -1102 1372 4302
rect 1288 -1180 1372 -1102
rect -1264 -1199 -680 -1180
rect -1264 -1245 -1097 -1199
rect -769 -1245 -680 -1199
rect -1264 -1264 -680 -1245
rect 788 -1199 1372 -1180
rect 788 -1245 877 -1199
rect 1205 -1245 1372 -1199
rect 788 -1264 1372 -1245
<< labels >>
flabel ndiffc 50 1832 50 1832 0 FreeSans 400 0 0 0 E
flabel metal1 214 -102 214 -102 0 FreeSans 400 0 0 0 B
flabel psubdiffcont 214 3301 214 3301 0 FreeSans 400 0 0 0 B
flabel metal1 -104 -99 -104 -99 0 FreeSans 400 0 0 0 B
flabel metal1 361 -248 361 -248 0 FreeSans 400 0 0 0 C
flabel metal1 362 3453 362 3453 0 FreeSans 400 0 0 0 C
flabel metal1 -248 -248 -248 -248 0 FreeSans 400 0 0 0 C
flabel metal1 -1223 -1221 -1223 -1221 0 FreeSans 400 0 0 0 S
flabel metal1 -1223 -1221 -1223 -1221 0 FreeSans 400 0 0 0 S
flabel metal1 1328 -1221 1328 -1221 0 FreeSans 400 0 0 0 S
flabel metal1 1328 -1221 1328 -1221 0 FreeSans 400 0 0 0 S
flabel metal1 1330 4422 1330 4422 0 FreeSans 400 0 0 0 S
<< properties >>
string GDS_END 25004
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_pr/gds/npn_00p54x16p00.gds
string GDS_START 112
string gencell npn_00p54x16p00
<< end >>
