magic
tech gf180mcuA
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 453 534 1094
<< pwell >>
rect -86 -86 534 453
<< metal1 >>
rect 0 918 448 1098
rect 50 589 96 918
rect 254 578 306 740
rect 50 90 96 271
rect 0 -90 448 90
<< obsm1 >>
rect 175 366 320 412
rect 274 263 320 366
<< labels >>
rlabel metal1 s 254 578 306 740 6 Z
port 1 nsew default output
rlabel metal1 s 50 589 96 918 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 0 918 448 1098 6 VDD
port 2 nsew power bidirectional abutment
rlabel nwell s -86 453 534 1094 6 VNW
port 3 nsew power bidirectional
rlabel pwell s -86 -86 534 453 6 VPW
port 4 nsew ground bidirectional
rlabel metal1 s 0 -90 448 90 8 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 50 90 96 271 6 VSS
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 448 1008
string LEFclass core TIEHIGH
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 443306
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 441202
<< end >>
