magic
tech gf180mcuA
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 407 3894 870
rect -86 352 575 407
rect 943 352 3894 407
<< pwell >>
rect 575 352 943 407
rect -86 -86 3894 352
<< mvnmos >>
rect 124 68 244 232
rect 348 68 468 232
rect 572 68 692 232
rect 1064 68 1184 232
rect 1288 68 1408 232
rect 1512 68 1632 232
rect 1736 68 1856 232
rect 1960 68 2080 232
rect 2184 68 2304 232
rect 2408 68 2528 232
rect 2632 68 2752 232
rect 2856 68 2976 232
rect 3080 68 3200 232
rect 3304 68 3424 232
rect 3528 68 3648 232
<< mvpmos >>
rect 172 527 272 716
rect 376 527 476 716
rect 660 527 760 716
rect 1144 481 1244 716
rect 1348 481 1448 716
rect 1552 481 1652 716
rect 1756 481 1856 716
rect 1960 481 2060 716
rect 2164 481 2264 716
rect 2368 481 2468 716
rect 2572 481 2672 716
rect 2776 481 2876 716
rect 2980 481 3080 716
rect 3184 481 3284 716
rect 3388 481 3488 716
<< mvndiff >>
rect 752 274 824 287
rect 752 232 765 274
rect 36 219 124 232
rect 36 173 49 219
rect 95 173 124 219
rect 36 68 124 173
rect 244 128 348 232
rect 244 82 273 128
rect 319 82 348 128
rect 244 68 348 82
rect 468 152 572 232
rect 468 106 497 152
rect 543 106 572 152
rect 468 68 572 106
rect 692 228 765 232
rect 811 228 824 274
rect 692 68 824 228
rect 932 95 1064 232
rect 932 49 945 95
rect 991 68 1064 95
rect 1184 219 1288 232
rect 1184 173 1213 219
rect 1259 173 1288 219
rect 1184 68 1288 173
rect 1408 127 1512 232
rect 1408 81 1437 127
rect 1483 81 1512 127
rect 1408 68 1512 81
rect 1632 219 1736 232
rect 1632 173 1661 219
rect 1707 173 1736 219
rect 1632 68 1736 173
rect 1856 127 1960 232
rect 1856 81 1885 127
rect 1931 81 1960 127
rect 1856 68 1960 81
rect 2080 219 2184 232
rect 2080 173 2109 219
rect 2155 173 2184 219
rect 2080 68 2184 173
rect 2304 127 2408 232
rect 2304 81 2333 127
rect 2379 81 2408 127
rect 2304 68 2408 81
rect 2528 219 2632 232
rect 2528 173 2557 219
rect 2603 173 2632 219
rect 2528 68 2632 173
rect 2752 127 2856 232
rect 2752 81 2781 127
rect 2827 81 2856 127
rect 2752 68 2856 81
rect 2976 219 3080 232
rect 2976 173 3005 219
rect 3051 173 3080 219
rect 2976 68 3080 173
rect 3200 127 3304 232
rect 3200 81 3229 127
rect 3275 81 3304 127
rect 3200 68 3304 81
rect 3424 219 3528 232
rect 3424 173 3453 219
rect 3499 173 3528 219
rect 3424 68 3528 173
rect 3648 127 3736 232
rect 3648 81 3677 127
rect 3723 81 3736 127
rect 3648 68 3736 81
rect 991 49 1004 68
rect 932 36 1004 49
<< mvpdiff >>
rect 84 602 172 716
rect 84 556 97 602
rect 143 556 172 602
rect 84 527 172 556
rect 272 698 376 716
rect 272 652 301 698
rect 347 652 376 698
rect 272 527 376 652
rect 476 678 660 716
rect 476 632 547 678
rect 593 632 660 678
rect 476 527 660 632
rect 760 586 848 716
rect 760 540 789 586
rect 835 540 848 586
rect 760 527 848 540
rect 1056 703 1144 716
rect 1056 657 1069 703
rect 1115 657 1144 703
rect 1056 481 1144 657
rect 1244 665 1348 716
rect 1244 525 1273 665
rect 1319 525 1348 665
rect 1244 481 1348 525
rect 1448 703 1552 716
rect 1448 657 1477 703
rect 1523 657 1552 703
rect 1448 481 1552 657
rect 1652 665 1756 716
rect 1652 525 1681 665
rect 1727 525 1756 665
rect 1652 481 1756 525
rect 1856 703 1960 716
rect 1856 657 1885 703
rect 1931 657 1960 703
rect 1856 481 1960 657
rect 2060 665 2164 716
rect 2060 525 2089 665
rect 2135 525 2164 665
rect 2060 481 2164 525
rect 2264 703 2368 716
rect 2264 657 2293 703
rect 2339 657 2368 703
rect 2264 481 2368 657
rect 2468 665 2572 716
rect 2468 525 2497 665
rect 2543 525 2572 665
rect 2468 481 2572 525
rect 2672 703 2776 716
rect 2672 657 2701 703
rect 2747 657 2776 703
rect 2672 481 2776 657
rect 2876 665 2980 716
rect 2876 525 2905 665
rect 2951 525 2980 665
rect 2876 481 2980 525
rect 3080 703 3184 716
rect 3080 657 3109 703
rect 3155 657 3184 703
rect 3080 481 3184 657
rect 3284 665 3388 716
rect 3284 525 3313 665
rect 3359 525 3388 665
rect 3284 481 3388 525
rect 3488 703 3576 716
rect 3488 657 3517 703
rect 3563 657 3576 703
rect 3488 481 3576 657
<< mvndiffc >>
rect 49 173 95 219
rect 273 82 319 128
rect 497 106 543 152
rect 765 228 811 274
rect 945 49 991 95
rect 1213 173 1259 219
rect 1437 81 1483 127
rect 1661 173 1707 219
rect 1885 81 1931 127
rect 2109 173 2155 219
rect 2333 81 2379 127
rect 2557 173 2603 219
rect 2781 81 2827 127
rect 3005 173 3051 219
rect 3229 81 3275 127
rect 3453 173 3499 219
rect 3677 81 3723 127
<< mvpdiffc >>
rect 97 556 143 602
rect 301 652 347 698
rect 547 632 593 678
rect 789 540 835 586
rect 1069 657 1115 703
rect 1273 525 1319 665
rect 1477 657 1523 703
rect 1681 525 1727 665
rect 1885 657 1931 703
rect 2089 525 2135 665
rect 2293 657 2339 703
rect 2497 525 2543 665
rect 2701 657 2747 703
rect 2905 525 2951 665
rect 3109 657 3155 703
rect 3313 525 3359 665
rect 3517 657 3563 703
<< polysilicon >>
rect 172 716 272 760
rect 376 716 476 760
rect 660 716 760 760
rect 1144 716 1244 760
rect 1348 716 1448 760
rect 1552 716 1652 760
rect 1756 716 1856 760
rect 1960 716 2060 760
rect 2164 716 2264 760
rect 2368 716 2468 760
rect 2572 716 2672 760
rect 2776 716 2876 760
rect 2980 716 3080 760
rect 3184 716 3284 760
rect 3388 716 3488 760
rect 172 413 272 527
rect 376 413 476 527
rect 660 493 760 527
rect 660 447 673 493
rect 719 447 760 493
rect 660 434 760 447
rect 1144 415 1244 481
rect 124 412 612 413
rect 124 366 185 412
rect 231 373 612 412
rect 1144 399 1171 415
rect 231 366 244 373
rect 124 232 244 366
rect 572 324 612 373
rect 1064 369 1171 399
rect 1217 399 1244 415
rect 1348 415 1448 481
rect 1348 399 1375 415
rect 1217 369 1375 399
rect 1421 399 1448 415
rect 1552 415 1652 481
rect 1552 399 1579 415
rect 1421 369 1579 399
rect 1625 399 1652 415
rect 1756 415 1856 481
rect 1756 399 1783 415
rect 1625 369 1783 399
rect 1829 369 1856 415
rect 1960 439 2060 481
rect 1960 393 2001 439
rect 2047 420 2060 439
rect 2164 439 2264 481
rect 2164 420 2190 439
rect 2047 393 2190 420
rect 2236 420 2264 439
rect 2368 439 2468 481
rect 2368 420 2395 439
rect 2236 393 2395 420
rect 2441 420 2468 439
rect 2572 420 2672 481
rect 2776 420 2876 481
rect 2980 439 3080 481
rect 2980 420 3021 439
rect 2441 393 3021 420
rect 3067 420 3080 439
rect 3184 439 3284 481
rect 3184 420 3225 439
rect 3067 393 3225 420
rect 3271 420 3284 439
rect 3388 439 3488 481
rect 3388 420 3429 439
rect 3271 393 3429 420
rect 3475 393 3488 439
rect 1960 380 3488 393
rect 1064 349 1856 369
rect 348 311 468 324
rect 348 265 385 311
rect 431 265 468 311
rect 348 232 468 265
rect 572 232 692 324
rect 1064 232 1184 349
rect 1288 232 1408 349
rect 1512 232 1632 349
rect 1736 232 1856 349
rect 1960 319 3648 332
rect 1960 273 1995 319
rect 2041 292 2219 319
rect 2041 273 2080 292
rect 1960 232 2080 273
rect 2184 273 2219 292
rect 2265 292 2444 319
rect 2265 273 2304 292
rect 2184 232 2304 273
rect 2408 273 2444 292
rect 2490 292 3094 319
rect 2490 273 2528 292
rect 2408 232 2528 273
rect 2632 232 2752 292
rect 2856 232 2976 292
rect 3080 273 3094 292
rect 3140 292 3318 319
rect 3140 273 3200 292
rect 3080 232 3200 273
rect 3304 273 3318 292
rect 3364 292 3541 319
rect 3364 273 3424 292
rect 3304 232 3424 273
rect 3528 273 3541 292
rect 3587 273 3648 319
rect 3528 232 3648 273
rect 124 24 244 68
rect 348 24 468 68
rect 572 24 692 68
rect 1064 24 1184 68
rect 1288 24 1408 68
rect 1512 24 1632 68
rect 1736 24 1856 68
rect 1960 24 2080 68
rect 2184 24 2304 68
rect 2408 24 2528 68
rect 2632 24 2752 68
rect 2856 24 2976 68
rect 3080 24 3200 68
rect 3304 24 3424 68
rect 3528 24 3648 68
<< polycontact >>
rect 673 447 719 493
rect 185 366 231 412
rect 1171 369 1217 415
rect 1375 369 1421 415
rect 1579 369 1625 415
rect 1783 369 1829 415
rect 2001 393 2047 439
rect 2190 393 2236 439
rect 2395 393 2441 439
rect 3021 393 3067 439
rect 3225 393 3271 439
rect 3429 393 3475 439
rect 385 265 431 311
rect 1995 273 2041 319
rect 2219 273 2265 319
rect 2444 273 2490 319
rect 3094 273 3140 319
rect 3318 273 3364 319
rect 3541 273 3587 319
<< metal1 >>
rect 0 724 3808 844
rect 290 698 358 724
rect 290 652 301 698
rect 347 652 358 698
rect 1058 703 1126 724
rect 536 632 547 678
rect 593 632 965 678
rect 1058 657 1069 703
rect 1115 657 1126 703
rect 1466 703 1534 724
rect 1273 665 1319 676
rect 84 556 97 602
rect 143 556 431 602
rect 385 504 431 556
rect 778 540 789 586
rect 835 540 846 586
rect 385 493 730 504
rect 385 447 673 493
rect 719 447 730 493
rect 109 412 335 437
rect 109 366 185 412
rect 231 366 335 412
rect 109 355 335 366
rect 385 311 431 447
rect 778 401 846 540
rect 38 219 431 265
rect 641 355 846 401
rect 919 552 965 632
rect 919 525 1273 552
rect 1466 657 1477 703
rect 1523 657 1534 703
rect 1874 703 1942 724
rect 1681 665 1727 676
rect 1319 525 1681 552
rect 1874 657 1885 703
rect 1931 657 1942 703
rect 2282 703 2350 724
rect 2078 665 2146 676
rect 1727 525 1997 552
rect 919 506 1997 525
rect 38 173 49 219
rect 95 173 106 219
rect 38 170 106 173
rect 641 152 687 355
rect 919 309 965 506
rect 1951 439 1997 506
rect 2078 525 2089 665
rect 2135 553 2146 665
rect 2282 657 2293 703
rect 2339 657 2350 703
rect 2690 703 2758 724
rect 2486 665 2554 676
rect 2486 553 2497 665
rect 2135 525 2497 553
rect 2543 553 2554 665
rect 2690 657 2701 703
rect 2747 657 2758 703
rect 3098 703 3166 724
rect 2894 665 2962 676
rect 2894 553 2905 665
rect 2543 525 2905 553
rect 2951 553 2962 665
rect 3098 657 3109 703
rect 3155 657 3166 703
rect 3506 703 3574 724
rect 3302 665 3370 676
rect 3302 553 3313 665
rect 2951 525 3313 553
rect 3359 525 3370 665
rect 3506 657 3517 703
rect 3563 657 3574 703
rect 2078 485 3370 525
rect 1015 415 1886 424
rect 1015 369 1171 415
rect 1217 369 1375 415
rect 1421 369 1579 415
rect 1625 369 1783 415
rect 1829 369 1886 415
rect 1951 393 2001 439
rect 2047 393 2190 439
rect 2236 393 2395 439
rect 2441 393 2452 439
rect 1015 360 1886 369
rect 754 274 965 309
rect 754 228 765 274
rect 811 263 965 274
rect 1951 273 1995 319
rect 2041 273 2219 319
rect 2265 273 2444 319
rect 2490 273 2504 319
rect 811 228 822 263
rect 1951 219 1997 273
rect 2684 227 2814 485
rect 3010 393 3021 439
rect 3067 393 3225 439
rect 3271 393 3429 439
rect 3475 393 3486 439
rect 3083 273 3094 319
rect 3140 273 3318 319
rect 3364 273 3541 319
rect 3587 273 3598 319
rect 1139 187 1213 219
rect 843 173 1213 187
rect 1259 173 1661 219
rect 1707 173 1997 219
rect 2080 219 3510 227
rect 2080 173 2109 219
rect 2155 173 2557 219
rect 2603 173 3005 219
rect 3051 173 3453 219
rect 3499 173 3510 219
rect 843 152 1189 173
rect 262 128 330 131
rect 262 82 273 128
rect 319 82 330 128
rect 478 106 497 152
rect 543 141 1189 152
rect 543 106 888 141
rect 262 60 330 82
rect 934 60 945 95
rect 0 49 945 60
rect 991 60 1002 95
rect 1426 81 1437 127
rect 1483 81 1494 127
rect 1426 60 1494 81
rect 1874 81 1885 127
rect 1931 81 1942 127
rect 1874 60 1942 81
rect 2322 81 2333 127
rect 2379 81 2390 127
rect 2322 60 2390 81
rect 2770 81 2781 127
rect 2827 81 2838 127
rect 2770 60 2838 81
rect 3218 81 3229 127
rect 3275 81 3286 127
rect 3218 60 3286 81
rect 3666 81 3677 127
rect 3723 81 3734 127
rect 3666 60 3734 81
rect 991 49 3808 60
rect 0 -60 3808 49
<< labels >>
flabel metal1 s 3302 553 3370 676 0 FreeSans 400 0 0 0 Z
port 3 nsew default output
flabel metal1 s 109 355 335 437 0 FreeSans 600 0 0 0 EN
port 1 nsew default input
flabel metal1 s 1015 360 1886 424 0 FreeSans 400 0 0 0 I
port 2 nsew default input
flabel metal1 s 262 127 330 131 0 FreeSans 400 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel metal1 s 0 724 3808 844 0 FreeSans 400 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 5 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 6 nsew ground bidirectional
rlabel metal1 s 2894 553 2962 676 1 Z
port 3 nsew default output
rlabel metal1 s 2486 553 2554 676 1 Z
port 3 nsew default output
rlabel metal1 s 2078 553 2146 676 1 Z
port 3 nsew default output
rlabel metal1 s 2078 485 3370 553 1 Z
port 3 nsew default output
rlabel metal1 s 2684 227 2814 485 1 Z
port 3 nsew default output
rlabel metal1 s 2080 173 3510 227 1 Z
port 3 nsew default output
rlabel metal1 s 3506 657 3574 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3098 657 3166 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2690 657 2758 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2282 657 2350 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1874 657 1942 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1466 657 1534 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1058 657 1126 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 290 657 358 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 290 652 358 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3666 95 3734 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3218 95 3286 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2770 95 2838 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2322 95 2390 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1874 95 1942 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1426 95 1494 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 95 330 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3666 60 3734 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3218 60 3286 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2770 60 2838 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2322 60 2390 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1874 60 1942 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1426 60 1494 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 934 60 1002 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 60 330 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3808 60 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3808 784
string GDS_END 1417210
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1408920
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
