magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 377 5462 870
rect -86 352 1291 377
rect 1974 352 2726 377
rect 3918 352 5462 377
<< pwell >>
rect 1291 352 1974 377
rect 2726 352 3918 377
rect -86 -86 5462 352
<< metal1 >>
rect 0 724 5376 844
rect 252 569 320 724
rect 1075 577 1121 724
rect 1518 670 1586 724
rect 2602 689 2670 724
rect 3240 689 3312 724
rect 141 119 206 430
rect 273 60 319 228
rect 365 119 430 430
rect 681 353 878 438
rect 1026 353 1326 431
rect 1110 60 1156 205
rect 1573 60 1619 209
rect 4093 583 4139 724
rect 2756 60 2828 183
rect 4121 242 4228 439
rect 4526 594 4594 724
rect 4505 353 4686 431
rect 5011 506 5057 724
rect 5172 501 5264 676
rect 5172 441 5311 501
rect 4372 60 4440 215
rect 5251 232 5311 441
rect 5011 60 5057 232
rect 5151 131 5311 232
rect 0 -60 5376 60
<< obsm1 >>
rect 49 523 95 608
rect 654 549 1015 595
rect 1217 632 1472 678
rect 969 531 1015 549
rect 1217 531 1263 632
rect 1426 624 1472 632
rect 1641 632 1967 678
rect 2253 643 2556 678
rect 2716 643 3194 678
rect 3358 643 3655 678
rect 2253 632 3655 643
rect 1641 624 1687 632
rect 1426 578 1687 624
rect 49 477 571 523
rect 969 484 1263 531
rect 1322 524 1368 578
rect 1322 477 1707 524
rect 49 156 95 477
rect 525 307 571 477
rect 926 307 972 350
rect 525 261 972 307
rect 1018 252 1248 298
rect 1389 255 1435 477
rect 1661 382 1707 477
rect 1777 407 1823 569
rect 1921 497 1967 632
rect 2510 597 2762 632
rect 3148 597 3404 632
rect 2160 459 2206 574
rect 2336 551 2440 555
rect 2832 551 2920 556
rect 2336 505 2920 551
rect 2992 551 3080 556
rect 3472 551 3558 556
rect 2992 505 3558 551
rect 2160 413 3181 459
rect 1777 360 2081 407
rect 1018 215 1064 252
rect 650 169 1064 215
rect 1202 152 1248 252
rect 1367 198 1435 255
rect 1481 259 1736 306
rect 1481 152 1527 259
rect 1202 106 1527 152
rect 1690 152 1736 259
rect 1830 198 1898 360
rect 1985 152 2031 196
rect 1690 106 2031 152
rect 2209 124 2255 413
rect 3265 367 3333 505
rect 3609 407 3655 632
rect 3705 632 4047 678
rect 2325 275 2371 340
rect 2459 321 3333 367
rect 3705 361 3751 632
rect 3909 445 3955 567
rect 4001 537 4047 632
rect 4185 632 4462 678
rect 4185 537 4231 632
rect 4001 491 4231 537
rect 2325 229 2920 275
rect 2874 152 2920 229
rect 3265 198 3333 321
rect 3388 152 3434 349
rect 3489 315 3751 361
rect 3797 399 4037 445
rect 3489 198 3557 315
rect 3797 244 3843 399
rect 3714 198 3843 244
rect 3889 152 3935 353
rect 2874 106 3935 152
rect 3991 192 4037 399
rect 4286 431 4354 586
rect 4416 548 4462 632
rect 4640 632 4898 678
rect 4640 548 4686 632
rect 4416 502 4686 548
rect 4280 385 4354 431
rect 4280 192 4326 385
rect 4413 307 4459 440
rect 4738 307 4806 586
rect 4852 412 4898 632
rect 4867 320 5156 366
rect 4867 307 4913 320
rect 4413 261 4913 307
rect 3991 143 4326 192
rect 4867 156 4913 261
<< labels >>
rlabel metal1 s 681 353 878 438 6 D
port 1 nsew default input
rlabel metal1 s 4505 353 4686 431 6 RN
port 2 nsew default input
rlabel metal1 s 141 119 206 430 6 SE
port 3 nsew default input
rlabel metal1 s 4121 242 4228 439 6 SETN
port 4 nsew default input
rlabel metal1 s 365 119 430 430 6 SI
port 5 nsew default input
rlabel metal1 s 1026 353 1326 431 6 CLK
port 6 nsew clock input
rlabel metal1 s 5151 131 5311 232 6 Q
port 7 nsew default output
rlabel metal1 s 5251 232 5311 441 6 Q
port 7 nsew default output
rlabel metal1 s 5172 441 5311 501 6 Q
port 7 nsew default output
rlabel metal1 s 5172 501 5264 676 6 Q
port 7 nsew default output
rlabel metal1 s 5011 506 5057 724 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4526 594 4594 724 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4093 583 4139 724 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3240 689 3312 724 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 2602 689 2670 724 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1518 670 1586 724 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1075 577 1121 724 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 252 569 320 724 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 724 5376 844 6 VDD
port 8 nsew power bidirectional abutment
rlabel nwell s 3918 352 5462 377 6 VNW
port 9 nsew power bidirectional
rlabel nwell s 1974 352 2726 377 6 VNW
port 9 nsew power bidirectional
rlabel nwell s -86 352 1291 377 6 VNW
port 9 nsew power bidirectional
rlabel nwell s -86 377 5462 870 6 VNW
port 9 nsew power bidirectional
rlabel pwell s -86 -86 5462 352 6 VPW
port 10 nsew ground bidirectional
rlabel pwell s 2726 352 3918 377 6 VPW
port 10 nsew ground bidirectional
rlabel pwell s 1291 352 1974 377 6 VPW
port 10 nsew ground bidirectional
rlabel metal1 s 0 -60 5376 60 8 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 5011 60 5057 232 6 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 4372 60 4440 215 6 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 2756 60 2828 183 6 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 1573 60 1619 209 6 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 1110 60 1156 205 6 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 273 60 319 228 6 VSS
port 11 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 5376 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 256132
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 244294
<< end >>
