magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 377 3110 870
rect -86 352 228 377
rect 2011 352 3110 377
<< pwell >>
rect -86 -86 3110 352
<< mvnmos >>
rect 124 68 244 232
rect 392 93 512 257
rect 616 93 736 257
rect 840 93 960 257
rect 1064 93 1184 257
rect 1288 93 1408 257
rect 1512 93 1632 257
rect 1736 93 1856 257
rect 2004 68 2124 232
rect 2228 68 2348 232
rect 2452 68 2572 232
rect 2676 68 2796 232
<< mvpmos >>
rect 124 497 224 716
rect 412 497 512 716
rect 616 497 716 716
rect 860 497 960 716
rect 1064 497 1164 716
rect 1308 497 1408 716
rect 1512 497 1612 716
rect 1736 497 1836 716
rect 2044 525 2144 716
rect 2248 525 2348 716
rect 2452 525 2552 716
rect 2656 525 2756 716
<< mvndiff >>
rect 304 244 392 257
rect 304 232 317 244
rect 36 152 124 232
rect 36 106 49 152
rect 95 106 124 152
rect 36 68 124 106
rect 244 198 317 232
rect 363 198 392 244
rect 244 93 392 198
rect 512 152 616 257
rect 512 106 541 152
rect 587 106 616 152
rect 512 93 616 106
rect 736 244 840 257
rect 736 198 765 244
rect 811 198 840 244
rect 736 93 840 198
rect 960 152 1064 257
rect 960 106 989 152
rect 1035 106 1064 152
rect 960 93 1064 106
rect 1184 244 1288 257
rect 1184 198 1213 244
rect 1259 198 1288 244
rect 1184 93 1288 198
rect 1408 152 1512 257
rect 1408 106 1437 152
rect 1483 106 1512 152
rect 1408 93 1512 106
rect 1632 244 1736 257
rect 1632 198 1661 244
rect 1707 198 1736 244
rect 1632 93 1736 198
rect 1856 232 1936 257
rect 1856 152 2004 232
rect 1856 106 1885 152
rect 1931 106 2004 152
rect 1856 93 2004 106
rect 244 68 324 93
rect 1924 68 2004 93
rect 2124 171 2228 232
rect 2124 125 2153 171
rect 2199 125 2228 171
rect 2124 68 2228 125
rect 2348 171 2452 232
rect 2348 125 2377 171
rect 2423 125 2452 171
rect 2348 68 2452 125
rect 2572 171 2676 232
rect 2572 125 2601 171
rect 2647 125 2676 171
rect 2572 68 2676 125
rect 2796 171 2884 232
rect 2796 125 2825 171
rect 2871 125 2884 171
rect 2796 68 2884 125
<< mvpdiff >>
rect 36 639 124 716
rect 36 593 49 639
rect 95 593 124 639
rect 36 497 124 593
rect 224 497 412 716
rect 512 639 616 716
rect 512 593 541 639
rect 587 593 616 639
rect 512 497 616 593
rect 716 497 860 716
rect 960 703 1064 716
rect 960 657 989 703
rect 1035 657 1064 703
rect 960 497 1064 657
rect 1164 497 1308 716
rect 1408 639 1512 716
rect 1408 593 1437 639
rect 1483 593 1512 639
rect 1408 497 1512 593
rect 1612 497 1736 716
rect 1836 639 2044 716
rect 1836 593 1969 639
rect 2015 593 2044 639
rect 1836 525 2044 593
rect 2144 639 2248 716
rect 2144 593 2173 639
rect 2219 593 2248 639
rect 2144 525 2248 593
rect 2348 639 2452 716
rect 2348 593 2377 639
rect 2423 593 2452 639
rect 2348 525 2452 593
rect 2552 639 2656 716
rect 2552 593 2581 639
rect 2627 593 2656 639
rect 2552 525 2656 593
rect 2756 639 2844 716
rect 2756 593 2785 639
rect 2831 593 2844 639
rect 2756 525 2844 593
rect 1836 497 1916 525
<< mvndiffc >>
rect 49 106 95 152
rect 317 198 363 244
rect 541 106 587 152
rect 765 198 811 244
rect 989 106 1035 152
rect 1213 198 1259 244
rect 1437 106 1483 152
rect 1661 198 1707 244
rect 1885 106 1931 152
rect 2153 125 2199 171
rect 2377 125 2423 171
rect 2601 125 2647 171
rect 2825 125 2871 171
<< mvpdiffc >>
rect 49 593 95 639
rect 541 593 587 639
rect 989 657 1035 703
rect 1437 593 1483 639
rect 1969 593 2015 639
rect 2173 593 2219 639
rect 2377 593 2423 639
rect 2581 593 2627 639
rect 2785 593 2831 639
<< polysilicon >>
rect 124 716 224 760
rect 412 716 512 760
rect 616 716 716 760
rect 860 716 960 760
rect 1064 716 1164 760
rect 1308 716 1408 760
rect 1512 716 1612 760
rect 1736 716 1836 760
rect 2044 716 2144 760
rect 2248 716 2348 760
rect 2452 716 2552 760
rect 2656 716 2756 760
rect 124 415 224 497
rect 124 369 145 415
rect 191 408 224 415
rect 412 414 512 497
rect 191 369 244 408
rect 412 394 439 414
rect 124 232 244 369
rect 392 368 439 394
rect 485 394 512 414
rect 616 414 716 497
rect 616 394 643 414
rect 485 368 643 394
rect 689 394 716 414
rect 860 428 960 497
rect 860 394 887 428
rect 689 368 736 394
rect 392 348 736 368
rect 392 257 512 348
rect 616 257 736 348
rect 840 382 887 394
rect 933 394 960 428
rect 1064 428 1164 497
rect 1064 394 1091 428
rect 933 382 1091 394
rect 1137 394 1164 428
rect 1308 394 1408 497
rect 1512 394 1612 497
rect 1736 428 1836 497
rect 1137 382 1184 394
rect 840 348 1184 382
rect 840 257 960 348
rect 1064 257 1184 348
rect 1288 348 1632 394
rect 1288 336 1408 348
rect 1288 290 1325 336
rect 1371 290 1408 336
rect 1288 257 1408 290
rect 1512 336 1632 348
rect 1512 290 1549 336
rect 1595 290 1632 336
rect 1512 257 1632 290
rect 1736 382 1763 428
rect 1809 394 1836 428
rect 2044 415 2144 525
rect 2044 394 2071 415
rect 1809 382 1856 394
rect 1736 257 1856 382
rect 2004 369 2071 394
rect 2117 394 2144 415
rect 2248 415 2348 525
rect 2248 394 2275 415
rect 2117 369 2275 394
rect 2321 394 2348 415
rect 2452 415 2552 525
rect 2452 394 2479 415
rect 2321 369 2479 394
rect 2525 394 2552 415
rect 2656 415 2756 525
rect 2656 394 2683 415
rect 2525 369 2683 394
rect 2729 394 2756 415
rect 2729 369 2796 394
rect 2004 348 2796 369
rect 2004 232 2124 348
rect 2228 232 2348 348
rect 2452 232 2572 348
rect 2676 232 2796 348
rect 124 24 244 68
rect 392 24 512 93
rect 616 24 736 93
rect 840 24 960 93
rect 1064 24 1184 93
rect 1288 24 1408 93
rect 1512 24 1632 93
rect 1736 24 1856 93
rect 2004 24 2124 68
rect 2228 24 2348 68
rect 2452 24 2572 68
rect 2676 24 2796 68
<< polycontact >>
rect 145 369 191 415
rect 439 368 485 414
rect 643 368 689 414
rect 887 382 933 428
rect 1091 382 1137 428
rect 1325 290 1371 336
rect 1549 290 1595 336
rect 1763 382 1809 428
rect 2071 369 2117 415
rect 2275 369 2321 415
rect 2479 369 2525 415
rect 2683 369 2729 415
<< metal1 >>
rect 0 724 3024 844
rect 49 639 95 724
rect 978 703 1046 724
rect 978 657 989 703
rect 1035 657 1046 703
rect 49 582 95 593
rect 217 639 928 648
rect 217 593 541 639
rect 587 611 928 639
rect 1096 639 1923 648
rect 1096 611 1437 639
rect 587 593 1437 611
rect 1483 593 1923 639
rect 217 584 1923 593
rect 882 565 1142 584
rect 1877 536 1923 584
rect 1969 639 2015 724
rect 1969 582 2015 593
rect 2173 639 2219 650
rect 2173 536 2219 593
rect 2377 639 2423 724
rect 2377 582 2423 593
rect 2581 639 2627 650
rect 2581 536 2627 593
rect 2785 639 2831 724
rect 2785 582 2831 593
rect 136 472 820 536
rect 136 415 200 472
rect 774 428 820 472
rect 1877 472 2627 536
rect 136 369 145 415
rect 191 369 200 415
rect 136 339 200 369
rect 306 414 716 424
rect 306 368 439 414
rect 485 368 643 414
rect 689 368 716 414
rect 774 382 887 428
rect 933 382 1091 428
rect 1137 382 1763 428
rect 1809 382 1828 428
rect 306 360 716 368
rect 670 336 716 360
rect 670 290 1325 336
rect 1371 290 1549 336
rect 1595 290 1614 336
rect 1877 244 1923 472
rect 2004 415 2910 424
rect 2004 369 2071 415
rect 2117 369 2275 415
rect 2321 369 2479 415
rect 2525 369 2683 415
rect 2729 369 2910 415
rect 2004 360 2910 369
rect 304 198 317 244
rect 363 198 765 244
rect 811 198 1213 244
rect 1259 198 1661 244
rect 1707 198 1923 244
rect 2030 232 2871 278
rect 2030 152 2076 232
rect 36 106 49 152
rect 95 106 541 152
rect 587 106 989 152
rect 1035 106 1437 152
rect 1483 106 1885 152
rect 1931 106 2076 152
rect 2153 171 2199 182
rect 2153 60 2199 125
rect 2377 171 2423 232
rect 2377 114 2423 125
rect 2601 171 2647 182
rect 2601 60 2647 125
rect 2825 171 2871 232
rect 2825 114 2871 125
rect 0 -60 3024 60
<< labels >>
flabel metal1 s 2004 360 2910 424 0 FreeSans 400 0 0 0 B
port 3 nsew default input
flabel metal1 s 0 724 3024 844 0 FreeSans 400 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 2601 60 2647 182 0 FreeSans 400 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel metal1 s 306 360 716 424 0 FreeSans 400 0 0 0 A1
port 1 nsew default input
flabel metal1 s 2581 648 2627 650 0 FreeSans 400 0 0 0 ZN
port 4 nsew default output
flabel metal1 s 136 472 820 536 0 FreeSans 400 0 0 0 A2
port 2 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 6 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 670 336 716 360 1 A1
port 1 nsew default input
rlabel metal1 s 670 290 1614 336 1 A1
port 1 nsew default input
rlabel metal1 s 774 428 820 472 1 A2
port 2 nsew default input
rlabel metal1 s 136 428 200 472 1 A2
port 2 nsew default input
rlabel metal1 s 774 382 1828 428 1 A2
port 2 nsew default input
rlabel metal1 s 136 382 200 428 1 A2
port 2 nsew default input
rlabel metal1 s 136 339 200 382 1 A2
port 2 nsew default input
rlabel metal1 s 2173 648 2219 650 1 ZN
port 4 nsew default output
rlabel metal1 s 2581 611 2627 648 1 ZN
port 4 nsew default output
rlabel metal1 s 2173 611 2219 648 1 ZN
port 4 nsew default output
rlabel metal1 s 1096 611 1923 648 1 ZN
port 4 nsew default output
rlabel metal1 s 217 611 928 648 1 ZN
port 4 nsew default output
rlabel metal1 s 2581 584 2627 611 1 ZN
port 4 nsew default output
rlabel metal1 s 2173 584 2219 611 1 ZN
port 4 nsew default output
rlabel metal1 s 217 584 1923 611 1 ZN
port 4 nsew default output
rlabel metal1 s 2581 565 2627 584 1 ZN
port 4 nsew default output
rlabel metal1 s 2173 565 2219 584 1 ZN
port 4 nsew default output
rlabel metal1 s 1877 565 1923 584 1 ZN
port 4 nsew default output
rlabel metal1 s 882 565 1142 584 1 ZN
port 4 nsew default output
rlabel metal1 s 2581 536 2627 565 1 ZN
port 4 nsew default output
rlabel metal1 s 2173 536 2219 565 1 ZN
port 4 nsew default output
rlabel metal1 s 1877 536 1923 565 1 ZN
port 4 nsew default output
rlabel metal1 s 1877 472 2627 536 1 ZN
port 4 nsew default output
rlabel metal1 s 1877 244 1923 472 1 ZN
port 4 nsew default output
rlabel metal1 s 304 198 1923 244 1 ZN
port 4 nsew default output
rlabel metal1 s 2785 657 2831 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2377 657 2423 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1969 657 2015 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 978 657 1046 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 49 657 95 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2785 582 2831 657 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2377 582 2423 657 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1969 582 2015 657 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 49 582 95 657 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2153 60 2199 182 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3024 60 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3024 784
string GDS_END 20336
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 14704
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
