magic
tech gf180mcuA
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -1730 9497 11766 10481
rect -1730 -15 -500 9497
rect 10573 -15 11766 9497
rect -1730 -583 11766 -15
<< psubdiff >>
rect -458 8756 10536 9430
rect -458 8300 -118 8756
rect -458 54 -396 8300
rect -150 322 -118 8300
rect 10146 8322 10536 8756
rect 10146 8300 10541 8322
rect 10146 322 10173 8300
rect -150 300 10173 322
rect -150 54 11 300
rect 10057 54 10173 300
rect 10519 54 10541 8300
rect -458 32 10541 54
<< nsubdiff >>
rect -1647 10376 11683 10398
rect -1647 10330 -436 10376
rect 10510 10330 11683 10376
rect -1647 10272 11683 10330
rect -1647 10226 -436 10272
rect 10510 10226 11683 10272
rect -1647 10168 11683 10226
rect -1647 10122 -436 10168
rect 10510 10122 11683 10168
rect -1647 10064 11683 10122
rect -1647 10018 -436 10064
rect 10510 10018 11683 10064
rect -1647 9960 11683 10018
rect -1647 9914 -436 9960
rect 10510 9914 11683 9960
rect -1647 9856 11683 9914
rect -1647 9810 -436 9856
rect 10510 9810 11683 9856
rect -1647 9752 11683 9810
rect -1647 9706 -436 9752
rect 10510 9706 11683 9752
rect -1647 9648 11683 9706
rect -1647 9602 -436 9648
rect 10510 9602 11683 9648
rect -1647 9580 11683 9602
rect -1647 8368 -583 9580
rect -1647 -478 -1587 8368
rect -1541 -478 -1483 8368
rect -1437 -478 -1379 8368
rect -1333 -478 -1275 8368
rect -1229 -478 -1171 8368
rect -1125 -478 -1067 8368
rect -1021 -478 -963 8368
rect -917 -478 -859 8368
rect -813 -478 -755 8368
rect -709 -478 -651 8368
rect -605 -98 -583 8368
rect 10656 8368 11683 9580
rect 10656 -98 10678 8368
rect -605 -120 10678 -98
rect -605 -166 -436 -120
rect 10510 -166 10678 -120
rect -605 -224 10678 -166
rect -605 -270 -436 -224
rect 10510 -270 10678 -224
rect -605 -328 10678 -270
rect -605 -374 -436 -328
rect 10510 -374 10678 -328
rect -605 -432 10678 -374
rect -605 -478 -436 -432
rect 10510 -478 10678 -432
rect 10724 -478 10782 8368
rect 10828 -478 10886 8368
rect 10932 -478 10990 8368
rect 11036 -478 11094 8368
rect 11140 -478 11198 8368
rect 11244 -478 11302 8368
rect 11348 -478 11406 8368
rect 11452 -478 11510 8368
rect 11556 -478 11614 8368
rect 11660 -478 11683 8368
rect -1647 -500 11683 -478
<< psubdiffcont >>
rect -396 54 -150 8300
rect 11 54 10057 300
rect 10173 54 10519 8300
<< nsubdiffcont >>
rect -436 10330 10510 10376
rect -436 10226 10510 10272
rect -436 10122 10510 10168
rect -436 10018 10510 10064
rect -436 9914 10510 9960
rect -436 9810 10510 9856
rect -436 9706 10510 9752
rect -436 9602 10510 9648
rect -1587 -478 -1541 8368
rect -1483 -478 -1437 8368
rect -1379 -478 -1333 8368
rect -1275 -478 -1229 8368
rect -1171 -478 -1125 8368
rect -1067 -478 -1021 8368
rect -963 -478 -917 8368
rect -859 -478 -813 8368
rect -755 -478 -709 8368
rect -651 -478 -605 8368
rect -436 -166 10510 -120
rect -436 -270 10510 -224
rect -436 -374 10510 -328
rect -436 -478 10510 -432
rect 10678 -478 10724 8368
rect 10782 -478 10828 8368
rect 10886 -478 10932 8368
rect 10990 -478 11036 8368
rect 11094 -478 11140 8368
rect 11198 -478 11244 8368
rect 11302 -478 11348 8368
rect 11406 -478 11452 8368
rect 11510 -478 11556 8368
rect 11614 -478 11660 8368
<< metal1 >>
rect -447 10376 10521 10387
rect -447 10330 -436 10376
rect 10510 10330 10521 10376
rect -447 10272 10521 10330
rect -447 10226 -436 10272
rect 10510 10226 10521 10272
rect -447 10168 10521 10226
rect -447 10122 -436 10168
rect 10510 10122 10521 10168
rect -447 10064 10521 10122
rect -447 10018 -436 10064
rect 10510 10018 10521 10064
rect -447 9960 10521 10018
rect -447 9914 -436 9960
rect 10510 9914 10521 9960
rect -447 9856 10521 9914
rect -447 9810 -436 9856
rect 10510 9810 10521 9856
rect -447 9752 10521 9810
rect -447 9706 -436 9752
rect 10510 9706 10521 9752
rect -447 9648 10521 9706
rect -447 9602 -436 9648
rect 10510 9602 10521 9648
rect -447 9591 10521 9602
rect -1598 8368 -594 8388
rect -1598 -478 -1587 8368
rect -1541 -478 -1483 8368
rect -1437 -478 -1379 8368
rect -1333 -478 -1275 8368
rect -1229 -478 -1171 8368
rect -1125 -478 -1067 8368
rect -1021 -478 -963 8368
rect -917 -478 -859 8368
rect -813 -478 -755 8368
rect -709 -478 -651 8368
rect -605 -109 -594 8368
rect -457 8300 111 8396
rect -457 54 -396 8300
rect -150 311 111 8300
rect 9962 8300 10530 8397
rect 9962 311 10173 8300
rect -150 300 10173 311
rect -150 54 11 300
rect 10057 54 10173 300
rect 10519 54 10530 8300
rect -457 43 10530 54
rect 10666 8368 11670 8410
rect 10666 -109 10678 8368
rect -605 -120 10678 -109
rect -605 -166 -436 -120
rect 10510 -166 10678 -120
rect -605 -224 10678 -166
rect -605 -270 -436 -224
rect 10510 -270 10678 -224
rect -605 -328 10678 -270
rect -605 -374 -436 -328
rect 10510 -374 10678 -328
rect -605 -432 10678 -374
rect -605 -478 -436 -432
rect 10510 -478 10678 -432
rect 10724 -478 10782 8368
rect 10828 -478 10886 8368
rect 10932 -478 10990 8368
rect 11036 -478 11094 8368
rect 11140 -478 11198 8368
rect 11244 -478 11302 8368
rect 11348 -478 11406 8368
rect 11452 -478 11510 8368
rect 11556 -478 11614 8368
rect 11660 -478 11670 8368
rect -1598 -489 11670 -478
use M1_NWELL_CDNS_40661956134476  M1_NWELL_CDNS_40661956134476_0
timestamp 1698431365
transform 1 0 5037 0 1 -299
box 0 0 1 1
use M1_NWELL_CDNS_40661956134477  M1_NWELL_CDNS_40661956134477_0
timestamp 1698431365
transform 1 0 5037 0 1 9989
box 0 0 1 1
use M1_PSUB_CDNS_40661956134475  M1_PSUB_CDNS_40661956134475_0
timestamp 1698431365
transform 1 0 -273 0 1 4177
box 0 0 1 1
use M1_PSUB_CDNS_40661956134478  M1_PSUB_CDNS_40661956134478_0
timestamp 1698431365
transform 1 0 10346 0 1 4177
box 0 0 1 1
use M1_PSUB_CDNS_40661956134479  M1_PSUB_CDNS_40661956134479_0
timestamp 1698431365
transform 0 -1 5034 1 0 177
box 0 0 1 1
<< properties >>
string GDS_END 2841230
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 2702260
<< end >>
