magic
tech gf180mcuD
magscale 1 10
timestamp 1698431365
<< metal1 >>
rect 3621 1336 3945 1348
rect 3621 1284 3633 1336
rect 3685 1284 3757 1336
rect 3809 1284 3881 1336
rect 3933 1284 3945 1336
rect 3621 1212 3945 1284
rect 3621 1160 3633 1212
rect 3685 1160 3757 1212
rect 3809 1160 3881 1212
rect 3933 1160 3945 1212
rect 3621 1088 3945 1160
rect 3621 1036 3633 1088
rect 3685 1036 3757 1088
rect 3809 1036 3881 1088
rect 3933 1036 3945 1088
rect 3621 964 3945 1036
rect 3621 912 3633 964
rect 3685 912 3757 964
rect 3809 912 3881 964
rect 3933 912 3945 964
rect 3621 840 3945 912
rect 3621 788 3633 840
rect 3685 788 3757 840
rect 3809 788 3881 840
rect 3933 788 3945 840
rect 3621 716 3945 788
rect 3621 664 3633 716
rect 3685 664 3757 716
rect 3809 664 3881 716
rect 3933 664 3945 716
rect 3621 652 3945 664
rect 4721 436 5045 448
rect 4721 384 4733 436
rect 4785 384 4857 436
rect 4909 384 4981 436
rect 5033 384 5045 436
rect 4721 312 5045 384
rect 4721 260 4733 312
rect 4785 260 4857 312
rect 4909 260 4981 312
rect 5033 260 5045 312
rect 4721 188 5045 260
rect 4721 136 4733 188
rect 4785 136 4857 188
rect 4909 136 4981 188
rect 5033 150 5045 188
rect 5033 136 5611 150
rect 4721 64 5611 136
rect 4721 12 4733 64
rect 4785 12 4857 64
rect 4909 12 4981 64
rect 5033 50 5611 64
rect 5033 12 5045 50
rect 4721 -60 5045 12
rect 4721 -112 4733 -60
rect 4785 -112 4857 -60
rect 4909 -112 4981 -60
rect 5033 -112 5045 -60
rect 4721 -184 5045 -112
rect 4721 -236 4733 -184
rect 4785 -236 4857 -184
rect 4909 -236 4981 -184
rect 5033 -236 5045 -184
rect 4721 -248 5045 -236
<< via1 >>
rect 3633 1284 3685 1336
rect 3757 1284 3809 1336
rect 3881 1284 3933 1336
rect 3633 1160 3685 1212
rect 3757 1160 3809 1212
rect 3881 1160 3933 1212
rect 3633 1036 3685 1088
rect 3757 1036 3809 1088
rect 3881 1036 3933 1088
rect 3633 912 3685 964
rect 3757 912 3809 964
rect 3881 912 3933 964
rect 3633 788 3685 840
rect 3757 788 3809 840
rect 3881 788 3933 840
rect 3633 664 3685 716
rect 3757 664 3809 716
rect 3881 664 3933 716
rect 4733 384 4785 436
rect 4857 384 4909 436
rect 4981 384 5033 436
rect 4733 260 4785 312
rect 4857 260 4909 312
rect 4981 260 5033 312
rect 4733 136 4785 188
rect 4857 136 4909 188
rect 4981 136 5033 188
rect 4733 12 4785 64
rect 4857 12 4909 64
rect 4981 12 5033 64
rect 4733 -112 4785 -60
rect 4857 -112 4909 -60
rect 4981 -112 5033 -60
rect 4733 -236 4785 -184
rect 4857 -236 4909 -184
rect 4981 -236 5033 -184
<< metal2 >>
rect 3621 1338 3945 1348
rect 3621 1282 3631 1338
rect 3687 1282 3755 1338
rect 3811 1282 3879 1338
rect 3935 1282 3945 1338
rect 3621 1214 3945 1282
rect 3621 1158 3631 1214
rect 3687 1158 3755 1214
rect 3811 1158 3879 1214
rect 3935 1158 3945 1214
rect 3621 1090 3945 1158
rect 3621 1034 3631 1090
rect 3687 1034 3755 1090
rect 3811 1034 3879 1090
rect 3935 1034 3945 1090
rect 3621 966 3945 1034
rect 3621 910 3631 966
rect 3687 910 3755 966
rect 3811 910 3879 966
rect 3935 910 3945 966
rect 3621 842 3945 910
rect 3621 786 3631 842
rect 3687 786 3755 842
rect 3811 786 3879 842
rect 3935 786 3945 842
rect 3621 718 3945 786
rect 3621 662 3631 718
rect 3687 662 3755 718
rect 3811 662 3879 718
rect 3935 662 3945 718
rect 3621 652 3945 662
rect 4721 438 5045 448
rect 4721 382 4731 438
rect 4787 382 4855 438
rect 4911 382 4979 438
rect 5035 382 5045 438
rect 4721 314 5045 382
rect 4721 258 4731 314
rect 4787 258 4855 314
rect 4911 258 4979 314
rect 5035 258 5045 314
rect 4721 190 5045 258
rect 4721 134 4731 190
rect 4787 134 4855 190
rect 4911 134 4979 190
rect 5035 134 5045 190
rect 4721 66 5045 134
rect 4721 10 4731 66
rect 4787 10 4855 66
rect 4911 10 4979 66
rect 5035 10 5045 66
rect 4721 -58 5045 10
rect 4721 -114 4731 -58
rect 4787 -114 4855 -58
rect 4911 -114 4979 -58
rect 5035 -114 5045 -58
rect 4721 -182 5045 -114
rect 4721 -238 4731 -182
rect 4787 -238 4855 -182
rect 4911 -238 4979 -182
rect 5035 -238 5045 -182
rect 4721 -248 5045 -238
<< via2 >>
rect 3631 1336 3687 1338
rect 3631 1284 3633 1336
rect 3633 1284 3685 1336
rect 3685 1284 3687 1336
rect 3631 1282 3687 1284
rect 3755 1336 3811 1338
rect 3755 1284 3757 1336
rect 3757 1284 3809 1336
rect 3809 1284 3811 1336
rect 3755 1282 3811 1284
rect 3879 1336 3935 1338
rect 3879 1284 3881 1336
rect 3881 1284 3933 1336
rect 3933 1284 3935 1336
rect 3879 1282 3935 1284
rect 3631 1212 3687 1214
rect 3631 1160 3633 1212
rect 3633 1160 3685 1212
rect 3685 1160 3687 1212
rect 3631 1158 3687 1160
rect 3755 1212 3811 1214
rect 3755 1160 3757 1212
rect 3757 1160 3809 1212
rect 3809 1160 3811 1212
rect 3755 1158 3811 1160
rect 3879 1212 3935 1214
rect 3879 1160 3881 1212
rect 3881 1160 3933 1212
rect 3933 1160 3935 1212
rect 3879 1158 3935 1160
rect 3631 1088 3687 1090
rect 3631 1036 3633 1088
rect 3633 1036 3685 1088
rect 3685 1036 3687 1088
rect 3631 1034 3687 1036
rect 3755 1088 3811 1090
rect 3755 1036 3757 1088
rect 3757 1036 3809 1088
rect 3809 1036 3811 1088
rect 3755 1034 3811 1036
rect 3879 1088 3935 1090
rect 3879 1036 3881 1088
rect 3881 1036 3933 1088
rect 3933 1036 3935 1088
rect 3879 1034 3935 1036
rect 3631 964 3687 966
rect 3631 912 3633 964
rect 3633 912 3685 964
rect 3685 912 3687 964
rect 3631 910 3687 912
rect 3755 964 3811 966
rect 3755 912 3757 964
rect 3757 912 3809 964
rect 3809 912 3811 964
rect 3755 910 3811 912
rect 3879 964 3935 966
rect 3879 912 3881 964
rect 3881 912 3933 964
rect 3933 912 3935 964
rect 3879 910 3935 912
rect 3631 840 3687 842
rect 3631 788 3633 840
rect 3633 788 3685 840
rect 3685 788 3687 840
rect 3631 786 3687 788
rect 3755 840 3811 842
rect 3755 788 3757 840
rect 3757 788 3809 840
rect 3809 788 3811 840
rect 3755 786 3811 788
rect 3879 840 3935 842
rect 3879 788 3881 840
rect 3881 788 3933 840
rect 3933 788 3935 840
rect 3879 786 3935 788
rect 3631 716 3687 718
rect 3631 664 3633 716
rect 3633 664 3685 716
rect 3685 664 3687 716
rect 3631 662 3687 664
rect 3755 716 3811 718
rect 3755 664 3757 716
rect 3757 664 3809 716
rect 3809 664 3811 716
rect 3755 662 3811 664
rect 3879 716 3935 718
rect 3879 664 3881 716
rect 3881 664 3933 716
rect 3933 664 3935 716
rect 3879 662 3935 664
rect 4731 436 4787 438
rect 4731 384 4733 436
rect 4733 384 4785 436
rect 4785 384 4787 436
rect 4731 382 4787 384
rect 4855 436 4911 438
rect 4855 384 4857 436
rect 4857 384 4909 436
rect 4909 384 4911 436
rect 4855 382 4911 384
rect 4979 436 5035 438
rect 4979 384 4981 436
rect 4981 384 5033 436
rect 5033 384 5035 436
rect 4979 382 5035 384
rect 4731 312 4787 314
rect 4731 260 4733 312
rect 4733 260 4785 312
rect 4785 260 4787 312
rect 4731 258 4787 260
rect 4855 312 4911 314
rect 4855 260 4857 312
rect 4857 260 4909 312
rect 4909 260 4911 312
rect 4855 258 4911 260
rect 4979 312 5035 314
rect 4979 260 4981 312
rect 4981 260 5033 312
rect 5033 260 5035 312
rect 4979 258 5035 260
rect 4731 188 4787 190
rect 4731 136 4733 188
rect 4733 136 4785 188
rect 4785 136 4787 188
rect 4731 134 4787 136
rect 4855 188 4911 190
rect 4855 136 4857 188
rect 4857 136 4909 188
rect 4909 136 4911 188
rect 4855 134 4911 136
rect 4979 188 5035 190
rect 4979 136 4981 188
rect 4981 136 5033 188
rect 5033 136 5035 188
rect 4979 134 5035 136
rect 4731 64 4787 66
rect 4731 12 4733 64
rect 4733 12 4785 64
rect 4785 12 4787 64
rect 4731 10 4787 12
rect 4855 64 4911 66
rect 4855 12 4857 64
rect 4857 12 4909 64
rect 4909 12 4911 64
rect 4855 10 4911 12
rect 4979 64 5035 66
rect 4979 12 4981 64
rect 4981 12 5033 64
rect 5033 12 5035 64
rect 4979 10 5035 12
rect 4731 -60 4787 -58
rect 4731 -112 4733 -60
rect 4733 -112 4785 -60
rect 4785 -112 4787 -60
rect 4731 -114 4787 -112
rect 4855 -60 4911 -58
rect 4855 -112 4857 -60
rect 4857 -112 4909 -60
rect 4909 -112 4911 -60
rect 4855 -114 4911 -112
rect 4979 -60 5035 -58
rect 4979 -112 4981 -60
rect 4981 -112 5033 -60
rect 5033 -112 5035 -60
rect 4979 -114 5035 -112
rect 4731 -184 4787 -182
rect 4731 -236 4733 -184
rect 4733 -236 4785 -184
rect 4785 -236 4787 -184
rect 4731 -238 4787 -236
rect 4855 -184 4911 -182
rect 4855 -236 4857 -184
rect 4857 -236 4909 -184
rect 4909 -236 4911 -184
rect 4855 -238 4911 -236
rect 4979 -184 5035 -182
rect 4979 -236 4981 -184
rect 4981 -236 5033 -184
rect 5033 -236 5035 -184
rect 4979 -238 5035 -236
<< metal3 >>
rect 3339 1338 4353 1350
rect 3339 1282 3631 1338
rect 3687 1282 3755 1338
rect 3811 1282 3879 1338
rect 3935 1282 4353 1338
rect 3339 1214 4353 1282
rect 3339 1158 3631 1214
rect 3687 1158 3755 1214
rect 3811 1158 3879 1214
rect 3935 1158 4353 1214
rect 3339 1150 4353 1158
rect 3339 1090 30290 1150
rect 3339 1034 3631 1090
rect 3687 1034 3755 1090
rect 3811 1034 3879 1090
rect 3935 1034 30290 1090
rect 3339 966 30290 1034
rect 3339 910 3631 966
rect 3687 910 3755 966
rect 3811 910 3879 966
rect 3935 910 30290 966
rect 3339 850 30290 910
rect 3339 842 4353 850
rect 3339 786 3631 842
rect 3687 786 3755 842
rect 3811 786 3879 842
rect 3935 786 4353 842
rect 3339 718 4353 786
rect 3339 662 3631 718
rect 3687 662 3755 718
rect 3811 662 3879 718
rect 3935 662 4353 718
rect 3339 650 4353 662
rect 3339 438 5045 450
rect 3339 382 4731 438
rect 4787 382 4855 438
rect 4911 382 4979 438
rect 5035 382 5045 438
rect 3339 314 5045 382
rect 3339 258 4731 314
rect 4787 258 4855 314
rect 4911 258 4979 314
rect 5035 258 5045 314
rect 3339 190 5045 258
rect 3339 134 4731 190
rect 4787 134 4855 190
rect 4911 134 4979 190
rect 5035 134 5045 190
rect 3339 66 5045 134
rect 3339 10 4731 66
rect 4787 10 4855 66
rect 4911 10 4979 66
rect 5035 10 5045 66
rect 3339 -58 5045 10
rect 3339 -114 4731 -58
rect 4787 -114 4855 -58
rect 4911 -114 4979 -58
rect 5035 -114 5045 -58
rect 3339 -182 5045 -114
rect 3339 -238 4731 -182
rect 4787 -238 4855 -182
rect 4911 -238 4979 -182
rect 5035 -238 5045 -182
rect 3339 -250 5045 -238
use M2_M14310589983284_64x8m81  M2_M14310589983284_64x8m81_0
timestamp 1698431365
transform 1 0 3783 0 1 1000
box 0 0 1 1
use M2_M14310589983284_64x8m81  M2_M14310589983284_64x8m81_1
timestamp 1698431365
transform 1 0 4883 0 1 100
box 0 0 1 1
use M3_M24310589983287_64x8m81  M3_M24310589983287_64x8m81_0
timestamp 1698431365
transform 1 0 4883 0 1 100
box 0 0 1 1
use M3_M24310589983287_64x8m81  M3_M24310589983287_64x8m81_1
timestamp 1698431365
transform 1 0 3783 0 1 1000
box 0 0 1 1
<< properties >>
string GDS_END 1624584
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 1624164
string path 25.225 0.500 16.695 0.500 
<< end >>
