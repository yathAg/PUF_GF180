magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< nwell >>
rect 85 29129 22775 29790
rect 85 29053 23905 29129
rect 1342 27025 23905 29053
rect 1342 25454 23709 27025
rect 1342 23867 23707 25454
rect 1216 17407 22310 19961
rect 22338 18379 23707 19961
rect 22338 17923 23923 18379
rect 22338 17407 23905 17923
rect 22338 17406 22926 17407
rect 22827 14326 23842 15917
rect 22992 9181 23846 10665
rect 22880 8391 23846 9181
rect 22992 8114 23846 8391
rect 22861 7037 23846 7493
<< pwell >>
rect 239 39263 23775 39295
rect 239 30119 23775 30151
<< mvnmos >>
rect 23332 22316 23452 23678
rect 23332 20312 23452 21674
rect 23292 17142 23412 17256
rect 23516 17142 23636 17256
rect 23243 13889 23363 14165
rect 23467 13889 23587 14165
rect 23247 10804 23367 12504
rect 23471 10804 23591 12504
<< mvpmos >>
rect 361 29194 834 29649
rect 980 29194 1453 29649
rect 1599 29194 2072 29649
rect 2218 29194 2691 29649
rect 2837 29194 3310 29649
rect 3456 29194 3929 29649
rect 4075 29194 4548 29649
rect 4694 29194 5167 29649
rect 5313 29194 5786 29649
rect 5932 29194 6405 29649
rect 6551 29194 7024 29649
rect 7170 29194 7643 29649
rect 7789 29194 8262 29649
rect 8408 29194 8881 29649
rect 9027 29194 9500 29649
rect 9646 29194 10119 29649
rect 10265 29194 10738 29649
rect 10884 29194 11357 29649
rect 11503 29194 11976 29649
rect 12122 29194 12595 29649
rect 12741 29194 13214 29649
rect 13360 29194 13833 29649
rect 13979 29194 14452 29649
rect 14598 29194 15071 29649
rect 15217 29194 15690 29649
rect 15836 29194 16309 29649
rect 16455 29194 16928 29649
rect 17074 29194 17547 29649
rect 17693 29194 18166 29649
rect 18312 29194 18785 29649
rect 18931 29194 19404 29649
rect 19550 29194 20023 29649
rect 20169 29194 20642 29649
rect 20788 29194 21261 29649
rect 21407 29194 21880 29649
rect 22026 29194 22499 29649
rect 23220 27950 23340 28632
rect 23444 27950 23564 28632
rect 23220 27175 23340 27857
rect 23444 27175 23564 27857
rect 23334 25594 23454 26956
rect 23332 24007 23452 25369
rect 23332 18457 23452 19819
rect 23263 17547 23383 17844
rect 23515 17547 23635 17844
rect 23243 14469 23363 15171
rect 23467 14469 23587 15171
rect 23247 8395 23367 10523
rect 23471 8395 23591 10523
<< mvndiff >>
rect 23244 23665 23332 23678
rect 23244 23619 23257 23665
rect 23303 23619 23332 23665
rect 23244 23557 23332 23619
rect 23244 23511 23257 23557
rect 23303 23511 23332 23557
rect 23244 23449 23332 23511
rect 23244 23403 23257 23449
rect 23303 23403 23332 23449
rect 23244 23341 23332 23403
rect 23244 23295 23257 23341
rect 23303 23295 23332 23341
rect 23244 23233 23332 23295
rect 23244 23187 23257 23233
rect 23303 23187 23332 23233
rect 23244 23125 23332 23187
rect 23244 23079 23257 23125
rect 23303 23079 23332 23125
rect 23244 23017 23332 23079
rect 23244 22971 23257 23017
rect 23303 22971 23332 23017
rect 23244 22910 23332 22971
rect 23244 22864 23257 22910
rect 23303 22864 23332 22910
rect 23244 22803 23332 22864
rect 23244 22757 23257 22803
rect 23303 22757 23332 22803
rect 23244 22696 23332 22757
rect 23244 22650 23257 22696
rect 23303 22650 23332 22696
rect 23244 22589 23332 22650
rect 23244 22543 23257 22589
rect 23303 22543 23332 22589
rect 23244 22482 23332 22543
rect 23244 22436 23257 22482
rect 23303 22436 23332 22482
rect 23244 22375 23332 22436
rect 23244 22329 23257 22375
rect 23303 22329 23332 22375
rect 23244 22316 23332 22329
rect 23452 23665 23540 23678
rect 23452 23619 23481 23665
rect 23527 23619 23540 23665
rect 23452 23557 23540 23619
rect 23452 23511 23481 23557
rect 23527 23511 23540 23557
rect 23452 23449 23540 23511
rect 23452 23403 23481 23449
rect 23527 23403 23540 23449
rect 23452 23341 23540 23403
rect 23452 23295 23481 23341
rect 23527 23295 23540 23341
rect 23452 23233 23540 23295
rect 23452 23187 23481 23233
rect 23527 23187 23540 23233
rect 23452 23125 23540 23187
rect 23452 23079 23481 23125
rect 23527 23079 23540 23125
rect 23452 23017 23540 23079
rect 23452 22971 23481 23017
rect 23527 22971 23540 23017
rect 23452 22910 23540 22971
rect 23452 22864 23481 22910
rect 23527 22864 23540 22910
rect 23452 22803 23540 22864
rect 23452 22757 23481 22803
rect 23527 22757 23540 22803
rect 23452 22696 23540 22757
rect 23452 22650 23481 22696
rect 23527 22650 23540 22696
rect 23452 22589 23540 22650
rect 23452 22543 23481 22589
rect 23527 22543 23540 22589
rect 23452 22482 23540 22543
rect 23452 22436 23481 22482
rect 23527 22436 23540 22482
rect 23452 22375 23540 22436
rect 23452 22329 23481 22375
rect 23527 22329 23540 22375
rect 23452 22316 23540 22329
rect 23244 21661 23332 21674
rect 23244 21615 23257 21661
rect 23303 21615 23332 21661
rect 23244 21553 23332 21615
rect 23244 21507 23257 21553
rect 23303 21507 23332 21553
rect 23244 21445 23332 21507
rect 23244 21399 23257 21445
rect 23303 21399 23332 21445
rect 23244 21337 23332 21399
rect 23244 21291 23257 21337
rect 23303 21291 23332 21337
rect 23244 21229 23332 21291
rect 23244 21183 23257 21229
rect 23303 21183 23332 21229
rect 23244 21121 23332 21183
rect 23244 21075 23257 21121
rect 23303 21075 23332 21121
rect 23244 21013 23332 21075
rect 23244 20967 23257 21013
rect 23303 20967 23332 21013
rect 23244 20906 23332 20967
rect 23244 20860 23257 20906
rect 23303 20860 23332 20906
rect 23244 20799 23332 20860
rect 23244 20753 23257 20799
rect 23303 20753 23332 20799
rect 23244 20692 23332 20753
rect 23244 20646 23257 20692
rect 23303 20646 23332 20692
rect 23244 20585 23332 20646
rect 23244 20539 23257 20585
rect 23303 20539 23332 20585
rect 23244 20478 23332 20539
rect 23244 20432 23257 20478
rect 23303 20432 23332 20478
rect 23244 20371 23332 20432
rect 23244 20325 23257 20371
rect 23303 20325 23332 20371
rect 23244 20312 23332 20325
rect 23452 21661 23540 21674
rect 23452 21615 23481 21661
rect 23527 21615 23540 21661
rect 23452 21553 23540 21615
rect 23452 21507 23481 21553
rect 23527 21507 23540 21553
rect 23452 21445 23540 21507
rect 23452 21399 23481 21445
rect 23527 21399 23540 21445
rect 23452 21337 23540 21399
rect 23452 21291 23481 21337
rect 23527 21291 23540 21337
rect 23452 21229 23540 21291
rect 23452 21183 23481 21229
rect 23527 21183 23540 21229
rect 23452 21121 23540 21183
rect 23452 21075 23481 21121
rect 23527 21075 23540 21121
rect 23452 21013 23540 21075
rect 23452 20967 23481 21013
rect 23527 20967 23540 21013
rect 23452 20906 23540 20967
rect 23452 20860 23481 20906
rect 23527 20860 23540 20906
rect 23452 20799 23540 20860
rect 23452 20753 23481 20799
rect 23527 20753 23540 20799
rect 23452 20692 23540 20753
rect 23452 20646 23481 20692
rect 23527 20646 23540 20692
rect 23452 20585 23540 20646
rect 23452 20539 23481 20585
rect 23527 20539 23540 20585
rect 23452 20478 23540 20539
rect 23452 20432 23481 20478
rect 23527 20432 23540 20478
rect 23452 20371 23540 20432
rect 23452 20325 23481 20371
rect 23527 20325 23540 20371
rect 23452 20312 23540 20325
rect 23204 17222 23292 17256
rect 23204 17176 23217 17222
rect 23263 17176 23292 17222
rect 23204 17142 23292 17176
rect 23412 17222 23516 17256
rect 23412 17176 23441 17222
rect 23487 17176 23516 17222
rect 23412 17142 23516 17176
rect 23636 17222 23724 17256
rect 23636 17176 23665 17222
rect 23711 17176 23724 17222
rect 23636 17142 23724 17176
rect 23155 14152 23243 14165
rect 23155 13902 23168 14152
rect 23214 13902 23243 14152
rect 23155 13889 23243 13902
rect 23363 14152 23467 14165
rect 23363 13902 23392 14152
rect 23438 13902 23467 14152
rect 23363 13889 23467 13902
rect 23587 14152 23675 14165
rect 23587 13902 23616 14152
rect 23662 13902 23675 14152
rect 23587 13889 23675 13902
rect 23159 12491 23247 12504
rect 23159 10817 23172 12491
rect 23218 10817 23247 12491
rect 23159 10804 23247 10817
rect 23367 12491 23471 12504
rect 23367 10817 23396 12491
rect 23442 10817 23471 12491
rect 23367 10804 23471 10817
rect 23591 12491 23679 12504
rect 23591 10817 23620 12491
rect 23666 10817 23679 12491
rect 23591 10804 23679 10817
<< mvpdiff >>
rect 221 29604 361 29649
rect 221 29558 265 29604
rect 311 29558 361 29604
rect 221 29286 361 29558
rect 221 29240 265 29286
rect 311 29240 361 29286
rect 221 29194 361 29240
rect 834 29604 980 29649
rect 834 29558 884 29604
rect 930 29558 980 29604
rect 834 29286 980 29558
rect 834 29240 884 29286
rect 930 29240 980 29286
rect 834 29194 980 29240
rect 1453 29604 1599 29649
rect 1453 29558 1503 29604
rect 1549 29558 1599 29604
rect 1453 29286 1599 29558
rect 1453 29240 1503 29286
rect 1549 29240 1599 29286
rect 1453 29194 1599 29240
rect 2072 29604 2218 29649
rect 2072 29558 2122 29604
rect 2168 29558 2218 29604
rect 2072 29286 2218 29558
rect 2072 29240 2122 29286
rect 2168 29240 2218 29286
rect 2072 29194 2218 29240
rect 2691 29604 2837 29649
rect 2691 29558 2741 29604
rect 2787 29558 2837 29604
rect 2691 29286 2837 29558
rect 2691 29240 2741 29286
rect 2787 29240 2837 29286
rect 2691 29194 2837 29240
rect 3310 29604 3456 29649
rect 3310 29558 3360 29604
rect 3406 29558 3456 29604
rect 3310 29286 3456 29558
rect 3310 29240 3360 29286
rect 3406 29240 3456 29286
rect 3310 29194 3456 29240
rect 3929 29604 4075 29649
rect 3929 29558 3979 29604
rect 4025 29558 4075 29604
rect 3929 29286 4075 29558
rect 3929 29240 3979 29286
rect 4025 29240 4075 29286
rect 3929 29194 4075 29240
rect 4548 29604 4694 29649
rect 4548 29558 4598 29604
rect 4644 29558 4694 29604
rect 4548 29286 4694 29558
rect 4548 29240 4598 29286
rect 4644 29240 4694 29286
rect 4548 29194 4694 29240
rect 5167 29604 5313 29649
rect 5167 29558 5217 29604
rect 5263 29558 5313 29604
rect 5167 29286 5313 29558
rect 5167 29240 5217 29286
rect 5263 29240 5313 29286
rect 5167 29194 5313 29240
rect 5786 29604 5932 29649
rect 5786 29558 5836 29604
rect 5882 29558 5932 29604
rect 5786 29286 5932 29558
rect 5786 29240 5836 29286
rect 5882 29240 5932 29286
rect 5786 29194 5932 29240
rect 6405 29604 6551 29649
rect 6405 29558 6455 29604
rect 6501 29558 6551 29604
rect 6405 29286 6551 29558
rect 6405 29240 6455 29286
rect 6501 29240 6551 29286
rect 6405 29194 6551 29240
rect 7024 29604 7170 29649
rect 7024 29558 7074 29604
rect 7120 29558 7170 29604
rect 7024 29286 7170 29558
rect 7024 29240 7074 29286
rect 7120 29240 7170 29286
rect 7024 29194 7170 29240
rect 7643 29604 7789 29649
rect 7643 29558 7693 29604
rect 7739 29558 7789 29604
rect 7643 29286 7789 29558
rect 7643 29240 7693 29286
rect 7739 29240 7789 29286
rect 7643 29194 7789 29240
rect 8262 29604 8408 29649
rect 8262 29558 8312 29604
rect 8358 29558 8408 29604
rect 8262 29286 8408 29558
rect 8262 29240 8312 29286
rect 8358 29240 8408 29286
rect 8262 29194 8408 29240
rect 8881 29604 9027 29649
rect 8881 29558 8931 29604
rect 8977 29558 9027 29604
rect 8881 29286 9027 29558
rect 8881 29240 8931 29286
rect 8977 29240 9027 29286
rect 8881 29194 9027 29240
rect 9500 29604 9646 29649
rect 9500 29558 9550 29604
rect 9596 29558 9646 29604
rect 9500 29286 9646 29558
rect 9500 29240 9550 29286
rect 9596 29240 9646 29286
rect 9500 29194 9646 29240
rect 10119 29604 10265 29649
rect 10119 29558 10169 29604
rect 10215 29558 10265 29604
rect 10119 29286 10265 29558
rect 10119 29240 10169 29286
rect 10215 29240 10265 29286
rect 10119 29194 10265 29240
rect 10738 29604 10884 29649
rect 10738 29558 10788 29604
rect 10834 29558 10884 29604
rect 10738 29286 10884 29558
rect 10738 29240 10788 29286
rect 10834 29240 10884 29286
rect 10738 29194 10884 29240
rect 11357 29604 11503 29649
rect 11357 29558 11407 29604
rect 11453 29558 11503 29604
rect 11357 29286 11503 29558
rect 11357 29240 11407 29286
rect 11453 29240 11503 29286
rect 11357 29194 11503 29240
rect 11976 29604 12122 29649
rect 11976 29558 12026 29604
rect 12072 29558 12122 29604
rect 11976 29286 12122 29558
rect 11976 29240 12026 29286
rect 12072 29240 12122 29286
rect 11976 29194 12122 29240
rect 12595 29604 12741 29649
rect 12595 29558 12645 29604
rect 12691 29558 12741 29604
rect 12595 29286 12741 29558
rect 12595 29240 12645 29286
rect 12691 29240 12741 29286
rect 12595 29194 12741 29240
rect 13214 29604 13360 29649
rect 13214 29558 13264 29604
rect 13310 29558 13360 29604
rect 13214 29286 13360 29558
rect 13214 29240 13264 29286
rect 13310 29240 13360 29286
rect 13214 29194 13360 29240
rect 13833 29604 13979 29649
rect 13833 29558 13883 29604
rect 13929 29558 13979 29604
rect 13833 29286 13979 29558
rect 13833 29240 13883 29286
rect 13929 29240 13979 29286
rect 13833 29194 13979 29240
rect 14452 29604 14598 29649
rect 14452 29558 14502 29604
rect 14548 29558 14598 29604
rect 14452 29286 14598 29558
rect 14452 29240 14502 29286
rect 14548 29240 14598 29286
rect 14452 29194 14598 29240
rect 15071 29604 15217 29649
rect 15071 29558 15121 29604
rect 15167 29558 15217 29604
rect 15071 29286 15217 29558
rect 15071 29240 15121 29286
rect 15167 29240 15217 29286
rect 15071 29194 15217 29240
rect 15690 29604 15836 29649
rect 15690 29558 15740 29604
rect 15786 29558 15836 29604
rect 15690 29286 15836 29558
rect 15690 29240 15740 29286
rect 15786 29240 15836 29286
rect 15690 29194 15836 29240
rect 16309 29604 16455 29649
rect 16309 29558 16359 29604
rect 16405 29558 16455 29604
rect 16309 29286 16455 29558
rect 16309 29240 16359 29286
rect 16405 29240 16455 29286
rect 16309 29194 16455 29240
rect 16928 29604 17074 29649
rect 16928 29558 16978 29604
rect 17024 29558 17074 29604
rect 16928 29286 17074 29558
rect 16928 29240 16978 29286
rect 17024 29240 17074 29286
rect 16928 29194 17074 29240
rect 17547 29604 17693 29649
rect 17547 29558 17597 29604
rect 17643 29558 17693 29604
rect 17547 29286 17693 29558
rect 17547 29240 17597 29286
rect 17643 29240 17693 29286
rect 17547 29194 17693 29240
rect 18166 29604 18312 29649
rect 18166 29558 18216 29604
rect 18262 29558 18312 29604
rect 18166 29286 18312 29558
rect 18166 29240 18216 29286
rect 18262 29240 18312 29286
rect 18166 29194 18312 29240
rect 18785 29604 18931 29649
rect 18785 29558 18835 29604
rect 18881 29558 18931 29604
rect 18785 29286 18931 29558
rect 18785 29240 18835 29286
rect 18881 29240 18931 29286
rect 18785 29194 18931 29240
rect 19404 29604 19550 29649
rect 19404 29558 19454 29604
rect 19500 29558 19550 29604
rect 19404 29286 19550 29558
rect 19404 29240 19454 29286
rect 19500 29240 19550 29286
rect 19404 29194 19550 29240
rect 20023 29604 20169 29649
rect 20023 29558 20073 29604
rect 20119 29558 20169 29604
rect 20023 29286 20169 29558
rect 20023 29240 20073 29286
rect 20119 29240 20169 29286
rect 20023 29194 20169 29240
rect 20642 29604 20788 29649
rect 20642 29558 20692 29604
rect 20738 29558 20788 29604
rect 20642 29286 20788 29558
rect 20642 29240 20692 29286
rect 20738 29240 20788 29286
rect 20642 29194 20788 29240
rect 21261 29604 21407 29649
rect 21261 29558 21311 29604
rect 21357 29558 21407 29604
rect 21261 29286 21407 29558
rect 21261 29240 21311 29286
rect 21357 29240 21407 29286
rect 21261 29194 21407 29240
rect 21880 29604 22026 29649
rect 21880 29558 21930 29604
rect 21976 29558 22026 29604
rect 21880 29286 22026 29558
rect 21880 29240 21930 29286
rect 21976 29240 22026 29286
rect 21880 29194 22026 29240
rect 22499 29604 22639 29649
rect 22499 29558 22549 29604
rect 22595 29558 22639 29604
rect 22499 29286 22639 29558
rect 22499 29240 22549 29286
rect 22595 29240 22639 29286
rect 22499 29194 22639 29240
rect 23052 28587 23220 28632
rect 23052 28541 23143 28587
rect 23189 28541 23220 28587
rect 23052 28405 23220 28541
rect 23052 28359 23143 28405
rect 23189 28359 23220 28405
rect 23052 28224 23220 28359
rect 23052 28178 23143 28224
rect 23189 28178 23220 28224
rect 23052 28042 23220 28178
rect 23052 27996 23143 28042
rect 23189 27996 23220 28042
rect 23052 27950 23220 27996
rect 23340 28587 23444 28632
rect 23340 28541 23369 28587
rect 23415 28541 23444 28587
rect 23340 28405 23444 28541
rect 23340 28359 23369 28405
rect 23415 28359 23444 28405
rect 23340 28224 23444 28359
rect 23340 28178 23369 28224
rect 23415 28178 23444 28224
rect 23340 28042 23444 28178
rect 23340 27996 23369 28042
rect 23415 27996 23444 28042
rect 23340 27950 23444 27996
rect 23564 28587 23769 28632
rect 23564 28541 23679 28587
rect 23725 28541 23769 28587
rect 23564 28405 23769 28541
rect 23564 28359 23679 28405
rect 23725 28359 23769 28405
rect 23564 28224 23769 28359
rect 23564 28178 23679 28224
rect 23725 28178 23769 28224
rect 23564 28042 23769 28178
rect 23564 27996 23679 28042
rect 23725 27996 23769 28042
rect 23564 27950 23769 27996
rect 23052 27811 23220 27857
rect 23052 27765 23143 27811
rect 23189 27765 23220 27811
rect 23052 27630 23220 27765
rect 23052 27584 23143 27630
rect 23189 27584 23220 27630
rect 23052 27449 23220 27584
rect 23052 27403 23143 27449
rect 23189 27403 23220 27449
rect 23052 27267 23220 27403
rect 23052 27221 23143 27267
rect 23189 27221 23220 27267
rect 23052 27175 23220 27221
rect 23340 27811 23444 27857
rect 23340 27765 23369 27811
rect 23415 27765 23444 27811
rect 23340 27630 23444 27765
rect 23340 27584 23369 27630
rect 23415 27584 23444 27630
rect 23340 27449 23444 27584
rect 23340 27403 23369 27449
rect 23415 27403 23444 27449
rect 23340 27267 23444 27403
rect 23340 27221 23369 27267
rect 23415 27221 23444 27267
rect 23340 27175 23444 27221
rect 23564 27811 23769 27857
rect 23564 27765 23679 27811
rect 23725 27765 23769 27811
rect 23564 27630 23769 27765
rect 23564 27584 23679 27630
rect 23725 27584 23769 27630
rect 23564 27449 23769 27584
rect 23564 27403 23679 27449
rect 23725 27403 23769 27449
rect 23564 27267 23769 27403
rect 23564 27221 23679 27267
rect 23725 27221 23769 27267
rect 23564 27175 23769 27221
rect 23246 26943 23334 26956
rect 23246 26897 23259 26943
rect 23305 26897 23334 26943
rect 23246 26835 23334 26897
rect 23246 26789 23259 26835
rect 23305 26789 23334 26835
rect 23246 26727 23334 26789
rect 23246 26681 23259 26727
rect 23305 26681 23334 26727
rect 23246 26619 23334 26681
rect 23246 26573 23259 26619
rect 23305 26573 23334 26619
rect 23246 26511 23334 26573
rect 23246 26465 23259 26511
rect 23305 26465 23334 26511
rect 23246 26403 23334 26465
rect 23246 26357 23259 26403
rect 23305 26357 23334 26403
rect 23246 26295 23334 26357
rect 23246 26249 23259 26295
rect 23305 26249 23334 26295
rect 23246 26188 23334 26249
rect 23246 26142 23259 26188
rect 23305 26142 23334 26188
rect 23246 26081 23334 26142
rect 23246 26035 23259 26081
rect 23305 26035 23334 26081
rect 23246 25974 23334 26035
rect 23246 25928 23259 25974
rect 23305 25928 23334 25974
rect 23246 25867 23334 25928
rect 23246 25821 23259 25867
rect 23305 25821 23334 25867
rect 23246 25760 23334 25821
rect 23246 25714 23259 25760
rect 23305 25714 23334 25760
rect 23246 25653 23334 25714
rect 23246 25607 23259 25653
rect 23305 25607 23334 25653
rect 23246 25594 23334 25607
rect 23454 26943 23542 26956
rect 23454 26897 23483 26943
rect 23529 26897 23542 26943
rect 23454 26835 23542 26897
rect 23454 26789 23483 26835
rect 23529 26789 23542 26835
rect 23454 26727 23542 26789
rect 23454 26681 23483 26727
rect 23529 26681 23542 26727
rect 23454 26619 23542 26681
rect 23454 26573 23483 26619
rect 23529 26573 23542 26619
rect 23454 26511 23542 26573
rect 23454 26465 23483 26511
rect 23529 26465 23542 26511
rect 23454 26403 23542 26465
rect 23454 26357 23483 26403
rect 23529 26357 23542 26403
rect 23454 26295 23542 26357
rect 23454 26249 23483 26295
rect 23529 26249 23542 26295
rect 23454 26188 23542 26249
rect 23454 26142 23483 26188
rect 23529 26142 23542 26188
rect 23454 26081 23542 26142
rect 23454 26035 23483 26081
rect 23529 26035 23542 26081
rect 23454 25974 23542 26035
rect 23454 25928 23483 25974
rect 23529 25928 23542 25974
rect 23454 25867 23542 25928
rect 23454 25821 23483 25867
rect 23529 25821 23542 25867
rect 23454 25760 23542 25821
rect 23454 25714 23483 25760
rect 23529 25714 23542 25760
rect 23454 25653 23542 25714
rect 23454 25607 23483 25653
rect 23529 25607 23542 25653
rect 23454 25594 23542 25607
rect 23244 25356 23332 25369
rect 23244 25310 23257 25356
rect 23303 25310 23332 25356
rect 23244 25248 23332 25310
rect 23244 25202 23257 25248
rect 23303 25202 23332 25248
rect 23244 25140 23332 25202
rect 23244 25094 23257 25140
rect 23303 25094 23332 25140
rect 23244 25032 23332 25094
rect 23244 24986 23257 25032
rect 23303 24986 23332 25032
rect 23244 24924 23332 24986
rect 23244 24878 23257 24924
rect 23303 24878 23332 24924
rect 23244 24816 23332 24878
rect 23244 24770 23257 24816
rect 23303 24770 23332 24816
rect 23244 24708 23332 24770
rect 23244 24662 23257 24708
rect 23303 24662 23332 24708
rect 23244 24601 23332 24662
rect 23244 24555 23257 24601
rect 23303 24555 23332 24601
rect 23244 24494 23332 24555
rect 23244 24448 23257 24494
rect 23303 24448 23332 24494
rect 23244 24387 23332 24448
rect 23244 24341 23257 24387
rect 23303 24341 23332 24387
rect 23244 24280 23332 24341
rect 23244 24234 23257 24280
rect 23303 24234 23332 24280
rect 23244 24173 23332 24234
rect 23244 24127 23257 24173
rect 23303 24127 23332 24173
rect 23244 24066 23332 24127
rect 23244 24020 23257 24066
rect 23303 24020 23332 24066
rect 23244 24007 23332 24020
rect 23452 25356 23540 25369
rect 23452 25310 23481 25356
rect 23527 25310 23540 25356
rect 23452 25248 23540 25310
rect 23452 25202 23481 25248
rect 23527 25202 23540 25248
rect 23452 25140 23540 25202
rect 23452 25094 23481 25140
rect 23527 25094 23540 25140
rect 23452 25032 23540 25094
rect 23452 24986 23481 25032
rect 23527 24986 23540 25032
rect 23452 24924 23540 24986
rect 23452 24878 23481 24924
rect 23527 24878 23540 24924
rect 23452 24816 23540 24878
rect 23452 24770 23481 24816
rect 23527 24770 23540 24816
rect 23452 24708 23540 24770
rect 23452 24662 23481 24708
rect 23527 24662 23540 24708
rect 23452 24601 23540 24662
rect 23452 24555 23481 24601
rect 23527 24555 23540 24601
rect 23452 24494 23540 24555
rect 23452 24448 23481 24494
rect 23527 24448 23540 24494
rect 23452 24387 23540 24448
rect 23452 24341 23481 24387
rect 23527 24341 23540 24387
rect 23452 24280 23540 24341
rect 23452 24234 23481 24280
rect 23527 24234 23540 24280
rect 23452 24173 23540 24234
rect 23452 24127 23481 24173
rect 23527 24127 23540 24173
rect 23452 24066 23540 24127
rect 23452 24020 23481 24066
rect 23527 24020 23540 24066
rect 23452 24007 23540 24020
rect 23244 19806 23332 19819
rect 23244 19760 23257 19806
rect 23303 19760 23332 19806
rect 23244 19698 23332 19760
rect 23244 19652 23257 19698
rect 23303 19652 23332 19698
rect 23244 19590 23332 19652
rect 23244 19544 23257 19590
rect 23303 19544 23332 19590
rect 23244 19482 23332 19544
rect 23244 19436 23257 19482
rect 23303 19436 23332 19482
rect 23244 19374 23332 19436
rect 23244 19328 23257 19374
rect 23303 19328 23332 19374
rect 23244 19266 23332 19328
rect 23244 19220 23257 19266
rect 23303 19220 23332 19266
rect 23244 19158 23332 19220
rect 23244 19112 23257 19158
rect 23303 19112 23332 19158
rect 23244 19051 23332 19112
rect 23244 19005 23257 19051
rect 23303 19005 23332 19051
rect 23244 18944 23332 19005
rect 23244 18898 23257 18944
rect 23303 18898 23332 18944
rect 23244 18837 23332 18898
rect 23244 18791 23257 18837
rect 23303 18791 23332 18837
rect 23244 18730 23332 18791
rect 23244 18684 23257 18730
rect 23303 18684 23332 18730
rect 23244 18623 23332 18684
rect 23244 18577 23257 18623
rect 23303 18577 23332 18623
rect 23244 18516 23332 18577
rect 23244 18470 23257 18516
rect 23303 18470 23332 18516
rect 23244 18457 23332 18470
rect 23452 19806 23540 19819
rect 23452 19760 23481 19806
rect 23527 19760 23540 19806
rect 23452 19698 23540 19760
rect 23452 19652 23481 19698
rect 23527 19652 23540 19698
rect 23452 19590 23540 19652
rect 23452 19544 23481 19590
rect 23527 19544 23540 19590
rect 23452 19482 23540 19544
rect 23452 19436 23481 19482
rect 23527 19436 23540 19482
rect 23452 19374 23540 19436
rect 23452 19328 23481 19374
rect 23527 19328 23540 19374
rect 23452 19266 23540 19328
rect 23452 19220 23481 19266
rect 23527 19220 23540 19266
rect 23452 19158 23540 19220
rect 23452 19112 23481 19158
rect 23527 19112 23540 19158
rect 23452 19051 23540 19112
rect 23452 19005 23481 19051
rect 23527 19005 23540 19051
rect 23452 18944 23540 19005
rect 23452 18898 23481 18944
rect 23527 18898 23540 18944
rect 23452 18837 23540 18898
rect 23452 18791 23481 18837
rect 23527 18791 23540 18837
rect 23452 18730 23540 18791
rect 23452 18684 23481 18730
rect 23527 18684 23540 18730
rect 23452 18623 23540 18684
rect 23452 18577 23481 18623
rect 23527 18577 23540 18623
rect 23452 18516 23540 18577
rect 23452 18470 23481 18516
rect 23527 18470 23540 18516
rect 23452 18457 23540 18470
rect 23082 17719 23263 17844
rect 23082 17673 23176 17719
rect 23222 17673 23263 17719
rect 23082 17547 23263 17673
rect 23383 17719 23515 17844
rect 23383 17673 23426 17719
rect 23472 17673 23515 17719
rect 23383 17547 23515 17673
rect 23635 17719 23769 17844
rect 23635 17673 23679 17719
rect 23725 17673 23769 17719
rect 23635 17547 23769 17673
rect 23155 15158 23243 15171
rect 23155 15112 23168 15158
rect 23214 15112 23243 15158
rect 23155 15053 23243 15112
rect 23155 15007 23168 15053
rect 23214 15007 23243 15053
rect 23155 14948 23243 15007
rect 23155 14902 23168 14948
rect 23214 14902 23243 14948
rect 23155 14843 23243 14902
rect 23155 14797 23168 14843
rect 23214 14797 23243 14843
rect 23155 14738 23243 14797
rect 23155 14692 23168 14738
rect 23214 14692 23243 14738
rect 23155 14633 23243 14692
rect 23155 14587 23168 14633
rect 23214 14587 23243 14633
rect 23155 14528 23243 14587
rect 23155 14482 23168 14528
rect 23214 14482 23243 14528
rect 23155 14469 23243 14482
rect 23363 15158 23467 15171
rect 23363 15112 23392 15158
rect 23438 15112 23467 15158
rect 23363 15053 23467 15112
rect 23363 15007 23392 15053
rect 23438 15007 23467 15053
rect 23363 14948 23467 15007
rect 23363 14902 23392 14948
rect 23438 14902 23467 14948
rect 23363 14843 23467 14902
rect 23363 14797 23392 14843
rect 23438 14797 23467 14843
rect 23363 14738 23467 14797
rect 23363 14692 23392 14738
rect 23438 14692 23467 14738
rect 23363 14633 23467 14692
rect 23363 14587 23392 14633
rect 23438 14587 23467 14633
rect 23363 14528 23467 14587
rect 23363 14482 23392 14528
rect 23438 14482 23467 14528
rect 23363 14469 23467 14482
rect 23587 15158 23675 15171
rect 23587 15112 23616 15158
rect 23662 15112 23675 15158
rect 23587 15053 23675 15112
rect 23587 15007 23616 15053
rect 23662 15007 23675 15053
rect 23587 14948 23675 15007
rect 23587 14902 23616 14948
rect 23662 14902 23675 14948
rect 23587 14843 23675 14902
rect 23587 14797 23616 14843
rect 23662 14797 23675 14843
rect 23587 14738 23675 14797
rect 23587 14692 23616 14738
rect 23662 14692 23675 14738
rect 23587 14633 23675 14692
rect 23587 14587 23616 14633
rect 23662 14587 23675 14633
rect 23587 14528 23675 14587
rect 23587 14482 23616 14528
rect 23662 14482 23675 14528
rect 23587 14469 23675 14482
rect 23159 10510 23247 10523
rect 23159 10464 23172 10510
rect 23218 10464 23247 10510
rect 23159 10407 23247 10464
rect 23159 10361 23172 10407
rect 23218 10361 23247 10407
rect 23159 10304 23247 10361
rect 23159 10258 23172 10304
rect 23218 10258 23247 10304
rect 23159 10201 23247 10258
rect 23159 10155 23172 10201
rect 23218 10155 23247 10201
rect 23159 10098 23247 10155
rect 23159 10052 23172 10098
rect 23218 10052 23247 10098
rect 23159 9995 23247 10052
rect 23159 9949 23172 9995
rect 23218 9949 23247 9995
rect 23159 9892 23247 9949
rect 23159 9846 23172 9892
rect 23218 9846 23247 9892
rect 23159 9789 23247 9846
rect 23159 9743 23172 9789
rect 23218 9743 23247 9789
rect 23159 9686 23247 9743
rect 23159 9640 23172 9686
rect 23218 9640 23247 9686
rect 23159 9583 23247 9640
rect 23159 9537 23172 9583
rect 23218 9537 23247 9583
rect 23159 9480 23247 9537
rect 23159 9434 23172 9480
rect 23218 9434 23247 9480
rect 23159 9377 23247 9434
rect 23159 9331 23172 9377
rect 23218 9331 23247 9377
rect 23159 9274 23247 9331
rect 23159 9228 23172 9274
rect 23218 9228 23247 9274
rect 23159 9171 23247 9228
rect 23159 9125 23172 9171
rect 23218 9125 23247 9171
rect 23159 9068 23247 9125
rect 23159 9022 23172 9068
rect 23218 9022 23247 9068
rect 23159 8965 23247 9022
rect 23159 8919 23172 8965
rect 23218 8919 23247 8965
rect 23159 8862 23247 8919
rect 23159 8408 23172 8862
rect 23218 8408 23247 8862
rect 23159 8395 23247 8408
rect 23367 10510 23471 10523
rect 23367 10464 23396 10510
rect 23442 10464 23471 10510
rect 23367 10407 23471 10464
rect 23367 10361 23396 10407
rect 23442 10361 23471 10407
rect 23367 10304 23471 10361
rect 23367 10258 23396 10304
rect 23442 10258 23471 10304
rect 23367 10201 23471 10258
rect 23367 10155 23396 10201
rect 23442 10155 23471 10201
rect 23367 10098 23471 10155
rect 23367 10052 23396 10098
rect 23442 10052 23471 10098
rect 23367 9995 23471 10052
rect 23367 9949 23396 9995
rect 23442 9949 23471 9995
rect 23367 9892 23471 9949
rect 23367 9846 23396 9892
rect 23442 9846 23471 9892
rect 23367 9789 23471 9846
rect 23367 9743 23396 9789
rect 23442 9743 23471 9789
rect 23367 9686 23471 9743
rect 23367 9640 23396 9686
rect 23442 9640 23471 9686
rect 23367 9583 23471 9640
rect 23367 9537 23396 9583
rect 23442 9537 23471 9583
rect 23367 9480 23471 9537
rect 23367 9434 23396 9480
rect 23442 9434 23471 9480
rect 23367 9377 23471 9434
rect 23367 9331 23396 9377
rect 23442 9331 23471 9377
rect 23367 9274 23471 9331
rect 23367 9228 23396 9274
rect 23442 9228 23471 9274
rect 23367 9171 23471 9228
rect 23367 9125 23396 9171
rect 23442 9125 23471 9171
rect 23367 9068 23471 9125
rect 23367 9022 23396 9068
rect 23442 9022 23471 9068
rect 23367 8965 23471 9022
rect 23367 8919 23396 8965
rect 23442 8919 23471 8965
rect 23367 8862 23471 8919
rect 23367 8408 23396 8862
rect 23442 8408 23471 8862
rect 23367 8395 23471 8408
rect 23591 10510 23679 10523
rect 23591 10464 23620 10510
rect 23666 10464 23679 10510
rect 23591 10407 23679 10464
rect 23591 10361 23620 10407
rect 23666 10361 23679 10407
rect 23591 10304 23679 10361
rect 23591 10258 23620 10304
rect 23666 10258 23679 10304
rect 23591 10201 23679 10258
rect 23591 10155 23620 10201
rect 23666 10155 23679 10201
rect 23591 10098 23679 10155
rect 23591 10052 23620 10098
rect 23666 10052 23679 10098
rect 23591 9995 23679 10052
rect 23591 9949 23620 9995
rect 23666 9949 23679 9995
rect 23591 9892 23679 9949
rect 23591 9846 23620 9892
rect 23666 9846 23679 9892
rect 23591 9789 23679 9846
rect 23591 9743 23620 9789
rect 23666 9743 23679 9789
rect 23591 9686 23679 9743
rect 23591 9640 23620 9686
rect 23666 9640 23679 9686
rect 23591 9583 23679 9640
rect 23591 9537 23620 9583
rect 23666 9537 23679 9583
rect 23591 9480 23679 9537
rect 23591 9434 23620 9480
rect 23666 9434 23679 9480
rect 23591 9377 23679 9434
rect 23591 9331 23620 9377
rect 23666 9331 23679 9377
rect 23591 9274 23679 9331
rect 23591 9228 23620 9274
rect 23666 9228 23679 9274
rect 23591 9171 23679 9228
rect 23591 9125 23620 9171
rect 23666 9125 23679 9171
rect 23591 9068 23679 9125
rect 23591 9022 23620 9068
rect 23666 9022 23679 9068
rect 23591 8965 23679 9022
rect 23591 8919 23620 8965
rect 23666 8919 23679 8965
rect 23591 8862 23679 8919
rect 23591 8408 23620 8862
rect 23666 8408 23679 8862
rect 23591 8395 23679 8408
<< mvndiffc >>
rect 23257 23619 23303 23665
rect 23257 23511 23303 23557
rect 23257 23403 23303 23449
rect 23257 23295 23303 23341
rect 23257 23187 23303 23233
rect 23257 23079 23303 23125
rect 23257 22971 23303 23017
rect 23257 22864 23303 22910
rect 23257 22757 23303 22803
rect 23257 22650 23303 22696
rect 23257 22543 23303 22589
rect 23257 22436 23303 22482
rect 23257 22329 23303 22375
rect 23481 23619 23527 23665
rect 23481 23511 23527 23557
rect 23481 23403 23527 23449
rect 23481 23295 23527 23341
rect 23481 23187 23527 23233
rect 23481 23079 23527 23125
rect 23481 22971 23527 23017
rect 23481 22864 23527 22910
rect 23481 22757 23527 22803
rect 23481 22650 23527 22696
rect 23481 22543 23527 22589
rect 23481 22436 23527 22482
rect 23481 22329 23527 22375
rect 23257 21615 23303 21661
rect 23257 21507 23303 21553
rect 23257 21399 23303 21445
rect 23257 21291 23303 21337
rect 23257 21183 23303 21229
rect 23257 21075 23303 21121
rect 23257 20967 23303 21013
rect 23257 20860 23303 20906
rect 23257 20753 23303 20799
rect 23257 20646 23303 20692
rect 23257 20539 23303 20585
rect 23257 20432 23303 20478
rect 23257 20325 23303 20371
rect 23481 21615 23527 21661
rect 23481 21507 23527 21553
rect 23481 21399 23527 21445
rect 23481 21291 23527 21337
rect 23481 21183 23527 21229
rect 23481 21075 23527 21121
rect 23481 20967 23527 21013
rect 23481 20860 23527 20906
rect 23481 20753 23527 20799
rect 23481 20646 23527 20692
rect 23481 20539 23527 20585
rect 23481 20432 23527 20478
rect 23481 20325 23527 20371
rect 23217 17176 23263 17222
rect 23441 17176 23487 17222
rect 23665 17176 23711 17222
rect 23168 13902 23214 14152
rect 23392 13902 23438 14152
rect 23616 13902 23662 14152
rect 23172 10817 23218 12491
rect 23396 10817 23442 12491
rect 23620 10817 23666 12491
<< mvpdiffc >>
rect 265 29558 311 29604
rect 265 29240 311 29286
rect 884 29558 930 29604
rect 884 29240 930 29286
rect 1503 29558 1549 29604
rect 1503 29240 1549 29286
rect 2122 29558 2168 29604
rect 2122 29240 2168 29286
rect 2741 29558 2787 29604
rect 2741 29240 2787 29286
rect 3360 29558 3406 29604
rect 3360 29240 3406 29286
rect 3979 29558 4025 29604
rect 3979 29240 4025 29286
rect 4598 29558 4644 29604
rect 4598 29240 4644 29286
rect 5217 29558 5263 29604
rect 5217 29240 5263 29286
rect 5836 29558 5882 29604
rect 5836 29240 5882 29286
rect 6455 29558 6501 29604
rect 6455 29240 6501 29286
rect 7074 29558 7120 29604
rect 7074 29240 7120 29286
rect 7693 29558 7739 29604
rect 7693 29240 7739 29286
rect 8312 29558 8358 29604
rect 8312 29240 8358 29286
rect 8931 29558 8977 29604
rect 8931 29240 8977 29286
rect 9550 29558 9596 29604
rect 9550 29240 9596 29286
rect 10169 29558 10215 29604
rect 10169 29240 10215 29286
rect 10788 29558 10834 29604
rect 10788 29240 10834 29286
rect 11407 29558 11453 29604
rect 11407 29240 11453 29286
rect 12026 29558 12072 29604
rect 12026 29240 12072 29286
rect 12645 29558 12691 29604
rect 12645 29240 12691 29286
rect 13264 29558 13310 29604
rect 13264 29240 13310 29286
rect 13883 29558 13929 29604
rect 13883 29240 13929 29286
rect 14502 29558 14548 29604
rect 14502 29240 14548 29286
rect 15121 29558 15167 29604
rect 15121 29240 15167 29286
rect 15740 29558 15786 29604
rect 15740 29240 15786 29286
rect 16359 29558 16405 29604
rect 16359 29240 16405 29286
rect 16978 29558 17024 29604
rect 16978 29240 17024 29286
rect 17597 29558 17643 29604
rect 17597 29240 17643 29286
rect 18216 29558 18262 29604
rect 18216 29240 18262 29286
rect 18835 29558 18881 29604
rect 18835 29240 18881 29286
rect 19454 29558 19500 29604
rect 19454 29240 19500 29286
rect 20073 29558 20119 29604
rect 20073 29240 20119 29286
rect 20692 29558 20738 29604
rect 20692 29240 20738 29286
rect 21311 29558 21357 29604
rect 21311 29240 21357 29286
rect 21930 29558 21976 29604
rect 21930 29240 21976 29286
rect 22549 29558 22595 29604
rect 22549 29240 22595 29286
rect 23143 28541 23189 28587
rect 23143 28359 23189 28405
rect 23143 28178 23189 28224
rect 23143 27996 23189 28042
rect 23369 28541 23415 28587
rect 23369 28359 23415 28405
rect 23369 28178 23415 28224
rect 23369 27996 23415 28042
rect 23679 28541 23725 28587
rect 23679 28359 23725 28405
rect 23679 28178 23725 28224
rect 23679 27996 23725 28042
rect 23143 27765 23189 27811
rect 23143 27584 23189 27630
rect 23143 27403 23189 27449
rect 23143 27221 23189 27267
rect 23369 27765 23415 27811
rect 23369 27584 23415 27630
rect 23369 27403 23415 27449
rect 23369 27221 23415 27267
rect 23679 27765 23725 27811
rect 23679 27584 23725 27630
rect 23679 27403 23725 27449
rect 23679 27221 23725 27267
rect 23259 26897 23305 26943
rect 23259 26789 23305 26835
rect 23259 26681 23305 26727
rect 23259 26573 23305 26619
rect 23259 26465 23305 26511
rect 23259 26357 23305 26403
rect 23259 26249 23305 26295
rect 23259 26142 23305 26188
rect 23259 26035 23305 26081
rect 23259 25928 23305 25974
rect 23259 25821 23305 25867
rect 23259 25714 23305 25760
rect 23259 25607 23305 25653
rect 23483 26897 23529 26943
rect 23483 26789 23529 26835
rect 23483 26681 23529 26727
rect 23483 26573 23529 26619
rect 23483 26465 23529 26511
rect 23483 26357 23529 26403
rect 23483 26249 23529 26295
rect 23483 26142 23529 26188
rect 23483 26035 23529 26081
rect 23483 25928 23529 25974
rect 23483 25821 23529 25867
rect 23483 25714 23529 25760
rect 23483 25607 23529 25653
rect 23257 25310 23303 25356
rect 23257 25202 23303 25248
rect 23257 25094 23303 25140
rect 23257 24986 23303 25032
rect 23257 24878 23303 24924
rect 23257 24770 23303 24816
rect 23257 24662 23303 24708
rect 23257 24555 23303 24601
rect 23257 24448 23303 24494
rect 23257 24341 23303 24387
rect 23257 24234 23303 24280
rect 23257 24127 23303 24173
rect 23257 24020 23303 24066
rect 23481 25310 23527 25356
rect 23481 25202 23527 25248
rect 23481 25094 23527 25140
rect 23481 24986 23527 25032
rect 23481 24878 23527 24924
rect 23481 24770 23527 24816
rect 23481 24662 23527 24708
rect 23481 24555 23527 24601
rect 23481 24448 23527 24494
rect 23481 24341 23527 24387
rect 23481 24234 23527 24280
rect 23481 24127 23527 24173
rect 23481 24020 23527 24066
rect 23257 19760 23303 19806
rect 23257 19652 23303 19698
rect 23257 19544 23303 19590
rect 23257 19436 23303 19482
rect 23257 19328 23303 19374
rect 23257 19220 23303 19266
rect 23257 19112 23303 19158
rect 23257 19005 23303 19051
rect 23257 18898 23303 18944
rect 23257 18791 23303 18837
rect 23257 18684 23303 18730
rect 23257 18577 23303 18623
rect 23257 18470 23303 18516
rect 23481 19760 23527 19806
rect 23481 19652 23527 19698
rect 23481 19544 23527 19590
rect 23481 19436 23527 19482
rect 23481 19328 23527 19374
rect 23481 19220 23527 19266
rect 23481 19112 23527 19158
rect 23481 19005 23527 19051
rect 23481 18898 23527 18944
rect 23481 18791 23527 18837
rect 23481 18684 23527 18730
rect 23481 18577 23527 18623
rect 23481 18470 23527 18516
rect 23176 17673 23222 17719
rect 23426 17673 23472 17719
rect 23679 17673 23725 17719
rect 23168 15112 23214 15158
rect 23168 15007 23214 15053
rect 23168 14902 23214 14948
rect 23168 14797 23214 14843
rect 23168 14692 23214 14738
rect 23168 14587 23214 14633
rect 23168 14482 23214 14528
rect 23392 15112 23438 15158
rect 23392 15007 23438 15053
rect 23392 14902 23438 14948
rect 23392 14797 23438 14843
rect 23392 14692 23438 14738
rect 23392 14587 23438 14633
rect 23392 14482 23438 14528
rect 23616 15112 23662 15158
rect 23616 15007 23662 15053
rect 23616 14902 23662 14948
rect 23616 14797 23662 14843
rect 23616 14692 23662 14738
rect 23616 14587 23662 14633
rect 23616 14482 23662 14528
rect 23172 10464 23218 10510
rect 23172 10361 23218 10407
rect 23172 10258 23218 10304
rect 23172 10155 23218 10201
rect 23172 10052 23218 10098
rect 23172 9949 23218 9995
rect 23172 9846 23218 9892
rect 23172 9743 23218 9789
rect 23172 9640 23218 9686
rect 23172 9537 23218 9583
rect 23172 9434 23218 9480
rect 23172 9331 23218 9377
rect 23172 9228 23218 9274
rect 23172 9125 23218 9171
rect 23172 9022 23218 9068
rect 23172 8919 23218 8965
rect 23172 8408 23218 8862
rect 23396 10464 23442 10510
rect 23396 10361 23442 10407
rect 23396 10258 23442 10304
rect 23396 10155 23442 10201
rect 23396 10052 23442 10098
rect 23396 9949 23442 9995
rect 23396 9846 23442 9892
rect 23396 9743 23442 9789
rect 23396 9640 23442 9686
rect 23396 9537 23442 9583
rect 23396 9434 23442 9480
rect 23396 9331 23442 9377
rect 23396 9228 23442 9274
rect 23396 9125 23442 9171
rect 23396 9022 23442 9068
rect 23396 8919 23442 8965
rect 23396 8408 23442 8862
rect 23620 10464 23666 10510
rect 23620 10361 23666 10407
rect 23620 10258 23666 10304
rect 23620 10155 23666 10201
rect 23620 10052 23666 10098
rect 23620 9949 23666 9995
rect 23620 9846 23666 9892
rect 23620 9743 23666 9789
rect 23620 9640 23666 9686
rect 23620 9537 23666 9583
rect 23620 9434 23666 9480
rect 23620 9331 23666 9377
rect 23620 9228 23666 9274
rect 23620 9125 23666 9171
rect 23620 9022 23666 9068
rect 23620 8919 23666 8965
rect 23620 8408 23666 8862
<< mvpsubdiff >>
rect 23622 22019 23782 22079
rect 23622 21973 23679 22019
rect 23725 21973 23782 22019
rect 23622 21913 23782 21973
rect 23228 16923 23688 16942
rect 23228 16877 23247 16923
rect 23669 16877 23688 16923
rect 23228 16858 23688 16877
rect 23176 13613 23652 13673
rect 23176 13567 23233 13613
rect 23279 13567 23391 13613
rect 23437 13567 23549 13613
rect 23595 13567 23652 13613
rect 23176 13507 23652 13567
<< mvnsubdiff >>
rect 23052 28924 23703 28981
rect 23052 28878 23211 28924
rect 23257 28878 23369 28924
rect 23415 28878 23527 28924
rect 23573 28878 23703 28924
rect 23052 28821 23703 28878
rect 23082 18174 23780 18231
rect 23082 18128 23205 18174
rect 23251 18128 23363 18174
rect 23409 18128 23521 18174
rect 23567 18128 23679 18174
rect 23725 18128 23780 18174
rect 23082 18071 23780 18128
rect 23121 15608 23593 15665
rect 23121 15562 23176 15608
rect 23222 15562 23334 15608
rect 23380 15562 23492 15608
rect 23538 15562 23593 15608
rect 23121 15505 23593 15562
rect 23004 7288 23159 7345
rect 23004 7242 23058 7288
rect 23104 7242 23159 7288
rect 23004 7185 23159 7242
rect 23548 7288 23703 7345
rect 23548 7242 23602 7288
rect 23648 7242 23703 7288
rect 23548 7185 23703 7242
<< mvpsubdiffcont >>
rect 23679 21973 23725 22019
rect 23247 16877 23669 16923
rect 23233 13567 23279 13613
rect 23391 13567 23437 13613
rect 23549 13567 23595 13613
<< mvnsubdiffcont >>
rect 23211 28878 23257 28924
rect 23369 28878 23415 28924
rect 23527 28878 23573 28924
rect 23205 18128 23251 18174
rect 23363 18128 23409 18174
rect 23521 18128 23567 18174
rect 23679 18128 23725 18174
rect 23176 15562 23222 15608
rect 23334 15562 23380 15608
rect 23492 15562 23538 15608
rect 23058 7242 23104 7288
rect 23602 7242 23648 7288
<< polysilicon >>
rect 50 39136 364 39155
rect 50 38996 69 39136
rect 115 39001 364 39136
rect 23648 39072 24018 39155
rect 23648 39026 23899 39072
rect 23945 39026 24018 39072
rect 23648 39001 24018 39026
rect 115 38996 134 39001
rect 50 38977 134 38996
rect 23826 38908 24018 39001
rect 23826 38862 23899 38908
rect 23945 38862 24018 38908
rect 23826 38816 24018 38862
rect 50 37477 364 37613
rect 50 37337 69 37477
rect 115 37459 364 37477
rect 23648 37512 24018 37613
rect 23648 37466 23899 37512
rect 23945 37466 24018 37512
rect 23648 37459 24018 37466
rect 115 37355 134 37459
rect 23826 37355 24018 37459
rect 115 37337 364 37355
rect 50 37201 364 37337
rect 23648 37348 24018 37355
rect 23648 37302 23899 37348
rect 23945 37302 24018 37348
rect 23648 37201 24018 37302
rect 50 35677 364 35813
rect 50 35537 69 35677
rect 115 35659 364 35677
rect 23648 35712 24018 35813
rect 23648 35666 23899 35712
rect 23945 35666 24018 35712
rect 23648 35659 24018 35666
rect 115 35555 134 35659
rect 23826 35555 24018 35659
rect 115 35537 364 35555
rect 50 35401 364 35537
rect 23648 35548 24018 35555
rect 23648 35502 23899 35548
rect 23945 35502 24018 35548
rect 23648 35401 24018 35502
rect 50 33877 364 34013
rect 50 33737 69 33877
rect 115 33859 364 33877
rect 23648 33912 24018 34013
rect 23648 33866 23899 33912
rect 23945 33866 24018 33912
rect 23648 33859 24018 33866
rect 115 33755 134 33859
rect 23826 33755 24018 33859
rect 115 33737 364 33755
rect 50 33601 364 33737
rect 23648 33748 24018 33755
rect 23648 33702 23899 33748
rect 23945 33702 24018 33748
rect 23648 33601 24018 33702
rect 50 32077 364 32213
rect 50 31937 69 32077
rect 115 32059 364 32077
rect 23648 32112 24018 32213
rect 23648 32066 23899 32112
rect 23945 32066 24018 32112
rect 23648 32059 24018 32066
rect 115 31955 134 32059
rect 23826 31955 24018 32059
rect 115 31937 364 31955
rect 50 31801 364 31937
rect 23648 31948 24018 31955
rect 23648 31902 23899 31948
rect 23945 31902 24018 31948
rect 23648 31801 24018 31902
rect 23826 30552 24018 30598
rect 23826 30506 23899 30552
rect 23945 30506 24018 30552
rect 50 30418 134 30437
rect 50 30278 69 30418
rect 115 30413 134 30418
rect 23826 30413 24018 30506
rect 115 30278 364 30413
rect 50 30259 364 30278
rect 23702 30388 24018 30413
rect 23702 30342 23899 30388
rect 23945 30342 24018 30388
rect 23702 30259 24018 30342
rect 361 29803 834 29858
rect 361 29757 414 29803
rect 460 29757 735 29803
rect 781 29757 834 29803
rect 361 29649 834 29757
rect 980 29803 1453 29858
rect 980 29757 1033 29803
rect 1079 29757 1354 29803
rect 1400 29757 1453 29803
rect 980 29649 1453 29757
rect 1599 29803 2072 29858
rect 1599 29757 1652 29803
rect 1698 29757 1973 29803
rect 2019 29757 2072 29803
rect 1599 29649 2072 29757
rect 2218 29803 2691 29858
rect 2218 29757 2271 29803
rect 2317 29757 2592 29803
rect 2638 29757 2691 29803
rect 2218 29649 2691 29757
rect 2837 29803 3310 29858
rect 2837 29757 2890 29803
rect 2936 29757 3211 29803
rect 3257 29757 3310 29803
rect 2837 29649 3310 29757
rect 3456 29803 3929 29858
rect 3456 29757 3509 29803
rect 3555 29757 3830 29803
rect 3876 29757 3929 29803
rect 3456 29649 3929 29757
rect 4075 29803 4548 29858
rect 4075 29757 4128 29803
rect 4174 29757 4449 29803
rect 4495 29757 4548 29803
rect 4075 29649 4548 29757
rect 4694 29803 5167 29858
rect 4694 29757 4747 29803
rect 4793 29757 5068 29803
rect 5114 29757 5167 29803
rect 4694 29649 5167 29757
rect 5313 29803 5786 29858
rect 5313 29757 5366 29803
rect 5412 29757 5687 29803
rect 5733 29757 5786 29803
rect 5313 29649 5786 29757
rect 5932 29803 6405 29858
rect 5932 29757 5985 29803
rect 6031 29757 6306 29803
rect 6352 29757 6405 29803
rect 5932 29649 6405 29757
rect 6551 29803 7024 29858
rect 6551 29757 6604 29803
rect 6650 29757 6925 29803
rect 6971 29757 7024 29803
rect 6551 29649 7024 29757
rect 7170 29803 7643 29858
rect 7170 29757 7223 29803
rect 7269 29757 7544 29803
rect 7590 29757 7643 29803
rect 7170 29649 7643 29757
rect 7789 29803 8262 29858
rect 7789 29757 7842 29803
rect 7888 29757 8163 29803
rect 8209 29757 8262 29803
rect 7789 29649 8262 29757
rect 8408 29803 8881 29858
rect 8408 29757 8461 29803
rect 8507 29757 8782 29803
rect 8828 29757 8881 29803
rect 8408 29649 8881 29757
rect 9027 29803 9500 29858
rect 9027 29757 9080 29803
rect 9126 29757 9401 29803
rect 9447 29757 9500 29803
rect 9027 29649 9500 29757
rect 9646 29803 10119 29858
rect 9646 29757 9699 29803
rect 9745 29757 10020 29803
rect 10066 29757 10119 29803
rect 9646 29649 10119 29757
rect 10265 29803 10738 29858
rect 10265 29757 10318 29803
rect 10364 29757 10639 29803
rect 10685 29757 10738 29803
rect 10265 29649 10738 29757
rect 10884 29803 11357 29858
rect 10884 29757 10937 29803
rect 10983 29757 11258 29803
rect 11304 29757 11357 29803
rect 10884 29649 11357 29757
rect 11503 29803 11976 29858
rect 11503 29757 11556 29803
rect 11602 29757 11877 29803
rect 11923 29757 11976 29803
rect 11503 29649 11976 29757
rect 12122 29803 12595 29858
rect 12122 29757 12175 29803
rect 12221 29757 12496 29803
rect 12542 29757 12595 29803
rect 12122 29649 12595 29757
rect 12741 29803 13214 29858
rect 12741 29757 12794 29803
rect 12840 29757 13115 29803
rect 13161 29757 13214 29803
rect 12741 29649 13214 29757
rect 13360 29803 13833 29858
rect 13360 29757 13413 29803
rect 13459 29757 13734 29803
rect 13780 29757 13833 29803
rect 13360 29649 13833 29757
rect 13979 29803 14452 29858
rect 13979 29757 14032 29803
rect 14078 29757 14353 29803
rect 14399 29757 14452 29803
rect 13979 29649 14452 29757
rect 14598 29803 15071 29858
rect 14598 29757 14651 29803
rect 14697 29757 14972 29803
rect 15018 29757 15071 29803
rect 14598 29649 15071 29757
rect 15217 29803 15690 29858
rect 15217 29757 15270 29803
rect 15316 29757 15591 29803
rect 15637 29757 15690 29803
rect 15217 29649 15690 29757
rect 15836 29803 16309 29858
rect 15836 29757 15889 29803
rect 15935 29757 16210 29803
rect 16256 29757 16309 29803
rect 15836 29649 16309 29757
rect 16455 29803 16928 29858
rect 16455 29757 16508 29803
rect 16554 29757 16829 29803
rect 16875 29757 16928 29803
rect 16455 29649 16928 29757
rect 17074 29803 17547 29858
rect 17074 29757 17127 29803
rect 17173 29757 17448 29803
rect 17494 29757 17547 29803
rect 17074 29649 17547 29757
rect 17693 29803 18166 29858
rect 17693 29757 17746 29803
rect 17792 29757 18067 29803
rect 18113 29757 18166 29803
rect 17693 29649 18166 29757
rect 18312 29803 18785 29858
rect 18312 29757 18365 29803
rect 18411 29757 18686 29803
rect 18732 29757 18785 29803
rect 18312 29649 18785 29757
rect 18931 29803 19404 29858
rect 18931 29757 18984 29803
rect 19030 29757 19305 29803
rect 19351 29757 19404 29803
rect 18931 29649 19404 29757
rect 19550 29803 20023 29858
rect 19550 29757 19603 29803
rect 19649 29757 19924 29803
rect 19970 29757 20023 29803
rect 19550 29649 20023 29757
rect 20169 29803 20642 29858
rect 20169 29757 20222 29803
rect 20268 29757 20543 29803
rect 20589 29757 20642 29803
rect 20169 29649 20642 29757
rect 20788 29803 21261 29858
rect 20788 29757 20841 29803
rect 20887 29757 21162 29803
rect 21208 29757 21261 29803
rect 20788 29649 21261 29757
rect 21407 29803 21880 29858
rect 21407 29757 21460 29803
rect 21506 29757 21781 29803
rect 21827 29757 21880 29803
rect 21407 29649 21880 29757
rect 22026 29803 22499 29858
rect 22026 29757 22079 29803
rect 22125 29757 22400 29803
rect 22446 29757 22499 29803
rect 22026 29649 22499 29757
rect 361 29112 834 29194
rect 980 29112 1453 29194
rect 1599 29112 2072 29194
rect 2218 29112 2691 29194
rect 2837 29112 3310 29194
rect 3456 29112 3929 29194
rect 4075 29112 4548 29194
rect 4694 29112 5167 29194
rect 5313 29112 5786 29194
rect 5932 29112 6405 29194
rect 6551 29112 7024 29194
rect 7170 29112 7643 29194
rect 7789 29112 8262 29194
rect 8408 29112 8881 29194
rect 9027 29112 9500 29194
rect 9646 29112 10119 29194
rect 10265 29112 10738 29194
rect 10884 29112 11357 29194
rect 11503 29112 11976 29194
rect 12122 29112 12595 29194
rect 12741 29112 13214 29194
rect 13360 29112 13833 29194
rect 13979 29112 14452 29194
rect 14598 29112 15071 29194
rect 15217 29112 15690 29194
rect 15836 29112 16309 29194
rect 16455 29112 16928 29194
rect 17074 29112 17547 29194
rect 17693 29112 18166 29194
rect 18312 29112 18785 29194
rect 18931 29112 19404 29194
rect 19550 29112 20023 29194
rect 20169 29112 20642 29194
rect 20788 29112 21261 29194
rect 21407 29112 21880 29194
rect 22026 29112 22499 29194
rect 23220 28632 23340 28705
rect 23444 28632 23564 28705
rect 23220 27857 23340 27950
rect 23444 27857 23564 27950
rect 23220 27115 23340 27175
rect 23444 27115 23564 27175
rect 23220 27093 23564 27115
rect 23220 27047 23328 27093
rect 23468 27047 23564 27093
rect 23220 27028 23564 27047
rect 23334 26956 23454 27028
rect 23334 25550 23454 25594
rect 23332 25369 23452 25413
rect 23332 23926 23452 24007
rect 23332 23880 23369 23926
rect 23415 23880 23452 23926
rect 23332 23861 23452 23880
rect 23332 23678 23452 23722
rect 23332 21674 23452 22316
rect 23332 20228 23452 20312
rect 23332 20182 23369 20228
rect 23415 20182 23452 20228
rect 23332 20163 23452 20182
rect 23332 19951 23452 19970
rect 23332 19905 23369 19951
rect 23415 19905 23452 19951
rect 23332 19819 23452 19905
rect 23332 18413 23452 18457
rect 23263 17984 23635 18003
rect 23263 17938 23426 17984
rect 23472 17938 23635 17984
rect 23263 17904 23635 17938
rect 23263 17844 23383 17904
rect 23515 17844 23635 17904
rect 23263 17360 23383 17547
rect 23515 17378 23635 17547
rect 23292 17329 23383 17360
rect 23516 17371 23635 17378
rect 23292 17256 23412 17329
rect 23516 17256 23636 17371
rect 23292 17069 23412 17142
rect 23516 17069 23636 17142
rect 23243 15171 23363 15215
rect 23467 15171 23587 15215
rect 23243 14409 23363 14469
rect 23467 14409 23587 14469
rect 23243 14393 23587 14409
rect 23243 14347 23876 14393
rect 23243 14301 23598 14347
rect 23644 14301 23756 14347
rect 23802 14301 23876 14347
rect 23243 14255 23876 14301
rect 23243 14246 23587 14255
rect 23243 14165 23363 14246
rect 23467 14165 23587 14246
rect 23243 13806 23363 13889
rect 23467 13806 23587 13889
rect 23247 12504 23367 12548
rect 23471 12504 23591 12548
rect 23247 10741 23367 10804
rect 23471 10741 23591 10804
rect 23247 10732 23591 10741
rect 22940 10686 23591 10732
rect 22940 10640 23014 10686
rect 23060 10640 23172 10686
rect 23218 10640 23591 10686
rect 22940 10594 23591 10640
rect 23247 10583 23591 10594
rect 23247 10523 23367 10583
rect 23471 10523 23591 10583
rect 23247 8351 23367 8395
rect 23471 8351 23591 8395
<< polycontact >>
rect 69 38996 115 39136
rect 23899 39026 23945 39072
rect 23899 38862 23945 38908
rect 69 37337 115 37477
rect 23899 37466 23945 37512
rect 23899 37302 23945 37348
rect 69 35537 115 35677
rect 23899 35666 23945 35712
rect 23899 35502 23945 35548
rect 69 33737 115 33877
rect 23899 33866 23945 33912
rect 23899 33702 23945 33748
rect 69 31937 115 32077
rect 23899 32066 23945 32112
rect 23899 31902 23945 31948
rect 23899 30506 23945 30552
rect 69 30278 115 30418
rect 23899 30342 23945 30388
rect 414 29757 460 29803
rect 735 29757 781 29803
rect 1033 29757 1079 29803
rect 1354 29757 1400 29803
rect 1652 29757 1698 29803
rect 1973 29757 2019 29803
rect 2271 29757 2317 29803
rect 2592 29757 2638 29803
rect 2890 29757 2936 29803
rect 3211 29757 3257 29803
rect 3509 29757 3555 29803
rect 3830 29757 3876 29803
rect 4128 29757 4174 29803
rect 4449 29757 4495 29803
rect 4747 29757 4793 29803
rect 5068 29757 5114 29803
rect 5366 29757 5412 29803
rect 5687 29757 5733 29803
rect 5985 29757 6031 29803
rect 6306 29757 6352 29803
rect 6604 29757 6650 29803
rect 6925 29757 6971 29803
rect 7223 29757 7269 29803
rect 7544 29757 7590 29803
rect 7842 29757 7888 29803
rect 8163 29757 8209 29803
rect 8461 29757 8507 29803
rect 8782 29757 8828 29803
rect 9080 29757 9126 29803
rect 9401 29757 9447 29803
rect 9699 29757 9745 29803
rect 10020 29757 10066 29803
rect 10318 29757 10364 29803
rect 10639 29757 10685 29803
rect 10937 29757 10983 29803
rect 11258 29757 11304 29803
rect 11556 29757 11602 29803
rect 11877 29757 11923 29803
rect 12175 29757 12221 29803
rect 12496 29757 12542 29803
rect 12794 29757 12840 29803
rect 13115 29757 13161 29803
rect 13413 29757 13459 29803
rect 13734 29757 13780 29803
rect 14032 29757 14078 29803
rect 14353 29757 14399 29803
rect 14651 29757 14697 29803
rect 14972 29757 15018 29803
rect 15270 29757 15316 29803
rect 15591 29757 15637 29803
rect 15889 29757 15935 29803
rect 16210 29757 16256 29803
rect 16508 29757 16554 29803
rect 16829 29757 16875 29803
rect 17127 29757 17173 29803
rect 17448 29757 17494 29803
rect 17746 29757 17792 29803
rect 18067 29757 18113 29803
rect 18365 29757 18411 29803
rect 18686 29757 18732 29803
rect 18984 29757 19030 29803
rect 19305 29757 19351 29803
rect 19603 29757 19649 29803
rect 19924 29757 19970 29803
rect 20222 29757 20268 29803
rect 20543 29757 20589 29803
rect 20841 29757 20887 29803
rect 21162 29757 21208 29803
rect 21460 29757 21506 29803
rect 21781 29757 21827 29803
rect 22079 29757 22125 29803
rect 22400 29757 22446 29803
rect 23328 27047 23468 27093
rect 23369 23880 23415 23926
rect 23369 20182 23415 20228
rect 23369 19905 23415 19951
rect 23426 17938 23472 17984
rect 23598 14301 23644 14347
rect 23756 14301 23802 14347
rect 23014 10640 23060 10686
rect 23172 10640 23218 10686
<< metal1 >>
rect 54 39136 130 39147
rect 54 39135 69 39136
rect 115 39135 130 39136
rect 54 38875 66 39135
rect 118 38875 130 39135
rect 54 38863 130 38875
rect 23858 39077 23982 39117
rect 23858 39025 23894 39077
rect 23946 39025 23982 39077
rect 23858 38908 23982 39025
rect 23858 38862 23899 38908
rect 23945 38862 23982 38908
rect 23858 38859 23982 38862
rect 23858 38807 23894 38859
rect 23946 38807 23982 38859
rect 23858 38767 23982 38807
rect 54 37537 130 37549
rect 54 37277 66 37537
rect 118 37277 130 37537
rect 54 37265 130 37277
rect 23858 37544 23982 37584
rect 23858 37492 23894 37544
rect 23946 37492 23982 37544
rect 23858 37466 23899 37492
rect 23945 37466 23982 37492
rect 23858 37348 23982 37466
rect 23858 37326 23899 37348
rect 23945 37326 23982 37348
rect 23858 37274 23894 37326
rect 23946 37274 23982 37326
rect 23858 37234 23982 37274
rect 54 35737 130 35749
rect 54 35477 66 35737
rect 118 35477 130 35737
rect 54 35465 130 35477
rect 23858 35740 23982 35780
rect 23858 35688 23894 35740
rect 23946 35688 23982 35740
rect 23858 35666 23899 35688
rect 23945 35666 23982 35688
rect 23858 35548 23982 35666
rect 23858 35522 23899 35548
rect 23945 35522 23982 35548
rect 23858 35470 23894 35522
rect 23946 35470 23982 35522
rect 23858 35430 23982 35470
rect 54 33937 130 33949
rect 54 33677 66 33937
rect 118 33677 130 33937
rect 54 33665 130 33677
rect 23858 33944 23982 33984
rect 23858 33892 23894 33944
rect 23946 33892 23982 33944
rect 23858 33866 23899 33892
rect 23945 33866 23982 33892
rect 23858 33748 23982 33866
rect 23858 33726 23899 33748
rect 23945 33726 23982 33748
rect 23858 33674 23894 33726
rect 23946 33674 23982 33726
rect 23858 33634 23982 33674
rect 54 32137 130 32149
rect 54 31877 66 32137
rect 118 31877 130 32137
rect 54 31865 130 31877
rect 23858 32140 23982 32180
rect 23858 32088 23894 32140
rect 23946 32088 23982 32140
rect 23858 32066 23899 32088
rect 23945 32066 23982 32088
rect 23858 31948 23982 32066
rect 23858 31922 23899 31948
rect 23945 31922 23982 31948
rect 23858 31870 23894 31922
rect 23946 31870 23982 31922
rect 23858 31830 23982 31870
rect 23858 30607 23982 30647
rect 23858 30555 23894 30607
rect 23946 30555 23982 30607
rect 23858 30552 23982 30555
rect 23858 30506 23899 30552
rect 23945 30506 23982 30552
rect 58 30418 126 30429
rect 58 30278 69 30418
rect 115 30278 126 30418
rect 23858 30389 23982 30506
rect 23858 30337 23894 30389
rect 23946 30337 23982 30389
rect 23858 30307 23982 30337
rect 23858 30297 24405 30307
rect 58 30267 126 30278
rect 1125 29890 1289 30213
rect 6525 29890 6689 30213
rect 11925 29890 12089 30213
rect 17325 29890 17489 30213
rect 22725 29997 22889 30213
rect 23945 30107 24405 30297
rect 22725 29985 22988 29997
rect 22725 29933 22800 29985
rect 22852 29933 22924 29985
rect 22976 29933 22988 29985
rect 22725 29890 22988 29933
rect 287 29878 25315 29890
rect 287 29826 948 29878
rect 1104 29826 11789 29878
rect 11945 29861 25315 29878
rect 11945 29826 22800 29861
rect 287 29809 22800 29826
rect 22852 29809 22924 29861
rect 22976 29809 25315 29861
rect 287 29803 25315 29809
rect 287 29757 414 29803
rect 460 29757 735 29803
rect 781 29757 1033 29803
rect 1079 29757 1354 29803
rect 1400 29757 1652 29803
rect 1698 29757 1973 29803
rect 2019 29757 2271 29803
rect 2317 29757 2592 29803
rect 2638 29757 2890 29803
rect 2936 29757 3211 29803
rect 3257 29757 3509 29803
rect 3555 29757 3830 29803
rect 3876 29757 4128 29803
rect 4174 29757 4449 29803
rect 4495 29757 4747 29803
rect 4793 29757 5068 29803
rect 5114 29757 5366 29803
rect 5412 29757 5687 29803
rect 5733 29757 5985 29803
rect 6031 29757 6306 29803
rect 6352 29757 6604 29803
rect 6650 29757 6925 29803
rect 6971 29757 7223 29803
rect 7269 29757 7544 29803
rect 7590 29757 7842 29803
rect 7888 29757 8163 29803
rect 8209 29757 8461 29803
rect 8507 29757 8782 29803
rect 8828 29757 9080 29803
rect 9126 29757 9401 29803
rect 9447 29757 9699 29803
rect 9745 29757 10020 29803
rect 10066 29757 10318 29803
rect 10364 29757 10639 29803
rect 10685 29757 10937 29803
rect 10983 29757 11258 29803
rect 11304 29757 11556 29803
rect 11602 29757 11877 29803
rect 11923 29757 12175 29803
rect 12221 29757 12496 29803
rect 12542 29757 12794 29803
rect 12840 29757 13115 29803
rect 13161 29757 13413 29803
rect 13459 29757 13734 29803
rect 13780 29757 14032 29803
rect 14078 29757 14353 29803
rect 14399 29757 14651 29803
rect 14697 29757 14972 29803
rect 15018 29757 15270 29803
rect 15316 29757 15591 29803
rect 15637 29757 15889 29803
rect 15935 29757 16210 29803
rect 16256 29757 16508 29803
rect 16554 29757 16829 29803
rect 16875 29757 17127 29803
rect 17173 29757 17448 29803
rect 17494 29757 17746 29803
rect 17792 29757 18067 29803
rect 18113 29757 18365 29803
rect 18411 29757 18686 29803
rect 18732 29757 18984 29803
rect 19030 29757 19305 29803
rect 19351 29757 19603 29803
rect 19649 29757 19924 29803
rect 19970 29757 20222 29803
rect 20268 29757 20543 29803
rect 20589 29757 20841 29803
rect 20887 29757 21162 29803
rect 21208 29757 21460 29803
rect 21506 29757 21781 29803
rect 21827 29757 22079 29803
rect 22125 29757 22400 29803
rect 22446 29757 25315 29803
rect 287 29720 25315 29757
rect 230 29604 346 29640
rect 230 29558 265 29604
rect 311 29558 346 29604
rect 230 29286 346 29558
rect 230 29240 265 29286
rect 311 29240 346 29286
rect 230 28890 346 29240
rect 849 29604 965 29640
rect 849 29558 884 29604
rect 930 29558 965 29604
rect 849 29286 965 29558
rect 849 29240 884 29286
rect 930 29240 965 29286
rect 849 28890 965 29240
rect 1468 29604 1584 29640
rect 1468 29558 1503 29604
rect 1549 29558 1584 29604
rect 1468 29286 1584 29558
rect 1468 29240 1503 29286
rect 1549 29240 1584 29286
rect 1468 28890 1584 29240
rect 2087 29604 2203 29640
rect 2087 29558 2122 29604
rect 2168 29558 2203 29604
rect 2087 29286 2203 29558
rect 2087 29240 2122 29286
rect 2168 29240 2203 29286
rect 2087 28890 2203 29240
rect 2706 29604 2822 29640
rect 2706 29558 2741 29604
rect 2787 29558 2822 29604
rect 2706 29286 2822 29558
rect 2706 29240 2741 29286
rect 2787 29240 2822 29286
rect 2706 28890 2822 29240
rect 3325 29604 3441 29640
rect 3325 29558 3360 29604
rect 3406 29558 3441 29604
rect 3325 29286 3441 29558
rect 3325 29240 3360 29286
rect 3406 29240 3441 29286
rect 3325 28890 3441 29240
rect 3944 29604 4060 29640
rect 3944 29558 3979 29604
rect 4025 29558 4060 29604
rect 3944 29286 4060 29558
rect 3944 29240 3979 29286
rect 4025 29240 4060 29286
rect 3944 28890 4060 29240
rect 4563 29604 4679 29640
rect 4563 29558 4598 29604
rect 4644 29558 4679 29604
rect 4563 29286 4679 29558
rect 4563 29240 4598 29286
rect 4644 29240 4679 29286
rect 4563 28890 4679 29240
rect 5182 29604 5298 29640
rect 5182 29558 5217 29604
rect 5263 29558 5298 29604
rect 5182 29286 5298 29558
rect 5182 29240 5217 29286
rect 5263 29240 5298 29286
rect 5182 28890 5298 29240
rect 5801 29604 5917 29640
rect 5801 29558 5836 29604
rect 5882 29558 5917 29604
rect 5801 29286 5917 29558
rect 5801 29240 5836 29286
rect 5882 29240 5917 29286
rect 5801 28890 5917 29240
rect 6420 29604 6536 29640
rect 6420 29558 6455 29604
rect 6501 29558 6536 29604
rect 6420 29286 6536 29558
rect 6420 29240 6455 29286
rect 6501 29240 6536 29286
rect 6420 28890 6536 29240
rect 7039 29604 7155 29640
rect 7039 29558 7074 29604
rect 7120 29558 7155 29604
rect 7039 29286 7155 29558
rect 7039 29240 7074 29286
rect 7120 29240 7155 29286
rect 7039 28890 7155 29240
rect 7658 29604 7774 29640
rect 7658 29558 7693 29604
rect 7739 29558 7774 29604
rect 7658 29286 7774 29558
rect 7658 29240 7693 29286
rect 7739 29240 7774 29286
rect 7658 28890 7774 29240
rect 8277 29604 8393 29640
rect 8277 29558 8312 29604
rect 8358 29558 8393 29604
rect 8277 29286 8393 29558
rect 8277 29240 8312 29286
rect 8358 29240 8393 29286
rect 8277 28890 8393 29240
rect 8896 29604 9012 29640
rect 8896 29558 8931 29604
rect 8977 29558 9012 29604
rect 8896 29286 9012 29558
rect 8896 29240 8931 29286
rect 8977 29240 9012 29286
rect 8896 28890 9012 29240
rect 9515 29604 9631 29640
rect 9515 29558 9550 29604
rect 9596 29558 9631 29604
rect 9515 29286 9631 29558
rect 9515 29240 9550 29286
rect 9596 29240 9631 29286
rect 9515 28890 9631 29240
rect 10134 29604 10250 29640
rect 10134 29558 10169 29604
rect 10215 29558 10250 29604
rect 10134 29286 10250 29558
rect 10134 29240 10169 29286
rect 10215 29240 10250 29286
rect 10134 28890 10250 29240
rect 10753 29604 10869 29640
rect 10753 29558 10788 29604
rect 10834 29558 10869 29604
rect 10753 29286 10869 29558
rect 10753 29240 10788 29286
rect 10834 29240 10869 29286
rect 10753 28890 10869 29240
rect 11372 29604 11488 29640
rect 11372 29558 11407 29604
rect 11453 29558 11488 29604
rect 11372 29286 11488 29558
rect 11372 29240 11407 29286
rect 11453 29240 11488 29286
rect 11372 28890 11488 29240
rect 11991 29604 12107 29640
rect 11991 29558 12026 29604
rect 12072 29558 12107 29604
rect 11991 29286 12107 29558
rect 11991 29240 12026 29286
rect 12072 29240 12107 29286
rect 11991 28890 12107 29240
rect 12610 29604 12726 29640
rect 12610 29558 12645 29604
rect 12691 29558 12726 29604
rect 12610 29286 12726 29558
rect 12610 29240 12645 29286
rect 12691 29240 12726 29286
rect 12610 28890 12726 29240
rect 13229 29604 13345 29640
rect 13229 29558 13264 29604
rect 13310 29558 13345 29604
rect 13229 29286 13345 29558
rect 13229 29240 13264 29286
rect 13310 29240 13345 29286
rect 13229 28890 13345 29240
rect 13848 29604 13964 29640
rect 13848 29558 13883 29604
rect 13929 29558 13964 29604
rect 13848 29286 13964 29558
rect 13848 29240 13883 29286
rect 13929 29240 13964 29286
rect 13848 28890 13964 29240
rect 14467 29604 14583 29640
rect 14467 29558 14502 29604
rect 14548 29558 14583 29604
rect 14467 29286 14583 29558
rect 14467 29240 14502 29286
rect 14548 29240 14583 29286
rect 14467 28890 14583 29240
rect 15086 29604 15202 29640
rect 15086 29558 15121 29604
rect 15167 29558 15202 29604
rect 15086 29286 15202 29558
rect 15086 29240 15121 29286
rect 15167 29240 15202 29286
rect 15086 28890 15202 29240
rect 15705 29604 15821 29640
rect 15705 29558 15740 29604
rect 15786 29558 15821 29604
rect 15705 29286 15821 29558
rect 15705 29240 15740 29286
rect 15786 29240 15821 29286
rect 15705 28890 15821 29240
rect 16324 29604 16440 29640
rect 16324 29558 16359 29604
rect 16405 29558 16440 29604
rect 16324 29286 16440 29558
rect 16324 29240 16359 29286
rect 16405 29240 16440 29286
rect 16324 28890 16440 29240
rect 16943 29604 17059 29640
rect 16943 29558 16978 29604
rect 17024 29558 17059 29604
rect 16943 29286 17059 29558
rect 16943 29240 16978 29286
rect 17024 29240 17059 29286
rect 16943 28890 17059 29240
rect 17562 29604 17678 29640
rect 17562 29558 17597 29604
rect 17643 29558 17678 29604
rect 17562 29286 17678 29558
rect 17562 29240 17597 29286
rect 17643 29240 17678 29286
rect 17562 28890 17678 29240
rect 18181 29604 18297 29640
rect 18181 29558 18216 29604
rect 18262 29558 18297 29604
rect 18181 29286 18297 29558
rect 18181 29240 18216 29286
rect 18262 29240 18297 29286
rect 18181 28890 18297 29240
rect 18800 29604 18916 29640
rect 18800 29558 18835 29604
rect 18881 29558 18916 29604
rect 18800 29286 18916 29558
rect 18800 29240 18835 29286
rect 18881 29240 18916 29286
rect 18800 28890 18916 29240
rect 19419 29604 19535 29640
rect 19419 29558 19454 29604
rect 19500 29558 19535 29604
rect 19419 29286 19535 29558
rect 19419 29240 19454 29286
rect 19500 29240 19535 29286
rect 19419 28890 19535 29240
rect 20038 29604 20154 29640
rect 20038 29558 20073 29604
rect 20119 29558 20154 29604
rect 20038 29286 20154 29558
rect 20038 29240 20073 29286
rect 20119 29240 20154 29286
rect 20038 28890 20154 29240
rect 20657 29604 20773 29640
rect 20657 29558 20692 29604
rect 20738 29558 20773 29604
rect 20657 29286 20773 29558
rect 20657 29240 20692 29286
rect 20738 29240 20773 29286
rect 20657 28890 20773 29240
rect 21276 29604 21392 29640
rect 21276 29558 21311 29604
rect 21357 29558 21392 29604
rect 21276 29286 21392 29558
rect 21276 29240 21311 29286
rect 21357 29240 21392 29286
rect 21276 28890 21392 29240
rect 21895 29604 22011 29640
rect 21895 29558 21930 29604
rect 21976 29558 22011 29604
rect 21895 29286 22011 29558
rect 21895 29240 21930 29286
rect 21976 29240 22011 29286
rect 21895 28890 22011 29240
rect 22514 29604 22630 29640
rect 22514 29558 22549 29604
rect 22595 29558 22630 29604
rect 22514 29286 22630 29558
rect 22514 29240 22549 29286
rect 22595 29240 22630 29286
rect 22514 28890 22630 29240
rect 230 28725 22630 28890
rect 23082 28962 23760 28986
rect 23082 28924 23369 28962
rect 23421 28924 23760 28962
rect 23082 28878 23211 28924
rect 23257 28878 23369 28924
rect 23421 28910 23527 28924
rect 23415 28878 23527 28910
rect 23573 28878 23760 28924
rect 23082 28776 23760 28878
rect 23082 28724 23369 28776
rect 23421 28724 23760 28776
rect 23082 28703 23760 28724
rect 23082 28587 23230 28703
rect 23082 28541 23143 28587
rect 23189 28541 23230 28587
rect 23082 28405 23230 28541
rect 23082 28359 23143 28405
rect 23189 28359 23230 28405
rect 23082 28224 23230 28359
rect 23082 28178 23143 28224
rect 23189 28178 23230 28224
rect 23082 28042 23230 28178
rect 23082 27996 23143 28042
rect 23189 27996 23230 28042
rect 23082 27811 23230 27996
rect 23335 28587 23450 28623
rect 23335 28541 23369 28587
rect 23415 28541 23450 28587
rect 23335 28405 23450 28541
rect 23335 28359 23369 28405
rect 23415 28372 23450 28405
rect 23335 28224 23386 28359
rect 23335 28178 23369 28224
rect 23438 28216 23450 28372
rect 23415 28178 23450 28216
rect 23335 28042 23450 28178
rect 23335 27996 23369 28042
rect 23415 27996 23450 28042
rect 23335 27959 23450 27996
rect 23555 28587 23760 28703
rect 23555 28541 23679 28587
rect 23725 28541 23760 28587
rect 23555 28405 23760 28541
rect 23555 28359 23679 28405
rect 23725 28359 23760 28405
rect 23555 28224 23760 28359
rect 23555 28178 23679 28224
rect 23725 28178 23760 28224
rect 23555 28042 23760 28178
rect 23555 27996 23679 28042
rect 23725 27996 23760 28042
rect 23082 27765 23143 27811
rect 23189 27765 23230 27811
rect 23082 27630 23230 27765
rect 23082 27584 23143 27630
rect 23189 27584 23230 27630
rect 23082 27449 23230 27584
rect 23082 27403 23143 27449
rect 23189 27403 23230 27449
rect 23082 27267 23230 27403
rect 23082 27221 23143 27267
rect 23189 27221 23230 27267
rect 23082 27184 23230 27221
rect 23335 27811 23450 27848
rect 23335 27765 23369 27811
rect 23415 27765 23450 27811
rect 23335 27630 23450 27765
rect 23335 27593 23369 27630
rect 23335 27437 23347 27593
rect 23415 27584 23450 27630
rect 23399 27449 23450 27584
rect 23335 27403 23369 27437
rect 23415 27403 23450 27449
rect 23335 27267 23450 27403
rect 23335 27221 23369 27267
rect 23415 27221 23450 27267
rect 23335 27184 23450 27221
rect 23555 27811 23760 27996
rect 23555 27765 23679 27811
rect 23725 27765 23760 27811
rect 23555 27630 23760 27765
rect 23555 27584 23679 27630
rect 23725 27584 23760 27630
rect 23555 27449 23760 27584
rect 23555 27403 23679 27449
rect 23725 27403 23760 27449
rect 23555 27267 23760 27403
rect 23555 27221 23679 27267
rect 23725 27221 23760 27267
rect 23555 27184 23760 27221
rect 22263 27031 22913 27105
rect 23249 27093 23624 27104
rect 23249 27047 23328 27093
rect 23468 27047 23624 27093
rect 23249 27030 23624 27047
rect 23259 26943 23305 26956
rect 23259 26835 23305 26897
rect 23259 26727 23305 26789
rect 23259 26619 23305 26681
rect 23259 26511 23305 26573
rect 23259 26417 23305 26465
rect 23144 26405 23305 26417
rect 23144 26249 23156 26405
rect 23208 26403 23305 26405
rect 23208 26357 23259 26403
rect 23208 26295 23305 26357
rect 23208 26249 23259 26295
rect 23144 26237 23305 26249
rect 23259 26188 23305 26237
rect 23259 26081 23305 26142
rect 23259 25974 23305 26035
rect 23259 25867 23305 25928
rect 23259 25760 23305 25821
rect 23259 25653 23305 25714
rect 23259 25594 23305 25607
rect 23483 26943 23529 26956
rect 23483 26835 23529 26897
rect 23483 26727 23529 26789
rect 23483 26619 23529 26681
rect 23483 26511 23529 26573
rect 23483 26417 23529 26465
rect 23483 26405 23644 26417
rect 23483 26403 23580 26405
rect 23529 26357 23580 26403
rect 23483 26295 23580 26357
rect 23529 26249 23580 26295
rect 23632 26249 23644 26405
rect 23483 26237 23644 26249
rect 23483 26188 23529 26237
rect 23483 26081 23529 26142
rect 23483 25974 23529 26035
rect 23483 25867 23529 25928
rect 23483 25760 23529 25821
rect 23483 25653 23529 25714
rect 23483 25594 23529 25607
rect 23153 25357 23635 25369
rect 23153 25356 23571 25357
rect 23153 25310 23257 25356
rect 23303 25310 23481 25356
rect 23527 25310 23571 25356
rect 23153 25248 23571 25310
rect 23153 25202 23257 25248
rect 23303 25202 23481 25248
rect 23527 25202 23571 25248
rect 23153 25201 23571 25202
rect 23623 25201 23635 25357
rect 23153 25189 23635 25201
rect 23153 25140 23632 25189
rect 23153 25094 23257 25140
rect 23303 25094 23481 25140
rect 23527 25094 23632 25140
rect 23153 25032 23632 25094
rect 23153 24986 23257 25032
rect 23303 24986 23481 25032
rect 23527 24986 23632 25032
rect 23153 24924 23632 24986
rect 23153 24878 23257 24924
rect 23303 24878 23481 24924
rect 23527 24878 23632 24924
rect 23153 24816 23632 24878
rect 23153 24770 23257 24816
rect 23303 24770 23481 24816
rect 23527 24770 23632 24816
rect 23153 24708 23632 24770
rect 23153 24662 23257 24708
rect 23303 24662 23481 24708
rect 23527 24662 23632 24708
rect 23153 24601 23632 24662
rect 23153 24555 23257 24601
rect 23303 24555 23481 24601
rect 23527 24555 23632 24601
rect 23153 24494 23632 24555
rect 23153 24448 23257 24494
rect 23303 24448 23481 24494
rect 23527 24448 23632 24494
rect 23153 24387 23632 24448
rect 23153 24341 23257 24387
rect 23303 24341 23481 24387
rect 23527 24341 23632 24387
rect 23153 24280 23632 24341
rect 23153 24234 23257 24280
rect 23303 24234 23481 24280
rect 23527 24234 23632 24280
rect 23153 24173 23632 24234
rect 23153 24127 23257 24173
rect 23303 24127 23481 24173
rect 23527 24127 23632 24173
rect 23153 24066 23632 24127
rect 23153 24020 23257 24066
rect 23303 24020 23481 24066
rect 23527 24020 23632 24066
rect 23153 24007 23632 24020
rect 23153 23678 23223 24007
rect 23302 23926 23483 23937
rect 23302 23922 23369 23926
rect 23302 23766 23349 23922
rect 23415 23880 23483 23926
rect 23401 23766 23483 23880
rect 23302 23754 23483 23766
rect 23561 23678 23632 24007
rect 23153 23665 23303 23678
rect 23153 23619 23257 23665
rect 23153 23557 23303 23619
rect 23153 23511 23257 23557
rect 23153 23449 23303 23511
rect 23153 23403 23257 23449
rect 23153 23341 23303 23403
rect 23153 23295 23257 23341
rect 23153 23233 23303 23295
rect 23153 23187 23257 23233
rect 23153 23125 23303 23187
rect 23153 23079 23257 23125
rect 23153 23017 23303 23079
rect 23153 22971 23257 23017
rect 23153 22910 23303 22971
rect 23153 22864 23257 22910
rect 23153 22803 23303 22864
rect 23153 22757 23257 22803
rect 23153 22696 23303 22757
rect 23153 22650 23257 22696
rect 23153 22589 23303 22650
rect 23153 22543 23257 22589
rect 23153 22482 23303 22543
rect 23153 22436 23257 22482
rect 23153 22416 23303 22436
rect 23481 23665 23632 23678
rect 23527 23619 23632 23665
rect 23481 23557 23632 23619
rect 23527 23511 23632 23557
rect 23481 23449 23632 23511
rect 23527 23403 23632 23449
rect 23481 23341 23632 23403
rect 23527 23295 23632 23341
rect 23481 23233 23632 23295
rect 23527 23187 23632 23233
rect 23481 23125 23632 23187
rect 23527 23079 23632 23125
rect 23481 23017 23632 23079
rect 23527 22971 23632 23017
rect 23481 22910 23632 22971
rect 23527 22864 23632 22910
rect 23481 22803 23632 22864
rect 23527 22757 23632 22803
rect 23481 22696 23632 22757
rect 23527 22650 23632 22696
rect 23481 22589 23632 22650
rect 23527 22543 23632 22589
rect 23481 22482 23632 22543
rect 23527 22436 23632 22482
rect 23153 22375 23338 22416
rect 23153 22329 23257 22375
rect 23303 22329 23338 22375
rect 23153 22326 23338 22329
rect 23245 22246 23338 22326
rect 23481 22375 23632 22436
rect 23527 22329 23632 22375
rect 23481 22316 23632 22329
rect 23245 22242 23657 22246
rect 23245 22222 23856 22242
rect 23245 22170 23578 22222
rect 23630 22170 23764 22222
rect 23816 22170 23856 22222
rect 23245 22150 23856 22170
rect 23245 22149 23657 22150
rect 23631 22065 23773 22070
rect 23082 22024 23773 22065
rect 23082 21972 23536 22024
rect 23588 22019 23773 22024
rect 23588 21973 23679 22019
rect 23725 21973 23773 22019
rect 23588 21972 23773 21973
rect 23082 21931 23773 21972
rect 23631 21922 23773 21931
rect 23141 21820 23654 21843
rect 23141 21768 23156 21820
rect 23208 21768 23654 21820
rect 23141 21746 23654 21768
rect 23561 21674 23654 21746
rect 23153 21661 23303 21674
rect 23153 21615 23257 21661
rect 23153 21553 23303 21615
rect 23153 21507 23257 21553
rect 23153 21445 23303 21507
rect 23153 21399 23257 21445
rect 23153 21337 23303 21399
rect 23153 21291 23257 21337
rect 23153 21229 23303 21291
rect 23153 21183 23257 21229
rect 23153 21121 23303 21183
rect 23153 21075 23257 21121
rect 23153 21013 23303 21075
rect 23153 20967 23257 21013
rect 23153 20906 23303 20967
rect 23153 20860 23257 20906
rect 23153 20799 23303 20860
rect 23153 20753 23257 20799
rect 23153 20692 23303 20753
rect 23153 20646 23257 20692
rect 23153 20585 23303 20646
rect 23153 20539 23257 20585
rect 23153 20478 23303 20539
rect 23153 20432 23257 20478
rect 23153 20371 23303 20432
rect 23153 20325 23257 20371
rect 23153 20312 23303 20325
rect 23481 21661 23654 21674
rect 23527 21615 23654 21661
rect 23481 21553 23654 21615
rect 23527 21507 23654 21553
rect 23481 21445 23654 21507
rect 23527 21399 23654 21445
rect 23481 21337 23654 21399
rect 23527 21291 23654 21337
rect 23481 21229 23654 21291
rect 23527 21183 23654 21229
rect 23481 21121 23654 21183
rect 23527 21075 23654 21121
rect 23481 21013 23654 21075
rect 23527 20967 23654 21013
rect 23481 20906 23654 20967
rect 23527 20860 23654 20906
rect 23481 20799 23654 20860
rect 23527 20753 23654 20799
rect 23481 20692 23654 20753
rect 23527 20646 23654 20692
rect 23481 20585 23654 20646
rect 23527 20539 23654 20585
rect 23481 20478 23654 20539
rect 23527 20432 23654 20478
rect 23481 20371 23654 20432
rect 23527 20325 23654 20371
rect 23481 20312 23654 20325
rect 23153 19819 23223 20312
rect 23302 20228 23483 20242
rect 23302 20182 23369 20228
rect 23415 20182 23483 20228
rect 23302 20179 23483 20182
rect 23302 20127 23364 20179
rect 23416 20127 23483 20179
rect 23302 20107 23483 20127
rect 23302 19984 23483 20027
rect 23302 19932 23314 19984
rect 23470 19932 23483 19984
rect 23302 19905 23369 19932
rect 23415 19905 23483 19932
rect 23302 19891 23483 19905
rect 23561 19819 23654 20312
rect 23153 19818 23303 19819
rect 23481 19818 23654 19819
rect 23153 19806 23654 19818
rect 23153 19760 23257 19806
rect 23303 19760 23481 19806
rect 23527 19760 23654 19806
rect 23153 19698 23654 19760
rect 23153 19652 23257 19698
rect 23303 19652 23481 19698
rect 23527 19652 23654 19698
rect 23153 19590 23654 19652
rect 23153 19544 23257 19590
rect 23303 19544 23481 19590
rect 23527 19544 23654 19590
rect 23153 19482 23654 19544
rect 23153 19436 23257 19482
rect 23303 19436 23481 19482
rect 23527 19436 23654 19482
rect 23153 19374 23654 19436
rect 23153 19328 23257 19374
rect 23303 19328 23481 19374
rect 23527 19328 23654 19374
rect 23153 19266 23654 19328
rect 23153 19220 23257 19266
rect 23303 19220 23481 19266
rect 23527 19220 23654 19266
rect 23153 19158 23654 19220
rect 23153 19112 23257 19158
rect 23303 19112 23481 19158
rect 23527 19112 23654 19158
rect 23153 19051 23654 19112
rect 23153 19005 23257 19051
rect 23303 19005 23481 19051
rect 23527 19005 23654 19051
rect 23153 18944 23654 19005
rect 23153 18898 23257 18944
rect 23303 18898 23481 18944
rect 23527 18898 23654 18944
rect 23153 18837 23654 18898
rect 23153 18791 23257 18837
rect 23303 18791 23481 18837
rect 23527 18791 23654 18837
rect 23153 18730 23654 18791
rect 23153 18684 23257 18730
rect 23303 18684 23481 18730
rect 23527 18684 23654 18730
rect 23153 18623 23654 18684
rect 23153 18577 23257 18623
rect 23303 18577 23481 18623
rect 23527 18577 23654 18623
rect 23153 18516 23654 18577
rect 23153 18470 23257 18516
rect 23303 18470 23481 18516
rect 23527 18470 23654 18516
rect 23153 18467 23654 18470
rect 23153 18457 23552 18467
rect 23153 18433 23338 18457
rect 22779 18313 23338 18433
rect 22779 16586 22895 18313
rect 23082 18183 23760 18211
rect 23082 18131 23139 18183
rect 23191 18174 23319 18183
rect 23371 18174 23760 18183
rect 23191 18131 23205 18174
rect 23082 18128 23205 18131
rect 23251 18131 23319 18174
rect 23251 18128 23363 18131
rect 23409 18128 23521 18174
rect 23567 18128 23679 18174
rect 23725 18128 23760 18174
rect 23082 18091 23760 18128
rect 23082 17835 23153 18091
rect 23518 18011 23760 18091
rect 23257 17988 23760 18011
rect 23257 17936 23295 17988
rect 23347 17984 23760 17988
rect 23347 17938 23426 17984
rect 23472 17938 23760 17984
rect 23347 17936 23760 17938
rect 23257 17914 23760 17936
rect 23082 17719 23256 17835
rect 23082 17673 23176 17719
rect 23222 17673 23256 17719
rect 23082 17556 23256 17673
rect 23379 17823 23507 17835
rect 23379 17719 23443 17823
rect 23379 17673 23426 17719
rect 23379 17667 23443 17673
rect 23495 17667 23507 17823
rect 23379 17556 23507 17667
rect 23645 17719 23759 17914
rect 23645 17673 23679 17719
rect 23725 17673 23759 17719
rect 23645 17556 23759 17673
rect 23082 17222 23263 17259
rect 23082 17176 23217 17222
rect 23082 17030 23263 17176
rect 23414 17222 23487 17556
rect 23414 17176 23441 17222
rect 23414 17139 23487 17176
rect 23645 17222 23760 17259
rect 23645 17176 23665 17222
rect 23711 17176 23760 17222
rect 23645 17030 23760 17176
rect 23082 16939 23760 17030
rect 23082 16923 23366 16939
rect 23418 16923 23760 16939
rect 23082 16877 23247 16923
rect 23669 16877 23760 16923
rect 23082 16835 23760 16877
rect 22779 16466 23910 16586
rect 23141 15609 23573 15645
rect 23141 15608 23216 15609
rect 23268 15608 23402 15609
rect 23141 15562 23176 15608
rect 23268 15562 23334 15608
rect 23380 15562 23402 15608
rect 23141 15557 23216 15562
rect 23268 15557 23402 15562
rect 23454 15608 23573 15609
rect 23454 15562 23492 15608
rect 23538 15562 23573 15608
rect 23454 15557 23573 15562
rect 23141 15525 23573 15557
rect 23168 15158 23214 15171
rect 23168 15053 23214 15112
rect 23144 15015 23168 15045
rect 23392 15158 23438 15171
rect 23392 15053 23438 15112
rect 23214 15015 23236 15045
rect 23144 14963 23164 15015
rect 23216 14963 23236 15015
rect 23144 14948 23236 14963
rect 23144 14902 23168 14948
rect 23214 14902 23236 14948
rect 23144 14843 23236 14902
rect 23144 14829 23168 14843
rect 23214 14829 23236 14843
rect 23144 14777 23164 14829
rect 23216 14777 23236 14829
rect 23616 15158 23662 15171
rect 23616 15053 23662 15112
rect 23392 14948 23438 15007
rect 23392 14843 23438 14902
rect 23392 14783 23438 14797
rect 23592 15015 23616 15045
rect 23662 15015 23684 15045
rect 23592 14963 23612 15015
rect 23664 14963 23684 15015
rect 23592 14948 23684 14963
rect 23592 14902 23616 14948
rect 23662 14902 23684 14948
rect 23592 14843 23684 14902
rect 23592 14829 23616 14843
rect 23662 14829 23684 14843
rect 23144 14738 23236 14777
rect 23144 14737 23168 14738
rect 23214 14737 23236 14738
rect 23356 14738 23473 14783
rect 23168 14633 23214 14692
rect 23168 14528 23214 14587
rect 23168 14469 23214 14482
rect 23356 14692 23392 14738
rect 23438 14692 23473 14738
rect 23592 14777 23612 14829
rect 23664 14777 23684 14829
rect 23592 14738 23684 14777
rect 23592 14737 23616 14738
rect 23356 14633 23473 14692
rect 23356 14587 23392 14633
rect 23438 14587 23473 14633
rect 23356 14528 23473 14587
rect 23356 14482 23392 14528
rect 23438 14482 23473 14528
rect 23356 14398 23473 14482
rect 23662 14737 23684 14738
rect 23616 14633 23662 14692
rect 23616 14528 23662 14587
rect 23616 14469 23662 14482
rect 22955 14323 23473 14398
rect 23793 14384 23910 16466
rect 22955 10723 23027 14323
rect 23168 14152 23214 14165
rect 23132 13902 23168 13938
rect 23356 14152 23473 14323
rect 23563 14347 23910 14384
rect 23563 14301 23598 14347
rect 23644 14301 23756 14347
rect 23802 14301 23910 14347
rect 23563 14264 23910 14301
rect 23356 14060 23392 14152
rect 23214 13902 23249 13938
rect 23132 13664 23249 13902
rect 23438 14060 23473 14152
rect 23616 14152 23662 14165
rect 23392 13889 23438 13902
rect 23580 13902 23616 13938
rect 23662 13902 23697 13938
rect 23580 13664 23697 13902
rect 23132 13613 23697 13664
rect 23132 13567 23233 13613
rect 23279 13567 23391 13613
rect 23437 13567 23549 13613
rect 23595 13567 23697 13613
rect 23132 13516 23697 13567
rect 23132 12576 23249 13516
rect 23132 12524 23169 12576
rect 23221 12524 23249 12576
rect 23132 12491 23249 12524
rect 23132 12390 23172 12491
rect 23218 12390 23249 12491
rect 23132 12338 23169 12390
rect 23221 12338 23249 12390
rect 23132 12038 23172 12338
rect 23218 12038 23249 12338
rect 23132 11986 23169 12038
rect 23221 11986 23249 12038
rect 23132 11852 23172 11986
rect 23218 11852 23249 11986
rect 23132 11800 23169 11852
rect 23221 11800 23249 11852
rect 23132 11719 23172 11800
rect 23149 11433 23172 11463
rect 23218 11719 23249 11800
rect 23356 12576 23486 12616
rect 23356 12524 23395 12576
rect 23447 12524 23486 12576
rect 23356 12491 23486 12524
rect 23356 12358 23396 12491
rect 23442 12358 23486 12491
rect 23356 12306 23395 12358
rect 23447 12306 23486 12358
rect 23356 12140 23396 12306
rect 23442 12140 23486 12306
rect 23356 12088 23395 12140
rect 23447 12088 23486 12140
rect 23356 11923 23396 12088
rect 23442 11923 23486 12088
rect 23356 11871 23395 11923
rect 23447 11871 23486 11923
rect 23356 11705 23396 11871
rect 23442 11705 23486 11871
rect 23580 12576 23697 13516
rect 23580 12524 23610 12576
rect 23662 12524 23697 12576
rect 23580 12491 23697 12524
rect 23580 12390 23620 12491
rect 23580 12338 23610 12390
rect 23580 12038 23620 12338
rect 23580 11986 23610 12038
rect 23580 11852 23620 11986
rect 23580 11800 23610 11852
rect 23580 11719 23620 11800
rect 23356 11653 23395 11705
rect 23447 11653 23486 11705
rect 23356 11487 23396 11653
rect 23442 11487 23486 11653
rect 23218 11433 23241 11463
rect 23149 11381 23169 11433
rect 23221 11381 23241 11433
rect 23149 11247 23172 11381
rect 23218 11247 23241 11381
rect 23149 11195 23169 11247
rect 23221 11195 23241 11247
rect 23149 11155 23172 11195
rect 23218 11155 23241 11195
rect 23356 11435 23395 11487
rect 23447 11435 23486 11487
rect 23356 11270 23396 11435
rect 23442 11270 23486 11435
rect 23356 11218 23395 11270
rect 23447 11218 23486 11270
rect 23172 10804 23218 10817
rect 23356 11052 23396 11218
rect 23442 11052 23486 11218
rect 23590 11433 23620 11463
rect 23666 11719 23697 12491
rect 23590 11381 23610 11433
rect 23590 11247 23620 11381
rect 23590 11195 23610 11247
rect 23590 11155 23620 11195
rect 23356 11000 23395 11052
rect 23447 11000 23486 11052
rect 23356 10835 23396 11000
rect 23442 10835 23486 11000
rect 23356 10783 23395 10835
rect 23447 10783 23486 10835
rect 23666 11155 23682 11463
rect 23620 10804 23666 10817
rect 22955 10686 23253 10723
rect 22955 10640 23014 10686
rect 23060 10640 23172 10686
rect 23218 10640 23253 10686
rect 22955 10603 23253 10640
rect 23356 10617 23486 10783
rect 23356 10565 23395 10617
rect 23447 10565 23486 10617
rect 23172 10510 23218 10523
rect 23172 10407 23218 10464
rect 23172 10304 23218 10361
rect 23172 10201 23218 10258
rect 23172 10098 23218 10155
rect 23172 9995 23218 10052
rect 23172 9892 23218 9949
rect 23172 9789 23218 9846
rect 23172 9686 23218 9743
rect 23172 9583 23218 9640
rect 23172 9480 23218 9537
rect 23172 9377 23218 9434
rect 23172 9274 23218 9331
rect 23172 9171 23218 9228
rect 23172 9068 23218 9125
rect 23172 8965 23218 9022
rect 23172 8862 23218 8919
rect 23137 8408 23172 8519
rect 23356 10510 23486 10565
rect 23356 10464 23396 10510
rect 23442 10464 23486 10510
rect 23356 10407 23486 10464
rect 23356 10399 23396 10407
rect 23442 10399 23486 10407
rect 23356 10347 23395 10399
rect 23447 10347 23486 10399
rect 23356 10304 23486 10347
rect 23356 10258 23396 10304
rect 23442 10258 23486 10304
rect 23356 10201 23486 10258
rect 23356 10182 23396 10201
rect 23442 10182 23486 10201
rect 23356 10130 23395 10182
rect 23447 10130 23486 10182
rect 23356 10098 23486 10130
rect 23356 10052 23396 10098
rect 23442 10052 23486 10098
rect 23356 9995 23486 10052
rect 23356 9964 23396 9995
rect 23442 9964 23486 9995
rect 23356 9912 23395 9964
rect 23447 9912 23486 9964
rect 23356 9892 23486 9912
rect 23356 9846 23396 9892
rect 23442 9846 23486 9892
rect 23356 9789 23486 9846
rect 23356 9746 23396 9789
rect 23442 9746 23486 9789
rect 23356 9694 23395 9746
rect 23447 9694 23486 9746
rect 23356 9686 23486 9694
rect 23356 9640 23396 9686
rect 23442 9640 23486 9686
rect 23356 9583 23486 9640
rect 23356 9537 23396 9583
rect 23442 9537 23486 9583
rect 23356 9529 23486 9537
rect 23356 9477 23395 9529
rect 23447 9477 23486 9529
rect 23356 9434 23396 9477
rect 23442 9434 23486 9477
rect 23356 9377 23486 9434
rect 23356 9331 23396 9377
rect 23442 9331 23486 9377
rect 23356 9311 23486 9331
rect 23356 9259 23395 9311
rect 23447 9259 23486 9311
rect 23356 9228 23396 9259
rect 23442 9228 23486 9259
rect 23356 9171 23486 9228
rect 23356 9125 23396 9171
rect 23442 9125 23486 9171
rect 23356 9093 23486 9125
rect 23356 9041 23395 9093
rect 23447 9041 23486 9093
rect 23356 9022 23396 9041
rect 23442 9022 23486 9041
rect 23356 8965 23486 9022
rect 23356 8919 23396 8965
rect 23442 8919 23486 8965
rect 23356 8876 23486 8919
rect 23356 8824 23395 8876
rect 23447 8824 23486 8876
rect 23356 8658 23396 8824
rect 23442 8658 23486 8824
rect 23356 8606 23395 8658
rect 23447 8606 23486 8658
rect 23218 8408 23253 8519
rect 23137 7774 23253 8408
rect 23137 7722 23173 7774
rect 23225 7722 23253 7774
rect 23137 7588 23253 7722
rect 23137 7536 23173 7588
rect 23225 7536 23253 7588
rect 23137 7402 23253 7536
rect 23137 7350 23173 7402
rect 23225 7350 23253 7402
rect 23137 7325 23253 7350
rect 23024 7288 23253 7325
rect 23024 7242 23058 7288
rect 23104 7242 23253 7288
rect 23024 7205 23253 7242
rect 23356 8441 23396 8606
rect 23442 8441 23486 8606
rect 23620 10510 23666 10523
rect 23620 10407 23666 10464
rect 23620 10304 23666 10361
rect 23620 10201 23666 10258
rect 23620 10098 23666 10155
rect 23620 9995 23666 10052
rect 23620 9892 23666 9949
rect 23620 9789 23666 9846
rect 23620 9686 23666 9743
rect 23620 9583 23666 9640
rect 23620 9480 23666 9537
rect 23620 9377 23666 9434
rect 23620 9274 23666 9331
rect 23620 9171 23666 9228
rect 23620 9068 23666 9125
rect 23620 8965 23666 9022
rect 23620 8862 23666 8919
rect 23356 8389 23395 8441
rect 23447 8389 23486 8441
rect 23356 8223 23486 8389
rect 23356 8171 23395 8223
rect 23447 8171 23486 8223
rect 23356 8005 23486 8171
rect 23356 7953 23395 8005
rect 23447 7953 23486 8005
rect 23356 7788 23486 7953
rect 23356 7736 23395 7788
rect 23447 7736 23486 7788
rect 23356 7570 23486 7736
rect 23356 7518 23395 7570
rect 23447 7518 23486 7570
rect 23356 7352 23486 7518
rect 23356 7300 23395 7352
rect 23447 7300 23486 7352
rect 23585 8408 23620 8519
rect 23666 8408 23701 8519
rect 23585 7774 23701 8408
rect 23585 7722 23615 7774
rect 23667 7722 23701 7774
rect 23585 7588 23701 7722
rect 23585 7536 23615 7588
rect 23667 7536 23701 7588
rect 23585 7402 23701 7536
rect 23585 7350 23615 7402
rect 23667 7350 23701 7402
rect 23585 7325 23701 7350
rect 23356 7042 23486 7300
rect 23568 7288 23701 7325
rect 23568 7242 23602 7288
rect 23648 7242 23701 7288
rect 23568 7205 23701 7242
rect 23308 5013 23530 7042
rect 23259 4973 23599 5013
rect 23259 4921 23297 4973
rect 23349 4921 23509 4973
rect 23561 4921 23599 4973
rect 23259 4755 23599 4921
rect 23259 4703 23297 4755
rect 23349 4703 23509 4755
rect 23561 4703 23599 4755
rect 23259 4662 23599 4703
<< via1 >>
rect 66 38996 69 39135
rect 69 38996 115 39135
rect 115 38996 118 39135
rect 66 38875 118 38996
rect 23894 39072 23946 39077
rect 23894 39026 23899 39072
rect 23899 39026 23945 39072
rect 23945 39026 23946 39072
rect 23894 39025 23946 39026
rect 23894 38807 23946 38859
rect 66 37477 118 37537
rect 66 37337 69 37477
rect 69 37337 115 37477
rect 115 37337 118 37477
rect 66 37277 118 37337
rect 23894 37512 23946 37544
rect 23894 37492 23899 37512
rect 23899 37492 23945 37512
rect 23945 37492 23946 37512
rect 23894 37302 23899 37326
rect 23899 37302 23945 37326
rect 23945 37302 23946 37326
rect 23894 37274 23946 37302
rect 66 35677 118 35737
rect 66 35537 69 35677
rect 69 35537 115 35677
rect 115 35537 118 35677
rect 66 35477 118 35537
rect 23894 35712 23946 35740
rect 23894 35688 23899 35712
rect 23899 35688 23945 35712
rect 23945 35688 23946 35712
rect 23894 35502 23899 35522
rect 23899 35502 23945 35522
rect 23945 35502 23946 35522
rect 23894 35470 23946 35502
rect 66 33877 118 33937
rect 66 33737 69 33877
rect 69 33737 115 33877
rect 115 33737 118 33877
rect 66 33677 118 33737
rect 23894 33912 23946 33944
rect 23894 33892 23899 33912
rect 23899 33892 23945 33912
rect 23945 33892 23946 33912
rect 23894 33702 23899 33726
rect 23899 33702 23945 33726
rect 23945 33702 23946 33726
rect 23894 33674 23946 33702
rect 66 32077 118 32137
rect 66 31937 69 32077
rect 69 31937 115 32077
rect 115 31937 118 32077
rect 66 31877 118 31937
rect 23894 32112 23946 32140
rect 23894 32088 23899 32112
rect 23899 32088 23945 32112
rect 23945 32088 23946 32112
rect 23894 31902 23899 31922
rect 23899 31902 23945 31922
rect 23945 31902 23946 31922
rect 23894 31870 23946 31902
rect 23894 30555 23946 30607
rect 23894 30388 23946 30389
rect 23894 30342 23899 30388
rect 23899 30342 23945 30388
rect 23945 30342 23946 30388
rect 23894 30337 23946 30342
rect 22800 29933 22852 29985
rect 22924 29933 22976 29985
rect 948 29826 1104 29878
rect 11789 29826 11945 29878
rect 22800 29809 22852 29861
rect 22924 29809 22976 29861
rect 23369 28924 23421 28962
rect 23369 28910 23415 28924
rect 23415 28910 23421 28924
rect 23369 28724 23421 28776
rect 23386 28359 23415 28372
rect 23415 28359 23438 28372
rect 23386 28224 23438 28359
rect 23386 28216 23415 28224
rect 23415 28216 23438 28224
rect 23347 27584 23369 27593
rect 23369 27584 23399 27593
rect 23347 27449 23399 27584
rect 23347 27437 23369 27449
rect 23369 27437 23399 27449
rect 23156 26249 23208 26405
rect 23580 26249 23632 26405
rect 23571 25201 23623 25357
rect 23349 23880 23369 23922
rect 23369 23880 23401 23922
rect 23349 23766 23401 23880
rect 23578 22170 23630 22222
rect 23764 22170 23816 22222
rect 23536 21972 23588 22024
rect 23156 21768 23208 21820
rect 23364 20127 23416 20179
rect 23314 19951 23470 19984
rect 23314 19932 23369 19951
rect 23369 19932 23415 19951
rect 23415 19932 23470 19951
rect 23139 18131 23191 18183
rect 23319 18174 23371 18183
rect 23319 18131 23363 18174
rect 23363 18131 23371 18174
rect 23295 17936 23347 17988
rect 23443 17719 23495 17823
rect 23443 17673 23472 17719
rect 23472 17673 23495 17719
rect 23443 17667 23495 17673
rect 23366 16923 23418 16939
rect 23366 16887 23418 16923
rect 23216 15608 23268 15609
rect 23216 15562 23222 15608
rect 23222 15562 23268 15608
rect 23216 15557 23268 15562
rect 23402 15557 23454 15609
rect 23164 15007 23168 15015
rect 23168 15007 23214 15015
rect 23214 15007 23216 15015
rect 23164 14963 23216 15007
rect 23164 14797 23168 14829
rect 23168 14797 23214 14829
rect 23214 14797 23216 14829
rect 23164 14777 23216 14797
rect 23612 15007 23616 15015
rect 23616 15007 23662 15015
rect 23662 15007 23664 15015
rect 23612 14963 23664 15007
rect 23612 14797 23616 14829
rect 23616 14797 23662 14829
rect 23662 14797 23664 14829
rect 23612 14777 23664 14797
rect 23169 12524 23221 12576
rect 23169 12338 23172 12390
rect 23172 12338 23218 12390
rect 23218 12338 23221 12390
rect 23169 11986 23172 12038
rect 23172 11986 23218 12038
rect 23218 11986 23221 12038
rect 23169 11800 23172 11852
rect 23172 11800 23218 11852
rect 23218 11800 23221 11852
rect 23395 12524 23447 12576
rect 23395 12306 23396 12358
rect 23396 12306 23442 12358
rect 23442 12306 23447 12358
rect 23395 12088 23396 12140
rect 23396 12088 23442 12140
rect 23442 12088 23447 12140
rect 23395 11871 23396 11923
rect 23396 11871 23442 11923
rect 23442 11871 23447 11923
rect 23610 12524 23662 12576
rect 23610 12338 23620 12390
rect 23620 12338 23662 12390
rect 23610 11986 23620 12038
rect 23620 11986 23662 12038
rect 23610 11800 23620 11852
rect 23620 11800 23662 11852
rect 23395 11653 23396 11705
rect 23396 11653 23442 11705
rect 23442 11653 23447 11705
rect 23169 11381 23172 11433
rect 23172 11381 23218 11433
rect 23218 11381 23221 11433
rect 23169 11195 23172 11247
rect 23172 11195 23218 11247
rect 23218 11195 23221 11247
rect 23395 11435 23396 11487
rect 23396 11435 23442 11487
rect 23442 11435 23447 11487
rect 23395 11218 23396 11270
rect 23396 11218 23442 11270
rect 23442 11218 23447 11270
rect 23610 11381 23620 11433
rect 23620 11381 23662 11433
rect 23610 11195 23620 11247
rect 23620 11195 23662 11247
rect 23395 11000 23396 11052
rect 23396 11000 23442 11052
rect 23442 11000 23447 11052
rect 23395 10817 23396 10835
rect 23396 10817 23442 10835
rect 23442 10817 23447 10835
rect 23395 10783 23447 10817
rect 23395 10565 23447 10617
rect 23395 10361 23396 10399
rect 23396 10361 23442 10399
rect 23442 10361 23447 10399
rect 23395 10347 23447 10361
rect 23395 10155 23396 10182
rect 23396 10155 23442 10182
rect 23442 10155 23447 10182
rect 23395 10130 23447 10155
rect 23395 9949 23396 9964
rect 23396 9949 23442 9964
rect 23442 9949 23447 9964
rect 23395 9912 23447 9949
rect 23395 9743 23396 9746
rect 23396 9743 23442 9746
rect 23442 9743 23447 9746
rect 23395 9694 23447 9743
rect 23395 9480 23447 9529
rect 23395 9477 23396 9480
rect 23396 9477 23442 9480
rect 23442 9477 23447 9480
rect 23395 9274 23447 9311
rect 23395 9259 23396 9274
rect 23396 9259 23442 9274
rect 23442 9259 23447 9274
rect 23395 9068 23447 9093
rect 23395 9041 23396 9068
rect 23396 9041 23442 9068
rect 23442 9041 23447 9068
rect 23395 8862 23447 8876
rect 23395 8824 23396 8862
rect 23396 8824 23442 8862
rect 23442 8824 23447 8862
rect 23395 8606 23396 8658
rect 23396 8606 23442 8658
rect 23442 8606 23447 8658
rect 23173 7722 23225 7774
rect 23173 7536 23225 7588
rect 23173 7350 23225 7402
rect 23395 8408 23396 8441
rect 23396 8408 23442 8441
rect 23442 8408 23447 8441
rect 23395 8389 23447 8408
rect 23395 8171 23447 8223
rect 23395 7953 23447 8005
rect 23395 7736 23447 7788
rect 23395 7518 23447 7570
rect 23395 7300 23447 7352
rect 23615 7722 23667 7774
rect 23615 7536 23667 7588
rect 23615 7350 23667 7402
rect 23297 4921 23349 4973
rect 23509 4921 23561 4973
rect 23297 4703 23349 4755
rect 23509 4703 23561 4755
<< metal2 >>
rect 54 39135 130 39147
rect 54 38875 66 39135
rect 118 38875 130 39135
rect 54 37537 130 38875
rect 54 37277 66 37537
rect 118 37277 130 37537
rect 54 35737 130 37277
rect 23857 39077 23982 39117
rect 23857 39025 23894 39077
rect 23946 39025 23982 39077
rect 23857 38859 23982 39025
rect 23857 38807 23894 38859
rect 23946 38807 23982 38859
rect 23857 37544 23982 38807
rect 23857 37492 23894 37544
rect 23946 37492 23982 37544
rect 23857 37326 23982 37492
rect 23857 37274 23894 37326
rect 23946 37274 23982 37326
rect 23857 37140 23982 37274
rect 54 35477 66 35737
rect 118 35477 130 35737
rect 54 33937 130 35477
rect 54 33677 66 33937
rect 118 33677 130 33937
rect 54 32137 130 33677
rect 54 31877 66 32137
rect 118 31877 130 32137
rect 54 30351 130 31877
rect 23857 35740 23982 36714
rect 23857 35688 23894 35740
rect 23946 35688 23982 35740
rect 23857 35522 23982 35688
rect 23857 35470 23894 35522
rect 23946 35470 23982 35522
rect 23857 33944 23982 35470
rect 23857 33892 23894 33944
rect 23946 33892 23982 33944
rect 23857 33726 23982 33892
rect 23857 33674 23894 33726
rect 23946 33674 23982 33726
rect 23857 32140 23982 33674
rect 23857 32088 23894 32140
rect 23946 32088 23982 32140
rect 23857 31922 23982 32088
rect 23857 31870 23894 31922
rect 23946 31870 23982 31922
rect 52 30341 130 30351
rect 52 30077 62 30341
rect 118 30106 130 30341
rect 118 30077 128 30106
rect 52 30067 128 30077
rect 976 29987 1077 31182
rect 976 29931 996 29987
rect 1052 29931 1077 29987
rect 976 29890 1077 29931
rect 936 29878 1116 29890
rect 936 29826 948 29878
rect 1104 29826 1116 29878
rect 936 29814 996 29826
rect 976 29799 996 29814
rect 1052 29814 1116 29826
rect 1052 29799 1077 29814
rect 976 29723 1077 29799
rect 976 29667 996 29723
rect 1052 29667 1077 29723
rect 976 29591 1077 29667
rect 976 29535 996 29591
rect 1052 29535 1077 29591
rect 976 29471 1077 29535
rect 1337 29071 1437 31182
rect 11777 29987 11877 31182
rect 11777 29931 11798 29987
rect 11854 29931 11877 29987
rect 11777 29890 11877 29931
rect 11777 29878 11957 29890
rect 11777 29826 11789 29878
rect 11945 29826 11957 29878
rect 11777 29799 11798 29826
rect 11854 29814 11957 29826
rect 11854 29799 11877 29814
rect 11777 29723 11877 29799
rect 11777 29667 11798 29723
rect 11854 29667 11877 29723
rect 11777 29591 11877 29667
rect 11777 29535 11798 29591
rect 11854 29535 11877 29591
rect 11777 29471 11877 29535
rect 1337 29015 1358 29071
rect 1414 29015 1437 29071
rect 1337 28939 1437 29015
rect 1337 28883 1358 28939
rect 1414 28883 1437 28939
rect 1337 28807 1437 28883
rect 1337 28751 1358 28807
rect 1414 28751 1437 28807
rect 1337 28675 1437 28751
rect 1337 28619 1358 28675
rect 1414 28619 1437 28675
rect 1337 28543 1437 28619
rect 1337 28487 1358 28543
rect 1414 28487 1437 28543
rect 1337 28411 1437 28487
rect 1337 28355 1358 28411
rect 1414 28355 1437 28411
rect 1337 28279 1437 28355
rect 1337 28223 1358 28279
rect 1414 28223 1437 28279
rect 1337 28147 1437 28223
rect 1337 28091 1358 28147
rect 1414 28091 1437 28147
rect 1337 28015 1437 28091
rect 1337 27959 1358 28015
rect 1414 27959 1437 28015
rect 1337 27883 1437 27959
rect 1337 27827 1358 27883
rect 1414 27827 1437 27883
rect 1337 27751 1437 27827
rect 1337 27695 1358 27751
rect 1414 27695 1437 27751
rect 1337 27619 1437 27695
rect 1337 27563 1358 27619
rect 1414 27563 1437 27619
rect 1337 27527 1437 27563
rect 12137 29071 12237 31182
rect 12137 29015 12158 29071
rect 12214 29015 12237 29071
rect 12137 28939 12237 29015
rect 12137 28883 12158 28939
rect 12214 28883 12237 28939
rect 12137 28807 12237 28883
rect 12137 28751 12158 28807
rect 12214 28751 12237 28807
rect 12137 28675 12237 28751
rect 12137 28619 12158 28675
rect 12214 28619 12237 28675
rect 12137 28543 12237 28619
rect 12137 28487 12158 28543
rect 12214 28487 12237 28543
rect 12137 28411 12237 28487
rect 12137 28355 12158 28411
rect 12214 28355 12237 28411
rect 12137 28279 12237 28355
rect 12137 28223 12158 28279
rect 12214 28223 12237 28279
rect 12137 28147 12237 28223
rect 12137 28091 12158 28147
rect 12214 28091 12237 28147
rect 12137 28015 12237 28091
rect 12137 27959 12158 28015
rect 12214 27959 12237 28015
rect 12137 27883 12237 27959
rect 12137 27827 12158 27883
rect 12214 27827 12237 27883
rect 12137 27751 12237 27827
rect 12137 27695 12158 27751
rect 12214 27695 12237 27751
rect 12137 27619 12237 27695
rect 12137 27563 12158 27619
rect 12214 27563 12237 27619
rect 12137 27527 12237 27563
rect 22577 29071 22677 31182
rect 22937 29997 23037 31182
rect 23857 30879 23982 31870
rect 23858 30607 23982 30647
rect 23858 30555 23894 30607
rect 23946 30555 23982 30607
rect 22788 29987 23037 29997
rect 22788 29985 22958 29987
rect 22788 29933 22800 29985
rect 22852 29933 22924 29985
rect 22788 29931 22958 29933
rect 23014 29931 23037 29987
rect 22788 29861 23037 29931
rect 22788 29809 22800 29861
rect 22852 29809 22924 29861
rect 22976 29855 23037 29861
rect 22788 29799 22958 29809
rect 23014 29799 23037 29855
rect 22788 29797 23037 29799
rect 22577 29015 22598 29071
rect 22654 29015 22677 29071
rect 22577 28939 22677 29015
rect 22577 28883 22598 28939
rect 22654 28883 22677 28939
rect 22577 28807 22677 28883
rect 22577 28751 22598 28807
rect 22654 28751 22677 28807
rect 22577 28675 22677 28751
rect 22577 28619 22598 28675
rect 22654 28619 22677 28675
rect 22577 28543 22677 28619
rect 22577 28487 22598 28543
rect 22654 28487 22677 28543
rect 22577 28411 22677 28487
rect 22577 28355 22598 28411
rect 22654 28355 22677 28411
rect 22577 28279 22677 28355
rect 22577 28223 22598 28279
rect 22654 28223 22677 28279
rect 22577 28147 22677 28223
rect 22577 28091 22598 28147
rect 22654 28091 22677 28147
rect 22577 28015 22677 28091
rect 22577 27959 22598 28015
rect 22654 27959 22677 28015
rect 22577 27883 22677 27959
rect 22577 27827 22598 27883
rect 22654 27827 22677 27883
rect 22577 27751 22677 27827
rect 22577 27695 22598 27751
rect 22654 27695 22677 27751
rect 22577 27619 22677 27695
rect 22577 27563 22598 27619
rect 22654 27563 22677 27619
rect 22577 27527 22677 27563
rect 22937 29723 23037 29797
rect 22937 29667 22958 29723
rect 23014 29667 23037 29723
rect 22937 29591 23037 29667
rect 22937 29535 22958 29591
rect 23014 29535 23037 29591
rect 22937 27527 23037 29535
rect 23197 29350 23317 30533
rect 23154 29252 23317 29350
rect 23497 29350 23617 30533
rect 23858 30472 23982 30555
rect 23857 30389 23982 30472
rect 23857 30337 23894 30389
rect 23946 30337 23982 30389
rect 23857 30297 23982 30337
rect 23497 29252 23625 29350
rect 23154 27543 23210 29252
rect 23328 28964 23456 28986
rect 23328 28908 23367 28964
rect 23423 28908 23456 28964
rect 23328 28778 23456 28908
rect 23328 28722 23367 28778
rect 23423 28722 23456 28778
rect 23328 28703 23456 28722
rect 23374 28372 23450 28384
rect 23374 28216 23386 28372
rect 23438 28322 23450 28372
rect 23569 28322 23625 29252
rect 23438 28266 23625 28322
rect 23438 28216 23450 28266
rect 23374 28204 23450 28216
rect 23335 27593 23411 27605
rect 23335 27543 23347 27593
rect 23154 27487 23347 27543
rect 23154 26417 23210 27487
rect 23335 27437 23347 27487
rect 23399 27437 23411 27593
rect 23335 27425 23411 27437
rect 23569 26417 23625 28266
rect 23144 26405 23220 26417
rect 23144 26249 23156 26405
rect 23208 26249 23220 26405
rect 23144 26237 23220 26249
rect 23568 26405 23644 26417
rect 23568 26249 23580 26405
rect 23632 26249 23644 26405
rect 23568 26237 23644 26249
rect 23154 21832 23210 26237
rect 23569 25369 23625 26237
rect 23559 25357 23635 25369
rect 23559 25201 23571 25357
rect 23623 25201 23635 25357
rect 23559 25189 23635 25201
rect 23337 23922 23413 23934
rect 23337 23766 23349 23922
rect 23401 23766 23413 23922
rect 23337 23754 23413 23766
rect 23144 21820 23220 21832
rect 23144 21768 23156 21820
rect 23208 21768 23220 21820
rect 23144 21756 23220 21768
rect 23347 21571 23403 23754
rect 23569 22344 23625 25189
rect 23548 22222 23856 22242
rect 23548 22170 23578 22222
rect 23630 22170 23764 22222
rect 23816 22170 23856 22222
rect 23548 22150 23856 22170
rect 23497 22026 23626 22065
rect 23497 21970 23534 22026
rect 23590 21970 23626 22026
rect 23497 21931 23626 21970
rect 23498 21808 23626 21931
rect 23498 21752 23534 21808
rect 23590 21752 23626 21808
rect 23498 21714 23626 21752
rect 23347 21515 23621 21571
rect 23129 20179 23452 20203
rect 23129 20127 23364 20179
rect 23416 20127 23452 20179
rect 23129 20106 23452 20127
rect 23129 18612 23221 20106
rect 23565 19996 23621 21515
rect 23302 19984 23621 19996
rect 23302 19932 23314 19984
rect 23470 19932 23621 19984
rect 23302 19920 23621 19932
rect 23129 18515 23320 18612
rect 23227 18206 23320 18515
rect 23101 18185 23409 18206
rect 23101 18129 23137 18185
rect 23193 18129 23317 18185
rect 23373 18129 23409 18185
rect 23101 18109 23409 18129
rect 23227 18011 23320 18109
rect 23227 17988 23386 18011
rect 23227 17936 23295 17988
rect 23347 17936 23386 17988
rect 23227 17914 23386 17936
rect 23565 17835 23621 19920
rect 23431 17823 23621 17835
rect 23431 17667 23443 17823
rect 23495 17779 23621 17823
rect 23495 17667 23507 17779
rect 23431 17655 23507 17667
rect 23328 16941 23456 17037
rect 23328 16885 23364 16941
rect 23420 16885 23456 16941
rect 23328 16808 23456 16885
rect 23768 16758 23856 22150
rect 23186 15611 23494 15629
rect 23186 15555 23214 15611
rect 23270 15555 23400 15611
rect 23456 15555 23494 15611
rect 23186 15537 23494 15555
rect 23144 15017 23236 15045
rect 23144 14961 23162 15017
rect 23218 14961 23236 15017
rect 23144 14831 23236 14961
rect 23144 14775 23162 14831
rect 23218 14775 23236 14831
rect 23144 14737 23236 14775
rect 23592 15017 23684 15045
rect 23592 14961 23610 15017
rect 23666 14961 23684 15017
rect 23592 14831 23684 14961
rect 23592 14775 23610 14831
rect 23666 14775 23684 14831
rect 23592 14737 23684 14775
rect 23149 12578 23241 12606
rect 23149 12522 23167 12578
rect 23223 12522 23241 12578
rect 23149 12392 23241 12522
rect 23149 12336 23167 12392
rect 23223 12336 23241 12392
rect 23149 12298 23241 12336
rect 23356 12576 23486 12616
rect 23356 12524 23395 12576
rect 23447 12524 23486 12576
rect 23356 12358 23486 12524
rect 23356 12306 23395 12358
rect 23447 12306 23486 12358
rect 23356 12140 23486 12306
rect 23590 12578 23682 12606
rect 23590 12522 23608 12578
rect 23664 12522 23682 12578
rect 23590 12392 23682 12522
rect 23590 12336 23608 12392
rect 23664 12336 23682 12392
rect 23590 12298 23682 12336
rect 23356 12088 23395 12140
rect 23447 12088 23486 12140
rect 23149 12040 23241 12068
rect 23149 11984 23167 12040
rect 23223 11984 23241 12040
rect 23149 11854 23241 11984
rect 23149 11798 23167 11854
rect 23223 11798 23241 11854
rect 23149 11760 23241 11798
rect 23356 11923 23486 12088
rect 23356 11871 23395 11923
rect 23447 11871 23486 11923
rect 23356 11705 23486 11871
rect 23590 12040 23682 12068
rect 23590 11984 23608 12040
rect 23664 11984 23682 12040
rect 23590 11854 23682 11984
rect 23590 11798 23608 11854
rect 23664 11798 23682 11854
rect 23590 11760 23682 11798
rect 23356 11653 23395 11705
rect 23447 11653 23486 11705
rect 23356 11487 23486 11653
rect 23149 11435 23241 11463
rect 23149 11379 23167 11435
rect 23223 11379 23241 11435
rect 23149 11249 23241 11379
rect 23149 11193 23167 11249
rect 23223 11193 23241 11249
rect 23149 11155 23241 11193
rect 23356 11435 23395 11487
rect 23447 11435 23486 11487
rect 23356 11270 23486 11435
rect 23356 11218 23395 11270
rect 23447 11218 23486 11270
rect 23356 11052 23486 11218
rect 23590 11435 23682 11463
rect 23590 11379 23608 11435
rect 23664 11379 23682 11435
rect 23590 11249 23682 11379
rect 23590 11193 23608 11249
rect 23664 11193 23682 11249
rect 23590 11155 23682 11193
rect 23356 11000 23395 11052
rect 23447 11000 23486 11052
rect 23356 10835 23486 11000
rect 23356 10783 23395 10835
rect 23447 10783 23486 10835
rect 23356 10617 23486 10783
rect 23356 10565 23395 10617
rect 23447 10565 23486 10617
rect 23356 10399 23486 10565
rect 23356 10347 23395 10399
rect 23447 10347 23486 10399
rect 23356 10182 23486 10347
rect 23356 10130 23395 10182
rect 23447 10130 23486 10182
rect 23356 9964 23486 10130
rect 23356 9912 23395 9964
rect 23447 9912 23486 9964
rect 23356 9746 23486 9912
rect 23356 9694 23395 9746
rect 23447 9694 23486 9746
rect 23356 9529 23486 9694
rect 23356 9477 23395 9529
rect 23447 9477 23486 9529
rect 23356 9311 23486 9477
rect 23356 9259 23395 9311
rect 23447 9259 23486 9311
rect 23356 9093 23486 9259
rect 23356 9041 23395 9093
rect 23447 9041 23486 9093
rect 23356 8876 23486 9041
rect 23356 8824 23395 8876
rect 23447 8824 23486 8876
rect 23356 8658 23486 8824
rect 23356 8606 23395 8658
rect 23447 8606 23486 8658
rect 23356 8441 23486 8606
rect 23356 8389 23395 8441
rect 23447 8389 23486 8441
rect 23356 8223 23486 8389
rect 23356 8171 23395 8223
rect 23447 8171 23486 8223
rect 23356 8005 23486 8171
rect 23356 7953 23395 8005
rect 23447 7953 23486 8005
rect 23153 7776 23245 7804
rect 23153 7720 23171 7776
rect 23227 7720 23245 7776
rect 23153 7590 23245 7720
rect 23153 7534 23171 7590
rect 23227 7534 23245 7590
rect 23153 7404 23245 7534
rect 23153 7348 23171 7404
rect 23227 7348 23245 7404
rect 23153 7310 23245 7348
rect 23356 7788 23486 7953
rect 23356 7736 23395 7788
rect 23447 7736 23486 7788
rect 23356 7570 23486 7736
rect 23356 7518 23395 7570
rect 23447 7518 23486 7570
rect 23356 7352 23486 7518
rect 23356 7300 23395 7352
rect 23447 7300 23486 7352
rect 23595 7776 23687 7804
rect 23595 7720 23613 7776
rect 23669 7720 23687 7776
rect 23595 7590 23687 7720
rect 23595 7534 23613 7590
rect 23669 7534 23687 7590
rect 23595 7404 23687 7534
rect 23595 7348 23613 7404
rect 23669 7348 23687 7404
rect 23595 7310 23687 7348
rect 23356 5014 23486 7300
rect 23259 4975 23599 5014
rect 23259 4919 23295 4975
rect 23351 4919 23507 4975
rect 23563 4919 23599 4975
rect 23259 4757 23599 4919
rect 23259 4701 23295 4757
rect 23351 4701 23507 4757
rect 23563 4701 23599 4757
rect 23259 4662 23599 4701
<< via2 >>
rect 62 30077 118 30341
rect 996 29931 1052 29987
rect 996 29826 1052 29855
rect 996 29799 1052 29826
rect 996 29667 1052 29723
rect 996 29535 1052 29591
rect 11798 29931 11854 29987
rect 11798 29826 11854 29855
rect 11798 29799 11854 29826
rect 11798 29667 11854 29723
rect 11798 29535 11854 29591
rect 1358 29015 1414 29071
rect 1358 28883 1414 28939
rect 1358 28751 1414 28807
rect 1358 28619 1414 28675
rect 1358 28487 1414 28543
rect 1358 28355 1414 28411
rect 1358 28223 1414 28279
rect 1358 28091 1414 28147
rect 1358 27959 1414 28015
rect 1358 27827 1414 27883
rect 1358 27695 1414 27751
rect 1358 27563 1414 27619
rect 12158 29015 12214 29071
rect 12158 28883 12214 28939
rect 12158 28751 12214 28807
rect 12158 28619 12214 28675
rect 12158 28487 12214 28543
rect 12158 28355 12214 28411
rect 12158 28223 12214 28279
rect 12158 28091 12214 28147
rect 12158 27959 12214 28015
rect 12158 27827 12214 27883
rect 12158 27695 12214 27751
rect 12158 27563 12214 27619
rect 22958 29985 23014 29987
rect 22958 29933 22976 29985
rect 22976 29933 23014 29985
rect 22958 29931 23014 29933
rect 22958 29809 22976 29855
rect 22976 29809 23014 29855
rect 22958 29799 23014 29809
rect 22598 29015 22654 29071
rect 22598 28883 22654 28939
rect 22598 28751 22654 28807
rect 22598 28619 22654 28675
rect 22598 28487 22654 28543
rect 22598 28355 22654 28411
rect 22598 28223 22654 28279
rect 22598 28091 22654 28147
rect 22598 27959 22654 28015
rect 22598 27827 22654 27883
rect 22598 27695 22654 27751
rect 22598 27563 22654 27619
rect 22958 29667 23014 29723
rect 22958 29535 23014 29591
rect 23367 28962 23423 28964
rect 23367 28910 23369 28962
rect 23369 28910 23421 28962
rect 23421 28910 23423 28962
rect 23367 28908 23423 28910
rect 23367 28776 23423 28778
rect 23367 28724 23369 28776
rect 23369 28724 23421 28776
rect 23421 28724 23423 28776
rect 23367 28722 23423 28724
rect 23534 22024 23590 22026
rect 23534 21972 23536 22024
rect 23536 21972 23588 22024
rect 23588 21972 23590 22024
rect 23534 21970 23590 21972
rect 23534 21752 23590 21808
rect 23137 18183 23193 18185
rect 23137 18131 23139 18183
rect 23139 18131 23191 18183
rect 23191 18131 23193 18183
rect 23137 18129 23193 18131
rect 23317 18183 23373 18185
rect 23317 18131 23319 18183
rect 23319 18131 23371 18183
rect 23371 18131 23373 18183
rect 23317 18129 23373 18131
rect 23364 16939 23420 16941
rect 23364 16887 23366 16939
rect 23366 16887 23418 16939
rect 23418 16887 23420 16939
rect 23364 16885 23420 16887
rect 23214 15609 23270 15611
rect 23214 15557 23216 15609
rect 23216 15557 23268 15609
rect 23268 15557 23270 15609
rect 23214 15555 23270 15557
rect 23400 15609 23456 15611
rect 23400 15557 23402 15609
rect 23402 15557 23454 15609
rect 23454 15557 23456 15609
rect 23400 15555 23456 15557
rect 23162 15015 23218 15017
rect 23162 14963 23164 15015
rect 23164 14963 23216 15015
rect 23216 14963 23218 15015
rect 23162 14961 23218 14963
rect 23162 14829 23218 14831
rect 23162 14777 23164 14829
rect 23164 14777 23216 14829
rect 23216 14777 23218 14829
rect 23162 14775 23218 14777
rect 23610 15015 23666 15017
rect 23610 14963 23612 15015
rect 23612 14963 23664 15015
rect 23664 14963 23666 15015
rect 23610 14961 23666 14963
rect 23610 14829 23666 14831
rect 23610 14777 23612 14829
rect 23612 14777 23664 14829
rect 23664 14777 23666 14829
rect 23610 14775 23666 14777
rect 23167 12576 23223 12578
rect 23167 12524 23169 12576
rect 23169 12524 23221 12576
rect 23221 12524 23223 12576
rect 23167 12522 23223 12524
rect 23167 12390 23223 12392
rect 23167 12338 23169 12390
rect 23169 12338 23221 12390
rect 23221 12338 23223 12390
rect 23167 12336 23223 12338
rect 23608 12576 23664 12578
rect 23608 12524 23610 12576
rect 23610 12524 23662 12576
rect 23662 12524 23664 12576
rect 23608 12522 23664 12524
rect 23608 12390 23664 12392
rect 23608 12338 23610 12390
rect 23610 12338 23662 12390
rect 23662 12338 23664 12390
rect 23608 12336 23664 12338
rect 23167 12038 23223 12040
rect 23167 11986 23169 12038
rect 23169 11986 23221 12038
rect 23221 11986 23223 12038
rect 23167 11984 23223 11986
rect 23167 11852 23223 11854
rect 23167 11800 23169 11852
rect 23169 11800 23221 11852
rect 23221 11800 23223 11852
rect 23167 11798 23223 11800
rect 23608 12038 23664 12040
rect 23608 11986 23610 12038
rect 23610 11986 23662 12038
rect 23662 11986 23664 12038
rect 23608 11984 23664 11986
rect 23608 11852 23664 11854
rect 23608 11800 23610 11852
rect 23610 11800 23662 11852
rect 23662 11800 23664 11852
rect 23608 11798 23664 11800
rect 23167 11433 23223 11435
rect 23167 11381 23169 11433
rect 23169 11381 23221 11433
rect 23221 11381 23223 11433
rect 23167 11379 23223 11381
rect 23167 11247 23223 11249
rect 23167 11195 23169 11247
rect 23169 11195 23221 11247
rect 23221 11195 23223 11247
rect 23167 11193 23223 11195
rect 23608 11433 23664 11435
rect 23608 11381 23610 11433
rect 23610 11381 23662 11433
rect 23662 11381 23664 11433
rect 23608 11379 23664 11381
rect 23608 11247 23664 11249
rect 23608 11195 23610 11247
rect 23610 11195 23662 11247
rect 23662 11195 23664 11247
rect 23608 11193 23664 11195
rect 23171 7774 23227 7776
rect 23171 7722 23173 7774
rect 23173 7722 23225 7774
rect 23225 7722 23227 7774
rect 23171 7720 23227 7722
rect 23171 7588 23227 7590
rect 23171 7536 23173 7588
rect 23173 7536 23225 7588
rect 23225 7536 23227 7588
rect 23171 7534 23227 7536
rect 23171 7402 23227 7404
rect 23171 7350 23173 7402
rect 23173 7350 23225 7402
rect 23225 7350 23227 7402
rect 23171 7348 23227 7350
rect 23613 7774 23669 7776
rect 23613 7722 23615 7774
rect 23615 7722 23667 7774
rect 23667 7722 23669 7774
rect 23613 7720 23669 7722
rect 23613 7588 23669 7590
rect 23613 7536 23615 7588
rect 23615 7536 23667 7588
rect 23667 7536 23669 7588
rect 23613 7534 23669 7536
rect 23613 7402 23669 7404
rect 23613 7350 23615 7402
rect 23615 7350 23667 7402
rect 23667 7350 23669 7402
rect 23613 7348 23669 7350
rect 23295 4973 23351 4975
rect 23295 4921 23297 4973
rect 23297 4921 23349 4973
rect 23349 4921 23351 4973
rect 23295 4919 23351 4921
rect 23507 4973 23563 4975
rect 23507 4921 23509 4973
rect 23509 4921 23561 4973
rect 23561 4921 23563 4973
rect 23507 4919 23563 4921
rect 23295 4755 23351 4757
rect 23295 4703 23297 4755
rect 23297 4703 23349 4755
rect 23349 4703 23351 4755
rect 23295 4701 23351 4703
rect 23507 4755 23563 4757
rect 23507 4703 23509 4755
rect 23509 4703 23561 4755
rect 23561 4703 23563 4755
rect 23507 4701 23563 4703
<< metal3 >>
rect -1 39107 23681 39307
rect -1 30537 23681 30897
rect 38 30341 128 30351
rect 38 30077 62 30341
rect 118 30279 128 30341
rect 118 30139 23681 30279
rect 118 30077 128 30139
rect 38 30067 128 30077
rect 800 29987 24087 29997
rect 800 29943 996 29987
rect -1 29931 996 29943
rect 1052 29931 11798 29987
rect 11854 29931 22958 29987
rect 23014 29931 24087 29987
rect -1 29855 24087 29931
rect -1 29799 996 29855
rect 1052 29799 11798 29855
rect 11854 29799 22958 29855
rect 23014 29799 24087 29855
rect -1 29723 24087 29799
rect -1 29667 996 29723
rect 1052 29667 11798 29723
rect 11854 29667 22958 29723
rect 23014 29667 24087 29723
rect -1 29591 24087 29667
rect -1 29535 996 29591
rect 1052 29535 11798 29591
rect 11854 29535 22958 29591
rect 23014 29535 24087 29591
rect -1 29517 24087 29535
rect -1 29471 1243 29517
rect 22636 29105 24206 29106
rect 800 29071 24206 29105
rect 800 29015 1358 29071
rect 1414 29015 12158 29071
rect 12214 29015 22598 29071
rect 22654 29015 24206 29071
rect 800 28964 24206 29015
rect 800 28939 23367 28964
rect 800 28883 1358 28939
rect 1414 28883 12158 28939
rect 12214 28883 22598 28939
rect 22654 28908 23367 28939
rect 23423 28908 24206 28964
rect 22654 28883 24206 28908
rect 800 28807 24206 28883
rect 800 28751 1358 28807
rect 1414 28751 12158 28807
rect 12214 28751 22598 28807
rect 22654 28778 24206 28807
rect 22654 28751 23367 28778
rect 800 28722 23367 28751
rect 23423 28722 24206 28778
rect 800 28675 24206 28722
rect 800 28619 1358 28675
rect 1414 28619 12158 28675
rect 12214 28619 22598 28675
rect 22654 28619 24206 28675
rect 800 28543 24206 28619
rect 800 28487 1358 28543
rect 1414 28487 12158 28543
rect 12214 28487 22598 28543
rect 22654 28487 24206 28543
rect 800 28411 24206 28487
rect 800 28355 1358 28411
rect 1414 28355 12158 28411
rect 12214 28355 22598 28411
rect 22654 28355 24206 28411
rect 800 28279 24206 28355
rect 800 28223 1358 28279
rect 1414 28223 12158 28279
rect 12214 28223 22598 28279
rect 22654 28223 24206 28279
rect 800 28147 24206 28223
rect 800 28091 1358 28147
rect 1414 28091 12158 28147
rect 12214 28091 22598 28147
rect 22654 28091 24206 28147
rect 800 28015 24206 28091
rect 800 27959 1358 28015
rect 1414 27959 12158 28015
rect 12214 27959 22598 28015
rect 22654 27959 24206 28015
rect 800 27883 24206 27959
rect 800 27827 1358 27883
rect 1414 27827 12158 27883
rect 12214 27827 22598 27883
rect 22654 27827 24206 27883
rect 800 27751 24206 27827
rect 800 27695 1358 27751
rect 1414 27695 12158 27751
rect 12214 27695 22598 27751
rect 22654 27695 24206 27751
rect 800 27619 24206 27695
rect 800 27563 1358 27619
rect 1414 27563 12158 27619
rect 12214 27563 22598 27619
rect 22654 27563 24206 27619
rect 800 27297 24206 27563
rect 800 27296 24087 27297
rect 22691 22026 24206 23296
rect 22691 21970 23534 22026
rect 23590 21970 24206 22026
rect 22691 21808 24206 21970
rect 22691 21752 23534 21808
rect 23590 21752 24206 21808
rect 22691 21415 24206 21752
rect 22586 21304 24206 21305
rect 1314 21090 24206 21304
rect 1314 21089 23252 21090
rect 22586 20983 24206 20984
rect 1314 20768 24206 20983
rect 1314 20767 23252 20768
rect 22586 20661 24206 20662
rect 1314 20447 24206 20661
rect 1314 20446 23252 20447
rect 22586 20339 24206 20340
rect 1314 20125 24206 20339
rect 1314 20124 23252 20125
rect 1314 19433 23939 19648
rect 1314 19432 23252 19433
rect 1314 19111 23939 19326
rect 1314 19110 23252 19111
rect 1314 18789 23939 19004
rect 22586 18682 23939 18683
rect 1314 18467 23939 18682
rect 1314 18185 24206 18361
rect 1314 18129 23137 18185
rect 23193 18129 23317 18185
rect 23373 18129 24206 18185
rect 1314 17919 24206 18129
rect 1314 17918 23252 17919
rect 1314 16941 24206 17263
rect 1314 16885 23364 16941
rect 23420 16885 24206 16941
rect 1314 16808 24206 16885
rect 1314 16807 23252 16808
rect 1314 15611 23710 15720
rect 1314 15555 23214 15611
rect 23270 15555 23400 15611
rect 23456 15555 23710 15611
rect 1314 15017 23710 15555
rect 1314 14961 23162 15017
rect 23218 14961 23610 15017
rect 23666 14961 23710 15017
rect 1314 14831 23710 14961
rect 1314 14775 23162 14831
rect 23218 14775 23610 14831
rect 23666 14775 23710 14831
rect 1314 12997 23710 14775
rect 1314 12996 23252 12997
rect 1314 12578 23710 12711
rect 1314 12522 23167 12578
rect 23223 12522 23608 12578
rect 23664 12522 23710 12578
rect 1314 12392 23710 12522
rect 1314 12336 23167 12392
rect 23223 12336 23608 12392
rect 23664 12336 23710 12392
rect 1314 12040 23710 12336
rect 1314 11984 23167 12040
rect 23223 11984 23608 12040
rect 23664 11984 23710 12040
rect 1314 11854 23710 11984
rect 1314 11798 23167 11854
rect 23223 11798 23608 11854
rect 23664 11798 23710 11854
rect 1314 11435 23710 11798
rect 1314 11379 23167 11435
rect 23223 11379 23608 11435
rect 23664 11379 23710 11435
rect 1314 11249 23710 11379
rect 1314 11193 23167 11249
rect 23223 11193 23608 11249
rect 23664 11193 23710 11249
rect 1314 9309 23710 11193
rect 1314 9308 23252 9309
rect 22658 9158 23710 9160
rect 1262 8442 23710 9158
rect 22658 7827 23710 7828
rect 1262 7776 24488 7827
rect 1262 7720 23171 7776
rect 23227 7720 23613 7776
rect 23669 7720 24488 7776
rect 1262 7590 24488 7720
rect 1262 7534 23171 7590
rect 23227 7534 23613 7590
rect 23669 7534 24488 7590
rect 1262 7404 24488 7534
rect 1262 7348 23171 7404
rect 23227 7348 23613 7404
rect 23669 7348 24488 7404
rect 1262 7016 24488 7348
rect 1314 5154 23971 6474
rect 1165 4929 22567 5005
rect 23259 4975 23599 5014
rect 23259 4919 23295 4975
rect 23351 4919 23507 4975
rect 23563 4919 23599 4975
rect 23259 4758 23599 4919
rect 1165 4757 23599 4758
rect 1165 4701 23295 4757
rect 23351 4701 23507 4757
rect 23563 4701 23599 4757
rect 1165 4662 23599 4701
rect 1314 3133 24166 4495
rect 1314 1961 24276 2576
rect 1314 1286 23252 1855
rect 1314 747 24089 1179
rect 1314 155 24508 610
rect 1277 -959 24602 -504
rect 1277 -1599 23252 -1247
rect 1277 -2041 23252 -1953
rect 1277 -2517 23252 -2165
rect 1277 -3242 23252 -2787
use col_64a_64x8m81  col_64a_64x8m81_0
timestamp 1698431365
transform 1 0 907 0 1 31107
box -1997 -68 23144 7268
use dcap_103_novia_64x8m81  dcap_103_novia_64x8m81_0
array 0 35 619 0 0 0
timestamp 1698431365
transform 1 0 288 0 1 29009
box 0 0 1 1
use M2_M1$$43374636_64x8m81  M2_M1$$43374636_64x8m81_0
timestamp 1698431365
transform 1 0 23429 0 1 4838
box 0 0 1 1
use M2_M1431058998320_64x8m81  M2_M1431058998320_64x8m81_0
timestamp 1698431365
transform -1 0 11867 0 -1 29852
box 0 0 1 1
use M2_M1431058998320_64x8m81  M2_M1431058998320_64x8m81_1
timestamp 1698431365
transform -1 0 1026 0 -1 29852
box 0 0 1 1
use M2_M14310589983225_64x8m81  M2_M14310589983225_64x8m81_0
timestamp 1698431365
transform -1 0 22888 0 -1 29897
box 0 0 1 1
use M3_M2$$201416748_64x8m81  M3_M2$$201416748_64x8m81_0
timestamp 1698431365
transform 1 0 23429 0 1 4838
box 0 0 1 1
use M3_M24310589983226_64x8m81  M3_M24310589983226_64x8m81_0
timestamp 1698431365
transform 1 0 1024 0 1 29761
box 0 0 1 1
use M3_M24310589983226_64x8m81  M3_M24310589983226_64x8m81_1
timestamp 1698431365
transform 1 0 11826 0 1 29761
box 0 0 1 1
use M3_M24310589983226_64x8m81  M3_M24310589983226_64x8m81_2
timestamp 1698431365
transform 1 0 22986 0 1 29761
box 0 0 1 1
use M3_M24310589983227_64x8m81  M3_M24310589983227_64x8m81_0
timestamp 1698431365
transform 1 0 12186 0 1 28317
box 0 0 1 1
use M3_M24310589983227_64x8m81  M3_M24310589983227_64x8m81_1
timestamp 1698431365
transform 1 0 22626 0 1 28317
box 0 0 1 1
use M3_M24310589983227_64x8m81  M3_M24310589983227_64x8m81_2
timestamp 1698431365
transform 1 0 1386 0 1 28317
box 0 0 1 1
use rdummy_64x4_64x8m81  rdummy_64x4_64x8m81_0
timestamp 1698431365
transform 1 0 307 0 1 30207
box -217 -22942 23616 9068
use saout_m2_64x8m81  saout_m2_64x8m81_0
timestamp 1698431365
transform 1 0 11820 0 1 -1
box -269 -3393 7633 31140
use saout_m2_64x8m81  saout_m2_64x8m81_1
timestamp 1698431365
transform 1 0 1020 0 1 -1
box -269 -3393 7633 31140
use saout_R_m2_64x8m81  saout_R_m2_64x8m81_0
timestamp 1698431365
transform -1 0 12194 0 1 6
box -269 -3400 7633 31133
use saout_R_m2_64x8m81  saout_R_m2_64x8m81_1
timestamp 1698431365
transform -1 0 22994 0 1 6
box -269 -3400 7633 31133
<< labels >>
rlabel metal1 s 7342 15928 7342 15928 4 pcb[6]
port 1 nsew
rlabel metal1 s 5921 15928 5921 15928 4 pcb[7]
port 2 nsew
rlabel metal1 s 18209 15928 18209 15928 4 pcb[4]
port 3 nsew
rlabel metal1 s 1827 18163 1827 18163 4 vdd
port 4 nsew
flabel metal1 s 22465 -3332 22465 -3332 0 FreeSans 600 0 0 0 WEN[4]
port 5 nsew
flabel metal1 s 1584 -3332 1584 -3332 0 FreeSans 600 0 0 0 WEN[7]
port 6 nsew
rlabel metal1 s 16588 15928 16588 15928 4 pcb[5]
port 7 nsew
flabel metal1 s 12358 -3332 12358 -3332 0 FreeSans 600 0 0 0 WEN[5]
port 8 nsew
flabel metal1 s 11643 -3332 11643 -3332 0 FreeSans 600 0 0 0 WEN[6]
port 9 nsew
rlabel metal3 s 1607 36968 1607 36968 4 WL[6]
port 10 nsew
rlabel metal3 s 1607 36068 1607 36068 4 WL[5]
port 11 nsew
rlabel metal3 s 1777 1467 1777 1467 4 men
port 12 nsew
rlabel metal3 s 1704 18914 1704 18914 4 ypass[1]
port 13 nsew
rlabel metal3 s 1704 19231 1704 19231 4 ypass[2]
port 14 nsew
rlabel metal3 s 1704 19548 1704 19548 4 ypass[3]
port 15 nsew
rlabel metal3 s 1704 20204 1704 20204 4 ypass[4]
port 16 nsew
rlabel metal3 s 1704 20528 1704 20528 4 ypass[5]
port 17 nsew
rlabel metal3 s 1704 20845 1704 20845 4 ypass[6]
port 18 nsew
rlabel metal3 s 1774 1467 1774 1467 4 men
port 12 nsew
rlabel metal3 s 1592 38757 1592 38757 4 DWL
port 19 nsew
rlabel metal3 s 1346 4726 1346 4726 4 tblhl
port 20 nsew
flabel metal3 s 1659 -2004 1659 -2004 0 FreeSans 1000 0 0 0 GWEN
port 21 nsew
flabel metal3 s 1659 -3019 1659 -3019 0 FreeSans 448 0 0 0 VDD
port 22 nsew
rlabel metal3 s 1777 8832 1777 8832 4 VDD
port 22 nsew
rlabel metal3 s 1777 5806 1777 5806 4 VSS
port 23 nsew
flabel metal3 s 1659 -781 1659 -781 0 FreeSans 448 0 0 0 VDD
port 22 nsew
flabel metal3 s 1659 -2347 1659 -2347 0 FreeSans 448 0 0 0 VSS
port 23 nsew
rlabel metal3 s 240 30277 240 30277 4 VSS
port 23 nsew
rlabel metal3 s 1777 39217 1777 39217 4 VSS
port 23 nsew
rlabel metal3 s 1777 1466 1777 1466 4 men
port 12 nsew
rlabel metal3 s 1704 18591 1704 18591 4 ypass[0]
port 24 nsew
rlabel metal3 s 1775 1466 1775 1466 4 men
port 12 nsew
rlabel metal3 s 1346 4983 1346 4983 4 GWE
port 25 nsew
rlabel metal3 s 1608 31568 1608 31568 4 WL[0]
port 26 nsew
rlabel metal3 s 1608 33368 1608 33368 4 WL[2]
port 27 nsew
rlabel metal3 s 1608 34268 1608 34268 4 WL[3]
port 28 nsew
rlabel metal3 s 1608 35168 1608 35168 4 WL[4]
port 29 nsew
rlabel metal3 s 1608 37868 1608 37868 4 WL[7]
port 30 nsew
rlabel metal3 s 1608 32468 1608 32468 4 WL[1]
port 31 nsew
rlabel metal3 s 1705 21162 1705 21162 4 ypass[7]
port 32 nsew
rlabel metal3 s 1777 1466 1777 1466 4 men
port 12 nsew
rlabel metal3 s 1775 1466 1775 1466 4 men
port 12 nsew
flabel metal3 s 1659 -1446 1659 -1446 0 FreeSans 448 0 0 0 VSS
port 23 nsew
flabel metal3 s 1659 390 1659 390 0 FreeSans 448 0 0 0 VDD
port 22 nsew
flabel metal3 s 1659 3623 1659 3623 0 FreeSans 448 0 0 0 VDD
port 22 nsew
flabel metal3 s 1659 7598 1659 7598 0 FreeSans 448 0 0 0 VDD
port 22 nsew
flabel metal3 s 1659 14001 1659 14001 0 FreeSans 448 0 0 0 VDD
port 22 nsew
flabel metal3 s 1659 18106 1659 18106 0 FreeSans 448 0 0 0 VDD
port 22 nsew
flabel metal3 s 1659 28191 1659 28191 0 FreeSans 448 0 0 0 VDD
port 22 nsew
flabel metal3 s 315 29699 315 29699 0 FreeSans 448 0 0 0 VSS
port 23 nsew
flabel metal3 s 1659 23123 1659 23123 0 FreeSans 448 0 0 0 VSS
port 23 nsew
flabel metal3 s 1659 16976 1659 16976 0 FreeSans 448 0 0 0 VSS
port 23 nsew
flabel metal3 s 1659 12236 1659 12236 0 FreeSans 448 0 0 0 VSS
port 23 nsew
flabel metal3 s 1659 6155 1659 6155 0 FreeSans 448 0 0 0 VSS
port 23 nsew
flabel metal3 s 1659 2247 1659 2247 0 FreeSans 448 0 0 0 VSS
port 23 nsew
flabel metal3 s 1659 949 1659 949 0 FreeSans 448 0 0 0 VSS
port 23 nsew
rlabel metal2 s 1523 104 1523 104 4 din[4]
port 33 nsew
rlabel metal2 s 22489 104 22489 104 4 din[7]
port 34 nsew
rlabel metal2 s 10837 138 10837 138 4 q[5]
port 35 nsew
rlabel metal2 s 13166 104 13166 104 4 q[6]
port 36 nsew
rlabel metal2 s 21642 104 21642 104 4 q[7]
port 37 nsew
rlabel metal2 s 11684 104 11684 104 4 din[5]
port 38 nsew
rlabel metal2 s 12319 104 12319 104 4 din[6]
port 39 nsew
rlabel metal2 s 2377 104 2377 104 4 q[4]
port 40 nsew
<< properties >>
string GDS_END 2231102
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 2220982
<< end >>
