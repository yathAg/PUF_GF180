magic
tech gf180mcuA
magscale 1 10
timestamp 1698431365
<< metal3 >>
rect -1997 57030 22836 57390
rect -1997 56010 22836 56370
rect -1997 55230 22836 55590
rect -1997 54210 22836 54570
rect -1997 53430 22836 53790
rect -1997 52410 22836 52770
rect -1997 51630 22836 51990
rect -1997 50610 22836 50970
rect -1997 49830 22836 50190
rect -1997 48810 22836 49170
rect -1997 48030 22836 48390
rect -1997 47010 22836 47370
rect -1997 46230 22836 46590
rect -1997 45210 22836 45570
rect -1997 44430 22836 44790
rect -1997 43410 22836 43770
rect -1997 42630 22836 42990
rect -1997 41610 22836 41970
rect -1997 40830 22836 41190
rect -1997 39810 22836 40170
rect -1997 39030 22836 39390
rect -1997 38010 22836 38370
rect -1997 37230 22836 37590
rect -1997 36210 22836 36570
rect -1997 35430 22836 35790
rect -1997 34410 22836 34770
rect -1997 33630 22836 33990
rect -1997 32610 22836 32970
rect -1997 31830 22836 32190
rect -1997 30810 22836 31170
rect -1997 30030 22836 30390
rect -1997 29010 22836 29370
rect -1997 28230 22836 28590
rect -1997 27210 22836 27570
rect -1997 26430 22836 26790
rect -1997 25410 22836 25770
rect -1997 24630 22836 24990
rect -1997 23610 22836 23970
rect -1997 22830 22836 23190
rect -1997 21810 22836 22170
rect -1997 21030 22836 21390
rect -1997 20010 22836 20370
rect -1997 19230 22836 19590
rect -1997 18210 22836 18570
rect -1997 17430 22836 17790
rect -1997 16410 22836 16770
rect -1997 15630 22836 15990
rect -1997 14610 22836 14970
rect -1997 13830 22836 14190
rect -1997 12810 22836 13170
rect -1997 12030 22836 12390
rect -1997 11010 22836 11370
rect -1997 10230 22836 10590
rect -1997 9210 22836 9570
rect -1997 8430 22836 8790
rect -1997 7410 22836 7770
rect -1997 6630 22836 6990
rect -1997 5610 22836 5970
rect -1997 4830 22836 5190
rect -1997 3810 22836 4170
rect -1997 3030 22836 3390
rect -1997 2010 22836 2370
rect -1997 1230 22836 1590
rect -1997 210 22836 570
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_0
timestamp 1698431365
transform -1 0 18000 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1
timestamp 1698431365
transform -1 0 18000 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_2
timestamp 1698431365
transform -1 0 18000 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_3
timestamp 1698431365
transform -1 0 17400 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_4
timestamp 1698431365
transform -1 0 17400 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_5
timestamp 1698431365
transform -1 0 17400 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_6
timestamp 1698431365
transform -1 0 18000 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_7
timestamp 1698431365
transform -1 0 17400 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_8
timestamp 1698431365
transform -1 0 21600 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_9
timestamp 1698431365
transform -1 0 17400 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_10
timestamp 1698431365
transform -1 0 21600 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_11
timestamp 1698431365
transform -1 0 21600 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_12
timestamp 1698431365
transform -1 0 21600 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_13
timestamp 1698431365
transform -1 0 21600 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_14
timestamp 1698431365
transform -1 0 21600 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_15
timestamp 1698431365
transform -1 0 21600 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_16
timestamp 1698431365
transform -1 0 18600 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_17
timestamp 1698431365
transform -1 0 19200 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_18
timestamp 1698431365
transform -1 0 19200 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_19
timestamp 1698431365
transform -1 0 19200 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_20
timestamp 1698431365
transform -1 0 19200 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_21
timestamp 1698431365
transform -1 0 19200 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_22
timestamp 1698431365
transform -1 0 19200 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_23
timestamp 1698431365
transform -1 0 19200 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_24
timestamp 1698431365
transform -1 0 18600 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_25
timestamp 1698431365
transform -1 0 18000 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_26
timestamp 1698431365
transform -1 0 18600 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_27
timestamp 1698431365
transform -1 0 18000 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_28
timestamp 1698431365
transform -1 0 18600 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_29
timestamp 1698431365
transform -1 0 18600 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_30
timestamp 1698431365
transform -1 0 17400 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_31
timestamp 1698431365
transform -1 0 17400 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_32
timestamp 1698431365
transform -1 0 18600 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_33
timestamp 1698431365
transform -1 0 18600 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_34
timestamp 1698431365
transform -1 0 20400 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_35
timestamp 1698431365
transform -1 0 20400 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_36
timestamp 1698431365
transform -1 0 19800 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_37
timestamp 1698431365
transform -1 0 19800 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_38
timestamp 1698431365
transform -1 0 19800 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_39
timestamp 1698431365
transform -1 0 19800 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_40
timestamp 1698431365
transform -1 0 21000 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_41
timestamp 1698431365
transform -1 0 21000 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_42
timestamp 1698431365
transform -1 0 21000 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_43
timestamp 1698431365
transform -1 0 21000 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_44
timestamp 1698431365
transform -1 0 21000 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_45
timestamp 1698431365
transform -1 0 21000 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_46
timestamp 1698431365
transform -1 0 21000 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_47
timestamp 1698431365
transform -1 0 19800 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_48
timestamp 1698431365
transform -1 0 19800 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_49
timestamp 1698431365
transform -1 0 19800 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_50
timestamp 1698431365
transform -1 0 18000 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_51
timestamp 1698431365
transform -1 0 20400 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_52
timestamp 1698431365
transform -1 0 20400 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_53
timestamp 1698431365
transform -1 0 20400 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_54
timestamp 1698431365
transform -1 0 20400 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_55
timestamp 1698431365
transform -1 0 20400 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_56
timestamp 1698431365
transform 1 0 11400 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_57
timestamp 1698431365
transform 1 0 11400 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_58
timestamp 1698431365
transform 1 0 11400 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_59
timestamp 1698431365
transform 1 0 11400 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_60
timestamp 1698431365
transform 1 0 11400 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_61
timestamp 1698431365
transform 1 0 11400 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_62
timestamp 1698431365
transform 1 0 11400 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_63
timestamp 1698431365
transform 1 0 12000 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_64
timestamp 1698431365
transform 1 0 12000 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_65
timestamp 1698431365
transform 1 0 12000 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_66
timestamp 1698431365
transform 1 0 15000 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_67
timestamp 1698431365
transform 1 0 14400 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_68
timestamp 1698431365
transform 1 0 15000 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_69
timestamp 1698431365
transform 1 0 15000 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_70
timestamp 1698431365
transform 1 0 15000 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_71
timestamp 1698431365
transform 1 0 15000 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_72
timestamp 1698431365
transform 1 0 12600 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_73
timestamp 1698431365
transform 1 0 12600 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_74
timestamp 1698431365
transform 1 0 12600 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_75
timestamp 1698431365
transform 1 0 12600 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_76
timestamp 1698431365
transform 1 0 14400 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_77
timestamp 1698431365
transform 1 0 14400 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_78
timestamp 1698431365
transform 1 0 14400 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_79
timestamp 1698431365
transform 1 0 14400 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_80
timestamp 1698431365
transform 1 0 14400 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_81
timestamp 1698431365
transform 1 0 14400 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_82
timestamp 1698431365
transform 1 0 12600 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_83
timestamp 1698431365
transform 1 0 15000 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_84
timestamp 1698431365
transform 1 0 13800 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_85
timestamp 1698431365
transform 1 0 13800 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_86
timestamp 1698431365
transform 1 0 13800 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_87
timestamp 1698431365
transform 1 0 13800 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_88
timestamp 1698431365
transform 1 0 13800 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_89
timestamp 1698431365
transform 1 0 15000 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_90
timestamp 1698431365
transform 1 0 15600 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_91
timestamp 1698431365
transform 1 0 15600 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_92
timestamp 1698431365
transform 1 0 15600 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_93
timestamp 1698431365
transform 1 0 15600 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_94
timestamp 1698431365
transform 1 0 15600 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_95
timestamp 1698431365
transform 1 0 15600 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_96
timestamp 1698431365
transform 1 0 15600 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_97
timestamp 1698431365
transform 1 0 13800 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_98
timestamp 1698431365
transform 1 0 13800 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_99
timestamp 1698431365
transform 1 0 13200 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_100
timestamp 1698431365
transform 1 0 13200 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_101
timestamp 1698431365
transform 1 0 13200 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_102
timestamp 1698431365
transform 1 0 13200 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_103
timestamp 1698431365
transform 1 0 13200 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_104
timestamp 1698431365
transform 1 0 13200 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_105
timestamp 1698431365
transform 1 0 13200 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_106
timestamp 1698431365
transform 1 0 12000 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_107
timestamp 1698431365
transform 1 0 12000 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_108
timestamp 1698431365
transform 1 0 12000 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_109
timestamp 1698431365
transform 1 0 12000 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_110
timestamp 1698431365
transform 1 0 12600 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_111
timestamp 1698431365
transform 1 0 12600 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_112
timestamp 1698431365
transform 1 0 15600 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_113
timestamp 1698431365
transform 1 0 11400 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_114
timestamp 1698431365
transform 1 0 15600 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_115
timestamp 1698431365
transform 1 0 15600 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_116
timestamp 1698431365
transform 1 0 15600 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_117
timestamp 1698431365
transform 1 0 13200 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_118
timestamp 1698431365
transform 1 0 15600 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_119
timestamp 1698431365
transform 1 0 13200 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_120
timestamp 1698431365
transform 1 0 11400 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_121
timestamp 1698431365
transform 1 0 11400 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_122
timestamp 1698431365
transform 1 0 13200 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_123
timestamp 1698431365
transform 1 0 15000 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_124
timestamp 1698431365
transform 1 0 15000 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_125
timestamp 1698431365
transform 1 0 13200 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_126
timestamp 1698431365
transform 1 0 13200 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_127
timestamp 1698431365
transform 1 0 12000 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_128
timestamp 1698431365
transform 1 0 12000 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_129
timestamp 1698431365
transform 1 0 15000 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_130
timestamp 1698431365
transform 1 0 15000 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_131
timestamp 1698431365
transform 1 0 15000 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_132
timestamp 1698431365
transform 1 0 15000 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_133
timestamp 1698431365
transform 1 0 13200 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_134
timestamp 1698431365
transform 1 0 15600 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_135
timestamp 1698431365
transform 1 0 12000 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_136
timestamp 1698431365
transform 1 0 12600 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_137
timestamp 1698431365
transform 1 0 14400 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_138
timestamp 1698431365
transform 1 0 14400 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_139
timestamp 1698431365
transform 1 0 14400 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_140
timestamp 1698431365
transform 1 0 14400 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_141
timestamp 1698431365
transform 1 0 14400 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_142
timestamp 1698431365
transform 1 0 14400 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_143
timestamp 1698431365
transform 1 0 11400 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_144
timestamp 1698431365
transform 1 0 11400 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_145
timestamp 1698431365
transform 1 0 12600 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_146
timestamp 1698431365
transform 1 0 12600 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_147
timestamp 1698431365
transform 1 0 12600 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_148
timestamp 1698431365
transform 1 0 12600 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_149
timestamp 1698431365
transform 1 0 12600 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_150
timestamp 1698431365
transform 1 0 13800 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_151
timestamp 1698431365
transform 1 0 13800 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_152
timestamp 1698431365
transform 1 0 13800 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_153
timestamp 1698431365
transform 1 0 13800 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_154
timestamp 1698431365
transform 1 0 13800 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_155
timestamp 1698431365
transform 1 0 13800 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_156
timestamp 1698431365
transform 1 0 12000 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_157
timestamp 1698431365
transform 1 0 12000 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_158
timestamp 1698431365
transform 1 0 12000 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_159
timestamp 1698431365
transform 1 0 11400 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_160
timestamp 1698431365
transform -1 0 18000 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_161
timestamp 1698431365
transform -1 0 20400 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_162
timestamp 1698431365
transform -1 0 18000 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_163
timestamp 1698431365
transform -1 0 18000 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_164
timestamp 1698431365
transform -1 0 18000 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_165
timestamp 1698431365
transform -1 0 18000 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_166
timestamp 1698431365
transform -1 0 18000 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_167
timestamp 1698431365
transform -1 0 20400 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_168
timestamp 1698431365
transform -1 0 19800 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_169
timestamp 1698431365
transform -1 0 19800 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_170
timestamp 1698431365
transform -1 0 18600 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_171
timestamp 1698431365
transform -1 0 17400 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_172
timestamp 1698431365
transform -1 0 17400 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_173
timestamp 1698431365
transform -1 0 17400 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_174
timestamp 1698431365
transform -1 0 17400 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_175
timestamp 1698431365
transform -1 0 17400 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_176
timestamp 1698431365
transform -1 0 17400 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_177
timestamp 1698431365
transform -1 0 18600 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_178
timestamp 1698431365
transform -1 0 18600 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_179
timestamp 1698431365
transform -1 0 18600 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_180
timestamp 1698431365
transform -1 0 18600 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_181
timestamp 1698431365
transform -1 0 18600 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_182
timestamp 1698431365
transform -1 0 19800 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_183
timestamp 1698431365
transform -1 0 21600 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_184
timestamp 1698431365
transform -1 0 21600 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_185
timestamp 1698431365
transform -1 0 21600 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_186
timestamp 1698431365
transform -1 0 21600 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_187
timestamp 1698431365
transform -1 0 21600 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_188
timestamp 1698431365
transform -1 0 21600 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_189
timestamp 1698431365
transform -1 0 19800 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_190
timestamp 1698431365
transform -1 0 19800 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_191
timestamp 1698431365
transform -1 0 19800 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_192
timestamp 1698431365
transform -1 0 20400 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_193
timestamp 1698431365
transform -1 0 21000 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_194
timestamp 1698431365
transform -1 0 21000 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_195
timestamp 1698431365
transform -1 0 21000 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_196
timestamp 1698431365
transform -1 0 21000 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_197
timestamp 1698431365
transform -1 0 21000 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_198
timestamp 1698431365
transform -1 0 21000 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_199
timestamp 1698431365
transform -1 0 20400 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_200
timestamp 1698431365
transform -1 0 20400 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_201
timestamp 1698431365
transform -1 0 20400 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_202
timestamp 1698431365
transform -1 0 19200 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_203
timestamp 1698431365
transform -1 0 19200 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_204
timestamp 1698431365
transform -1 0 19200 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_205
timestamp 1698431365
transform -1 0 19200 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_206
timestamp 1698431365
transform -1 0 19200 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_207
timestamp 1698431365
transform -1 0 19200 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_208
timestamp 1698431365
transform -1 0 18000 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_209
timestamp 1698431365
transform -1 0 18000 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_210
timestamp 1698431365
transform -1 0 17400 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_211
timestamp 1698431365
transform -1 0 17400 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_212
timestamp 1698431365
transform 1 0 13800 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_213
timestamp 1698431365
transform 1 0 13800 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_214
timestamp 1698431365
transform 1 0 11400 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_215
timestamp 1698431365
transform 1 0 11400 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_216
timestamp 1698431365
transform -1 0 21600 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_217
timestamp 1698431365
transform -1 0 21600 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_218
timestamp 1698431365
transform 1 0 14400 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_219
timestamp 1698431365
transform 1 0 14400 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_220
timestamp 1698431365
transform -1 0 21000 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_221
timestamp 1698431365
transform -1 0 21000 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_222
timestamp 1698431365
transform -1 0 19200 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_223
timestamp 1698431365
transform -1 0 19200 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_224
timestamp 1698431365
transform 1 0 12600 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_225
timestamp 1698431365
transform 1 0 12600 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_226
timestamp 1698431365
transform -1 0 18600 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_227
timestamp 1698431365
transform -1 0 18600 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_228
timestamp 1698431365
transform 1 0 15000 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_229
timestamp 1698431365
transform 1 0 15000 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_230
timestamp 1698431365
transform -1 0 20400 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_231
timestamp 1698431365
transform -1 0 20400 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_232
timestamp 1698431365
transform 1 0 12000 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_233
timestamp 1698431365
transform 1 0 12000 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_234
timestamp 1698431365
transform -1 0 19800 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_235
timestamp 1698431365
transform -1 0 19800 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_236
timestamp 1698431365
transform 1 0 13200 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_237
timestamp 1698431365
transform 1 0 13200 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_238
timestamp 1698431365
transform 1 0 15600 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_239
timestamp 1698431365
transform 1 0 15600 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_240
timestamp 1698431365
transform -1 0 9600 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_241
timestamp 1698431365
transform -1 0 9600 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_242
timestamp 1698431365
transform -1 0 9600 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_243
timestamp 1698431365
transform -1 0 9600 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_244
timestamp 1698431365
transform -1 0 9600 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_245
timestamp 1698431365
transform -1 0 9600 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_246
timestamp 1698431365
transform -1 0 9600 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_247
timestamp 1698431365
transform -1 0 10800 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_248
timestamp 1698431365
transform -1 0 10800 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_249
timestamp 1698431365
transform -1 0 10800 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_250
timestamp 1698431365
transform -1 0 7800 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_251
timestamp 1698431365
transform -1 0 7800 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_252
timestamp 1698431365
transform -1 0 7800 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_253
timestamp 1698431365
transform -1 0 7800 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_254
timestamp 1698431365
transform -1 0 7800 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_255
timestamp 1698431365
transform -1 0 7800 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_256
timestamp 1698431365
transform -1 0 7800 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_257
timestamp 1698431365
transform -1 0 6600 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_258
timestamp 1698431365
transform -1 0 6600 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_259
timestamp 1698431365
transform -1 0 6600 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_260
timestamp 1698431365
transform -1 0 6600 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_261
timestamp 1698431365
transform -1 0 6600 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_262
timestamp 1698431365
transform -1 0 6600 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_263
timestamp 1698431365
transform -1 0 6600 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_264
timestamp 1698431365
transform -1 0 10800 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_265
timestamp 1698431365
transform -1 0 10800 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_266
timestamp 1698431365
transform -1 0 10800 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_267
timestamp 1698431365
transform -1 0 10800 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_268
timestamp 1698431365
transform -1 0 10200 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_269
timestamp 1698431365
transform -1 0 10200 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_270
timestamp 1698431365
transform -1 0 10200 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_271
timestamp 1698431365
transform -1 0 10200 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_272
timestamp 1698431365
transform -1 0 10200 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_273
timestamp 1698431365
transform -1 0 10200 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_274
timestamp 1698431365
transform -1 0 10200 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_275
timestamp 1698431365
transform -1 0 8400 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_276
timestamp 1698431365
transform -1 0 8400 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_277
timestamp 1698431365
transform -1 0 8400 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_278
timestamp 1698431365
transform -1 0 9000 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_279
timestamp 1698431365
transform -1 0 9000 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_280
timestamp 1698431365
transform -1 0 9000 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_281
timestamp 1698431365
transform -1 0 9000 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_282
timestamp 1698431365
transform -1 0 7200 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_283
timestamp 1698431365
transform -1 0 7200 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_284
timestamp 1698431365
transform -1 0 7200 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_285
timestamp 1698431365
transform -1 0 7200 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_286
timestamp 1698431365
transform -1 0 7200 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_287
timestamp 1698431365
transform -1 0 7200 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_288
timestamp 1698431365
transform -1 0 7200 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_289
timestamp 1698431365
transform -1 0 9000 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_290
timestamp 1698431365
transform -1 0 9000 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_291
timestamp 1698431365
transform -1 0 9000 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_292
timestamp 1698431365
transform -1 0 8400 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_293
timestamp 1698431365
transform -1 0 8400 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_294
timestamp 1698431365
transform -1 0 8400 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_295
timestamp 1698431365
transform -1 0 8400 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_296
timestamp 1698431365
transform 1 0 1800 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_297
timestamp 1698431365
transform 1 0 600 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_298
timestamp 1698431365
transform 1 0 600 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_299
timestamp 1698431365
transform 1 0 600 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_300
timestamp 1698431365
transform 1 0 2400 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_301
timestamp 1698431365
transform 1 0 2400 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_302
timestamp 1698431365
transform 1 0 2400 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_303
timestamp 1698431365
transform 1 0 2400 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_304
timestamp 1698431365
transform 1 0 2400 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_305
timestamp 1698431365
transform 1 0 2400 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_306
timestamp 1698431365
transform 1 0 600 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_307
timestamp 1698431365
transform 1 0 600 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_308
timestamp 1698431365
transform 1 0 600 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_309
timestamp 1698431365
transform 1 0 1200 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_310
timestamp 1698431365
transform 1 0 1200 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_311
timestamp 1698431365
transform 1 0 1200 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_312
timestamp 1698431365
transform 1 0 4800 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_313
timestamp 1698431365
transform 1 0 4800 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_314
timestamp 1698431365
transform 1 0 4800 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_315
timestamp 1698431365
transform 1 0 4800 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_316
timestamp 1698431365
transform 1 0 4800 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_317
timestamp 1698431365
transform 1 0 4800 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_318
timestamp 1698431365
transform 1 0 4800 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_319
timestamp 1698431365
transform 1 0 1200 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_320
timestamp 1698431365
transform 1 0 1200 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_321
timestamp 1698431365
transform 1 0 4200 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_322
timestamp 1698431365
transform 1 0 4200 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_323
timestamp 1698431365
transform 1 0 4200 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_324
timestamp 1698431365
transform 1 0 4200 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_325
timestamp 1698431365
transform 1 0 4200 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_326
timestamp 1698431365
transform 1 0 1200 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_327
timestamp 1698431365
transform 1 0 3000 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_328
timestamp 1698431365
transform 1 0 3000 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_329
timestamp 1698431365
transform 1 0 3000 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_330
timestamp 1698431365
transform 1 0 3000 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_331
timestamp 1698431365
transform 1 0 4200 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_332
timestamp 1698431365
transform 1 0 4200 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_333
timestamp 1698431365
transform 1 0 3000 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_334
timestamp 1698431365
transform 1 0 3000 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_335
timestamp 1698431365
transform 1 0 3000 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_336
timestamp 1698431365
transform 1 0 3600 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_337
timestamp 1698431365
transform 1 0 3600 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_338
timestamp 1698431365
transform 1 0 3600 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_339
timestamp 1698431365
transform 1 0 3600 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_340
timestamp 1698431365
transform 1 0 3600 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_341
timestamp 1698431365
transform 1 0 2400 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_342
timestamp 1698431365
transform 1 0 3600 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_343
timestamp 1698431365
transform 1 0 3600 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_344
timestamp 1698431365
transform 1 0 1200 0 1 10800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_345
timestamp 1698431365
transform 1 0 1800 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_346
timestamp 1698431365
transform 1 0 600 0 1 1800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_347
timestamp 1698431365
transform 1 0 1800 0 1 0
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_348
timestamp 1698431365
transform 1 0 1800 0 1 3600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_349
timestamp 1698431365
transform 1 0 1800 0 1 5400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_350
timestamp 1698431365
transform 1 0 1800 0 1 7200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_351
timestamp 1698431365
transform 1 0 1800 0 1 9000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_352
timestamp 1698431365
transform 1 0 1200 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_353
timestamp 1698431365
transform 1 0 1200 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_354
timestamp 1698431365
transform 1 0 1200 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_355
timestamp 1698431365
transform 1 0 4800 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_356
timestamp 1698431365
transform 1 0 4800 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_357
timestamp 1698431365
transform 1 0 4800 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_358
timestamp 1698431365
transform 1 0 4800 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_359
timestamp 1698431365
transform 1 0 4800 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_360
timestamp 1698431365
transform 1 0 2400 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_361
timestamp 1698431365
transform 1 0 2400 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_362
timestamp 1698431365
transform 1 0 2400 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_363
timestamp 1698431365
transform 1 0 2400 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_364
timestamp 1698431365
transform 1 0 2400 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_365
timestamp 1698431365
transform 1 0 2400 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_366
timestamp 1698431365
transform 1 0 3600 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_367
timestamp 1698431365
transform 1 0 3600 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_368
timestamp 1698431365
transform 1 0 3600 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_369
timestamp 1698431365
transform 1 0 3600 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_370
timestamp 1698431365
transform 1 0 3600 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_371
timestamp 1698431365
transform 1 0 1200 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_372
timestamp 1698431365
transform 1 0 1200 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_373
timestamp 1698431365
transform 1 0 4800 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_374
timestamp 1698431365
transform 1 0 600 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_375
timestamp 1698431365
transform 1 0 600 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_376
timestamp 1698431365
transform 1 0 600 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_377
timestamp 1698431365
transform 1 0 600 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_378
timestamp 1698431365
transform 1 0 3600 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_379
timestamp 1698431365
transform 1 0 1800 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_380
timestamp 1698431365
transform 1 0 4200 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_381
timestamp 1698431365
transform 1 0 4200 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_382
timestamp 1698431365
transform 1 0 4200 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_383
timestamp 1698431365
transform 1 0 4200 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_384
timestamp 1698431365
transform 1 0 4200 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_385
timestamp 1698431365
transform 1 0 4200 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_386
timestamp 1698431365
transform 1 0 3000 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_387
timestamp 1698431365
transform 1 0 3000 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_388
timestamp 1698431365
transform 1 0 3000 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_389
timestamp 1698431365
transform 1 0 3000 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_390
timestamp 1698431365
transform 1 0 3000 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_391
timestamp 1698431365
transform 1 0 3000 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_392
timestamp 1698431365
transform 1 0 600 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_393
timestamp 1698431365
transform 1 0 600 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_394
timestamp 1698431365
transform 1 0 1800 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_395
timestamp 1698431365
transform 1 0 1800 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_396
timestamp 1698431365
transform 1 0 1800 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_397
timestamp 1698431365
transform 1 0 1800 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_398
timestamp 1698431365
transform 1 0 1800 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_399
timestamp 1698431365
transform 1 0 1200 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_400
timestamp 1698431365
transform -1 0 10200 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_401
timestamp 1698431365
transform -1 0 10200 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_402
timestamp 1698431365
transform -1 0 10200 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_403
timestamp 1698431365
transform -1 0 10200 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_404
timestamp 1698431365
transform -1 0 10200 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_405
timestamp 1698431365
transform -1 0 10200 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_406
timestamp 1698431365
transform -1 0 10800 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_407
timestamp 1698431365
transform -1 0 10800 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_408
timestamp 1698431365
transform -1 0 10800 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_409
timestamp 1698431365
transform -1 0 8400 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_410
timestamp 1698431365
transform -1 0 8400 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_411
timestamp 1698431365
transform -1 0 7200 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_412
timestamp 1698431365
transform -1 0 7200 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_413
timestamp 1698431365
transform -1 0 7200 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_414
timestamp 1698431365
transform -1 0 7200 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_415
timestamp 1698431365
transform -1 0 7200 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_416
timestamp 1698431365
transform -1 0 7200 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_417
timestamp 1698431365
transform -1 0 8400 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_418
timestamp 1698431365
transform -1 0 8400 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_419
timestamp 1698431365
transform -1 0 8400 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_420
timestamp 1698431365
transform -1 0 8400 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_421
timestamp 1698431365
transform -1 0 6600 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_422
timestamp 1698431365
transform -1 0 6600 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_423
timestamp 1698431365
transform -1 0 6600 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_424
timestamp 1698431365
transform -1 0 6600 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_425
timestamp 1698431365
transform -1 0 6600 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_426
timestamp 1698431365
transform -1 0 6600 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_427
timestamp 1698431365
transform -1 0 10800 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_428
timestamp 1698431365
transform -1 0 10800 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_429
timestamp 1698431365
transform -1 0 10800 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_430
timestamp 1698431365
transform -1 0 7800 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_431
timestamp 1698431365
transform -1 0 9600 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_432
timestamp 1698431365
transform -1 0 9600 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_433
timestamp 1698431365
transform -1 0 9600 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_434
timestamp 1698431365
transform -1 0 9600 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_435
timestamp 1698431365
transform -1 0 9600 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_436
timestamp 1698431365
transform -1 0 9600 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_437
timestamp 1698431365
transform -1 0 7800 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_438
timestamp 1698431365
transform -1 0 7800 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_439
timestamp 1698431365
transform -1 0 7800 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_440
timestamp 1698431365
transform -1 0 7800 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_441
timestamp 1698431365
transform -1 0 9000 0 1 16200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_442
timestamp 1698431365
transform -1 0 9000 0 1 18000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_443
timestamp 1698431365
transform -1 0 9000 0 1 19800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_444
timestamp 1698431365
transform -1 0 9000 0 1 21600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_445
timestamp 1698431365
transform -1 0 9000 0 1 23400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_446
timestamp 1698431365
transform -1 0 9000 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_447
timestamp 1698431365
transform -1 0 7800 0 1 25200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_448
timestamp 1698431365
transform 1 0 2400 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_449
timestamp 1698431365
transform 1 0 2400 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_450
timestamp 1698431365
transform -1 0 7200 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_451
timestamp 1698431365
transform -1 0 7200 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_452
timestamp 1698431365
transform 1 0 4200 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_453
timestamp 1698431365
transform 1 0 4200 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_454
timestamp 1698431365
transform -1 0 6600 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_455
timestamp 1698431365
transform -1 0 6600 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_456
timestamp 1698431365
transform 1 0 600 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_457
timestamp 1698431365
transform 1 0 600 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_458
timestamp 1698431365
transform -1 0 9600 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_459
timestamp 1698431365
transform -1 0 9600 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_460
timestamp 1698431365
transform 1 0 4800 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_461
timestamp 1698431365
transform 1 0 4800 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_462
timestamp 1698431365
transform -1 0 9000 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_463
timestamp 1698431365
transform -1 0 9000 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_464
timestamp 1698431365
transform 1 0 3000 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_465
timestamp 1698431365
transform -1 0 8400 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_466
timestamp 1698431365
transform -1 0 8400 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_467
timestamp 1698431365
transform 1 0 3000 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_468
timestamp 1698431365
transform -1 0 7800 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_469
timestamp 1698431365
transform -1 0 7800 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_470
timestamp 1698431365
transform 1 0 1800 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_471
timestamp 1698431365
transform 1 0 1800 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_472
timestamp 1698431365
transform 1 0 1200 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_473
timestamp 1698431365
transform -1 0 10800 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_474
timestamp 1698431365
transform -1 0 10800 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_475
timestamp 1698431365
transform 1 0 1200 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_476
timestamp 1698431365
transform 1 0 3600 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_477
timestamp 1698431365
transform 1 0 3600 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_478
timestamp 1698431365
transform -1 0 10200 0 1 12600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_479
timestamp 1698431365
transform -1 0 10200 0 1 14400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_480
timestamp 1698431365
transform -1 0 7200 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_481
timestamp 1698431365
transform -1 0 9000 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_482
timestamp 1698431365
transform -1 0 7800 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_483
timestamp 1698431365
transform -1 0 10200 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_484
timestamp 1698431365
transform -1 0 8400 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_485
timestamp 1698431365
transform -1 0 10200 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_486
timestamp 1698431365
transform -1 0 10800 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_487
timestamp 1698431365
transform -1 0 10800 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_488
timestamp 1698431365
transform -1 0 10800 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_489
timestamp 1698431365
transform -1 0 10800 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_490
timestamp 1698431365
transform -1 0 9000 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_491
timestamp 1698431365
transform -1 0 9000 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_492
timestamp 1698431365
transform -1 0 9000 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_493
timestamp 1698431365
transform -1 0 9000 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_494
timestamp 1698431365
transform -1 0 9000 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_495
timestamp 1698431365
transform -1 0 6600 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_496
timestamp 1698431365
transform -1 0 6600 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_497
timestamp 1698431365
transform -1 0 6600 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_498
timestamp 1698431365
transform -1 0 6600 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_499
timestamp 1698431365
transform -1 0 6600 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_500
timestamp 1698431365
transform -1 0 6600 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_501
timestamp 1698431365
transform -1 0 10800 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_502
timestamp 1698431365
transform -1 0 10200 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_503
timestamp 1698431365
transform -1 0 10200 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_504
timestamp 1698431365
transform -1 0 10200 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_505
timestamp 1698431365
transform -1 0 10800 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_506
timestamp 1698431365
transform -1 0 10200 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_507
timestamp 1698431365
transform -1 0 7800 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_508
timestamp 1698431365
transform -1 0 7800 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_509
timestamp 1698431365
transform -1 0 7800 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_510
timestamp 1698431365
transform -1 0 9600 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_511
timestamp 1698431365
transform -1 0 8400 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_512
timestamp 1698431365
transform -1 0 7800 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_513
timestamp 1698431365
transform -1 0 9600 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_514
timestamp 1698431365
transform -1 0 9600 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_515
timestamp 1698431365
transform -1 0 9600 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_516
timestamp 1698431365
transform -1 0 9600 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_517
timestamp 1698431365
transform -1 0 9600 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_518
timestamp 1698431365
transform -1 0 7800 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_519
timestamp 1698431365
transform -1 0 8400 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_520
timestamp 1698431365
transform -1 0 8400 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_521
timestamp 1698431365
transform -1 0 7200 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_522
timestamp 1698431365
transform -1 0 8400 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_523
timestamp 1698431365
transform -1 0 8400 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_524
timestamp 1698431365
transform -1 0 7200 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_525
timestamp 1698431365
transform -1 0 7200 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_526
timestamp 1698431365
transform -1 0 7200 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_527
timestamp 1698431365
transform -1 0 7200 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_528
timestamp 1698431365
transform 1 0 4800 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_529
timestamp 1698431365
transform 1 0 3600 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_530
timestamp 1698431365
transform 1 0 1200 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_531
timestamp 1698431365
transform 1 0 1800 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_532
timestamp 1698431365
transform 1 0 1800 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_533
timestamp 1698431365
transform 1 0 1800 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_534
timestamp 1698431365
transform 1 0 1800 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_535
timestamp 1698431365
transform 1 0 1800 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_536
timestamp 1698431365
transform 1 0 1800 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_537
timestamp 1698431365
transform 1 0 3000 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_538
timestamp 1698431365
transform 1 0 2400 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_539
timestamp 1698431365
transform 1 0 4200 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_540
timestamp 1698431365
transform 1 0 2400 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_541
timestamp 1698431365
transform 1 0 2400 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_542
timestamp 1698431365
transform 1 0 2400 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_543
timestamp 1698431365
transform 1 0 2400 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_544
timestamp 1698431365
transform 1 0 2400 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_545
timestamp 1698431365
transform 1 0 4200 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_546
timestamp 1698431365
transform 1 0 1200 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_547
timestamp 1698431365
transform 1 0 3000 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_548
timestamp 1698431365
transform 1 0 3000 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_549
timestamp 1698431365
transform 1 0 3000 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_550
timestamp 1698431365
transform 1 0 3000 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_551
timestamp 1698431365
transform 1 0 3000 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_552
timestamp 1698431365
transform 1 0 600 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_553
timestamp 1698431365
transform 1 0 1200 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_554
timestamp 1698431365
transform 1 0 4200 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_555
timestamp 1698431365
transform 1 0 1200 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_556
timestamp 1698431365
transform 1 0 600 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_557
timestamp 1698431365
transform 1 0 600 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_558
timestamp 1698431365
transform 1 0 600 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_559
timestamp 1698431365
transform 1 0 600 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_560
timestamp 1698431365
transform 1 0 600 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_561
timestamp 1698431365
transform 1 0 1200 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_562
timestamp 1698431365
transform 1 0 1200 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_563
timestamp 1698431365
transform 1 0 3600 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_564
timestamp 1698431365
transform 1 0 4200 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_565
timestamp 1698431365
transform 1 0 3600 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_566
timestamp 1698431365
transform 1 0 3600 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_567
timestamp 1698431365
transform 1 0 4800 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_568
timestamp 1698431365
transform 1 0 4800 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_569
timestamp 1698431365
transform 1 0 4800 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_570
timestamp 1698431365
transform 1 0 4800 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_571
timestamp 1698431365
transform 1 0 4800 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_572
timestamp 1698431365
transform 1 0 3600 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_573
timestamp 1698431365
transform 1 0 3600 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_574
timestamp 1698431365
transform 1 0 4200 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_575
timestamp 1698431365
transform 1 0 4200 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_576
timestamp 1698431365
transform 1 0 3600 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_577
timestamp 1698431365
transform 1 0 3600 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_578
timestamp 1698431365
transform 1 0 1800 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_579
timestamp 1698431365
transform 1 0 1800 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_580
timestamp 1698431365
transform 1 0 1800 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_581
timestamp 1698431365
transform 1 0 1800 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_582
timestamp 1698431365
transform 1 0 1800 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_583
timestamp 1698431365
transform 1 0 1800 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_584
timestamp 1698431365
transform 1 0 1800 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_585
timestamp 1698431365
transform 1 0 3600 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_586
timestamp 1698431365
transform 1 0 3600 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_587
timestamp 1698431365
transform 1 0 2400 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_588
timestamp 1698431365
transform 1 0 2400 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_589
timestamp 1698431365
transform 1 0 2400 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_590
timestamp 1698431365
transform 1 0 2400 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_591
timestamp 1698431365
transform 1 0 2400 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_592
timestamp 1698431365
transform 1 0 2400 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_593
timestamp 1698431365
transform 1 0 2400 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_594
timestamp 1698431365
transform 1 0 3600 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_595
timestamp 1698431365
transform 1 0 3600 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_596
timestamp 1698431365
transform 1 0 4200 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_597
timestamp 1698431365
transform 1 0 4200 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_598
timestamp 1698431365
transform 1 0 3600 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_599
timestamp 1698431365
transform 1 0 600 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_600
timestamp 1698431365
transform 1 0 600 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_601
timestamp 1698431365
transform 1 0 600 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_602
timestamp 1698431365
transform 1 0 600 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_603
timestamp 1698431365
transform 1 0 4200 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_604
timestamp 1698431365
transform 1 0 4200 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_605
timestamp 1698431365
transform 1 0 600 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_606
timestamp 1698431365
transform 1 0 600 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_607
timestamp 1698431365
transform 1 0 600 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_608
timestamp 1698431365
transform 1 0 1200 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_609
timestamp 1698431365
transform 1 0 1200 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_610
timestamp 1698431365
transform 1 0 4200 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_611
timestamp 1698431365
transform 1 0 1200 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_612
timestamp 1698431365
transform 1 0 1200 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_613
timestamp 1698431365
transform 1 0 4800 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_614
timestamp 1698431365
transform 1 0 4800 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_615
timestamp 1698431365
transform 1 0 4800 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_616
timestamp 1698431365
transform 1 0 4800 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_617
timestamp 1698431365
transform 1 0 4800 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_618
timestamp 1698431365
transform 1 0 4800 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_619
timestamp 1698431365
transform 1 0 4800 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_620
timestamp 1698431365
transform 1 0 1200 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_621
timestamp 1698431365
transform 1 0 1200 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_622
timestamp 1698431365
transform 1 0 3000 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_623
timestamp 1698431365
transform 1 0 3000 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_624
timestamp 1698431365
transform 1 0 3000 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_625
timestamp 1698431365
transform 1 0 3000 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_626
timestamp 1698431365
transform 1 0 3000 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_627
timestamp 1698431365
transform 1 0 3000 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_628
timestamp 1698431365
transform 1 0 3000 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_629
timestamp 1698431365
transform 1 0 4200 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_630
timestamp 1698431365
transform 1 0 4200 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_631
timestamp 1698431365
transform 1 0 1200 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_632
timestamp 1698431365
transform -1 0 7800 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_633
timestamp 1698431365
transform -1 0 7800 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_634
timestamp 1698431365
transform -1 0 7800 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_635
timestamp 1698431365
transform -1 0 7800 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_636
timestamp 1698431365
transform -1 0 7800 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_637
timestamp 1698431365
transform -1 0 10200 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_638
timestamp 1698431365
transform -1 0 7200 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_639
timestamp 1698431365
transform -1 0 7200 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_640
timestamp 1698431365
transform -1 0 7200 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_641
timestamp 1698431365
transform -1 0 7200 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_642
timestamp 1698431365
transform -1 0 7200 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_643
timestamp 1698431365
transform -1 0 7200 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_644
timestamp 1698431365
transform -1 0 7200 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_645
timestamp 1698431365
transform -1 0 10200 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_646
timestamp 1698431365
transform -1 0 10800 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_647
timestamp 1698431365
transform -1 0 10800 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_648
timestamp 1698431365
transform -1 0 6600 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_649
timestamp 1698431365
transform -1 0 6600 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_650
timestamp 1698431365
transform -1 0 6600 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_651
timestamp 1698431365
transform -1 0 6600 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_652
timestamp 1698431365
transform -1 0 6600 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_653
timestamp 1698431365
transform -1 0 6600 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_654
timestamp 1698431365
transform -1 0 6600 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_655
timestamp 1698431365
transform -1 0 10800 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_656
timestamp 1698431365
transform -1 0 10800 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_657
timestamp 1698431365
transform -1 0 9600 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_658
timestamp 1698431365
transform -1 0 9600 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_659
timestamp 1698431365
transform -1 0 9600 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_660
timestamp 1698431365
transform -1 0 9600 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_661
timestamp 1698431365
transform -1 0 9600 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_662
timestamp 1698431365
transform -1 0 9600 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_663
timestamp 1698431365
transform -1 0 9600 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_664
timestamp 1698431365
transform -1 0 10800 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_665
timestamp 1698431365
transform -1 0 10800 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_666
timestamp 1698431365
transform -1 0 9000 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_667
timestamp 1698431365
transform -1 0 9000 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_668
timestamp 1698431365
transform -1 0 9000 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_669
timestamp 1698431365
transform -1 0 9000 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_670
timestamp 1698431365
transform -1 0 9000 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_671
timestamp 1698431365
transform -1 0 9000 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_672
timestamp 1698431365
transform -1 0 9000 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_673
timestamp 1698431365
transform -1 0 10800 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_674
timestamp 1698431365
transform -1 0 10200 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_675
timestamp 1698431365
transform -1 0 10200 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_676
timestamp 1698431365
transform -1 0 10200 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_677
timestamp 1698431365
transform -1 0 8400 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_678
timestamp 1698431365
transform -1 0 8400 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_679
timestamp 1698431365
transform -1 0 8400 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_680
timestamp 1698431365
transform -1 0 8400 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_681
timestamp 1698431365
transform -1 0 8400 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_682
timestamp 1698431365
transform -1 0 8400 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_683
timestamp 1698431365
transform -1 0 8400 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_684
timestamp 1698431365
transform -1 0 10200 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_685
timestamp 1698431365
transform -1 0 10200 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_686
timestamp 1698431365
transform -1 0 7800 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_687
timestamp 1698431365
transform -1 0 7800 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_688
timestamp 1698431365
transform 1 0 1800 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_689
timestamp 1698431365
transform 1 0 1800 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_690
timestamp 1698431365
transform 1 0 2400 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_691
timestamp 1698431365
transform 1 0 2400 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_692
timestamp 1698431365
transform -1 0 7200 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_693
timestamp 1698431365
transform -1 0 7200 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_694
timestamp 1698431365
transform -1 0 6600 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_695
timestamp 1698431365
transform -1 0 6600 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_696
timestamp 1698431365
transform -1 0 9600 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_697
timestamp 1698431365
transform -1 0 9600 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_698
timestamp 1698431365
transform -1 0 9000 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_699
timestamp 1698431365
transform -1 0 9000 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_700
timestamp 1698431365
transform 1 0 4200 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_701
timestamp 1698431365
transform 1 0 4200 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_702
timestamp 1698431365
transform -1 0 8400 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_703
timestamp 1698431365
transform -1 0 8400 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_704
timestamp 1698431365
transform -1 0 7800 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_705
timestamp 1698431365
transform -1 0 7800 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_706
timestamp 1698431365
transform -1 0 10800 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_707
timestamp 1698431365
transform -1 0 10800 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_708
timestamp 1698431365
transform -1 0 10200 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_709
timestamp 1698431365
transform -1 0 10200 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_710
timestamp 1698431365
transform 1 0 4800 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_711
timestamp 1698431365
transform 1 0 4800 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_712
timestamp 1698431365
transform 1 0 3000 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_713
timestamp 1698431365
transform 1 0 3000 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_714
timestamp 1698431365
transform 1 0 3600 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_715
timestamp 1698431365
transform 1 0 3600 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_716
timestamp 1698431365
transform 1 0 600 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_717
timestamp 1698431365
transform 1 0 600 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_718
timestamp 1698431365
transform 1 0 1200 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_719
timestamp 1698431365
transform 1 0 1200 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_720
timestamp 1698431365
transform -1 0 17400 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_721
timestamp 1698431365
transform -1 0 21000 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_722
timestamp 1698431365
transform -1 0 18000 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_723
timestamp 1698431365
transform -1 0 18600 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_724
timestamp 1698431365
transform -1 0 20400 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_725
timestamp 1698431365
transform -1 0 20400 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_726
timestamp 1698431365
transform -1 0 19800 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_727
timestamp 1698431365
transform -1 0 19800 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_728
timestamp 1698431365
transform -1 0 18000 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_729
timestamp 1698431365
transform -1 0 18000 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_730
timestamp 1698431365
transform -1 0 18000 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_731
timestamp 1698431365
transform -1 0 18000 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_732
timestamp 1698431365
transform -1 0 18600 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_733
timestamp 1698431365
transform -1 0 18600 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_734
timestamp 1698431365
transform -1 0 18600 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_735
timestamp 1698431365
transform -1 0 18600 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_736
timestamp 1698431365
transform -1 0 18000 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_737
timestamp 1698431365
transform -1 0 21000 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_738
timestamp 1698431365
transform -1 0 17400 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_739
timestamp 1698431365
transform -1 0 17400 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_740
timestamp 1698431365
transform -1 0 17400 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_741
timestamp 1698431365
transform -1 0 17400 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_742
timestamp 1698431365
transform -1 0 17400 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_743
timestamp 1698431365
transform -1 0 21000 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_744
timestamp 1698431365
transform -1 0 21000 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_745
timestamp 1698431365
transform -1 0 21000 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_746
timestamp 1698431365
transform -1 0 21000 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_747
timestamp 1698431365
transform -1 0 18600 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_748
timestamp 1698431365
transform -1 0 19800 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_749
timestamp 1698431365
transform -1 0 19200 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_750
timestamp 1698431365
transform -1 0 19800 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_751
timestamp 1698431365
transform -1 0 20400 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_752
timestamp 1698431365
transform -1 0 19200 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_753
timestamp 1698431365
transform -1 0 19200 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_754
timestamp 1698431365
transform -1 0 19200 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_755
timestamp 1698431365
transform -1 0 19200 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_756
timestamp 1698431365
transform -1 0 19200 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_757
timestamp 1698431365
transform -1 0 19800 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_758
timestamp 1698431365
transform -1 0 19800 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_759
timestamp 1698431365
transform -1 0 21600 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_760
timestamp 1698431365
transform -1 0 20400 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_761
timestamp 1698431365
transform -1 0 20400 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_762
timestamp 1698431365
transform -1 0 21600 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_763
timestamp 1698431365
transform -1 0 21600 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_764
timestamp 1698431365
transform -1 0 21600 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_765
timestamp 1698431365
transform -1 0 21600 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_766
timestamp 1698431365
transform -1 0 21600 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_767
timestamp 1698431365
transform -1 0 20400 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_768
timestamp 1698431365
transform 1 0 15000 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_769
timestamp 1698431365
transform 1 0 11400 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_770
timestamp 1698431365
transform 1 0 15000 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_771
timestamp 1698431365
transform 1 0 15000 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_772
timestamp 1698431365
transform 1 0 13800 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_773
timestamp 1698431365
transform 1 0 13800 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_774
timestamp 1698431365
transform 1 0 12600 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_775
timestamp 1698431365
transform 1 0 12600 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_776
timestamp 1698431365
transform 1 0 12600 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_777
timestamp 1698431365
transform 1 0 12600 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_778
timestamp 1698431365
transform 1 0 11400 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_779
timestamp 1698431365
transform 1 0 12600 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_780
timestamp 1698431365
transform 1 0 13200 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_781
timestamp 1698431365
transform 1 0 13200 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_782
timestamp 1698431365
transform 1 0 15600 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_783
timestamp 1698431365
transform 1 0 15600 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_784
timestamp 1698431365
transform 1 0 15600 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_785
timestamp 1698431365
transform 1 0 15600 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_786
timestamp 1698431365
transform 1 0 15600 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_787
timestamp 1698431365
transform 1 0 13200 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_788
timestamp 1698431365
transform 1 0 11400 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_789
timestamp 1698431365
transform 1 0 11400 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_790
timestamp 1698431365
transform 1 0 11400 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_791
timestamp 1698431365
transform 1 0 11400 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_792
timestamp 1698431365
transform 1 0 13200 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_793
timestamp 1698431365
transform 1 0 12600 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_794
timestamp 1698431365
transform 1 0 13200 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_795
timestamp 1698431365
transform 1 0 14400 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_796
timestamp 1698431365
transform 1 0 14400 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_797
timestamp 1698431365
transform 1 0 14400 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_798
timestamp 1698431365
transform 1 0 14400 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_799
timestamp 1698431365
transform 1 0 14400 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_800
timestamp 1698431365
transform 1 0 13800 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_801
timestamp 1698431365
transform 1 0 12000 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_802
timestamp 1698431365
transform 1 0 12000 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_803
timestamp 1698431365
transform 1 0 12000 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_804
timestamp 1698431365
transform 1 0 13800 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_805
timestamp 1698431365
transform 1 0 13800 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_806
timestamp 1698431365
transform 1 0 13800 0 1 36000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_807
timestamp 1698431365
transform 1 0 14400 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_808
timestamp 1698431365
transform 1 0 13200 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_809
timestamp 1698431365
transform 1 0 12000 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_810
timestamp 1698431365
transform 1 0 15600 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_811
timestamp 1698431365
transform 1 0 15000 0 1 30600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_812
timestamp 1698431365
transform 1 0 15000 0 1 32400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_813
timestamp 1698431365
transform 1 0 12000 0 1 37800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_814
timestamp 1698431365
transform 1 0 12000 0 1 39600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_815
timestamp 1698431365
transform 1 0 15000 0 1 34200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_816
timestamp 1698431365
transform 1 0 12000 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_817
timestamp 1698431365
transform 1 0 12000 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_818
timestamp 1698431365
transform 1 0 12600 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_819
timestamp 1698431365
transform 1 0 15000 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_820
timestamp 1698431365
transform 1 0 15000 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_821
timestamp 1698431365
transform 1 0 15000 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_822
timestamp 1698431365
transform 1 0 15000 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_823
timestamp 1698431365
transform 1 0 15000 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_824
timestamp 1698431365
transform 1 0 15000 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_825
timestamp 1698431365
transform 1 0 15000 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_826
timestamp 1698431365
transform 1 0 12600 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_827
timestamp 1698431365
transform 1 0 12000 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_828
timestamp 1698431365
transform 1 0 12000 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_829
timestamp 1698431365
transform 1 0 12600 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_830
timestamp 1698431365
transform 1 0 15600 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_831
timestamp 1698431365
transform 1 0 15600 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_832
timestamp 1698431365
transform 1 0 15600 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_833
timestamp 1698431365
transform 1 0 15600 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_834
timestamp 1698431365
transform 1 0 15600 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_835
timestamp 1698431365
transform 1 0 15600 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_836
timestamp 1698431365
transform 1 0 11400 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_837
timestamp 1698431365
transform 1 0 11400 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_838
timestamp 1698431365
transform 1 0 11400 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_839
timestamp 1698431365
transform 1 0 11400 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_840
timestamp 1698431365
transform 1 0 11400 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_841
timestamp 1698431365
transform 1 0 11400 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_842
timestamp 1698431365
transform 1 0 11400 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_843
timestamp 1698431365
transform 1 0 15600 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_844
timestamp 1698431365
transform 1 0 12600 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_845
timestamp 1698431365
transform 1 0 12000 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_846
timestamp 1698431365
transform 1 0 12000 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_847
timestamp 1698431365
transform 1 0 12600 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_848
timestamp 1698431365
transform 1 0 13800 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_849
timestamp 1698431365
transform 1 0 13800 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_850
timestamp 1698431365
transform 1 0 13800 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_851
timestamp 1698431365
transform 1 0 13800 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_852
timestamp 1698431365
transform 1 0 13800 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_853
timestamp 1698431365
transform 1 0 13800 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_854
timestamp 1698431365
transform 1 0 13800 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_855
timestamp 1698431365
transform 1 0 13200 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_856
timestamp 1698431365
transform 1 0 12000 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_857
timestamp 1698431365
transform 1 0 13200 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_858
timestamp 1698431365
transform 1 0 13200 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_859
timestamp 1698431365
transform 1 0 13200 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_860
timestamp 1698431365
transform 1 0 14400 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_861
timestamp 1698431365
transform 1 0 14400 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_862
timestamp 1698431365
transform 1 0 14400 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_863
timestamp 1698431365
transform 1 0 14400 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_864
timestamp 1698431365
transform 1 0 14400 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_865
timestamp 1698431365
transform 1 0 14400 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_866
timestamp 1698431365
transform 1 0 14400 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_867
timestamp 1698431365
transform 1 0 13200 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_868
timestamp 1698431365
transform 1 0 13200 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_869
timestamp 1698431365
transform 1 0 13200 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_870
timestamp 1698431365
transform 1 0 12600 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_871
timestamp 1698431365
transform 1 0 12600 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_872
timestamp 1698431365
transform -1 0 18000 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_873
timestamp 1698431365
transform -1 0 18000 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_874
timestamp 1698431365
transform -1 0 18000 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_875
timestamp 1698431365
transform -1 0 18000 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_876
timestamp 1698431365
transform -1 0 18000 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_877
timestamp 1698431365
transform -1 0 18000 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_878
timestamp 1698431365
transform -1 0 18000 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_879
timestamp 1698431365
transform -1 0 19800 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_880
timestamp 1698431365
transform -1 0 19800 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_881
timestamp 1698431365
transform -1 0 19800 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_882
timestamp 1698431365
transform -1 0 19800 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_883
timestamp 1698431365
transform -1 0 17400 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_884
timestamp 1698431365
transform -1 0 17400 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_885
timestamp 1698431365
transform -1 0 17400 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_886
timestamp 1698431365
transform -1 0 17400 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_887
timestamp 1698431365
transform -1 0 17400 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_888
timestamp 1698431365
transform -1 0 17400 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_889
timestamp 1698431365
transform -1 0 17400 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_890
timestamp 1698431365
transform -1 0 19800 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_891
timestamp 1698431365
transform -1 0 21600 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_892
timestamp 1698431365
transform -1 0 21600 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_893
timestamp 1698431365
transform -1 0 21600 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_894
timestamp 1698431365
transform -1 0 21600 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_895
timestamp 1698431365
transform -1 0 21600 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_896
timestamp 1698431365
transform -1 0 21600 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_897
timestamp 1698431365
transform -1 0 21600 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_898
timestamp 1698431365
transform -1 0 21000 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_899
timestamp 1698431365
transform -1 0 21000 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_900
timestamp 1698431365
transform -1 0 21000 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_901
timestamp 1698431365
transform -1 0 21000 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_902
timestamp 1698431365
transform -1 0 21000 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_903
timestamp 1698431365
transform -1 0 21000 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_904
timestamp 1698431365
transform -1 0 21000 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_905
timestamp 1698431365
transform -1 0 19200 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_906
timestamp 1698431365
transform -1 0 19200 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_907
timestamp 1698431365
transform -1 0 19200 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_908
timestamp 1698431365
transform -1 0 19200 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_909
timestamp 1698431365
transform -1 0 19200 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_910
timestamp 1698431365
transform -1 0 19200 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_911
timestamp 1698431365
transform -1 0 19200 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_912
timestamp 1698431365
transform -1 0 18600 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_913
timestamp 1698431365
transform -1 0 18600 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_914
timestamp 1698431365
transform -1 0 18600 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_915
timestamp 1698431365
transform -1 0 18600 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_916
timestamp 1698431365
transform -1 0 18600 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_917
timestamp 1698431365
transform -1 0 18600 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_918
timestamp 1698431365
transform -1 0 18600 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_919
timestamp 1698431365
transform -1 0 20400 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_920
timestamp 1698431365
transform -1 0 20400 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_921
timestamp 1698431365
transform -1 0 20400 0 1 48600
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_922
timestamp 1698431365
transform -1 0 20400 0 1 50400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_923
timestamp 1698431365
transform -1 0 20400 0 1 52200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_924
timestamp 1698431365
transform -1 0 20400 0 1 54000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_925
timestamp 1698431365
transform -1 0 20400 0 1 55800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_926
timestamp 1698431365
transform -1 0 19800 0 1 45000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_927
timestamp 1698431365
transform -1 0 19800 0 1 46800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_928
timestamp 1698431365
transform -1 0 18000 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_929
timestamp 1698431365
transform -1 0 18000 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_930
timestamp 1698431365
transform -1 0 17400 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_931
timestamp 1698431365
transform -1 0 17400 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_932
timestamp 1698431365
transform 1 0 11400 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_933
timestamp 1698431365
transform 1 0 11400 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_934
timestamp 1698431365
transform -1 0 21600 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_935
timestamp 1698431365
transform -1 0 21600 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_936
timestamp 1698431365
transform -1 0 21000 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_937
timestamp 1698431365
transform -1 0 21000 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_938
timestamp 1698431365
transform 1 0 12000 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_939
timestamp 1698431365
transform 1 0 12000 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_940
timestamp 1698431365
transform -1 0 19200 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_941
timestamp 1698431365
transform -1 0 19200 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_942
timestamp 1698431365
transform -1 0 18600 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_943
timestamp 1698431365
transform -1 0 18600 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_944
timestamp 1698431365
transform -1 0 20400 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_945
timestamp 1698431365
transform -1 0 20400 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_946
timestamp 1698431365
transform -1 0 19800 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_947
timestamp 1698431365
transform -1 0 19800 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_948
timestamp 1698431365
transform 1 0 15000 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_949
timestamp 1698431365
transform 1 0 15000 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_950
timestamp 1698431365
transform 1 0 15600 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_951
timestamp 1698431365
transform 1 0 15600 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_952
timestamp 1698431365
transform 1 0 13800 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_953
timestamp 1698431365
transform 1 0 13800 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_954
timestamp 1698431365
transform 1 0 14400 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_955
timestamp 1698431365
transform 1 0 14400 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_956
timestamp 1698431365
transform 1 0 12600 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_957
timestamp 1698431365
transform 1 0 12600 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_958
timestamp 1698431365
transform 1 0 13200 0 1 41400
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_959
timestamp 1698431365
transform 1 0 13200 0 1 43200
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_960
timestamp 1698431365
transform -1 0 18000 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_961
timestamp 1698431365
transform -1 0 18000 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_962
timestamp 1698431365
transform -1 0 17400 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_963
timestamp 1698431365
transform -1 0 17400 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_964
timestamp 1698431365
transform -1 0 7200 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_965
timestamp 1698431365
transform -1 0 7200 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_966
timestamp 1698431365
transform -1 0 6600 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_967
timestamp 1698431365
transform -1 0 6600 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_968
timestamp 1698431365
transform -1 0 9600 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_969
timestamp 1698431365
transform -1 0 9600 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_970
timestamp 1698431365
transform -1 0 9000 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_971
timestamp 1698431365
transform -1 0 9000 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_972
timestamp 1698431365
transform -1 0 8400 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_973
timestamp 1698431365
transform -1 0 8400 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_974
timestamp 1698431365
transform -1 0 7800 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_975
timestamp 1698431365
transform -1 0 7800 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_976
timestamp 1698431365
transform -1 0 10800 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_977
timestamp 1698431365
transform -1 0 10800 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_978
timestamp 1698431365
transform -1 0 10200 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_979
timestamp 1698431365
transform -1 0 10200 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_980
timestamp 1698431365
transform -1 0 21600 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_981
timestamp 1698431365
transform -1 0 21600 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_982
timestamp 1698431365
transform -1 0 21000 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_983
timestamp 1698431365
transform -1 0 21000 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_984
timestamp 1698431365
transform -1 0 19200 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_985
timestamp 1698431365
transform -1 0 19200 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_986
timestamp 1698431365
transform -1 0 18600 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_987
timestamp 1698431365
transform -1 0 18600 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_988
timestamp 1698431365
transform -1 0 20400 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_989
timestamp 1698431365
transform -1 0 20400 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_990
timestamp 1698431365
transform -1 0 19800 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_991
timestamp 1698431365
transform -1 0 19800 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_992
timestamp 1698431365
transform 1 0 1800 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_993
timestamp 1698431365
transform 1 0 1800 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_994
timestamp 1698431365
transform 1 0 2400 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_995
timestamp 1698431365
transform 1 0 2400 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_996
timestamp 1698431365
transform 1 0 4200 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_997
timestamp 1698431365
transform 1 0 4200 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_998
timestamp 1698431365
transform 1 0 4800 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_999
timestamp 1698431365
transform 1 0 4800 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1000
timestamp 1698431365
transform 1 0 3000 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1001
timestamp 1698431365
transform 1 0 3000 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1002
timestamp 1698431365
transform 1 0 3600 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1003
timestamp 1698431365
transform 1 0 3600 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1004
timestamp 1698431365
transform 1 0 600 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1005
timestamp 1698431365
transform 1 0 600 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1006
timestamp 1698431365
transform 1 0 1200 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1007
timestamp 1698431365
transform 1 0 1200 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1008
timestamp 1698431365
transform 1 0 15000 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1009
timestamp 1698431365
transform 1 0 15000 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1010
timestamp 1698431365
transform 1 0 15600 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1011
timestamp 1698431365
transform 1 0 15600 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1012
timestamp 1698431365
transform 1 0 13800 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1013
timestamp 1698431365
transform 1 0 13800 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1014
timestamp 1698431365
transform 1 0 14400 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1015
timestamp 1698431365
transform 1 0 14400 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1016
timestamp 1698431365
transform 1 0 12600 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1017
timestamp 1698431365
transform 1 0 12600 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1018
timestamp 1698431365
transform 1 0 13200 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1019
timestamp 1698431365
transform 1 0 13200 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1020
timestamp 1698431365
transform 1 0 11400 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1021
timestamp 1698431365
transform 1 0 11400 0 1 28800
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1022
timestamp 1698431365
transform 1 0 12000 0 1 27000
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1023
timestamp 1698431365
transform 1 0 12000 0 1 28800
box -68 -68 668 1868
use 018SRAM_strap1_2x_512x8m81  018SRAM_strap1_2x_512x8m81_0
array 0 0 0 0 31 1800
timestamp 1698431365
transform -1 0 16800 0 1 900
box -68 -968 668 968
use 018SRAM_strap1_2x_512x8m81  018SRAM_strap1_2x_512x8m81_1
array 0 0 0 0 31 1800
timestamp 1698431365
transform -1 0 11400 0 1 900
box -68 -968 668 968
use 018SRAM_strap1_2x_512x8m81  018SRAM_strap1_2x_512x8m81_2
array 0 0 0 0 31 1800
timestamp 1698431365
transform -1 0 6000 0 1 900
box -68 -968 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_0
timestamp 1698431365
transform 1 0 21600 0 1 9900
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_1
timestamp 1698431365
transform 1 0 21600 0 -1 13500
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_2
timestamp 1698431365
transform 1 0 21600 0 -1 11700
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_3
timestamp 1698431365
transform 1 0 21600 0 -1 9900
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_4
timestamp 1698431365
transform 1 0 21600 0 -1 8100
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_5
timestamp 1698431365
transform 1 0 21600 0 -1 6300
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_6
timestamp 1698431365
transform 1 0 21600 0 -1 4500
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_7
timestamp 1698431365
transform 1 0 21600 0 -1 2700
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_8
timestamp 1698431365
transform 1 0 21600 0 -1 900
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_9
timestamp 1698431365
transform 1 0 21600 0 1 900
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_10
timestamp 1698431365
transform 1 0 21600 0 1 2700
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_11
timestamp 1698431365
transform 1 0 21600 0 1 4500
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_12
timestamp 1698431365
transform 1 0 21600 0 1 6300
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_13
timestamp 1698431365
transform 1 0 21600 0 1 11700
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_14
timestamp 1698431365
transform 1 0 21600 0 1 8100
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_15
timestamp 1698431365
transform 1 0 21600 0 1 15300
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_16
timestamp 1698431365
transform 1 0 21600 0 1 17100
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_17
timestamp 1698431365
transform 1 0 21600 0 1 18900
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_18
timestamp 1698431365
transform 1 0 21600 0 1 20700
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_19
timestamp 1698431365
transform 1 0 21600 0 1 22500
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_20
timestamp 1698431365
transform 1 0 21600 0 1 24300
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_21
timestamp 1698431365
transform 1 0 21600 0 1 26100
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_22
timestamp 1698431365
transform 1 0 21600 0 -1 27900
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_23
timestamp 1698431365
transform 1 0 21600 0 -1 26100
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_24
timestamp 1698431365
transform 1 0 21600 0 -1 24300
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_25
timestamp 1698431365
transform 1 0 21600 0 -1 22500
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_26
timestamp 1698431365
transform 1 0 21600 0 -1 20700
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_27
timestamp 1698431365
transform 1 0 21600 0 -1 18900
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_28
timestamp 1698431365
transform 1 0 21600 0 -1 17100
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_29
timestamp 1698431365
transform 1 0 21600 0 1 13500
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_30
timestamp 1698431365
transform 1 0 21600 0 -1 15300
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_31
timestamp 1698431365
transform -1 0 600 0 -1 8100
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_32
timestamp 1698431365
transform -1 0 600 0 -1 6300
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_33
timestamp 1698431365
transform -1 0 600 0 -1 4500
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_34
timestamp 1698431365
transform -1 0 600 0 -1 2700
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_35
timestamp 1698431365
transform -1 0 600 0 -1 900
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_36
timestamp 1698431365
transform -1 0 600 0 1 900
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_37
timestamp 1698431365
transform -1 0 600 0 1 2700
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_38
timestamp 1698431365
transform -1 0 600 0 1 4500
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_39
timestamp 1698431365
transform -1 0 600 0 1 6300
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_40
timestamp 1698431365
transform -1 0 600 0 1 8100
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_41
timestamp 1698431365
transform -1 0 600 0 1 9900
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_42
timestamp 1698431365
transform -1 0 600 0 1 11700
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_43
timestamp 1698431365
transform -1 0 600 0 -1 13500
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_44
timestamp 1698431365
transform -1 0 600 0 -1 11700
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_45
timestamp 1698431365
transform -1 0 600 0 -1 9900
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_46
timestamp 1698431365
transform -1 0 600 0 1 24300
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_47
timestamp 1698431365
transform -1 0 600 0 1 26100
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_48
timestamp 1698431365
transform -1 0 600 0 -1 27900
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_49
timestamp 1698431365
transform -1 0 600 0 -1 26100
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_50
timestamp 1698431365
transform -1 0 600 0 1 15300
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_51
timestamp 1698431365
transform -1 0 600 0 1 17100
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_52
timestamp 1698431365
transform -1 0 600 0 1 18900
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_53
timestamp 1698431365
transform -1 0 600 0 1 20700
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_54
timestamp 1698431365
transform -1 0 600 0 1 22500
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_55
timestamp 1698431365
transform -1 0 600 0 -1 24300
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_56
timestamp 1698431365
transform -1 0 600 0 -1 22500
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_57
timestamp 1698431365
transform -1 0 600 0 -1 20700
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_58
timestamp 1698431365
transform -1 0 600 0 -1 18900
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_59
timestamp 1698431365
transform -1 0 600 0 -1 17100
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_60
timestamp 1698431365
transform -1 0 600 0 1 13500
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_61
timestamp 1698431365
transform -1 0 600 0 -1 15300
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_62
timestamp 1698431365
transform -1 0 600 0 1 31500
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_63
timestamp 1698431365
transform -1 0 600 0 1 33300
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_64
timestamp 1698431365
transform -1 0 600 0 1 35100
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_65
timestamp 1698431365
transform -1 0 600 0 -1 33300
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_66
timestamp 1698431365
transform -1 0 600 0 -1 31500
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_67
timestamp 1698431365
transform -1 0 600 0 1 29700
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_68
timestamp 1698431365
transform -1 0 600 0 -1 42300
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_69
timestamp 1698431365
transform -1 0 600 0 -1 40500
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_70
timestamp 1698431365
transform -1 0 600 0 -1 38700
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_71
timestamp 1698431365
transform -1 0 600 0 1 36900
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_72
timestamp 1698431365
transform -1 0 600 0 1 38700
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_73
timestamp 1698431365
transform -1 0 600 0 1 40500
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_74
timestamp 1698431365
transform -1 0 600 0 -1 36900
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_75
timestamp 1698431365
transform -1 0 600 0 -1 35100
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_76
timestamp 1698431365
transform -1 0 600 0 1 54900
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_77
timestamp 1698431365
transform -1 0 600 0 1 56700
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_78
timestamp 1698431365
transform -1 0 600 0 -1 49500
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_79
timestamp 1698431365
transform -1 0 600 0 -1 47700
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_80
timestamp 1698431365
transform -1 0 600 0 -1 54900
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_81
timestamp 1698431365
transform -1 0 600 0 -1 53100
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_82
timestamp 1698431365
transform -1 0 600 0 -1 45900
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_83
timestamp 1698431365
transform -1 0 600 0 -1 56700
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_84
timestamp 1698431365
transform -1 0 600 0 1 44100
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_85
timestamp 1698431365
transform -1 0 600 0 1 45900
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_86
timestamp 1698431365
transform -1 0 600 0 1 47700
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_87
timestamp 1698431365
transform -1 0 600 0 1 49500
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_88
timestamp 1698431365
transform -1 0 600 0 1 51300
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_89
timestamp 1698431365
transform -1 0 600 0 1 53100
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_90
timestamp 1698431365
transform -1 0 600 0 -1 51300
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_91
timestamp 1698431365
transform -1 0 600 0 1 42300
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_92
timestamp 1698431365
transform -1 0 600 0 -1 44100
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_93
timestamp 1698431365
transform 1 0 21600 0 1 35100
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_94
timestamp 1698431365
transform 1 0 21600 0 -1 40500
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_95
timestamp 1698431365
transform 1 0 21600 0 -1 38700
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_96
timestamp 1698431365
transform 1 0 21600 0 -1 36900
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_97
timestamp 1698431365
transform 1 0 21600 0 1 36900
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_98
timestamp 1698431365
transform 1 0 21600 0 -1 35100
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_99
timestamp 1698431365
transform 1 0 21600 0 -1 42300
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_100
timestamp 1698431365
transform 1 0 21600 0 -1 33300
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_101
timestamp 1698431365
transform 1 0 21600 0 -1 31500
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_102
timestamp 1698431365
transform 1 0 21600 0 1 31500
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_103
timestamp 1698431365
transform 1 0 21600 0 1 33300
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_104
timestamp 1698431365
transform 1 0 21600 0 1 29700
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_105
timestamp 1698431365
transform 1 0 21600 0 1 38700
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_106
timestamp 1698431365
transform 1 0 21600 0 1 40500
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_107
timestamp 1698431365
transform 1 0 21600 0 1 56700
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_108
timestamp 1698431365
transform 1 0 21600 0 1 44100
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_109
timestamp 1698431365
transform 1 0 21600 0 1 45900
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_110
timestamp 1698431365
transform 1 0 21600 0 1 47700
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_111
timestamp 1698431365
transform 1 0 21600 0 1 49500
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_112
timestamp 1698431365
transform 1 0 21600 0 1 51300
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_113
timestamp 1698431365
transform 1 0 21600 0 -1 56700
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_114
timestamp 1698431365
transform 1 0 21600 0 -1 54900
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_115
timestamp 1698431365
transform 1 0 21600 0 -1 53100
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_116
timestamp 1698431365
transform 1 0 21600 0 -1 51300
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_117
timestamp 1698431365
transform 1 0 21600 0 -1 49500
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_118
timestamp 1698431365
transform 1 0 21600 0 -1 47700
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_119
timestamp 1698431365
transform 1 0 21600 0 -1 45900
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_120
timestamp 1698431365
transform 1 0 21600 0 1 54900
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_121
timestamp 1698431365
transform 1 0 21600 0 1 53100
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_122
timestamp 1698431365
transform 1 0 21600 0 1 42300
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_123
timestamp 1698431365
transform 1 0 21600 0 -1 44100
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_124
timestamp 1698431365
transform -1 0 600 0 1 27900
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_125
timestamp 1698431365
transform -1 0 600 0 -1 29700
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_126
timestamp 1698431365
transform 1 0 21600 0 -1 29700
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_127
timestamp 1698431365
transform 1 0 21600 0 1 27900
box -68 -68 668 968
<< labels >>
rlabel metal2 s 11793 231 11793 231 4 bb[7]
rlabel metal2 s 12381 231 12381 231 4 bb[6]
rlabel metal2 s 12187 231 12187 231 4 b[6]
rlabel metal2 s 12785 231 12785 231 4 b[5]
rlabel metal2 s 12978 231 12978 231 4 bb[5]
rlabel metal2 s 13595 231 13595 231 4 bb[4]
rlabel metal2 s 13402 231 13402 231 4 b[4]
rlabel metal2 s 14181 231 14181 231 4 bb[3]
rlabel metal2 s 13987 231 13987 231 4 b[3]
rlabel metal2 s 14787 231 14787 231 4 bb[2]
rlabel metal2 s 14593 231 14593 231 4 b[2]
rlabel metal2 s 15385 231 15385 231 4 bb[1]
rlabel metal2 s 15191 231 15191 231 4 b[1]
rlabel metal2 s 15983 231 15983 231 4 bb[0]
rlabel metal2 s 15789 231 15789 231 4 b[0]
rlabel metal2 s 11600 231 11600 231 4 b[7]
rlabel metal2 s 302 -20 302 -20 4 VDD
rlabel metal2 s 21898 -20 21898 -20 4 VDD
rlabel metal3 21534 53558 21534 53558 4 WL[59]
rlabel metal3 21534 54458 21534 54458 4 WL[60]
rlabel metal3 21534 55358 21534 55358 4 WL[61]
rlabel metal3 21534 50858 21534 50858 4 WL[56]
rlabel metal3 21534 56258 21534 56258 4 WL[62]
rlabel metal3 21534 57158 21534 57158 4 WL[63]
rlabel metal3 21534 51758 21534 51758 4 WL[57]
rlabel metal3 21534 52658 21534 52658 4 WL[58]
rlabel metal3 20464 50865 20464 50865 4 WL[56]
rlabel metal3 20464 51765 20464 51765 4 WL[57]
rlabel metal3 20464 52665 20464 52665 4 WL[58]
rlabel metal3 20464 53565 20464 53565 4 WL[59]
rlabel metal3 20464 54465 20464 54465 4 WL[60]
rlabel metal3 20464 55365 20464 55365 4 WL[61]
rlabel metal3 20464 56265 20464 56265 4 WL[62]
rlabel metal3 20464 57149 20464 57149 4 WL[63]
rlabel metal3 21591 57162 21591 57162 4 WL[63]
rlabel metal3 21591 56262 21591 56262 4 WL[62]
rlabel metal3 21591 55362 21591 55362 4 WL[61]
rlabel metal3 21591 54462 21591 54462 4 WL[60]
rlabel metal3 21591 53562 21591 53562 4 WL[59]
rlabel metal3 21591 52662 21591 52662 4 WL[58]
rlabel metal3 21591 51762 21591 51762 4 WL[57]
rlabel metal3 21591 50862 21591 50862 4 WL[56]
rlabel metal3 20991 57162 20991 57162 4 WL[63]
rlabel metal3 20991 56262 20991 56262 4 WL[62]
rlabel metal3 20991 55362 20991 55362 4 WL[61]
rlabel metal3 20991 54462 20991 54462 4 WL[60]
rlabel metal3 20991 53562 20991 53562 4 WL[59]
rlabel metal3 20991 52662 20991 52662 4 WL[58]
rlabel metal3 20991 51762 20991 51762 4 WL[57]
rlabel metal3 20991 50862 20991 50862 4 WL[56]
rlabel metal3 19191 57162 19191 57162 4 WL[63]
rlabel metal3 19191 56262 19191 56262 4 WL[62]
rlabel metal3 19191 55362 19191 55362 4 WL[61]
rlabel metal3 19191 54462 19191 54462 4 WL[60]
rlabel metal3 19191 53562 19191 53562 4 WL[59]
rlabel metal3 19191 52662 19191 52662 4 WL[58]
rlabel metal3 19191 51762 19191 51762 4 WL[57]
rlabel metal3 19191 50862 19191 50862 4 WL[56]
rlabel metal3 19264 50865 19264 50865 4 WL[56]
rlabel metal3 19264 51765 19264 51765 4 WL[57]
rlabel metal3 19264 52665 19264 52665 4 WL[58]
rlabel metal3 19264 53565 19264 53565 4 WL[59]
rlabel metal3 19264 54465 19264 54465 4 WL[60]
rlabel metal3 19264 55365 19264 55365 4 WL[61]
rlabel metal3 19264 56265 19264 56265 4 WL[62]
rlabel metal3 19264 57149 19264 57149 4 WL[63]
rlabel metal3 20391 57162 20391 57162 4 WL[63]
rlabel metal3 20391 56262 20391 56262 4 WL[62]
rlabel metal3 20391 55362 20391 55362 4 WL[61]
rlabel metal3 20391 54462 20391 54462 4 WL[60]
rlabel metal3 20391 53562 20391 53562 4 WL[59]
rlabel metal3 20391 52662 20391 52662 4 WL[58]
rlabel metal3 20391 51762 20391 51762 4 WL[57]
rlabel metal3 20391 50862 20391 50862 4 WL[56]
rlabel metal3 19791 57162 19791 57162 4 WL[63]
rlabel metal3 19791 56262 19791 56262 4 WL[62]
rlabel metal3 19791 55362 19791 55362 4 WL[61]
rlabel metal3 19791 54462 19791 54462 4 WL[60]
rlabel metal3 19791 53562 19791 53562 4 WL[59]
rlabel metal3 19791 52662 19791 52662 4 WL[58]
rlabel metal3 19791 51762 19791 51762 4 WL[57]
rlabel metal3 19791 50862 19791 50862 4 WL[56]
rlabel metal3 17391 57162 17391 57162 4 WL[63]
rlabel metal3 16864 52665 16864 52665 4 WL[58]
rlabel metal3 16864 50865 16864 50865 4 WL[56]
rlabel metal3 17391 50862 17391 50862 4 WL[56]
rlabel metal3 17391 51762 17391 51762 4 WL[57]
rlabel metal3 17391 54462 17391 54462 4 WL[60]
rlabel metal3 16864 51765 16864 51765 4 WL[57]
rlabel metal3 16864 53565 16864 53565 4 WL[59]
rlabel metal3 18591 57162 18591 57162 4 WL[63]
rlabel metal3 18591 56262 18591 56262 4 WL[62]
rlabel metal3 18591 55362 18591 55362 4 WL[61]
rlabel metal3 18591 54462 18591 54462 4 WL[60]
rlabel metal3 18591 53562 18591 53562 4 WL[59]
rlabel metal3 18591 52662 18591 52662 4 WL[58]
rlabel metal3 18591 51762 18591 51762 4 WL[57]
rlabel metal3 18591 50862 18591 50862 4 WL[56]
rlabel metal3 17391 56262 17391 56262 4 WL[62]
rlabel metal3 17391 52662 17391 52662 4 WL[58]
rlabel metal3 17391 53562 17391 53562 4 WL[59]
rlabel metal3 17391 55362 17391 55362 4 WL[61]
rlabel metal3 17991 55362 17991 55362 4 WL[61]
rlabel metal3 17991 56262 17991 56262 4 WL[62]
rlabel metal3 17991 54462 17991 54462 4 WL[60]
rlabel metal3 17991 53562 17991 53562 4 WL[59]
rlabel metal3 17991 52662 17991 52662 4 WL[58]
rlabel metal3 17991 51762 17991 51762 4 WL[57]
rlabel metal3 17991 50862 17991 50862 4 WL[56]
rlabel metal3 17991 57162 17991 57162 4 WL[63]
rlabel metal3 16864 57149 16864 57149 4 WL[63]
rlabel metal3 16864 56265 16864 56265 4 WL[62]
rlabel metal3 16864 55365 16864 55365 4 WL[61]
rlabel metal3 16864 54465 16864 54465 4 WL[60]
rlabel metal3 18064 50865 18064 50865 4 WL[56]
rlabel metal3 18064 51765 18064 51765 4 WL[57]
rlabel metal3 18064 52665 18064 52665 4 WL[58]
rlabel metal3 18064 53565 18064 53565 4 WL[59]
rlabel metal3 18064 54465 18064 54465 4 WL[60]
rlabel metal3 18064 55365 18064 55365 4 WL[61]
rlabel metal3 18064 56265 18064 56265 4 WL[62]
rlabel metal3 18064 57149 18064 57149 4 WL[63]
rlabel metal3 17391 43662 17391 43662 4 WL[48]
rlabel metal3 17391 44562 17391 44562 4 WL[49]
rlabel metal3 17391 45462 17391 45462 4 WL[50]
rlabel metal3 17391 46362 17391 46362 4 WL[51]
rlabel metal3 16864 43665 16864 43665 4 WL[48]
rlabel metal3 16864 44565 16864 44565 4 WL[49]
rlabel metal3 16864 45465 16864 45465 4 WL[50]
rlabel metal3 16864 46365 16864 46365 4 WL[51]
rlabel metal3 18591 49962 18591 49962 4 WL[55]
rlabel metal3 18591 49062 18591 49062 4 WL[54]
rlabel metal3 18591 48162 18591 48162 4 WL[53]
rlabel metal3 18591 47262 18591 47262 4 WL[52]
rlabel metal3 18591 46362 18591 46362 4 WL[51]
rlabel metal3 18591 45462 18591 45462 4 WL[50]
rlabel metal3 18591 44562 18591 44562 4 WL[49]
rlabel metal3 18591 43662 18591 43662 4 WL[48]
rlabel metal3 18064 43665 18064 43665 4 WL[48]
rlabel metal3 18064 44565 18064 44565 4 WL[49]
rlabel metal3 18064 45465 18064 45465 4 WL[50]
rlabel metal3 18064 46365 18064 46365 4 WL[51]
rlabel metal3 18064 47265 18064 47265 4 WL[52]
rlabel metal3 18064 48165 18064 48165 4 WL[53]
rlabel metal3 18064 49065 18064 49065 4 WL[54]
rlabel metal3 18064 49965 18064 49965 4 WL[55]
rlabel metal3 17391 47262 17391 47262 4 WL[52]
rlabel metal3 17991 49062 17991 49062 4 WL[54]
rlabel metal3 17991 48162 17991 48162 4 WL[53]
rlabel metal3 16864 49965 16864 49965 4 WL[55]
rlabel metal3 17391 48162 17391 48162 4 WL[53]
rlabel metal3 17991 47262 17991 47262 4 WL[52]
rlabel metal3 17391 49062 17391 49062 4 WL[54]
rlabel metal3 17391 49962 17391 49962 4 WL[55]
rlabel metal3 17991 44562 17991 44562 4 WL[49]
rlabel metal3 17991 43662 17991 43662 4 WL[48]
rlabel metal3 17991 46362 17991 46362 4 WL[51]
rlabel metal3 16864 49065 16864 49065 4 WL[54]
rlabel metal3 16864 48165 16864 48165 4 WL[53]
rlabel metal3 16864 47265 16864 47265 4 WL[52]
rlabel metal3 17991 49962 17991 49962 4 WL[55]
rlabel metal3 17991 45462 17991 45462 4 WL[50]
rlabel metal3 20991 49962 20991 49962 4 WL[55]
rlabel metal3 20991 49062 20991 49062 4 WL[54]
rlabel metal3 20991 48162 20991 48162 4 WL[53]
rlabel metal3 20991 47262 20991 47262 4 WL[52]
rlabel metal3 20991 46362 20991 46362 4 WL[51]
rlabel metal3 20991 45462 20991 45462 4 WL[50]
rlabel metal3 20991 44562 20991 44562 4 WL[49]
rlabel metal3 20991 43662 20991 43662 4 WL[48]
rlabel metal3 20464 43665 20464 43665 4 WL[48]
rlabel metal3 20464 44565 20464 44565 4 WL[49]
rlabel metal3 20464 45465 20464 45465 4 WL[50]
rlabel metal3 20464 46365 20464 46365 4 WL[51]
rlabel metal3 20464 47265 20464 47265 4 WL[52]
rlabel metal3 20464 48165 20464 48165 4 WL[53]
rlabel metal3 20464 49065 20464 49065 4 WL[54]
rlabel metal3 20464 49965 20464 49965 4 WL[55]
rlabel metal3 19264 43665 19264 43665 4 WL[48]
rlabel metal3 19264 44565 19264 44565 4 WL[49]
rlabel metal3 19264 45465 19264 45465 4 WL[50]
rlabel metal3 19264 46365 19264 46365 4 WL[51]
rlabel metal3 19264 47265 19264 47265 4 WL[52]
rlabel metal3 19264 48165 19264 48165 4 WL[53]
rlabel metal3 19264 49065 19264 49065 4 WL[54]
rlabel metal3 19264 49965 19264 49965 4 WL[55]
rlabel metal3 21591 49962 21591 49962 4 WL[55]
rlabel metal3 21591 49062 21591 49062 4 WL[54]
rlabel metal3 21591 48162 21591 48162 4 WL[53]
rlabel metal3 21591 47262 21591 47262 4 WL[52]
rlabel metal3 21591 46362 21591 46362 4 WL[51]
rlabel metal3 21591 45462 21591 45462 4 WL[50]
rlabel metal3 21591 44562 21591 44562 4 WL[49]
rlabel metal3 21591 43662 21591 43662 4 WL[48]
rlabel metal3 21534 43658 21534 43658 4 WL[48]
rlabel metal3 21534 48158 21534 48158 4 WL[53]
rlabel metal3 21534 46358 21534 46358 4 WL[51]
rlabel metal3 21534 49958 21534 49958 4 WL[55]
rlabel metal3 21534 47258 21534 47258 4 WL[52]
rlabel metal3 21534 49058 21534 49058 4 WL[54]
rlabel metal3 21534 44558 21534 44558 4 WL[49]
rlabel metal3 21534 45458 21534 45458 4 WL[50]
rlabel metal3 20391 49962 20391 49962 4 WL[55]
rlabel metal3 20391 49062 20391 49062 4 WL[54]
rlabel metal3 20391 48162 20391 48162 4 WL[53]
rlabel metal3 20391 47262 20391 47262 4 WL[52]
rlabel metal3 20391 46362 20391 46362 4 WL[51]
rlabel metal3 20391 45462 20391 45462 4 WL[50]
rlabel metal3 20391 44562 20391 44562 4 WL[49]
rlabel metal3 20391 43662 20391 43662 4 WL[48]
rlabel metal3 19191 49962 19191 49962 4 WL[55]
rlabel metal3 19191 49062 19191 49062 4 WL[54]
rlabel metal3 19191 48162 19191 48162 4 WL[53]
rlabel metal3 19191 47262 19191 47262 4 WL[52]
rlabel metal3 19191 46362 19191 46362 4 WL[51]
rlabel metal3 19191 45462 19191 45462 4 WL[50]
rlabel metal3 19191 44562 19191 44562 4 WL[49]
rlabel metal3 19191 43662 19191 43662 4 WL[48]
rlabel metal3 19791 49962 19791 49962 4 WL[55]
rlabel metal3 19791 49062 19791 49062 4 WL[54]
rlabel metal3 19791 48162 19791 48162 4 WL[53]
rlabel metal3 19791 47262 19791 47262 4 WL[52]
rlabel metal3 19791 46362 19791 46362 4 WL[51]
rlabel metal3 19791 45462 19791 45462 4 WL[50]
rlabel metal3 19791 44562 19791 44562 4 WL[49]
rlabel metal3 19791 43662 19791 43662 4 WL[48]
rlabel metal3 16136 50865 16136 50865 4 WL[56]
rlabel metal3 16136 51765 16136 51765 4 WL[57]
rlabel metal3 16136 52665 16136 52665 4 WL[58]
rlabel metal3 16136 53565 16136 53565 4 WL[59]
rlabel metal3 16136 54465 16136 54465 4 WL[60]
rlabel metal3 16136 55365 16136 55365 4 WL[61]
rlabel metal3 16136 56265 16136 56265 4 WL[62]
rlabel metal3 16136 57149 16136 57149 4 WL[63]
rlabel metal3 15009 57162 15009 57162 4 WL[63]
rlabel metal3 15009 56262 15009 56262 4 WL[62]
rlabel metal3 15009 55362 15009 55362 4 WL[61]
rlabel metal3 15009 54462 15009 54462 4 WL[60]
rlabel metal3 15009 53562 15009 53562 4 WL[59]
rlabel metal3 15009 52662 15009 52662 4 WL[58]
rlabel metal3 15009 51762 15009 51762 4 WL[57]
rlabel metal3 15009 50862 15009 50862 4 WL[56]
rlabel metal3 15609 57162 15609 57162 4 WL[63]
rlabel metal3 15609 56262 15609 56262 4 WL[62]
rlabel metal3 15609 55362 15609 55362 4 WL[61]
rlabel metal3 15609 54462 15609 54462 4 WL[60]
rlabel metal3 15609 53562 15609 53562 4 WL[59]
rlabel metal3 15609 52662 15609 52662 4 WL[58]
rlabel metal3 15609 51762 15609 51762 4 WL[57]
rlabel metal3 15609 50862 15609 50862 4 WL[56]
rlabel metal3 14936 50865 14936 50865 4 WL[56]
rlabel metal3 14936 51765 14936 51765 4 WL[57]
rlabel metal3 14936 52665 14936 52665 4 WL[58]
rlabel metal3 14936 53565 14936 53565 4 WL[59]
rlabel metal3 14936 54465 14936 54465 4 WL[60]
rlabel metal3 14936 55365 14936 55365 4 WL[61]
rlabel metal3 14936 56265 14936 56265 4 WL[62]
rlabel metal3 14936 57149 14936 57149 4 WL[63]
rlabel metal3 13809 57162 13809 57162 4 WL[63]
rlabel metal3 13809 56262 13809 56262 4 WL[62]
rlabel metal3 13809 55362 13809 55362 4 WL[61]
rlabel metal3 13809 54462 13809 54462 4 WL[60]
rlabel metal3 13809 53562 13809 53562 4 WL[59]
rlabel metal3 13809 52662 13809 52662 4 WL[58]
rlabel metal3 13809 51762 13809 51762 4 WL[57]
rlabel metal3 13809 50862 13809 50862 4 WL[56]
rlabel metal3 14409 57162 14409 57162 4 WL[63]
rlabel metal3 14409 56262 14409 56262 4 WL[62]
rlabel metal3 14409 55362 14409 55362 4 WL[61]
rlabel metal3 14409 54462 14409 54462 4 WL[60]
rlabel metal3 14409 53562 14409 53562 4 WL[59]
rlabel metal3 14409 52662 14409 52662 4 WL[58]
rlabel metal3 14409 51762 14409 51762 4 WL[57]
rlabel metal3 14409 50862 14409 50862 4 WL[56]
rlabel metal3 13736 50865 13736 50865 4 WL[56]
rlabel metal3 13736 51765 13736 51765 4 WL[57]
rlabel metal3 13736 52665 13736 52665 4 WL[58]
rlabel metal3 13736 53565 13736 53565 4 WL[59]
rlabel metal3 13736 54465 13736 54465 4 WL[60]
rlabel metal3 13736 55365 13736 55365 4 WL[61]
rlabel metal3 13736 56265 13736 56265 4 WL[62]
rlabel metal3 13736 57149 13736 57149 4 WL[63]
rlabel metal3 11466 50858 11466 50858 4 WL[56]
rlabel metal3 11466 51758 11466 51758 4 WL[57]
rlabel metal3 11466 52658 11466 52658 4 WL[58]
rlabel metal3 11466 53558 11466 53558 4 WL[59]
rlabel metal3 11466 54458 11466 54458 4 WL[60]
rlabel metal3 11466 55358 11466 55358 4 WL[61]
rlabel metal3 11466 56258 11466 56258 4 WL[62]
rlabel metal3 11466 57158 11466 57158 4 WL[63]
rlabel metal3 12609 57162 12609 57162 4 WL[63]
rlabel metal3 12609 56262 12609 56262 4 WL[62]
rlabel metal3 12609 55362 12609 55362 4 WL[61]
rlabel metal3 12609 54462 12609 54462 4 WL[60]
rlabel metal3 12609 53562 12609 53562 4 WL[59]
rlabel metal3 12609 52662 12609 52662 4 WL[58]
rlabel metal3 12609 51762 12609 51762 4 WL[57]
rlabel metal3 12609 50862 12609 50862 4 WL[56]
rlabel metal3 13209 57162 13209 57162 4 WL[63]
rlabel metal3 13209 56262 13209 56262 4 WL[62]
rlabel metal3 13209 55362 13209 55362 4 WL[61]
rlabel metal3 13209 54462 13209 54462 4 WL[60]
rlabel metal3 13209 53562 13209 53562 4 WL[59]
rlabel metal3 13209 52662 13209 52662 4 WL[58]
rlabel metal3 13209 51762 13209 51762 4 WL[57]
rlabel metal3 13209 50862 13209 50862 4 WL[56]
rlabel metal3 12536 50865 12536 50865 4 WL[56]
rlabel metal3 12536 51765 12536 51765 4 WL[57]
rlabel metal3 12536 52665 12536 52665 4 WL[58]
rlabel metal3 12536 53565 12536 53565 4 WL[59]
rlabel metal3 12536 54465 12536 54465 4 WL[60]
rlabel metal3 12536 55365 12536 55365 4 WL[61]
rlabel metal3 12536 56265 12536 56265 4 WL[62]
rlabel metal3 12536 57149 12536 57149 4 WL[63]
rlabel metal3 11409 57162 11409 57162 4 WL[63]
rlabel metal3 11409 56262 11409 56262 4 WL[62]
rlabel metal3 11409 55362 11409 55362 4 WL[61]
rlabel metal3 11409 54462 11409 54462 4 WL[60]
rlabel metal3 11409 53562 11409 53562 4 WL[59]
rlabel metal3 11409 52662 11409 52662 4 WL[58]
rlabel metal3 11409 51762 11409 51762 4 WL[57]
rlabel metal3 11409 50862 11409 50862 4 WL[56]
rlabel metal3 12009 57162 12009 57162 4 WL[63]
rlabel metal3 12009 56262 12009 56262 4 WL[62]
rlabel metal3 12009 55362 12009 55362 4 WL[61]
rlabel metal3 12009 54462 12009 54462 4 WL[60]
rlabel metal3 12009 53562 12009 53562 4 WL[59]
rlabel metal3 12009 52662 12009 52662 4 WL[58]
rlabel metal3 12009 51762 12009 51762 4 WL[57]
rlabel metal3 12009 50862 12009 50862 4 WL[56]
rlabel metal3 12536 43665 12536 43665 4 WL[48]
rlabel metal3 12536 44565 12536 44565 4 WL[49]
rlabel metal3 12536 45465 12536 45465 4 WL[50]
rlabel metal3 12536 46365 12536 46365 4 WL[51]
rlabel metal3 12536 47265 12536 47265 4 WL[52]
rlabel metal3 12536 48165 12536 48165 4 WL[53]
rlabel metal3 12536 49065 12536 49065 4 WL[54]
rlabel metal3 12536 49965 12536 49965 4 WL[55]
rlabel metal3 12609 49962 12609 49962 4 WL[55]
rlabel metal3 12609 49062 12609 49062 4 WL[54]
rlabel metal3 12609 48162 12609 48162 4 WL[53]
rlabel metal3 12609 47262 12609 47262 4 WL[52]
rlabel metal3 12609 46362 12609 46362 4 WL[51]
rlabel metal3 12609 45462 12609 45462 4 WL[50]
rlabel metal3 12609 44562 12609 44562 4 WL[49]
rlabel metal3 12609 43662 12609 43662 4 WL[48]
rlabel metal3 11466 43658 11466 43658 4 WL[48]
rlabel metal3 11466 44558 11466 44558 4 WL[49]
rlabel metal3 11466 45458 11466 45458 4 WL[50]
rlabel metal3 11466 46358 11466 46358 4 WL[51]
rlabel metal3 11466 47258 11466 47258 4 WL[52]
rlabel metal3 11466 48158 11466 48158 4 WL[53]
rlabel metal3 11466 49058 11466 49058 4 WL[54]
rlabel metal3 11466 49958 11466 49958 4 WL[55]
rlabel metal3 11409 49962 11409 49962 4 WL[55]
rlabel metal3 11409 49062 11409 49062 4 WL[54]
rlabel metal3 11409 48162 11409 48162 4 WL[53]
rlabel metal3 11409 47262 11409 47262 4 WL[52]
rlabel metal3 11409 46362 11409 46362 4 WL[51]
rlabel metal3 11409 45462 11409 45462 4 WL[50]
rlabel metal3 11409 44562 11409 44562 4 WL[49]
rlabel metal3 11409 43662 11409 43662 4 WL[48]
rlabel metal3 13209 49962 13209 49962 4 WL[55]
rlabel metal3 13209 49062 13209 49062 4 WL[54]
rlabel metal3 13209 48162 13209 48162 4 WL[53]
rlabel metal3 13209 47262 13209 47262 4 WL[52]
rlabel metal3 13209 46362 13209 46362 4 WL[51]
rlabel metal3 13209 45462 13209 45462 4 WL[50]
rlabel metal3 13209 44562 13209 44562 4 WL[49]
rlabel metal3 13209 43662 13209 43662 4 WL[48]
rlabel metal3 12009 49962 12009 49962 4 WL[55]
rlabel metal3 12009 49062 12009 49062 4 WL[54]
rlabel metal3 12009 48162 12009 48162 4 WL[53]
rlabel metal3 12009 47262 12009 47262 4 WL[52]
rlabel metal3 12009 46362 12009 46362 4 WL[51]
rlabel metal3 12009 45462 12009 45462 4 WL[50]
rlabel metal3 12009 44562 12009 44562 4 WL[49]
rlabel metal3 12009 43662 12009 43662 4 WL[48]
rlabel metal3 15609 49962 15609 49962 4 WL[55]
rlabel metal3 15609 49062 15609 49062 4 WL[54]
rlabel metal3 15609 48162 15609 48162 4 WL[53]
rlabel metal3 15609 47262 15609 47262 4 WL[52]
rlabel metal3 15609 46362 15609 46362 4 WL[51]
rlabel metal3 15609 45462 15609 45462 4 WL[50]
rlabel metal3 15609 44562 15609 44562 4 WL[49]
rlabel metal3 15609 43662 15609 43662 4 WL[48]
rlabel metal3 14409 49962 14409 49962 4 WL[55]
rlabel metal3 14409 49062 14409 49062 4 WL[54]
rlabel metal3 14409 48162 14409 48162 4 WL[53]
rlabel metal3 14409 47262 14409 47262 4 WL[52]
rlabel metal3 14409 46362 14409 46362 4 WL[51]
rlabel metal3 14409 45462 14409 45462 4 WL[50]
rlabel metal3 14409 44562 14409 44562 4 WL[49]
rlabel metal3 14409 43662 14409 43662 4 WL[48]
rlabel metal3 13736 43665 13736 43665 4 WL[48]
rlabel metal3 13736 44565 13736 44565 4 WL[49]
rlabel metal3 13736 45465 13736 45465 4 WL[50]
rlabel metal3 13736 46365 13736 46365 4 WL[51]
rlabel metal3 13736 47265 13736 47265 4 WL[52]
rlabel metal3 13736 48165 13736 48165 4 WL[53]
rlabel metal3 13736 49065 13736 49065 4 WL[54]
rlabel metal3 13736 49965 13736 49965 4 WL[55]
rlabel metal3 14936 43665 14936 43665 4 WL[48]
rlabel metal3 14936 44565 14936 44565 4 WL[49]
rlabel metal3 14936 45465 14936 45465 4 WL[50]
rlabel metal3 14936 46365 14936 46365 4 WL[51]
rlabel metal3 14936 47265 14936 47265 4 WL[52]
rlabel metal3 14936 48165 14936 48165 4 WL[53]
rlabel metal3 14936 49065 14936 49065 4 WL[54]
rlabel metal3 14936 49965 14936 49965 4 WL[55]
rlabel metal3 15009 49962 15009 49962 4 WL[55]
rlabel metal3 15009 49062 15009 49062 4 WL[54]
rlabel metal3 15009 48162 15009 48162 4 WL[53]
rlabel metal3 15009 47262 15009 47262 4 WL[52]
rlabel metal3 15009 46362 15009 46362 4 WL[51]
rlabel metal3 15009 45462 15009 45462 4 WL[50]
rlabel metal3 15009 44562 15009 44562 4 WL[49]
rlabel metal3 15009 43662 15009 43662 4 WL[48]
rlabel metal3 16136 43665 16136 43665 4 WL[48]
rlabel metal3 16136 44565 16136 44565 4 WL[49]
rlabel metal3 16136 45465 16136 45465 4 WL[50]
rlabel metal3 16136 46365 16136 46365 4 WL[51]
rlabel metal3 16136 47265 16136 47265 4 WL[52]
rlabel metal3 16136 48165 16136 48165 4 WL[53]
rlabel metal3 16136 49065 16136 49065 4 WL[54]
rlabel metal3 16136 49965 16136 49965 4 WL[55]
rlabel metal3 13809 49962 13809 49962 4 WL[55]
rlabel metal3 13809 49062 13809 49062 4 WL[54]
rlabel metal3 13809 48162 13809 48162 4 WL[53]
rlabel metal3 13809 47262 13809 47262 4 WL[52]
rlabel metal3 13809 46362 13809 46362 4 WL[51]
rlabel metal3 13809 45462 13809 45462 4 WL[50]
rlabel metal3 13809 44562 13809 44562 4 WL[49]
rlabel metal3 13809 43662 13809 43662 4 WL[48]
rlabel metal3 14409 42762 14409 42762 4 WL[47]
rlabel metal3 14409 41862 14409 41862 4 WL[46]
rlabel metal3 14409 40962 14409 40962 4 WL[45]
rlabel metal3 14409 40062 14409 40062 4 WL[44]
rlabel metal3 14409 39162 14409 39162 4 WL[43]
rlabel metal3 14409 38262 14409 38262 4 WL[42]
rlabel metal3 14409 37362 14409 37362 4 WL[41]
rlabel metal3 14409 36462 14409 36462 4 WL[40]
rlabel metal3 13736 36465 13736 36465 4 WL[40]
rlabel metal3 13736 37365 13736 37365 4 WL[41]
rlabel metal3 13736 38265 13736 38265 4 WL[42]
rlabel metal3 13736 39165 13736 39165 4 WL[43]
rlabel metal3 13736 40065 13736 40065 4 WL[44]
rlabel metal3 13736 40965 13736 40965 4 WL[45]
rlabel metal3 13736 41865 13736 41865 4 WL[46]
rlabel metal3 13736 42765 13736 42765 4 WL[47]
rlabel metal3 15609 42762 15609 42762 4 WL[47]
rlabel metal3 15609 41862 15609 41862 4 WL[46]
rlabel metal3 15609 40962 15609 40962 4 WL[45]
rlabel metal3 15609 40062 15609 40062 4 WL[44]
rlabel metal3 15609 39162 15609 39162 4 WL[43]
rlabel metal3 15609 38262 15609 38262 4 WL[42]
rlabel metal3 15609 37362 15609 37362 4 WL[41]
rlabel metal3 15609 36462 15609 36462 4 WL[40]
rlabel metal3 14936 36465 14936 36465 4 WL[40]
rlabel metal3 14936 37365 14936 37365 4 WL[41]
rlabel metal3 14936 38265 14936 38265 4 WL[42]
rlabel metal3 14936 39165 14936 39165 4 WL[43]
rlabel metal3 14936 40065 14936 40065 4 WL[44]
rlabel metal3 14936 40965 14936 40965 4 WL[45]
rlabel metal3 14936 41865 14936 41865 4 WL[46]
rlabel metal3 14936 42765 14936 42765 4 WL[47]
rlabel metal3 16136 36465 16136 36465 4 WL[40]
rlabel metal3 16136 37365 16136 37365 4 WL[41]
rlabel metal3 16136 38265 16136 38265 4 WL[42]
rlabel metal3 16136 39165 16136 39165 4 WL[43]
rlabel metal3 16136 40065 16136 40065 4 WL[44]
rlabel metal3 16136 40965 16136 40965 4 WL[45]
rlabel metal3 16136 41865 16136 41865 4 WL[46]
rlabel metal3 16136 42765 16136 42765 4 WL[47]
rlabel metal3 15009 42762 15009 42762 4 WL[47]
rlabel metal3 15009 41862 15009 41862 4 WL[46]
rlabel metal3 15009 40962 15009 40962 4 WL[45]
rlabel metal3 15009 40062 15009 40062 4 WL[44]
rlabel metal3 15009 39162 15009 39162 4 WL[43]
rlabel metal3 15009 38262 15009 38262 4 WL[42]
rlabel metal3 15009 37362 15009 37362 4 WL[41]
rlabel metal3 15009 36462 15009 36462 4 WL[40]
rlabel metal3 13809 42762 13809 42762 4 WL[47]
rlabel metal3 13809 41862 13809 41862 4 WL[46]
rlabel metal3 13809 40962 13809 40962 4 WL[45]
rlabel metal3 13809 40062 13809 40062 4 WL[44]
rlabel metal3 13809 39162 13809 39162 4 WL[43]
rlabel metal3 13809 38262 13809 38262 4 WL[42]
rlabel metal3 13809 37362 13809 37362 4 WL[41]
rlabel metal3 13809 36462 13809 36462 4 WL[40]
rlabel metal3 13209 38262 13209 38262 4 WL[42]
rlabel metal3 13209 37362 13209 37362 4 WL[41]
rlabel metal3 13209 36462 13209 36462 4 WL[40]
rlabel metal3 12536 36465 12536 36465 4 WL[40]
rlabel metal3 12536 37365 12536 37365 4 WL[41]
rlabel metal3 12536 38265 12536 38265 4 WL[42]
rlabel metal3 12536 39165 12536 39165 4 WL[43]
rlabel metal3 12536 40065 12536 40065 4 WL[44]
rlabel metal3 12536 40965 12536 40965 4 WL[45]
rlabel metal3 12536 41865 12536 41865 4 WL[46]
rlabel metal3 12536 42765 12536 42765 4 WL[47]
rlabel metal3 12609 39162 12609 39162 4 WL[43]
rlabel metal3 12609 38262 12609 38262 4 WL[42]
rlabel metal3 12609 37362 12609 37362 4 WL[41]
rlabel metal3 12609 36462 12609 36462 4 WL[40]
rlabel metal3 11466 42758 11466 42758 4 WL[47]
rlabel metal3 11466 39158 11466 39158 4 WL[43]
rlabel metal3 11466 40058 11466 40058 4 WL[44]
rlabel metal3 11466 40958 11466 40958 4 WL[45]
rlabel metal3 11466 41858 11466 41858 4 WL[46]
rlabel metal3 12609 42762 12609 42762 4 WL[47]
rlabel metal3 12609 41862 12609 41862 4 WL[46]
rlabel metal3 12609 40962 12609 40962 4 WL[45]
rlabel metal3 12609 40062 12609 40062 4 WL[44]
rlabel metal3 13209 42762 13209 42762 4 WL[47]
rlabel metal3 13209 41862 13209 41862 4 WL[46]
rlabel metal3 13209 40962 13209 40962 4 WL[45]
rlabel metal3 13209 40062 13209 40062 4 WL[44]
rlabel metal3 13209 39162 13209 39162 4 WL[43]
rlabel metal3 11409 42762 11409 42762 4 WL[47]
rlabel metal3 11409 41862 11409 41862 4 WL[46]
rlabel metal3 11409 40962 11409 40962 4 WL[45]
rlabel metal3 11409 40062 11409 40062 4 WL[44]
rlabel metal3 11409 39162 11409 39162 4 WL[43]
rlabel metal3 11409 38262 11409 38262 4 WL[42]
rlabel metal3 11409 37362 11409 37362 4 WL[41]
rlabel metal3 11409 36462 11409 36462 4 WL[40]
rlabel metal3 11466 36458 11466 36458 4 WL[40]
rlabel metal3 11466 37358 11466 37358 4 WL[41]
rlabel metal3 11466 38258 11466 38258 4 WL[42]
rlabel metal3 12009 42762 12009 42762 4 WL[47]
rlabel metal3 12009 41862 12009 41862 4 WL[46]
rlabel metal3 12009 40962 12009 40962 4 WL[45]
rlabel metal3 12009 40062 12009 40062 4 WL[44]
rlabel metal3 12009 39162 12009 39162 4 WL[43]
rlabel metal3 12009 38262 12009 38262 4 WL[42]
rlabel metal3 12009 37362 12009 37362 4 WL[41]
rlabel metal3 12009 36462 12009 36462 4 WL[40]
rlabel metal3 13209 31062 13209 31062 4 WL[34]
rlabel metal3 13209 30162 13209 30162 4 WL[33]
rlabel metal3 13209 29262 13209 29262 4 WL[32]
rlabel metal3 12536 34665 12536 34665 4 WL[38]
rlabel metal3 13209 35562 13209 35562 4 WL[39]
rlabel metal3 13209 34662 13209 34662 4 WL[38]
rlabel metal3 s 13266 29718 13266 29718 4 VSS
rlabel metal3 s 13266 28793 13266 28793 4 VDD
rlabel metal3 12536 35565 12536 35565 4 WL[39]
rlabel metal3 12536 29265 12536 29265 4 WL[32]
rlabel metal3 12536 30165 12536 30165 4 WL[33]
rlabel metal3 12536 31065 12536 31065 4 WL[34]
rlabel metal3 12536 31965 12536 31965 4 WL[35]
rlabel metal3 12536 32865 12536 32865 4 WL[36]
rlabel metal3 12536 33765 12536 33765 4 WL[37]
rlabel metal3 12609 31062 12609 31062 4 WL[34]
rlabel metal3 12609 30162 12609 30162 4 WL[33]
rlabel metal3 12609 29262 12609 29262 4 WL[32]
rlabel metal3 12609 35562 12609 35562 4 WL[39]
rlabel metal3 12609 34662 12609 34662 4 WL[38]
rlabel metal3 11409 33762 11409 33762 4 WL[37]
rlabel metal3 11409 32862 11409 32862 4 WL[36]
rlabel metal3 11409 31962 11409 31962 4 WL[35]
rlabel metal3 11409 31062 11409 31062 4 WL[34]
rlabel metal3 11409 30162 11409 30162 4 WL[33]
rlabel metal3 11409 29262 11409 29262 4 WL[32]
rlabel metal3 11409 35562 11409 35562 4 WL[39]
rlabel metal3 11409 34662 11409 34662 4 WL[38]
rlabel metal3 s 11466 29718 11466 29718 4 VSS
rlabel metal3 s 11466 28793 11466 28793 4 VDD
rlabel metal3 11466 34658 11466 34658 4 WL[38]
rlabel metal3 11466 35558 11466 35558 4 WL[39]
rlabel metal3 11466 31958 11466 31958 4 WL[35]
rlabel metal3 11466 32858 11466 32858 4 WL[36]
rlabel metal3 11466 33758 11466 33758 4 WL[37]
rlabel metal3 s 12666 29718 12666 29718 4 VSS
rlabel metal3 s 12666 28793 12666 28793 4 VDD
rlabel metal3 11466 29258 11466 29258 4 WL[32]
rlabel metal3 11466 30158 11466 30158 4 WL[33]
rlabel metal3 12609 33762 12609 33762 4 WL[37]
rlabel metal3 11466 31058 11466 31058 4 WL[34]
rlabel metal3 12609 32862 12609 32862 4 WL[36]
rlabel metal3 12609 31962 12609 31962 4 WL[35]
rlabel metal3 13209 33762 13209 33762 4 WL[37]
rlabel metal3 13209 32862 13209 32862 4 WL[36]
rlabel metal3 13209 31962 13209 31962 4 WL[35]
rlabel metal3 12009 33762 12009 33762 4 WL[37]
rlabel metal3 12009 32862 12009 32862 4 WL[36]
rlabel metal3 12009 31962 12009 31962 4 WL[35]
rlabel metal3 12009 31062 12009 31062 4 WL[34]
rlabel metal3 12009 30162 12009 30162 4 WL[33]
rlabel metal3 12009 29262 12009 29262 4 WL[32]
rlabel metal3 12009 35562 12009 35562 4 WL[39]
rlabel metal3 12009 34662 12009 34662 4 WL[38]
rlabel metal3 s 12066 29718 12066 29718 4 VSS
rlabel metal3 s 12066 28793 12066 28793 4 VDD
rlabel metal3 14936 32865 14936 32865 4 WL[36]
rlabel metal3 14936 33765 14936 33765 4 WL[37]
rlabel metal3 14409 33762 14409 33762 4 WL[37]
rlabel metal3 14409 32862 14409 32862 4 WL[36]
rlabel metal3 14409 31962 14409 31962 4 WL[35]
rlabel metal3 14409 31062 14409 31062 4 WL[34]
rlabel metal3 14409 30162 14409 30162 4 WL[33]
rlabel metal3 14409 29262 14409 29262 4 WL[32]
rlabel metal3 13809 33762 13809 33762 4 WL[37]
rlabel metal3 13809 32862 13809 32862 4 WL[36]
rlabel metal3 13809 31962 13809 31962 4 WL[35]
rlabel metal3 13809 31062 13809 31062 4 WL[34]
rlabel metal3 14409 35562 14409 35562 4 WL[39]
rlabel metal3 14409 34662 14409 34662 4 WL[38]
rlabel metal3 s 14466 29718 14466 29718 4 VSS
rlabel metal3 16136 34665 16136 34665 4 WL[38]
rlabel metal3 s 14466 28793 14466 28793 4 VDD
rlabel metal3 13736 35565 13736 35565 4 WL[39]
rlabel metal3 13736 29265 13736 29265 4 WL[32]
rlabel metal3 13736 30165 13736 30165 4 WL[33]
rlabel metal3 13736 31065 13736 31065 4 WL[34]
rlabel metal3 13736 31965 13736 31965 4 WL[35]
rlabel metal3 13736 32865 13736 32865 4 WL[36]
rlabel metal3 13736 33765 13736 33765 4 WL[37]
rlabel metal3 15609 33762 15609 33762 4 WL[37]
rlabel metal3 15609 32862 15609 32862 4 WL[36]
rlabel metal3 15609 31962 15609 31962 4 WL[35]
rlabel metal3 15609 31062 15609 31062 4 WL[34]
rlabel metal3 15609 30162 15609 30162 4 WL[33]
rlabel metal3 15609 29262 15609 29262 4 WL[32]
rlabel metal3 13809 30162 13809 30162 4 WL[33]
rlabel metal3 13809 29262 13809 29262 4 WL[32]
rlabel metal3 13809 35562 13809 35562 4 WL[39]
rlabel metal3 13809 34662 13809 34662 4 WL[38]
rlabel metal3 s 13866 29718 13866 29718 4 VSS
rlabel metal3 s 13866 28793 13866 28793 4 VDD
rlabel metal3 s 15066 29718 15066 29718 4 VSS
rlabel metal3 s 15066 28793 15066 28793 4 VDD
rlabel metal3 13736 34665 13736 34665 4 WL[38]
rlabel metal3 15609 35562 15609 35562 4 WL[39]
rlabel metal3 16136 35565 16136 35565 4 WL[39]
rlabel metal3 16136 29265 16136 29265 4 WL[32]
rlabel metal3 16136 30165 16136 30165 4 WL[33]
rlabel metal3 16136 31065 16136 31065 4 WL[34]
rlabel metal3 16136 31965 16136 31965 4 WL[35]
rlabel metal3 16136 32865 16136 32865 4 WL[36]
rlabel metal3 14936 34665 14936 34665 4 WL[38]
rlabel metal3 16136 33765 16136 33765 4 WL[37]
rlabel metal3 15609 34662 15609 34662 4 WL[38]
rlabel metal3 s 15666 29718 15666 29718 4 VSS
rlabel metal3 s 15666 28793 15666 28793 4 VDD
rlabel metal3 14936 35565 14936 35565 4 WL[39]
rlabel metal3 14936 29265 14936 29265 4 WL[32]
rlabel metal3 14936 30165 14936 30165 4 WL[33]
rlabel metal3 14936 31065 14936 31065 4 WL[34]
rlabel metal3 15009 33762 15009 33762 4 WL[37]
rlabel metal3 15009 32862 15009 32862 4 WL[36]
rlabel metal3 15009 31962 15009 31962 4 WL[35]
rlabel metal3 15009 31062 15009 31062 4 WL[34]
rlabel metal3 14936 31965 14936 31965 4 WL[35]
rlabel metal3 15009 30162 15009 30162 4 WL[33]
rlabel metal3 15009 29262 15009 29262 4 WL[32]
rlabel metal3 15009 35562 15009 35562 4 WL[39]
rlabel metal3 15009 34662 15009 34662 4 WL[38]
rlabel metal3 19791 40962 19791 40962 4 WL[45]
rlabel metal3 19791 40062 19791 40062 4 WL[44]
rlabel metal3 19791 39162 19791 39162 4 WL[43]
rlabel metal3 19791 38262 19791 38262 4 WL[42]
rlabel metal3 19791 37362 19791 37362 4 WL[41]
rlabel metal3 19791 36462 19791 36462 4 WL[40]
rlabel metal3 21534 38258 21534 38258 4 WL[42]
rlabel metal3 20991 42762 20991 42762 4 WL[47]
rlabel metal3 20991 41862 20991 41862 4 WL[46]
rlabel metal3 20991 40962 20991 40962 4 WL[45]
rlabel metal3 20991 40062 20991 40062 4 WL[44]
rlabel metal3 20991 39162 20991 39162 4 WL[43]
rlabel metal3 20991 38262 20991 38262 4 WL[42]
rlabel metal3 20991 37362 20991 37362 4 WL[41]
rlabel metal3 20991 36462 20991 36462 4 WL[40]
rlabel metal3 21534 40058 21534 40058 4 WL[44]
rlabel metal3 21534 42758 21534 42758 4 WL[47]
rlabel metal3 20464 36465 20464 36465 4 WL[40]
rlabel metal3 20464 37365 20464 37365 4 WL[41]
rlabel metal3 20464 38265 20464 38265 4 WL[42]
rlabel metal3 20464 39165 20464 39165 4 WL[43]
rlabel metal3 20464 40065 20464 40065 4 WL[44]
rlabel metal3 19191 42762 19191 42762 4 WL[47]
rlabel metal3 19191 41862 19191 41862 4 WL[46]
rlabel metal3 19191 40962 19191 40962 4 WL[45]
rlabel metal3 19191 40062 19191 40062 4 WL[44]
rlabel metal3 19191 39162 19191 39162 4 WL[43]
rlabel metal3 19191 38262 19191 38262 4 WL[42]
rlabel metal3 19191 37362 19191 37362 4 WL[41]
rlabel metal3 19191 36462 19191 36462 4 WL[40]
rlabel metal3 20464 40965 20464 40965 4 WL[45]
rlabel metal3 20464 41865 20464 41865 4 WL[46]
rlabel metal3 20464 42765 20464 42765 4 WL[47]
rlabel metal3 21534 36458 21534 36458 4 WL[40]
rlabel metal3 19264 36465 19264 36465 4 WL[40]
rlabel metal3 19264 37365 19264 37365 4 WL[41]
rlabel metal3 19264 38265 19264 38265 4 WL[42]
rlabel metal3 19264 39165 19264 39165 4 WL[43]
rlabel metal3 19264 40065 19264 40065 4 WL[44]
rlabel metal3 19264 40965 19264 40965 4 WL[45]
rlabel metal3 19264 41865 19264 41865 4 WL[46]
rlabel metal3 19264 42765 19264 42765 4 WL[47]
rlabel metal3 21534 41858 21534 41858 4 WL[46]
rlabel metal3 21534 40958 21534 40958 4 WL[45]
rlabel metal3 21534 37358 21534 37358 4 WL[41]
rlabel metal3 21534 39158 21534 39158 4 WL[43]
rlabel metal3 21591 42762 21591 42762 4 WL[47]
rlabel metal3 21591 41862 21591 41862 4 WL[46]
rlabel metal3 21591 40962 21591 40962 4 WL[45]
rlabel metal3 21591 40062 21591 40062 4 WL[44]
rlabel metal3 21591 39162 21591 39162 4 WL[43]
rlabel metal3 21591 38262 21591 38262 4 WL[42]
rlabel metal3 21591 37362 21591 37362 4 WL[41]
rlabel metal3 21591 36462 21591 36462 4 WL[40]
rlabel metal3 20391 42762 20391 42762 4 WL[47]
rlabel metal3 20391 41862 20391 41862 4 WL[46]
rlabel metal3 20391 40962 20391 40962 4 WL[45]
rlabel metal3 20391 40062 20391 40062 4 WL[44]
rlabel metal3 20391 39162 20391 39162 4 WL[43]
rlabel metal3 20391 38262 20391 38262 4 WL[42]
rlabel metal3 20391 37362 20391 37362 4 WL[41]
rlabel metal3 20391 36462 20391 36462 4 WL[40]
rlabel metal3 19791 42762 19791 42762 4 WL[47]
rlabel metal3 19791 41862 19791 41862 4 WL[46]
rlabel metal3 18064 42765 18064 42765 4 WL[47]
rlabel metal3 17991 42762 17991 42762 4 WL[47]
rlabel metal3 16864 40965 16864 40965 4 WL[45]
rlabel metal3 16864 41865 16864 41865 4 WL[46]
rlabel metal3 16864 42765 16864 42765 4 WL[47]
rlabel metal3 17391 42762 17391 42762 4 WL[47]
rlabel metal3 18064 36465 18064 36465 4 WL[40]
rlabel metal3 17991 40962 17991 40962 4 WL[45]
rlabel metal3 18064 37365 18064 37365 4 WL[41]
rlabel metal3 18064 38265 18064 38265 4 WL[42]
rlabel metal3 18064 39165 18064 39165 4 WL[43]
rlabel metal3 17991 41862 17991 41862 4 WL[46]
rlabel metal3 16864 37365 16864 37365 4 WL[41]
rlabel metal3 16864 38265 16864 38265 4 WL[42]
rlabel metal3 16864 36465 16864 36465 4 WL[40]
rlabel metal3 17391 36462 17391 36462 4 WL[40]
rlabel metal3 17391 37362 17391 37362 4 WL[41]
rlabel metal3 17391 39162 17391 39162 4 WL[43]
rlabel metal3 17391 40062 17391 40062 4 WL[44]
rlabel metal3 17391 40962 17391 40962 4 WL[45]
rlabel metal3 16864 40065 16864 40065 4 WL[44]
rlabel metal3 18064 40065 18064 40065 4 WL[44]
rlabel metal3 18591 42762 18591 42762 4 WL[47]
rlabel metal3 18591 41862 18591 41862 4 WL[46]
rlabel metal3 18591 40962 18591 40962 4 WL[45]
rlabel metal3 18591 40062 18591 40062 4 WL[44]
rlabel metal3 18591 39162 18591 39162 4 WL[43]
rlabel metal3 18591 38262 18591 38262 4 WL[42]
rlabel metal3 18591 37362 18591 37362 4 WL[41]
rlabel metal3 18591 36462 18591 36462 4 WL[40]
rlabel metal3 16864 39165 16864 39165 4 WL[43]
rlabel metal3 17391 41862 17391 41862 4 WL[46]
rlabel metal3 17391 38262 17391 38262 4 WL[42]
rlabel metal3 17991 36462 17991 36462 4 WL[40]
rlabel metal3 17991 37362 17991 37362 4 WL[41]
rlabel metal3 17991 38262 17991 38262 4 WL[42]
rlabel metal3 17991 40062 17991 40062 4 WL[44]
rlabel metal3 17991 39162 17991 39162 4 WL[43]
rlabel metal3 18064 40965 18064 40965 4 WL[45]
rlabel metal3 18064 41865 18064 41865 4 WL[46]
rlabel metal3 16864 31965 16864 31965 4 WL[35]
rlabel metal3 16864 35565 16864 35565 4 WL[39]
rlabel metal3 17391 34662 17391 34662 4 WL[38]
rlabel metal3 18064 34665 18064 34665 4 WL[38]
rlabel metal3 17391 29262 17391 29262 4 WL[32]
rlabel metal3 16864 31065 16864 31065 4 WL[34]
rlabel metal3 16864 32865 16864 32865 4 WL[36]
rlabel metal3 16864 30165 16864 30165 4 WL[33]
rlabel metal3 17991 32862 17991 32862 4 WL[36]
rlabel metal3 17391 30162 17391 30162 4 WL[33]
rlabel metal3 17391 31062 17391 31062 4 WL[34]
rlabel metal3 17391 31962 17391 31962 4 WL[35]
rlabel metal3 17391 32862 17391 32862 4 WL[36]
rlabel metal3 17391 33762 17391 33762 4 WL[37]
rlabel metal3 s 17334 28793 17334 28793 4 VDD
rlabel metal3 17991 31062 17991 31062 4 WL[34]
rlabel metal3 s 17934 28793 17934 28793 4 VDD
rlabel metal3 18064 35565 18064 35565 4 WL[39]
rlabel metal3 18064 29265 18064 29265 4 WL[32]
rlabel metal3 18064 30165 18064 30165 4 WL[33]
rlabel metal3 18064 31065 18064 31065 4 WL[34]
rlabel metal3 18064 31965 18064 31965 4 WL[35]
rlabel metal3 17991 35562 17991 35562 4 WL[39]
rlabel metal3 17991 30162 17991 30162 4 WL[33]
rlabel metal3 16864 34665 16864 34665 4 WL[38]
rlabel metal3 17991 34662 17991 34662 4 WL[38]
rlabel metal3 18591 33762 18591 33762 4 WL[37]
rlabel metal3 18591 32862 18591 32862 4 WL[36]
rlabel metal3 18591 31962 18591 31962 4 WL[35]
rlabel metal3 18591 31062 18591 31062 4 WL[34]
rlabel metal3 18591 30162 18591 30162 4 WL[33]
rlabel metal3 18591 29262 18591 29262 4 WL[32]
rlabel metal3 18591 35562 18591 35562 4 WL[39]
rlabel metal3 18591 34662 18591 34662 4 WL[38]
rlabel metal3 s 18534 29718 18534 29718 4 VSS
rlabel metal3 s 17334 29718 17334 29718 4 VSS
rlabel metal3 s 18534 28793 18534 28793 4 VDD
rlabel metal3 16864 33765 16864 33765 4 WL[37]
rlabel metal3 18064 32865 18064 32865 4 WL[36]
rlabel metal3 16864 29265 16864 29265 4 WL[32]
rlabel metal3 18064 33765 18064 33765 4 WL[37]
rlabel metal3 s 17934 29718 17934 29718 4 VSS
rlabel metal3 17991 31962 17991 31962 4 WL[35]
rlabel metal3 17991 33762 17991 33762 4 WL[37]
rlabel metal3 17391 35562 17391 35562 4 WL[39]
rlabel metal3 17991 29262 17991 29262 4 WL[32]
rlabel metal3 19191 31062 19191 31062 4 WL[34]
rlabel metal3 19191 30162 19191 30162 4 WL[33]
rlabel metal3 19191 29262 19191 29262 4 WL[32]
rlabel metal3 19191 35562 19191 35562 4 WL[39]
rlabel metal3 19191 34662 19191 34662 4 WL[38]
rlabel metal3 s 19134 29718 19134 29718 4 VSS
rlabel metal3 s 19134 28793 19134 28793 4 VDD
rlabel metal3 19791 34662 19791 34662 4 WL[38]
rlabel metal3 20464 34665 20464 34665 4 WL[38]
rlabel metal3 s 19734 29718 19734 29718 4 VSS
rlabel metal3 s 19734 28793 19734 28793 4 VDD
rlabel metal3 21534 33758 21534 33758 4 WL[37]
rlabel metal3 21534 29258 21534 29258 4 WL[32]
rlabel metal3 21534 30158 21534 30158 4 WL[33]
rlabel metal3 19791 33762 19791 33762 4 WL[37]
rlabel metal3 19791 32862 19791 32862 4 WL[36]
rlabel metal3 19791 31962 19791 31962 4 WL[35]
rlabel metal3 21534 31958 21534 31958 4 WL[35]
rlabel metal3 21534 35558 21534 35558 4 WL[39]
rlabel metal3 19791 31062 19791 31062 4 WL[34]
rlabel metal3 20991 33762 20991 33762 4 WL[37]
rlabel metal3 19264 34665 19264 34665 4 WL[38]
rlabel metal3 20991 32862 20991 32862 4 WL[36]
rlabel metal3 21534 31058 21534 31058 4 WL[34]
rlabel metal3 20464 35565 20464 35565 4 WL[39]
rlabel metal3 20464 29265 20464 29265 4 WL[32]
rlabel metal3 20464 30165 20464 30165 4 WL[33]
rlabel metal3 20464 31065 20464 31065 4 WL[34]
rlabel metal3 20464 31965 20464 31965 4 WL[35]
rlabel metal3 20464 32865 20464 32865 4 WL[36]
rlabel metal3 20464 33765 20464 33765 4 WL[37]
rlabel metal3 20991 31962 20991 31962 4 WL[35]
rlabel metal3 20991 31062 20991 31062 4 WL[34]
rlabel metal3 20991 30162 20991 30162 4 WL[33]
rlabel metal3 21591 33762 21591 33762 4 WL[37]
rlabel metal3 21591 32862 21591 32862 4 WL[36]
rlabel metal3 21591 31962 21591 31962 4 WL[35]
rlabel metal3 21591 31062 21591 31062 4 WL[34]
rlabel metal3 20991 29262 20991 29262 4 WL[32]
rlabel metal3 20991 35562 20991 35562 4 WL[39]
rlabel metal3 20991 34662 20991 34662 4 WL[38]
rlabel metal3 21534 32858 21534 32858 4 WL[36]
rlabel metal3 21534 34658 21534 34658 4 WL[38]
rlabel metal3 s 20934 29718 20934 29718 4 VSS
rlabel metal3 s 20934 28793 20934 28793 4 VDD
rlabel metal3 19791 30162 19791 30162 4 WL[33]
rlabel metal3 20391 33762 20391 33762 4 WL[37]
rlabel metal3 20391 32862 20391 32862 4 WL[36]
rlabel metal3 20391 31962 20391 31962 4 WL[35]
rlabel metal3 20391 31062 20391 31062 4 WL[34]
rlabel metal3 20391 30162 20391 30162 4 WL[33]
rlabel metal3 20391 29262 20391 29262 4 WL[32]
rlabel metal3 20391 35562 20391 35562 4 WL[39]
rlabel metal3 20391 34662 20391 34662 4 WL[38]
rlabel metal3 s 20334 29718 20334 29718 4 VSS
rlabel metal3 s 20334 28793 20334 28793 4 VDD
rlabel metal3 21591 30162 21591 30162 4 WL[33]
rlabel metal3 21591 29262 21591 29262 4 WL[32]
rlabel metal3 21591 35562 21591 35562 4 WL[39]
rlabel metal3 21591 34662 21591 34662 4 WL[38]
rlabel metal3 s 21534 29718 21534 29718 4 VSS
rlabel metal3 s 21534 28793 21534 28793 4 VDD
rlabel metal3 19791 29262 19791 29262 4 WL[32]
rlabel metal3 19791 35562 19791 35562 4 WL[39]
rlabel metal3 19264 35565 19264 35565 4 WL[39]
rlabel metal3 19264 29265 19264 29265 4 WL[32]
rlabel metal3 19264 30165 19264 30165 4 WL[33]
rlabel metal3 19264 31065 19264 31065 4 WL[34]
rlabel metal3 19264 31965 19264 31965 4 WL[35]
rlabel metal3 19264 32865 19264 32865 4 WL[36]
rlabel metal3 19264 33765 19264 33765 4 WL[37]
rlabel metal3 19191 33762 19191 33762 4 WL[37]
rlabel metal3 19191 32862 19191 32862 4 WL[36]
rlabel metal3 19191 31962 19191 31962 4 WL[35]
rlabel metal3 10734 56258 10734 56258 4 WL[62]
rlabel metal3 9591 57162 9591 57162 4 WL[63]
rlabel metal3 9591 56262 9591 56262 4 WL[62]
rlabel metal3 9591 55362 9591 55362 4 WL[61]
rlabel metal3 9591 54462 9591 54462 4 WL[60]
rlabel metal3 9591 53562 9591 53562 4 WL[59]
rlabel metal3 9591 52662 9591 52662 4 WL[58]
rlabel metal3 9591 51762 9591 51762 4 WL[57]
rlabel metal3 9591 50862 9591 50862 4 WL[56]
rlabel metal3 8991 57162 8991 57162 4 WL[63]
rlabel metal3 8991 56262 8991 56262 4 WL[62]
rlabel metal3 8991 55362 8991 55362 4 WL[61]
rlabel metal3 8991 54462 8991 54462 4 WL[60]
rlabel metal3 8991 53562 8991 53562 4 WL[59]
rlabel metal3 8991 52662 8991 52662 4 WL[58]
rlabel metal3 8991 51762 8991 51762 4 WL[57]
rlabel metal3 8991 50862 8991 50862 4 WL[56]
rlabel metal3 9664 50865 9664 50865 4 WL[56]
rlabel metal3 9664 51765 9664 51765 4 WL[57]
rlabel metal3 9664 52665 9664 52665 4 WL[58]
rlabel metal3 9664 53565 9664 53565 4 WL[59]
rlabel metal3 9664 54465 9664 54465 4 WL[60]
rlabel metal3 9664 55365 9664 55365 4 WL[61]
rlabel metal3 9664 56265 9664 56265 4 WL[62]
rlabel metal3 9664 57149 9664 57149 4 WL[63]
rlabel metal3 10791 57162 10791 57162 4 WL[63]
rlabel metal3 10791 56262 10791 56262 4 WL[62]
rlabel metal3 10791 55362 10791 55362 4 WL[61]
rlabel metal3 10791 54462 10791 54462 4 WL[60]
rlabel metal3 10791 53562 10791 53562 4 WL[59]
rlabel metal3 10791 52662 10791 52662 4 WL[58]
rlabel metal3 10791 51762 10791 51762 4 WL[57]
rlabel metal3 10791 50862 10791 50862 4 WL[56]
rlabel metal3 10191 57162 10191 57162 4 WL[63]
rlabel metal3 10191 56262 10191 56262 4 WL[62]
rlabel metal3 10191 55362 10191 55362 4 WL[61]
rlabel metal3 10191 54462 10191 54462 4 WL[60]
rlabel metal3 10191 53562 10191 53562 4 WL[59]
rlabel metal3 10191 52662 10191 52662 4 WL[58]
rlabel metal3 10191 51762 10191 51762 4 WL[57]
rlabel metal3 10191 50862 10191 50862 4 WL[56]
rlabel metal3 10734 57158 10734 57158 4 WL[63]
rlabel metal3 10734 53558 10734 53558 4 WL[59]
rlabel metal3 10734 54458 10734 54458 4 WL[60]
rlabel metal3 10734 50858 10734 50858 4 WL[56]
rlabel metal3 10734 51758 10734 51758 4 WL[57]
rlabel metal3 10734 55358 10734 55358 4 WL[61]
rlabel metal3 10734 52658 10734 52658 4 WL[58]
rlabel metal3 7264 51765 7264 51765 4 WL[57]
rlabel metal3 7264 52665 7264 52665 4 WL[58]
rlabel metal3 7264 53565 7264 53565 4 WL[59]
rlabel metal3 7264 54465 7264 54465 4 WL[60]
rlabel metal3 7264 55365 7264 55365 4 WL[61]
rlabel metal3 7264 56265 7264 56265 4 WL[62]
rlabel metal3 7264 57149 7264 57149 4 WL[63]
rlabel metal3 8391 57162 8391 57162 4 WL[63]
rlabel metal3 8391 56262 8391 56262 4 WL[62]
rlabel metal3 8391 55362 8391 55362 4 WL[61]
rlabel metal3 8391 54462 8391 54462 4 WL[60]
rlabel metal3 8391 53562 8391 53562 4 WL[59]
rlabel metal3 8391 52662 8391 52662 4 WL[58]
rlabel metal3 8391 51762 8391 51762 4 WL[57]
rlabel metal3 8391 50862 8391 50862 4 WL[56]
rlabel metal3 7791 57162 7791 57162 4 WL[63]
rlabel metal3 7791 56262 7791 56262 4 WL[62]
rlabel metal3 7791 55362 7791 55362 4 WL[61]
rlabel metal3 7791 54462 7791 54462 4 WL[60]
rlabel metal3 7791 53562 7791 53562 4 WL[59]
rlabel metal3 7791 52662 7791 52662 4 WL[58]
rlabel metal3 7791 51762 7791 51762 4 WL[57]
rlabel metal3 7791 50862 7791 50862 4 WL[56]
rlabel metal3 6591 55362 6591 55362 4 WL[61]
rlabel metal3 6591 54462 6591 54462 4 WL[60]
rlabel metal3 6591 53562 6591 53562 4 WL[59]
rlabel metal3 6591 52662 6591 52662 4 WL[58]
rlabel metal3 6591 51762 6591 51762 4 WL[57]
rlabel metal3 6591 50862 6591 50862 4 WL[56]
rlabel metal3 8464 50865 8464 50865 4 WL[56]
rlabel metal3 8464 51765 8464 51765 4 WL[57]
rlabel metal3 8464 52665 8464 52665 4 WL[58]
rlabel metal3 8464 53565 8464 53565 4 WL[59]
rlabel metal3 8464 54465 8464 54465 4 WL[60]
rlabel metal3 8464 55365 8464 55365 4 WL[61]
rlabel metal3 8464 56265 8464 56265 4 WL[62]
rlabel metal3 8464 57149 8464 57149 4 WL[63]
rlabel metal3 6064 57149 6064 57149 4 WL[63]
rlabel metal3 6064 55365 6064 55365 4 WL[61]
rlabel metal3 6064 54465 6064 54465 4 WL[60]
rlabel metal3 6064 52665 6064 52665 4 WL[58]
rlabel metal3 6064 51765 6064 51765 4 WL[57]
rlabel metal3 6064 50865 6064 50865 4 WL[56]
rlabel metal3 7191 52662 7191 52662 4 WL[58]
rlabel metal3 7191 54462 7191 54462 4 WL[60]
rlabel metal3 7191 56262 7191 56262 4 WL[62]
rlabel metal3 7191 50862 7191 50862 4 WL[56]
rlabel metal3 6064 53565 6064 53565 4 WL[59]
rlabel metal3 7191 51762 7191 51762 4 WL[57]
rlabel metal3 7191 53562 7191 53562 4 WL[59]
rlabel metal3 7191 55362 7191 55362 4 WL[61]
rlabel metal3 7191 57162 7191 57162 4 WL[63]
rlabel metal3 6591 57162 6591 57162 4 WL[63]
rlabel metal3 6591 56262 6591 56262 4 WL[62]
rlabel metal3 6064 56265 6064 56265 4 WL[62]
rlabel metal3 7264 50865 7264 50865 4 WL[56]
rlabel metal3 8391 49062 8391 49062 4 WL[54]
rlabel metal3 8391 48162 8391 48162 4 WL[53]
rlabel metal3 8391 47262 8391 47262 4 WL[52]
rlabel metal3 8391 46362 8391 46362 4 WL[51]
rlabel metal3 8391 45462 8391 45462 4 WL[50]
rlabel metal3 8391 44562 8391 44562 4 WL[49]
rlabel metal3 8391 43662 8391 43662 4 WL[48]
rlabel metal3 7191 43662 7191 43662 4 WL[48]
rlabel metal3 7191 44562 7191 44562 4 WL[49]
rlabel metal3 7191 45462 7191 45462 4 WL[50]
rlabel metal3 7191 46362 7191 46362 4 WL[51]
rlabel metal3 7191 47262 7191 47262 4 WL[52]
rlabel metal3 7191 48162 7191 48162 4 WL[53]
rlabel metal3 7191 49062 7191 49062 4 WL[54]
rlabel metal3 7191 49962 7191 49962 4 WL[55]
rlabel metal3 7791 49962 7791 49962 4 WL[55]
rlabel metal3 7791 49062 7791 49062 4 WL[54]
rlabel metal3 7791 48162 7791 48162 4 WL[53]
rlabel metal3 7791 47262 7791 47262 4 WL[52]
rlabel metal3 7791 46362 7791 46362 4 WL[51]
rlabel metal3 7791 45462 7791 45462 4 WL[50]
rlabel metal3 7791 44562 7791 44562 4 WL[49]
rlabel metal3 7791 43662 7791 43662 4 WL[48]
rlabel metal3 6591 49962 6591 49962 4 WL[55]
rlabel metal3 6591 49062 6591 49062 4 WL[54]
rlabel metal3 6591 48162 6591 48162 4 WL[53]
rlabel metal3 6591 47262 6591 47262 4 WL[52]
rlabel metal3 6591 46362 6591 46362 4 WL[51]
rlabel metal3 6591 45462 6591 45462 4 WL[50]
rlabel metal3 6591 44562 6591 44562 4 WL[49]
rlabel metal3 6591 43662 6591 43662 4 WL[48]
rlabel metal3 7264 43665 7264 43665 4 WL[48]
rlabel metal3 7264 44565 7264 44565 4 WL[49]
rlabel metal3 7264 45465 7264 45465 4 WL[50]
rlabel metal3 7264 46365 7264 46365 4 WL[51]
rlabel metal3 7264 47265 7264 47265 4 WL[52]
rlabel metal3 7264 48165 7264 48165 4 WL[53]
rlabel metal3 7264 49065 7264 49065 4 WL[54]
rlabel metal3 7264 49965 7264 49965 4 WL[55]
rlabel metal3 8464 43665 8464 43665 4 WL[48]
rlabel metal3 8464 44565 8464 44565 4 WL[49]
rlabel metal3 8464 45465 8464 45465 4 WL[50]
rlabel metal3 8464 46365 8464 46365 4 WL[51]
rlabel metal3 8464 47265 8464 47265 4 WL[52]
rlabel metal3 8464 48165 8464 48165 4 WL[53]
rlabel metal3 8464 49065 8464 49065 4 WL[54]
rlabel metal3 8464 49965 8464 49965 4 WL[55]
rlabel metal3 6064 49965 6064 49965 4 WL[55]
rlabel metal3 6064 49065 6064 49065 4 WL[54]
rlabel metal3 6064 48165 6064 48165 4 WL[53]
rlabel metal3 6064 47265 6064 47265 4 WL[52]
rlabel metal3 6064 46365 6064 46365 4 WL[51]
rlabel metal3 6064 45465 6064 45465 4 WL[50]
rlabel metal3 6064 44565 6064 44565 4 WL[49]
rlabel metal3 6064 43665 6064 43665 4 WL[48]
rlabel metal3 8391 49962 8391 49962 4 WL[55]
rlabel metal3 8991 49062 8991 49062 4 WL[54]
rlabel metal3 8991 48162 8991 48162 4 WL[53]
rlabel metal3 8991 47262 8991 47262 4 WL[52]
rlabel metal3 8991 46362 8991 46362 4 WL[51]
rlabel metal3 8991 45462 8991 45462 4 WL[50]
rlabel metal3 8991 44562 8991 44562 4 WL[49]
rlabel metal3 8991 43662 8991 43662 4 WL[48]
rlabel metal3 10791 49962 10791 49962 4 WL[55]
rlabel metal3 10791 49062 10791 49062 4 WL[54]
rlabel metal3 10791 48162 10791 48162 4 WL[53]
rlabel metal3 10791 47262 10791 47262 4 WL[52]
rlabel metal3 10791 46362 10791 46362 4 WL[51]
rlabel metal3 10791 45462 10791 45462 4 WL[50]
rlabel metal3 10791 44562 10791 44562 4 WL[49]
rlabel metal3 10791 43662 10791 43662 4 WL[48]
rlabel metal3 9664 43665 9664 43665 4 WL[48]
rlabel metal3 9664 44565 9664 44565 4 WL[49]
rlabel metal3 9664 45465 9664 45465 4 WL[50]
rlabel metal3 9664 46365 9664 46365 4 WL[51]
rlabel metal3 9664 47265 9664 47265 4 WL[52]
rlabel metal3 9664 48165 9664 48165 4 WL[53]
rlabel metal3 9664 49065 9664 49065 4 WL[54]
rlabel metal3 9664 49965 9664 49965 4 WL[55]
rlabel metal3 10191 49962 10191 49962 4 WL[55]
rlabel metal3 10191 49062 10191 49062 4 WL[54]
rlabel metal3 10191 48162 10191 48162 4 WL[53]
rlabel metal3 10191 47262 10191 47262 4 WL[52]
rlabel metal3 10191 46362 10191 46362 4 WL[51]
rlabel metal3 10191 45462 10191 45462 4 WL[50]
rlabel metal3 10191 44562 10191 44562 4 WL[49]
rlabel metal3 10191 43662 10191 43662 4 WL[48]
rlabel metal3 9591 49962 9591 49962 4 WL[55]
rlabel metal3 9591 49062 9591 49062 4 WL[54]
rlabel metal3 9591 48162 9591 48162 4 WL[53]
rlabel metal3 10734 49958 10734 49958 4 WL[55]
rlabel metal3 10734 46358 10734 46358 4 WL[51]
rlabel metal3 9591 47262 9591 47262 4 WL[52]
rlabel metal3 9591 46362 9591 46362 4 WL[51]
rlabel metal3 10734 47258 10734 47258 4 WL[52]
rlabel metal3 10734 43658 10734 43658 4 WL[48]
rlabel metal3 10734 44558 10734 44558 4 WL[49]
rlabel metal3 10734 48158 10734 48158 4 WL[53]
rlabel metal3 9591 45462 9591 45462 4 WL[50]
rlabel metal3 9591 44562 9591 44562 4 WL[49]
rlabel metal3 9591 43662 9591 43662 4 WL[48]
rlabel metal3 10734 45458 10734 45458 4 WL[50]
rlabel metal3 10734 49058 10734 49058 4 WL[54]
rlabel metal3 8991 49962 8991 49962 4 WL[55]
rlabel metal3 4136 50865 4136 50865 4 WL[56]
rlabel metal3 4136 51765 4136 51765 4 WL[57]
rlabel metal3 4136 52665 4136 52665 4 WL[58]
rlabel metal3 4136 53565 4136 53565 4 WL[59]
rlabel metal3 4136 54465 4136 54465 4 WL[60]
rlabel metal3 4136 55365 4136 55365 4 WL[61]
rlabel metal3 4136 56265 4136 56265 4 WL[62]
rlabel metal3 4136 57149 4136 57149 4 WL[63]
rlabel metal3 5336 50865 5336 50865 4 WL[56]
rlabel metal3 5336 51765 5336 51765 4 WL[57]
rlabel metal3 5336 52665 5336 52665 4 WL[58]
rlabel metal3 5336 53565 5336 53565 4 WL[59]
rlabel metal3 5336 54465 5336 54465 4 WL[60]
rlabel metal3 5336 55365 5336 55365 4 WL[61]
rlabel metal3 5336 56265 5336 56265 4 WL[62]
rlabel metal3 5336 57149 5336 57149 4 WL[63]
rlabel metal3 4209 57162 4209 57162 4 WL[63]
rlabel metal3 4209 56262 4209 56262 4 WL[62]
rlabel metal3 4209 55362 4209 55362 4 WL[61]
rlabel metal3 4209 54462 4209 54462 4 WL[60]
rlabel metal3 4209 53562 4209 53562 4 WL[59]
rlabel metal3 4209 52662 4209 52662 4 WL[58]
rlabel metal3 4209 51762 4209 51762 4 WL[57]
rlabel metal3 4209 50862 4209 50862 4 WL[56]
rlabel metal3 4809 57162 4809 57162 4 WL[63]
rlabel metal3 4809 56262 4809 56262 4 WL[62]
rlabel metal3 4809 55362 4809 55362 4 WL[61]
rlabel metal3 4809 54462 4809 54462 4 WL[60]
rlabel metal3 4809 53562 4809 53562 4 WL[59]
rlabel metal3 4809 52662 4809 52662 4 WL[58]
rlabel metal3 4809 51762 4809 51762 4 WL[57]
rlabel metal3 4809 50862 4809 50862 4 WL[56]
rlabel metal3 3609 57162 3609 57162 4 WL[63]
rlabel metal3 3609 56262 3609 56262 4 WL[62]
rlabel metal3 3609 55362 3609 55362 4 WL[61]
rlabel metal3 3609 54462 3609 54462 4 WL[60]
rlabel metal3 3609 53562 3609 53562 4 WL[59]
rlabel metal3 3609 52662 3609 52662 4 WL[58]
rlabel metal3 3609 51762 3609 51762 4 WL[57]
rlabel metal3 3609 50862 3609 50862 4 WL[56]
rlabel metal3 3009 50862 3009 50862 4 WL[56]
rlabel metal3 2409 56262 2409 56262 4 WL[62]
rlabel metal3 2409 55362 2409 55362 4 WL[61]
rlabel metal3 2409 54462 2409 54462 4 WL[60]
rlabel metal3 2409 53562 2409 53562 4 WL[59]
rlabel metal3 2409 52662 2409 52662 4 WL[58]
rlabel metal3 2409 51762 2409 51762 4 WL[57]
rlabel metal3 2409 50862 2409 50862 4 WL[56]
rlabel metal3 666 57158 666 57158 4 WL[63]
rlabel metal3 2936 50865 2936 50865 4 WL[56]
rlabel metal3 2936 51765 2936 51765 4 WL[57]
rlabel metal3 2936 52665 2936 52665 4 WL[58]
rlabel metal3 2936 53565 2936 53565 4 WL[59]
rlabel metal3 2936 54465 2936 54465 4 WL[60]
rlabel metal3 2936 55365 2936 55365 4 WL[61]
rlabel metal3 2936 56265 2936 56265 4 WL[62]
rlabel metal3 2936 57149 2936 57149 4 WL[63]
rlabel metal3 1809 57162 1809 57162 4 WL[63]
rlabel metal3 1809 56262 1809 56262 4 WL[62]
rlabel metal3 1809 55362 1809 55362 4 WL[61]
rlabel metal3 1809 54462 1809 54462 4 WL[60]
rlabel metal3 1809 53562 1809 53562 4 WL[59]
rlabel metal3 1809 52662 1809 52662 4 WL[58]
rlabel metal3 1809 51762 1809 51762 4 WL[57]
rlabel metal3 1809 50862 1809 50862 4 WL[56]
rlabel metal3 2409 57162 2409 57162 4 WL[63]
rlabel metal3 3009 57162 3009 57162 4 WL[63]
rlabel metal3 3009 56262 3009 56262 4 WL[62]
rlabel metal3 3009 55362 3009 55362 4 WL[61]
rlabel metal3 3009 54462 3009 54462 4 WL[60]
rlabel metal3 3009 53562 3009 53562 4 WL[59]
rlabel metal3 3009 52662 3009 52662 4 WL[58]
rlabel metal3 3009 51762 3009 51762 4 WL[57]
rlabel metal3 1736 50865 1736 50865 4 WL[56]
rlabel metal3 1736 51765 1736 51765 4 WL[57]
rlabel metal3 1736 52665 1736 52665 4 WL[58]
rlabel metal3 1736 53565 1736 53565 4 WL[59]
rlabel metal3 1736 54465 1736 54465 4 WL[60]
rlabel metal3 1736 55365 1736 55365 4 WL[61]
rlabel metal3 1736 56265 1736 56265 4 WL[62]
rlabel metal3 1736 57149 1736 57149 4 WL[63]
rlabel metal3 609 57162 609 57162 4 WL[63]
rlabel metal3 609 56262 609 56262 4 WL[62]
rlabel metal3 609 55362 609 55362 4 WL[61]
rlabel metal3 609 54462 609 54462 4 WL[60]
rlabel metal3 609 53562 609 53562 4 WL[59]
rlabel metal3 609 52662 609 52662 4 WL[58]
rlabel metal3 609 51762 609 51762 4 WL[57]
rlabel metal3 609 50862 609 50862 4 WL[56]
rlabel metal3 666 52658 666 52658 4 WL[58]
rlabel metal3 666 50858 666 50858 4 WL[56]
rlabel metal3 666 51758 666 51758 4 WL[57]
rlabel metal3 666 55358 666 55358 4 WL[61]
rlabel metal3 1209 57162 1209 57162 4 WL[63]
rlabel metal3 1209 56262 1209 56262 4 WL[62]
rlabel metal3 1209 55362 1209 55362 4 WL[61]
rlabel metal3 1209 54462 1209 54462 4 WL[60]
rlabel metal3 1209 53562 1209 53562 4 WL[59]
rlabel metal3 1209 52662 1209 52662 4 WL[58]
rlabel metal3 666 53558 666 53558 4 WL[59]
rlabel metal3 1209 51762 1209 51762 4 WL[57]
rlabel metal3 1209 50862 1209 50862 4 WL[56]
rlabel metal3 666 54458 666 54458 4 WL[60]
rlabel metal3 666 56258 666 56258 4 WL[62]
rlabel metal3 3009 43662 3009 43662 4 WL[48]
rlabel metal3 2409 46362 2409 46362 4 WL[51]
rlabel metal3 2409 45462 2409 45462 4 WL[50]
rlabel metal3 2409 44562 2409 44562 4 WL[49]
rlabel metal3 2409 43662 2409 43662 4 WL[48]
rlabel metal3 1809 48162 1809 48162 4 WL[53]
rlabel metal3 666 43658 666 43658 4 WL[48]
rlabel metal3 666 44558 666 44558 4 WL[49]
rlabel metal3 2936 43665 2936 43665 4 WL[48]
rlabel metal3 1736 43665 1736 43665 4 WL[48]
rlabel metal3 1736 44565 1736 44565 4 WL[49]
rlabel metal3 1736 45465 1736 45465 4 WL[50]
rlabel metal3 1736 46365 1736 46365 4 WL[51]
rlabel metal3 1736 47265 1736 47265 4 WL[52]
rlabel metal3 1736 48165 1736 48165 4 WL[53]
rlabel metal3 1736 49065 1736 49065 4 WL[54]
rlabel metal3 1736 49965 1736 49965 4 WL[55]
rlabel metal3 3009 49962 3009 49962 4 WL[55]
rlabel metal3 2936 44565 2936 44565 4 WL[49]
rlabel metal3 2936 45465 2936 45465 4 WL[50]
rlabel metal3 2936 46365 2936 46365 4 WL[51]
rlabel metal3 2936 47265 2936 47265 4 WL[52]
rlabel metal3 2936 48165 2936 48165 4 WL[53]
rlabel metal3 2936 49065 2936 49065 4 WL[54]
rlabel metal3 2936 49965 2936 49965 4 WL[55]
rlabel metal3 1809 47262 1809 47262 4 WL[52]
rlabel metal3 1809 46362 1809 46362 4 WL[51]
rlabel metal3 1809 45462 1809 45462 4 WL[50]
rlabel metal3 1809 44562 1809 44562 4 WL[49]
rlabel metal3 1809 43662 1809 43662 4 WL[48]
rlabel metal3 1209 47262 1209 47262 4 WL[52]
rlabel metal3 1209 46362 1209 46362 4 WL[51]
rlabel metal3 1209 45462 1209 45462 4 WL[50]
rlabel metal3 609 49962 609 49962 4 WL[55]
rlabel metal3 666 49058 666 49058 4 WL[54]
rlabel metal3 1209 44562 1209 44562 4 WL[49]
rlabel metal3 609 49062 609 49062 4 WL[54]
rlabel metal3 666 49958 666 49958 4 WL[55]
rlabel metal3 1209 43662 1209 43662 4 WL[48]
rlabel metal3 1209 48162 1209 48162 4 WL[53]
rlabel metal3 1809 49962 1809 49962 4 WL[55]
rlabel metal3 666 45458 666 45458 4 WL[50]
rlabel metal3 609 48162 609 48162 4 WL[53]
rlabel metal3 609 47262 609 47262 4 WL[52]
rlabel metal3 609 46362 609 46362 4 WL[51]
rlabel metal3 609 45462 609 45462 4 WL[50]
rlabel metal3 609 44562 609 44562 4 WL[49]
rlabel metal3 609 43662 609 43662 4 WL[48]
rlabel metal3 1809 49062 1809 49062 4 WL[54]
rlabel metal3 2409 49962 2409 49962 4 WL[55]
rlabel metal3 2409 49062 2409 49062 4 WL[54]
rlabel metal3 2409 48162 2409 48162 4 WL[53]
rlabel metal3 2409 47262 2409 47262 4 WL[52]
rlabel metal3 3009 49062 3009 49062 4 WL[54]
rlabel metal3 3009 48162 3009 48162 4 WL[53]
rlabel metal3 3009 47262 3009 47262 4 WL[52]
rlabel metal3 3009 46362 3009 46362 4 WL[51]
rlabel metal3 1209 49962 1209 49962 4 WL[55]
rlabel metal3 666 46358 666 46358 4 WL[51]
rlabel metal3 666 47258 666 47258 4 WL[52]
rlabel metal3 666 48158 666 48158 4 WL[53]
rlabel metal3 3009 45462 3009 45462 4 WL[50]
rlabel metal3 3009 44562 3009 44562 4 WL[49]
rlabel metal3 1209 49062 1209 49062 4 WL[54]
rlabel metal3 4809 44562 4809 44562 4 WL[49]
rlabel metal3 4809 43662 4809 43662 4 WL[48]
rlabel metal3 5336 43665 5336 43665 4 WL[48]
rlabel metal3 5336 44565 5336 44565 4 WL[49]
rlabel metal3 5336 45465 5336 45465 4 WL[50]
rlabel metal3 5336 46365 5336 46365 4 WL[51]
rlabel metal3 5336 47265 5336 47265 4 WL[52]
rlabel metal3 5336 48165 5336 48165 4 WL[53]
rlabel metal3 5336 49065 5336 49065 4 WL[54]
rlabel metal3 5336 49965 5336 49965 4 WL[55]
rlabel metal3 4209 49962 4209 49962 4 WL[55]
rlabel metal3 4209 49062 4209 49062 4 WL[54]
rlabel metal3 4209 48162 4209 48162 4 WL[53]
rlabel metal3 4209 47262 4209 47262 4 WL[52]
rlabel metal3 4209 46362 4209 46362 4 WL[51]
rlabel metal3 4209 45462 4209 45462 4 WL[50]
rlabel metal3 4209 44562 4209 44562 4 WL[49]
rlabel metal3 3609 49962 3609 49962 4 WL[55]
rlabel metal3 3609 49062 3609 49062 4 WL[54]
rlabel metal3 3609 48162 3609 48162 4 WL[53]
rlabel metal3 3609 47262 3609 47262 4 WL[52]
rlabel metal3 3609 46362 3609 46362 4 WL[51]
rlabel metal3 3609 45462 3609 45462 4 WL[50]
rlabel metal3 3609 44562 3609 44562 4 WL[49]
rlabel metal3 3609 43662 3609 43662 4 WL[48]
rlabel metal3 4209 43662 4209 43662 4 WL[48]
rlabel metal3 4136 44565 4136 44565 4 WL[49]
rlabel metal3 4136 45465 4136 45465 4 WL[50]
rlabel metal3 4136 46365 4136 46365 4 WL[51]
rlabel metal3 4136 47265 4136 47265 4 WL[52]
rlabel metal3 4136 48165 4136 48165 4 WL[53]
rlabel metal3 4136 49065 4136 49065 4 WL[54]
rlabel metal3 4136 49965 4136 49965 4 WL[55]
rlabel metal3 4136 43665 4136 43665 4 WL[48]
rlabel metal3 4809 49962 4809 49962 4 WL[55]
rlabel metal3 4809 49062 4809 49062 4 WL[54]
rlabel metal3 4809 48162 4809 48162 4 WL[53]
rlabel metal3 4809 47262 4809 47262 4 WL[52]
rlabel metal3 4809 46362 4809 46362 4 WL[51]
rlabel metal3 4809 45462 4809 45462 4 WL[50]
rlabel metal3 3609 42762 3609 42762 4 WL[47]
rlabel metal3 3609 41862 3609 41862 4 WL[46]
rlabel metal3 3609 40962 3609 40962 4 WL[45]
rlabel metal3 3609 40062 3609 40062 4 WL[44]
rlabel metal3 3609 39162 3609 39162 4 WL[43]
rlabel metal3 3609 38262 3609 38262 4 WL[42]
rlabel metal3 3609 37362 3609 37362 4 WL[41]
rlabel metal3 3609 36462 3609 36462 4 WL[40]
rlabel metal3 5336 36465 5336 36465 4 WL[40]
rlabel metal3 5336 37365 5336 37365 4 WL[41]
rlabel metal3 5336 38265 5336 38265 4 WL[42]
rlabel metal3 5336 39165 5336 39165 4 WL[43]
rlabel metal3 5336 40065 5336 40065 4 WL[44]
rlabel metal3 5336 40965 5336 40965 4 WL[45]
rlabel metal3 5336 41865 5336 41865 4 WL[46]
rlabel metal3 5336 42765 5336 42765 4 WL[47]
rlabel metal3 4136 36465 4136 36465 4 WL[40]
rlabel metal3 4136 37365 4136 37365 4 WL[41]
rlabel metal3 4136 38265 4136 38265 4 WL[42]
rlabel metal3 4136 39165 4136 39165 4 WL[43]
rlabel metal3 4136 40065 4136 40065 4 WL[44]
rlabel metal3 4136 40965 4136 40965 4 WL[45]
rlabel metal3 4136 41865 4136 41865 4 WL[46]
rlabel metal3 4136 42765 4136 42765 4 WL[47]
rlabel metal3 4209 42762 4209 42762 4 WL[47]
rlabel metal3 4209 41862 4209 41862 4 WL[46]
rlabel metal3 4209 40962 4209 40962 4 WL[45]
rlabel metal3 4209 40062 4209 40062 4 WL[44]
rlabel metal3 4209 39162 4209 39162 4 WL[43]
rlabel metal3 4209 38262 4209 38262 4 WL[42]
rlabel metal3 4209 37362 4209 37362 4 WL[41]
rlabel metal3 4209 36462 4209 36462 4 WL[40]
rlabel metal3 4809 42762 4809 42762 4 WL[47]
rlabel metal3 4809 41862 4809 41862 4 WL[46]
rlabel metal3 4809 40962 4809 40962 4 WL[45]
rlabel metal3 4809 40062 4809 40062 4 WL[44]
rlabel metal3 4809 39162 4809 39162 4 WL[43]
rlabel metal3 4809 38262 4809 38262 4 WL[42]
rlabel metal3 4809 37362 4809 37362 4 WL[41]
rlabel metal3 4809 36462 4809 36462 4 WL[40]
rlabel metal3 1736 38265 1736 38265 4 WL[42]
rlabel metal3 1736 39165 1736 39165 4 WL[43]
rlabel metal3 1736 40065 1736 40065 4 WL[44]
rlabel metal3 1736 40965 1736 40965 4 WL[45]
rlabel metal3 1736 41865 1736 41865 4 WL[46]
rlabel metal3 1736 42765 1736 42765 4 WL[47]
rlabel metal3 1809 42762 1809 42762 4 WL[47]
rlabel metal3 1809 41862 1809 41862 4 WL[46]
rlabel metal3 1809 40962 1809 40962 4 WL[45]
rlabel metal3 1809 40062 1809 40062 4 WL[44]
rlabel metal3 1809 39162 1809 39162 4 WL[43]
rlabel metal3 609 42762 609 42762 4 WL[47]
rlabel metal3 609 41862 609 41862 4 WL[46]
rlabel metal3 609 40962 609 40962 4 WL[45]
rlabel metal3 609 40062 609 40062 4 WL[44]
rlabel metal3 609 39162 609 39162 4 WL[43]
rlabel metal3 609 38262 609 38262 4 WL[42]
rlabel metal3 609 37362 609 37362 4 WL[41]
rlabel metal3 609 36462 609 36462 4 WL[40]
rlabel metal3 1809 38262 1809 38262 4 WL[42]
rlabel metal3 1809 37362 1809 37362 4 WL[41]
rlabel metal3 1809 36462 1809 36462 4 WL[40]
rlabel metal3 666 36458 666 36458 4 WL[40]
rlabel metal3 666 40958 666 40958 4 WL[45]
rlabel metal3 666 40058 666 40058 4 WL[44]
rlabel metal3 1736 36465 1736 36465 4 WL[40]
rlabel metal3 1736 37365 1736 37365 4 WL[41]
rlabel metal3 2936 36465 2936 36465 4 WL[40]
rlabel metal3 2936 37365 2936 37365 4 WL[41]
rlabel metal3 2936 38265 2936 38265 4 WL[42]
rlabel metal3 2936 39165 2936 39165 4 WL[43]
rlabel metal3 2936 40065 2936 40065 4 WL[44]
rlabel metal3 2936 40965 2936 40965 4 WL[45]
rlabel metal3 2936 41865 2936 41865 4 WL[46]
rlabel metal3 1209 42762 1209 42762 4 WL[47]
rlabel metal3 1209 41862 1209 41862 4 WL[46]
rlabel metal3 1209 40962 1209 40962 4 WL[45]
rlabel metal3 1209 40062 1209 40062 4 WL[44]
rlabel metal3 1209 39162 1209 39162 4 WL[43]
rlabel metal3 1209 38262 1209 38262 4 WL[42]
rlabel metal3 1209 37362 1209 37362 4 WL[41]
rlabel metal3 1209 36462 1209 36462 4 WL[40]
rlabel metal3 2936 42765 2936 42765 4 WL[47]
rlabel metal3 666 37358 666 37358 4 WL[41]
rlabel metal3 2409 42762 2409 42762 4 WL[47]
rlabel metal3 2409 41862 2409 41862 4 WL[46]
rlabel metal3 2409 40962 2409 40962 4 WL[45]
rlabel metal3 2409 40062 2409 40062 4 WL[44]
rlabel metal3 2409 39162 2409 39162 4 WL[43]
rlabel metal3 2409 38262 2409 38262 4 WL[42]
rlabel metal3 2409 37362 2409 37362 4 WL[41]
rlabel metal3 2409 36462 2409 36462 4 WL[40]
rlabel metal3 3009 42762 3009 42762 4 WL[47]
rlabel metal3 3009 41862 3009 41862 4 WL[46]
rlabel metal3 3009 40962 3009 40962 4 WL[45]
rlabel metal3 3009 40062 3009 40062 4 WL[44]
rlabel metal3 3009 39162 3009 39162 4 WL[43]
rlabel metal3 3009 38262 3009 38262 4 WL[42]
rlabel metal3 3009 37362 3009 37362 4 WL[41]
rlabel metal3 3009 36462 3009 36462 4 WL[40]
rlabel metal3 666 38258 666 38258 4 WL[42]
rlabel metal3 666 39158 666 39158 4 WL[43]
rlabel metal3 666 41858 666 41858 4 WL[46]
rlabel metal3 666 42758 666 42758 4 WL[47]
rlabel metal3 2936 32865 2936 32865 4 WL[36]
rlabel metal3 2936 33765 2936 33765 4 WL[37]
rlabel metal3 1809 31962 1809 31962 4 WL[35]
rlabel metal3 2936 34665 2936 34665 4 WL[38]
rlabel metal3 1809 31062 1809 31062 4 WL[34]
rlabel metal3 1809 29262 1809 29262 4 WL[32]
rlabel metal3 1809 35562 1809 35562 4 WL[39]
rlabel metal3 1809 34662 1809 34662 4 WL[38]
rlabel metal3 s 1866 29718 1866 29718 4 VSS
rlabel metal3 1736 34665 1736 34665 4 WL[38]
rlabel metal3 666 29258 666 29258 4 WL[32]
rlabel metal3 2936 35565 2936 35565 4 WL[39]
rlabel metal3 666 31958 666 31958 4 WL[35]
rlabel metal3 666 35558 666 35558 4 WL[39]
rlabel metal3 666 30158 666 30158 4 WL[33]
rlabel metal3 1736 35565 1736 35565 4 WL[39]
rlabel metal3 1736 29265 1736 29265 4 WL[32]
rlabel metal3 609 33762 609 33762 4 WL[37]
rlabel metal3 1209 33762 1209 33762 4 WL[37]
rlabel metal3 1209 32862 1209 32862 4 WL[36]
rlabel metal3 1209 31962 1209 31962 4 WL[35]
rlabel metal3 1209 31062 1209 31062 4 WL[34]
rlabel metal3 1209 30162 1209 30162 4 WL[33]
rlabel metal3 1209 29262 1209 29262 4 WL[32]
rlabel metal3 1209 35562 1209 35562 4 WL[39]
rlabel metal3 1209 34662 1209 34662 4 WL[38]
rlabel metal3 s 1266 29718 1266 29718 4 VSS
rlabel metal3 s 1266 28793 1266 28793 4 VDD
rlabel metal3 609 32862 609 32862 4 WL[36]
rlabel metal3 609 31962 609 31962 4 WL[35]
rlabel metal3 609 31062 609 31062 4 WL[34]
rlabel metal3 1736 30165 1736 30165 4 WL[33]
rlabel metal3 1809 30162 1809 30162 4 WL[33]
rlabel metal3 1736 31065 1736 31065 4 WL[34]
rlabel metal3 1736 31965 1736 31965 4 WL[35]
rlabel metal3 1736 32865 1736 32865 4 WL[36]
rlabel metal3 1736 33765 1736 33765 4 WL[37]
rlabel metal3 1809 33762 1809 33762 4 WL[37]
rlabel metal3 2409 33762 2409 33762 4 WL[37]
rlabel metal3 2409 32862 2409 32862 4 WL[36]
rlabel metal3 1809 32862 1809 32862 4 WL[36]
rlabel metal3 609 30162 609 30162 4 WL[33]
rlabel metal3 609 29262 609 29262 4 WL[32]
rlabel metal3 609 35562 609 35562 4 WL[39]
rlabel metal3 609 34662 609 34662 4 WL[38]
rlabel metal3 s 666 29718 666 29718 4 VSS
rlabel metal3 s 666 28793 666 28793 4 VDD
rlabel metal3 s 1866 28793 1866 28793 4 VDD
rlabel metal3 3009 33762 3009 33762 4 WL[37]
rlabel metal3 3009 32862 3009 32862 4 WL[36]
rlabel metal3 3009 31962 3009 31962 4 WL[35]
rlabel metal3 3009 31062 3009 31062 4 WL[34]
rlabel metal3 666 31058 666 31058 4 WL[34]
rlabel metal3 666 34658 666 34658 4 WL[38]
rlabel metal3 3009 30162 3009 30162 4 WL[33]
rlabel metal3 3009 29262 3009 29262 4 WL[32]
rlabel metal3 3009 35562 3009 35562 4 WL[39]
rlabel metal3 3009 34662 3009 34662 4 WL[38]
rlabel metal3 666 32858 666 32858 4 WL[36]
rlabel metal3 666 33758 666 33758 4 WL[37]
rlabel metal3 s 3066 29718 3066 29718 4 VSS
rlabel metal3 s 3066 28793 3066 28793 4 VDD
rlabel metal3 2936 29265 2936 29265 4 WL[32]
rlabel metal3 2936 30165 2936 30165 4 WL[33]
rlabel metal3 2409 31962 2409 31962 4 WL[35]
rlabel metal3 2409 31062 2409 31062 4 WL[34]
rlabel metal3 2936 31065 2936 31065 4 WL[34]
rlabel metal3 2936 31965 2936 31965 4 WL[35]
rlabel metal3 2409 30162 2409 30162 4 WL[33]
rlabel metal3 2409 29262 2409 29262 4 WL[32]
rlabel metal3 2409 35562 2409 35562 4 WL[39]
rlabel metal3 2409 34662 2409 34662 4 WL[38]
rlabel metal3 s 2466 29718 2466 29718 4 VSS
rlabel metal3 s 2466 28793 2466 28793 4 VDD
rlabel metal3 4809 30162 4809 30162 4 WL[33]
rlabel metal3 4809 29262 4809 29262 4 WL[32]
rlabel metal3 4809 35562 4809 35562 4 WL[39]
rlabel metal3 4809 34662 4809 34662 4 WL[38]
rlabel metal3 s 4866 29718 4866 29718 4 VSS
rlabel metal3 s 4866 28793 4866 28793 4 VDD
rlabel metal3 4136 35565 4136 35565 4 WL[39]
rlabel metal3 4209 33762 4209 33762 4 WL[37]
rlabel metal3 4209 32862 4209 32862 4 WL[36]
rlabel metal3 4209 31962 4209 31962 4 WL[35]
rlabel metal3 4209 31062 4209 31062 4 WL[34]
rlabel metal3 4209 30162 4209 30162 4 WL[33]
rlabel metal3 4209 29262 4209 29262 4 WL[32]
rlabel metal3 4209 35562 4209 35562 4 WL[39]
rlabel metal3 4209 34662 4209 34662 4 WL[38]
rlabel metal3 s 4266 29718 4266 29718 4 VSS
rlabel metal3 s 4266 28793 4266 28793 4 VDD
rlabel metal3 5336 34665 5336 34665 4 WL[38]
rlabel metal3 4136 29265 4136 29265 4 WL[32]
rlabel metal3 4136 30165 4136 30165 4 WL[33]
rlabel metal3 4136 31065 4136 31065 4 WL[34]
rlabel metal3 s 3666 29718 3666 29718 4 VSS
rlabel metal3 4136 31965 4136 31965 4 WL[35]
rlabel metal3 4136 34665 4136 34665 4 WL[38]
rlabel metal3 4136 32865 4136 32865 4 WL[36]
rlabel metal3 4136 33765 4136 33765 4 WL[37]
rlabel metal3 s 3666 28793 3666 28793 4 VDD
rlabel metal3 3609 33762 3609 33762 4 WL[37]
rlabel metal3 3609 32862 3609 32862 4 WL[36]
rlabel metal3 5336 35565 5336 35565 4 WL[39]
rlabel metal3 5336 29265 5336 29265 4 WL[32]
rlabel metal3 5336 30165 5336 30165 4 WL[33]
rlabel metal3 5336 31065 5336 31065 4 WL[34]
rlabel metal3 5336 31965 5336 31965 4 WL[35]
rlabel metal3 5336 32865 5336 32865 4 WL[36]
rlabel metal3 5336 33765 5336 33765 4 WL[37]
rlabel metal3 3609 31962 3609 31962 4 WL[35]
rlabel metal3 3609 31062 3609 31062 4 WL[34]
rlabel metal3 3609 30162 3609 30162 4 WL[33]
rlabel metal3 3609 29262 3609 29262 4 WL[32]
rlabel metal3 3609 35562 3609 35562 4 WL[39]
rlabel metal3 3609 34662 3609 34662 4 WL[38]
rlabel metal3 4809 33762 4809 33762 4 WL[37]
rlabel metal3 4809 32862 4809 32862 4 WL[36]
rlabel metal3 4809 31962 4809 31962 4 WL[35]
rlabel metal3 4809 31062 4809 31062 4 WL[34]
rlabel metal3 9664 36465 9664 36465 4 WL[40]
rlabel metal3 9664 37365 9664 37365 4 WL[41]
rlabel metal3 9664 38265 9664 38265 4 WL[42]
rlabel metal3 9664 39165 9664 39165 4 WL[43]
rlabel metal3 9664 40065 9664 40065 4 WL[44]
rlabel metal3 9664 40965 9664 40965 4 WL[45]
rlabel metal3 9664 41865 9664 41865 4 WL[46]
rlabel metal3 9664 42765 9664 42765 4 WL[47]
rlabel metal3 9591 42762 9591 42762 4 WL[47]
rlabel metal3 9591 41862 9591 41862 4 WL[46]
rlabel metal3 9591 40962 9591 40962 4 WL[45]
rlabel metal3 9591 40062 9591 40062 4 WL[44]
rlabel metal3 9591 39162 9591 39162 4 WL[43]
rlabel metal3 9591 38262 9591 38262 4 WL[42]
rlabel metal3 9591 37362 9591 37362 4 WL[41]
rlabel metal3 9591 36462 9591 36462 4 WL[40]
rlabel metal3 10791 42762 10791 42762 4 WL[47]
rlabel metal3 10791 41862 10791 41862 4 WL[46]
rlabel metal3 10791 40962 10791 40962 4 WL[45]
rlabel metal3 10791 40062 10791 40062 4 WL[44]
rlabel metal3 10791 39162 10791 39162 4 WL[43]
rlabel metal3 10791 38262 10791 38262 4 WL[42]
rlabel metal3 10791 37362 10791 37362 4 WL[41]
rlabel metal3 10791 36462 10791 36462 4 WL[40]
rlabel metal3 10191 42762 10191 42762 4 WL[47]
rlabel metal3 10191 41862 10191 41862 4 WL[46]
rlabel metal3 10191 40962 10191 40962 4 WL[45]
rlabel metal3 10191 40062 10191 40062 4 WL[44]
rlabel metal3 10191 39162 10191 39162 4 WL[43]
rlabel metal3 10191 38262 10191 38262 4 WL[42]
rlabel metal3 10191 37362 10191 37362 4 WL[41]
rlabel metal3 10191 36462 10191 36462 4 WL[40]
rlabel metal3 10734 36458 10734 36458 4 WL[40]
rlabel metal3 10734 42758 10734 42758 4 WL[47]
rlabel metal3 10734 39158 10734 39158 4 WL[43]
rlabel metal3 10734 40058 10734 40058 4 WL[44]
rlabel metal3 10734 37358 10734 37358 4 WL[41]
rlabel metal3 10734 40958 10734 40958 4 WL[45]
rlabel metal3 8991 42762 8991 42762 4 WL[47]
rlabel metal3 8991 41862 8991 41862 4 WL[46]
rlabel metal3 8991 40962 8991 40962 4 WL[45]
rlabel metal3 8991 40062 8991 40062 4 WL[44]
rlabel metal3 8991 39162 8991 39162 4 WL[43]
rlabel metal3 8991 38262 8991 38262 4 WL[42]
rlabel metal3 8991 37362 8991 37362 4 WL[41]
rlabel metal3 8991 36462 8991 36462 4 WL[40]
rlabel metal3 10734 38258 10734 38258 4 WL[42]
rlabel metal3 10734 41858 10734 41858 4 WL[46]
rlabel metal3 8464 38265 8464 38265 4 WL[42]
rlabel metal3 7791 42762 7791 42762 4 WL[47]
rlabel metal3 7791 41862 7791 41862 4 WL[46]
rlabel metal3 7791 40962 7791 40962 4 WL[45]
rlabel metal3 7791 40062 7791 40062 4 WL[44]
rlabel metal3 7791 39162 7791 39162 4 WL[43]
rlabel metal3 7791 38262 7791 38262 4 WL[42]
rlabel metal3 7791 37362 7791 37362 4 WL[41]
rlabel metal3 7791 36462 7791 36462 4 WL[40]
rlabel metal3 8464 39165 8464 39165 4 WL[43]
rlabel metal3 8464 40065 8464 40065 4 WL[44]
rlabel metal3 8464 40965 8464 40965 4 WL[45]
rlabel metal3 8464 41865 8464 41865 4 WL[46]
rlabel metal3 8464 42765 8464 42765 4 WL[47]
rlabel metal3 6591 39162 6591 39162 4 WL[43]
rlabel metal3 6591 38262 6591 38262 4 WL[42]
rlabel metal3 6591 37362 6591 37362 4 WL[41]
rlabel metal3 6591 36462 6591 36462 4 WL[40]
rlabel metal3 8391 42762 8391 42762 4 WL[47]
rlabel metal3 8391 41862 8391 41862 4 WL[46]
rlabel metal3 8391 40962 8391 40962 4 WL[45]
rlabel metal3 8391 40062 8391 40062 4 WL[44]
rlabel metal3 8391 39162 8391 39162 4 WL[43]
rlabel metal3 8391 38262 8391 38262 4 WL[42]
rlabel metal3 8391 37362 8391 37362 4 WL[41]
rlabel metal3 8391 36462 8391 36462 4 WL[40]
rlabel metal3 7191 37362 7191 37362 4 WL[41]
rlabel metal3 6064 37365 6064 37365 4 WL[41]
rlabel metal3 6064 39165 6064 39165 4 WL[43]
rlabel metal3 6064 41865 6064 41865 4 WL[46]
rlabel metal3 6064 38265 6064 38265 4 WL[42]
rlabel metal3 6064 36465 6064 36465 4 WL[40]
rlabel metal3 7191 36462 7191 36462 4 WL[40]
rlabel metal3 7191 38262 7191 38262 4 WL[42]
rlabel metal3 7191 39162 7191 39162 4 WL[43]
rlabel metal3 7264 36465 7264 36465 4 WL[40]
rlabel metal3 7264 37365 7264 37365 4 WL[41]
rlabel metal3 6064 42765 6064 42765 4 WL[47]
rlabel metal3 7191 40062 7191 40062 4 WL[44]
rlabel metal3 7191 40962 7191 40962 4 WL[45]
rlabel metal3 7191 41862 7191 41862 4 WL[46]
rlabel metal3 7264 38265 7264 38265 4 WL[42]
rlabel metal3 7264 39165 7264 39165 4 WL[43]
rlabel metal3 7264 40065 7264 40065 4 WL[44]
rlabel metal3 7191 42762 7191 42762 4 WL[47]
rlabel metal3 6064 40965 6064 40965 4 WL[45]
rlabel metal3 7264 40965 7264 40965 4 WL[45]
rlabel metal3 7264 41865 7264 41865 4 WL[46]
rlabel metal3 7264 42765 7264 42765 4 WL[47]
rlabel metal3 6064 40065 6064 40065 4 WL[44]
rlabel metal3 6591 42762 6591 42762 4 WL[47]
rlabel metal3 6591 41862 6591 41862 4 WL[46]
rlabel metal3 6591 40962 6591 40962 4 WL[45]
rlabel metal3 6591 40062 6591 40062 4 WL[44]
rlabel metal3 8464 36465 8464 36465 4 WL[40]
rlabel metal3 8464 37365 8464 37365 4 WL[41]
rlabel metal3 7791 31962 7791 31962 4 WL[35]
rlabel metal3 7791 31062 7791 31062 4 WL[34]
rlabel metal3 7791 30162 7791 30162 4 WL[33]
rlabel metal3 7791 29262 7791 29262 4 WL[32]
rlabel metal3 7791 35562 7791 35562 4 WL[39]
rlabel metal3 7791 34662 7791 34662 4 WL[38]
rlabel metal3 s 7734 29718 7734 29718 4 VSS
rlabel metal3 s 7734 28793 7734 28793 4 VDD
rlabel metal3 8391 31062 8391 31062 4 WL[34]
rlabel metal3 8391 30162 8391 30162 4 WL[33]
rlabel metal3 8391 29262 8391 29262 4 WL[32]
rlabel metal3 8391 35562 8391 35562 4 WL[39]
rlabel metal3 8391 34662 8391 34662 4 WL[38]
rlabel metal3 s 8334 29718 8334 29718 4 VSS
rlabel metal3 s 8334 28793 8334 28793 4 VDD
rlabel metal3 6591 34662 6591 34662 4 WL[38]
rlabel metal3 s 6534 29718 6534 29718 4 VSS
rlabel metal3 s 7134 29718 7134 29718 4 VSS
rlabel metal3 6064 34665 6064 34665 4 WL[38]
rlabel metal3 s 6534 28793 6534 28793 4 VDD
rlabel metal3 s 7134 28793 7134 28793 4 VDD
rlabel metal3 7191 35562 7191 35562 4 WL[39]
rlabel metal3 7191 34662 7191 34662 4 WL[38]
rlabel metal3 8464 34665 8464 34665 4 WL[38]
rlabel metal3 6591 31962 6591 31962 4 WL[35]
rlabel metal3 6591 31062 6591 31062 4 WL[34]
rlabel metal3 6591 30162 6591 30162 4 WL[33]
rlabel metal3 6591 29262 6591 29262 4 WL[32]
rlabel metal3 6591 35562 6591 35562 4 WL[39]
rlabel metal3 8464 33765 8464 33765 4 WL[37]
rlabel metal3 7264 32865 7264 32865 4 WL[36]
rlabel metal3 7191 29262 7191 29262 4 WL[32]
rlabel metal3 7264 33765 7264 33765 4 WL[37]
rlabel metal3 7264 34665 7264 34665 4 WL[38]
rlabel metal3 7264 30165 7264 30165 4 WL[33]
rlabel metal3 7264 31065 7264 31065 4 WL[34]
rlabel metal3 7264 31965 7264 31965 4 WL[35]
rlabel metal3 8391 33762 8391 33762 4 WL[37]
rlabel metal3 8391 32862 8391 32862 4 WL[36]
rlabel metal3 8464 35565 8464 35565 4 WL[39]
rlabel metal3 8464 29265 8464 29265 4 WL[32]
rlabel metal3 8464 30165 8464 30165 4 WL[33]
rlabel metal3 8464 31065 8464 31065 4 WL[34]
rlabel metal3 8464 31965 8464 31965 4 WL[35]
rlabel metal3 8464 32865 8464 32865 4 WL[36]
rlabel metal3 6591 33762 6591 33762 4 WL[37]
rlabel metal3 6591 32862 6591 32862 4 WL[36]
rlabel metal3 8391 31962 8391 31962 4 WL[35]
rlabel metal3 7791 33762 7791 33762 4 WL[37]
rlabel metal3 7791 32862 7791 32862 4 WL[36]
rlabel metal3 7191 33762 7191 33762 4 WL[37]
rlabel metal3 6064 33765 6064 33765 4 WL[37]
rlabel metal3 6064 32865 6064 32865 4 WL[36]
rlabel metal3 6064 31965 6064 31965 4 WL[35]
rlabel metal3 6064 31065 6064 31065 4 WL[34]
rlabel metal3 7191 32862 7191 32862 4 WL[36]
rlabel metal3 6064 30165 6064 30165 4 WL[33]
rlabel metal3 6064 29265 6064 29265 4 WL[32]
rlabel metal3 6064 35565 6064 35565 4 WL[39]
rlabel metal3 7191 31962 7191 31962 4 WL[35]
rlabel metal3 7191 31062 7191 31062 4 WL[34]
rlabel metal3 7191 30162 7191 30162 4 WL[33]
rlabel metal3 7264 35565 7264 35565 4 WL[39]
rlabel metal3 7264 29265 7264 29265 4 WL[32]
rlabel metal3 10734 31058 10734 31058 4 WL[34]
rlabel metal3 10734 35558 10734 35558 4 WL[39]
rlabel metal3 9664 31965 9664 31965 4 WL[35]
rlabel metal3 9664 32865 9664 32865 4 WL[36]
rlabel metal3 9664 33765 9664 33765 4 WL[37]
rlabel metal3 9591 31962 9591 31962 4 WL[35]
rlabel metal3 9591 31062 9591 31062 4 WL[34]
rlabel metal3 9591 30162 9591 30162 4 WL[33]
rlabel metal3 9591 29262 9591 29262 4 WL[32]
rlabel metal3 9591 35562 9591 35562 4 WL[39]
rlabel metal3 9591 34662 9591 34662 4 WL[38]
rlabel metal3 10791 33762 10791 33762 4 WL[37]
rlabel metal3 10791 32862 10791 32862 4 WL[36]
rlabel metal3 10734 33758 10734 33758 4 WL[37]
rlabel metal3 10791 31962 10791 31962 4 WL[35]
rlabel metal3 10791 31062 10791 31062 4 WL[34]
rlabel metal3 10791 30162 10791 30162 4 WL[33]
rlabel metal3 10791 29262 10791 29262 4 WL[32]
rlabel metal3 10791 35562 10791 35562 4 WL[39]
rlabel metal3 10791 34662 10791 34662 4 WL[38]
rlabel metal3 10191 33762 10191 33762 4 WL[37]
rlabel metal3 10191 32862 10191 32862 4 WL[36]
rlabel metal3 10734 34658 10734 34658 4 WL[38]
rlabel metal3 10191 31962 10191 31962 4 WL[35]
rlabel metal3 10191 31062 10191 31062 4 WL[34]
rlabel metal3 10734 32858 10734 32858 4 WL[36]
rlabel metal3 10191 30162 10191 30162 4 WL[33]
rlabel metal3 10191 29262 10191 29262 4 WL[32]
rlabel metal3 10734 30158 10734 30158 4 WL[33]
rlabel metal3 10734 31958 10734 31958 4 WL[35]
rlabel metal3 10191 35562 10191 35562 4 WL[39]
rlabel metal3 10191 34662 10191 34662 4 WL[38]
rlabel metal3 s 10134 29718 10134 29718 4 VSS
rlabel metal3 8991 33762 8991 33762 4 WL[37]
rlabel metal3 8991 32862 8991 32862 4 WL[36]
rlabel metal3 8991 31962 8991 31962 4 WL[35]
rlabel metal3 8991 31062 8991 31062 4 WL[34]
rlabel metal3 s 10134 28793 10134 28793 4 VDD
rlabel metal3 s 10734 29718 10734 29718 4 VSS
rlabel metal3 s 9534 29718 9534 29718 4 VSS
rlabel metal3 s 9534 28793 9534 28793 4 VDD
rlabel metal3 s 10734 28793 10734 28793 4 VDD
rlabel metal3 8991 30162 8991 30162 4 WL[33]
rlabel metal3 8991 29262 8991 29262 4 WL[32]
rlabel metal3 9664 35565 9664 35565 4 WL[39]
rlabel metal3 9664 29265 9664 29265 4 WL[32]
rlabel metal3 9591 33762 9591 33762 4 WL[37]
rlabel metal3 9591 32862 9591 32862 4 WL[36]
rlabel metal3 9664 30165 9664 30165 4 WL[33]
rlabel metal3 10734 29258 10734 29258 4 WL[32]
rlabel metal3 8991 35562 8991 35562 4 WL[39]
rlabel metal3 8991 34662 8991 34662 4 WL[38]
rlabel metal3 s 8934 29718 8934 29718 4 VSS
rlabel metal3 s 8934 28793 8934 28793 4 VDD
rlabel metal3 9664 34665 9664 34665 4 WL[38]
rlabel metal3 9664 31065 9664 31065 4 WL[34]
rlabel metal3 8479 23860 8479 23860 4 WL[26]
rlabel metal3 8479 24760 8479 24760 4 WL[27]
rlabel metal3 8479 25660 8479 25660 4 WL[28]
rlabel metal3 8479 26560 8479 26560 4 WL[29]
rlabel metal3 8479 27460 8479 27460 4 WL[30]
rlabel metal3 8479 28360 8479 28360 4 WL[31]
rlabel metal3 9679 23860 9679 23860 4 WL[26]
rlabel metal3 9679 24760 9679 24760 4 WL[27]
rlabel metal3 9679 25660 9679 25660 4 WL[28]
rlabel metal3 9679 26560 9679 26560 4 WL[29]
rlabel metal3 9679 27460 9679 27460 4 WL[30]
rlabel metal3 9679 28360 9679 28360 4 WL[31]
rlabel metal3 9679 22060 9679 22060 4 WL[24]
rlabel metal3 9679 22960 9679 22960 4 WL[25]
rlabel metal3 8479 22060 8479 22060 4 WL[24]
rlabel metal3 8479 22960 8479 22960 4 WL[25]
rlabel metal3 10719 22060 10719 22060 4 WL[24]
rlabel metal3 10777 22960 10777 22960 4 WL[25]
rlabel metal3 10777 22060 10777 22060 4 WL[24]
rlabel metal3 10777 28360 10777 28360 4 WL[31]
rlabel metal3 10777 27460 10777 27460 4 WL[30]
rlabel metal3 10777 26560 10777 26560 4 WL[29]
rlabel metal3 10777 25660 10777 25660 4 WL[28]
rlabel metal3 10777 24760 10777 24760 4 WL[27]
rlabel metal3 10777 23860 10777 23860 4 WL[26]
rlabel metal3 9577 22960 9577 22960 4 WL[25]
rlabel metal3 9577 22060 9577 22060 4 WL[24]
rlabel metal3 10177 22960 10177 22960 4 WL[25]
rlabel metal3 10177 22060 10177 22060 4 WL[24]
rlabel metal3 10177 28360 10177 28360 4 WL[31]
rlabel metal3 10177 27460 10177 27460 4 WL[30]
rlabel metal3 10177 26560 10177 26560 4 WL[29]
rlabel metal3 10177 25660 10177 25660 4 WL[28]
rlabel metal3 10177 24760 10177 24760 4 WL[27]
rlabel metal3 10177 23860 10177 23860 4 WL[26]
rlabel metal3 9577 28360 9577 28360 4 WL[31]
rlabel metal3 9577 27460 9577 27460 4 WL[30]
rlabel metal3 9577 26560 9577 26560 4 WL[29]
rlabel metal3 9577 25660 9577 25660 4 WL[28]
rlabel metal3 9577 24760 9577 24760 4 WL[27]
rlabel metal3 9577 23860 9577 23860 4 WL[26]
rlabel metal3 10719 22960 10719 22960 4 WL[25]
rlabel metal3 8977 22960 8977 22960 4 WL[25]
rlabel metal3 8977 22060 8977 22060 4 WL[24]
rlabel metal3 8977 28360 8977 28360 4 WL[31]
rlabel metal3 8977 27460 8977 27460 4 WL[30]
rlabel metal3 8977 26560 8977 26560 4 WL[29]
rlabel metal3 8977 25660 8977 25660 4 WL[28]
rlabel metal3 8977 24760 8977 24760 4 WL[27]
rlabel metal3 8977 23860 8977 23860 4 WL[26]
rlabel metal3 10719 23860 10719 23860 4 WL[26]
rlabel metal3 10719 24760 10719 24760 4 WL[27]
rlabel metal3 10719 25660 10719 25660 4 WL[28]
rlabel metal3 10719 26560 10719 26560 4 WL[29]
rlabel metal3 10719 27460 10719 27460 4 WL[30]
rlabel metal3 10719 28360 10719 28360 4 WL[31]
rlabel metal3 7177 24760 7177 24760 4 WL[27]
rlabel metal3 7177 22060 7177 22060 4 WL[24]
rlabel metal3 6577 28360 6577 28360 4 WL[31]
rlabel metal3 6577 27460 6577 27460 4 WL[30]
rlabel metal3 6577 26560 6577 26560 4 WL[29]
rlabel metal3 6079 22960 6079 22960 4 WL[25]
rlabel metal3 6079 22060 6079 22060 4 WL[24]
rlabel metal3 6577 22960 6577 22960 4 WL[25]
rlabel metal3 6577 22060 6577 22060 4 WL[24]
rlabel metal3 7177 23860 7177 23860 4 WL[26]
rlabel metal3 7777 22960 7777 22960 4 WL[25]
rlabel metal3 6577 25660 6577 25660 4 WL[28]
rlabel metal3 6577 24760 6577 24760 4 WL[27]
rlabel metal3 6577 23860 6577 23860 4 WL[26]
rlabel metal3 7177 22960 7177 22960 4 WL[25]
rlabel metal3 7777 22060 7777 22060 4 WL[24]
rlabel metal3 6079 28360 6079 28360 4 WL[31]
rlabel metal3 6079 27460 6079 27460 4 WL[30]
rlabel metal3 7777 28360 7777 28360 4 WL[31]
rlabel metal3 7777 27460 7777 27460 4 WL[30]
rlabel metal3 7777 26560 7777 26560 4 WL[29]
rlabel metal3 7777 25660 7777 25660 4 WL[28]
rlabel metal3 7777 24760 7777 24760 4 WL[27]
rlabel metal3 7777 23860 7777 23860 4 WL[26]
rlabel metal3 7279 23860 7279 23860 4 WL[26]
rlabel metal3 7279 24760 7279 24760 4 WL[27]
rlabel metal3 7279 25660 7279 25660 4 WL[28]
rlabel metal3 7279 26560 7279 26560 4 WL[29]
rlabel metal3 7279 27460 7279 27460 4 WL[30]
rlabel metal3 7279 28360 7279 28360 4 WL[31]
rlabel metal3 7279 22060 7279 22060 4 WL[24]
rlabel metal3 7279 22960 7279 22960 4 WL[25]
rlabel metal3 6079 25660 6079 25660 4 WL[28]
rlabel metal3 6079 23860 6079 23860 4 WL[26]
rlabel metal3 7177 28360 7177 28360 4 WL[31]
rlabel metal3 7177 27460 7177 27460 4 WL[30]
rlabel metal3 7177 26560 7177 26560 4 WL[29]
rlabel metal3 7177 25660 7177 25660 4 WL[28]
rlabel metal3 6079 26560 6079 26560 4 WL[29]
rlabel metal3 6079 24760 6079 24760 4 WL[27]
rlabel metal3 8377 22960 8377 22960 4 WL[25]
rlabel metal3 8377 22060 8377 22060 4 WL[24]
rlabel metal3 8377 28360 8377 28360 4 WL[31]
rlabel metal3 8377 27460 8377 27460 4 WL[30]
rlabel metal3 8377 26560 8377 26560 4 WL[29]
rlabel metal3 8377 25660 8377 25660 4 WL[28]
rlabel metal3 8377 24760 8377 24760 4 WL[27]
rlabel metal3 8377 23860 8377 23860 4 WL[26]
rlabel metal3 6079 18460 6079 18460 4 WL[20]
rlabel metal3 7777 18460 7777 18460 4 WL[20]
rlabel metal3 7177 19360 7177 19360 4 WL[21]
rlabel metal3 7777 17560 7777 17560 4 WL[19]
rlabel metal3 6577 21160 6577 21160 4 WL[23]
rlabel metal3 6577 20260 6577 20260 4 WL[22]
rlabel metal3 6577 19360 6577 19360 4 WL[21]
rlabel metal3 6577 18460 6577 18460 4 WL[20]
rlabel metal3 6577 17560 6577 17560 4 WL[19]
rlabel metal3 7177 20260 7177 20260 4 WL[22]
rlabel metal3 6577 16660 6577 16660 4 WL[18]
rlabel metal3 6577 15760 6577 15760 4 WL[17]
rlabel metal3 6577 14860 6577 14860 4 WL[16]
rlabel metal3 7279 14860 7279 14860 4 WL[16]
rlabel metal3 7279 15760 7279 15760 4 WL[17]
rlabel metal3 7279 16660 7279 16660 4 WL[18]
rlabel metal3 7279 17560 7279 17560 4 WL[19]
rlabel metal3 7279 18460 7279 18460 4 WL[20]
rlabel metal3 7279 19360 7279 19360 4 WL[21]
rlabel metal3 7279 20260 7279 20260 4 WL[22]
rlabel metal3 7279 21160 7279 21160 4 WL[23]
rlabel metal3 7777 16660 7777 16660 4 WL[18]
rlabel metal3 7777 15760 7777 15760 4 WL[17]
rlabel metal3 7777 14860 7777 14860 4 WL[16]
rlabel metal3 7777 21160 7777 21160 4 WL[23]
rlabel metal3 6079 14860 6079 14860 4 WL[16]
rlabel metal3 7777 20260 7777 20260 4 WL[22]
rlabel metal3 6079 21160 6079 21160 4 WL[23]
rlabel metal3 7177 21160 7177 21160 4 WL[23]
rlabel metal3 7777 19360 7777 19360 4 WL[21]
rlabel metal3 6079 17560 6079 17560 4 WL[19]
rlabel metal3 6079 16660 6079 16660 4 WL[18]
rlabel metal3 6079 15760 6079 15760 4 WL[17]
rlabel metal3 6079 20260 6079 20260 4 WL[22]
rlabel metal3 8377 21160 8377 21160 4 WL[23]
rlabel metal3 8377 20260 8377 20260 4 WL[22]
rlabel metal3 8377 19360 8377 19360 4 WL[21]
rlabel metal3 8377 18460 8377 18460 4 WL[20]
rlabel metal3 8377 17560 8377 17560 4 WL[19]
rlabel metal3 8377 16660 8377 16660 4 WL[18]
rlabel metal3 8377 15760 8377 15760 4 WL[17]
rlabel metal3 8377 14860 8377 14860 4 WL[16]
rlabel metal3 7177 18460 7177 18460 4 WL[20]
rlabel metal3 7177 17560 7177 17560 4 WL[19]
rlabel metal3 7177 15760 7177 15760 4 WL[17]
rlabel metal3 7177 16660 7177 16660 4 WL[18]
rlabel metal3 7177 14860 7177 14860 4 WL[16]
rlabel metal3 6079 19360 6079 19360 4 WL[21]
rlabel metal3 8977 19360 8977 19360 4 WL[21]
rlabel metal3 8977 18460 8977 18460 4 WL[20]
rlabel metal3 8977 17560 8977 17560 4 WL[19]
rlabel metal3 8977 16660 8977 16660 4 WL[18]
rlabel metal3 8977 15760 8977 15760 4 WL[17]
rlabel metal3 8977 14860 8977 14860 4 WL[16]
rlabel metal3 9577 15760 9577 15760 4 WL[17]
rlabel metal3 9577 14860 9577 14860 4 WL[16]
rlabel metal3 8479 21160 8479 21160 4 WL[23]
rlabel metal3 9679 16660 9679 16660 4 WL[18]
rlabel metal3 10177 21160 10177 21160 4 WL[23]
rlabel metal3 10177 20260 10177 20260 4 WL[22]
rlabel metal3 10177 19360 10177 19360 4 WL[21]
rlabel metal3 10177 18460 10177 18460 4 WL[20]
rlabel metal3 10177 17560 10177 17560 4 WL[19]
rlabel metal3 10177 16660 10177 16660 4 WL[18]
rlabel metal3 10177 15760 10177 15760 4 WL[17]
rlabel metal3 10177 14860 10177 14860 4 WL[16]
rlabel metal3 9679 17560 9679 17560 4 WL[19]
rlabel metal3 9679 18460 9679 18460 4 WL[20]
rlabel metal3 10719 17560 10719 17560 4 WL[19]
rlabel metal3 10719 16660 10719 16660 4 WL[18]
rlabel metal3 9679 19360 9679 19360 4 WL[21]
rlabel metal3 10777 21160 10777 21160 4 WL[23]
rlabel metal3 10777 20260 10777 20260 4 WL[22]
rlabel metal3 10777 19360 10777 19360 4 WL[21]
rlabel metal3 10777 18460 10777 18460 4 WL[20]
rlabel metal3 10777 17560 10777 17560 4 WL[19]
rlabel metal3 10719 20260 10719 20260 4 WL[22]
rlabel metal3 10719 14860 10719 14860 4 WL[16]
rlabel metal3 10777 16660 10777 16660 4 WL[18]
rlabel metal3 10777 15760 10777 15760 4 WL[17]
rlabel metal3 10719 19360 10719 19360 4 WL[21]
rlabel metal3 10777 14860 10777 14860 4 WL[16]
rlabel metal3 9679 20260 9679 20260 4 WL[22]
rlabel metal3 9679 21160 9679 21160 4 WL[23]
rlabel metal3 9679 14860 9679 14860 4 WL[16]
rlabel metal3 9679 15760 9679 15760 4 WL[17]
rlabel metal3 8479 14860 8479 14860 4 WL[16]
rlabel metal3 8479 15760 8479 15760 4 WL[17]
rlabel metal3 8479 16660 8479 16660 4 WL[18]
rlabel metal3 8479 17560 8479 17560 4 WL[19]
rlabel metal3 8479 18460 8479 18460 4 WL[20]
rlabel metal3 10719 18460 10719 18460 4 WL[20]
rlabel metal3 8479 19360 8479 19360 4 WL[21]
rlabel metal3 8479 20260 8479 20260 4 WL[22]
rlabel metal3 9577 21160 9577 21160 4 WL[23]
rlabel metal3 9577 20260 9577 20260 4 WL[22]
rlabel metal3 9577 19360 9577 19360 4 WL[21]
rlabel metal3 9577 18460 9577 18460 4 WL[20]
rlabel metal3 10719 21160 10719 21160 4 WL[23]
rlabel metal3 10719 15760 10719 15760 4 WL[17]
rlabel metal3 9577 17560 9577 17560 4 WL[19]
rlabel metal3 9577 16660 9577 16660 4 WL[18]
rlabel metal3 8977 21160 8977 21160 4 WL[23]
rlabel metal3 8977 20260 8977 20260 4 WL[22]
rlabel metal3 4121 23860 4121 23860 4 WL[26]
rlabel metal3 4121 24760 4121 24760 4 WL[27]
rlabel metal3 4121 25660 4121 25660 4 WL[28]
rlabel metal3 4121 26560 4121 26560 4 WL[29]
rlabel metal3 4121 27460 4121 27460 4 WL[30]
rlabel metal3 4121 28360 4121 28360 4 WL[31]
rlabel metal3 4121 22060 4121 22060 4 WL[24]
rlabel metal3 4121 22960 4121 22960 4 WL[25]
rlabel metal3 5321 22060 5321 22060 4 WL[24]
rlabel metal3 5321 22960 5321 22960 4 WL[25]
rlabel metal3 4223 22960 4223 22960 4 WL[25]
rlabel metal3 4223 22060 4223 22060 4 WL[24]
rlabel metal3 3623 22960 3623 22960 4 WL[25]
rlabel metal3 3623 22060 3623 22060 4 WL[24]
rlabel metal3 3623 28360 3623 28360 4 WL[31]
rlabel metal3 3623 27460 3623 27460 4 WL[30]
rlabel metal3 3623 26560 3623 26560 4 WL[29]
rlabel metal3 3623 25660 3623 25660 4 WL[28]
rlabel metal3 3623 24760 3623 24760 4 WL[27]
rlabel metal3 3623 23860 3623 23860 4 WL[26]
rlabel metal3 4223 28360 4223 28360 4 WL[31]
rlabel metal3 4223 27460 4223 27460 4 WL[30]
rlabel metal3 4223 26560 4223 26560 4 WL[29]
rlabel metal3 4223 25660 4223 25660 4 WL[28]
rlabel metal3 4223 24760 4223 24760 4 WL[27]
rlabel metal3 4223 23860 4223 23860 4 WL[26]
rlabel metal3 5321 23860 5321 23860 4 WL[26]
rlabel metal3 5321 24760 5321 24760 4 WL[27]
rlabel metal3 5321 25660 5321 25660 4 WL[28]
rlabel metal3 5321 26560 5321 26560 4 WL[29]
rlabel metal3 5321 27460 5321 27460 4 WL[30]
rlabel metal3 5321 28360 5321 28360 4 WL[31]
rlabel metal3 4823 22960 4823 22960 4 WL[25]
rlabel metal3 4823 22060 4823 22060 4 WL[24]
rlabel metal3 4823 28360 4823 28360 4 WL[31]
rlabel metal3 4823 27460 4823 27460 4 WL[30]
rlabel metal3 4823 26560 4823 26560 4 WL[29]
rlabel metal3 4823 25660 4823 25660 4 WL[28]
rlabel metal3 4823 24760 4823 24760 4 WL[27]
rlabel metal3 4823 23860 4823 23860 4 WL[26]
rlabel metal3 1721 26560 1721 26560 4 WL[29]
rlabel metal3 1721 27460 1721 27460 4 WL[30]
rlabel metal3 1721 28360 1721 28360 4 WL[31]
rlabel metal3 1721 22060 1721 22060 4 WL[24]
rlabel metal3 1721 22960 1721 22960 4 WL[25]
rlabel metal3 1823 27460 1823 27460 4 WL[30]
rlabel metal3 1823 26560 1823 26560 4 WL[29]
rlabel metal3 1823 25660 1823 25660 4 WL[28]
rlabel metal3 2423 22060 2423 22060 4 WL[24]
rlabel metal3 2921 23860 2921 23860 4 WL[26]
rlabel metal3 2921 24760 2921 24760 4 WL[27]
rlabel metal3 2921 25660 2921 25660 4 WL[28]
rlabel metal3 2921 26560 2921 26560 4 WL[29]
rlabel metal3 2921 27460 2921 27460 4 WL[30]
rlabel metal3 2921 28360 2921 28360 4 WL[31]
rlabel metal3 3023 28360 3023 28360 4 WL[31]
rlabel metal3 3023 27460 3023 27460 4 WL[30]
rlabel metal3 3023 26560 3023 26560 4 WL[29]
rlabel metal3 3023 25660 3023 25660 4 WL[28]
rlabel metal3 3023 24760 3023 24760 4 WL[27]
rlabel metal3 1823 24760 1823 24760 4 WL[27]
rlabel metal3 1823 23860 1823 23860 4 WL[26]
rlabel metal3 2423 28360 2423 28360 4 WL[31]
rlabel metal3 2423 27460 2423 27460 4 WL[30]
rlabel metal3 2423 26560 2423 26560 4 WL[29]
rlabel metal3 2423 25660 2423 25660 4 WL[28]
rlabel metal3 2423 24760 2423 24760 4 WL[27]
rlabel metal3 2423 23860 2423 23860 4 WL[26]
rlabel metal3 3023 23860 3023 23860 4 WL[26]
rlabel metal3 1223 23860 1223 23860 4 WL[26]
rlabel metal3 681 24760 681 24760 4 WL[27]
rlabel metal3 1223 24760 1223 24760 4 WL[27]
rlabel metal3 681 23860 681 23860 4 WL[26]
rlabel metal3 681 22960 681 22960 4 WL[25]
rlabel metal3 681 22060 681 22060 4 WL[24]
rlabel metal3 3023 22960 3023 22960 4 WL[25]
rlabel metal3 623 22960 623 22960 4 WL[25]
rlabel metal3 623 22060 623 22060 4 WL[24]
rlabel metal3 2921 22060 2921 22060 4 WL[24]
rlabel metal3 2921 22960 2921 22960 4 WL[25]
rlabel metal3 623 28360 623 28360 4 WL[31]
rlabel metal3 623 27460 623 27460 4 WL[30]
rlabel metal3 623 26560 623 26560 4 WL[29]
rlabel metal3 623 25660 623 25660 4 WL[28]
rlabel metal3 623 24760 623 24760 4 WL[27]
rlabel metal3 623 23860 623 23860 4 WL[26]
rlabel metal3 3023 22060 3023 22060 4 WL[24]
rlabel metal3 1823 28360 1823 28360 4 WL[31]
rlabel metal3 2423 22960 2423 22960 4 WL[25]
rlabel metal3 1721 23860 1721 23860 4 WL[26]
rlabel metal3 1721 24760 1721 24760 4 WL[27]
rlabel metal3 1721 25660 1721 25660 4 WL[28]
rlabel metal3 1223 22960 1223 22960 4 WL[25]
rlabel metal3 1223 22060 1223 22060 4 WL[24]
rlabel metal3 681 28360 681 28360 4 WL[31]
rlabel metal3 681 27460 681 27460 4 WL[30]
rlabel metal3 681 26560 681 26560 4 WL[29]
rlabel metal3 1223 28360 1223 28360 4 WL[31]
rlabel metal3 1223 27460 1223 27460 4 WL[30]
rlabel metal3 1223 26560 1223 26560 4 WL[29]
rlabel metal3 1223 25660 1223 25660 4 WL[28]
rlabel metal3 681 25660 681 25660 4 WL[28]
rlabel metal3 1823 22960 1823 22960 4 WL[25]
rlabel metal3 1823 22060 1823 22060 4 WL[24]
rlabel metal3 1721 19360 1721 19360 4 WL[21]
rlabel metal3 1721 20260 1721 20260 4 WL[22]
rlabel metal3 1721 21160 1721 21160 4 WL[23]
rlabel metal3 681 20260 681 20260 4 WL[22]
rlabel metal3 3023 21160 3023 21160 4 WL[23]
rlabel metal3 2423 19360 2423 19360 4 WL[21]
rlabel metal3 623 21160 623 21160 4 WL[23]
rlabel metal3 2921 14860 2921 14860 4 WL[16]
rlabel metal3 2921 15760 2921 15760 4 WL[17]
rlabel metal3 2921 16660 2921 16660 4 WL[18]
rlabel metal3 2921 17560 2921 17560 4 WL[19]
rlabel metal3 2921 18460 2921 18460 4 WL[20]
rlabel metal3 2921 19360 2921 19360 4 WL[21]
rlabel metal3 623 20260 623 20260 4 WL[22]
rlabel metal3 623 19360 623 19360 4 WL[21]
rlabel metal3 623 18460 623 18460 4 WL[20]
rlabel metal3 623 17560 623 17560 4 WL[19]
rlabel metal3 623 16660 623 16660 4 WL[18]
rlabel metal3 623 15760 623 15760 4 WL[17]
rlabel metal3 623 14860 623 14860 4 WL[16]
rlabel metal3 2921 20260 2921 20260 4 WL[22]
rlabel metal3 2921 21160 2921 21160 4 WL[23]
rlabel metal3 2423 18460 2423 18460 4 WL[20]
rlabel metal3 2423 17560 2423 17560 4 WL[19]
rlabel metal3 2423 16660 2423 16660 4 WL[18]
rlabel metal3 2423 15760 2423 15760 4 WL[17]
rlabel metal3 2423 14860 2423 14860 4 WL[16]
rlabel metal3 3023 20260 3023 20260 4 WL[22]
rlabel metal3 3023 19360 3023 19360 4 WL[21]
rlabel metal3 3023 18460 3023 18460 4 WL[20]
rlabel metal3 3023 17560 3023 17560 4 WL[19]
rlabel metal3 3023 16660 3023 16660 4 WL[18]
rlabel metal3 3023 15760 3023 15760 4 WL[17]
rlabel metal3 3023 14860 3023 14860 4 WL[16]
rlabel metal3 681 19360 681 19360 4 WL[21]
rlabel metal3 681 18460 681 18460 4 WL[20]
rlabel metal3 681 17560 681 17560 4 WL[19]
rlabel metal3 2423 21160 2423 21160 4 WL[23]
rlabel metal3 1223 21160 1223 21160 4 WL[23]
rlabel metal3 1223 20260 1223 20260 4 WL[22]
rlabel metal3 1223 19360 1223 19360 4 WL[21]
rlabel metal3 1223 18460 1223 18460 4 WL[20]
rlabel metal3 1223 17560 1223 17560 4 WL[19]
rlabel metal3 1223 16660 1223 16660 4 WL[18]
rlabel metal3 2423 20260 2423 20260 4 WL[22]
rlabel metal3 681 16660 681 16660 4 WL[18]
rlabel metal3 681 15760 681 15760 4 WL[17]
rlabel metal3 1223 15760 1223 15760 4 WL[17]
rlabel metal3 1223 14860 1223 14860 4 WL[16]
rlabel metal3 681 14860 681 14860 4 WL[16]
rlabel metal3 681 21160 681 21160 4 WL[23]
rlabel metal3 1721 14860 1721 14860 4 WL[16]
rlabel metal3 1721 15760 1721 15760 4 WL[17]
rlabel metal3 1721 16660 1721 16660 4 WL[18]
rlabel metal3 1721 17560 1721 17560 4 WL[19]
rlabel metal3 1721 18460 1721 18460 4 WL[20]
rlabel metal3 1823 21160 1823 21160 4 WL[23]
rlabel metal3 1823 20260 1823 20260 4 WL[22]
rlabel metal3 1823 19360 1823 19360 4 WL[21]
rlabel metal3 1823 18460 1823 18460 4 WL[20]
rlabel metal3 1823 17560 1823 17560 4 WL[19]
rlabel metal3 1823 16660 1823 16660 4 WL[18]
rlabel metal3 1823 15760 1823 15760 4 WL[17]
rlabel metal3 1823 14860 1823 14860 4 WL[16]
rlabel metal3 4121 21160 4121 21160 4 WL[23]
rlabel metal3 4121 14860 4121 14860 4 WL[16]
rlabel metal3 4121 15760 4121 15760 4 WL[17]
rlabel metal3 5321 14860 5321 14860 4 WL[16]
rlabel metal3 5321 15760 5321 15760 4 WL[17]
rlabel metal3 4223 21160 4223 21160 4 WL[23]
rlabel metal3 4223 20260 4223 20260 4 WL[22]
rlabel metal3 4223 19360 4223 19360 4 WL[21]
rlabel metal3 4223 18460 4223 18460 4 WL[20]
rlabel metal3 4223 17560 4223 17560 4 WL[19]
rlabel metal3 4223 16660 4223 16660 4 WL[18]
rlabel metal3 4223 15760 4223 15760 4 WL[17]
rlabel metal3 4823 21160 4823 21160 4 WL[23]
rlabel metal3 4823 20260 4823 20260 4 WL[22]
rlabel metal3 4823 19360 4823 19360 4 WL[21]
rlabel metal3 5321 16660 5321 16660 4 WL[18]
rlabel metal3 5321 17560 5321 17560 4 WL[19]
rlabel metal3 3623 21160 3623 21160 4 WL[23]
rlabel metal3 3623 20260 3623 20260 4 WL[22]
rlabel metal3 3623 19360 3623 19360 4 WL[21]
rlabel metal3 3623 18460 3623 18460 4 WL[20]
rlabel metal3 3623 17560 3623 17560 4 WL[19]
rlabel metal3 3623 16660 3623 16660 4 WL[18]
rlabel metal3 3623 15760 3623 15760 4 WL[17]
rlabel metal3 3623 14860 3623 14860 4 WL[16]
rlabel metal3 4223 14860 4223 14860 4 WL[16]
rlabel metal3 5321 18460 5321 18460 4 WL[20]
rlabel metal3 5321 19360 5321 19360 4 WL[21]
rlabel metal3 5321 20260 5321 20260 4 WL[22]
rlabel metal3 5321 21160 5321 21160 4 WL[23]
rlabel metal3 4121 16660 4121 16660 4 WL[18]
rlabel metal3 4823 18460 4823 18460 4 WL[20]
rlabel metal3 4823 17560 4823 17560 4 WL[19]
rlabel metal3 4823 16660 4823 16660 4 WL[18]
rlabel metal3 4121 17560 4121 17560 4 WL[19]
rlabel metal3 4121 18460 4121 18460 4 WL[20]
rlabel metal3 4121 19360 4121 19360 4 WL[21]
rlabel metal3 4121 20260 4121 20260 4 WL[22]
rlabel metal3 4823 15760 4823 15760 4 WL[17]
rlabel metal3 4823 14860 4823 14860 4 WL[16]
rlabel metal3 3623 13960 3623 13960 4 WL[15]
rlabel metal3 3623 13060 3623 13060 4 WL[14]
rlabel metal3 3623 12160 3623 12160 4 WL[13]
rlabel metal3 3623 11260 3623 11260 4 WL[12]
rlabel metal3 3623 10360 3623 10360 4 WL[11]
rlabel metal3 3623 9460 3623 9460 4 WL[10]
rlabel metal3 3623 8560 3623 8560 4 WL[9]
rlabel metal3 3623 7660 3623 7660 4 WL[8]
rlabel metal3 4223 13960 4223 13960 4 WL[15]
rlabel metal3 4223 13060 4223 13060 4 WL[14]
rlabel metal3 4223 12160 4223 12160 4 WL[13]
rlabel metal3 4223 11260 4223 11260 4 WL[12]
rlabel metal3 4223 10360 4223 10360 4 WL[11]
rlabel metal3 4223 9460 4223 9460 4 WL[10]
rlabel metal3 4223 8560 4223 8560 4 WL[9]
rlabel metal3 4223 7660 4223 7660 4 WL[8]
rlabel metal3 4121 7660 4121 7660 4 WL[8]
rlabel metal3 4121 8560 4121 8560 4 WL[9]
rlabel metal3 4121 9460 4121 9460 4 WL[10]
rlabel metal3 4121 10360 4121 10360 4 WL[11]
rlabel metal3 4121 11260 4121 11260 4 WL[12]
rlabel metal3 4121 12160 4121 12160 4 WL[13]
rlabel metal3 4121 13060 4121 13060 4 WL[14]
rlabel metal3 4121 13960 4121 13960 4 WL[15]
rlabel metal3 5321 7660 5321 7660 4 WL[8]
rlabel metal3 5321 8560 5321 8560 4 WL[9]
rlabel metal3 5321 9460 5321 9460 4 WL[10]
rlabel metal3 5321 10360 5321 10360 4 WL[11]
rlabel metal3 4823 13960 4823 13960 4 WL[15]
rlabel metal3 4823 13060 4823 13060 4 WL[14]
rlabel metal3 4823 12160 4823 12160 4 WL[13]
rlabel metal3 4823 11260 4823 11260 4 WL[12]
rlabel metal3 4823 10360 4823 10360 4 WL[11]
rlabel metal3 4823 9460 4823 9460 4 WL[10]
rlabel metal3 4823 8560 4823 8560 4 WL[9]
rlabel metal3 4823 7660 4823 7660 4 WL[8]
rlabel metal3 5321 11260 5321 11260 4 WL[12]
rlabel metal3 5321 12160 5321 12160 4 WL[13]
rlabel metal3 5321 13060 5321 13060 4 WL[14]
rlabel metal3 5321 13960 5321 13960 4 WL[15]
rlabel metal3 3023 11260 3023 11260 4 WL[12]
rlabel metal3 3023 10360 3023 10360 4 WL[11]
rlabel metal3 3023 9460 3023 9460 4 WL[10]
rlabel metal3 3023 8560 3023 8560 4 WL[9]
rlabel metal3 3023 7660 3023 7660 4 WL[8]
rlabel metal3 1823 12160 1823 12160 4 WL[13]
rlabel metal3 1823 11260 1823 11260 4 WL[12]
rlabel metal3 1823 10360 1823 10360 4 WL[11]
rlabel metal3 1823 9460 1823 9460 4 WL[10]
rlabel metal3 681 11260 681 11260 4 WL[12]
rlabel metal3 623 13960 623 13960 4 WL[15]
rlabel metal3 623 13060 623 13060 4 WL[14]
rlabel metal3 623 12160 623 12160 4 WL[13]
rlabel metal3 2921 7660 2921 7660 4 WL[8]
rlabel metal3 2921 8560 2921 8560 4 WL[9]
rlabel metal3 2921 9460 2921 9460 4 WL[10]
rlabel metal3 623 11260 623 11260 4 WL[12]
rlabel metal3 623 10360 623 10360 4 WL[11]
rlabel metal3 623 9460 623 9460 4 WL[10]
rlabel metal3 623 8560 623 8560 4 WL[9]
rlabel metal3 623 7660 623 7660 4 WL[8]
rlabel metal3 2921 10360 2921 10360 4 WL[11]
rlabel metal3 2921 11260 2921 11260 4 WL[12]
rlabel metal3 2921 12160 2921 12160 4 WL[13]
rlabel metal3 2921 13060 2921 13060 4 WL[14]
rlabel metal3 2921 13960 2921 13960 4 WL[15]
rlabel metal3 1721 12160 1721 12160 4 WL[13]
rlabel metal3 1721 13060 1721 13060 4 WL[14]
rlabel metal3 1721 13960 1721 13960 4 WL[15]
rlabel metal3 681 13960 681 13960 4 WL[15]
rlabel metal3 681 13060 681 13060 4 WL[14]
rlabel metal3 2423 13960 2423 13960 4 WL[15]
rlabel metal3 2423 13060 2423 13060 4 WL[14]
rlabel metal3 2423 12160 2423 12160 4 WL[13]
rlabel metal3 2423 11260 2423 11260 4 WL[12]
rlabel metal3 2423 10360 2423 10360 4 WL[11]
rlabel metal3 2423 9460 2423 9460 4 WL[10]
rlabel metal3 681 10360 681 10360 4 WL[11]
rlabel metal3 681 12160 681 12160 4 WL[13]
rlabel metal3 681 8560 681 8560 4 WL[9]
rlabel metal3 1721 7660 1721 7660 4 WL[8]
rlabel metal3 1721 8560 1721 8560 4 WL[9]
rlabel metal3 1721 9460 1721 9460 4 WL[10]
rlabel metal3 1721 10360 1721 10360 4 WL[11]
rlabel metal3 681 7660 681 7660 4 WL[8]
rlabel metal3 2423 8560 2423 8560 4 WL[9]
rlabel metal3 2423 7660 2423 7660 4 WL[8]
rlabel metal3 1721 11260 1721 11260 4 WL[12]
rlabel metal3 3023 13960 3023 13960 4 WL[15]
rlabel metal3 3023 13060 3023 13060 4 WL[14]
rlabel metal3 3023 12160 3023 12160 4 WL[13]
rlabel metal3 681 9460 681 9460 4 WL[10]
rlabel metal3 1823 8560 1823 8560 4 WL[9]
rlabel metal3 1823 7660 1823 7660 4 WL[8]
rlabel metal3 1223 13960 1223 13960 4 WL[15]
rlabel metal3 1223 13060 1223 13060 4 WL[14]
rlabel metal3 1223 12160 1223 12160 4 WL[13]
rlabel metal3 1223 11260 1223 11260 4 WL[12]
rlabel metal3 1223 10360 1223 10360 4 WL[11]
rlabel metal3 1223 9460 1223 9460 4 WL[10]
rlabel metal3 1223 8560 1223 8560 4 WL[9]
rlabel metal3 1223 7660 1223 7660 4 WL[8]
rlabel metal3 1823 13960 1823 13960 4 WL[15]
rlabel metal3 1823 13060 1823 13060 4 WL[14]
rlabel metal3 s 1866 -7 1866 -7 4 VDD
rlabel metal3 2921 4960 2921 4960 4 WL[5]
rlabel metal3 2921 5860 2921 5860 4 WL[6]
rlabel metal3 2921 6760 2921 6760 4 WL[7]
rlabel metal3 1223 1360 1223 1360 4 WL[1]
rlabel metal3 s 2466 918 2466 918 4 VSS
rlabel metal3 2423 2260 2423 2260 4 WL[2]
rlabel metal3 2423 1360 2423 1360 4 WL[1]
rlabel metal3 2423 460 2423 460 4 WL[0]
rlabel metal3 1721 460 1721 460 4 WL[0]
rlabel metal3 1721 1360 1721 1360 4 WL[1]
rlabel metal3 1721 2260 1721 2260 4 WL[2]
rlabel metal3 623 6760 623 6760 4 WL[7]
rlabel metal3 1721 3160 1721 3160 4 WL[3]
rlabel metal3 1823 3160 1823 3160 4 WL[3]
rlabel metal3 1721 4060 1721 4060 4 WL[4]
rlabel metal3 1721 4960 1721 4960 4 WL[5]
rlabel metal3 1721 5860 1721 5860 4 WL[6]
rlabel metal3 623 5860 623 5860 4 WL[6]
rlabel metal3 623 4960 623 4960 4 WL[5]
rlabel metal3 623 4060 623 4060 4 WL[4]
rlabel metal3 623 3160 623 3160 4 WL[3]
rlabel metal3 623 2260 623 2260 4 WL[2]
rlabel metal3 623 1360 623 1360 4 WL[1]
rlabel metal3 623 460 623 460 4 WL[0]
rlabel metal3 1721 6760 1721 6760 4 WL[7]
rlabel metal3 s 1266 -11 1266 -11 4 VDD
rlabel metal3 681 4960 681 4960 4 WL[5]
rlabel metal3 s 1266 918 1266 918 4 VSS
rlabel metal3 s 1266 -7 1266 -7 4 VDD
rlabel metal3 3023 6760 3023 6760 4 WL[7]
rlabel metal3 3023 5860 3023 5860 4 WL[6]
rlabel metal3 3023 4960 3023 4960 4 WL[5]
rlabel metal3 s 1734 907 1734 907 4 VSS
rlabel metal3 s 1734 5 1734 5 4 VDD
rlabel metal3 3023 4060 3023 4060 4 WL[4]
rlabel metal3 s 666 918 666 918 4 VSS
rlabel metal3 s 2466 -11 2466 -11 4 VDD
rlabel metal3 s 666 -11 666 -11 4 VDD
rlabel metal3 s 666 918 666 918 4 VSS
rlabel metal3 s 666 -7 666 -7 4 VDD
rlabel metal3 s 2466 918 2466 918 4 VSS
rlabel metal3 s 2466 -7 2466 -7 4 VDD
rlabel metal3 s 1266 918 1266 918 4 VSS
rlabel metal3 3023 3160 3023 3160 4 WL[3]
rlabel metal3 3023 2260 3023 2260 4 WL[2]
rlabel metal3 3023 1360 3023 1360 4 WL[1]
rlabel metal3 s 2934 907 2934 907 4 VSS
rlabel metal3 s 2934 5 2934 5 4 VDD
rlabel metal3 s 1866 918 1866 918 4 VSS
rlabel metal3 3023 460 3023 460 4 WL[0]
rlabel metal3 681 6760 681 6760 4 WL[7]
rlabel metal3 681 5860 681 5860 4 WL[6]
rlabel metal3 681 2260 681 2260 4 WL[2]
rlabel metal3 1823 2260 1823 2260 4 WL[2]
rlabel metal3 s 666 920 666 920 4 VSS
rlabel metal3 2423 6760 2423 6760 4 WL[7]
rlabel metal3 2423 5860 2423 5860 4 WL[6]
rlabel metal3 2423 4960 2423 4960 4 WL[5]
rlabel metal3 2423 4060 2423 4060 4 WL[4]
rlabel metal3 2423 3160 2423 3160 4 WL[3]
rlabel metal3 1823 1360 1823 1360 4 WL[1]
rlabel metal3 1823 460 1823 460 4 WL[0]
rlabel metal3 s 3066 918 3066 918 4 VSS
rlabel metal3 681 1360 681 1360 4 WL[1]
rlabel metal3 681 460 681 460 4 WL[0]
rlabel metal3 1223 460 1223 460 4 WL[0]
rlabel metal3 s 1866 -11 1866 -11 4 VDD
rlabel metal3 s 1866 918 1866 918 4 VSS
rlabel metal3 1823 5860 1823 5860 4 WL[6]
rlabel metal3 681 4060 681 4060 4 WL[4]
rlabel metal3 681 3160 681 3160 4 WL[3]
rlabel metal3 1823 6760 1823 6760 4 WL[7]
rlabel metal3 2921 460 2921 460 4 WL[0]
rlabel metal3 2921 1360 2921 1360 4 WL[1]
rlabel metal3 2921 2260 2921 2260 4 WL[2]
rlabel metal3 2921 3160 2921 3160 4 WL[3]
rlabel metal3 2921 4060 2921 4060 4 WL[4]
rlabel metal3 s 3066 -11 3066 -11 4 VDD
rlabel metal3 s 3066 918 3066 918 4 VSS
rlabel metal3 s 3066 -7 3066 -7 4 VDD
rlabel metal3 1223 6760 1223 6760 4 WL[7]
rlabel metal3 1223 5860 1223 5860 4 WL[6]
rlabel metal3 1223 4960 1223 4960 4 WL[5]
rlabel metal3 1223 4060 1223 4060 4 WL[4]
rlabel metal3 1223 3160 1223 3160 4 WL[3]
rlabel metal3 1223 2260 1223 2260 4 WL[2]
rlabel metal3 1823 4960 1823 4960 4 WL[5]
rlabel metal3 1823 4060 1823 4060 4 WL[4]
rlabel metal3 5321 6760 5321 6760 4 WL[7]
rlabel metal3 4223 4960 4223 4960 4 WL[5]
rlabel metal3 4223 4060 4223 4060 4 WL[4]
rlabel metal3 4223 3160 4223 3160 4 WL[3]
rlabel metal3 4223 2260 4223 2260 4 WL[2]
rlabel metal3 4223 1360 4223 1360 4 WL[1]
rlabel metal3 4823 6760 4823 6760 4 WL[7]
rlabel metal3 4823 5860 4823 5860 4 WL[6]
rlabel metal3 4223 460 4223 460 4 WL[0]
rlabel metal3 3623 460 3623 460 4 WL[0]
rlabel metal3 5321 460 5321 460 4 WL[0]
rlabel metal3 4823 4960 4823 4960 4 WL[5]
rlabel metal3 4823 4060 4823 4060 4 WL[4]
rlabel metal3 4823 3160 4823 3160 4 WL[3]
rlabel metal3 4823 2260 4823 2260 4 WL[2]
rlabel metal3 4823 1360 4823 1360 4 WL[1]
rlabel metal3 4823 460 4823 460 4 WL[0]
rlabel metal3 s 4266 -11 4266 -11 4 VDD
rlabel metal3 s 4266 918 4266 918 4 VSS
rlabel metal3 s 4266 -7 4266 -7 4 VDD
rlabel metal3 s 4134 907 4134 907 4 VSS
rlabel metal3 s 4866 918 4866 918 4 VSS
rlabel metal3 s 4134 5 4134 5 4 VDD
rlabel metal3 s 4866 -7 4866 -7 4 VDD
rlabel metal3 s 4866 -11 4866 -11 4 VDD
rlabel metal3 s 4866 918 4866 918 4 VSS
rlabel metal3 3623 6760 3623 6760 4 WL[7]
rlabel metal3 3623 5860 3623 5860 4 WL[6]
rlabel metal3 3623 4960 3623 4960 4 WL[5]
rlabel metal3 5321 1360 5321 1360 4 WL[1]
rlabel metal3 5321 2260 5321 2260 4 WL[2]
rlabel metal3 5321 3160 5321 3160 4 WL[3]
rlabel metal3 3623 4060 3623 4060 4 WL[4]
rlabel metal3 3623 3160 3623 3160 4 WL[3]
rlabel metal3 s 3666 -11 3666 -11 4 VDD
rlabel metal3 4121 5860 4121 5860 4 WL[6]
rlabel metal3 s 3666 918 3666 918 4 VSS
rlabel metal3 s 4266 918 4266 918 4 VSS
rlabel metal3 3623 2260 3623 2260 4 WL[2]
rlabel metal3 s 5334 907 5334 907 4 VSS
rlabel metal3 s 5334 5 5334 5 4 VDD
rlabel metal3 s 3666 918 3666 918 4 VSS
rlabel metal3 4121 6760 4121 6760 4 WL[7]
rlabel metal3 s 3666 -7 3666 -7 4 VDD
rlabel metal3 3623 1360 3623 1360 4 WL[1]
rlabel metal3 4223 6760 4223 6760 4 WL[7]
rlabel metal3 4223 5860 4223 5860 4 WL[6]
rlabel metal3 4121 460 4121 460 4 WL[0]
rlabel metal3 4121 1360 4121 1360 4 WL[1]
rlabel metal3 4121 2260 4121 2260 4 WL[2]
rlabel metal3 4121 3160 4121 3160 4 WL[3]
rlabel metal3 4121 4060 4121 4060 4 WL[4]
rlabel metal3 4121 4960 4121 4960 4 WL[5]
rlabel metal3 5321 4060 5321 4060 4 WL[4]
rlabel metal3 5321 4960 5321 4960 4 WL[5]
rlabel metal3 5321 5860 5321 5860 4 WL[6]
rlabel metal3 10719 7660 10719 7660 4 WL[8]
rlabel metal3 8479 7660 8479 7660 4 WL[8]
rlabel metal3 8479 8560 8479 8560 4 WL[9]
rlabel metal3 8977 13960 8977 13960 4 WL[15]
rlabel metal3 8977 13060 8977 13060 4 WL[14]
rlabel metal3 8977 12160 8977 12160 4 WL[13]
rlabel metal3 8977 11260 8977 11260 4 WL[12]
rlabel metal3 8977 10360 8977 10360 4 WL[11]
rlabel metal3 8977 9460 8977 9460 4 WL[10]
rlabel metal3 8977 8560 8977 8560 4 WL[9]
rlabel metal3 8977 7660 8977 7660 4 WL[8]
rlabel metal3 10719 8560 10719 8560 4 WL[9]
rlabel metal3 8479 9460 8479 9460 4 WL[10]
rlabel metal3 8479 10360 8479 10360 4 WL[11]
rlabel metal3 10777 13960 10777 13960 4 WL[15]
rlabel metal3 10777 13060 10777 13060 4 WL[14]
rlabel metal3 10777 12160 10777 12160 4 WL[13]
rlabel metal3 10777 11260 10777 11260 4 WL[12]
rlabel metal3 10777 10360 10777 10360 4 WL[11]
rlabel metal3 10777 9460 10777 9460 4 WL[10]
rlabel metal3 10777 8560 10777 8560 4 WL[9]
rlabel metal3 10777 7660 10777 7660 4 WL[8]
rlabel metal3 8479 11260 8479 11260 4 WL[12]
rlabel metal3 8479 12160 8479 12160 4 WL[13]
rlabel metal3 8479 13060 8479 13060 4 WL[14]
rlabel metal3 8479 13960 8479 13960 4 WL[15]
rlabel metal3 10719 12160 10719 12160 4 WL[13]
rlabel metal3 10719 13960 10719 13960 4 WL[15]
rlabel metal3 9679 7660 9679 7660 4 WL[8]
rlabel metal3 9679 8560 9679 8560 4 WL[9]
rlabel metal3 9679 9460 9679 9460 4 WL[10]
rlabel metal3 9679 10360 9679 10360 4 WL[11]
rlabel metal3 9679 11260 9679 11260 4 WL[12]
rlabel metal3 9679 12160 9679 12160 4 WL[13]
rlabel metal3 9679 13060 9679 13060 4 WL[14]
rlabel metal3 9577 13960 9577 13960 4 WL[15]
rlabel metal3 9577 13060 9577 13060 4 WL[14]
rlabel metal3 9577 12160 9577 12160 4 WL[13]
rlabel metal3 9577 11260 9577 11260 4 WL[12]
rlabel metal3 9577 10360 9577 10360 4 WL[11]
rlabel metal3 9577 9460 9577 9460 4 WL[10]
rlabel metal3 9577 8560 9577 8560 4 WL[9]
rlabel metal3 9577 7660 9577 7660 4 WL[8]
rlabel metal3 9679 13960 9679 13960 4 WL[15]
rlabel metal3 10719 9460 10719 9460 4 WL[10]
rlabel metal3 10719 10360 10719 10360 4 WL[11]
rlabel metal3 10719 11260 10719 11260 4 WL[12]
rlabel metal3 10719 13060 10719 13060 4 WL[14]
rlabel metal3 10177 13960 10177 13960 4 WL[15]
rlabel metal3 10177 13060 10177 13060 4 WL[14]
rlabel metal3 10177 12160 10177 12160 4 WL[13]
rlabel metal3 10177 11260 10177 11260 4 WL[12]
rlabel metal3 10177 10360 10177 10360 4 WL[11]
rlabel metal3 10177 9460 10177 9460 4 WL[10]
rlabel metal3 10177 8560 10177 8560 4 WL[9]
rlabel metal3 10177 7660 10177 7660 4 WL[8]
rlabel metal3 7177 12160 7177 12160 4 WL[13]
rlabel metal3 7177 13060 7177 13060 4 WL[14]
rlabel metal3 7177 10360 7177 10360 4 WL[11]
rlabel metal3 7177 11260 7177 11260 4 WL[12]
rlabel metal3 6079 13960 6079 13960 4 WL[15]
rlabel metal3 6079 12160 6079 12160 4 WL[13]
rlabel metal3 6079 11260 6079 11260 4 WL[12]
rlabel metal3 6079 9460 6079 9460 4 WL[10]
rlabel metal3 6079 8560 6079 8560 4 WL[9]
rlabel metal3 6079 13060 6079 13060 4 WL[14]
rlabel metal3 6079 7660 6079 7660 4 WL[8]
rlabel metal3 7777 10360 7777 10360 4 WL[11]
rlabel metal3 7777 9460 7777 9460 4 WL[10]
rlabel metal3 7777 8560 7777 8560 4 WL[9]
rlabel metal3 6577 9460 6577 9460 4 WL[10]
rlabel metal3 7177 9460 7177 9460 4 WL[10]
rlabel metal3 7177 13960 7177 13960 4 WL[15]
rlabel metal3 7777 13960 7777 13960 4 WL[15]
rlabel metal3 7777 7660 7777 7660 4 WL[8]
rlabel metal3 7177 8560 7177 8560 4 WL[9]
rlabel metal3 7777 13060 7777 13060 4 WL[14]
rlabel metal3 6577 13960 6577 13960 4 WL[15]
rlabel metal3 6577 13060 6577 13060 4 WL[14]
rlabel metal3 6577 12160 6577 12160 4 WL[13]
rlabel metal3 6577 11260 6577 11260 4 WL[12]
rlabel metal3 6577 10360 6577 10360 4 WL[11]
rlabel metal3 6577 8560 6577 8560 4 WL[9]
rlabel metal3 6577 7660 6577 7660 4 WL[8]
rlabel metal3 8377 13960 8377 13960 4 WL[15]
rlabel metal3 8377 13060 8377 13060 4 WL[14]
rlabel metal3 8377 12160 8377 12160 4 WL[13]
rlabel metal3 8377 11260 8377 11260 4 WL[12]
rlabel metal3 8377 10360 8377 10360 4 WL[11]
rlabel metal3 8377 9460 8377 9460 4 WL[10]
rlabel metal3 8377 8560 8377 8560 4 WL[9]
rlabel metal3 8377 7660 8377 7660 4 WL[8]
rlabel metal3 7279 7660 7279 7660 4 WL[8]
rlabel metal3 7279 8560 7279 8560 4 WL[9]
rlabel metal3 7279 9460 7279 9460 4 WL[10]
rlabel metal3 7279 10360 7279 10360 4 WL[11]
rlabel metal3 7279 11260 7279 11260 4 WL[12]
rlabel metal3 7279 12160 7279 12160 4 WL[13]
rlabel metal3 7279 13060 7279 13060 4 WL[14]
rlabel metal3 7279 13960 7279 13960 4 WL[15]
rlabel metal3 7177 7660 7177 7660 4 WL[8]
rlabel metal3 6079 10360 6079 10360 4 WL[11]
rlabel metal3 7777 12160 7777 12160 4 WL[13]
rlabel metal3 7777 11260 7777 11260 4 WL[12]
rlabel metal3 s 8466 5 8466 5 4 VDD
rlabel metal3 7777 5860 7777 5860 4 WL[6]
rlabel metal3 s 7134 918 7134 918 4 VSS
rlabel metal3 7777 2260 7777 2260 4 WL[2]
rlabel metal3 7777 1360 7777 1360 4 WL[1]
rlabel metal3 6079 6760 6079 6760 4 WL[7]
rlabel metal3 6079 5860 6079 5860 4 WL[6]
rlabel metal3 7177 4960 7177 4960 4 WL[5]
rlabel metal3 s 7266 907 7266 907 4 VSS
rlabel metal3 s 7266 5 7266 5 4 VDD
rlabel metal3 s 8334 918 8334 918 4 VSS
rlabel metal3 6079 4960 6079 4960 4 WL[5]
rlabel metal3 6079 4060 6079 4060 4 WL[4]
rlabel metal3 6079 3160 6079 3160 4 WL[3]
rlabel metal3 7177 5860 7177 5860 4 WL[6]
rlabel metal3 6079 2260 6079 2260 4 WL[2]
rlabel metal3 6079 1360 6079 1360 4 WL[1]
rlabel metal3 6079 460 6079 460 4 WL[0]
rlabel metal3 7177 2260 7177 2260 4 WL[2]
rlabel metal3 7177 1360 7177 1360 4 WL[1]
rlabel metal3 7279 460 7279 460 4 WL[0]
rlabel metal3 7279 1360 7279 1360 4 WL[1]
rlabel metal3 7177 4060 7177 4060 4 WL[4]
rlabel metal3 7279 2260 7279 2260 4 WL[2]
rlabel metal3 7279 3160 7279 3160 4 WL[3]
rlabel metal3 7279 4060 7279 4060 4 WL[4]
rlabel metal3 7279 4960 7279 4960 4 WL[5]
rlabel metal3 7279 5860 7279 5860 4 WL[6]
rlabel metal3 7279 6760 7279 6760 4 WL[7]
rlabel metal3 s 6534 -11 6534 -11 4 VDD
rlabel metal3 s 6534 918 6534 918 4 VSS
rlabel metal3 s 6534 -7 6534 -7 4 VDD
rlabel metal3 s 6066 5 6066 5 4 VDD
rlabel metal3 7777 460 7777 460 4 WL[0]
rlabel metal3 s 6066 907 6066 907 4 VSS
rlabel metal3 7177 460 7177 460 4 WL[0]
rlabel metal3 s 7734 -11 7734 -11 4 VDD
rlabel metal3 6577 6760 6577 6760 4 WL[7]
rlabel metal3 6577 5860 6577 5860 4 WL[6]
rlabel metal3 6577 4960 6577 4960 4 WL[5]
rlabel metal3 6577 4060 6577 4060 4 WL[4]
rlabel metal3 s 7734 918 7734 918 4 VSS
rlabel metal3 s 7134 -11 7134 -11 4 VDD
rlabel metal3 8377 6760 8377 6760 4 WL[7]
rlabel metal3 8377 5860 8377 5860 4 WL[6]
rlabel metal3 8377 4960 8377 4960 4 WL[5]
rlabel metal3 8377 4060 8377 4060 4 WL[4]
rlabel metal3 8377 3160 8377 3160 4 WL[3]
rlabel metal3 8377 2260 8377 2260 4 WL[2]
rlabel metal3 8377 1360 8377 1360 4 WL[1]
rlabel metal3 8377 460 8377 460 4 WL[0]
rlabel metal3 7777 4060 7777 4060 4 WL[4]
rlabel metal3 7777 3160 7777 3160 4 WL[3]
rlabel metal3 s 7134 918 7134 918 4 VSS
rlabel metal3 s 6534 918 6534 918 4 VSS
rlabel metal3 s 7134 -7 7134 -7 4 VDD
rlabel metal3 6577 3160 6577 3160 4 WL[3]
rlabel metal3 6577 2260 6577 2260 4 WL[2]
rlabel metal3 6577 1360 6577 1360 4 WL[1]
rlabel metal3 s 7734 -7 7734 -7 4 VDD
rlabel metal3 7777 4960 7777 4960 4 WL[5]
rlabel metal3 7177 6760 7177 6760 4 WL[7]
rlabel metal3 7177 3160 7177 3160 4 WL[3]
rlabel metal3 s 8334 -11 8334 -11 4 VDD
rlabel metal3 s 8334 918 8334 918 4 VSS
rlabel metal3 s 8334 -7 8334 -7 4 VDD
rlabel metal3 6577 460 6577 460 4 WL[0]
rlabel metal3 7777 6760 7777 6760 4 WL[7]
rlabel metal3 s 7734 918 7734 918 4 VSS
rlabel metal3 s 8466 907 8466 907 4 VSS
rlabel metal3 9679 4960 9679 4960 4 WL[5]
rlabel metal3 9577 3160 9577 3160 4 WL[3]
rlabel metal3 9679 5860 9679 5860 4 WL[6]
rlabel metal3 8479 6760 8479 6760 4 WL[7]
rlabel metal3 9577 2260 9577 2260 4 WL[2]
rlabel metal3 s 8934 918 8934 918 4 VSS
rlabel metal3 9679 6760 9679 6760 4 WL[7]
rlabel metal3 8977 6760 8977 6760 4 WL[7]
rlabel metal3 8977 5860 8977 5860 4 WL[6]
rlabel metal3 8977 4960 8977 4960 4 WL[5]
rlabel metal3 10719 460 10719 460 4 WL[0]
rlabel metal3 10719 3160 10719 3160 4 WL[3]
rlabel metal3 8977 4060 8977 4060 4 WL[4]
rlabel metal3 8977 3160 8977 3160 4 WL[3]
rlabel metal3 8977 2260 8977 2260 4 WL[2]
rlabel metal3 10719 4960 10719 4960 4 WL[5]
rlabel metal3 8977 1360 8977 1360 4 WL[1]
rlabel metal3 8977 460 8977 460 4 WL[0]
rlabel metal3 9577 1360 9577 1360 4 WL[1]
rlabel metal3 8479 3160 8479 3160 4 WL[3]
rlabel metal3 8479 4060 8479 4060 4 WL[4]
rlabel metal3 9577 460 9577 460 4 WL[0]
rlabel metal3 10719 6760 10719 6760 4 WL[7]
rlabel metal3 9577 4060 9577 4060 4 WL[4]
rlabel metal3 10719 2260 10719 2260 4 WL[2]
rlabel metal3 10719 4060 10719 4060 4 WL[4]
rlabel metal3 9577 6760 9577 6760 4 WL[7]
rlabel metal3 9577 5860 9577 5860 4 WL[6]
rlabel metal3 9577 4960 9577 4960 4 WL[5]
rlabel metal3 s 9534 918 9534 918 4 VSS
rlabel metal3 s 10134 -11 10134 -11 4 VDD
rlabel metal3 9679 460 9679 460 4 WL[0]
rlabel metal3 9679 1360 9679 1360 4 WL[1]
rlabel metal3 8479 460 8479 460 4 WL[0]
rlabel metal3 8479 1360 8479 1360 4 WL[1]
rlabel metal3 s 10734 -11 10734 -11 4 VDD
rlabel metal3 s 10734 918 10734 918 4 VSS
rlabel metal3 s 10734 -7 10734 -7 4 VDD
rlabel metal3 s 10134 918 10134 918 4 VSS
rlabel metal3 8479 2260 8479 2260 4 WL[2]
rlabel metal3 s 8934 -11 8934 -11 4 VDD
rlabel metal3 s 8934 918 8934 918 4 VSS
rlabel metal3 s 8934 -7 8934 -7 4 VDD
rlabel metal3 s 10734 920 10734 920 4 VSS
rlabel metal3 s 9666 907 9666 907 4 VSS
rlabel metal3 s 10134 918 10134 918 4 VSS
rlabel metal3 8479 4960 8479 4960 4 WL[5]
rlabel metal3 s 9666 5 9666 5 4 VDD
rlabel metal3 10719 5860 10719 5860 4 WL[6]
rlabel metal3 s 10134 -7 10134 -7 4 VDD
rlabel metal3 s 10734 918 10734 918 4 VSS
rlabel metal3 10719 1360 10719 1360 4 WL[1]
rlabel metal3 10777 6760 10777 6760 4 WL[7]
rlabel metal3 10777 5860 10777 5860 4 WL[6]
rlabel metal3 9679 2260 9679 2260 4 WL[2]
rlabel metal3 10777 4960 10777 4960 4 WL[5]
rlabel metal3 10777 4060 10777 4060 4 WL[4]
rlabel metal3 10777 3160 10777 3160 4 WL[3]
rlabel metal3 10777 2260 10777 2260 4 WL[2]
rlabel metal3 10777 1360 10777 1360 4 WL[1]
rlabel metal3 10777 460 10777 460 4 WL[0]
rlabel metal3 9679 3160 9679 3160 4 WL[3]
rlabel metal3 8479 5860 8479 5860 4 WL[6]
rlabel metal3 s 9534 -11 9534 -11 4 VDD
rlabel metal3 s 9534 918 9534 918 4 VSS
rlabel metal3 s 9534 -7 9534 -7 4 VDD
rlabel metal3 9679 4060 9679 4060 4 WL[4]
rlabel metal3 10177 6760 10177 6760 4 WL[7]
rlabel metal3 10177 5860 10177 5860 4 WL[6]
rlabel metal3 10177 4960 10177 4960 4 WL[5]
rlabel metal3 10177 4060 10177 4060 4 WL[4]
rlabel metal3 10177 3160 10177 3160 4 WL[3]
rlabel metal3 10177 2260 10177 2260 4 WL[2]
rlabel metal3 10177 1360 10177 1360 4 WL[1]
rlabel metal3 10177 460 10177 460 4 WL[0]
rlabel metal3 21577 24760 21577 24760 4 WL[27]
rlabel metal3 21577 23860 21577 23860 4 WL[26]
rlabel metal3 19777 22960 19777 22960 4 WL[25]
rlabel metal3 19777 22060 19777 22060 4 WL[24]
rlabel metal3 19777 28360 19777 28360 4 WL[31]
rlabel metal3 19777 27460 19777 27460 4 WL[30]
rlabel metal3 19777 26560 19777 26560 4 WL[29]
rlabel metal3 19777 25660 19777 25660 4 WL[28]
rlabel metal3 19777 24760 19777 24760 4 WL[27]
rlabel metal3 19777 23860 19777 23860 4 WL[26]
rlabel metal3 21519 22960 21519 22960 4 WL[25]
rlabel metal3 20977 22960 20977 22960 4 WL[25]
rlabel metal3 20977 22060 20977 22060 4 WL[24]
rlabel metal3 20977 28360 20977 28360 4 WL[31]
rlabel metal3 20977 27460 20977 27460 4 WL[30]
rlabel metal3 20977 26560 20977 26560 4 WL[29]
rlabel metal3 20977 25660 20977 25660 4 WL[28]
rlabel metal3 20977 24760 20977 24760 4 WL[27]
rlabel metal3 20977 23860 20977 23860 4 WL[26]
rlabel metal3 21519 26560 21519 26560 4 WL[29]
rlabel metal3 21519 27460 21519 27460 4 WL[30]
rlabel metal3 20479 23860 20479 23860 4 WL[26]
rlabel metal3 20479 24760 20479 24760 4 WL[27]
rlabel metal3 20479 25660 20479 25660 4 WL[28]
rlabel metal3 20479 26560 20479 26560 4 WL[29]
rlabel metal3 20479 27460 20479 27460 4 WL[30]
rlabel metal3 20479 28360 20479 28360 4 WL[31]
rlabel metal3 19177 22960 19177 22960 4 WL[25]
rlabel metal3 19177 22060 19177 22060 4 WL[24]
rlabel metal3 19177 28360 19177 28360 4 WL[31]
rlabel metal3 19177 27460 19177 27460 4 WL[30]
rlabel metal3 19177 26560 19177 26560 4 WL[29]
rlabel metal3 19177 25660 19177 25660 4 WL[28]
rlabel metal3 19177 24760 19177 24760 4 WL[27]
rlabel metal3 19177 23860 19177 23860 4 WL[26]
rlabel metal3 20479 22060 20479 22060 4 WL[24]
rlabel metal3 20479 22960 20479 22960 4 WL[25]
rlabel metal3 21519 28360 21519 28360 4 WL[31]
rlabel metal3 21519 22060 21519 22060 4 WL[24]
rlabel metal3 21519 23860 21519 23860 4 WL[26]
rlabel metal3 19279 23860 19279 23860 4 WL[26]
rlabel metal3 19279 24760 19279 24760 4 WL[27]
rlabel metal3 19279 25660 19279 25660 4 WL[28]
rlabel metal3 19279 26560 19279 26560 4 WL[29]
rlabel metal3 19279 27460 19279 27460 4 WL[30]
rlabel metal3 19279 28360 19279 28360 4 WL[31]
rlabel metal3 21519 24760 21519 24760 4 WL[27]
rlabel metal3 21519 25660 21519 25660 4 WL[28]
rlabel metal3 19279 22060 19279 22060 4 WL[24]
rlabel metal3 19279 22960 19279 22960 4 WL[25]
rlabel metal3 21577 22960 21577 22960 4 WL[25]
rlabel metal3 21577 22060 21577 22060 4 WL[24]
rlabel metal3 20377 22960 20377 22960 4 WL[25]
rlabel metal3 20377 22060 20377 22060 4 WL[24]
rlabel metal3 20377 28360 20377 28360 4 WL[31]
rlabel metal3 20377 27460 20377 27460 4 WL[30]
rlabel metal3 20377 26560 20377 26560 4 WL[29]
rlabel metal3 20377 25660 20377 25660 4 WL[28]
rlabel metal3 20377 24760 20377 24760 4 WL[27]
rlabel metal3 20377 23860 20377 23860 4 WL[26]
rlabel metal3 21577 28360 21577 28360 4 WL[31]
rlabel metal3 21577 27460 21577 27460 4 WL[30]
rlabel metal3 21577 26560 21577 26560 4 WL[29]
rlabel metal3 21577 25660 21577 25660 4 WL[28]
rlabel metal3 18577 28360 18577 28360 4 WL[31]
rlabel metal3 18577 27460 18577 27460 4 WL[30]
rlabel metal3 18577 26560 18577 26560 4 WL[29]
rlabel metal3 18577 25660 18577 25660 4 WL[28]
rlabel metal3 18577 24760 18577 24760 4 WL[27]
rlabel metal3 18577 23860 18577 23860 4 WL[26]
rlabel metal3 16879 26560 16879 26560 4 WL[29]
rlabel metal3 17977 22960 17977 22960 4 WL[25]
rlabel metal3 17977 24760 17977 24760 4 WL[27]
rlabel metal3 17977 26560 17977 26560 4 WL[29]
rlabel metal3 17977 25660 17977 25660 4 WL[28]
rlabel metal3 16879 22060 16879 22060 4 WL[24]
rlabel metal3 16879 23860 16879 23860 4 WL[26]
rlabel metal3 17977 23860 17977 23860 4 WL[26]
rlabel metal3 17377 24760 17377 24760 4 WL[27]
rlabel metal3 18079 23860 18079 23860 4 WL[26]
rlabel metal3 18079 24760 18079 24760 4 WL[27]
rlabel metal3 17377 22060 17377 22060 4 WL[24]
rlabel metal3 16879 27460 16879 27460 4 WL[30]
rlabel metal3 16879 22960 16879 22960 4 WL[25]
rlabel metal3 16879 25660 16879 25660 4 WL[28]
rlabel metal3 17377 27460 17377 27460 4 WL[30]
rlabel metal3 17377 23860 17377 23860 4 WL[26]
rlabel metal3 17377 25660 17377 25660 4 WL[28]
rlabel metal3 18079 25660 18079 25660 4 WL[28]
rlabel metal3 18079 26560 18079 26560 4 WL[29]
rlabel metal3 18079 27460 18079 27460 4 WL[30]
rlabel metal3 18079 28360 18079 28360 4 WL[31]
rlabel metal3 17977 28360 17977 28360 4 WL[31]
rlabel metal3 17377 26560 17377 26560 4 WL[29]
rlabel metal3 16879 28360 16879 28360 4 WL[31]
rlabel metal3 18079 22060 18079 22060 4 WL[24]
rlabel metal3 18079 22960 18079 22960 4 WL[25]
rlabel metal3 17377 28360 17377 28360 4 WL[31]
rlabel metal3 17977 27460 17977 27460 4 WL[30]
rlabel metal3 16879 24760 16879 24760 4 WL[27]
rlabel metal3 17977 22060 17977 22060 4 WL[24]
rlabel metal3 18577 22960 18577 22960 4 WL[25]
rlabel metal3 18577 22060 18577 22060 4 WL[24]
rlabel metal3 17377 22960 17377 22960 4 WL[25]
rlabel metal3 18079 16660 18079 16660 4 WL[18]
rlabel metal3 16879 19360 16879 19360 4 WL[21]
rlabel metal3 18079 17560 18079 17560 4 WL[19]
rlabel metal3 18079 18460 18079 18460 4 WL[20]
rlabel metal3 17377 14860 17377 14860 4 WL[16]
rlabel metal3 17377 15760 17377 15760 4 WL[17]
rlabel metal3 17377 16660 17377 16660 4 WL[18]
rlabel metal3 17377 17560 17377 17560 4 WL[19]
rlabel metal3 18079 19360 18079 19360 4 WL[21]
rlabel metal3 17377 21160 17377 21160 4 WL[23]
rlabel metal3 18079 20260 18079 20260 4 WL[22]
rlabel metal3 18079 21160 18079 21160 4 WL[23]
rlabel metal3 16879 20260 16879 20260 4 WL[22]
rlabel metal3 18577 21160 18577 21160 4 WL[23]
rlabel metal3 18577 20260 18577 20260 4 WL[22]
rlabel metal3 17377 18460 17377 18460 4 WL[20]
rlabel metal3 18577 19360 18577 19360 4 WL[21]
rlabel metal3 17977 17560 17977 17560 4 WL[19]
rlabel metal3 18577 18460 18577 18460 4 WL[20]
rlabel metal3 18577 17560 18577 17560 4 WL[19]
rlabel metal3 18577 16660 18577 16660 4 WL[18]
rlabel metal3 18577 15760 18577 15760 4 WL[17]
rlabel metal3 18577 14860 18577 14860 4 WL[16]
rlabel metal3 17377 19360 17377 19360 4 WL[21]
rlabel metal3 17977 19360 17977 19360 4 WL[21]
rlabel metal3 17977 16660 17977 16660 4 WL[18]
rlabel metal3 17977 21160 17977 21160 4 WL[23]
rlabel metal3 17977 20260 17977 20260 4 WL[22]
rlabel metal3 16879 18460 16879 18460 4 WL[20]
rlabel metal3 17977 18460 17977 18460 4 WL[20]
rlabel metal3 16879 14860 16879 14860 4 WL[16]
rlabel metal3 17377 20260 17377 20260 4 WL[22]
rlabel metal3 16879 17560 16879 17560 4 WL[19]
rlabel metal3 17977 14860 17977 14860 4 WL[16]
rlabel metal3 16879 21160 16879 21160 4 WL[23]
rlabel metal3 17977 15760 17977 15760 4 WL[17]
rlabel metal3 16879 16660 16879 16660 4 WL[18]
rlabel metal3 18079 14860 18079 14860 4 WL[16]
rlabel metal3 16879 15760 16879 15760 4 WL[17]
rlabel metal3 18079 15760 18079 15760 4 WL[17]
rlabel metal3 20479 21160 20479 21160 4 WL[23]
rlabel metal3 20977 14860 20977 14860 4 WL[16]
rlabel metal3 19777 18460 19777 18460 4 WL[20]
rlabel metal3 19777 17560 19777 17560 4 WL[19]
rlabel metal3 19279 14860 19279 14860 4 WL[16]
rlabel metal3 19279 15760 19279 15760 4 WL[17]
rlabel metal3 19279 16660 19279 16660 4 WL[18]
rlabel metal3 19279 17560 19279 17560 4 WL[19]
rlabel metal3 19279 18460 19279 18460 4 WL[20]
rlabel metal3 19279 19360 19279 19360 4 WL[21]
rlabel metal3 19279 20260 19279 20260 4 WL[22]
rlabel metal3 19279 21160 19279 21160 4 WL[23]
rlabel metal3 21519 17560 21519 17560 4 WL[19]
rlabel metal3 21519 20260 21519 20260 4 WL[22]
rlabel metal3 21519 14860 21519 14860 4 WL[16]
rlabel metal3 19777 16660 19777 16660 4 WL[18]
rlabel metal3 19777 15760 19777 15760 4 WL[17]
rlabel metal3 21519 19360 21519 19360 4 WL[21]
rlabel metal3 19777 14860 19777 14860 4 WL[16]
rlabel metal3 21519 16660 21519 16660 4 WL[18]
rlabel metal3 21519 18460 21519 18460 4 WL[20]
rlabel metal3 19777 21160 19777 21160 4 WL[23]
rlabel metal3 21519 21160 21519 21160 4 WL[23]
rlabel metal3 19777 20260 19777 20260 4 WL[22]
rlabel metal3 21519 15760 21519 15760 4 WL[17]
rlabel metal3 19777 19360 19777 19360 4 WL[21]
rlabel metal3 20977 21160 20977 21160 4 WL[23]
rlabel metal3 19177 21160 19177 21160 4 WL[23]
rlabel metal3 19177 20260 19177 20260 4 WL[22]
rlabel metal3 19177 19360 19177 19360 4 WL[21]
rlabel metal3 21577 21160 21577 21160 4 WL[23]
rlabel metal3 21577 20260 21577 20260 4 WL[22]
rlabel metal3 21577 19360 21577 19360 4 WL[21]
rlabel metal3 21577 18460 21577 18460 4 WL[20]
rlabel metal3 21577 17560 21577 17560 4 WL[19]
rlabel metal3 21577 16660 21577 16660 4 WL[18]
rlabel metal3 21577 15760 21577 15760 4 WL[17]
rlabel metal3 21577 14860 21577 14860 4 WL[16]
rlabel metal3 19177 18460 19177 18460 4 WL[20]
rlabel metal3 19177 17560 19177 17560 4 WL[19]
rlabel metal3 20377 21160 20377 21160 4 WL[23]
rlabel metal3 20377 20260 20377 20260 4 WL[22]
rlabel metal3 20377 19360 20377 19360 4 WL[21]
rlabel metal3 20377 18460 20377 18460 4 WL[20]
rlabel metal3 20377 17560 20377 17560 4 WL[19]
rlabel metal3 20377 16660 20377 16660 4 WL[18]
rlabel metal3 20377 15760 20377 15760 4 WL[17]
rlabel metal3 20377 14860 20377 14860 4 WL[16]
rlabel metal3 19177 16660 19177 16660 4 WL[18]
rlabel metal3 19177 15760 19177 15760 4 WL[17]
rlabel metal3 19177 14860 19177 14860 4 WL[16]
rlabel metal3 20977 20260 20977 20260 4 WL[22]
rlabel metal3 20977 19360 20977 19360 4 WL[21]
rlabel metal3 20977 18460 20977 18460 4 WL[20]
rlabel metal3 20977 17560 20977 17560 4 WL[19]
rlabel metal3 20977 16660 20977 16660 4 WL[18]
rlabel metal3 20977 15760 20977 15760 4 WL[17]
rlabel metal3 20479 14860 20479 14860 4 WL[16]
rlabel metal3 20479 15760 20479 15760 4 WL[17]
rlabel metal3 20479 16660 20479 16660 4 WL[18]
rlabel metal3 20479 17560 20479 17560 4 WL[19]
rlabel metal3 20479 18460 20479 18460 4 WL[20]
rlabel metal3 20479 19360 20479 19360 4 WL[21]
rlabel metal3 20479 20260 20479 20260 4 WL[22]
rlabel metal3 14423 26560 14423 26560 4 WL[29]
rlabel metal3 14423 25660 14423 25660 4 WL[28]
rlabel metal3 14423 24760 14423 24760 4 WL[27]
rlabel metal3 14423 23860 14423 23860 4 WL[26]
rlabel metal3 16121 22060 16121 22060 4 WL[24]
rlabel metal3 16121 22960 16121 22960 4 WL[25]
rlabel metal3 15623 22960 15623 22960 4 WL[25]
rlabel metal3 15623 22060 15623 22060 4 WL[24]
rlabel metal3 15623 28360 15623 28360 4 WL[31]
rlabel metal3 15623 27460 15623 27460 4 WL[30]
rlabel metal3 15623 26560 15623 26560 4 WL[29]
rlabel metal3 15623 25660 15623 25660 4 WL[28]
rlabel metal3 15623 24760 15623 24760 4 WL[27]
rlabel metal3 15623 23860 15623 23860 4 WL[26]
rlabel metal3 16121 23860 16121 23860 4 WL[26]
rlabel metal3 16121 24760 16121 24760 4 WL[27]
rlabel metal3 14921 23860 14921 23860 4 WL[26]
rlabel metal3 14921 24760 14921 24760 4 WL[27]
rlabel metal3 14921 25660 14921 25660 4 WL[28]
rlabel metal3 14921 26560 14921 26560 4 WL[29]
rlabel metal3 14921 27460 14921 27460 4 WL[30]
rlabel metal3 14921 28360 14921 28360 4 WL[31]
rlabel metal3 16121 25660 16121 25660 4 WL[28]
rlabel metal3 16121 26560 16121 26560 4 WL[29]
rlabel metal3 14921 22060 14921 22060 4 WL[24]
rlabel metal3 14921 22960 14921 22960 4 WL[25]
rlabel metal3 16121 27460 16121 27460 4 WL[30]
rlabel metal3 16121 28360 16121 28360 4 WL[31]
rlabel metal3 15023 22960 15023 22960 4 WL[25]
rlabel metal3 15023 22060 15023 22060 4 WL[24]
rlabel metal3 13823 22960 13823 22960 4 WL[25]
rlabel metal3 13823 22060 13823 22060 4 WL[24]
rlabel metal3 13823 28360 13823 28360 4 WL[31]
rlabel metal3 13823 27460 13823 27460 4 WL[30]
rlabel metal3 13823 26560 13823 26560 4 WL[29]
rlabel metal3 13823 25660 13823 25660 4 WL[28]
rlabel metal3 13823 24760 13823 24760 4 WL[27]
rlabel metal3 13823 23860 13823 23860 4 WL[26]
rlabel metal3 15023 28360 15023 28360 4 WL[31]
rlabel metal3 15023 27460 15023 27460 4 WL[30]
rlabel metal3 15023 26560 15023 26560 4 WL[29]
rlabel metal3 15023 25660 15023 25660 4 WL[28]
rlabel metal3 15023 24760 15023 24760 4 WL[27]
rlabel metal3 15023 23860 15023 23860 4 WL[26]
rlabel metal3 14423 22960 14423 22960 4 WL[25]
rlabel metal3 14423 22060 14423 22060 4 WL[24]
rlabel metal3 14423 28360 14423 28360 4 WL[31]
rlabel metal3 14423 27460 14423 27460 4 WL[30]
rlabel metal3 13223 22060 13223 22060 4 WL[24]
rlabel metal3 13721 28360 13721 28360 4 WL[31]
rlabel metal3 13721 23860 13721 23860 4 WL[26]
rlabel metal3 13223 28360 13223 28360 4 WL[31]
rlabel metal3 13223 27460 13223 27460 4 WL[30]
rlabel metal3 13223 26560 13223 26560 4 WL[29]
rlabel metal3 13223 25660 13223 25660 4 WL[28]
rlabel metal3 13223 24760 13223 24760 4 WL[27]
rlabel metal3 13223 23860 13223 23860 4 WL[26]
rlabel metal3 13721 24760 13721 24760 4 WL[27]
rlabel metal3 13721 25660 13721 25660 4 WL[28]
rlabel metal3 11481 22060 11481 22060 4 WL[24]
rlabel metal3 12521 23860 12521 23860 4 WL[26]
rlabel metal3 12521 24760 12521 24760 4 WL[27]
rlabel metal3 12521 25660 12521 25660 4 WL[28]
rlabel metal3 12521 26560 12521 26560 4 WL[29]
rlabel metal3 12521 27460 12521 27460 4 WL[30]
rlabel metal3 12521 28360 12521 28360 4 WL[31]
rlabel metal3 11481 22960 11481 22960 4 WL[25]
rlabel metal3 12521 22060 12521 22060 4 WL[24]
rlabel metal3 12521 22960 12521 22960 4 WL[25]
rlabel metal3 13721 22060 13721 22060 4 WL[24]
rlabel metal3 13721 22960 13721 22960 4 WL[25]
rlabel metal3 11481 28360 11481 28360 4 WL[31]
rlabel metal3 11423 22960 11423 22960 4 WL[25]
rlabel metal3 11423 22060 11423 22060 4 WL[24]
rlabel metal3 11481 27460 11481 27460 4 WL[30]
rlabel metal3 11481 26560 11481 26560 4 WL[29]
rlabel metal3 11481 25660 11481 25660 4 WL[28]
rlabel metal3 12623 22960 12623 22960 4 WL[25]
rlabel metal3 12623 22060 12623 22060 4 WL[24]
rlabel metal3 11423 28360 11423 28360 4 WL[31]
rlabel metal3 11423 27460 11423 27460 4 WL[30]
rlabel metal3 11423 26560 11423 26560 4 WL[29]
rlabel metal3 11423 25660 11423 25660 4 WL[28]
rlabel metal3 11423 24760 11423 24760 4 WL[27]
rlabel metal3 11423 23860 11423 23860 4 WL[26]
rlabel metal3 11481 24760 11481 24760 4 WL[27]
rlabel metal3 12623 28360 12623 28360 4 WL[31]
rlabel metal3 12623 27460 12623 27460 4 WL[30]
rlabel metal3 12623 26560 12623 26560 4 WL[29]
rlabel metal3 12623 25660 12623 25660 4 WL[28]
rlabel metal3 12623 24760 12623 24760 4 WL[27]
rlabel metal3 12623 23860 12623 23860 4 WL[26]
rlabel metal3 11481 23860 11481 23860 4 WL[26]
rlabel metal3 13721 26560 13721 26560 4 WL[29]
rlabel metal3 12023 22960 12023 22960 4 WL[25]
rlabel metal3 12023 22060 12023 22060 4 WL[24]
rlabel metal3 12023 28360 12023 28360 4 WL[31]
rlabel metal3 12023 27460 12023 27460 4 WL[30]
rlabel metal3 12023 26560 12023 26560 4 WL[29]
rlabel metal3 12023 25660 12023 25660 4 WL[28]
rlabel metal3 12023 24760 12023 24760 4 WL[27]
rlabel metal3 12023 23860 12023 23860 4 WL[26]
rlabel metal3 13721 27460 13721 27460 4 WL[30]
rlabel metal3 13223 22960 13223 22960 4 WL[25]
rlabel metal3 12521 19360 12521 19360 4 WL[21]
rlabel metal3 12521 20260 12521 20260 4 WL[22]
rlabel metal3 12521 21160 12521 21160 4 WL[23]
rlabel metal3 12623 21160 12623 21160 4 WL[23]
rlabel metal3 13223 21160 13223 21160 4 WL[23]
rlabel metal3 13223 20260 13223 20260 4 WL[22]
rlabel metal3 13223 19360 13223 19360 4 WL[21]
rlabel metal3 13223 18460 13223 18460 4 WL[20]
rlabel metal3 13223 17560 13223 17560 4 WL[19]
rlabel metal3 13223 16660 13223 16660 4 WL[18]
rlabel metal3 11423 21160 11423 21160 4 WL[23]
rlabel metal3 11423 20260 11423 20260 4 WL[22]
rlabel metal3 11423 19360 11423 19360 4 WL[21]
rlabel metal3 11423 18460 11423 18460 4 WL[20]
rlabel metal3 11423 17560 11423 17560 4 WL[19]
rlabel metal3 11423 16660 11423 16660 4 WL[18]
rlabel metal3 11423 15760 11423 15760 4 WL[17]
rlabel metal3 11423 14860 11423 14860 4 WL[16]
rlabel metal3 13223 15760 13223 15760 4 WL[17]
rlabel metal3 13223 14860 13223 14860 4 WL[16]
rlabel metal3 12623 20260 12623 20260 4 WL[22]
rlabel metal3 12623 19360 12623 19360 4 WL[21]
rlabel metal3 12623 18460 12623 18460 4 WL[20]
rlabel metal3 12623 17560 12623 17560 4 WL[19]
rlabel metal3 12623 16660 12623 16660 4 WL[18]
rlabel metal3 12623 15760 12623 15760 4 WL[17]
rlabel metal3 12623 14860 12623 14860 4 WL[16]
rlabel metal3 11481 16660 11481 16660 4 WL[18]
rlabel metal3 11481 15760 11481 15760 4 WL[17]
rlabel metal3 13721 14860 13721 14860 4 WL[16]
rlabel metal3 13721 15760 13721 15760 4 WL[17]
rlabel metal3 11481 21160 11481 21160 4 WL[23]
rlabel metal3 11481 20260 11481 20260 4 WL[22]
rlabel metal3 13721 16660 13721 16660 4 WL[18]
rlabel metal3 13721 17560 13721 17560 4 WL[19]
rlabel metal3 13721 18460 13721 18460 4 WL[20]
rlabel metal3 13721 19360 13721 19360 4 WL[21]
rlabel metal3 13721 20260 13721 20260 4 WL[22]
rlabel metal3 13721 21160 13721 21160 4 WL[23]
rlabel metal3 11481 19360 11481 19360 4 WL[21]
rlabel metal3 12023 21160 12023 21160 4 WL[23]
rlabel metal3 12023 20260 12023 20260 4 WL[22]
rlabel metal3 12023 19360 12023 19360 4 WL[21]
rlabel metal3 12023 18460 12023 18460 4 WL[20]
rlabel metal3 12023 17560 12023 17560 4 WL[19]
rlabel metal3 12023 16660 12023 16660 4 WL[18]
rlabel metal3 12023 15760 12023 15760 4 WL[17]
rlabel metal3 12023 14860 12023 14860 4 WL[16]
rlabel metal3 11481 18460 11481 18460 4 WL[20]
rlabel metal3 11481 17560 11481 17560 4 WL[19]
rlabel metal3 11481 14860 11481 14860 4 WL[16]
rlabel metal3 12521 14860 12521 14860 4 WL[16]
rlabel metal3 12521 15760 12521 15760 4 WL[17]
rlabel metal3 12521 16660 12521 16660 4 WL[18]
rlabel metal3 12521 17560 12521 17560 4 WL[19]
rlabel metal3 12521 18460 12521 18460 4 WL[20]
rlabel metal3 14921 19360 14921 19360 4 WL[21]
rlabel metal3 16121 18460 16121 18460 4 WL[20]
rlabel metal3 14921 20260 14921 20260 4 WL[22]
rlabel metal3 15623 18460 15623 18460 4 WL[20]
rlabel metal3 15623 17560 15623 17560 4 WL[19]
rlabel metal3 15623 16660 15623 16660 4 WL[18]
rlabel metal3 15623 15760 15623 15760 4 WL[17]
rlabel metal3 15623 14860 15623 14860 4 WL[16]
rlabel metal3 16121 21160 16121 21160 4 WL[23]
rlabel metal3 16121 19360 16121 19360 4 WL[21]
rlabel metal3 15023 21160 15023 21160 4 WL[23]
rlabel metal3 15023 20260 15023 20260 4 WL[22]
rlabel metal3 15023 19360 15023 19360 4 WL[21]
rlabel metal3 15023 18460 15023 18460 4 WL[20]
rlabel metal3 15023 17560 15023 17560 4 WL[19]
rlabel metal3 15023 16660 15023 16660 4 WL[18]
rlabel metal3 15023 15760 15023 15760 4 WL[17]
rlabel metal3 15023 14860 15023 14860 4 WL[16]
rlabel metal3 16121 15760 16121 15760 4 WL[17]
rlabel metal3 16121 20260 16121 20260 4 WL[22]
rlabel metal3 15623 21160 15623 21160 4 WL[23]
rlabel metal3 13823 21160 13823 21160 4 WL[23]
rlabel metal3 14423 21160 14423 21160 4 WL[23]
rlabel metal3 14423 20260 14423 20260 4 WL[22]
rlabel metal3 14423 19360 14423 19360 4 WL[21]
rlabel metal3 13823 20260 13823 20260 4 WL[22]
rlabel metal3 13823 19360 13823 19360 4 WL[21]
rlabel metal3 13823 18460 13823 18460 4 WL[20]
rlabel metal3 13823 17560 13823 17560 4 WL[19]
rlabel metal3 13823 16660 13823 16660 4 WL[18]
rlabel metal3 13823 15760 13823 15760 4 WL[17]
rlabel metal3 13823 14860 13823 14860 4 WL[16]
rlabel metal3 16121 16660 16121 16660 4 WL[18]
rlabel metal3 16121 17560 16121 17560 4 WL[19]
rlabel metal3 15623 20260 15623 20260 4 WL[22]
rlabel metal3 14423 18460 14423 18460 4 WL[20]
rlabel metal3 14423 17560 14423 17560 4 WL[19]
rlabel metal3 14423 16660 14423 16660 4 WL[18]
rlabel metal3 14423 15760 14423 15760 4 WL[17]
rlabel metal3 14423 14860 14423 14860 4 WL[16]
rlabel metal3 14921 21160 14921 21160 4 WL[23]
rlabel metal3 15623 19360 15623 19360 4 WL[21]
rlabel metal3 14921 14860 14921 14860 4 WL[16]
rlabel metal3 14921 15760 14921 15760 4 WL[17]
rlabel metal3 16121 14860 16121 14860 4 WL[16]
rlabel metal3 14921 16660 14921 16660 4 WL[18]
rlabel metal3 14921 17560 14921 17560 4 WL[19]
rlabel metal3 14921 18460 14921 18460 4 WL[20]
rlabel metal3 16121 8560 16121 8560 4 WL[9]
rlabel metal3 16121 9460 16121 9460 4 WL[10]
rlabel metal3 16121 10360 16121 10360 4 WL[11]
rlabel metal3 16121 11260 16121 11260 4 WL[12]
rlabel metal3 16121 12160 16121 12160 4 WL[13]
rlabel metal3 16121 13060 16121 13060 4 WL[14]
rlabel metal3 16121 13960 16121 13960 4 WL[15]
rlabel metal3 15623 13960 15623 13960 4 WL[15]
rlabel metal3 15623 13060 15623 13060 4 WL[14]
rlabel metal3 15623 12160 15623 12160 4 WL[13]
rlabel metal3 15623 11260 15623 11260 4 WL[12]
rlabel metal3 15623 10360 15623 10360 4 WL[11]
rlabel metal3 15623 9460 15623 9460 4 WL[10]
rlabel metal3 13823 13960 13823 13960 4 WL[15]
rlabel metal3 13823 13060 13823 13060 4 WL[14]
rlabel metal3 13823 12160 13823 12160 4 WL[13]
rlabel metal3 13823 11260 13823 11260 4 WL[12]
rlabel metal3 13823 10360 13823 10360 4 WL[11]
rlabel metal3 13823 9460 13823 9460 4 WL[10]
rlabel metal3 13823 8560 13823 8560 4 WL[9]
rlabel metal3 13823 7660 13823 7660 4 WL[8]
rlabel metal3 15623 8560 15623 8560 4 WL[9]
rlabel metal3 15623 7660 15623 7660 4 WL[8]
rlabel metal3 15023 13960 15023 13960 4 WL[15]
rlabel metal3 15023 13060 15023 13060 4 WL[14]
rlabel metal3 15023 12160 15023 12160 4 WL[13]
rlabel metal3 15023 11260 15023 11260 4 WL[12]
rlabel metal3 14423 13960 14423 13960 4 WL[15]
rlabel metal3 14423 13060 14423 13060 4 WL[14]
rlabel metal3 14423 12160 14423 12160 4 WL[13]
rlabel metal3 14423 11260 14423 11260 4 WL[12]
rlabel metal3 14423 10360 14423 10360 4 WL[11]
rlabel metal3 14423 9460 14423 9460 4 WL[10]
rlabel metal3 14423 8560 14423 8560 4 WL[9]
rlabel metal3 14423 7660 14423 7660 4 WL[8]
rlabel metal3 15023 10360 15023 10360 4 WL[11]
rlabel metal3 15023 9460 15023 9460 4 WL[10]
rlabel metal3 15023 8560 15023 8560 4 WL[9]
rlabel metal3 15023 7660 15023 7660 4 WL[8]
rlabel metal3 14921 7660 14921 7660 4 WL[8]
rlabel metal3 14921 8560 14921 8560 4 WL[9]
rlabel metal3 14921 9460 14921 9460 4 WL[10]
rlabel metal3 14921 10360 14921 10360 4 WL[11]
rlabel metal3 14921 11260 14921 11260 4 WL[12]
rlabel metal3 14921 12160 14921 12160 4 WL[13]
rlabel metal3 14921 13060 14921 13060 4 WL[14]
rlabel metal3 14921 13960 14921 13960 4 WL[15]
rlabel metal3 16121 7660 16121 7660 4 WL[8]
rlabel metal3 12623 7660 12623 7660 4 WL[8]
rlabel metal3 12623 13960 12623 13960 4 WL[15]
rlabel metal3 12623 13060 12623 13060 4 WL[14]
rlabel metal3 12623 12160 12623 12160 4 WL[13]
rlabel metal3 13223 13960 13223 13960 4 WL[15]
rlabel metal3 13223 13060 13223 13060 4 WL[14]
rlabel metal3 12521 7660 12521 7660 4 WL[8]
rlabel metal3 12521 8560 12521 8560 4 WL[9]
rlabel metal3 12521 9460 12521 9460 4 WL[10]
rlabel metal3 12521 10360 12521 10360 4 WL[11]
rlabel metal3 12521 11260 12521 11260 4 WL[12]
rlabel metal3 12521 12160 12521 12160 4 WL[13]
rlabel metal3 12521 13060 12521 13060 4 WL[14]
rlabel metal3 12521 13960 12521 13960 4 WL[15]
rlabel metal3 13223 12160 13223 12160 4 WL[13]
rlabel metal3 13223 11260 13223 11260 4 WL[12]
rlabel metal3 13223 10360 13223 10360 4 WL[11]
rlabel metal3 13223 9460 13223 9460 4 WL[10]
rlabel metal3 13223 8560 13223 8560 4 WL[9]
rlabel metal3 13223 7660 13223 7660 4 WL[8]
rlabel metal3 11481 11260 11481 11260 4 WL[12]
rlabel metal3 11481 10360 11481 10360 4 WL[11]
rlabel metal3 11481 9460 11481 9460 4 WL[10]
rlabel metal3 11423 13960 11423 13960 4 WL[15]
rlabel metal3 11423 13060 11423 13060 4 WL[14]
rlabel metal3 11423 12160 11423 12160 4 WL[13]
rlabel metal3 11423 11260 11423 11260 4 WL[12]
rlabel metal3 11423 10360 11423 10360 4 WL[11]
rlabel metal3 11423 9460 11423 9460 4 WL[10]
rlabel metal3 11423 8560 11423 8560 4 WL[9]
rlabel metal3 11423 7660 11423 7660 4 WL[8]
rlabel metal3 13721 7660 13721 7660 4 WL[8]
rlabel metal3 13721 8560 13721 8560 4 WL[9]
rlabel metal3 13721 9460 13721 9460 4 WL[10]
rlabel metal3 13721 10360 13721 10360 4 WL[11]
rlabel metal3 13721 11260 13721 11260 4 WL[12]
rlabel metal3 13721 12160 13721 12160 4 WL[13]
rlabel metal3 13721 13060 13721 13060 4 WL[14]
rlabel metal3 13721 13960 13721 13960 4 WL[15]
rlabel metal3 11481 8560 11481 8560 4 WL[9]
rlabel metal3 11481 7660 11481 7660 4 WL[8]
rlabel metal3 12623 11260 12623 11260 4 WL[12]
rlabel metal3 12623 10360 12623 10360 4 WL[11]
rlabel metal3 12623 9460 12623 9460 4 WL[10]
rlabel metal3 11481 13960 11481 13960 4 WL[15]
rlabel metal3 11481 13060 11481 13060 4 WL[14]
rlabel metal3 11481 12160 11481 12160 4 WL[13]
rlabel metal3 12023 13960 12023 13960 4 WL[15]
rlabel metal3 12023 13060 12023 13060 4 WL[14]
rlabel metal3 12023 12160 12023 12160 4 WL[13]
rlabel metal3 12023 11260 12023 11260 4 WL[12]
rlabel metal3 12023 10360 12023 10360 4 WL[11]
rlabel metal3 12023 9460 12023 9460 4 WL[10]
rlabel metal3 12023 8560 12023 8560 4 WL[9]
rlabel metal3 12023 7660 12023 7660 4 WL[8]
rlabel metal3 12623 8560 12623 8560 4 WL[9]
rlabel metal3 s 12534 5 12534 5 4 VDD
rlabel metal3 s 11466 918 11466 918 4 VSS
rlabel metal3 s 13266 -7 13266 -7 4 VDD
rlabel metal3 11481 6760 11481 6760 4 WL[7]
rlabel metal3 11481 5860 11481 5860 4 WL[6]
rlabel metal3 13721 460 13721 460 4 WL[0]
rlabel metal3 13721 1360 13721 1360 4 WL[1]
rlabel metal3 13721 2260 13721 2260 4 WL[2]
rlabel metal3 13721 3160 13721 3160 4 WL[3]
rlabel metal3 13721 4060 13721 4060 4 WL[4]
rlabel metal3 13721 4960 13721 4960 4 WL[5]
rlabel metal3 13721 5860 13721 5860 4 WL[6]
rlabel metal3 12623 3160 12623 3160 4 WL[3]
rlabel metal3 12623 2260 12623 2260 4 WL[2]
rlabel metal3 12623 1360 12623 1360 4 WL[1]
rlabel metal3 12623 460 12623 460 4 WL[0]
rlabel metal3 s 12666 -11 12666 -11 4 VDD
rlabel metal3 s 12666 918 12666 918 4 VSS
rlabel metal3 s 12666 -7 12666 -7 4 VDD
rlabel metal3 13223 6760 13223 6760 4 WL[7]
rlabel metal3 11423 6760 11423 6760 4 WL[7]
rlabel metal3 11423 5860 11423 5860 4 WL[6]
rlabel metal3 11423 4960 11423 4960 4 WL[5]
rlabel metal3 11423 4060 11423 4060 4 WL[4]
rlabel metal3 11423 3160 11423 3160 4 WL[3]
rlabel metal3 11423 2260 11423 2260 4 WL[2]
rlabel metal3 11423 1360 11423 1360 4 WL[1]
rlabel metal3 11423 460 11423 460 4 WL[0]
rlabel metal3 13721 6760 13721 6760 4 WL[7]
rlabel metal3 13223 5860 13223 5860 4 WL[6]
rlabel metal3 13223 4960 13223 4960 4 WL[5]
rlabel metal3 12521 460 12521 460 4 WL[0]
rlabel metal3 12521 1360 12521 1360 4 WL[1]
rlabel metal3 12521 2260 12521 2260 4 WL[2]
rlabel metal3 12521 3160 12521 3160 4 WL[3]
rlabel metal3 12521 4060 12521 4060 4 WL[4]
rlabel metal3 12521 4960 12521 4960 4 WL[5]
rlabel metal3 12521 5860 12521 5860 4 WL[6]
rlabel metal3 12521 6760 12521 6760 4 WL[7]
rlabel metal3 13223 4060 13223 4060 4 WL[4]
rlabel metal3 13223 3160 13223 3160 4 WL[3]
rlabel metal3 13223 2260 13223 2260 4 WL[2]
rlabel metal3 s 11466 -11 11466 -11 4 VDD
rlabel metal3 s 11466 918 11466 918 4 VSS
rlabel metal3 s 11466 -7 11466 -7 4 VDD
rlabel metal3 s 12066 918 12066 918 4 VSS
rlabel metal3 11481 4960 11481 4960 4 WL[5]
rlabel metal3 11481 4060 11481 4060 4 WL[4]
rlabel metal3 11481 3160 11481 3160 4 WL[3]
rlabel metal3 11481 2260 11481 2260 4 WL[2]
rlabel metal3 11481 1360 11481 1360 4 WL[1]
rlabel metal3 11481 460 11481 460 4 WL[0]
rlabel metal3 13223 1360 13223 1360 4 WL[1]
rlabel metal3 13223 460 13223 460 4 WL[0]
rlabel metal3 12623 6760 12623 6760 4 WL[7]
rlabel metal3 s 13266 918 13266 918 4 VSS
rlabel metal3 12623 5860 12623 5860 4 WL[6]
rlabel metal3 s 11466 920 11466 920 4 VSS
rlabel metal3 s 11466 2 11466 2 4 VDD
rlabel metal3 12623 4960 12623 4960 4 WL[5]
rlabel metal3 12623 4060 12623 4060 4 WL[4]
rlabel metal3 s 13266 -11 13266 -11 4 VDD
rlabel metal3 s 13266 918 13266 918 4 VSS
rlabel metal3 12023 6760 12023 6760 4 WL[7]
rlabel metal3 12023 5860 12023 5860 4 WL[6]
rlabel metal3 12023 4960 12023 4960 4 WL[5]
rlabel metal3 12023 4060 12023 4060 4 WL[4]
rlabel metal3 12023 3160 12023 3160 4 WL[3]
rlabel metal3 12023 2260 12023 2260 4 WL[2]
rlabel metal3 12023 1360 12023 1360 4 WL[1]
rlabel metal3 12023 460 12023 460 4 WL[0]
rlabel metal3 s 12666 918 12666 918 4 VSS
rlabel metal3 s 12066 -11 12066 -11 4 VDD
rlabel metal3 s 12066 918 12066 918 4 VSS
rlabel metal3 s 12066 -7 12066 -7 4 VDD
rlabel metal3 s 12534 907 12534 907 4 VSS
rlabel metal3 13823 4960 13823 4960 4 WL[5]
rlabel metal3 13823 4060 13823 4060 4 WL[4]
rlabel metal3 15023 6760 15023 6760 4 WL[7]
rlabel metal3 15023 5860 15023 5860 4 WL[6]
rlabel metal3 s 14466 -11 14466 -11 4 VDD
rlabel metal3 s 14466 918 14466 918 4 VSS
rlabel metal3 s 14466 -7 14466 -7 4 VDD
rlabel metal3 15023 4960 15023 4960 4 WL[5]
rlabel metal3 15023 4060 15023 4060 4 WL[4]
rlabel metal3 15023 3160 15023 3160 4 WL[3]
rlabel metal3 13823 3160 13823 3160 4 WL[3]
rlabel metal3 13823 2260 13823 2260 4 WL[2]
rlabel metal3 15023 2260 15023 2260 4 WL[2]
rlabel metal3 13823 1360 13823 1360 4 WL[1]
rlabel metal3 14921 460 14921 460 4 WL[0]
rlabel metal3 14921 1360 14921 1360 4 WL[1]
rlabel metal3 14921 2260 14921 2260 4 WL[2]
rlabel metal3 15023 1360 15023 1360 4 WL[1]
rlabel metal3 14921 3160 14921 3160 4 WL[3]
rlabel metal3 15023 460 15023 460 4 WL[0]
rlabel metal3 14921 4060 14921 4060 4 WL[4]
rlabel metal3 14921 4960 14921 4960 4 WL[5]
rlabel metal3 14921 5860 14921 5860 4 WL[6]
rlabel metal3 14921 6760 14921 6760 4 WL[7]
rlabel metal3 13823 460 13823 460 4 WL[0]
rlabel metal3 13823 6760 13823 6760 4 WL[7]
rlabel metal3 13823 5860 13823 5860 4 WL[6]
rlabel metal3 15623 6760 15623 6760 4 WL[7]
rlabel metal3 15623 5860 15623 5860 4 WL[6]
rlabel metal3 16121 460 16121 460 4 WL[0]
rlabel metal3 16121 1360 16121 1360 4 WL[1]
rlabel metal3 16121 2260 16121 2260 4 WL[2]
rlabel metal3 s 15066 -11 15066 -11 4 VDD
rlabel metal3 s 15066 918 15066 918 4 VSS
rlabel metal3 s 14934 907 14934 907 4 VSS
rlabel metal3 s 14934 5 14934 5 4 VDD
rlabel metal3 s 13866 918 13866 918 4 VSS
rlabel metal3 s 15066 -7 15066 -7 4 VDD
rlabel metal3 15623 4960 15623 4960 4 WL[5]
rlabel metal3 15623 4060 15623 4060 4 WL[4]
rlabel metal3 15623 3160 15623 3160 4 WL[3]
rlabel metal3 15623 2260 15623 2260 4 WL[2]
rlabel metal3 15623 1360 15623 1360 4 WL[1]
rlabel metal3 s 13866 -11 13866 -11 4 VDD
rlabel metal3 s 15666 -11 15666 -11 4 VDD
rlabel metal3 s 15666 918 15666 918 4 VSS
rlabel metal3 s 13866 918 13866 918 4 VSS
rlabel metal3 s 13866 -7 13866 -7 4 VDD
rlabel metal3 14423 6760 14423 6760 4 WL[7]
rlabel metal3 14423 5860 14423 5860 4 WL[6]
rlabel metal3 14423 4960 14423 4960 4 WL[5]
rlabel metal3 14423 4060 14423 4060 4 WL[4]
rlabel metal3 14423 3160 14423 3160 4 WL[3]
rlabel metal3 14423 2260 14423 2260 4 WL[2]
rlabel metal3 16121 3160 16121 3160 4 WL[3]
rlabel metal3 s 15666 918 15666 918 4 VSS
rlabel metal3 16121 4060 16121 4060 4 WL[4]
rlabel metal3 s 13734 907 13734 907 4 VSS
rlabel metal3 s 13734 5 13734 5 4 VDD
rlabel metal3 14423 1360 14423 1360 4 WL[1]
rlabel metal3 s 16134 907 16134 907 4 VSS
rlabel metal3 s 16134 5 16134 5 4 VDD
rlabel metal3 s 15066 918 15066 918 4 VSS
rlabel metal3 16121 4960 16121 4960 4 WL[5]
rlabel metal3 16121 5860 16121 5860 4 WL[6]
rlabel metal3 14423 460 14423 460 4 WL[0]
rlabel metal3 s 15666 -7 15666 -7 4 VDD
rlabel metal3 s 14466 918 14466 918 4 VSS
rlabel metal3 16121 6760 16121 6760 4 WL[7]
rlabel metal3 15623 460 15623 460 4 WL[0]
rlabel metal3 20479 11260 20479 11260 4 WL[12]
rlabel metal3 20479 12160 20479 12160 4 WL[13]
rlabel metal3 20479 13060 20479 13060 4 WL[14]
rlabel metal3 19279 12160 19279 12160 4 WL[13]
rlabel metal3 19279 13060 19279 13060 4 WL[14]
rlabel metal3 19279 13960 19279 13960 4 WL[15]
rlabel metal3 20479 13960 20479 13960 4 WL[15]
rlabel metal3 21519 13060 21519 13060 4 WL[14]
rlabel metal3 21519 13960 21519 13960 4 WL[15]
rlabel metal3 21519 8560 21519 8560 4 WL[9]
rlabel metal3 21519 7660 21519 7660 4 WL[8]
rlabel metal3 19777 13960 19777 13960 4 WL[15]
rlabel metal3 19777 13060 19777 13060 4 WL[14]
rlabel metal3 19777 12160 19777 12160 4 WL[13]
rlabel metal3 19777 11260 19777 11260 4 WL[12]
rlabel metal3 19777 10360 19777 10360 4 WL[11]
rlabel metal3 21519 9460 21519 9460 4 WL[10]
rlabel metal3 21519 10360 21519 10360 4 WL[11]
rlabel metal3 21519 11260 21519 11260 4 WL[12]
rlabel metal3 21519 12160 21519 12160 4 WL[13]
rlabel metal3 19777 9460 19777 9460 4 WL[10]
rlabel metal3 19777 8560 19777 8560 4 WL[9]
rlabel metal3 19777 7660 19777 7660 4 WL[8]
rlabel metal3 21577 13960 21577 13960 4 WL[15]
rlabel metal3 21577 13060 21577 13060 4 WL[14]
rlabel metal3 21577 12160 21577 12160 4 WL[13]
rlabel metal3 21577 11260 21577 11260 4 WL[12]
rlabel metal3 21577 10360 21577 10360 4 WL[11]
rlabel metal3 21577 9460 21577 9460 4 WL[10]
rlabel metal3 21577 8560 21577 8560 4 WL[9]
rlabel metal3 21577 7660 21577 7660 4 WL[8]
rlabel metal3 19177 13960 19177 13960 4 WL[15]
rlabel metal3 19177 13060 19177 13060 4 WL[14]
rlabel metal3 19177 12160 19177 12160 4 WL[13]
rlabel metal3 19177 11260 19177 11260 4 WL[12]
rlabel metal3 19177 10360 19177 10360 4 WL[11]
rlabel metal3 20977 13960 20977 13960 4 WL[15]
rlabel metal3 20977 13060 20977 13060 4 WL[14]
rlabel metal3 19177 9460 19177 9460 4 WL[10]
rlabel metal3 19177 8560 19177 8560 4 WL[9]
rlabel metal3 19177 7660 19177 7660 4 WL[8]
rlabel metal3 20377 13960 20377 13960 4 WL[15]
rlabel metal3 20377 13060 20377 13060 4 WL[14]
rlabel metal3 20377 12160 20377 12160 4 WL[13]
rlabel metal3 20377 11260 20377 11260 4 WL[12]
rlabel metal3 20377 10360 20377 10360 4 WL[11]
rlabel metal3 20377 9460 20377 9460 4 WL[10]
rlabel metal3 20377 8560 20377 8560 4 WL[9]
rlabel metal3 20377 7660 20377 7660 4 WL[8]
rlabel metal3 20479 7660 20479 7660 4 WL[8]
rlabel metal3 20479 8560 20479 8560 4 WL[9]
rlabel metal3 20977 12160 20977 12160 4 WL[13]
rlabel metal3 20977 11260 20977 11260 4 WL[12]
rlabel metal3 20977 10360 20977 10360 4 WL[11]
rlabel metal3 20479 9460 20479 9460 4 WL[10]
rlabel metal3 20479 10360 20479 10360 4 WL[11]
rlabel metal3 20977 9460 20977 9460 4 WL[10]
rlabel metal3 20977 8560 20977 8560 4 WL[9]
rlabel metal3 20977 7660 20977 7660 4 WL[8]
rlabel metal3 19279 7660 19279 7660 4 WL[8]
rlabel metal3 19279 8560 19279 8560 4 WL[9]
rlabel metal3 19279 9460 19279 9460 4 WL[10]
rlabel metal3 19279 10360 19279 10360 4 WL[11]
rlabel metal3 19279 11260 19279 11260 4 WL[12]
rlabel metal3 17977 11260 17977 11260 4 WL[12]
rlabel metal3 17977 13960 17977 13960 4 WL[15]
rlabel metal3 17977 13060 17977 13060 4 WL[14]
rlabel metal3 17377 10360 17377 10360 4 WL[11]
rlabel metal3 16879 13060 16879 13060 4 WL[14]
rlabel metal3 18079 9460 18079 9460 4 WL[10]
rlabel metal3 16879 11260 16879 11260 4 WL[12]
rlabel metal3 18079 10360 18079 10360 4 WL[11]
rlabel metal3 18079 11260 18079 11260 4 WL[12]
rlabel metal3 16879 12160 16879 12160 4 WL[13]
rlabel metal3 17377 12160 17377 12160 4 WL[13]
rlabel metal3 18079 12160 18079 12160 4 WL[13]
rlabel metal3 17377 13960 17377 13960 4 WL[15]
rlabel metal3 16879 10360 16879 10360 4 WL[11]
rlabel metal3 18079 13060 18079 13060 4 WL[14]
rlabel metal3 18079 7660 18079 7660 4 WL[8]
rlabel metal3 16879 7660 16879 7660 4 WL[8]
rlabel metal3 18079 8560 18079 8560 4 WL[9]
rlabel metal3 18079 13960 18079 13960 4 WL[15]
rlabel metal3 16879 8560 16879 8560 4 WL[9]
rlabel metal3 17977 10360 17977 10360 4 WL[11]
rlabel metal3 17977 12160 17977 12160 4 WL[13]
rlabel metal3 18577 13960 18577 13960 4 WL[15]
rlabel metal3 18577 13060 18577 13060 4 WL[14]
rlabel metal3 18577 12160 18577 12160 4 WL[13]
rlabel metal3 16879 9460 16879 9460 4 WL[10]
rlabel metal3 16879 13960 16879 13960 4 WL[15]
rlabel metal3 17377 9460 17377 9460 4 WL[10]
rlabel metal3 17977 9460 17977 9460 4 WL[10]
rlabel metal3 17977 8560 17977 8560 4 WL[9]
rlabel metal3 17377 11260 17377 11260 4 WL[12]
rlabel metal3 17377 13060 17377 13060 4 WL[14]
rlabel metal3 17377 7660 17377 7660 4 WL[8]
rlabel metal3 17377 8560 17377 8560 4 WL[9]
rlabel metal3 17977 7660 17977 7660 4 WL[8]
rlabel metal3 18577 11260 18577 11260 4 WL[12]
rlabel metal3 18577 10360 18577 10360 4 WL[11]
rlabel metal3 18577 9460 18577 9460 4 WL[10]
rlabel metal3 18577 8560 18577 8560 4 WL[9]
rlabel metal3 18577 7660 18577 7660 4 WL[8]
rlabel metal3 s 17334 -7 17334 -7 4 VDD
rlabel metal3 s 17934 -11 17934 -11 4 VDD
rlabel metal3 17377 1360 17377 1360 4 WL[1]
rlabel metal3 s 17334 918 17334 918 4 VSS
rlabel metal3 17377 3160 17377 3160 4 WL[3]
rlabel metal3 17977 1360 17977 1360 4 WL[1]
rlabel metal3 17377 4060 17377 4060 4 WL[4]
rlabel metal3 18079 460 18079 460 4 WL[0]
rlabel metal3 16879 5860 16879 5860 4 WL[6]
rlabel metal3 17977 5860 17977 5860 4 WL[6]
rlabel metal3 16879 6760 16879 6760 4 WL[7]
rlabel metal3 s 17334 918 17334 918 4 VSS
rlabel metal3 s 17934 918 17934 918 4 VSS
rlabel metal3 17977 4960 17977 4960 4 WL[5]
rlabel metal3 s 17334 -11 17334 -11 4 VDD
rlabel metal3 16879 4960 16879 4960 4 WL[5]
rlabel metal3 s 16866 5 16866 5 4 VDD
rlabel metal3 17977 6760 17977 6760 4 WL[7]
rlabel metal3 s 17934 -7 17934 -7 4 VDD
rlabel metal3 18079 1360 18079 1360 4 WL[1]
rlabel metal3 18079 2260 18079 2260 4 WL[2]
rlabel metal3 18079 3160 18079 3160 4 WL[3]
rlabel metal3 s 18534 918 18534 918 4 VSS
rlabel metal3 17377 4960 17377 4960 4 WL[5]
rlabel metal3 18079 4060 18079 4060 4 WL[4]
rlabel metal3 18079 4960 18079 4960 4 WL[5]
rlabel metal3 s 18066 907 18066 907 4 VSS
rlabel metal3 s 18066 5 18066 5 4 VDD
rlabel metal3 18079 5860 18079 5860 4 WL[6]
rlabel metal3 18079 6760 18079 6760 4 WL[7]
rlabel metal3 16879 1360 16879 1360 4 WL[1]
rlabel metal3 s 18534 -11 18534 -11 4 VDD
rlabel metal3 s 18534 918 18534 918 4 VSS
rlabel metal3 s 18534 -7 18534 -7 4 VDD
rlabel metal3 17977 3160 17977 3160 4 WL[3]
rlabel metal3 16879 4060 16879 4060 4 WL[4]
rlabel metal3 17977 460 17977 460 4 WL[0]
rlabel metal3 17377 5860 17377 5860 4 WL[6]
rlabel metal3 17377 6760 17377 6760 4 WL[7]
rlabel metal3 s 17934 918 17934 918 4 VSS
rlabel metal3 16879 2260 16879 2260 4 WL[2]
rlabel metal3 17377 2260 17377 2260 4 WL[2]
rlabel metal3 18577 6760 18577 6760 4 WL[7]
rlabel metal3 18577 5860 18577 5860 4 WL[6]
rlabel metal3 18577 4960 18577 4960 4 WL[5]
rlabel metal3 18577 4060 18577 4060 4 WL[4]
rlabel metal3 18577 3160 18577 3160 4 WL[3]
rlabel metal3 18577 2260 18577 2260 4 WL[2]
rlabel metal3 s 16866 907 16866 907 4 VSS
rlabel metal3 17977 2260 17977 2260 4 WL[2]
rlabel metal3 18577 1360 18577 1360 4 WL[1]
rlabel metal3 18577 460 18577 460 4 WL[0]
rlabel metal3 17977 4060 17977 4060 4 WL[4]
rlabel metal3 16879 3160 16879 3160 4 WL[3]
rlabel metal3 16879 460 16879 460 4 WL[0]
rlabel metal3 17377 460 17377 460 4 WL[0]
rlabel metal3 21519 6760 21519 6760 4 WL[7]
rlabel metal3 s 19734 918 19734 918 4 VSS
rlabel metal3 s 19734 -7 19734 -7 4 VDD
rlabel metal3 21519 460 21519 460 4 WL[0]
rlabel metal3 s 21534 920 21534 920 4 VSS
rlabel metal3 s 21534 -7 21534 -7 4 VDD
rlabel metal3 s 20934 -11 20934 -11 4 VDD
rlabel metal3 21519 2260 21519 2260 4 WL[2]
rlabel metal3 s 20934 918 20934 918 4 VSS
rlabel metal3 21519 4960 21519 4960 4 WL[5]
rlabel metal3 20977 3160 20977 3160 4 WL[3]
rlabel metal3 20977 4060 20977 4060 4 WL[4]
rlabel metal3 21519 4060 21519 4060 4 WL[4]
rlabel metal3 21577 6760 21577 6760 4 WL[7]
rlabel metal3 21577 5860 21577 5860 4 WL[6]
rlabel metal3 19177 6760 19177 6760 4 WL[7]
rlabel metal3 19177 5860 19177 5860 4 WL[6]
rlabel metal3 19177 4960 19177 4960 4 WL[5]
rlabel metal3 21577 4960 21577 4960 4 WL[5]
rlabel metal3 19177 4060 19177 4060 4 WL[4]
rlabel metal3 21577 4060 21577 4060 4 WL[4]
rlabel metal3 21577 3160 21577 3160 4 WL[3]
rlabel metal3 21577 2260 21577 2260 4 WL[2]
rlabel metal3 21577 1360 21577 1360 4 WL[1]
rlabel metal3 21577 460 21577 460 4 WL[0]
rlabel metal3 s 20934 -7 20934 -7 4 VDD
rlabel metal3 20977 2260 20977 2260 4 WL[2]
rlabel metal3 20377 6760 20377 6760 4 WL[7]
rlabel metal3 20377 5860 20377 5860 4 WL[6]
rlabel metal3 20377 4960 20377 4960 4 WL[5]
rlabel metal3 20377 4060 20377 4060 4 WL[4]
rlabel metal3 20377 3160 20377 3160 4 WL[3]
rlabel metal3 20377 2260 20377 2260 4 WL[2]
rlabel metal3 20377 1360 20377 1360 4 WL[1]
rlabel metal3 20377 460 20377 460 4 WL[0]
rlabel metal3 19177 3160 19177 3160 4 WL[3]
rlabel metal3 19177 2260 19177 2260 4 WL[2]
rlabel metal3 19177 1360 19177 1360 4 WL[1]
rlabel metal3 19177 460 19177 460 4 WL[0]
rlabel metal3 20479 4060 20479 4060 4 WL[4]
rlabel metal3 20479 4960 20479 4960 4 WL[5]
rlabel metal3 21519 1360 21519 1360 4 WL[1]
rlabel metal3 21519 3160 21519 3160 4 WL[3]
rlabel metal3 20977 1360 20977 1360 4 WL[1]
rlabel metal3 s 19134 918 19134 918 4 VSS
rlabel metal3 s 19134 -7 19134 -7 4 VDD
rlabel metal3 20479 5860 20479 5860 4 WL[6]
rlabel metal3 20479 6760 20479 6760 4 WL[7]
rlabel metal3 20479 460 20479 460 4 WL[0]
rlabel metal3 20479 1360 20479 1360 4 WL[1]
rlabel metal3 20479 2260 20479 2260 4 WL[2]
rlabel metal3 19777 6760 19777 6760 4 WL[7]
rlabel metal3 19777 5860 19777 5860 4 WL[6]
rlabel metal3 20479 3160 20479 3160 4 WL[3]
rlabel metal3 s 21534 -11 21534 -11 4 VDD
rlabel metal3 19777 4960 19777 4960 4 WL[5]
rlabel metal3 19777 4060 19777 4060 4 WL[4]
rlabel metal3 19777 3160 19777 3160 4 WL[3]
rlabel metal3 s 19266 907 19266 907 4 VSS
rlabel metal3 s 19134 -11 19134 -11 4 VDD
rlabel metal3 s 19266 5 19266 5 4 VDD
rlabel metal3 19777 2260 19777 2260 4 WL[2]
rlabel metal3 s 21534 918 21534 918 4 VSS
rlabel metal3 s 20334 918 20334 918 4 VSS
rlabel metal3 s 20934 918 20934 918 4 VSS
rlabel metal3 20977 6760 20977 6760 4 WL[7]
rlabel metal3 s 20466 907 20466 907 4 VSS
rlabel metal3 s 20466 5 20466 5 4 VDD
rlabel metal3 19777 1360 19777 1360 4 WL[1]
rlabel metal3 s 21534 918 21534 918 4 VSS
rlabel metal3 21519 5860 21519 5860 4 WL[6]
rlabel metal3 19279 460 19279 460 4 WL[0]
rlabel metal3 19279 1360 19279 1360 4 WL[1]
rlabel metal3 19279 2260 19279 2260 4 WL[2]
rlabel metal3 19279 3160 19279 3160 4 WL[3]
rlabel metal3 s 20334 -11 20334 -11 4 VDD
rlabel metal3 19279 4060 19279 4060 4 WL[4]
rlabel metal3 19279 4960 19279 4960 4 WL[5]
rlabel metal3 19279 5860 19279 5860 4 WL[6]
rlabel metal3 19279 6760 19279 6760 4 WL[7]
rlabel metal3 19777 460 19777 460 4 WL[0]
rlabel metal3 20977 460 20977 460 4 WL[0]
rlabel metal3 s 20334 918 20334 918 4 VSS
rlabel metal3 s 20334 -7 20334 -7 4 VDD
rlabel metal3 20977 4960 20977 4960 4 WL[5]
rlabel metal3 s 19134 918 19134 918 4 VSS
rlabel metal3 s 19734 -11 19734 -11 4 VDD
rlabel metal3 20977 5860 20977 5860 4 WL[6]
rlabel metal3 s 19734 918 19734 918 4 VSS
rlabel metal3 s 685 41859 685 41859 4 WL[46]
port 1 nsew
rlabel metal3 s 685 31959 685 31959 4 WL[35]
port 2 nsew
rlabel metal3 s 685 30159 685 30159 4 WL[33]
port 3 nsew
rlabel metal3 s 685 44559 685 44559 4 WL[49]
port 4 nsew
rlabel metal3 s 685 40959 685 40959 4 WL[45]
port 5 nsew
rlabel metal3 s 685 36459 685 36459 4 WL[40]
port 6 nsew
rlabel metal3 s 685 35559 685 35559 4 WL[39]
port 7 nsew
rlabel metal3 s 685 29259 685 29259 4 WL[32]
port 8 nsew
rlabel metal3 s 685 49059 685 49059 4 WL[54]
port 9 nsew
rlabel metal3 s 685 34659 685 34659 4 WL[38]
port 10 nsew
rlabel metal3 s 685 33759 685 33759 4 WL[37]
port 11 nsew
rlabel metal3 s 685 40059 685 40059 4 WL[44]
port 12 nsew
rlabel metal3 s 685 43659 685 43659 4 WL[48]
port 13 nsew
rlabel metal3 s 685 31059 685 31059 4 WL[34]
port 14 nsew
rlabel metal3 s 685 32859 685 32859 4 WL[36]
port 15 nsew
rlabel metal3 s 685 39159 685 39159 4 WL[43]
port 16 nsew
rlabel metal3 s 685 42759 685 42759 4 WL[47]
port 17 nsew
rlabel metal3 s 685 48159 685 48159 4 WL[53]
port 18 nsew
rlabel metal3 s 685 45459 685 45459 4 WL[50]
port 19 nsew
rlabel metal3 s 685 41859 685 41859 4 WL[46]
port 1 nsew
rlabel metal3 s 685 38259 685 38259 4 WL[42]
port 20 nsew
rlabel metal3 s 685 47259 685 47259 4 WL[52]
port 21 nsew
rlabel metal3 s 685 55359 685 55359 4 WL[61]
port 22 nsew
rlabel metal3 s 685 46359 685 46359 4 WL[51]
port 23 nsew
rlabel metal3 s 685 37359 685 37359 4 WL[41]
port 24 nsew
rlabel metal3 s 685 46359 685 46359 4 WL[51]
port 23 nsew
rlabel metal3 s 685 29259 685 29259 4 WL[32]
port 8 nsew
rlabel metal3 s 685 37359 685 37359 4 WL[41]
port 24 nsew
rlabel metal3 s 685 34659 685 34659 4 WL[38]
port 10 nsew
rlabel metal3 s 685 32859 685 32859 4 WL[36]
port 15 nsew
rlabel metal3 s 685 57159 685 57159 4 WL[63]
port 25 nsew
rlabel metal3 s 685 52659 685 52659 4 WL[58]
port 26 nsew
rlabel metal3 s 685 56259 685 56259 4 WL[62]
port 27 nsew
rlabel metal3 s 685 38259 685 38259 4 WL[42]
port 20 nsew
rlabel metal3 s 685 53559 685 53559 4 WL[59]
port 28 nsew
rlabel metal3 s 685 40959 685 40959 4 WL[45]
port 5 nsew
rlabel metal3 s 685 50859 685 50859 4 WL[56]
port 29 nsew
rlabel metal3 s 685 39159 685 39159 4 WL[43]
port 16 nsew
rlabel metal3 s 685 40059 685 40059 4 WL[44]
port 12 nsew
rlabel metal3 s 685 36459 685 36459 4 WL[40]
port 6 nsew
rlabel metal3 s 685 33759 685 33759 4 WL[37]
port 11 nsew
rlabel metal3 s 685 31959 685 31959 4 WL[35]
port 2 nsew
rlabel metal3 s 685 35559 685 35559 4 WL[39]
port 7 nsew
rlabel metal3 s 685 31059 685 31059 4 WL[34]
port 14 nsew
rlabel metal3 s 685 30159 685 30159 4 WL[33]
port 3 nsew
rlabel metal3 s 685 50859 685 50859 4 WL[56]
port 29 nsew
rlabel metal3 s 685 51759 685 51759 4 WL[57]
port 30 nsew
rlabel metal3 s 685 52659 685 52659 4 WL[58]
port 26 nsew
rlabel metal3 s 685 53559 685 53559 4 WL[59]
port 28 nsew
rlabel metal3 s 685 54459 685 54459 4 WL[60]
port 31 nsew
rlabel metal3 s 685 56259 685 56259 4 WL[62]
port 27 nsew
rlabel metal3 s 685 57159 685 57159 4 WL[63]
port 25 nsew
rlabel metal3 s 685 43659 685 43659 4 WL[48]
port 13 nsew
rlabel metal3 s 685 44559 685 44559 4 WL[49]
port 4 nsew
rlabel metal3 s 685 45459 685 45459 4 WL[50]
port 19 nsew
rlabel metal3 s 685 47259 685 47259 4 WL[52]
port 21 nsew
rlabel metal3 s 685 48159 685 48159 4 WL[53]
port 18 nsew
rlabel metal3 s 685 49059 685 49059 4 WL[54]
port 9 nsew
rlabel metal3 s 685 42759 685 42759 4 WL[47]
port 17 nsew
rlabel metal3 s 685 49959 685 49959 4 WL[55]
port 32 nsew
rlabel metal3 s 685 49959 685 49959 4 WL[55]
port 32 nsew
rlabel metal3 s 685 55359 685 55359 4 WL[61]
port 22 nsew
rlabel metal3 s 685 54459 685 54459 4 WL[60]
port 31 nsew
rlabel metal3 s 685 51759 685 51759 4 WL[57]
port 30 nsew
rlabel metal3 s 701 5862 701 5862 4 WL[6]
port 33 nsew
rlabel metal3 s 701 26562 701 26562 4 WL[29]
port 34 nsew
rlabel metal3 s 701 17562 701 17562 4 WL[19]
port 35 nsew
rlabel metal3 s 701 6762 701 6762 4 WL[7]
port 36 nsew
rlabel metal3 s 701 7662 701 7662 4 WL[8]
port 37 nsew
rlabel metal3 s 701 21162 701 21162 4 WL[23]
port 38 nsew
rlabel metal3 s 701 18462 701 18462 4 WL[20]
port 39 nsew
rlabel metal3 s 701 24762 701 24762 4 WL[27]
port 40 nsew
rlabel metal3 s 701 22962 701 22962 4 WL[25]
port 41 nsew
rlabel metal3 s 701 8562 701 8562 4 WL[9]
port 42 nsew
rlabel metal3 s 701 1362 701 1362 4 WL[1]
port 43 nsew
rlabel metal3 s 701 20262 701 20262 4 WL[22]
port 44 nsew
rlabel metal3 s 701 27462 701 27462 4 WL[30]
port 45 nsew
rlabel metal3 s 701 26562 701 26562 4 WL[29]
port 34 nsew
rlabel metal3 s 701 22962 701 22962 4 WL[25]
port 41 nsew
rlabel metal3 s 701 22062 701 22062 4 WL[24]
port 46 nsew
rlabel metal3 s 701 21162 701 21162 4 WL[23]
port 38 nsew
rlabel metal3 s 701 20262 701 20262 4 WL[22]
port 44 nsew
rlabel metal3 s 701 18462 701 18462 4 WL[20]
port 39 nsew
rlabel metal3 s 701 24762 701 24762 4 WL[27]
port 40 nsew
rlabel metal3 s 701 27462 701 27462 4 WL[30]
port 45 nsew
rlabel metal3 s 701 16662 701 16662 4 WL[18]
port 47 nsew
rlabel metal3 s 701 7662 701 7662 4 WL[8]
port 37 nsew
rlabel metal3 s 701 28362 701 28362 4 WL[31]
port 48 nsew
rlabel metal3 s 701 9462 701 9462 4 WL[10]
port 49 nsew
rlabel metal3 s 701 12162 701 12162 4 WL[13]
port 50 nsew
rlabel metal3 s 701 13062 701 13062 4 WL[14]
port 51 nsew
rlabel metal3 s 701 14862 701 14862 4 WL[16]
port 52 nsew
rlabel metal3 s 701 15762 701 15762 4 WL[17]
port 53 nsew
rlabel metal3 s 701 23862 701 23862 4 WL[26]
port 54 nsew
rlabel metal3 s 701 17562 701 17562 4 WL[19]
port 35 nsew
rlabel metal3 s 701 23862 701 23862 4 WL[26]
port 54 nsew
rlabel metal3 s 701 10362 701 10362 4 WL[11]
port 55 nsew
rlabel metal3 s 701 13962 701 13962 4 WL[15]
port 56 nsew
rlabel metal3 s 701 8562 701 8562 4 WL[9]
port 42 nsew
rlabel metal3 s 701 462 701 462 4 WL[0]
port 57 nsew
rlabel metal3 s 701 2262 701 2262 4 WL[2]
port 58 nsew
rlabel metal3 s 701 25662 701 25662 4 WL[28]
port 59 nsew
rlabel metal3 s 701 11262 701 11262 4 WL[12]
port 60 nsew
rlabel metal3 s 701 19362 701 19362 4 WL[21]
port 61 nsew
rlabel metal3 s 701 9462 701 9462 4 WL[10]
port 49 nsew
rlabel metal3 s 701 10362 701 10362 4 WL[11]
port 55 nsew
rlabel metal3 s 701 5862 701 5862 4 WL[6]
port 33 nsew
rlabel metal3 s 701 4062 701 4062 4 WL[4]
port 62 nsew
rlabel metal3 s 701 3162 701 3162 4 WL[3]
port 63 nsew
rlabel metal3 s 701 4062 701 4062 4 WL[4]
port 62 nsew
rlabel metal3 s 701 25662 701 25662 4 WL[28]
port 59 nsew
rlabel metal3 s 701 13062 701 13062 4 WL[14]
port 51 nsew
rlabel metal3 s 701 13962 701 13962 4 WL[15]
port 56 nsew
rlabel metal3 s 701 16662 701 16662 4 WL[18]
port 47 nsew
rlabel metal3 s 701 1362 701 1362 4 WL[1]
port 43 nsew
rlabel metal3 s 701 462 701 462 4 WL[0]
port 57 nsew
rlabel metal3 s 701 2262 701 2262 4 WL[2]
port 58 nsew
rlabel metal3 s 701 3162 701 3162 4 WL[3]
port 63 nsew
rlabel metal3 s 701 4962 701 4962 4 WL[5]
port 64 nsew
rlabel metal3 s 701 11262 701 11262 4 WL[12]
port 60 nsew
rlabel metal3 s 701 28362 701 28362 4 WL[31]
port 48 nsew
rlabel metal3 s 701 12162 701 12162 4 WL[13]
port 50 nsew
rlabel metal3 s 701 14862 701 14862 4 WL[16]
port 52 nsew
rlabel metal3 s 701 19362 701 19362 4 WL[21]
port 61 nsew
rlabel metal3 s 701 22062 701 22062 4 WL[24]
port 46 nsew
rlabel metal3 s 701 4962 701 4962 4 WL[5]
port 64 nsew
rlabel metal3 s 701 15762 701 15762 4 WL[17]
port 53 nsew
rlabel metal3 s 701 6762 701 6762 4 WL[7]
port 36 nsew
<< properties >>
string GDS_END 2433720
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 2111642
<< end >>
