magic
tech gf180mcuB
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 453 3670 1094
<< pwell >>
rect -86 -86 3670 453
<< mvnmos >>
rect 128 175 248 333
rect 352 175 472 333
rect 720 170 840 310
rect 944 170 1064 310
rect 1168 170 1288 310
rect 1336 170 1456 310
rect 1592 170 1712 310
rect 1816 170 1936 310
rect 2040 170 2160 310
rect 2264 170 2384 310
rect 2488 170 2608 310
rect 2712 170 2832 310
rect 2972 170 3092 328
rect 3340 69 3460 333
<< mvpmos >>
rect 128 573 228 849
rect 332 573 432 849
rect 724 593 824 793
rect 928 593 1028 793
rect 1132 593 1232 793
rect 1336 593 1436 793
rect 1540 593 1640 793
rect 1888 630 1988 830
rect 2092 630 2192 830
rect 2296 630 2396 830
rect 2500 630 2600 830
rect 2792 630 2892 826
rect 2996 630 3096 826
rect 3344 573 3444 939
<< mvndiff >>
rect 40 320 128 333
rect 40 274 53 320
rect 99 274 128 320
rect 40 175 128 274
rect 248 234 352 333
rect 248 188 277 234
rect 323 188 352 234
rect 248 175 352 188
rect 472 320 560 333
rect 472 274 501 320
rect 547 274 560 320
rect 2892 310 2972 328
rect 472 175 560 274
rect 632 229 720 310
rect 632 183 645 229
rect 691 183 720 229
rect 632 170 720 183
rect 840 297 944 310
rect 840 251 869 297
rect 915 251 944 297
rect 840 170 944 251
rect 1064 297 1168 310
rect 1064 251 1093 297
rect 1139 251 1168 297
rect 1064 170 1168 251
rect 1288 170 1336 310
rect 1456 170 1592 310
rect 1712 229 1816 310
rect 1712 183 1741 229
rect 1787 183 1816 229
rect 1712 170 1816 183
rect 1936 297 2040 310
rect 1936 251 1965 297
rect 2011 251 2040 297
rect 1936 170 2040 251
rect 2160 297 2264 310
rect 2160 251 2189 297
rect 2235 251 2264 297
rect 2160 170 2264 251
rect 2384 297 2488 310
rect 2384 251 2413 297
rect 2459 251 2488 297
rect 2384 170 2488 251
rect 2608 229 2712 310
rect 2608 183 2637 229
rect 2683 183 2712 229
rect 2608 170 2712 183
rect 2832 170 2972 310
rect 3092 315 3180 328
rect 3092 269 3121 315
rect 3167 269 3180 315
rect 3092 170 3180 269
rect 3252 320 3340 333
rect 3252 180 3265 320
rect 3311 180 3340 320
rect 3252 69 3340 180
rect 3460 222 3548 333
rect 3460 82 3489 222
rect 3535 82 3548 222
rect 3460 69 3548 82
<< mvpdiff >>
rect 40 726 128 849
rect 40 586 53 726
rect 99 586 128 726
rect 40 573 128 586
rect 228 836 332 849
rect 228 696 257 836
rect 303 696 332 836
rect 228 573 332 696
rect 432 726 520 849
rect 2660 895 2732 908
rect 2660 849 2673 895
rect 2719 849 2732 895
rect 2660 830 2732 849
rect 1800 817 1888 830
rect 432 586 461 726
rect 507 586 520 726
rect 636 780 724 793
rect 636 734 649 780
rect 695 734 724 780
rect 636 593 724 734
rect 824 746 928 793
rect 824 606 853 746
rect 899 606 928 746
rect 824 593 928 606
rect 1028 746 1132 793
rect 1028 606 1057 746
rect 1103 606 1132 746
rect 1028 593 1132 606
rect 1232 780 1336 793
rect 1232 640 1261 780
rect 1307 640 1336 780
rect 1232 593 1336 640
rect 1436 780 1540 793
rect 1436 734 1465 780
rect 1511 734 1540 780
rect 1436 593 1540 734
rect 1640 780 1728 793
rect 1640 640 1669 780
rect 1715 640 1728 780
rect 1640 593 1728 640
rect 1800 677 1813 817
rect 1859 677 1888 817
rect 1800 630 1888 677
rect 1988 783 2092 830
rect 1988 643 2017 783
rect 2063 643 2092 783
rect 1988 630 2092 643
rect 2192 783 2296 830
rect 2192 643 2221 783
rect 2267 643 2296 783
rect 2192 630 2296 643
rect 2396 689 2500 830
rect 2396 643 2425 689
rect 2471 643 2500 689
rect 2396 630 2500 643
rect 2600 826 2732 830
rect 2600 630 2792 826
rect 2892 689 2996 826
rect 2892 643 2921 689
rect 2967 643 2996 689
rect 2892 630 2996 643
rect 3096 813 3184 826
rect 3096 673 3125 813
rect 3171 673 3184 813
rect 3096 630 3184 673
rect 3256 726 3344 939
rect 432 573 520 586
rect 3256 586 3269 726
rect 3315 586 3344 726
rect 3256 573 3344 586
rect 3444 926 3532 939
rect 3444 786 3473 926
rect 3519 786 3532 926
rect 3444 573 3532 786
<< mvndiffc >>
rect 53 274 99 320
rect 277 188 323 234
rect 501 274 547 320
rect 645 183 691 229
rect 869 251 915 297
rect 1093 251 1139 297
rect 1741 183 1787 229
rect 1965 251 2011 297
rect 2189 251 2235 297
rect 2413 251 2459 297
rect 2637 183 2683 229
rect 3121 269 3167 315
rect 3265 180 3311 320
rect 3489 82 3535 222
<< mvpdiffc >>
rect 53 586 99 726
rect 257 696 303 836
rect 2673 849 2719 895
rect 461 586 507 726
rect 649 734 695 780
rect 853 606 899 746
rect 1057 606 1103 746
rect 1261 640 1307 780
rect 1465 734 1511 780
rect 1669 640 1715 780
rect 1813 677 1859 817
rect 2017 643 2063 783
rect 2221 643 2267 783
rect 2425 643 2471 689
rect 2921 643 2967 689
rect 3125 673 3171 813
rect 3269 586 3315 726
rect 3473 786 3519 926
<< polysilicon >>
rect 332 933 2192 973
rect 3344 939 3444 983
rect 128 849 228 893
rect 332 849 432 933
rect 928 872 1028 885
rect 724 793 824 837
rect 928 826 941 872
rect 987 826 1028 872
rect 928 793 1028 826
rect 1132 793 1232 933
rect 1336 793 1436 837
rect 1540 793 1640 837
rect 1888 830 1988 874
rect 2092 830 2192 933
rect 2296 830 2396 874
rect 2500 830 2600 874
rect 2792 826 2892 870
rect 2996 826 3096 870
rect 128 487 228 573
rect 128 441 142 487
rect 188 441 228 487
rect 128 377 228 441
rect 332 452 432 573
rect 332 406 345 452
rect 391 406 432 452
rect 332 393 432 406
rect 724 523 824 593
rect 724 477 737 523
rect 783 477 824 523
rect 128 333 248 377
rect 352 333 472 393
rect 724 354 824 477
rect 928 501 1028 593
rect 1132 549 1232 593
rect 928 461 1288 501
rect 1168 389 1288 461
rect 720 310 840 354
rect 944 310 1064 354
rect 1168 343 1181 389
rect 1227 343 1288 389
rect 1168 310 1288 343
rect 1336 481 1436 593
rect 1540 549 1640 593
rect 1336 435 1377 481
rect 1423 435 1436 481
rect 1336 354 1436 435
rect 1592 354 1640 549
rect 1888 583 1988 630
rect 1888 537 1901 583
rect 1947 537 1988 583
rect 1888 370 1988 537
rect 2092 490 2192 630
rect 2296 597 2396 630
rect 2296 551 2309 597
rect 2355 551 2396 597
rect 2296 538 2396 551
rect 2500 530 2600 630
rect 2092 450 2384 490
rect 2040 389 2160 402
rect 1336 310 1456 354
rect 1592 310 1712 354
rect 1816 310 1936 370
rect 2040 343 2057 389
rect 2103 343 2160 389
rect 2040 310 2160 343
rect 2264 310 2384 450
rect 2500 484 2541 530
rect 2587 484 2600 530
rect 2500 354 2600 484
rect 2792 402 2892 630
rect 2996 597 3096 630
rect 2996 551 3013 597
rect 3059 551 3096 597
rect 2996 539 3096 551
rect 2712 389 2832 402
rect 2488 310 2608 354
rect 2712 343 2773 389
rect 2819 343 2832 389
rect 2996 372 3092 539
rect 3344 507 3444 573
rect 3150 494 3444 507
rect 3150 448 3163 494
rect 3209 448 3444 494
rect 3150 435 3444 448
rect 2712 310 2832 343
rect 2972 328 3092 372
rect 3340 377 3444 435
rect 3340 333 3460 377
rect 128 131 248 175
rect 352 78 472 175
rect 720 126 840 170
rect 944 78 1064 170
rect 1168 126 1288 170
rect 1336 126 1456 170
rect 352 38 1064 78
rect 1592 78 1712 170
rect 1816 126 1936 170
rect 2040 126 2160 170
rect 2264 126 2384 170
rect 2488 126 2608 170
rect 2712 78 2832 170
rect 2972 126 3092 170
rect 1592 38 2832 78
rect 3340 25 3460 69
<< polycontact >>
rect 941 826 987 872
rect 142 441 188 487
rect 345 406 391 452
rect 737 477 783 523
rect 1181 343 1227 389
rect 1377 435 1423 481
rect 1901 537 1947 583
rect 2309 551 2355 597
rect 2057 343 2103 389
rect 2541 484 2587 530
rect 3013 551 3059 597
rect 2773 343 2819 389
rect 3163 448 3209 494
<< metal1 >>
rect 0 926 3584 1098
rect 0 918 3473 926
rect 257 836 303 918
rect 53 726 99 737
rect 649 780 695 918
rect 257 685 303 696
rect 461 726 507 737
rect 99 588 286 634
rect 53 575 99 586
rect 132 487 194 542
rect 132 441 142 487
rect 188 441 194 487
rect 132 430 194 441
rect 240 452 286 588
rect 649 723 695 734
rect 741 826 941 872
rect 987 826 998 872
rect 741 677 787 826
rect 1261 780 1307 791
rect 507 631 787 677
rect 853 746 915 757
rect 507 586 547 631
rect 240 406 345 452
rect 391 406 402 452
rect 240 337 286 406
rect 42 320 286 337
rect 42 274 53 320
rect 99 291 286 320
rect 461 320 547 586
rect 899 606 915 746
rect 656 523 783 542
rect 656 477 737 523
rect 656 466 783 477
rect 99 274 217 291
rect 461 274 501 320
rect 461 263 547 274
rect 853 297 915 606
rect 853 251 869 297
rect 277 234 323 245
rect 853 240 915 251
rect 1057 746 1103 757
rect 1465 780 1511 918
rect 1813 817 1859 918
rect 2673 895 2719 918
rect 2673 838 2719 849
rect 1465 723 1511 734
rect 1669 780 1715 791
rect 1307 640 1669 675
rect 3125 813 3171 918
rect 1813 666 1859 677
rect 2017 783 2063 794
rect 1261 629 1715 640
rect 1057 583 1103 606
rect 1057 537 1901 583
rect 1947 537 1958 583
rect 1057 308 1104 537
rect 2017 492 2063 643
rect 1971 481 2063 492
rect 1366 435 1377 481
rect 1423 446 2063 481
rect 2189 792 2267 794
rect 2189 783 3059 792
rect 2189 643 2221 783
rect 2267 746 3059 783
rect 2189 632 2267 643
rect 2413 689 2471 700
rect 2413 643 2425 689
rect 1423 435 2011 446
rect 1170 343 1181 389
rect 1227 343 1919 389
rect 1057 297 1139 308
rect 1057 251 1093 297
rect 1057 240 1139 251
rect 277 90 323 188
rect 645 229 691 240
rect 645 90 691 183
rect 1741 229 1787 240
rect 1741 90 1787 183
rect 1873 194 1919 343
rect 1965 297 2011 435
rect 1965 240 2011 251
rect 2057 389 2103 400
rect 2057 194 2103 343
rect 2189 297 2235 632
rect 2189 240 2235 251
rect 2297 551 2309 597
rect 2355 551 2366 597
rect 2297 194 2366 551
rect 2413 297 2471 643
rect 2921 689 2967 700
rect 2921 530 2967 643
rect 3013 597 3059 746
rect 3519 918 3584 926
rect 3473 775 3519 786
rect 3125 662 3171 673
rect 3269 726 3330 737
rect 3013 540 3059 551
rect 3315 586 3330 726
rect 2530 484 2541 530
rect 2587 494 2967 530
rect 2587 484 3163 494
rect 2530 448 3163 484
rect 3209 448 3220 494
rect 2773 389 2876 400
rect 2819 343 2876 389
rect 2773 332 2876 343
rect 2459 251 2471 297
rect 2413 240 2471 251
rect 2830 318 2876 332
rect 2830 242 3014 318
rect 3121 315 3167 448
rect 3269 438 3330 586
rect 3121 258 3167 269
rect 3265 320 3330 438
rect 1873 148 2366 194
rect 2637 229 2683 240
rect 2637 90 2683 183
rect 3311 180 3330 320
rect 3265 169 3330 180
rect 3489 222 3535 233
rect 0 82 3489 90
rect 3535 82 3584 90
rect 0 -90 3584 82
<< labels >>
flabel metal1 s 132 430 194 542 0 FreeSans 200 0 0 0 CLK
port 3 nsew clock input
flabel metal1 s 656 466 783 542 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 3269 438 3330 737 0 FreeSans 200 0 0 0 Q
port 4 nsew default output
flabel metal1 s 2773 332 2876 400 0 FreeSans 200 0 0 0 RN
port 2 nsew default input
flabel metal1 s 0 918 3584 1098 0 FreeSans 200 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 277 240 323 245 0 FreeSans 200 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 6 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 2830 318 2876 332 1 RN
port 2 nsew default input
rlabel metal1 s 2830 242 3014 318 1 RN
port 2 nsew default input
rlabel metal1 s 3265 169 3330 438 1 Q
port 4 nsew default output
rlabel metal1 s 3473 838 3519 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3125 838 3171 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2673 838 2719 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1813 838 1859 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1465 838 1511 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 649 838 695 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 257 838 303 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3473 775 3519 838 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3125 775 3171 838 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1813 775 1859 838 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1465 775 1511 838 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 649 775 695 838 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 257 775 303 838 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3125 723 3171 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1813 723 1859 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1465 723 1511 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 649 723 695 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 257 723 303 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3125 685 3171 723 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1813 685 1859 723 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 257 685 303 723 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3125 666 3171 685 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1813 666 1859 685 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3125 662 3171 666 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2637 233 2683 240 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1741 233 1787 240 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 645 233 691 240 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 277 233 323 240 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3489 90 3535 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2637 90 2683 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1741 90 1787 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 645 90 691 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 277 90 323 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 3584 90 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3584 1008
string GDS_END 613628
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 604760
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
