magic
tech gf180mcuA
magscale 1 5
timestamp 1698431365
use 018SRAM_cell1_512x8m81  018SRAM_cell1_512x8m81_0
timestamp 1698431365
transform 1 0 0 0 -1 450
box -34 -34 334 484
use 018SRAM_cell1_512x8m81  018SRAM_cell1_512x8m81_1
timestamp 1698431365
transform 1 0 0 0 1 450
box -34 -34 334 484
<< properties >>
string GDS_END 515242
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 515140
<< end >>
