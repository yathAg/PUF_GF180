magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -530 4793 759 5011
rect -530 3964 4955 4793
rect -530 3963 4957 3964
rect -530 2692 5176 3963
rect -530 2672 4573 2692
rect -89 2671 2557 2672
rect 2599 2671 4573 2672
rect 2600 2602 4573 2671
rect -530 656 1442 713
rect 3582 679 4118 694
rect 3582 656 5175 679
rect -530 55 5175 656
rect -530 -24 1442 55
<< mvnmos >>
rect 159 5223 279 5451
rect 383 5223 503 5451
rect 1074 5006 1194 5460
rect 1298 5006 1418 5460
rect 1522 5006 1642 5460
rect 1746 5006 1866 5460
rect 1970 5006 2090 5460
rect 2483 5006 2603 5460
rect 2707 5006 2827 5460
rect 2931 5006 3051 5460
rect 3155 5006 3275 5460
rect 3379 5006 3499 5460
rect 3892 5006 4012 5460
rect 4116 5006 4236 5460
rect 4340 5006 4460 5460
rect 4564 5006 4684 5460
rect 390 1847 510 2301
rect 614 1847 734 2301
rect 838 1847 958 2301
rect 1062 1847 1182 2301
rect 1286 1847 1406 2301
rect 1510 1847 1630 2301
rect 1734 1847 1854 2301
rect 2182 1729 2302 2301
rect 2406 1729 2526 2301
rect 2630 1729 2750 2301
rect 2854 1729 2974 2301
rect 3078 1729 3198 2301
rect 3302 1729 3422 2301
rect 3750 1779 3870 2301
rect 3974 1779 4094 2301
rect 171 855 291 1083
rect 395 855 515 1083
rect 619 855 739 1083
rect 843 855 963 1083
rect 1067 855 1187 1083
rect 1616 884 1736 1004
rect 1840 884 1960 1004
rect 2341 884 2461 1004
rect 2565 884 2685 1004
rect 3065 884 3185 1004
rect 3289 884 3409 1004
rect 3790 884 3910 1004
rect 4251 818 4371 1106
<< mvpmos >>
rect 159 4189 279 4871
rect 383 4189 503 4871
rect 1074 4198 1194 4652
rect 1298 4198 1418 4652
rect 1522 4198 1642 4652
rect 1746 4198 1866 4652
rect 2548 4090 2668 4634
rect 2772 4090 2892 4634
rect 2996 4090 3116 4634
rect 3220 4090 3340 4634
rect 3444 4090 3564 4634
rect 3668 4090 3788 4634
rect 3892 4090 4012 4634
rect 4116 4090 4236 4634
rect 4340 4090 4460 4634
rect 4564 4090 4684 4634
rect 166 2811 286 3629
rect 390 2811 510 3629
rect 614 2811 734 3629
rect 838 2811 958 3629
rect 1062 2811 1182 3629
rect 1286 2811 1406 3629
rect 1510 2811 1630 3629
rect 1734 2811 1854 3629
rect 1958 2811 2078 3629
rect 2182 2811 2302 3629
rect 2854 2742 2974 3650
rect 3078 2742 3198 3650
rect 3302 2742 3422 3650
rect 3750 2742 3870 3650
rect 3974 2742 4094 3650
rect 4198 2742 4318 3650
rect 171 118 291 572
rect 395 118 515 572
rect 619 118 739 572
rect 843 118 963 572
rect 1067 118 1187 572
rect 1616 296 1736 536
rect 1840 296 1960 536
rect 2341 296 2461 536
rect 2565 296 2685 536
rect 3065 296 3185 536
rect 3289 296 3409 536
rect 3790 334 3910 574
rect 4251 197 4371 539
rect 4475 197 4595 539
<< mvndiff >>
rect 71 5438 159 5451
rect 71 5392 84 5438
rect 130 5392 159 5438
rect 71 5282 159 5392
rect 71 5236 84 5282
rect 130 5236 159 5282
rect 71 5223 159 5236
rect 279 5438 383 5451
rect 279 5392 308 5438
rect 354 5392 383 5438
rect 279 5282 383 5392
rect 279 5236 308 5282
rect 354 5236 383 5282
rect 279 5223 383 5236
rect 503 5438 591 5451
rect 503 5392 532 5438
rect 578 5392 591 5438
rect 503 5282 591 5392
rect 503 5236 532 5282
rect 578 5236 591 5282
rect 503 5223 591 5236
rect 986 5447 1074 5460
rect 986 5401 999 5447
rect 1045 5401 1074 5447
rect 986 5320 1074 5401
rect 986 5274 999 5320
rect 1045 5274 1074 5320
rect 986 5193 1074 5274
rect 986 5147 999 5193
rect 1045 5147 1074 5193
rect 986 5065 1074 5147
rect 986 5019 999 5065
rect 1045 5019 1074 5065
rect 986 5006 1074 5019
rect 1194 5447 1298 5460
rect 1194 5401 1223 5447
rect 1269 5401 1298 5447
rect 1194 5320 1298 5401
rect 1194 5274 1223 5320
rect 1269 5274 1298 5320
rect 1194 5193 1298 5274
rect 1194 5147 1223 5193
rect 1269 5147 1298 5193
rect 1194 5065 1298 5147
rect 1194 5019 1223 5065
rect 1269 5019 1298 5065
rect 1194 5006 1298 5019
rect 1418 5447 1522 5460
rect 1418 5401 1447 5447
rect 1493 5401 1522 5447
rect 1418 5320 1522 5401
rect 1418 5274 1447 5320
rect 1493 5274 1522 5320
rect 1418 5193 1522 5274
rect 1418 5147 1447 5193
rect 1493 5147 1522 5193
rect 1418 5065 1522 5147
rect 1418 5019 1447 5065
rect 1493 5019 1522 5065
rect 1418 5006 1522 5019
rect 1642 5447 1746 5460
rect 1642 5401 1671 5447
rect 1717 5401 1746 5447
rect 1642 5320 1746 5401
rect 1642 5274 1671 5320
rect 1717 5274 1746 5320
rect 1642 5193 1746 5274
rect 1642 5147 1671 5193
rect 1717 5147 1746 5193
rect 1642 5065 1746 5147
rect 1642 5019 1671 5065
rect 1717 5019 1746 5065
rect 1642 5006 1746 5019
rect 1866 5447 1970 5460
rect 1866 5401 1895 5447
rect 1941 5401 1970 5447
rect 1866 5320 1970 5401
rect 1866 5274 1895 5320
rect 1941 5274 1970 5320
rect 1866 5193 1970 5274
rect 1866 5147 1895 5193
rect 1941 5147 1970 5193
rect 1866 5065 1970 5147
rect 1866 5019 1895 5065
rect 1941 5019 1970 5065
rect 1866 5006 1970 5019
rect 2090 5447 2178 5460
rect 2090 5401 2119 5447
rect 2165 5401 2178 5447
rect 2090 5320 2178 5401
rect 2090 5274 2119 5320
rect 2165 5274 2178 5320
rect 2090 5193 2178 5274
rect 2090 5147 2119 5193
rect 2165 5147 2178 5193
rect 2090 5065 2178 5147
rect 2090 5019 2119 5065
rect 2165 5019 2178 5065
rect 2090 5006 2178 5019
rect 2395 5447 2483 5460
rect 2395 5401 2408 5447
rect 2454 5401 2483 5447
rect 2395 5320 2483 5401
rect 2395 5274 2408 5320
rect 2454 5274 2483 5320
rect 2395 5193 2483 5274
rect 2395 5147 2408 5193
rect 2454 5147 2483 5193
rect 2395 5065 2483 5147
rect 2395 5019 2408 5065
rect 2454 5019 2483 5065
rect 2395 5006 2483 5019
rect 2603 5447 2707 5460
rect 2603 5401 2632 5447
rect 2678 5401 2707 5447
rect 2603 5320 2707 5401
rect 2603 5274 2632 5320
rect 2678 5274 2707 5320
rect 2603 5193 2707 5274
rect 2603 5147 2632 5193
rect 2678 5147 2707 5193
rect 2603 5065 2707 5147
rect 2603 5019 2632 5065
rect 2678 5019 2707 5065
rect 2603 5006 2707 5019
rect 2827 5447 2931 5460
rect 2827 5401 2856 5447
rect 2902 5401 2931 5447
rect 2827 5320 2931 5401
rect 2827 5274 2856 5320
rect 2902 5274 2931 5320
rect 2827 5193 2931 5274
rect 2827 5147 2856 5193
rect 2902 5147 2931 5193
rect 2827 5065 2931 5147
rect 2827 5019 2856 5065
rect 2902 5019 2931 5065
rect 2827 5006 2931 5019
rect 3051 5447 3155 5460
rect 3051 5401 3080 5447
rect 3126 5401 3155 5447
rect 3051 5320 3155 5401
rect 3051 5274 3080 5320
rect 3126 5274 3155 5320
rect 3051 5193 3155 5274
rect 3051 5147 3080 5193
rect 3126 5147 3155 5193
rect 3051 5065 3155 5147
rect 3051 5019 3080 5065
rect 3126 5019 3155 5065
rect 3051 5006 3155 5019
rect 3275 5447 3379 5460
rect 3275 5401 3304 5447
rect 3350 5401 3379 5447
rect 3275 5320 3379 5401
rect 3275 5274 3304 5320
rect 3350 5274 3379 5320
rect 3275 5193 3379 5274
rect 3275 5147 3304 5193
rect 3350 5147 3379 5193
rect 3275 5065 3379 5147
rect 3275 5019 3304 5065
rect 3350 5019 3379 5065
rect 3275 5006 3379 5019
rect 3499 5447 3587 5460
rect 3499 5401 3528 5447
rect 3574 5401 3587 5447
rect 3499 5320 3587 5401
rect 3499 5274 3528 5320
rect 3574 5274 3587 5320
rect 3499 5193 3587 5274
rect 3499 5147 3528 5193
rect 3574 5147 3587 5193
rect 3499 5065 3587 5147
rect 3499 5019 3528 5065
rect 3574 5019 3587 5065
rect 3499 5006 3587 5019
rect 3804 5447 3892 5460
rect 3804 5401 3817 5447
rect 3863 5401 3892 5447
rect 3804 5320 3892 5401
rect 3804 5274 3817 5320
rect 3863 5274 3892 5320
rect 3804 5193 3892 5274
rect 3804 5147 3817 5193
rect 3863 5147 3892 5193
rect 3804 5065 3892 5147
rect 3804 5019 3817 5065
rect 3863 5019 3892 5065
rect 3804 5006 3892 5019
rect 4012 5447 4116 5460
rect 4012 5401 4041 5447
rect 4087 5401 4116 5447
rect 4012 5320 4116 5401
rect 4012 5274 4041 5320
rect 4087 5274 4116 5320
rect 4012 5193 4116 5274
rect 4012 5147 4041 5193
rect 4087 5147 4116 5193
rect 4012 5065 4116 5147
rect 4012 5019 4041 5065
rect 4087 5019 4116 5065
rect 4012 5006 4116 5019
rect 4236 5447 4340 5460
rect 4236 5401 4265 5447
rect 4311 5401 4340 5447
rect 4236 5320 4340 5401
rect 4236 5274 4265 5320
rect 4311 5274 4340 5320
rect 4236 5193 4340 5274
rect 4236 5147 4265 5193
rect 4311 5147 4340 5193
rect 4236 5065 4340 5147
rect 4236 5019 4265 5065
rect 4311 5019 4340 5065
rect 4236 5006 4340 5019
rect 4460 5447 4564 5460
rect 4460 5401 4489 5447
rect 4535 5401 4564 5447
rect 4460 5320 4564 5401
rect 4460 5274 4489 5320
rect 4535 5274 4564 5320
rect 4460 5193 4564 5274
rect 4460 5147 4489 5193
rect 4535 5147 4564 5193
rect 4460 5065 4564 5147
rect 4460 5019 4489 5065
rect 4535 5019 4564 5065
rect 4460 5006 4564 5019
rect 4684 5447 4772 5460
rect 4684 5401 4713 5447
rect 4759 5401 4772 5447
rect 4684 5320 4772 5401
rect 4684 5274 4713 5320
rect 4759 5274 4772 5320
rect 4684 5193 4772 5274
rect 4684 5147 4713 5193
rect 4759 5147 4772 5193
rect 4684 5065 4772 5147
rect 4684 5019 4713 5065
rect 4759 5019 4772 5065
rect 4684 5006 4772 5019
rect 302 2288 390 2301
rect 302 2242 315 2288
rect 361 2242 390 2288
rect 302 2160 390 2242
rect 302 2114 315 2160
rect 361 2114 390 2160
rect 302 2033 390 2114
rect 302 1987 315 2033
rect 361 1987 390 2033
rect 302 1906 390 1987
rect 302 1860 315 1906
rect 361 1860 390 1906
rect 302 1847 390 1860
rect 510 2288 614 2301
rect 510 2242 539 2288
rect 585 2242 614 2288
rect 510 2160 614 2242
rect 510 2114 539 2160
rect 585 2114 614 2160
rect 510 2033 614 2114
rect 510 1987 539 2033
rect 585 1987 614 2033
rect 510 1906 614 1987
rect 510 1860 539 1906
rect 585 1860 614 1906
rect 510 1847 614 1860
rect 734 2288 838 2301
rect 734 2242 763 2288
rect 809 2242 838 2288
rect 734 2160 838 2242
rect 734 2114 763 2160
rect 809 2114 838 2160
rect 734 2033 838 2114
rect 734 1987 763 2033
rect 809 1987 838 2033
rect 734 1906 838 1987
rect 734 1860 763 1906
rect 809 1860 838 1906
rect 734 1847 838 1860
rect 958 2288 1062 2301
rect 958 2242 987 2288
rect 1033 2242 1062 2288
rect 958 2160 1062 2242
rect 958 2114 987 2160
rect 1033 2114 1062 2160
rect 958 2033 1062 2114
rect 958 1987 987 2033
rect 1033 1987 1062 2033
rect 958 1906 1062 1987
rect 958 1860 987 1906
rect 1033 1860 1062 1906
rect 958 1847 1062 1860
rect 1182 2288 1286 2301
rect 1182 2242 1211 2288
rect 1257 2242 1286 2288
rect 1182 2160 1286 2242
rect 1182 2114 1211 2160
rect 1257 2114 1286 2160
rect 1182 2033 1286 2114
rect 1182 1987 1211 2033
rect 1257 1987 1286 2033
rect 1182 1906 1286 1987
rect 1182 1860 1211 1906
rect 1257 1860 1286 1906
rect 1182 1847 1286 1860
rect 1406 2288 1510 2301
rect 1406 2242 1435 2288
rect 1481 2242 1510 2288
rect 1406 2160 1510 2242
rect 1406 2114 1435 2160
rect 1481 2114 1510 2160
rect 1406 2033 1510 2114
rect 1406 1987 1435 2033
rect 1481 1987 1510 2033
rect 1406 1906 1510 1987
rect 1406 1860 1435 1906
rect 1481 1860 1510 1906
rect 1406 1847 1510 1860
rect 1630 2288 1734 2301
rect 1630 2242 1659 2288
rect 1705 2242 1734 2288
rect 1630 2160 1734 2242
rect 1630 2114 1659 2160
rect 1705 2114 1734 2160
rect 1630 2033 1734 2114
rect 1630 1987 1659 2033
rect 1705 1987 1734 2033
rect 1630 1906 1734 1987
rect 1630 1860 1659 1906
rect 1705 1860 1734 1906
rect 1630 1847 1734 1860
rect 1854 2288 1942 2301
rect 1854 2242 1883 2288
rect 1929 2242 1942 2288
rect 1854 2160 1942 2242
rect 1854 2114 1883 2160
rect 1929 2114 1942 2160
rect 1854 2033 1942 2114
rect 1854 1987 1883 2033
rect 1929 1987 1942 2033
rect 1854 1906 1942 1987
rect 1854 1860 1883 1906
rect 1929 1860 1942 1906
rect 1854 1847 1942 1860
rect 2094 2288 2182 2301
rect 2094 1742 2107 2288
rect 2153 1742 2182 2288
rect 2094 1729 2182 1742
rect 2302 2288 2406 2301
rect 2302 1742 2331 2288
rect 2377 1742 2406 2288
rect 2302 1729 2406 1742
rect 2526 2288 2630 2301
rect 2526 1742 2555 2288
rect 2601 1742 2630 2288
rect 2526 1729 2630 1742
rect 2750 2288 2854 2301
rect 2750 1742 2779 2288
rect 2825 1742 2854 2288
rect 2750 1729 2854 1742
rect 2974 2288 3078 2301
rect 2974 1742 3003 2288
rect 3049 1742 3078 2288
rect 2974 1729 3078 1742
rect 3198 2288 3302 2301
rect 3198 1742 3227 2288
rect 3273 1742 3302 2288
rect 3198 1729 3302 1742
rect 3422 2288 3510 2301
rect 3422 1742 3451 2288
rect 3497 1742 3510 2288
rect 3662 2288 3750 2301
rect 3662 2242 3675 2288
rect 3721 2242 3750 2288
rect 3662 2175 3750 2242
rect 3662 2129 3675 2175
rect 3721 2129 3750 2175
rect 3662 2062 3750 2129
rect 3662 2016 3675 2062
rect 3721 2016 3750 2062
rect 3662 1950 3750 2016
rect 3662 1904 3675 1950
rect 3721 1904 3750 1950
rect 3662 1838 3750 1904
rect 3662 1792 3675 1838
rect 3721 1792 3750 1838
rect 3662 1779 3750 1792
rect 3870 2288 3974 2301
rect 3870 2242 3899 2288
rect 3945 2242 3974 2288
rect 3870 2175 3974 2242
rect 3870 2129 3899 2175
rect 3945 2129 3974 2175
rect 3870 2062 3974 2129
rect 3870 2016 3899 2062
rect 3945 2016 3974 2062
rect 3870 1950 3974 2016
rect 3870 1904 3899 1950
rect 3945 1904 3974 1950
rect 3870 1838 3974 1904
rect 3870 1792 3899 1838
rect 3945 1792 3974 1838
rect 3870 1779 3974 1792
rect 4094 2288 4182 2301
rect 4094 2242 4123 2288
rect 4169 2242 4182 2288
rect 4094 2175 4182 2242
rect 4094 2129 4123 2175
rect 4169 2129 4182 2175
rect 4094 2062 4182 2129
rect 4094 2016 4123 2062
rect 4169 2016 4182 2062
rect 4094 1950 4182 2016
rect 4094 1904 4123 1950
rect 4169 1904 4182 1950
rect 4094 1838 4182 1904
rect 4094 1792 4123 1838
rect 4169 1792 4182 1838
rect 4094 1779 4182 1792
rect 3422 1729 3510 1742
rect 4163 1093 4251 1106
rect 83 1070 171 1083
rect 83 1024 96 1070
rect 142 1024 171 1070
rect 83 914 171 1024
rect 83 868 96 914
rect 142 868 171 914
rect 83 855 171 868
rect 291 1070 395 1083
rect 291 1024 320 1070
rect 366 1024 395 1070
rect 291 914 395 1024
rect 291 868 320 914
rect 366 868 395 914
rect 291 855 395 868
rect 515 1070 619 1083
rect 515 1024 544 1070
rect 590 1024 619 1070
rect 515 914 619 1024
rect 515 868 544 914
rect 590 868 619 914
rect 515 855 619 868
rect 739 1070 843 1083
rect 739 1024 768 1070
rect 814 1024 843 1070
rect 739 914 843 1024
rect 739 868 768 914
rect 814 868 843 914
rect 739 855 843 868
rect 963 1070 1067 1083
rect 963 1024 992 1070
rect 1038 1024 1067 1070
rect 963 914 1067 1024
rect 963 868 992 914
rect 1038 868 1067 914
rect 963 855 1067 868
rect 1187 1070 1275 1083
rect 1187 1024 1216 1070
rect 1262 1024 1275 1070
rect 1187 914 1275 1024
rect 4163 1047 4176 1093
rect 4222 1047 4251 1093
rect 1187 868 1216 914
rect 1262 868 1275 914
rect 1528 967 1616 1004
rect 1528 921 1541 967
rect 1587 921 1616 967
rect 1528 884 1616 921
rect 1736 967 1840 1004
rect 1736 921 1765 967
rect 1811 921 1840 967
rect 1736 884 1840 921
rect 1960 967 2048 1004
rect 1960 921 1989 967
rect 2035 921 2048 967
rect 1960 884 2048 921
rect 2253 967 2341 1004
rect 2253 921 2266 967
rect 2312 921 2341 967
rect 2253 884 2341 921
rect 2461 967 2565 1004
rect 2461 921 2490 967
rect 2536 921 2565 967
rect 2461 884 2565 921
rect 2685 967 2773 1004
rect 2685 921 2714 967
rect 2760 921 2773 967
rect 2685 884 2773 921
rect 2977 967 3065 1004
rect 2977 921 2990 967
rect 3036 921 3065 967
rect 2977 884 3065 921
rect 3185 967 3289 1004
rect 3185 921 3214 967
rect 3260 921 3289 967
rect 3185 884 3289 921
rect 3409 967 3497 1004
rect 3409 921 3438 967
rect 3484 921 3497 967
rect 3409 884 3497 921
rect 3702 967 3790 1004
rect 3702 921 3715 967
rect 3761 921 3790 967
rect 3702 884 3790 921
rect 3910 967 3998 1004
rect 3910 921 3939 967
rect 3985 921 3998 967
rect 3910 884 3998 921
rect 4163 985 4251 1047
rect 4163 939 4176 985
rect 4222 939 4251 985
rect 1187 855 1275 868
rect 4163 877 4251 939
rect 4163 831 4176 877
rect 4222 831 4251 877
rect 4163 818 4251 831
rect 4371 1093 4459 1106
rect 4371 1047 4400 1093
rect 4446 1047 4459 1093
rect 4371 985 4459 1047
rect 4371 939 4400 985
rect 4446 939 4459 985
rect 4371 877 4459 939
rect 4371 831 4400 877
rect 4446 831 4459 877
rect 4371 818 4459 831
<< mvpdiff >>
rect 71 4858 159 4871
rect 71 4202 84 4858
rect 130 4202 159 4858
rect 71 4189 159 4202
rect 279 4858 383 4871
rect 279 4202 308 4858
rect 354 4202 383 4858
rect 279 4189 383 4202
rect 503 4858 591 4871
rect 503 4202 532 4858
rect 578 4202 591 4858
rect 503 4189 591 4202
rect 986 4639 1074 4652
rect 986 4593 999 4639
rect 1045 4593 1074 4639
rect 986 4512 1074 4593
rect 986 4466 999 4512
rect 1045 4466 1074 4512
rect 986 4385 1074 4466
rect 986 4339 999 4385
rect 1045 4339 1074 4385
rect 986 4257 1074 4339
rect 986 4211 999 4257
rect 1045 4211 1074 4257
rect 986 4198 1074 4211
rect 1194 4639 1298 4652
rect 1194 4593 1223 4639
rect 1269 4593 1298 4639
rect 1194 4512 1298 4593
rect 1194 4466 1223 4512
rect 1269 4466 1298 4512
rect 1194 4385 1298 4466
rect 1194 4339 1223 4385
rect 1269 4339 1298 4385
rect 1194 4257 1298 4339
rect 1194 4211 1223 4257
rect 1269 4211 1298 4257
rect 1194 4198 1298 4211
rect 1418 4639 1522 4652
rect 1418 4593 1447 4639
rect 1493 4593 1522 4639
rect 1418 4512 1522 4593
rect 1418 4466 1447 4512
rect 1493 4466 1522 4512
rect 1418 4385 1522 4466
rect 1418 4339 1447 4385
rect 1493 4339 1522 4385
rect 1418 4257 1522 4339
rect 1418 4211 1447 4257
rect 1493 4211 1522 4257
rect 1418 4198 1522 4211
rect 1642 4639 1746 4652
rect 1642 4593 1671 4639
rect 1717 4593 1746 4639
rect 1642 4512 1746 4593
rect 1642 4466 1671 4512
rect 1717 4466 1746 4512
rect 1642 4385 1746 4466
rect 1642 4339 1671 4385
rect 1717 4339 1746 4385
rect 1642 4257 1746 4339
rect 1642 4211 1671 4257
rect 1717 4211 1746 4257
rect 1642 4198 1746 4211
rect 1866 4639 1954 4652
rect 1866 4593 1895 4639
rect 1941 4593 1954 4639
rect 1866 4512 1954 4593
rect 1866 4466 1895 4512
rect 1941 4466 1954 4512
rect 1866 4385 1954 4466
rect 1866 4339 1895 4385
rect 1941 4339 1954 4385
rect 2460 4621 2548 4634
rect 2460 4575 2473 4621
rect 2519 4575 2548 4621
rect 2460 4503 2548 4575
rect 2460 4457 2473 4503
rect 2519 4457 2548 4503
rect 2460 4385 2548 4457
rect 1866 4257 1954 4339
rect 1866 4211 1895 4257
rect 1941 4211 1954 4257
rect 1866 4198 1954 4211
rect 2460 4339 2473 4385
rect 2519 4339 2548 4385
rect 2460 4267 2548 4339
rect 2460 4221 2473 4267
rect 2519 4221 2548 4267
rect 2460 4149 2548 4221
rect 2460 4103 2473 4149
rect 2519 4103 2548 4149
rect 2460 4090 2548 4103
rect 2668 4621 2772 4634
rect 2668 4575 2697 4621
rect 2743 4575 2772 4621
rect 2668 4503 2772 4575
rect 2668 4457 2697 4503
rect 2743 4457 2772 4503
rect 2668 4385 2772 4457
rect 2668 4339 2697 4385
rect 2743 4339 2772 4385
rect 2668 4267 2772 4339
rect 2668 4221 2697 4267
rect 2743 4221 2772 4267
rect 2668 4149 2772 4221
rect 2668 4103 2697 4149
rect 2743 4103 2772 4149
rect 2668 4090 2772 4103
rect 2892 4621 2996 4634
rect 2892 4575 2921 4621
rect 2967 4575 2996 4621
rect 2892 4503 2996 4575
rect 2892 4457 2921 4503
rect 2967 4457 2996 4503
rect 2892 4385 2996 4457
rect 2892 4339 2921 4385
rect 2967 4339 2996 4385
rect 2892 4267 2996 4339
rect 2892 4221 2921 4267
rect 2967 4221 2996 4267
rect 2892 4149 2996 4221
rect 2892 4103 2921 4149
rect 2967 4103 2996 4149
rect 2892 4090 2996 4103
rect 3116 4621 3220 4634
rect 3116 4575 3145 4621
rect 3191 4575 3220 4621
rect 3116 4503 3220 4575
rect 3116 4457 3145 4503
rect 3191 4457 3220 4503
rect 3116 4385 3220 4457
rect 3116 4339 3145 4385
rect 3191 4339 3220 4385
rect 3116 4267 3220 4339
rect 3116 4221 3145 4267
rect 3191 4221 3220 4267
rect 3116 4149 3220 4221
rect 3116 4103 3145 4149
rect 3191 4103 3220 4149
rect 3116 4090 3220 4103
rect 3340 4621 3444 4634
rect 3340 4575 3369 4621
rect 3415 4575 3444 4621
rect 3340 4503 3444 4575
rect 3340 4457 3369 4503
rect 3415 4457 3444 4503
rect 3340 4385 3444 4457
rect 3340 4339 3369 4385
rect 3415 4339 3444 4385
rect 3340 4267 3444 4339
rect 3340 4221 3369 4267
rect 3415 4221 3444 4267
rect 3340 4149 3444 4221
rect 3340 4103 3369 4149
rect 3415 4103 3444 4149
rect 3340 4090 3444 4103
rect 3564 4621 3668 4634
rect 3564 4575 3593 4621
rect 3639 4575 3668 4621
rect 3564 4503 3668 4575
rect 3564 4457 3593 4503
rect 3639 4457 3668 4503
rect 3564 4385 3668 4457
rect 3564 4339 3593 4385
rect 3639 4339 3668 4385
rect 3564 4267 3668 4339
rect 3564 4221 3593 4267
rect 3639 4221 3668 4267
rect 3564 4149 3668 4221
rect 3564 4103 3593 4149
rect 3639 4103 3668 4149
rect 3564 4090 3668 4103
rect 3788 4621 3892 4634
rect 3788 4575 3817 4621
rect 3863 4575 3892 4621
rect 3788 4503 3892 4575
rect 3788 4457 3817 4503
rect 3863 4457 3892 4503
rect 3788 4385 3892 4457
rect 3788 4339 3817 4385
rect 3863 4339 3892 4385
rect 3788 4267 3892 4339
rect 3788 4221 3817 4267
rect 3863 4221 3892 4267
rect 3788 4149 3892 4221
rect 3788 4103 3817 4149
rect 3863 4103 3892 4149
rect 3788 4090 3892 4103
rect 4012 4621 4116 4634
rect 4012 4575 4041 4621
rect 4087 4575 4116 4621
rect 4012 4503 4116 4575
rect 4012 4457 4041 4503
rect 4087 4457 4116 4503
rect 4012 4385 4116 4457
rect 4012 4339 4041 4385
rect 4087 4339 4116 4385
rect 4012 4267 4116 4339
rect 4012 4221 4041 4267
rect 4087 4221 4116 4267
rect 4012 4149 4116 4221
rect 4012 4103 4041 4149
rect 4087 4103 4116 4149
rect 4012 4090 4116 4103
rect 4236 4621 4340 4634
rect 4236 4575 4265 4621
rect 4311 4575 4340 4621
rect 4236 4503 4340 4575
rect 4236 4457 4265 4503
rect 4311 4457 4340 4503
rect 4236 4385 4340 4457
rect 4236 4339 4265 4385
rect 4311 4339 4340 4385
rect 4236 4267 4340 4339
rect 4236 4221 4265 4267
rect 4311 4221 4340 4267
rect 4236 4149 4340 4221
rect 4236 4103 4265 4149
rect 4311 4103 4340 4149
rect 4236 4090 4340 4103
rect 4460 4621 4564 4634
rect 4460 4575 4489 4621
rect 4535 4575 4564 4621
rect 4460 4503 4564 4575
rect 4460 4457 4489 4503
rect 4535 4457 4564 4503
rect 4460 4385 4564 4457
rect 4460 4339 4489 4385
rect 4535 4339 4564 4385
rect 4460 4267 4564 4339
rect 4460 4221 4489 4267
rect 4535 4221 4564 4267
rect 4460 4149 4564 4221
rect 4460 4103 4489 4149
rect 4535 4103 4564 4149
rect 4460 4090 4564 4103
rect 4684 4621 4772 4634
rect 4684 4575 4713 4621
rect 4759 4575 4772 4621
rect 4684 4503 4772 4575
rect 4684 4457 4713 4503
rect 4759 4457 4772 4503
rect 4684 4385 4772 4457
rect 4684 4339 4713 4385
rect 4759 4339 4772 4385
rect 4684 4267 4772 4339
rect 4684 4221 4713 4267
rect 4759 4221 4772 4267
rect 4684 4149 4772 4221
rect 4684 4103 4713 4149
rect 4759 4103 4772 4149
rect 4684 4090 4772 4103
rect 2766 3637 2854 3650
rect 78 3616 166 3629
rect 78 3570 91 3616
rect 137 3570 166 3616
rect 78 3509 166 3570
rect 78 3463 91 3509
rect 137 3463 166 3509
rect 78 3402 166 3463
rect 78 3356 91 3402
rect 137 3356 166 3402
rect 78 3295 166 3356
rect 78 3249 91 3295
rect 137 3249 166 3295
rect 78 3188 166 3249
rect 78 3142 91 3188
rect 137 3142 166 3188
rect 78 3082 166 3142
rect 78 3036 91 3082
rect 137 3036 166 3082
rect 78 2976 166 3036
rect 78 2930 91 2976
rect 137 2930 166 2976
rect 78 2870 166 2930
rect 78 2824 91 2870
rect 137 2824 166 2870
rect 78 2811 166 2824
rect 286 3616 390 3629
rect 286 3570 315 3616
rect 361 3570 390 3616
rect 286 3509 390 3570
rect 286 3463 315 3509
rect 361 3463 390 3509
rect 286 3402 390 3463
rect 286 3356 315 3402
rect 361 3356 390 3402
rect 286 3295 390 3356
rect 286 3249 315 3295
rect 361 3249 390 3295
rect 286 3188 390 3249
rect 286 3142 315 3188
rect 361 3142 390 3188
rect 286 3082 390 3142
rect 286 3036 315 3082
rect 361 3036 390 3082
rect 286 2976 390 3036
rect 286 2930 315 2976
rect 361 2930 390 2976
rect 286 2870 390 2930
rect 286 2824 315 2870
rect 361 2824 390 2870
rect 286 2811 390 2824
rect 510 3616 614 3629
rect 510 3570 539 3616
rect 585 3570 614 3616
rect 510 3509 614 3570
rect 510 3463 539 3509
rect 585 3463 614 3509
rect 510 3402 614 3463
rect 510 3356 539 3402
rect 585 3356 614 3402
rect 510 3295 614 3356
rect 510 3249 539 3295
rect 585 3249 614 3295
rect 510 3188 614 3249
rect 510 3142 539 3188
rect 585 3142 614 3188
rect 510 3082 614 3142
rect 510 3036 539 3082
rect 585 3036 614 3082
rect 510 2976 614 3036
rect 510 2930 539 2976
rect 585 2930 614 2976
rect 510 2870 614 2930
rect 510 2824 539 2870
rect 585 2824 614 2870
rect 510 2811 614 2824
rect 734 3616 838 3629
rect 734 3570 763 3616
rect 809 3570 838 3616
rect 734 3509 838 3570
rect 734 3463 763 3509
rect 809 3463 838 3509
rect 734 3402 838 3463
rect 734 3356 763 3402
rect 809 3356 838 3402
rect 734 3295 838 3356
rect 734 3249 763 3295
rect 809 3249 838 3295
rect 734 3188 838 3249
rect 734 3142 763 3188
rect 809 3142 838 3188
rect 734 3082 838 3142
rect 734 3036 763 3082
rect 809 3036 838 3082
rect 734 2976 838 3036
rect 734 2930 763 2976
rect 809 2930 838 2976
rect 734 2870 838 2930
rect 734 2824 763 2870
rect 809 2824 838 2870
rect 734 2811 838 2824
rect 958 3616 1062 3629
rect 958 3570 987 3616
rect 1033 3570 1062 3616
rect 958 3509 1062 3570
rect 958 3463 987 3509
rect 1033 3463 1062 3509
rect 958 3402 1062 3463
rect 958 3356 987 3402
rect 1033 3356 1062 3402
rect 958 3295 1062 3356
rect 958 3249 987 3295
rect 1033 3249 1062 3295
rect 958 3188 1062 3249
rect 958 3142 987 3188
rect 1033 3142 1062 3188
rect 958 3082 1062 3142
rect 958 3036 987 3082
rect 1033 3036 1062 3082
rect 958 2976 1062 3036
rect 958 2930 987 2976
rect 1033 2930 1062 2976
rect 958 2870 1062 2930
rect 958 2824 987 2870
rect 1033 2824 1062 2870
rect 958 2811 1062 2824
rect 1182 3616 1286 3629
rect 1182 3570 1211 3616
rect 1257 3570 1286 3616
rect 1182 3509 1286 3570
rect 1182 3463 1211 3509
rect 1257 3463 1286 3509
rect 1182 3402 1286 3463
rect 1182 3356 1211 3402
rect 1257 3356 1286 3402
rect 1182 3295 1286 3356
rect 1182 3249 1211 3295
rect 1257 3249 1286 3295
rect 1182 3188 1286 3249
rect 1182 3142 1211 3188
rect 1257 3142 1286 3188
rect 1182 3082 1286 3142
rect 1182 3036 1211 3082
rect 1257 3036 1286 3082
rect 1182 2976 1286 3036
rect 1182 2930 1211 2976
rect 1257 2930 1286 2976
rect 1182 2870 1286 2930
rect 1182 2824 1211 2870
rect 1257 2824 1286 2870
rect 1182 2811 1286 2824
rect 1406 3616 1510 3629
rect 1406 3570 1435 3616
rect 1481 3570 1510 3616
rect 1406 3509 1510 3570
rect 1406 3463 1435 3509
rect 1481 3463 1510 3509
rect 1406 3402 1510 3463
rect 1406 3356 1435 3402
rect 1481 3356 1510 3402
rect 1406 3295 1510 3356
rect 1406 3249 1435 3295
rect 1481 3249 1510 3295
rect 1406 3188 1510 3249
rect 1406 3142 1435 3188
rect 1481 3142 1510 3188
rect 1406 3082 1510 3142
rect 1406 3036 1435 3082
rect 1481 3036 1510 3082
rect 1406 2976 1510 3036
rect 1406 2930 1435 2976
rect 1481 2930 1510 2976
rect 1406 2870 1510 2930
rect 1406 2824 1435 2870
rect 1481 2824 1510 2870
rect 1406 2811 1510 2824
rect 1630 3616 1734 3629
rect 1630 3570 1659 3616
rect 1705 3570 1734 3616
rect 1630 3509 1734 3570
rect 1630 3463 1659 3509
rect 1705 3463 1734 3509
rect 1630 3402 1734 3463
rect 1630 3356 1659 3402
rect 1705 3356 1734 3402
rect 1630 3295 1734 3356
rect 1630 3249 1659 3295
rect 1705 3249 1734 3295
rect 1630 3188 1734 3249
rect 1630 3142 1659 3188
rect 1705 3142 1734 3188
rect 1630 3082 1734 3142
rect 1630 3036 1659 3082
rect 1705 3036 1734 3082
rect 1630 2976 1734 3036
rect 1630 2930 1659 2976
rect 1705 2930 1734 2976
rect 1630 2870 1734 2930
rect 1630 2824 1659 2870
rect 1705 2824 1734 2870
rect 1630 2811 1734 2824
rect 1854 3616 1958 3629
rect 1854 3570 1883 3616
rect 1929 3570 1958 3616
rect 1854 3509 1958 3570
rect 1854 3463 1883 3509
rect 1929 3463 1958 3509
rect 1854 3402 1958 3463
rect 1854 3356 1883 3402
rect 1929 3356 1958 3402
rect 1854 3295 1958 3356
rect 1854 3249 1883 3295
rect 1929 3249 1958 3295
rect 1854 3188 1958 3249
rect 1854 3142 1883 3188
rect 1929 3142 1958 3188
rect 1854 3082 1958 3142
rect 1854 3036 1883 3082
rect 1929 3036 1958 3082
rect 1854 2976 1958 3036
rect 1854 2930 1883 2976
rect 1929 2930 1958 2976
rect 1854 2870 1958 2930
rect 1854 2824 1883 2870
rect 1929 2824 1958 2870
rect 1854 2811 1958 2824
rect 2078 3616 2182 3629
rect 2078 3570 2107 3616
rect 2153 3570 2182 3616
rect 2078 3509 2182 3570
rect 2078 3463 2107 3509
rect 2153 3463 2182 3509
rect 2078 3402 2182 3463
rect 2078 3356 2107 3402
rect 2153 3356 2182 3402
rect 2078 3295 2182 3356
rect 2078 3249 2107 3295
rect 2153 3249 2182 3295
rect 2078 3188 2182 3249
rect 2078 3142 2107 3188
rect 2153 3142 2182 3188
rect 2078 3082 2182 3142
rect 2078 3036 2107 3082
rect 2153 3036 2182 3082
rect 2078 2976 2182 3036
rect 2078 2930 2107 2976
rect 2153 2930 2182 2976
rect 2078 2870 2182 2930
rect 2078 2824 2107 2870
rect 2153 2824 2182 2870
rect 2078 2811 2182 2824
rect 2302 3616 2390 3629
rect 2302 3570 2331 3616
rect 2377 3570 2390 3616
rect 2302 3509 2390 3570
rect 2302 3463 2331 3509
rect 2377 3463 2390 3509
rect 2302 3402 2390 3463
rect 2302 3356 2331 3402
rect 2377 3356 2390 3402
rect 2302 3295 2390 3356
rect 2302 3249 2331 3295
rect 2377 3249 2390 3295
rect 2302 3188 2390 3249
rect 2302 3142 2331 3188
rect 2377 3142 2390 3188
rect 2302 3082 2390 3142
rect 2302 3036 2331 3082
rect 2377 3036 2390 3082
rect 2302 2976 2390 3036
rect 2302 2930 2331 2976
rect 2377 2930 2390 2976
rect 2302 2870 2390 2930
rect 2302 2824 2331 2870
rect 2377 2824 2390 2870
rect 2302 2811 2390 2824
rect 2766 3591 2779 3637
rect 2825 3591 2854 3637
rect 2766 3532 2854 3591
rect 2766 3486 2779 3532
rect 2825 3486 2854 3532
rect 2766 3427 2854 3486
rect 2766 3381 2779 3427
rect 2825 3381 2854 3427
rect 2766 3322 2854 3381
rect 2766 3276 2779 3322
rect 2825 3276 2854 3322
rect 2766 3217 2854 3276
rect 2766 3171 2779 3217
rect 2825 3171 2854 3217
rect 2766 3113 2854 3171
rect 2766 3067 2779 3113
rect 2825 3067 2854 3113
rect 2766 3009 2854 3067
rect 2766 2963 2779 3009
rect 2825 2963 2854 3009
rect 2766 2905 2854 2963
rect 2766 2859 2779 2905
rect 2825 2859 2854 2905
rect 2766 2801 2854 2859
rect 2766 2755 2779 2801
rect 2825 2755 2854 2801
rect 2766 2742 2854 2755
rect 2974 3637 3078 3650
rect 2974 3591 3003 3637
rect 3049 3591 3078 3637
rect 2974 3532 3078 3591
rect 2974 3486 3003 3532
rect 3049 3486 3078 3532
rect 2974 3427 3078 3486
rect 2974 3381 3003 3427
rect 3049 3381 3078 3427
rect 2974 3322 3078 3381
rect 2974 3276 3003 3322
rect 3049 3276 3078 3322
rect 2974 3217 3078 3276
rect 2974 3171 3003 3217
rect 3049 3171 3078 3217
rect 2974 3113 3078 3171
rect 2974 3067 3003 3113
rect 3049 3067 3078 3113
rect 2974 3009 3078 3067
rect 2974 2963 3003 3009
rect 3049 2963 3078 3009
rect 2974 2905 3078 2963
rect 2974 2859 3003 2905
rect 3049 2859 3078 2905
rect 2974 2801 3078 2859
rect 2974 2755 3003 2801
rect 3049 2755 3078 2801
rect 2974 2742 3078 2755
rect 3198 3637 3302 3650
rect 3198 3591 3227 3637
rect 3273 3591 3302 3637
rect 3198 3532 3302 3591
rect 3198 3486 3227 3532
rect 3273 3486 3302 3532
rect 3198 3427 3302 3486
rect 3198 3381 3227 3427
rect 3273 3381 3302 3427
rect 3198 3322 3302 3381
rect 3198 3276 3227 3322
rect 3273 3276 3302 3322
rect 3198 3217 3302 3276
rect 3198 3171 3227 3217
rect 3273 3171 3302 3217
rect 3198 3113 3302 3171
rect 3198 3067 3227 3113
rect 3273 3067 3302 3113
rect 3198 3009 3302 3067
rect 3198 2963 3227 3009
rect 3273 2963 3302 3009
rect 3198 2905 3302 2963
rect 3198 2859 3227 2905
rect 3273 2859 3302 2905
rect 3198 2801 3302 2859
rect 3198 2755 3227 2801
rect 3273 2755 3302 2801
rect 3198 2742 3302 2755
rect 3422 3637 3510 3650
rect 3422 3591 3451 3637
rect 3497 3591 3510 3637
rect 3422 3532 3510 3591
rect 3422 3486 3451 3532
rect 3497 3486 3510 3532
rect 3422 3427 3510 3486
rect 3422 3381 3451 3427
rect 3497 3381 3510 3427
rect 3422 3322 3510 3381
rect 3422 3276 3451 3322
rect 3497 3276 3510 3322
rect 3422 3217 3510 3276
rect 3422 3171 3451 3217
rect 3497 3171 3510 3217
rect 3422 3113 3510 3171
rect 3422 3067 3451 3113
rect 3497 3067 3510 3113
rect 3422 3009 3510 3067
rect 3422 2963 3451 3009
rect 3497 2963 3510 3009
rect 3422 2905 3510 2963
rect 3422 2859 3451 2905
rect 3497 2859 3510 2905
rect 3422 2801 3510 2859
rect 3422 2755 3451 2801
rect 3497 2755 3510 2801
rect 3422 2742 3510 2755
rect 3662 3637 3750 3650
rect 3662 3591 3675 3637
rect 3721 3591 3750 3637
rect 3662 3532 3750 3591
rect 3662 3486 3675 3532
rect 3721 3486 3750 3532
rect 3662 3427 3750 3486
rect 3662 3381 3675 3427
rect 3721 3381 3750 3427
rect 3662 3322 3750 3381
rect 3662 3276 3675 3322
rect 3721 3276 3750 3322
rect 3662 3217 3750 3276
rect 3662 3171 3675 3217
rect 3721 3171 3750 3217
rect 3662 3113 3750 3171
rect 3662 3067 3675 3113
rect 3721 3067 3750 3113
rect 3662 3009 3750 3067
rect 3662 2963 3675 3009
rect 3721 2963 3750 3009
rect 3662 2905 3750 2963
rect 3662 2859 3675 2905
rect 3721 2859 3750 2905
rect 3662 2801 3750 2859
rect 3662 2755 3675 2801
rect 3721 2755 3750 2801
rect 3662 2742 3750 2755
rect 3870 3637 3974 3650
rect 3870 3591 3899 3637
rect 3945 3591 3974 3637
rect 3870 3532 3974 3591
rect 3870 3486 3899 3532
rect 3945 3486 3974 3532
rect 3870 3427 3974 3486
rect 3870 3381 3899 3427
rect 3945 3381 3974 3427
rect 3870 3322 3974 3381
rect 3870 3276 3899 3322
rect 3945 3276 3974 3322
rect 3870 3217 3974 3276
rect 3870 3171 3899 3217
rect 3945 3171 3974 3217
rect 3870 3113 3974 3171
rect 3870 3067 3899 3113
rect 3945 3067 3974 3113
rect 3870 3009 3974 3067
rect 3870 2963 3899 3009
rect 3945 2963 3974 3009
rect 3870 2905 3974 2963
rect 3870 2859 3899 2905
rect 3945 2859 3974 2905
rect 3870 2801 3974 2859
rect 3870 2755 3899 2801
rect 3945 2755 3974 2801
rect 3870 2742 3974 2755
rect 4094 3637 4198 3650
rect 4094 3591 4123 3637
rect 4169 3591 4198 3637
rect 4094 3532 4198 3591
rect 4094 3486 4123 3532
rect 4169 3486 4198 3532
rect 4094 3427 4198 3486
rect 4094 3381 4123 3427
rect 4169 3381 4198 3427
rect 4094 3322 4198 3381
rect 4094 3276 4123 3322
rect 4169 3276 4198 3322
rect 4094 3217 4198 3276
rect 4094 3171 4123 3217
rect 4169 3171 4198 3217
rect 4094 3113 4198 3171
rect 4094 3067 4123 3113
rect 4169 3067 4198 3113
rect 4094 3009 4198 3067
rect 4094 2963 4123 3009
rect 4169 2963 4198 3009
rect 4094 2905 4198 2963
rect 4094 2859 4123 2905
rect 4169 2859 4198 2905
rect 4094 2801 4198 2859
rect 4094 2755 4123 2801
rect 4169 2755 4198 2801
rect 4094 2742 4198 2755
rect 4318 3637 4406 3650
rect 4318 3591 4347 3637
rect 4393 3591 4406 3637
rect 4318 3532 4406 3591
rect 4318 3486 4347 3532
rect 4393 3486 4406 3532
rect 4318 3427 4406 3486
rect 4318 3381 4347 3427
rect 4393 3381 4406 3427
rect 4318 3322 4406 3381
rect 4318 3276 4347 3322
rect 4393 3276 4406 3322
rect 4318 3217 4406 3276
rect 4318 3171 4347 3217
rect 4393 3171 4406 3217
rect 4318 3113 4406 3171
rect 4318 3067 4347 3113
rect 4393 3067 4406 3113
rect 4318 3009 4406 3067
rect 4318 2963 4347 3009
rect 4393 2963 4406 3009
rect 4318 2905 4406 2963
rect 4318 2859 4347 2905
rect 4393 2859 4406 2905
rect 4318 2801 4406 2859
rect 4318 2755 4347 2801
rect 4393 2755 4406 2801
rect 4318 2742 4406 2755
rect 83 559 171 572
rect 83 513 96 559
rect 142 513 171 559
rect 83 432 171 513
rect 83 386 96 432
rect 142 386 171 432
rect 83 305 171 386
rect 83 259 96 305
rect 142 259 171 305
rect 83 177 171 259
rect 83 131 96 177
rect 142 131 171 177
rect 83 118 171 131
rect 291 559 395 572
rect 291 513 320 559
rect 366 513 395 559
rect 291 432 395 513
rect 291 386 320 432
rect 366 386 395 432
rect 291 305 395 386
rect 291 259 320 305
rect 366 259 395 305
rect 291 177 395 259
rect 291 131 320 177
rect 366 131 395 177
rect 291 118 395 131
rect 515 559 619 572
rect 515 513 544 559
rect 590 513 619 559
rect 515 432 619 513
rect 515 386 544 432
rect 590 386 619 432
rect 515 305 619 386
rect 515 259 544 305
rect 590 259 619 305
rect 515 177 619 259
rect 515 131 544 177
rect 590 131 619 177
rect 515 118 619 131
rect 739 559 843 572
rect 739 513 768 559
rect 814 513 843 559
rect 739 432 843 513
rect 739 386 768 432
rect 814 386 843 432
rect 739 305 843 386
rect 739 259 768 305
rect 814 259 843 305
rect 739 177 843 259
rect 739 131 768 177
rect 814 131 843 177
rect 739 118 843 131
rect 963 559 1067 572
rect 963 513 992 559
rect 1038 513 1067 559
rect 963 432 1067 513
rect 963 386 992 432
rect 1038 386 1067 432
rect 963 305 1067 386
rect 963 259 992 305
rect 1038 259 1067 305
rect 963 177 1067 259
rect 963 131 992 177
rect 1038 131 1067 177
rect 963 118 1067 131
rect 1187 559 1275 572
rect 1187 513 1216 559
rect 1262 513 1275 559
rect 3702 561 3790 574
rect 1187 432 1275 513
rect 1187 386 1216 432
rect 1262 386 1275 432
rect 1187 305 1275 386
rect 1187 259 1216 305
rect 1262 259 1275 305
rect 1528 523 1616 536
rect 1528 477 1541 523
rect 1587 477 1616 523
rect 1528 355 1616 477
rect 1528 309 1541 355
rect 1587 309 1616 355
rect 1528 296 1616 309
rect 1736 523 1840 536
rect 1736 477 1765 523
rect 1811 477 1840 523
rect 1736 355 1840 477
rect 1736 309 1765 355
rect 1811 309 1840 355
rect 1736 296 1840 309
rect 1960 523 2048 536
rect 1960 477 1989 523
rect 2035 477 2048 523
rect 1960 355 2048 477
rect 1960 309 1989 355
rect 2035 309 2048 355
rect 1960 296 2048 309
rect 2253 523 2341 536
rect 2253 477 2266 523
rect 2312 477 2341 523
rect 2253 355 2341 477
rect 2253 309 2266 355
rect 2312 309 2341 355
rect 2253 296 2341 309
rect 2461 523 2565 536
rect 2461 477 2490 523
rect 2536 477 2565 523
rect 2461 355 2565 477
rect 2461 309 2490 355
rect 2536 309 2565 355
rect 2461 296 2565 309
rect 2685 523 2773 536
rect 2685 477 2714 523
rect 2760 477 2773 523
rect 2685 355 2773 477
rect 2685 309 2714 355
rect 2760 309 2773 355
rect 2685 296 2773 309
rect 2977 523 3065 536
rect 2977 477 2990 523
rect 3036 477 3065 523
rect 2977 355 3065 477
rect 2977 309 2990 355
rect 3036 309 3065 355
rect 2977 296 3065 309
rect 3185 523 3289 536
rect 3185 477 3214 523
rect 3260 477 3289 523
rect 3185 355 3289 477
rect 3185 309 3214 355
rect 3260 309 3289 355
rect 3185 296 3289 309
rect 3409 523 3497 536
rect 3409 477 3438 523
rect 3484 477 3497 523
rect 3409 355 3497 477
rect 3409 309 3438 355
rect 3484 309 3497 355
rect 3702 515 3715 561
rect 3761 515 3790 561
rect 3702 393 3790 515
rect 3702 347 3715 393
rect 3761 347 3790 393
rect 3702 334 3790 347
rect 3910 561 3998 574
rect 3910 515 3939 561
rect 3985 515 3998 561
rect 3910 393 3998 515
rect 3910 347 3939 393
rect 3985 347 3998 393
rect 3910 334 3998 347
rect 4163 526 4251 539
rect 4163 480 4176 526
rect 4222 480 4251 526
rect 4163 391 4251 480
rect 4163 345 4176 391
rect 4222 345 4251 391
rect 3409 296 3497 309
rect 1187 177 1275 259
rect 4163 256 4251 345
rect 4163 210 4176 256
rect 4222 210 4251 256
rect 4163 197 4251 210
rect 4371 526 4475 539
rect 4371 480 4400 526
rect 4446 480 4475 526
rect 4371 391 4475 480
rect 4371 345 4400 391
rect 4446 345 4475 391
rect 4371 256 4475 345
rect 4371 210 4400 256
rect 4446 210 4475 256
rect 4371 197 4475 210
rect 4595 526 4683 539
rect 4595 480 4624 526
rect 4670 480 4683 526
rect 4595 391 4683 480
rect 4595 345 4624 391
rect 4670 345 4683 391
rect 4595 256 4683 345
rect 4595 210 4624 256
rect 4670 210 4683 256
rect 4595 197 4683 210
rect 1187 131 1216 177
rect 1262 131 1275 177
rect 1187 118 1275 131
<< mvndiffc >>
rect 84 5392 130 5438
rect 84 5236 130 5282
rect 308 5392 354 5438
rect 308 5236 354 5282
rect 532 5392 578 5438
rect 532 5236 578 5282
rect 999 5401 1045 5447
rect 999 5274 1045 5320
rect 999 5147 1045 5193
rect 999 5019 1045 5065
rect 1223 5401 1269 5447
rect 1223 5274 1269 5320
rect 1223 5147 1269 5193
rect 1223 5019 1269 5065
rect 1447 5401 1493 5447
rect 1447 5274 1493 5320
rect 1447 5147 1493 5193
rect 1447 5019 1493 5065
rect 1671 5401 1717 5447
rect 1671 5274 1717 5320
rect 1671 5147 1717 5193
rect 1671 5019 1717 5065
rect 1895 5401 1941 5447
rect 1895 5274 1941 5320
rect 1895 5147 1941 5193
rect 1895 5019 1941 5065
rect 2119 5401 2165 5447
rect 2119 5274 2165 5320
rect 2119 5147 2165 5193
rect 2119 5019 2165 5065
rect 2408 5401 2454 5447
rect 2408 5274 2454 5320
rect 2408 5147 2454 5193
rect 2408 5019 2454 5065
rect 2632 5401 2678 5447
rect 2632 5274 2678 5320
rect 2632 5147 2678 5193
rect 2632 5019 2678 5065
rect 2856 5401 2902 5447
rect 2856 5274 2902 5320
rect 2856 5147 2902 5193
rect 2856 5019 2902 5065
rect 3080 5401 3126 5447
rect 3080 5274 3126 5320
rect 3080 5147 3126 5193
rect 3080 5019 3126 5065
rect 3304 5401 3350 5447
rect 3304 5274 3350 5320
rect 3304 5147 3350 5193
rect 3304 5019 3350 5065
rect 3528 5401 3574 5447
rect 3528 5274 3574 5320
rect 3528 5147 3574 5193
rect 3528 5019 3574 5065
rect 3817 5401 3863 5447
rect 3817 5274 3863 5320
rect 3817 5147 3863 5193
rect 3817 5019 3863 5065
rect 4041 5401 4087 5447
rect 4041 5274 4087 5320
rect 4041 5147 4087 5193
rect 4041 5019 4087 5065
rect 4265 5401 4311 5447
rect 4265 5274 4311 5320
rect 4265 5147 4311 5193
rect 4265 5019 4311 5065
rect 4489 5401 4535 5447
rect 4489 5274 4535 5320
rect 4489 5147 4535 5193
rect 4489 5019 4535 5065
rect 4713 5401 4759 5447
rect 4713 5274 4759 5320
rect 4713 5147 4759 5193
rect 4713 5019 4759 5065
rect 315 2242 361 2288
rect 315 2114 361 2160
rect 315 1987 361 2033
rect 315 1860 361 1906
rect 539 2242 585 2288
rect 539 2114 585 2160
rect 539 1987 585 2033
rect 539 1860 585 1906
rect 763 2242 809 2288
rect 763 2114 809 2160
rect 763 1987 809 2033
rect 763 1860 809 1906
rect 987 2242 1033 2288
rect 987 2114 1033 2160
rect 987 1987 1033 2033
rect 987 1860 1033 1906
rect 1211 2242 1257 2288
rect 1211 2114 1257 2160
rect 1211 1987 1257 2033
rect 1211 1860 1257 1906
rect 1435 2242 1481 2288
rect 1435 2114 1481 2160
rect 1435 1987 1481 2033
rect 1435 1860 1481 1906
rect 1659 2242 1705 2288
rect 1659 2114 1705 2160
rect 1659 1987 1705 2033
rect 1659 1860 1705 1906
rect 1883 2242 1929 2288
rect 1883 2114 1929 2160
rect 1883 1987 1929 2033
rect 1883 1860 1929 1906
rect 2107 1742 2153 2288
rect 2331 1742 2377 2288
rect 2555 1742 2601 2288
rect 2779 1742 2825 2288
rect 3003 1742 3049 2288
rect 3227 1742 3273 2288
rect 3451 1742 3497 2288
rect 3675 2242 3721 2288
rect 3675 2129 3721 2175
rect 3675 2016 3721 2062
rect 3675 1904 3721 1950
rect 3675 1792 3721 1838
rect 3899 2242 3945 2288
rect 3899 2129 3945 2175
rect 3899 2016 3945 2062
rect 3899 1904 3945 1950
rect 3899 1792 3945 1838
rect 4123 2242 4169 2288
rect 4123 2129 4169 2175
rect 4123 2016 4169 2062
rect 4123 1904 4169 1950
rect 4123 1792 4169 1838
rect 96 1024 142 1070
rect 96 868 142 914
rect 320 1024 366 1070
rect 320 868 366 914
rect 544 1024 590 1070
rect 544 868 590 914
rect 768 1024 814 1070
rect 768 868 814 914
rect 992 1024 1038 1070
rect 992 868 1038 914
rect 1216 1024 1262 1070
rect 4176 1047 4222 1093
rect 1216 868 1262 914
rect 1541 921 1587 967
rect 1765 921 1811 967
rect 1989 921 2035 967
rect 2266 921 2312 967
rect 2490 921 2536 967
rect 2714 921 2760 967
rect 2990 921 3036 967
rect 3214 921 3260 967
rect 3438 921 3484 967
rect 3715 921 3761 967
rect 3939 921 3985 967
rect 4176 939 4222 985
rect 4176 831 4222 877
rect 4400 1047 4446 1093
rect 4400 939 4446 985
rect 4400 831 4446 877
<< mvpdiffc >>
rect 84 4202 130 4858
rect 308 4202 354 4858
rect 532 4202 578 4858
rect 999 4593 1045 4639
rect 999 4466 1045 4512
rect 999 4339 1045 4385
rect 999 4211 1045 4257
rect 1223 4593 1269 4639
rect 1223 4466 1269 4512
rect 1223 4339 1269 4385
rect 1223 4211 1269 4257
rect 1447 4593 1493 4639
rect 1447 4466 1493 4512
rect 1447 4339 1493 4385
rect 1447 4211 1493 4257
rect 1671 4593 1717 4639
rect 1671 4466 1717 4512
rect 1671 4339 1717 4385
rect 1671 4211 1717 4257
rect 1895 4593 1941 4639
rect 1895 4466 1941 4512
rect 1895 4339 1941 4385
rect 2473 4575 2519 4621
rect 2473 4457 2519 4503
rect 1895 4211 1941 4257
rect 2473 4339 2519 4385
rect 2473 4221 2519 4267
rect 2473 4103 2519 4149
rect 2697 4575 2743 4621
rect 2697 4457 2743 4503
rect 2697 4339 2743 4385
rect 2697 4221 2743 4267
rect 2697 4103 2743 4149
rect 2921 4575 2967 4621
rect 2921 4457 2967 4503
rect 2921 4339 2967 4385
rect 2921 4221 2967 4267
rect 2921 4103 2967 4149
rect 3145 4575 3191 4621
rect 3145 4457 3191 4503
rect 3145 4339 3191 4385
rect 3145 4221 3191 4267
rect 3145 4103 3191 4149
rect 3369 4575 3415 4621
rect 3369 4457 3415 4503
rect 3369 4339 3415 4385
rect 3369 4221 3415 4267
rect 3369 4103 3415 4149
rect 3593 4575 3639 4621
rect 3593 4457 3639 4503
rect 3593 4339 3639 4385
rect 3593 4221 3639 4267
rect 3593 4103 3639 4149
rect 3817 4575 3863 4621
rect 3817 4457 3863 4503
rect 3817 4339 3863 4385
rect 3817 4221 3863 4267
rect 3817 4103 3863 4149
rect 4041 4575 4087 4621
rect 4041 4457 4087 4503
rect 4041 4339 4087 4385
rect 4041 4221 4087 4267
rect 4041 4103 4087 4149
rect 4265 4575 4311 4621
rect 4265 4457 4311 4503
rect 4265 4339 4311 4385
rect 4265 4221 4311 4267
rect 4265 4103 4311 4149
rect 4489 4575 4535 4621
rect 4489 4457 4535 4503
rect 4489 4339 4535 4385
rect 4489 4221 4535 4267
rect 4489 4103 4535 4149
rect 4713 4575 4759 4621
rect 4713 4457 4759 4503
rect 4713 4339 4759 4385
rect 4713 4221 4759 4267
rect 4713 4103 4759 4149
rect 91 3570 137 3616
rect 91 3463 137 3509
rect 91 3356 137 3402
rect 91 3249 137 3295
rect 91 3142 137 3188
rect 91 3036 137 3082
rect 91 2930 137 2976
rect 91 2824 137 2870
rect 315 3570 361 3616
rect 315 3463 361 3509
rect 315 3356 361 3402
rect 315 3249 361 3295
rect 315 3142 361 3188
rect 315 3036 361 3082
rect 315 2930 361 2976
rect 315 2824 361 2870
rect 539 3570 585 3616
rect 539 3463 585 3509
rect 539 3356 585 3402
rect 539 3249 585 3295
rect 539 3142 585 3188
rect 539 3036 585 3082
rect 539 2930 585 2976
rect 539 2824 585 2870
rect 763 3570 809 3616
rect 763 3463 809 3509
rect 763 3356 809 3402
rect 763 3249 809 3295
rect 763 3142 809 3188
rect 763 3036 809 3082
rect 763 2930 809 2976
rect 763 2824 809 2870
rect 987 3570 1033 3616
rect 987 3463 1033 3509
rect 987 3356 1033 3402
rect 987 3249 1033 3295
rect 987 3142 1033 3188
rect 987 3036 1033 3082
rect 987 2930 1033 2976
rect 987 2824 1033 2870
rect 1211 3570 1257 3616
rect 1211 3463 1257 3509
rect 1211 3356 1257 3402
rect 1211 3249 1257 3295
rect 1211 3142 1257 3188
rect 1211 3036 1257 3082
rect 1211 2930 1257 2976
rect 1211 2824 1257 2870
rect 1435 3570 1481 3616
rect 1435 3463 1481 3509
rect 1435 3356 1481 3402
rect 1435 3249 1481 3295
rect 1435 3142 1481 3188
rect 1435 3036 1481 3082
rect 1435 2930 1481 2976
rect 1435 2824 1481 2870
rect 1659 3570 1705 3616
rect 1659 3463 1705 3509
rect 1659 3356 1705 3402
rect 1659 3249 1705 3295
rect 1659 3142 1705 3188
rect 1659 3036 1705 3082
rect 1659 2930 1705 2976
rect 1659 2824 1705 2870
rect 1883 3570 1929 3616
rect 1883 3463 1929 3509
rect 1883 3356 1929 3402
rect 1883 3249 1929 3295
rect 1883 3142 1929 3188
rect 1883 3036 1929 3082
rect 1883 2930 1929 2976
rect 1883 2824 1929 2870
rect 2107 3570 2153 3616
rect 2107 3463 2153 3509
rect 2107 3356 2153 3402
rect 2107 3249 2153 3295
rect 2107 3142 2153 3188
rect 2107 3036 2153 3082
rect 2107 2930 2153 2976
rect 2107 2824 2153 2870
rect 2331 3570 2377 3616
rect 2331 3463 2377 3509
rect 2331 3356 2377 3402
rect 2331 3249 2377 3295
rect 2331 3142 2377 3188
rect 2331 3036 2377 3082
rect 2331 2930 2377 2976
rect 2331 2824 2377 2870
rect 2779 3591 2825 3637
rect 2779 3486 2825 3532
rect 2779 3381 2825 3427
rect 2779 3276 2825 3322
rect 2779 3171 2825 3217
rect 2779 3067 2825 3113
rect 2779 2963 2825 3009
rect 2779 2859 2825 2905
rect 2779 2755 2825 2801
rect 3003 3591 3049 3637
rect 3003 3486 3049 3532
rect 3003 3381 3049 3427
rect 3003 3276 3049 3322
rect 3003 3171 3049 3217
rect 3003 3067 3049 3113
rect 3003 2963 3049 3009
rect 3003 2859 3049 2905
rect 3003 2755 3049 2801
rect 3227 3591 3273 3637
rect 3227 3486 3273 3532
rect 3227 3381 3273 3427
rect 3227 3276 3273 3322
rect 3227 3171 3273 3217
rect 3227 3067 3273 3113
rect 3227 2963 3273 3009
rect 3227 2859 3273 2905
rect 3227 2755 3273 2801
rect 3451 3591 3497 3637
rect 3451 3486 3497 3532
rect 3451 3381 3497 3427
rect 3451 3276 3497 3322
rect 3451 3171 3497 3217
rect 3451 3067 3497 3113
rect 3451 2963 3497 3009
rect 3451 2859 3497 2905
rect 3451 2755 3497 2801
rect 3675 3591 3721 3637
rect 3675 3486 3721 3532
rect 3675 3381 3721 3427
rect 3675 3276 3721 3322
rect 3675 3171 3721 3217
rect 3675 3067 3721 3113
rect 3675 2963 3721 3009
rect 3675 2859 3721 2905
rect 3675 2755 3721 2801
rect 3899 3591 3945 3637
rect 3899 3486 3945 3532
rect 3899 3381 3945 3427
rect 3899 3276 3945 3322
rect 3899 3171 3945 3217
rect 3899 3067 3945 3113
rect 3899 2963 3945 3009
rect 3899 2859 3945 2905
rect 3899 2755 3945 2801
rect 4123 3591 4169 3637
rect 4123 3486 4169 3532
rect 4123 3381 4169 3427
rect 4123 3276 4169 3322
rect 4123 3171 4169 3217
rect 4123 3067 4169 3113
rect 4123 2963 4169 3009
rect 4123 2859 4169 2905
rect 4123 2755 4169 2801
rect 4347 3591 4393 3637
rect 4347 3486 4393 3532
rect 4347 3381 4393 3427
rect 4347 3276 4393 3322
rect 4347 3171 4393 3217
rect 4347 3067 4393 3113
rect 4347 2963 4393 3009
rect 4347 2859 4393 2905
rect 4347 2755 4393 2801
rect 96 513 142 559
rect 96 386 142 432
rect 96 259 142 305
rect 96 131 142 177
rect 320 513 366 559
rect 320 386 366 432
rect 320 259 366 305
rect 320 131 366 177
rect 544 513 590 559
rect 544 386 590 432
rect 544 259 590 305
rect 544 131 590 177
rect 768 513 814 559
rect 768 386 814 432
rect 768 259 814 305
rect 768 131 814 177
rect 992 513 1038 559
rect 992 386 1038 432
rect 992 259 1038 305
rect 992 131 1038 177
rect 1216 513 1262 559
rect 1216 386 1262 432
rect 1216 259 1262 305
rect 1541 477 1587 523
rect 1541 309 1587 355
rect 1765 477 1811 523
rect 1765 309 1811 355
rect 1989 477 2035 523
rect 1989 309 2035 355
rect 2266 477 2312 523
rect 2266 309 2312 355
rect 2490 477 2536 523
rect 2490 309 2536 355
rect 2714 477 2760 523
rect 2714 309 2760 355
rect 2990 477 3036 523
rect 2990 309 3036 355
rect 3214 477 3260 523
rect 3214 309 3260 355
rect 3438 477 3484 523
rect 3438 309 3484 355
rect 3715 515 3761 561
rect 3715 347 3761 393
rect 3939 515 3985 561
rect 3939 347 3985 393
rect 4176 480 4222 526
rect 4176 345 4222 391
rect 4176 210 4222 256
rect 4400 480 4446 526
rect 4400 345 4446 391
rect 4400 210 4446 256
rect 4624 480 4670 526
rect 4624 345 4670 391
rect 4624 210 4670 256
rect 1216 131 1262 177
<< psubdiff >>
rect -352 5539 -268 5558
rect -352 5211 -333 5539
rect -287 5211 -268 5539
rect -352 5192 -268 5211
rect -389 2191 86 2250
rect -389 2145 -333 2191
rect -287 2145 -175 2191
rect -129 2145 -17 2191
rect 29 2145 86 2191
rect -389 2027 86 2145
rect -389 1981 -333 2027
rect -287 1981 -175 2027
rect -129 1981 -17 2027
rect 29 1981 86 2027
rect -389 1922 86 1981
rect 4560 2191 5035 2250
rect 4560 2145 4616 2191
rect 4662 2145 4774 2191
rect 4820 2145 4932 2191
rect 4978 2145 5035 2191
rect 4560 2027 5035 2145
rect 4560 1981 4616 2027
rect 4662 1981 4774 2027
rect 4820 1981 4932 2027
rect 4978 1981 5035 2027
rect 4560 1922 5035 1981
rect -468 1088 -151 1148
rect -468 1042 -412 1088
rect -366 1042 -254 1088
rect -208 1042 -151 1088
rect -468 983 -151 1042
rect 4718 1088 5035 1148
rect 4718 1042 4774 1088
rect 4820 1042 4932 1088
rect 4978 1042 5035 1088
rect 4718 983 5035 1042
<< nsubdiff >>
rect -387 3759 -232 3816
rect -387 3713 -333 3759
rect -287 3713 -232 3759
rect 4720 3759 5033 3816
rect -387 3596 -232 3713
rect 4720 3713 4774 3759
rect 4820 3713 4932 3759
rect 4978 3713 5033 3759
rect -387 3550 -333 3596
rect -287 3550 -232 3596
rect -387 3433 -232 3550
rect -387 3387 -333 3433
rect -287 3387 -232 3433
rect -387 3269 -232 3387
rect -387 3223 -333 3269
rect -287 3223 -232 3269
rect -387 3106 -232 3223
rect -387 3060 -333 3106
rect -287 3060 -232 3106
rect -387 2943 -232 3060
rect -387 2897 -333 2943
rect -287 2897 -232 2943
rect -387 2840 -232 2897
rect 4720 3596 5033 3713
rect 4720 3550 4774 3596
rect 4820 3550 4932 3596
rect 4978 3550 5033 3596
rect 4720 3433 5033 3550
rect 4720 3387 4774 3433
rect 4820 3387 4932 3433
rect 4978 3387 5033 3433
rect 4720 3269 5033 3387
rect 4720 3223 4774 3269
rect 4820 3223 4932 3269
rect 4978 3223 5033 3269
rect 4720 3106 5033 3223
rect 4720 3060 4774 3106
rect 4820 3060 4932 3106
rect 4978 3060 5033 3106
rect 4720 2943 5033 3060
rect 4720 2897 4774 2943
rect 4820 2897 4932 2943
rect 4978 2897 5033 2943
rect 4720 2840 5033 2897
rect -387 388 -232 445
rect -387 342 -333 388
rect -287 342 -232 388
rect -387 285 -232 342
<< psubdiffcont >>
rect -333 5211 -287 5539
rect -333 2145 -287 2191
rect -175 2145 -129 2191
rect -17 2145 29 2191
rect -333 1981 -287 2027
rect -175 1981 -129 2027
rect -17 1981 29 2027
rect 4616 2145 4662 2191
rect 4774 2145 4820 2191
rect 4932 2145 4978 2191
rect 4616 1981 4662 2027
rect 4774 1981 4820 2027
rect 4932 1981 4978 2027
rect -412 1042 -366 1088
rect -254 1042 -208 1088
rect 4774 1042 4820 1088
rect 4932 1042 4978 1088
<< nsubdiffcont >>
rect -333 3713 -287 3759
rect 4774 3713 4820 3759
rect 4932 3713 4978 3759
rect -333 3550 -287 3596
rect -333 3387 -287 3433
rect -333 3223 -287 3269
rect -333 3060 -287 3106
rect -333 2897 -287 2943
rect 4774 3550 4820 3596
rect 4932 3550 4978 3596
rect 4774 3387 4820 3433
rect 4932 3387 4978 3433
rect 4774 3223 4820 3269
rect 4932 3223 4978 3269
rect 4774 3060 4820 3106
rect 4932 3060 4978 3106
rect 4774 2897 4820 2943
rect 4932 2897 4978 2943
rect -333 342 -287 388
<< polysilicon >>
rect 159 5451 279 5523
rect 383 5451 503 5523
rect 1074 5460 1194 5532
rect 1298 5460 1418 5532
rect 1522 5460 1642 5532
rect 1746 5460 1866 5532
rect 1970 5460 2090 5532
rect 2270 5520 3499 5580
rect 159 4871 279 5223
rect 383 4871 503 5223
rect 1074 4934 1194 5006
rect 1298 4934 1418 5006
rect 1522 4934 1642 5006
rect 1746 4934 1866 5006
rect 1970 4934 2090 5006
rect 661 4888 2090 4934
rect 661 4842 735 4888
rect 781 4873 2090 4888
rect 781 4842 854 4873
rect 661 4796 854 4842
rect 1074 4652 1194 4873
rect 1298 4652 1418 4873
rect 1522 4652 1642 4873
rect 2270 4772 2328 5520
rect 2483 5460 2603 5520
rect 2707 5460 2827 5520
rect 2931 5460 3051 5520
rect 3155 5460 3275 5520
rect 3379 5460 3499 5520
rect 3892 5460 4012 5532
rect 4116 5460 4236 5532
rect 4340 5460 4460 5532
rect 4564 5460 4684 5532
rect 2483 4932 2603 5006
rect 2707 4932 2827 5006
rect 2931 4932 3051 5006
rect 3155 4932 3275 5006
rect 3379 4932 3499 5006
rect 3892 4834 4012 5006
rect 1746 4712 2328 4772
rect 1746 4652 1866 4712
rect 2014 4683 2328 4712
rect 2548 4788 4012 4834
rect 2548 4742 2623 4788
rect 2669 4742 2781 4788
rect 2827 4742 2939 4788
rect 2985 4742 3097 4788
rect 3143 4742 3255 4788
rect 3301 4759 4012 4788
rect 4116 4759 4236 5006
rect 4340 4759 4460 5006
rect 4564 4759 4684 5006
rect 3301 4742 4684 4759
rect 2548 4698 4684 4742
rect 2548 4696 3376 4698
rect 2014 4607 2206 4683
rect 2548 4634 2668 4696
rect 2772 4634 2892 4696
rect 2996 4634 3116 4696
rect 3220 4634 3340 4696
rect 3444 4634 3564 4698
rect 3668 4634 3788 4698
rect 3892 4634 4012 4698
rect 4116 4634 4236 4698
rect 4340 4634 4460 4698
rect 4564 4634 4684 4698
rect 2014 4561 2087 4607
rect 2133 4561 2206 4607
rect 2014 4443 2206 4561
rect 2014 4397 2087 4443
rect 2133 4397 2206 4443
rect 2014 4351 2206 4397
rect 159 4118 279 4189
rect 383 4118 503 4189
rect 1074 4125 1194 4198
rect 1298 4125 1418 4198
rect 1522 4125 1642 4198
rect 1746 4125 1866 4198
rect 159 4072 503 4118
rect 159 4026 298 4072
rect 344 4026 503 4072
rect 159 3980 503 4026
rect 2548 4016 2668 4090
rect 2772 4016 2892 4090
rect 2996 4016 3116 4090
rect 3220 4016 3340 4090
rect 3444 4016 3564 4090
rect 3668 4016 3788 4090
rect 3892 4016 4012 4090
rect 4116 4016 4236 4090
rect 4340 4016 4460 4090
rect 4564 4016 4684 4090
rect 2796 3788 2974 3807
rect 2796 3742 2815 3788
rect 2955 3742 2974 3788
rect 2796 3723 2974 3742
rect 166 3629 286 3703
rect 390 3629 510 3703
rect 614 3629 734 3703
rect 838 3629 958 3703
rect 1062 3629 1182 3703
rect 1286 3629 1406 3703
rect 1510 3629 1630 3703
rect 1734 3629 1854 3703
rect 1958 3629 2078 3703
rect 2182 3629 2302 3703
rect 2854 3650 2974 3723
rect 3078 3650 3198 3723
rect 3302 3650 3422 3723
rect 3750 3650 3870 3723
rect 3974 3650 4094 3723
rect 4198 3650 4318 3723
rect 166 2749 286 2811
rect 390 2749 510 2811
rect 614 2749 734 2811
rect 838 2749 958 2811
rect 1062 2749 1182 2811
rect 1286 2749 1406 2811
rect 1510 2749 1630 2811
rect 1734 2749 1854 2811
rect 1958 2749 2078 2811
rect 2182 2749 2302 2811
rect 166 2709 2302 2749
rect 166 2690 2477 2709
rect 166 2688 2318 2690
rect 390 2301 510 2688
rect 614 2301 734 2688
rect 838 2301 958 2688
rect 1062 2301 1182 2688
rect 1286 2301 1406 2688
rect 1510 2301 1630 2688
rect 1734 2644 2318 2688
rect 2458 2644 2477 2690
rect 1734 2625 2477 2644
rect 1734 2301 1854 2625
rect 2182 2433 2302 2452
rect 2182 2387 2217 2433
rect 2263 2387 2302 2433
rect 2854 2422 2974 2742
rect 2182 2301 2302 2387
rect 2406 2301 2526 2374
rect 2630 2361 2974 2422
rect 2630 2301 2750 2361
rect 2854 2301 2974 2361
rect 3078 2301 3198 2742
rect 3302 2449 3422 2742
rect 3750 2671 3870 2742
rect 3974 2671 4094 2742
rect 4198 2671 4318 2742
rect 3750 2651 4318 2671
rect 3568 2632 4318 2651
rect 3568 2586 3587 2632
rect 3633 2611 4318 2632
rect 3633 2586 3870 2611
rect 3568 2568 3870 2586
rect 3568 2567 3652 2568
rect 3302 2403 3332 2449
rect 3378 2403 3422 2449
rect 3302 2301 3422 2403
rect 3750 2301 3870 2568
rect 3974 2301 4094 2611
rect 390 1774 510 1847
rect 614 1774 734 1847
rect 838 1774 958 1847
rect 1062 1774 1182 1847
rect 1286 1774 1406 1847
rect 1510 1774 1630 1847
rect 1734 1774 1854 1847
rect 3750 1735 3870 1779
rect 3974 1735 4094 1779
rect 2182 1656 2302 1729
rect 2406 1577 2526 1729
rect 2630 1656 2750 1729
rect 2854 1656 2974 1729
rect 2406 1576 2527 1577
rect 3078 1576 3198 1729
rect 3302 1656 3422 1729
rect 3751 1706 3870 1735
rect 3975 1706 4094 1735
rect 2406 1531 3198 1576
rect 2406 1516 2786 1531
rect 2713 1485 2786 1516
rect 2832 1516 3198 1531
rect 2832 1485 2905 1516
rect 2713 1440 2905 1485
rect 246 1336 439 1381
rect 246 1290 320 1336
rect 366 1290 439 1336
rect 246 1259 439 1290
rect 887 1336 1080 1381
rect 887 1290 961 1336
rect 1007 1290 1080 1336
rect 887 1259 1080 1290
rect 171 1198 1186 1259
rect 171 1083 291 1198
rect 395 1083 515 1198
rect 619 1083 739 1198
rect 843 1083 963 1198
rect 1067 1127 1186 1198
rect 4251 1150 4370 1177
rect 1067 1083 1187 1127
rect 4251 1106 4371 1150
rect 1616 1004 1736 1048
rect 1840 1004 1960 1048
rect 2341 1004 2461 1048
rect 2565 1004 2685 1048
rect 3065 1004 3185 1048
rect 3289 1004 3409 1048
rect 3790 1004 3910 1048
rect 171 572 291 855
rect 395 572 515 855
rect 619 572 739 855
rect 843 572 963 855
rect 1067 811 1187 855
rect 1067 616 1186 811
rect 1616 756 1736 884
rect 1305 737 1736 756
rect 1305 691 1324 737
rect 1370 691 1736 737
rect 1305 672 1736 691
rect 1067 572 1187 616
rect 1616 536 1736 672
rect 1840 796 1960 884
rect 2341 840 2461 884
rect 2341 815 2460 840
rect 1840 750 1859 796
rect 1905 750 1960 796
rect 1840 536 1960 750
rect 2029 796 2460 815
rect 2029 750 2048 796
rect 2094 750 2460 796
rect 2029 731 2460 750
rect 2340 683 2460 731
rect 2341 580 2460 683
rect 2565 735 2685 884
rect 3065 754 3185 884
rect 2565 689 2584 735
rect 2630 689 2685 735
rect 2341 536 2461 580
rect 2565 536 2685 689
rect 2796 735 3185 754
rect 2796 689 2815 735
rect 2861 689 3185 735
rect 2796 670 3185 689
rect 3065 536 3185 670
rect 3289 735 3409 884
rect 3790 754 3910 884
rect 3289 689 3308 735
rect 3354 689 3409 735
rect 3289 536 3409 689
rect 3495 735 3910 754
rect 3495 689 3514 735
rect 3560 689 3910 735
rect 4251 713 4371 818
rect 3495 670 3910 689
rect 3790 574 3910 670
rect 4188 694 4595 713
rect 4188 648 4207 694
rect 4253 648 4595 694
rect 4188 629 4595 648
rect 4251 539 4371 629
rect 4475 539 4595 629
rect 1616 252 1736 296
rect 1840 252 1960 296
rect 2341 252 2461 296
rect 2565 252 2685 296
rect 3065 252 3185 296
rect 3289 252 3409 296
rect 3790 273 3910 334
rect 4251 153 4371 197
rect 4475 153 4595 197
rect 4251 123 4370 153
rect 4475 123 4594 153
rect 171 74 291 118
rect 395 74 515 118
rect 619 74 739 118
rect 843 74 963 118
rect 1067 74 1187 118
rect 171 44 290 74
rect 395 44 514 74
rect 619 44 738 74
rect 843 44 962 74
rect 1067 44 1186 74
<< polycontact >>
rect 735 4842 781 4888
rect 2623 4742 2669 4788
rect 2781 4742 2827 4788
rect 2939 4742 2985 4788
rect 3097 4742 3143 4788
rect 3255 4742 3301 4788
rect 2087 4561 2133 4607
rect 2087 4397 2133 4443
rect 298 4026 344 4072
rect 2815 3742 2955 3788
rect 2318 2644 2458 2690
rect 2217 2387 2263 2433
rect 3587 2586 3633 2632
rect 3332 2403 3378 2449
rect 2786 1485 2832 1531
rect 320 1290 366 1336
rect 961 1290 1007 1336
rect 1324 691 1370 737
rect 1859 750 1905 796
rect 2048 750 2094 796
rect 2584 689 2630 735
rect 2815 689 2861 735
rect 3308 689 3354 735
rect 3514 689 3560 735
rect 4207 648 4253 694
<< metal1 >>
rect -356 5539 -264 5550
rect -356 5510 -333 5539
rect -287 5510 -264 5539
rect -356 5458 -336 5510
rect -284 5458 -264 5510
rect -356 5324 -333 5458
rect -287 5324 -264 5458
rect -356 5272 -336 5324
rect -284 5272 -264 5324
rect -356 5242 -333 5272
rect -344 5211 -333 5242
rect -287 5242 -264 5272
rect 13 5491 105 5531
rect 13 5439 33 5491
rect 85 5451 105 5491
rect 509 5491 601 5531
rect 85 5439 130 5451
rect 13 5438 130 5439
rect 13 5392 84 5438
rect 13 5305 130 5392
rect 13 5253 33 5305
rect 85 5282 130 5305
rect -287 5211 -276 5242
rect 13 5236 84 5253
rect 13 5223 130 5236
rect 308 5438 354 5451
rect 308 5282 354 5392
rect -344 5200 -276 5211
rect 308 5120 354 5236
rect 509 5439 529 5491
rect 581 5439 601 5491
rect 1190 5530 3574 5597
rect 999 5447 1045 5460
rect 1190 5451 1305 5530
rect 509 5438 601 5439
rect 509 5392 532 5438
rect 578 5392 601 5438
rect 509 5305 601 5392
rect 509 5253 529 5305
rect 581 5253 601 5305
rect 509 5236 532 5253
rect 578 5236 601 5253
rect 509 5223 601 5236
rect 973 5405 999 5445
rect 1189 5447 1305 5451
rect 973 5353 993 5405
rect 1045 5353 1065 5445
rect 973 5320 1065 5353
rect 973 5274 999 5320
rect 1045 5274 1065 5320
rect 973 5219 1065 5274
rect 1189 5401 1223 5447
rect 1269 5401 1305 5447
rect 1447 5447 1493 5460
rect 1189 5320 1305 5401
rect 1189 5274 1223 5320
rect 1269 5274 1305 5320
rect 1189 5268 1305 5274
rect 1412 5405 1447 5445
rect 1635 5447 1751 5530
rect 1412 5353 1432 5405
rect 1493 5401 1504 5445
rect 1484 5353 1504 5401
rect 1412 5320 1504 5353
rect 1412 5274 1447 5320
rect 1493 5274 1504 5320
rect 973 5167 993 5219
rect 973 5147 999 5167
rect 1045 5147 1065 5219
rect 973 5137 1065 5147
rect 1223 5193 1269 5268
rect 308 5045 763 5120
rect 84 4858 130 4871
rect 61 4369 84 4409
rect 308 4858 354 5045
rect 691 4924 763 5045
rect 999 5065 1045 5137
rect 999 5006 1045 5019
rect 1223 5065 1269 5147
rect 1412 5219 1504 5274
rect 1412 5167 1432 5219
rect 1484 5193 1504 5219
rect 1412 5147 1447 5167
rect 1493 5147 1504 5193
rect 1412 5137 1504 5147
rect 1635 5401 1671 5447
rect 1717 5401 1751 5447
rect 1895 5447 1941 5460
rect 1635 5320 1751 5401
rect 1635 5274 1671 5320
rect 1717 5274 1751 5320
rect 1635 5193 1751 5274
rect 1635 5147 1671 5193
rect 1717 5147 1751 5193
rect 1635 5145 1751 5147
rect 1878 5401 1895 5445
rect 2083 5447 2199 5530
rect 1941 5405 1970 5445
rect 1878 5353 1898 5401
rect 1950 5353 1970 5405
rect 1878 5320 1970 5353
rect 1878 5274 1895 5320
rect 1941 5274 1970 5320
rect 1878 5219 1970 5274
rect 1878 5193 1898 5219
rect 1878 5147 1895 5193
rect 1950 5167 1970 5219
rect 1941 5147 1970 5167
rect 1223 5006 1269 5019
rect 1447 5065 1493 5137
rect 1447 5006 1493 5019
rect 1671 5065 1717 5145
rect 1878 5137 1970 5147
rect 2083 5401 2119 5447
rect 2165 5401 2199 5447
rect 2083 5320 2199 5401
rect 2083 5274 2119 5320
rect 2165 5274 2199 5320
rect 2083 5193 2199 5274
rect 2083 5147 2119 5193
rect 2165 5147 2199 5193
rect 2083 5145 2199 5147
rect 2408 5447 2454 5460
rect 2408 5320 2454 5401
rect 2408 5193 2454 5274
rect 1671 5006 1717 5019
rect 1895 5065 1941 5137
rect 1895 5006 1941 5019
rect 2119 5065 2165 5145
rect 2119 5006 2165 5019
rect 2408 5065 2454 5147
rect 691 4888 815 4924
rect 130 4369 153 4409
rect 61 4317 81 4369
rect 133 4317 153 4369
rect 61 4202 84 4317
rect 130 4202 153 4317
rect 61 4183 153 4202
rect 532 4858 578 4871
rect 308 4189 354 4202
rect 509 4369 532 4409
rect 691 4842 735 4888
rect 781 4842 815 4888
rect 2408 4843 2454 5019
rect 2632 5447 2678 5530
rect 2632 5320 2678 5401
rect 2632 5193 2678 5274
rect 2632 5065 2678 5147
rect 2632 5006 2678 5019
rect 2856 5447 2902 5460
rect 2856 5320 2902 5401
rect 2856 5193 2902 5274
rect 2856 5065 2902 5147
rect 2856 4843 2902 5019
rect 3080 5447 3126 5530
rect 3080 5320 3126 5401
rect 3080 5193 3126 5274
rect 3080 5065 3126 5147
rect 3080 5006 3126 5019
rect 3304 5447 3350 5460
rect 3304 5320 3350 5401
rect 3304 5193 3350 5274
rect 3304 5065 3350 5147
rect 3304 4843 3350 5019
rect 3528 5447 3574 5530
rect 4007 5530 4569 5580
rect 3817 5447 3863 5460
rect 3528 5320 3574 5401
rect 3528 5193 3574 5274
rect 3528 5065 3574 5147
rect 3795 5405 3817 5445
rect 4007 5447 4123 5530
rect 3863 5405 3887 5445
rect 3795 5353 3815 5405
rect 3867 5353 3887 5405
rect 3795 5320 3887 5353
rect 3795 5274 3817 5320
rect 3863 5274 3887 5320
rect 3795 5219 3887 5274
rect 3795 5167 3815 5219
rect 3867 5167 3887 5219
rect 3795 5147 3817 5167
rect 3863 5147 3887 5167
rect 3795 5137 3887 5147
rect 4007 5401 4041 5447
rect 4087 5401 4123 5447
rect 4265 5447 4311 5460
rect 4007 5320 4123 5401
rect 4007 5274 4041 5320
rect 4087 5274 4123 5320
rect 4007 5193 4123 5274
rect 4007 5147 4041 5193
rect 4087 5147 4123 5193
rect 3528 5006 3574 5019
rect 3817 5065 3863 5137
rect 3817 5006 3863 5019
rect 4007 5065 4123 5147
rect 4241 5405 4265 5445
rect 4453 5447 4569 5530
rect 4311 5405 4333 5445
rect 4241 5353 4261 5405
rect 4313 5353 4333 5405
rect 4241 5320 4333 5353
rect 4241 5274 4265 5320
rect 4311 5274 4333 5320
rect 4241 5219 4333 5274
rect 4241 5167 4261 5219
rect 4313 5167 4333 5219
rect 4241 5147 4265 5167
rect 4311 5147 4333 5167
rect 4241 5137 4333 5147
rect 4453 5401 4489 5447
rect 4535 5401 4569 5447
rect 4713 5447 4759 5460
rect 4453 5320 4569 5401
rect 4453 5274 4489 5320
rect 4535 5274 4569 5320
rect 4453 5193 4569 5274
rect 4453 5147 4489 5193
rect 4535 5147 4569 5193
rect 4007 5019 4041 5065
rect 4087 5019 4123 5065
rect 691 4805 815 4842
rect 1187 4811 3350 4843
rect 1187 4759 2313 4811
rect 2365 4759 2493 4811
rect 2545 4788 3350 4811
rect 2545 4759 2623 4788
rect 1187 4742 2623 4759
rect 2669 4742 2781 4788
rect 2827 4742 2939 4788
rect 2985 4742 3097 4788
rect 3143 4742 3255 4788
rect 3301 4742 3350 4788
rect 1187 4723 3350 4742
rect 999 4639 1045 4652
rect 999 4512 1045 4593
rect 1187 4639 1303 4723
rect 1187 4593 1223 4639
rect 1269 4593 1303 4639
rect 1187 4512 1303 4593
rect 1187 4481 1223 4512
rect 999 4452 1045 4466
rect 1269 4481 1303 4512
rect 1447 4639 1493 4652
rect 1447 4512 1493 4593
rect 1635 4639 1751 4723
rect 2589 4705 3350 4723
rect 1635 4593 1671 4639
rect 1717 4593 1751 4639
rect 1635 4585 1751 4593
rect 1895 4639 1941 4652
rect 2054 4617 2166 4643
rect 975 4412 1067 4452
rect 578 4369 601 4409
rect 509 4317 529 4369
rect 581 4317 601 4369
rect 509 4202 532 4317
rect 578 4202 601 4317
rect 61 4131 81 4183
rect 133 4131 153 4183
rect 61 4101 153 4131
rect 509 4183 601 4202
rect 509 4131 529 4183
rect 581 4131 601 4183
rect 975 4360 995 4412
rect 1047 4360 1067 4412
rect 975 4339 999 4360
rect 1045 4339 1067 4360
rect 975 4257 1067 4339
rect 975 4226 999 4257
rect 1045 4226 1067 4257
rect 975 4174 995 4226
rect 1047 4174 1067 4226
rect 1223 4385 1269 4466
rect 1447 4409 1493 4466
rect 1671 4512 1717 4585
rect 1223 4257 1269 4339
rect 1223 4198 1269 4211
rect 1412 4385 1504 4409
rect 1412 4369 1447 4385
rect 1412 4317 1432 4369
rect 1493 4339 1504 4385
rect 1484 4317 1504 4339
rect 1412 4257 1504 4317
rect 1412 4211 1447 4257
rect 1493 4211 1504 4257
rect 975 4144 1067 4174
rect 1412 4183 1504 4211
rect 1671 4385 1717 4466
rect 1895 4512 1941 4593
rect 1895 4409 1941 4466
rect 2053 4607 2166 4617
rect 2053 4576 2087 4607
rect 2053 4524 2073 4576
rect 2133 4561 2166 4607
rect 2125 4524 2166 4561
rect 2053 4443 2166 4524
rect 1671 4257 1717 4339
rect 1671 4198 1717 4211
rect 1858 4385 1950 4409
rect 1858 4369 1895 4385
rect 1858 4317 1878 4369
rect 1941 4339 1950 4385
rect 1930 4317 1950 4339
rect 1858 4257 1950 4317
rect 2053 4397 2087 4443
rect 2133 4397 2166 4443
rect 2473 4621 2519 4634
rect 2473 4503 2519 4575
rect 2473 4434 2519 4457
rect 2697 4621 2743 4634
rect 2697 4503 2743 4575
rect 2053 4390 2166 4397
rect 2053 4338 2073 4390
rect 2125 4360 2166 4390
rect 2464 4394 2556 4434
rect 2464 4385 2484 4394
rect 2125 4338 2145 4360
rect 2053 4298 2145 4338
rect 2464 4339 2473 4385
rect 2536 4342 2556 4394
rect 2697 4385 2743 4457
rect 2921 4621 2967 4634
rect 2921 4503 2967 4575
rect 2921 4434 2967 4457
rect 3145 4621 3191 4634
rect 3145 4503 3191 4575
rect 2519 4339 2556 4342
rect 1858 4211 1895 4257
rect 1941 4211 1950 4257
rect 263 4072 378 4108
rect 509 4101 601 4131
rect 1412 4131 1432 4183
rect 1484 4131 1504 4183
rect 1412 4101 1504 4131
rect 1858 4183 1950 4211
rect 1858 4131 1878 4183
rect 1930 4131 1950 4183
rect 1858 4101 1950 4131
rect 2464 4267 2556 4339
rect 2464 4221 2473 4267
rect 2519 4221 2556 4267
rect 2464 4208 2556 4221
rect 2464 4156 2484 4208
rect 2536 4156 2556 4208
rect 2464 4149 2556 4156
rect 2464 4126 2473 4149
rect 2519 4126 2556 4149
rect 2665 4339 2697 4358
rect 2901 4394 2993 4434
rect 2743 4339 2781 4358
rect 2665 4267 2781 4339
rect 2665 4221 2697 4267
rect 2743 4221 2781 4267
rect 2665 4149 2781 4221
rect 2473 4090 2519 4103
rect 2665 4103 2697 4149
rect 2743 4103 2781 4149
rect 2901 4339 2921 4394
rect 2973 4342 2993 4394
rect 3145 4385 3191 4457
rect 3369 4621 3415 4634
rect 3369 4503 3415 4575
rect 3369 4434 3415 4457
rect 3593 4621 3639 4634
rect 3593 4503 3639 4575
rect 2967 4339 2993 4342
rect 2901 4267 2993 4339
rect 2901 4221 2921 4267
rect 2967 4221 2993 4267
rect 2901 4208 2993 4221
rect 2901 4156 2921 4208
rect 2973 4156 2993 4208
rect 2901 4149 2993 4156
rect 2901 4126 2921 4149
rect 263 4026 298 4072
rect 344 4026 378 4072
rect 263 4000 378 4026
rect 843 4000 1152 4022
rect -356 3962 -264 3992
rect -356 3910 -336 3962
rect -284 3910 -264 3962
rect 263 3948 881 4000
rect 933 3948 1061 4000
rect 1113 3948 1152 4000
rect 263 3925 1152 3948
rect 2665 4018 2781 4103
rect 2967 4126 2993 4149
rect 3111 4339 3145 4379
rect 3343 4394 3435 4434
rect 3191 4339 3227 4379
rect 3111 4267 3227 4339
rect 3111 4221 3145 4267
rect 3191 4221 3227 4267
rect 3111 4149 3227 4221
rect 2921 4090 2967 4103
rect 3111 4103 3145 4149
rect 3191 4103 3227 4149
rect 3343 4342 3363 4394
rect 3343 4339 3369 4342
rect 3415 4339 3435 4394
rect 3593 4385 3639 4457
rect 3817 4621 3863 4634
rect 3817 4503 3863 4575
rect 3817 4434 3863 4457
rect 4007 4621 4123 5019
rect 4265 5065 4311 5137
rect 4265 5006 4311 5019
rect 4453 5065 4569 5147
rect 4693 5353 4713 5445
rect 4759 5405 4785 5445
rect 4765 5353 4785 5405
rect 4693 5320 4785 5353
rect 4693 5274 4713 5320
rect 4759 5274 4785 5320
rect 4693 5219 4785 5274
rect 4693 5147 4713 5219
rect 4765 5167 4785 5219
rect 4759 5147 4785 5167
rect 4693 5137 4785 5147
rect 4453 5019 4489 5065
rect 4535 5019 4569 5065
rect 4007 4575 4041 4621
rect 4087 4575 4123 4621
rect 4007 4503 4123 4575
rect 4007 4457 4041 4503
rect 4087 4457 4123 4503
rect 3343 4267 3435 4339
rect 3343 4221 3369 4267
rect 3415 4221 3435 4267
rect 3343 4208 3435 4221
rect 3343 4156 3363 4208
rect 3415 4156 3435 4208
rect 3343 4149 3435 4156
rect 3343 4126 3369 4149
rect 3111 4018 3227 4103
rect 3415 4126 3435 4149
rect 3559 4339 3593 4379
rect 3797 4394 3889 4434
rect 3639 4339 3675 4379
rect 3559 4267 3675 4339
rect 3559 4221 3593 4267
rect 3639 4221 3675 4267
rect 3559 4149 3675 4221
rect 3369 4090 3415 4103
rect 3559 4103 3593 4149
rect 3639 4103 3675 4149
rect 3797 4339 3817 4394
rect 3869 4342 3889 4394
rect 3863 4339 3889 4342
rect 3797 4267 3889 4339
rect 3797 4221 3817 4267
rect 3863 4221 3889 4267
rect 3797 4208 3889 4221
rect 3797 4156 3817 4208
rect 3869 4156 3889 4208
rect 3797 4149 3889 4156
rect 3797 4126 3817 4149
rect 3559 4018 3675 4103
rect 3863 4126 3889 4149
rect 4007 4385 4123 4457
rect 4265 4621 4311 4634
rect 4265 4503 4311 4575
rect 4265 4434 4311 4457
rect 4453 4621 4569 5019
rect 4713 5065 4759 5137
rect 4713 5006 4759 5019
rect 4453 4575 4489 4621
rect 4535 4575 4569 4621
rect 4453 4503 4569 4575
rect 4453 4457 4489 4503
rect 4535 4457 4569 4503
rect 4007 4339 4041 4385
rect 4087 4339 4123 4385
rect 4007 4267 4123 4339
rect 4007 4221 4041 4267
rect 4087 4221 4123 4267
rect 4007 4149 4123 4221
rect 3817 4090 3863 4103
rect 4007 4103 4041 4149
rect 4087 4103 4123 4149
rect 4243 4394 4335 4434
rect 4243 4342 4263 4394
rect 4315 4342 4335 4394
rect 4243 4339 4265 4342
rect 4311 4339 4335 4342
rect 4243 4267 4335 4339
rect 4243 4221 4265 4267
rect 4311 4221 4335 4267
rect 4243 4208 4335 4221
rect 4243 4156 4263 4208
rect 4315 4156 4335 4208
rect 4243 4149 4335 4156
rect 4243 4126 4265 4149
rect 4007 4018 4123 4103
rect 4311 4126 4335 4149
rect 4453 4385 4569 4457
rect 4713 4621 4759 4634
rect 4713 4503 4759 4575
rect 4713 4434 4759 4457
rect 4453 4339 4489 4385
rect 4535 4339 4569 4385
rect 4453 4267 4569 4339
rect 4453 4221 4489 4267
rect 4535 4221 4569 4267
rect 4453 4149 4569 4221
rect 4265 4090 4311 4103
rect 4453 4103 4489 4149
rect 4535 4103 4569 4149
rect 4691 4394 4783 4434
rect 4691 4342 4711 4394
rect 4763 4342 4783 4394
rect 4691 4339 4713 4342
rect 4759 4339 4783 4342
rect 4691 4267 4783 4339
rect 4691 4221 4713 4267
rect 4759 4221 4783 4267
rect 4691 4208 4783 4221
rect 4691 4156 4711 4208
rect 4763 4156 4783 4208
rect 4691 4149 4783 4156
rect 4691 4126 4713 4149
rect 4453 4018 4569 4103
rect 4759 4126 4783 4149
rect 4713 4090 4759 4103
rect -356 3796 -264 3910
rect 2665 3898 4569 4018
rect 4909 3851 5001 3881
rect -367 3776 -252 3796
rect -367 3724 -336 3776
rect -284 3724 -252 3776
rect -367 3713 -333 3724
rect -287 3713 -252 3724
rect -367 3596 -252 3713
rect 54 3721 2412 3841
rect 2778 3796 3086 3818
rect 4909 3799 4929 3851
rect 4981 3799 5001 3851
rect 4909 3796 5001 3799
rect 2778 3788 2816 3796
rect 2868 3788 2996 3796
rect 2778 3742 2815 3788
rect 2955 3744 2996 3788
rect 3048 3744 3086 3796
rect 2955 3742 3086 3744
rect 2778 3722 3086 3742
rect 4739 3759 5013 3796
rect 54 3636 170 3721
rect -367 3550 -333 3596
rect -287 3550 -252 3596
rect -367 3433 -252 3550
rect -367 3387 -333 3433
rect -287 3387 -252 3433
rect -367 3384 -252 3387
rect -367 3332 -336 3384
rect -284 3332 -252 3384
rect -367 3269 -252 3332
rect 13 3616 170 3636
rect 13 3596 91 3616
rect 13 3544 33 3596
rect 85 3570 91 3596
rect 137 3570 170 3616
rect 85 3544 170 3570
rect 13 3509 170 3544
rect 13 3463 91 3509
rect 137 3463 170 3509
rect 13 3410 170 3463
rect 13 3358 33 3410
rect 85 3402 170 3410
rect 85 3358 91 3402
rect 13 3356 91 3358
rect 137 3356 170 3402
rect 13 3328 170 3356
rect 54 3325 170 3328
rect 315 3616 361 3629
rect 315 3509 361 3570
rect 315 3402 361 3463
rect 505 3616 620 3721
rect 505 3570 539 3616
rect 585 3570 620 3616
rect 505 3509 620 3570
rect 505 3463 539 3509
rect 585 3463 620 3509
rect 505 3402 620 3463
rect 505 3365 539 3402
rect -367 3223 -333 3269
rect -287 3223 -252 3269
rect -367 3198 -252 3223
rect -367 3146 -336 3198
rect -284 3146 -252 3198
rect -367 3106 -252 3146
rect -367 3060 -333 3106
rect -287 3060 -252 3106
rect -367 2943 -252 3060
rect -367 2897 -333 2943
rect -287 2897 -252 2943
rect -367 2860 -252 2897
rect 91 3295 137 3325
rect 91 3188 137 3249
rect 91 3082 137 3142
rect 91 2976 137 3036
rect 91 2870 137 2930
rect 315 3295 361 3356
rect 315 3188 361 3249
rect 315 3082 361 3142
rect 315 2976 361 3036
rect 315 2870 361 2930
rect 91 2811 137 2824
rect 281 2824 315 2866
rect 585 3365 620 3402
rect 763 3616 809 3629
rect 763 3509 809 3570
rect 763 3402 809 3463
rect 539 3295 585 3356
rect 539 3188 585 3249
rect 539 3082 585 3142
rect 539 2976 585 3036
rect 539 2870 585 2930
rect 361 2824 396 2866
rect 281 2633 396 2824
rect 953 3616 1068 3721
rect 953 3570 987 3616
rect 1033 3570 1068 3616
rect 953 3509 1068 3570
rect 953 3463 987 3509
rect 1033 3463 1068 3509
rect 953 3402 1068 3463
rect 953 3365 987 3402
rect 763 3295 809 3356
rect 763 3188 809 3249
rect 763 3082 809 3142
rect 763 2976 809 3036
rect 763 2870 809 2930
rect 539 2811 585 2824
rect 729 2824 763 2866
rect 1033 3365 1068 3402
rect 1211 3616 1257 3629
rect 1211 3509 1257 3570
rect 1211 3402 1257 3463
rect 987 3295 1033 3356
rect 987 3188 1033 3249
rect 987 3082 1033 3142
rect 987 2976 1033 3036
rect 987 2870 1033 2930
rect 809 2824 844 2866
rect 729 2633 844 2824
rect 1400 3616 1516 3721
rect 1400 3596 1435 3616
rect 1481 3596 1516 3616
rect 1400 3544 1432 3596
rect 1484 3544 1516 3596
rect 1400 3509 1516 3544
rect 1400 3463 1435 3509
rect 1481 3463 1516 3509
rect 1400 3410 1516 3463
rect 1400 3365 1432 3410
rect 1211 3295 1257 3356
rect 1412 3358 1432 3365
rect 1484 3365 1516 3410
rect 1659 3616 1705 3629
rect 1659 3509 1705 3570
rect 1659 3402 1705 3463
rect 1484 3358 1504 3365
rect 1412 3356 1435 3358
rect 1481 3356 1504 3358
rect 1412 3328 1504 3356
rect 1848 3616 1964 3721
rect 1848 3570 1883 3616
rect 1929 3570 1964 3616
rect 1848 3509 1964 3570
rect 1848 3463 1883 3509
rect 1929 3463 1964 3509
rect 1848 3402 1964 3463
rect 1848 3365 1883 3402
rect 1211 3188 1257 3249
rect 1211 3082 1257 3142
rect 1211 2976 1257 3036
rect 1211 2870 1257 2930
rect 987 2811 1033 2824
rect 1177 2824 1211 2866
rect 1435 3295 1481 3328
rect 1435 3188 1481 3249
rect 1435 3082 1481 3142
rect 1435 2976 1481 3036
rect 1435 2870 1481 2930
rect 1257 2824 1292 2866
rect 1177 2633 1292 2824
rect 1659 3295 1705 3356
rect 1659 3188 1705 3249
rect 1659 3082 1705 3142
rect 1659 2976 1705 3036
rect 1659 2870 1705 2930
rect 1435 2811 1481 2824
rect 1624 2824 1659 2866
rect 1929 3365 1964 3402
rect 2107 3616 2153 3629
rect 2107 3509 2153 3570
rect 2296 3616 2412 3721
rect 4739 3713 4774 3759
rect 4820 3713 4932 3759
rect 4978 3713 5013 3759
rect 4739 3665 5013 3713
rect 2296 3570 2331 3616
rect 2377 3570 2412 3616
rect 2779 3637 2825 3650
rect 2779 3575 2825 3591
rect 3003 3637 3049 3650
rect 2296 3553 2412 3570
rect 2296 3501 2317 3553
rect 2369 3509 2412 3553
rect 2296 3472 2331 3501
rect 2107 3402 2153 3463
rect 1883 3295 1929 3356
rect 2107 3336 2153 3356
rect 2297 3463 2331 3472
rect 2377 3472 2412 3509
rect 2776 3535 2868 3575
rect 2776 3532 2796 3535
rect 2776 3486 2779 3532
rect 2776 3483 2796 3486
rect 2848 3483 2868 3535
rect 2377 3463 2389 3472
rect 2297 3402 2389 3463
rect 2297 3367 2331 3402
rect 1883 3188 1929 3249
rect 1883 3082 1929 3142
rect 1883 2976 1929 3036
rect 1883 2870 1929 2930
rect 1705 2824 1740 2866
rect 1624 2719 1740 2824
rect 1883 2811 1929 2824
rect 2072 3295 2188 3336
rect 2072 3249 2107 3295
rect 2153 3249 2188 3295
rect 2297 3315 2317 3367
rect 2377 3356 2389 3402
rect 2369 3315 2389 3356
rect 2297 3295 2389 3315
rect 2297 3285 2331 3295
rect 2072 3188 2188 3249
rect 2072 3142 2107 3188
rect 2153 3142 2188 3188
rect 2072 3082 2188 3142
rect 2072 3036 2107 3082
rect 2153 3036 2188 3082
rect 2072 2976 2188 3036
rect 2072 2930 2107 2976
rect 2153 2930 2188 2976
rect 2072 2870 2188 2930
rect 2072 2824 2107 2870
rect 2153 2824 2188 2870
rect 2072 2719 2188 2824
rect 2377 3285 2389 3295
rect 2776 3427 2868 3483
rect 2776 3381 2779 3427
rect 2825 3381 2868 3427
rect 2776 3349 2868 3381
rect 2776 3322 2796 3349
rect 2776 3276 2779 3322
rect 2848 3297 2868 3349
rect 2825 3276 2868 3297
rect 2776 3267 2868 3276
rect 3003 3532 3049 3591
rect 3227 3637 3273 3650
rect 3227 3575 3273 3591
rect 3451 3637 3497 3650
rect 3003 3427 3049 3486
rect 3003 3322 3049 3381
rect 2331 3188 2377 3249
rect 2331 3082 2377 3142
rect 2331 2976 2377 3036
rect 2331 2870 2377 2930
rect 2331 2811 2377 2824
rect 2779 3217 2825 3267
rect 2779 3113 2825 3171
rect 2779 3009 2825 3067
rect 2779 2905 2825 2963
rect 2779 2801 2825 2859
rect 3003 3217 3049 3276
rect 3206 3535 3298 3575
rect 3206 3483 3226 3535
rect 3278 3483 3298 3535
rect 3206 3427 3298 3483
rect 3206 3381 3227 3427
rect 3273 3381 3298 3427
rect 3206 3349 3298 3381
rect 3206 3297 3226 3349
rect 3278 3297 3298 3349
rect 3206 3276 3227 3297
rect 3273 3276 3298 3297
rect 3206 3267 3298 3276
rect 3451 3532 3497 3591
rect 3675 3637 3721 3650
rect 3675 3575 3721 3591
rect 3899 3637 3945 3650
rect 3451 3427 3497 3486
rect 3451 3322 3497 3381
rect 3003 3113 3049 3171
rect 3003 3009 3049 3067
rect 3003 2905 3049 2963
rect 3003 2803 3049 2859
rect 3227 3217 3273 3267
rect 3227 3113 3273 3171
rect 3227 3009 3273 3067
rect 3227 2905 3273 2963
rect 2779 2742 2825 2755
rect 2968 2801 3084 2803
rect 2968 2755 3003 2801
rect 3049 2755 3084 2801
rect 1624 2633 2188 2719
rect 281 2599 2188 2633
rect 2294 2718 2592 2741
rect 2294 2690 2330 2718
rect 2382 2690 2592 2718
rect 2294 2644 2318 2690
rect 2458 2644 2592 2690
rect 2968 2672 3084 2755
rect 3227 2801 3273 2859
rect 3227 2742 3273 2755
rect 3451 3217 3497 3276
rect 3650 3535 3742 3575
rect 3650 3483 3670 3535
rect 3722 3483 3742 3535
rect 3650 3427 3742 3483
rect 3650 3381 3675 3427
rect 3721 3381 3742 3427
rect 3650 3349 3742 3381
rect 3650 3297 3670 3349
rect 3722 3297 3742 3349
rect 3650 3276 3675 3297
rect 3721 3276 3742 3297
rect 3650 3267 3742 3276
rect 3899 3532 3945 3591
rect 4123 3637 4169 3650
rect 4123 3575 4169 3591
rect 4347 3637 4393 3650
rect 3899 3427 3945 3486
rect 3899 3322 3945 3381
rect 3451 3113 3497 3171
rect 3451 3009 3497 3067
rect 3451 2905 3497 2963
rect 3451 2801 3497 2859
rect 3451 2672 3497 2755
rect 3675 3217 3721 3267
rect 3675 3113 3721 3171
rect 3675 3009 3721 3067
rect 3899 3217 3945 3276
rect 4100 3535 4192 3575
rect 4100 3483 4120 3535
rect 4172 3483 4192 3535
rect 4100 3427 4192 3483
rect 4100 3381 4123 3427
rect 4169 3381 4192 3427
rect 4100 3349 4192 3381
rect 4100 3297 4120 3349
rect 4172 3297 4192 3349
rect 4100 3276 4123 3297
rect 4169 3276 4192 3297
rect 4100 3267 4192 3276
rect 4347 3532 4393 3591
rect 4347 3427 4393 3486
rect 4347 3322 4393 3381
rect 3899 3113 3945 3171
rect 3899 3009 3945 3067
rect 4123 3217 4169 3267
rect 4123 3113 4169 3171
rect 4123 3009 4169 3067
rect 4347 3217 4393 3276
rect 4347 3113 4393 3171
rect 4347 3009 4393 3067
rect 4739 3613 4929 3665
rect 4981 3613 5013 3665
rect 4739 3596 5013 3613
rect 4739 3550 4774 3596
rect 4820 3550 4932 3596
rect 4978 3550 5013 3596
rect 4739 3433 5013 3550
rect 4739 3387 4774 3433
rect 4820 3387 4932 3433
rect 4978 3387 5013 3433
rect 4739 3384 5013 3387
rect 4739 3332 4929 3384
rect 4981 3332 5013 3384
rect 4739 3269 5013 3332
rect 4739 3223 4774 3269
rect 4820 3223 4932 3269
rect 4978 3223 5013 3269
rect 4739 3198 5013 3223
rect 4739 3146 4929 3198
rect 4981 3146 5013 3198
rect 4739 3106 5013 3146
rect 4739 3060 4774 3106
rect 4820 3060 4932 3106
rect 4978 3060 5013 3106
rect 3675 2905 3721 2963
rect 3675 2801 3721 2859
rect 3876 2923 3968 2963
rect 3876 2871 3896 2923
rect 3948 2871 3968 2923
rect 3876 2859 3899 2871
rect 3945 2859 3968 2871
rect 3876 2842 3968 2859
rect 4123 2905 4169 2963
rect 3675 2742 3721 2755
rect 3864 2801 3980 2842
rect 3864 2755 3899 2801
rect 3945 2755 3980 2801
rect 3864 2737 3980 2755
rect 4123 2801 4169 2859
rect 4123 2742 4169 2755
rect 4326 2923 4418 2963
rect 4326 2871 4346 2923
rect 4398 2871 4418 2923
rect 4326 2859 4347 2871
rect 4393 2859 4418 2871
rect 4739 2943 5013 3060
rect 4739 2897 4774 2943
rect 4820 2897 4932 2943
rect 4978 2897 5013 2943
rect 4739 2860 5013 2897
rect 4326 2801 4418 2859
rect 4326 2755 4347 2801
rect 4393 2755 4418 2801
rect 3864 2685 3896 2737
rect 3948 2685 3980 2737
rect 2968 2671 3085 2672
rect 3451 2671 3533 2672
rect 281 2513 1740 2599
rect 2294 2583 2592 2644
rect 2744 2632 3655 2671
rect 2744 2586 3587 2632
rect 3633 2586 3655 2632
rect 281 2288 396 2513
rect 281 2242 315 2288
rect 361 2242 396 2288
rect -356 2240 -264 2242
rect -380 2212 77 2240
rect -380 2160 -336 2212
rect -284 2191 77 2212
rect -284 2160 -175 2191
rect -380 2145 -333 2160
rect -287 2145 -175 2160
rect -129 2145 -17 2191
rect 29 2145 77 2191
rect 281 2187 396 2242
rect 539 2288 585 2301
rect -380 2027 77 2145
rect -380 2026 -333 2027
rect -287 2026 -175 2027
rect -380 1974 -336 2026
rect -284 1981 -175 2026
rect -129 1981 -17 2027
rect 29 1981 77 2027
rect -284 1974 77 1981
rect -380 1931 77 1974
rect 315 2160 361 2187
rect 539 2186 585 2242
rect 729 2288 844 2513
rect 729 2242 763 2288
rect 809 2242 844 2288
rect 729 2187 844 2242
rect 987 2288 1033 2301
rect 315 2033 361 2114
rect 315 1906 361 1987
rect 315 1847 361 1860
rect 505 2160 620 2186
rect 505 2114 539 2160
rect 585 2114 620 2160
rect 505 2033 620 2114
rect 505 1987 539 2033
rect 585 1987 620 2033
rect 505 1906 620 1987
rect 505 1860 539 1906
rect 585 1860 620 1906
rect 505 1762 620 1860
rect 763 2160 809 2187
rect 987 2186 1033 2242
rect 1177 2288 1292 2513
rect 1177 2242 1211 2288
rect 1257 2242 1292 2288
rect 1435 2288 1481 2301
rect 1177 2187 1292 2242
rect 1414 2242 1435 2251
rect 1624 2288 1740 2513
rect 2744 2552 3655 2586
rect 2181 2449 2489 2471
rect 2181 2433 2219 2449
rect 2181 2387 2217 2433
rect 2271 2397 2399 2449
rect 2451 2397 2489 2449
rect 2263 2387 2489 2397
rect 2181 2375 2489 2387
rect 1481 2242 1506 2251
rect 1414 2211 1506 2242
rect 763 2033 809 2114
rect 763 1906 809 1987
rect 763 1847 809 1860
rect 953 2160 1068 2186
rect 953 2114 987 2160
rect 1033 2114 1068 2160
rect 953 2033 1068 2114
rect 953 1987 987 2033
rect 1033 1987 1068 2033
rect 953 1906 1068 1987
rect 953 1860 987 1906
rect 1033 1860 1068 1906
rect 953 1762 1068 1860
rect 1211 2160 1257 2187
rect 1414 2186 1434 2211
rect 1211 2033 1257 2114
rect 1211 1906 1257 1987
rect 1211 1847 1257 1860
rect 1400 2159 1434 2186
rect 1486 2186 1506 2211
rect 1624 2242 1659 2288
rect 1705 2242 1740 2288
rect 1624 2187 1740 2242
rect 1883 2288 1929 2301
rect 2107 2288 2153 2301
rect 1486 2159 1516 2186
rect 1400 2114 1435 2159
rect 1481 2114 1516 2159
rect 1400 2033 1516 2114
rect 1400 2025 1435 2033
rect 1481 2025 1516 2033
rect 1400 1973 1434 2025
rect 1486 1973 1516 2025
rect 1400 1906 1516 1973
rect 1400 1860 1435 1906
rect 1481 1860 1516 1906
rect 1400 1762 1516 1860
rect 1659 2160 1705 2187
rect 1659 2033 1705 2114
rect 1883 2160 1929 2242
rect 1883 2035 1929 2114
rect 2082 2211 2107 2251
rect 2331 2288 2377 2301
rect 2153 2211 2174 2251
rect 2082 2159 2102 2211
rect 2154 2159 2174 2211
rect 1659 1906 1705 1987
rect 1659 1847 1705 1860
rect 1870 2033 1942 2035
rect 1870 1987 1883 2033
rect 1929 1987 1942 2033
rect 1870 1906 1942 1987
rect 2082 2025 2107 2159
rect 2153 2025 2174 2159
rect 2082 1973 2102 2025
rect 2154 1973 2174 2025
rect 2082 1943 2107 1973
rect 1870 1860 1883 1906
rect 1929 1860 1942 1906
rect 1870 1762 1942 1860
rect 505 1688 1942 1762
rect 2153 1943 2174 1973
rect 2107 1729 2153 1742
rect 2331 1729 2377 1742
rect 2555 2288 2601 2301
rect 2744 2288 2860 2552
rect 3083 2449 3391 2471
rect 3083 2397 3121 2449
rect 3173 2397 3301 2449
rect 3378 2403 3391 2449
rect 3353 2397 3391 2403
rect 3083 2375 3391 2397
rect 2744 1765 2779 2288
rect 2555 1729 2601 1742
rect 2825 1765 2860 2288
rect 3003 2288 3049 2301
rect 2779 1729 2825 1742
rect 3003 1729 3049 1742
rect 3227 2288 3273 2301
rect 3451 2288 3497 2301
rect 3430 2211 3451 2251
rect 3675 2288 3721 2301
rect 3497 2211 3522 2251
rect 3430 2159 3450 2211
rect 3502 2159 3522 2211
rect 3430 2025 3451 2159
rect 3497 2025 3522 2159
rect 3430 1973 3450 2025
rect 3502 1973 3522 2025
rect 3430 1943 3451 1973
rect 3227 1729 3273 1742
rect 3497 1943 3522 1973
rect 3652 2242 3675 2251
rect 3864 2288 3980 2685
rect 4326 2737 4418 2755
rect 4326 2685 4346 2737
rect 4398 2685 4418 2737
rect 4326 2655 4418 2685
rect 3721 2242 3744 2251
rect 3652 2211 3744 2242
rect 3652 2159 3672 2211
rect 3724 2159 3744 2211
rect 3864 2242 3899 2288
rect 3945 2242 3980 2288
rect 4123 2288 4169 2301
rect 3864 2175 3980 2242
rect 3864 2162 3899 2175
rect 3652 2129 3675 2159
rect 3721 2129 3744 2159
rect 3652 2062 3744 2129
rect 3652 2025 3675 2062
rect 3721 2025 3744 2062
rect 3652 1973 3672 2025
rect 3724 1973 3744 2025
rect 3652 1950 3744 1973
rect 3652 1943 3675 1950
rect 3721 1943 3744 1950
rect 3945 2162 3980 2175
rect 4098 2242 4123 2251
rect 4169 2242 4190 2251
rect 4098 2211 4190 2242
rect 4909 2240 5001 2242
rect 3899 2062 3945 2129
rect 3899 1950 3945 2016
rect 3675 1838 3721 1904
rect 3675 1779 3721 1792
rect 4098 2159 4118 2211
rect 4170 2159 4190 2211
rect 4098 2129 4123 2159
rect 4169 2129 4190 2159
rect 4098 2062 4190 2129
rect 4098 2025 4123 2062
rect 4169 2025 4190 2062
rect 4098 1973 4118 2025
rect 4170 1973 4190 2025
rect 4098 1950 4190 1973
rect 4098 1943 4123 1950
rect 3899 1838 3945 1904
rect 3899 1779 3945 1792
rect 4169 1943 4190 1950
rect 4569 2212 5026 2240
rect 4569 2191 4929 2212
rect 4569 2145 4616 2191
rect 4662 2145 4774 2191
rect 4820 2160 4929 2191
rect 4981 2160 5026 2212
rect 4820 2145 4932 2160
rect 4978 2145 5026 2160
rect 4569 2027 5026 2145
rect 4569 1981 4616 2027
rect 4662 1981 4774 2027
rect 4820 2026 4932 2027
rect 4978 2026 5026 2027
rect 4820 1981 4929 2026
rect 4569 1974 4929 1981
rect 4981 1974 5026 2026
rect 4569 1931 5026 1974
rect 4123 1838 4169 1904
rect 4123 1779 4169 1792
rect 4574 1786 4955 1826
rect 3451 1729 3497 1742
rect 4574 1734 4611 1786
rect 4663 1734 4823 1786
rect 4875 1734 4955 1786
rect 74 1568 414 1608
rect 864 1604 4470 1608
rect 74 1516 112 1568
rect 164 1516 324 1568
rect 376 1516 414 1568
rect 74 1390 414 1516
rect 860 1584 4470 1604
rect 860 1532 890 1584
rect 942 1532 1076 1584
rect 1128 1532 4191 1584
rect 4243 1532 4377 1584
rect 4429 1532 4470 1584
rect 860 1531 4470 1532
rect 860 1512 2786 1531
rect 864 1511 2786 1512
rect 2752 1485 2786 1511
rect 2832 1511 4470 1531
rect 4574 1568 4955 1734
rect 4574 1516 4611 1568
rect 4663 1516 4823 1568
rect 4875 1516 4955 1568
rect 2832 1485 2867 1511
rect 2752 1471 2867 1485
rect 4574 1391 4955 1516
rect 4574 1390 4956 1391
rect -374 1350 5025 1390
rect -374 1298 112 1350
rect 164 1336 324 1350
rect 376 1336 1983 1350
rect 164 1298 320 1336
rect 376 1298 961 1336
rect -374 1290 320 1298
rect 366 1290 961 1298
rect 1007 1298 1983 1336
rect 2035 1298 2193 1350
rect 2245 1298 2404 1350
rect 2456 1298 2615 1350
rect 2667 1298 2826 1350
rect 2878 1298 3037 1350
rect 3089 1298 3248 1350
rect 3300 1298 3459 1350
rect 3511 1298 3670 1350
rect 3722 1298 3881 1350
rect 3933 1298 4091 1350
rect 4143 1298 4611 1350
rect 4663 1298 4823 1350
rect 4875 1298 5025 1350
rect 1007 1290 5025 1298
rect -374 1253 5025 1290
rect -460 1108 -160 1139
rect -460 1088 -336 1108
rect -460 1042 -412 1088
rect -366 1056 -336 1088
rect -284 1088 -160 1108
rect -284 1056 -254 1088
rect -366 1042 -254 1056
rect -208 1042 -160 1088
rect -460 992 -160 1042
rect 72 1121 164 1161
rect 72 1069 92 1121
rect 144 1069 164 1121
rect 492 1121 584 1161
rect 72 1024 96 1069
rect 142 1024 164 1069
rect -356 991 -262 992
rect -356 922 -264 991
rect -356 870 -336 922
rect -284 870 -264 922
rect -356 830 -264 870
rect 72 935 164 1024
rect 72 883 92 935
rect 144 883 164 935
rect 72 868 96 883
rect 142 868 164 883
rect 72 842 164 868
rect 320 1070 366 1083
rect 320 914 366 1024
rect 320 762 366 868
rect 492 1069 512 1121
rect 564 1083 584 1121
rect 964 1121 1056 1161
rect 564 1070 590 1083
rect 492 1024 544 1069
rect 492 935 590 1024
rect 492 883 512 935
rect 564 914 590 935
rect 492 868 544 883
rect 492 855 590 868
rect 768 1070 814 1083
rect 768 914 814 1024
rect 492 842 584 855
rect 768 762 814 868
rect 964 1069 984 1121
rect 1036 1070 1056 1121
rect 964 1024 992 1069
rect 1038 1024 1056 1070
rect 964 935 1056 1024
rect 964 883 984 935
rect 1036 914 1056 935
rect 964 868 992 883
rect 1038 868 1056 914
rect 964 842 1056 868
rect 1216 1154 1604 1155
rect 1216 1132 1729 1154
rect 1216 1080 1459 1132
rect 1511 1080 1639 1132
rect 1691 1080 1729 1132
rect 1216 1070 1729 1080
rect 1262 1058 1729 1070
rect 1820 1121 1916 1161
rect 1820 1069 1840 1121
rect 1892 1069 1916 1121
rect 1216 914 1262 1024
rect 1216 762 1262 868
rect 1541 967 1587 1004
rect 1541 826 1587 921
rect 1765 967 1811 1004
rect 1765 884 1811 921
rect 1820 935 1916 1069
rect 2481 1121 2573 1161
rect 2481 1069 2501 1121
rect 2553 1069 2573 1121
rect 1820 883 1840 935
rect 1892 883 1916 935
rect 1989 967 2109 1004
rect 2266 978 2312 1004
rect 2035 921 2109 967
rect 1989 884 2109 921
rect 1820 842 1916 883
rect 1504 786 1596 826
rect 320 737 1413 762
rect 320 691 1324 737
rect 1370 691 1413 737
rect 320 643 1413 691
rect 1504 734 1524 786
rect 1576 734 1596 786
rect 1848 796 1916 842
rect 1848 750 1859 796
rect 1905 750 1916 796
rect 1848 739 1916 750
rect 2037 796 2109 884
rect 2037 750 2048 796
rect 2094 750 2109 796
rect 96 559 142 572
rect -356 515 -264 555
rect -356 463 -336 515
rect -284 463 -264 515
rect 96 502 142 513
rect 320 559 366 643
rect 732 642 814 643
rect 1180 642 1262 643
rect -356 425 -264 463
rect 72 472 164 502
rect -367 388 -252 425
rect -367 342 -333 388
rect -287 342 -252 388
rect -367 329 -252 342
rect -367 305 -336 329
rect -356 277 -336 305
rect -284 305 -252 329
rect 72 420 92 472
rect 144 420 164 472
rect 72 386 96 420
rect 142 386 164 420
rect 72 305 164 386
rect -284 277 -264 305
rect -356 247 -264 277
rect 72 286 96 305
rect 142 286 164 305
rect 72 234 92 286
rect 144 234 164 286
rect 72 194 164 234
rect 320 432 366 513
rect 544 559 590 572
rect 544 500 590 513
rect 768 559 814 642
rect 320 305 366 386
rect 96 177 142 194
rect 96 118 142 131
rect 320 177 366 259
rect 521 470 613 500
rect 521 418 541 470
rect 593 418 613 470
rect 521 386 544 418
rect 590 386 613 418
rect 521 305 613 386
rect 521 284 544 305
rect 590 284 613 305
rect 521 232 541 284
rect 593 232 613 284
rect 521 192 613 232
rect 768 432 814 513
rect 992 559 1038 572
rect 992 498 1038 513
rect 1216 559 1262 642
rect 768 305 814 386
rect 320 118 366 131
rect 544 177 590 192
rect 544 118 590 131
rect 768 177 814 259
rect 968 468 1060 498
rect 968 416 988 468
rect 1040 416 1060 468
rect 968 386 992 416
rect 1038 386 1060 416
rect 968 305 1060 386
rect 968 282 992 305
rect 1038 282 1060 305
rect 968 230 988 282
rect 1040 230 1060 282
rect 968 190 1060 230
rect 1216 432 1262 513
rect 1504 600 1596 734
rect 1504 548 1524 600
rect 1576 548 1596 600
rect 1504 523 1596 548
rect 1504 507 1541 523
rect 1216 305 1262 386
rect 1587 507 1596 523
rect 1765 523 1811 536
rect 1541 355 1587 477
rect 1765 435 1811 477
rect 1989 523 2035 536
rect 1541 296 1587 309
rect 1741 405 1833 435
rect 1741 353 1761 405
rect 1813 353 1833 405
rect 1741 309 1765 353
rect 1811 309 1833 353
rect 768 118 814 131
rect 992 177 1038 190
rect 992 118 1038 131
rect 1216 177 1262 259
rect 1216 118 1262 131
rect 1741 219 1833 309
rect 1989 355 2035 477
rect 2037 355 2109 750
rect 2228 967 2312 978
rect 2228 921 2266 967
rect 2228 884 2312 921
rect 2481 967 2573 1069
rect 3204 1121 3296 1161
rect 3204 1069 3224 1121
rect 3276 1069 3296 1121
rect 2481 921 2490 967
rect 2536 935 2573 967
rect 2228 746 2300 884
rect 2481 883 2501 921
rect 2553 883 2573 935
rect 2714 967 2760 1004
rect 2990 978 3036 1004
rect 2714 884 2760 921
rect 2481 842 2573 883
rect 2762 746 2834 978
rect 2950 967 3036 978
rect 2950 921 2990 967
rect 2950 884 3036 921
rect 3204 967 3296 1069
rect 3929 1121 4021 1161
rect 3929 1069 3949 1121
rect 4001 1069 4021 1121
rect 3204 921 3214 967
rect 3260 935 3296 967
rect 2950 858 3023 884
rect 2951 746 3023 858
rect 3204 883 3224 921
rect 3276 883 3296 935
rect 3204 842 3296 883
rect 3438 978 3484 1004
rect 3438 967 3571 978
rect 3484 921 3571 967
rect 3438 858 3571 921
rect 2228 735 2641 746
rect 2228 689 2584 735
rect 2630 689 2641 735
rect 2228 678 2641 689
rect 2762 735 2872 746
rect 2762 689 2815 735
rect 2861 689 2872 735
rect 2762 678 2872 689
rect 2951 735 3365 746
rect 2951 689 3308 735
rect 3354 689 3365 735
rect 2951 678 3365 689
rect 3503 735 3571 858
rect 3503 689 3514 735
rect 3560 689 3571 735
rect 2228 536 2300 678
rect 2228 523 2312 536
rect 2228 477 2266 523
rect 2228 355 2312 477
rect 2490 523 2536 536
rect 2490 435 2536 477
rect 2714 523 2760 536
rect 1989 296 2035 309
rect 2266 296 2312 309
rect 2466 405 2558 435
rect 2466 353 2486 405
rect 2538 353 2558 405
rect 2466 309 2490 353
rect 2536 309 2558 353
rect 1741 167 1761 219
rect 1813 167 1833 219
rect 1741 127 1833 167
rect 2466 219 2558 309
rect 2714 355 2760 477
rect 2762 355 2834 678
rect 2951 536 3023 678
rect 3503 536 3571 689
rect 2951 523 3036 536
rect 2951 477 2990 523
rect 2951 355 3036 477
rect 3214 523 3260 536
rect 3214 435 3260 477
rect 3438 523 3571 536
rect 3484 477 3571 523
rect 2951 347 2990 355
rect 2714 296 2760 309
rect 2990 296 3036 309
rect 3189 405 3281 435
rect 3189 353 3209 405
rect 3261 353 3281 405
rect 3189 309 3214 353
rect 3260 309 3281 353
rect 2466 167 2486 219
rect 2538 167 2558 219
rect 2466 127 2558 167
rect 3189 219 3281 309
rect 3438 355 3571 477
rect 3484 347 3571 355
rect 3715 967 3761 1004
rect 3715 561 3761 921
rect 3929 967 4021 1069
rect 3929 921 3939 967
rect 3985 935 4021 967
rect 3929 883 3949 921
rect 4001 883 4021 935
rect 3929 842 4021 883
rect 4153 1121 4245 1161
rect 4153 1069 4173 1121
rect 4225 1069 4245 1121
rect 4726 1108 5026 1139
rect 4400 1093 4446 1106
rect 4153 1047 4176 1069
rect 4222 1047 4245 1069
rect 4153 985 4245 1047
rect 4153 939 4176 985
rect 4222 939 4245 985
rect 4153 935 4245 939
rect 4153 883 4173 935
rect 4225 883 4245 935
rect 4153 877 4245 883
rect 4153 842 4176 877
rect 4222 842 4245 877
rect 4377 1053 4400 1093
rect 4446 1053 4469 1093
rect 4377 1001 4397 1053
rect 4449 1001 4469 1053
rect 4377 985 4469 1001
rect 4726 1088 4929 1108
rect 4726 1042 4774 1088
rect 4820 1056 4929 1088
rect 4981 1056 5026 1108
rect 4820 1042 4932 1056
rect 4978 1042 5026 1056
rect 4726 992 5026 1042
rect 4377 939 4400 985
rect 4446 939 4469 985
rect 4377 877 4469 939
rect 4377 867 4400 877
rect 4446 867 4469 877
rect 4176 818 4222 831
rect 4377 815 4397 867
rect 4449 815 4469 867
rect 4909 922 5001 992
rect 4909 870 4929 922
rect 4981 870 5001 922
rect 4909 830 5001 870
rect 4377 774 4469 815
rect 3979 694 4287 713
rect 3979 693 4207 694
rect 3979 641 4009 693
rect 4061 641 4195 693
rect 4253 648 4287 694
rect 4247 641 4287 648
rect 3979 621 4287 641
rect 3715 393 3761 515
rect 3715 334 3761 347
rect 3939 561 3985 574
rect 3939 435 3985 515
rect 4176 526 4222 539
rect 4176 435 4222 480
rect 4400 526 4446 774
rect 3939 405 4034 435
rect 3939 393 3962 405
rect 4014 353 4034 405
rect 3985 347 4034 353
rect 3939 334 4034 347
rect 3438 296 3484 309
rect 3189 167 3209 219
rect 3261 167 3281 219
rect 3189 127 3281 167
rect 3942 219 4034 334
rect 3942 167 3962 219
rect 4014 167 4034 219
rect 3942 127 4034 167
rect 4148 405 4240 435
rect 4148 353 4168 405
rect 4220 391 4240 405
rect 4148 345 4176 353
rect 4222 345 4240 391
rect 4148 256 4240 345
rect 4148 219 4176 256
rect 4148 167 4168 219
rect 4222 210 4240 256
rect 4220 167 4240 210
rect 4400 391 4446 480
rect 4624 526 4670 539
rect 4624 435 4670 480
rect 4400 256 4446 345
rect 4400 197 4446 210
rect 4601 405 4693 435
rect 4601 353 4621 405
rect 4673 353 4693 405
rect 4601 345 4624 353
rect 4670 345 4693 353
rect 4601 256 4693 345
rect 4601 219 4624 256
rect 4670 219 4693 256
rect 4148 127 4240 167
rect 4601 167 4621 219
rect 4673 167 4693 219
rect 4601 127 4693 167
<< via1 >>
rect -336 5458 -333 5510
rect -333 5458 -287 5510
rect -287 5458 -284 5510
rect -336 5272 -333 5324
rect -333 5272 -287 5324
rect -287 5272 -284 5324
rect 33 5439 85 5491
rect 33 5282 85 5305
rect 33 5253 84 5282
rect 84 5253 85 5282
rect 529 5439 581 5491
rect 529 5282 581 5305
rect 529 5253 532 5282
rect 532 5253 578 5282
rect 578 5253 581 5282
rect 993 5401 999 5405
rect 999 5401 1045 5405
rect 993 5353 1045 5401
rect 1432 5401 1447 5405
rect 1447 5401 1484 5405
rect 1432 5353 1484 5401
rect 993 5193 1045 5219
rect 993 5167 999 5193
rect 999 5167 1045 5193
rect 1432 5193 1484 5219
rect 1432 5167 1447 5193
rect 1447 5167 1484 5193
rect 1898 5401 1941 5405
rect 1941 5401 1950 5405
rect 1898 5353 1950 5401
rect 1898 5193 1950 5219
rect 1898 5167 1941 5193
rect 1941 5167 1950 5193
rect 81 4317 84 4369
rect 84 4317 130 4369
rect 130 4317 133 4369
rect 3815 5401 3817 5405
rect 3817 5401 3863 5405
rect 3863 5401 3867 5405
rect 3815 5353 3867 5401
rect 3815 5193 3867 5219
rect 3815 5167 3817 5193
rect 3817 5167 3863 5193
rect 3863 5167 3867 5193
rect 4261 5401 4265 5405
rect 4265 5401 4311 5405
rect 4311 5401 4313 5405
rect 4261 5353 4313 5401
rect 4261 5193 4313 5219
rect 4261 5167 4265 5193
rect 4265 5167 4311 5193
rect 4311 5167 4313 5193
rect 2313 4759 2365 4811
rect 2493 4759 2545 4811
rect 529 4317 532 4369
rect 532 4317 578 4369
rect 578 4317 581 4369
rect 81 4131 133 4183
rect 529 4131 581 4183
rect 995 4385 1047 4412
rect 995 4360 999 4385
rect 999 4360 1045 4385
rect 1045 4360 1047 4385
rect 995 4211 999 4226
rect 999 4211 1045 4226
rect 1045 4211 1047 4226
rect 995 4174 1047 4211
rect 1432 4339 1447 4369
rect 1447 4339 1484 4369
rect 1432 4317 1484 4339
rect 2073 4561 2087 4576
rect 2087 4561 2125 4576
rect 2073 4524 2125 4561
rect 1878 4339 1895 4369
rect 1895 4339 1930 4369
rect 1878 4317 1930 4339
rect 2073 4338 2125 4390
rect 2484 4385 2536 4394
rect 2484 4342 2519 4385
rect 2519 4342 2536 4385
rect 1432 4131 1484 4183
rect 1878 4131 1930 4183
rect 2484 4156 2536 4208
rect 2921 4385 2973 4394
rect 2921 4342 2967 4385
rect 2967 4342 2973 4385
rect 2921 4156 2973 4208
rect -336 3910 -284 3962
rect 881 3948 933 4000
rect 1061 3948 1113 4000
rect 3363 4385 3415 4394
rect 3363 4342 3369 4385
rect 3369 4342 3415 4385
rect 4713 5401 4759 5405
rect 4759 5401 4765 5405
rect 4713 5353 4765 5401
rect 4713 5193 4765 5219
rect 4713 5167 4759 5193
rect 4759 5167 4765 5193
rect 3363 4156 3415 4208
rect 3817 4385 3869 4394
rect 3817 4342 3863 4385
rect 3863 4342 3869 4385
rect 3817 4156 3869 4208
rect 4263 4385 4315 4394
rect 4263 4342 4265 4385
rect 4265 4342 4311 4385
rect 4311 4342 4315 4385
rect 4263 4156 4315 4208
rect 4711 4385 4763 4394
rect 4711 4342 4713 4385
rect 4713 4342 4759 4385
rect 4759 4342 4763 4385
rect 4711 4156 4763 4208
rect -336 3759 -284 3776
rect -336 3724 -333 3759
rect -333 3724 -287 3759
rect -287 3724 -284 3759
rect 4929 3799 4981 3851
rect 2816 3788 2868 3796
rect 2816 3744 2868 3788
rect 2996 3744 3048 3796
rect -336 3332 -284 3384
rect 33 3544 85 3596
rect 33 3358 85 3410
rect -336 3146 -284 3198
rect 1432 3570 1435 3596
rect 1435 3570 1481 3596
rect 1481 3570 1484 3596
rect 1432 3544 1484 3570
rect 1432 3402 1484 3410
rect 1432 3358 1435 3402
rect 1435 3358 1481 3402
rect 1481 3358 1484 3402
rect 2317 3509 2369 3553
rect 2317 3501 2331 3509
rect 2331 3501 2369 3509
rect 2796 3532 2848 3535
rect 2796 3486 2825 3532
rect 2825 3486 2848 3532
rect 2796 3483 2848 3486
rect 2317 3356 2331 3367
rect 2331 3356 2369 3367
rect 2317 3315 2369 3356
rect 2796 3322 2848 3349
rect 2796 3297 2825 3322
rect 2825 3297 2848 3322
rect 3226 3532 3278 3535
rect 3226 3486 3227 3532
rect 3227 3486 3273 3532
rect 3273 3486 3278 3532
rect 3226 3483 3278 3486
rect 3226 3322 3278 3349
rect 3226 3297 3227 3322
rect 3227 3297 3273 3322
rect 3273 3297 3278 3322
rect 2330 2690 2382 2718
rect 2330 2666 2382 2690
rect 3670 3532 3722 3535
rect 3670 3486 3675 3532
rect 3675 3486 3721 3532
rect 3721 3486 3722 3532
rect 3670 3483 3722 3486
rect 3670 3322 3722 3349
rect 3670 3297 3675 3322
rect 3675 3297 3721 3322
rect 3721 3297 3722 3322
rect 4120 3532 4172 3535
rect 4120 3486 4123 3532
rect 4123 3486 4169 3532
rect 4169 3486 4172 3532
rect 4120 3483 4172 3486
rect 4120 3322 4172 3349
rect 4120 3297 4123 3322
rect 4123 3297 4169 3322
rect 4169 3297 4172 3322
rect 4929 3613 4981 3665
rect 4929 3332 4981 3384
rect 4929 3146 4981 3198
rect 3896 2905 3948 2923
rect 3896 2871 3899 2905
rect 3899 2871 3945 2905
rect 3945 2871 3948 2905
rect 4346 2905 4398 2923
rect 4346 2871 4347 2905
rect 4347 2871 4393 2905
rect 4393 2871 4398 2905
rect 3896 2685 3948 2737
rect -336 2191 -284 2212
rect -336 2160 -333 2191
rect -333 2160 -287 2191
rect -287 2160 -284 2191
rect -336 1981 -333 2026
rect -333 1981 -287 2026
rect -287 1981 -284 2026
rect -336 1974 -284 1981
rect 2219 2433 2271 2449
rect 2219 2397 2263 2433
rect 2263 2397 2271 2433
rect 2399 2397 2451 2449
rect 1434 2160 1486 2211
rect 1434 2159 1435 2160
rect 1435 2159 1481 2160
rect 1481 2159 1486 2160
rect 1434 1987 1435 2025
rect 1435 1987 1481 2025
rect 1481 1987 1486 2025
rect 1434 1973 1486 1987
rect 2102 2159 2107 2211
rect 2107 2159 2153 2211
rect 2153 2159 2154 2211
rect 2102 1973 2107 2025
rect 2107 1973 2153 2025
rect 2153 1973 2154 2025
rect 3121 2397 3173 2449
rect 3301 2403 3332 2449
rect 3332 2403 3353 2449
rect 3301 2397 3353 2403
rect 3450 2159 3451 2211
rect 3451 2159 3497 2211
rect 3497 2159 3502 2211
rect 3450 1973 3451 2025
rect 3451 1973 3497 2025
rect 3497 1973 3502 2025
rect 4346 2685 4398 2737
rect 3672 2175 3724 2211
rect 3672 2159 3675 2175
rect 3675 2159 3721 2175
rect 3721 2159 3724 2175
rect 3672 2016 3675 2025
rect 3675 2016 3721 2025
rect 3721 2016 3724 2025
rect 3672 1973 3724 2016
rect 4118 2175 4170 2211
rect 4118 2159 4123 2175
rect 4123 2159 4169 2175
rect 4169 2159 4170 2175
rect 4118 2016 4123 2025
rect 4123 2016 4169 2025
rect 4169 2016 4170 2025
rect 4118 1973 4170 2016
rect 4929 2191 4981 2212
rect 4929 2160 4932 2191
rect 4932 2160 4978 2191
rect 4978 2160 4981 2191
rect 4929 1981 4932 2026
rect 4932 1981 4978 2026
rect 4978 1981 4981 2026
rect 4929 1974 4981 1981
rect 4611 1734 4663 1786
rect 4823 1734 4875 1786
rect 112 1516 164 1568
rect 324 1516 376 1568
rect 890 1532 942 1584
rect 1076 1532 1128 1584
rect 4191 1532 4243 1584
rect 4377 1532 4429 1584
rect 4611 1516 4663 1568
rect 4823 1516 4875 1568
rect 112 1298 164 1350
rect 324 1336 376 1350
rect 324 1298 366 1336
rect 366 1298 376 1336
rect 1983 1298 2035 1350
rect 2193 1298 2245 1350
rect 2404 1298 2456 1350
rect 2615 1298 2667 1350
rect 2826 1298 2878 1350
rect 3037 1298 3089 1350
rect 3248 1298 3300 1350
rect 3459 1298 3511 1350
rect 3670 1298 3722 1350
rect 3881 1298 3933 1350
rect 4091 1298 4143 1350
rect 4611 1298 4663 1350
rect 4823 1298 4875 1350
rect -336 1056 -284 1108
rect 92 1070 144 1121
rect 92 1069 96 1070
rect 96 1069 142 1070
rect 142 1069 144 1070
rect -336 870 -284 922
rect 92 914 144 935
rect 92 883 96 914
rect 96 883 142 914
rect 142 883 144 914
rect 512 1070 564 1121
rect 512 1069 544 1070
rect 544 1069 564 1070
rect 512 914 564 935
rect 512 883 544 914
rect 544 883 564 914
rect 984 1070 1036 1121
rect 984 1069 992 1070
rect 992 1069 1036 1070
rect 984 914 1036 935
rect 984 883 992 914
rect 992 883 1036 914
rect 1459 1080 1511 1132
rect 1639 1080 1691 1132
rect 1840 1069 1892 1121
rect 2501 1069 2553 1121
rect 1840 883 1892 935
rect 1524 734 1576 786
rect -336 463 -284 515
rect -336 277 -284 329
rect 92 432 144 472
rect 92 420 96 432
rect 96 420 142 432
rect 142 420 144 432
rect 92 259 96 286
rect 96 259 142 286
rect 142 259 144 286
rect 92 234 144 259
rect 541 432 593 470
rect 541 418 544 432
rect 544 418 590 432
rect 590 418 593 432
rect 541 259 544 284
rect 544 259 590 284
rect 590 259 593 284
rect 541 232 593 259
rect 988 432 1040 468
rect 988 416 992 432
rect 992 416 1038 432
rect 1038 416 1040 432
rect 988 259 992 282
rect 992 259 1038 282
rect 1038 259 1040 282
rect 988 230 1040 259
rect 1524 548 1576 600
rect 1761 355 1813 405
rect 1761 353 1765 355
rect 1765 353 1811 355
rect 1811 353 1813 355
rect 3224 1069 3276 1121
rect 2501 921 2536 935
rect 2536 921 2553 935
rect 2501 883 2553 921
rect 3949 1069 4001 1121
rect 3224 921 3260 935
rect 3260 921 3276 935
rect 3224 883 3276 921
rect 2486 355 2538 405
rect 2486 353 2490 355
rect 2490 353 2536 355
rect 2536 353 2538 355
rect 1761 167 1813 219
rect 3209 355 3261 405
rect 3209 353 3214 355
rect 3214 353 3260 355
rect 3260 353 3261 355
rect 2486 167 2538 219
rect 3949 921 3985 935
rect 3985 921 4001 935
rect 3949 883 4001 921
rect 4173 1093 4225 1121
rect 4173 1069 4176 1093
rect 4176 1069 4222 1093
rect 4222 1069 4225 1093
rect 4173 883 4225 935
rect 4397 1047 4400 1053
rect 4400 1047 4446 1053
rect 4446 1047 4449 1053
rect 4397 1001 4449 1047
rect 4929 1088 4981 1108
rect 4929 1056 4932 1088
rect 4932 1056 4978 1088
rect 4978 1056 4981 1088
rect 4397 831 4400 867
rect 4400 831 4446 867
rect 4446 831 4449 867
rect 4397 815 4449 831
rect 4929 870 4981 922
rect 4009 641 4061 693
rect 4195 648 4207 693
rect 4207 648 4247 693
rect 4195 641 4247 648
rect 3962 393 4014 405
rect 3962 353 3985 393
rect 3985 353 4014 393
rect 3209 167 3261 219
rect 3962 167 4014 219
rect 4168 391 4220 405
rect 4168 353 4176 391
rect 4176 353 4220 391
rect 4168 210 4176 219
rect 4176 210 4220 219
rect 4168 167 4220 210
rect 4621 391 4673 405
rect 4621 353 4624 391
rect 4624 353 4670 391
rect 4670 353 4673 391
rect 4621 210 4624 219
rect 4624 210 4670 219
rect 4670 210 4673 219
rect 4621 167 4673 210
<< metal2 >>
rect -356 5512 -264 5550
rect -356 5456 -338 5512
rect -282 5456 -264 5512
rect -356 5326 -264 5456
rect -356 5270 -338 5326
rect -282 5270 -264 5326
rect -356 5242 -264 5270
rect 13 5493 105 5531
rect 13 5437 31 5493
rect 87 5437 105 5493
rect 13 5307 105 5437
rect 13 5251 31 5307
rect 87 5251 105 5307
rect 13 5223 105 5251
rect 509 5493 601 5531
rect 509 5437 527 5493
rect 583 5437 601 5493
rect 509 5307 601 5437
rect 509 5251 527 5307
rect 583 5251 601 5307
rect 509 5223 601 5251
rect 973 5407 1065 5445
rect 973 5351 991 5407
rect 1047 5351 1065 5407
rect 973 5221 1065 5351
rect 973 5165 991 5221
rect 1047 5165 1065 5221
rect 973 5137 1065 5165
rect 1412 5407 1504 5445
rect 1412 5351 1430 5407
rect 1486 5351 1504 5407
rect 1412 5221 1504 5351
rect 1412 5165 1430 5221
rect 1486 5165 1504 5221
rect 1412 5137 1504 5165
rect 1878 5407 1970 5445
rect 1878 5351 1896 5407
rect 1952 5351 1970 5407
rect 1878 5221 1970 5351
rect 1878 5165 1896 5221
rect 1952 5165 1970 5221
rect 1878 5137 1970 5165
rect 3795 5407 3887 5445
rect 3795 5351 3813 5407
rect 3869 5351 3887 5407
rect 3795 5221 3887 5351
rect 3795 5165 3813 5221
rect 3869 5165 3887 5221
rect 3795 5137 3887 5165
rect 4241 5407 4333 5445
rect 4241 5351 4259 5407
rect 4315 5351 4333 5407
rect 4241 5221 4333 5351
rect 4241 5165 4259 5221
rect 4315 5165 4333 5221
rect 4241 5137 4333 5165
rect 4693 5407 4785 5445
rect 4693 5351 4711 5407
rect 4767 5351 4785 5407
rect 4693 5221 4785 5351
rect 4693 5165 4711 5221
rect 4767 5165 4785 5221
rect 4693 5137 4785 5165
rect 2275 4833 2364 4834
rect 2275 4811 2583 4833
rect 2275 4759 2313 4811
rect 2365 4759 2493 4811
rect 2545 4759 2583 4811
rect 2275 4737 2583 4759
rect 2053 4576 2146 4616
rect 2053 4524 2073 4576
rect 2125 4524 2146 4576
rect 975 4414 1067 4452
rect 61 4371 153 4409
rect 61 4315 79 4371
rect 135 4315 153 4371
rect 61 4185 153 4315
rect 61 4129 79 4185
rect 135 4129 153 4185
rect 61 4101 153 4129
rect 509 4371 601 4409
rect 509 4315 527 4371
rect 583 4315 601 4371
rect 509 4185 601 4315
rect 509 4129 527 4185
rect 583 4129 601 4185
rect 975 4358 993 4414
rect 1049 4358 1067 4414
rect 975 4228 1067 4358
rect 975 4172 993 4228
rect 1049 4172 1067 4228
rect 975 4144 1067 4172
rect 1412 4371 1504 4409
rect 1412 4315 1430 4371
rect 1486 4315 1504 4371
rect 1412 4185 1504 4315
rect 509 4101 601 4129
rect 1412 4129 1430 4185
rect 1486 4129 1504 4185
rect 1412 4101 1504 4129
rect 1858 4371 1950 4409
rect 1858 4315 1876 4371
rect 1932 4315 1950 4371
rect 1858 4185 1950 4315
rect 1858 4129 1876 4185
rect 1932 4129 1950 4185
rect 1858 4101 1950 4129
rect 2053 4390 2146 4524
rect 2053 4338 2073 4390
rect 2125 4338 2146 4390
rect 860 4000 1134 4040
rect -356 3964 -264 3992
rect -356 3908 -338 3964
rect -282 3908 -264 3964
rect -356 3778 -264 3908
rect -356 3722 -338 3778
rect -282 3722 -264 3778
rect -356 3684 -264 3722
rect 860 3948 881 4000
rect 933 3948 1061 4000
rect 1113 3948 1134 4000
rect 860 3907 1134 3948
rect 13 3598 105 3636
rect 13 3542 31 3598
rect 87 3542 105 3598
rect -356 3386 -264 3414
rect -356 3330 -338 3386
rect -282 3330 -264 3386
rect -356 3200 -264 3330
rect 13 3412 105 3542
rect 13 3356 31 3412
rect 87 3356 105 3412
rect 13 3328 105 3356
rect -356 3144 -338 3200
rect -282 3144 -264 3200
rect -356 3106 -264 3144
rect -356 2214 -264 2242
rect -356 2158 -338 2214
rect -282 2158 -264 2214
rect -356 2028 -264 2158
rect -356 1972 -338 2028
rect -282 1972 -264 2028
rect -356 1934 -264 1972
rect 199 1608 294 1609
rect 74 1570 414 1608
rect 74 1514 110 1570
rect 166 1514 322 1570
rect 378 1514 414 1570
rect 74 1352 414 1514
rect 860 1604 954 3907
rect 2053 3805 2146 4338
rect 2275 3997 2364 4737
rect 2464 4396 2556 4434
rect 2464 4340 2482 4396
rect 2538 4340 2556 4396
rect 2464 4210 2556 4340
rect 2464 4154 2482 4210
rect 2538 4154 2556 4210
rect 2464 4126 2556 4154
rect 2901 4396 2993 4434
rect 2901 4340 2919 4396
rect 2975 4340 2993 4396
rect 2901 4210 2993 4340
rect 2901 4154 2919 4210
rect 2975 4154 2993 4210
rect 2901 4126 2993 4154
rect 3343 4396 3435 4434
rect 3343 4340 3361 4396
rect 3417 4340 3435 4396
rect 3343 4210 3435 4340
rect 3343 4154 3361 4210
rect 3417 4154 3435 4210
rect 3343 4126 3435 4154
rect 3797 4396 3889 4434
rect 3797 4340 3815 4396
rect 3871 4340 3889 4396
rect 3797 4210 3889 4340
rect 3797 4154 3815 4210
rect 3871 4154 3889 4210
rect 3797 4126 3889 4154
rect 4243 4396 4335 4434
rect 4243 4340 4261 4396
rect 4317 4340 4335 4396
rect 4243 4210 4335 4340
rect 4243 4154 4261 4210
rect 4317 4154 4335 4210
rect 4243 4126 4335 4154
rect 4691 4396 4783 4434
rect 4691 4340 4709 4396
rect 4765 4340 4783 4396
rect 4691 4210 4783 4340
rect 4691 4154 4709 4210
rect 4765 4154 4783 4210
rect 4691 4126 4783 4154
rect 2275 3905 2867 3997
rect 2777 3818 2867 3905
rect 4909 3853 5001 3881
rect 2053 3708 2685 3805
rect 2777 3796 3086 3818
rect 2777 3744 2816 3796
rect 2868 3744 2996 3796
rect 3048 3744 3086 3796
rect 2777 3722 3086 3744
rect 4909 3797 4927 3853
rect 4983 3797 5001 3853
rect 2777 3721 2867 3722
rect 2590 3707 2685 3708
rect 1412 3598 1504 3636
rect 1412 3542 1430 3598
rect 1486 3542 1504 3598
rect 1412 3412 1504 3542
rect 1412 3356 1430 3412
rect 1486 3356 1504 3412
rect 1412 3328 1504 3356
rect 2297 3555 2389 3593
rect 2297 3499 2315 3555
rect 2371 3499 2389 3555
rect 2297 3369 2389 3499
rect 2297 3313 2315 3369
rect 2371 3313 2389 3369
rect 2297 3285 2389 3313
rect 2295 2738 2422 2739
rect 2189 2720 2497 2738
rect 2189 2664 2217 2720
rect 2273 2718 2403 2720
rect 2273 2666 2330 2718
rect 2382 2666 2403 2718
rect 2273 2664 2403 2666
rect 2459 2664 2497 2720
rect 2189 2646 2497 2664
rect 2591 2472 2685 3707
rect 4909 3667 5001 3797
rect 4909 3611 4927 3667
rect 4983 3611 5001 3667
rect 2776 3537 2868 3575
rect 2776 3481 2794 3537
rect 2850 3481 2868 3537
rect 2776 3351 2868 3481
rect 2776 3295 2794 3351
rect 2850 3295 2868 3351
rect 2776 3267 2868 3295
rect 3206 3537 3298 3575
rect 3206 3481 3224 3537
rect 3280 3481 3298 3537
rect 3206 3351 3298 3481
rect 3206 3295 3224 3351
rect 3280 3295 3298 3351
rect 3206 3267 3298 3295
rect 3650 3537 3742 3575
rect 3650 3481 3668 3537
rect 3724 3481 3742 3537
rect 3650 3351 3742 3481
rect 3650 3295 3668 3351
rect 3724 3295 3742 3351
rect 3650 3267 3742 3295
rect 4100 3537 4192 3575
rect 4909 3573 5001 3611
rect 4100 3481 4118 3537
rect 4174 3481 4192 3537
rect 4100 3351 4192 3481
rect 4100 3295 4118 3351
rect 4174 3295 4192 3351
rect 4100 3267 4192 3295
rect 4909 3386 5001 3414
rect 4909 3330 4927 3386
rect 4983 3330 5001 3386
rect 4909 3200 5001 3330
rect 4909 3144 4927 3200
rect 4983 3144 5001 3200
rect 4909 3106 5001 3144
rect 3876 2925 3968 2963
rect 3876 2869 3894 2925
rect 3950 2869 3968 2925
rect 3876 2739 3968 2869
rect 3876 2683 3894 2739
rect 3950 2683 3968 2739
rect 3876 2655 3968 2683
rect 4326 2925 4418 2963
rect 4326 2869 4344 2925
rect 4400 2869 4418 2925
rect 4326 2739 4418 2869
rect 4326 2683 4344 2739
rect 4400 2683 4418 2739
rect 4326 2655 4418 2683
rect 1635 2471 3280 2472
rect 1635 2449 3391 2471
rect 1635 2397 2219 2449
rect 2271 2397 2399 2449
rect 2451 2397 3121 2449
rect 3173 2397 3301 2449
rect 3353 2397 3391 2449
rect 1635 2375 3391 2397
rect 1414 2213 1506 2251
rect 1414 2157 1432 2213
rect 1488 2157 1506 2213
rect 1414 2027 1506 2157
rect 1414 1971 1432 2027
rect 1488 1971 1506 2027
rect 1414 1943 1506 1971
rect 860 1584 1168 1604
rect 860 1532 890 1584
rect 942 1532 1076 1584
rect 1128 1532 1168 1584
rect 860 1512 1168 1532
rect 860 1511 954 1512
rect 74 1296 110 1352
rect 166 1296 322 1352
rect 378 1296 414 1352
rect 74 1257 414 1296
rect 72 1150 164 1161
rect 492 1150 584 1161
rect 964 1150 1056 1161
rect 1421 1154 1510 1155
rect 1635 1154 1729 2375
rect 2082 2213 2174 2251
rect 2082 2157 2100 2213
rect 2156 2157 2174 2213
rect 2082 2027 2174 2157
rect 2082 1971 2100 2027
rect 2156 1971 2174 2027
rect 2082 1943 2174 1971
rect 3430 2213 3522 2251
rect 3430 2157 3448 2213
rect 3504 2157 3522 2213
rect 3430 2027 3522 2157
rect 3430 1971 3448 2027
rect 3504 1971 3522 2027
rect 3430 1943 3522 1971
rect 3652 2213 3744 2251
rect 3652 2157 3670 2213
rect 3726 2157 3744 2213
rect 3652 2027 3744 2157
rect 3652 1971 3670 2027
rect 3726 1971 3744 2027
rect 3652 1943 3744 1971
rect 4098 2213 4190 2251
rect 4098 2157 4116 2213
rect 4172 2157 4190 2213
rect 4098 2027 4190 2157
rect 4098 1971 4116 2027
rect 4172 1971 4190 2027
rect 4098 1943 4190 1971
rect 4909 2214 5001 2242
rect 4909 2158 4927 2214
rect 4983 2158 5001 2214
rect 4909 2028 5001 2158
rect 4909 1972 4927 2028
rect 4983 1972 5001 2028
rect 4909 1934 5001 1972
rect 4574 1788 4955 1826
rect 4574 1732 4609 1788
rect 4665 1732 4821 1788
rect 4877 1732 4955 1788
rect 4376 1604 4470 1608
rect 4161 1584 4470 1604
rect 4161 1532 4191 1584
rect 4243 1532 4377 1584
rect 4429 1532 4470 1584
rect 4161 1512 4470 1532
rect 1945 1352 4182 1390
rect 1945 1296 1981 1352
rect 2037 1296 2191 1352
rect 2247 1296 2402 1352
rect 2458 1296 2613 1352
rect 2669 1296 2824 1352
rect 2880 1296 3035 1352
rect 3091 1296 3246 1352
rect 3302 1296 3457 1352
rect 3513 1296 3668 1352
rect 3724 1296 3879 1352
rect 3935 1296 4089 1352
rect 4145 1296 4182 1352
rect 1945 1257 4182 1296
rect -356 1110 -264 1138
rect -356 1054 -338 1110
rect -282 1054 -264 1110
rect -356 924 -264 1054
rect -356 868 -338 924
rect -282 868 -264 924
rect -356 830 -264 868
rect 72 1121 165 1150
rect 72 1112 92 1121
rect 144 1112 165 1121
rect 72 1056 90 1112
rect 146 1056 165 1112
rect 72 935 165 1056
rect 72 926 92 935
rect 144 926 165 935
rect 72 870 90 926
rect 146 870 165 926
rect 72 831 165 870
rect 492 1121 585 1150
rect 492 1112 512 1121
rect 564 1112 585 1121
rect 492 1056 510 1112
rect 566 1056 585 1112
rect 492 935 585 1056
rect 492 926 512 935
rect 564 926 585 935
rect 492 870 510 926
rect 566 870 585 926
rect 492 831 585 870
rect 964 1121 1057 1150
rect 964 1112 984 1121
rect 1036 1112 1057 1121
rect 964 1056 982 1112
rect 1038 1056 1057 1112
rect 1421 1132 1729 1154
rect 1421 1080 1459 1132
rect 1511 1080 1639 1132
rect 1691 1080 1729 1132
rect 1421 1058 1729 1080
rect 1820 1150 1912 1161
rect 2481 1150 2573 1161
rect 3204 1150 3296 1161
rect 3929 1150 4021 1161
rect 4153 1150 4245 1161
rect 1820 1121 1913 1150
rect 1820 1112 1840 1121
rect 1892 1112 1913 1121
rect 964 935 1057 1056
rect 964 926 984 935
rect 1036 926 1057 935
rect 964 870 982 926
rect 1038 870 1057 926
rect 964 831 1057 870
rect 1820 1056 1838 1112
rect 1894 1056 1913 1112
rect 1820 935 1913 1056
rect 1820 926 1840 935
rect 1892 926 1913 935
rect 1820 870 1838 926
rect 1894 870 1913 926
rect 1820 831 1913 870
rect 2481 1121 2574 1150
rect 2481 1112 2501 1121
rect 2553 1112 2574 1121
rect 2481 1056 2499 1112
rect 2555 1056 2574 1112
rect 2481 935 2574 1056
rect 2481 926 2501 935
rect 2553 926 2574 935
rect 2481 870 2499 926
rect 2555 870 2574 926
rect 2481 831 2574 870
rect 3204 1121 3297 1150
rect 3204 1112 3224 1121
rect 3276 1112 3297 1121
rect 3204 1056 3222 1112
rect 3278 1056 3297 1112
rect 3204 935 3297 1056
rect 3204 926 3224 935
rect 3276 926 3297 935
rect 3204 870 3222 926
rect 3278 870 3297 926
rect 3204 831 3297 870
rect 3929 1121 4022 1150
rect 3929 1112 3949 1121
rect 4001 1112 4022 1121
rect 3929 1056 3947 1112
rect 4003 1056 4022 1112
rect 3929 935 4022 1056
rect 3929 926 3949 935
rect 4001 926 4022 935
rect 3929 870 3947 926
rect 4003 870 4022 926
rect 3929 831 4022 870
rect 4153 1121 4246 1150
rect 4153 1112 4173 1121
rect 4225 1112 4246 1121
rect 4153 1056 4171 1112
rect 4227 1056 4246 1112
rect 4153 935 4246 1056
rect 4153 926 4173 935
rect 4225 926 4246 935
rect 4153 870 4171 926
rect 4227 870 4246 926
rect 4153 831 4246 870
rect 4376 1053 4470 1512
rect 4574 1570 4955 1732
rect 4574 1514 4609 1570
rect 4665 1514 4821 1570
rect 4877 1514 4955 1570
rect 4574 1352 4955 1514
rect 4574 1296 4609 1352
rect 4665 1296 4821 1352
rect 4877 1296 4955 1352
rect 4574 1257 4955 1296
rect 4376 1001 4397 1053
rect 4449 1001 4470 1053
rect 4376 867 4470 1001
rect 1504 786 1596 826
rect 1504 734 1524 786
rect 1576 734 1596 786
rect 4376 815 4397 867
rect 4449 815 4470 867
rect 4909 1110 5001 1138
rect 4909 1054 4927 1110
rect 4983 1054 5001 1110
rect 4909 924 5001 1054
rect 4909 868 4927 924
rect 4983 868 5001 924
rect 4909 830 5001 868
rect 4376 777 4470 815
rect 4377 775 4469 777
rect 1504 717 1596 734
rect 1504 713 3989 717
rect 1504 693 4287 713
rect 1504 641 4009 693
rect 4061 641 4195 693
rect 4247 641 4287 693
rect 1504 621 4287 641
rect 1504 620 3989 621
rect 1504 600 1596 620
rect -356 517 -264 555
rect -356 461 -338 517
rect -282 461 -264 517
rect 1504 548 1524 600
rect 1576 548 1596 600
rect 1504 508 1596 548
rect -356 331 -264 461
rect -356 275 -338 331
rect -282 275 -264 331
rect -356 247 -264 275
rect 72 474 164 502
rect 72 418 90 474
rect 146 418 164 474
rect 72 288 164 418
rect 72 232 90 288
rect 146 232 164 288
rect 72 194 164 232
rect 521 472 613 500
rect 521 416 539 472
rect 595 416 613 472
rect 521 286 613 416
rect 521 230 539 286
rect 595 230 613 286
rect 521 192 613 230
rect 968 470 1060 498
rect 968 414 986 470
rect 1042 414 1060 470
rect 968 284 1060 414
rect 968 228 986 284
rect 1042 228 1060 284
rect 968 190 1060 228
rect 1741 407 1833 435
rect 1741 351 1759 407
rect 1815 351 1833 407
rect 1741 221 1833 351
rect 1741 165 1759 221
rect 1815 165 1833 221
rect 1741 127 1833 165
rect 2466 407 2558 435
rect 2466 351 2484 407
rect 2540 351 2558 407
rect 2466 221 2558 351
rect 2466 165 2484 221
rect 2540 165 2558 221
rect 2466 127 2558 165
rect 3189 407 3281 435
rect 3189 351 3207 407
rect 3263 351 3281 407
rect 3189 221 3281 351
rect 3189 165 3207 221
rect 3263 165 3281 221
rect 3189 127 3281 165
rect 3942 407 4034 435
rect 3942 351 3960 407
rect 4016 351 4034 407
rect 3942 221 4034 351
rect 3942 165 3960 221
rect 4016 165 4034 221
rect 3942 127 4034 165
rect 4148 407 4240 435
rect 4148 351 4166 407
rect 4222 351 4240 407
rect 4148 221 4240 351
rect 4148 165 4166 221
rect 4222 165 4240 221
rect 4148 127 4240 165
rect 4601 407 4693 435
rect 4601 351 4619 407
rect 4675 351 4693 407
rect 4601 221 4693 351
rect 4601 165 4619 221
rect 4675 165 4693 221
rect 4601 127 4693 165
<< via2 >>
rect -338 5510 -282 5512
rect -338 5458 -336 5510
rect -336 5458 -284 5510
rect -284 5458 -282 5510
rect -338 5456 -282 5458
rect -338 5324 -282 5326
rect -338 5272 -336 5324
rect -336 5272 -284 5324
rect -284 5272 -282 5324
rect -338 5270 -282 5272
rect 31 5491 87 5493
rect 31 5439 33 5491
rect 33 5439 85 5491
rect 85 5439 87 5491
rect 31 5437 87 5439
rect 31 5305 87 5307
rect 31 5253 33 5305
rect 33 5253 85 5305
rect 85 5253 87 5305
rect 31 5251 87 5253
rect 527 5491 583 5493
rect 527 5439 529 5491
rect 529 5439 581 5491
rect 581 5439 583 5491
rect 527 5437 583 5439
rect 527 5305 583 5307
rect 527 5253 529 5305
rect 529 5253 581 5305
rect 581 5253 583 5305
rect 527 5251 583 5253
rect 991 5405 1047 5407
rect 991 5353 993 5405
rect 993 5353 1045 5405
rect 1045 5353 1047 5405
rect 991 5351 1047 5353
rect 991 5219 1047 5221
rect 991 5167 993 5219
rect 993 5167 1045 5219
rect 1045 5167 1047 5219
rect 991 5165 1047 5167
rect 1430 5405 1486 5407
rect 1430 5353 1432 5405
rect 1432 5353 1484 5405
rect 1484 5353 1486 5405
rect 1430 5351 1486 5353
rect 1430 5219 1486 5221
rect 1430 5167 1432 5219
rect 1432 5167 1484 5219
rect 1484 5167 1486 5219
rect 1430 5165 1486 5167
rect 1896 5405 1952 5407
rect 1896 5353 1898 5405
rect 1898 5353 1950 5405
rect 1950 5353 1952 5405
rect 1896 5351 1952 5353
rect 1896 5219 1952 5221
rect 1896 5167 1898 5219
rect 1898 5167 1950 5219
rect 1950 5167 1952 5219
rect 1896 5165 1952 5167
rect 3813 5405 3869 5407
rect 3813 5353 3815 5405
rect 3815 5353 3867 5405
rect 3867 5353 3869 5405
rect 3813 5351 3869 5353
rect 3813 5219 3869 5221
rect 3813 5167 3815 5219
rect 3815 5167 3867 5219
rect 3867 5167 3869 5219
rect 3813 5165 3869 5167
rect 4259 5405 4315 5407
rect 4259 5353 4261 5405
rect 4261 5353 4313 5405
rect 4313 5353 4315 5405
rect 4259 5351 4315 5353
rect 4259 5219 4315 5221
rect 4259 5167 4261 5219
rect 4261 5167 4313 5219
rect 4313 5167 4315 5219
rect 4259 5165 4315 5167
rect 4711 5405 4767 5407
rect 4711 5353 4713 5405
rect 4713 5353 4765 5405
rect 4765 5353 4767 5405
rect 4711 5351 4767 5353
rect 4711 5219 4767 5221
rect 4711 5167 4713 5219
rect 4713 5167 4765 5219
rect 4765 5167 4767 5219
rect 4711 5165 4767 5167
rect 79 4369 135 4371
rect 79 4317 81 4369
rect 81 4317 133 4369
rect 133 4317 135 4369
rect 79 4315 135 4317
rect 79 4183 135 4185
rect 79 4131 81 4183
rect 81 4131 133 4183
rect 133 4131 135 4183
rect 79 4129 135 4131
rect 527 4369 583 4371
rect 527 4317 529 4369
rect 529 4317 581 4369
rect 581 4317 583 4369
rect 527 4315 583 4317
rect 527 4183 583 4185
rect 527 4131 529 4183
rect 529 4131 581 4183
rect 581 4131 583 4183
rect 527 4129 583 4131
rect 993 4412 1049 4414
rect 993 4360 995 4412
rect 995 4360 1047 4412
rect 1047 4360 1049 4412
rect 993 4358 1049 4360
rect 993 4226 1049 4228
rect 993 4174 995 4226
rect 995 4174 1047 4226
rect 1047 4174 1049 4226
rect 993 4172 1049 4174
rect 1430 4369 1486 4371
rect 1430 4317 1432 4369
rect 1432 4317 1484 4369
rect 1484 4317 1486 4369
rect 1430 4315 1486 4317
rect 1430 4183 1486 4185
rect 1430 4131 1432 4183
rect 1432 4131 1484 4183
rect 1484 4131 1486 4183
rect 1430 4129 1486 4131
rect 1876 4369 1932 4371
rect 1876 4317 1878 4369
rect 1878 4317 1930 4369
rect 1930 4317 1932 4369
rect 1876 4315 1932 4317
rect 1876 4183 1932 4185
rect 1876 4131 1878 4183
rect 1878 4131 1930 4183
rect 1930 4131 1932 4183
rect 1876 4129 1932 4131
rect -338 3962 -282 3964
rect -338 3910 -336 3962
rect -336 3910 -284 3962
rect -284 3910 -282 3962
rect -338 3908 -282 3910
rect -338 3776 -282 3778
rect -338 3724 -336 3776
rect -336 3724 -284 3776
rect -284 3724 -282 3776
rect -338 3722 -282 3724
rect 31 3596 87 3598
rect 31 3544 33 3596
rect 33 3544 85 3596
rect 85 3544 87 3596
rect 31 3542 87 3544
rect -338 3384 -282 3386
rect -338 3332 -336 3384
rect -336 3332 -284 3384
rect -284 3332 -282 3384
rect -338 3330 -282 3332
rect 31 3410 87 3412
rect 31 3358 33 3410
rect 33 3358 85 3410
rect 85 3358 87 3410
rect 31 3356 87 3358
rect -338 3198 -282 3200
rect -338 3146 -336 3198
rect -336 3146 -284 3198
rect -284 3146 -282 3198
rect -338 3144 -282 3146
rect -338 2212 -282 2214
rect -338 2160 -336 2212
rect -336 2160 -284 2212
rect -284 2160 -282 2212
rect -338 2158 -282 2160
rect -338 2026 -282 2028
rect -338 1974 -336 2026
rect -336 1974 -284 2026
rect -284 1974 -282 2026
rect -338 1972 -282 1974
rect 110 1568 166 1570
rect 110 1516 112 1568
rect 112 1516 164 1568
rect 164 1516 166 1568
rect 110 1514 166 1516
rect 322 1568 378 1570
rect 322 1516 324 1568
rect 324 1516 376 1568
rect 376 1516 378 1568
rect 322 1514 378 1516
rect 2482 4394 2538 4396
rect 2482 4342 2484 4394
rect 2484 4342 2536 4394
rect 2536 4342 2538 4394
rect 2482 4340 2538 4342
rect 2482 4208 2538 4210
rect 2482 4156 2484 4208
rect 2484 4156 2536 4208
rect 2536 4156 2538 4208
rect 2482 4154 2538 4156
rect 2919 4394 2975 4396
rect 2919 4342 2921 4394
rect 2921 4342 2973 4394
rect 2973 4342 2975 4394
rect 2919 4340 2975 4342
rect 2919 4208 2975 4210
rect 2919 4156 2921 4208
rect 2921 4156 2973 4208
rect 2973 4156 2975 4208
rect 2919 4154 2975 4156
rect 3361 4394 3417 4396
rect 3361 4342 3363 4394
rect 3363 4342 3415 4394
rect 3415 4342 3417 4394
rect 3361 4340 3417 4342
rect 3361 4208 3417 4210
rect 3361 4156 3363 4208
rect 3363 4156 3415 4208
rect 3415 4156 3417 4208
rect 3361 4154 3417 4156
rect 3815 4394 3871 4396
rect 3815 4342 3817 4394
rect 3817 4342 3869 4394
rect 3869 4342 3871 4394
rect 3815 4340 3871 4342
rect 3815 4208 3871 4210
rect 3815 4156 3817 4208
rect 3817 4156 3869 4208
rect 3869 4156 3871 4208
rect 3815 4154 3871 4156
rect 4261 4394 4317 4396
rect 4261 4342 4263 4394
rect 4263 4342 4315 4394
rect 4315 4342 4317 4394
rect 4261 4340 4317 4342
rect 4261 4208 4317 4210
rect 4261 4156 4263 4208
rect 4263 4156 4315 4208
rect 4315 4156 4317 4208
rect 4261 4154 4317 4156
rect 4709 4394 4765 4396
rect 4709 4342 4711 4394
rect 4711 4342 4763 4394
rect 4763 4342 4765 4394
rect 4709 4340 4765 4342
rect 4709 4208 4765 4210
rect 4709 4156 4711 4208
rect 4711 4156 4763 4208
rect 4763 4156 4765 4208
rect 4709 4154 4765 4156
rect 4927 3851 4983 3853
rect 4927 3799 4929 3851
rect 4929 3799 4981 3851
rect 4981 3799 4983 3851
rect 4927 3797 4983 3799
rect 1430 3596 1486 3598
rect 1430 3544 1432 3596
rect 1432 3544 1484 3596
rect 1484 3544 1486 3596
rect 1430 3542 1486 3544
rect 1430 3410 1486 3412
rect 1430 3358 1432 3410
rect 1432 3358 1484 3410
rect 1484 3358 1486 3410
rect 1430 3356 1486 3358
rect 2315 3553 2371 3555
rect 2315 3501 2317 3553
rect 2317 3501 2369 3553
rect 2369 3501 2371 3553
rect 2315 3499 2371 3501
rect 2315 3367 2371 3369
rect 2315 3315 2317 3367
rect 2317 3315 2369 3367
rect 2369 3315 2371 3367
rect 2315 3313 2371 3315
rect 2217 2664 2273 2720
rect 2403 2664 2459 2720
rect 4927 3665 4983 3667
rect 4927 3613 4929 3665
rect 4929 3613 4981 3665
rect 4981 3613 4983 3665
rect 4927 3611 4983 3613
rect 2794 3535 2850 3537
rect 2794 3483 2796 3535
rect 2796 3483 2848 3535
rect 2848 3483 2850 3535
rect 2794 3481 2850 3483
rect 2794 3349 2850 3351
rect 2794 3297 2796 3349
rect 2796 3297 2848 3349
rect 2848 3297 2850 3349
rect 2794 3295 2850 3297
rect 3224 3535 3280 3537
rect 3224 3483 3226 3535
rect 3226 3483 3278 3535
rect 3278 3483 3280 3535
rect 3224 3481 3280 3483
rect 3224 3349 3280 3351
rect 3224 3297 3226 3349
rect 3226 3297 3278 3349
rect 3278 3297 3280 3349
rect 3224 3295 3280 3297
rect 3668 3535 3724 3537
rect 3668 3483 3670 3535
rect 3670 3483 3722 3535
rect 3722 3483 3724 3535
rect 3668 3481 3724 3483
rect 3668 3349 3724 3351
rect 3668 3297 3670 3349
rect 3670 3297 3722 3349
rect 3722 3297 3724 3349
rect 3668 3295 3724 3297
rect 4118 3535 4174 3537
rect 4118 3483 4120 3535
rect 4120 3483 4172 3535
rect 4172 3483 4174 3535
rect 4118 3481 4174 3483
rect 4118 3349 4174 3351
rect 4118 3297 4120 3349
rect 4120 3297 4172 3349
rect 4172 3297 4174 3349
rect 4118 3295 4174 3297
rect 4927 3384 4983 3386
rect 4927 3332 4929 3384
rect 4929 3332 4981 3384
rect 4981 3332 4983 3384
rect 4927 3330 4983 3332
rect 4927 3198 4983 3200
rect 4927 3146 4929 3198
rect 4929 3146 4981 3198
rect 4981 3146 4983 3198
rect 4927 3144 4983 3146
rect 3894 2923 3950 2925
rect 3894 2871 3896 2923
rect 3896 2871 3948 2923
rect 3948 2871 3950 2923
rect 3894 2869 3950 2871
rect 3894 2737 3950 2739
rect 3894 2685 3896 2737
rect 3896 2685 3948 2737
rect 3948 2685 3950 2737
rect 3894 2683 3950 2685
rect 4344 2923 4400 2925
rect 4344 2871 4346 2923
rect 4346 2871 4398 2923
rect 4398 2871 4400 2923
rect 4344 2869 4400 2871
rect 4344 2737 4400 2739
rect 4344 2685 4346 2737
rect 4346 2685 4398 2737
rect 4398 2685 4400 2737
rect 4344 2683 4400 2685
rect 1432 2211 1488 2213
rect 1432 2159 1434 2211
rect 1434 2159 1486 2211
rect 1486 2159 1488 2211
rect 1432 2157 1488 2159
rect 1432 2025 1488 2027
rect 1432 1973 1434 2025
rect 1434 1973 1486 2025
rect 1486 1973 1488 2025
rect 1432 1971 1488 1973
rect 110 1350 166 1352
rect 110 1298 112 1350
rect 112 1298 164 1350
rect 164 1298 166 1350
rect 110 1296 166 1298
rect 322 1350 378 1352
rect 322 1298 324 1350
rect 324 1298 376 1350
rect 376 1298 378 1350
rect 322 1296 378 1298
rect 2100 2211 2156 2213
rect 2100 2159 2102 2211
rect 2102 2159 2154 2211
rect 2154 2159 2156 2211
rect 2100 2157 2156 2159
rect 2100 2025 2156 2027
rect 2100 1973 2102 2025
rect 2102 1973 2154 2025
rect 2154 1973 2156 2025
rect 2100 1971 2156 1973
rect 3448 2211 3504 2213
rect 3448 2159 3450 2211
rect 3450 2159 3502 2211
rect 3502 2159 3504 2211
rect 3448 2157 3504 2159
rect 3448 2025 3504 2027
rect 3448 1973 3450 2025
rect 3450 1973 3502 2025
rect 3502 1973 3504 2025
rect 3448 1971 3504 1973
rect 3670 2211 3726 2213
rect 3670 2159 3672 2211
rect 3672 2159 3724 2211
rect 3724 2159 3726 2211
rect 3670 2157 3726 2159
rect 3670 2025 3726 2027
rect 3670 1973 3672 2025
rect 3672 1973 3724 2025
rect 3724 1973 3726 2025
rect 3670 1971 3726 1973
rect 4116 2211 4172 2213
rect 4116 2159 4118 2211
rect 4118 2159 4170 2211
rect 4170 2159 4172 2211
rect 4116 2157 4172 2159
rect 4116 2025 4172 2027
rect 4116 1973 4118 2025
rect 4118 1973 4170 2025
rect 4170 1973 4172 2025
rect 4116 1971 4172 1973
rect 4927 2212 4983 2214
rect 4927 2160 4929 2212
rect 4929 2160 4981 2212
rect 4981 2160 4983 2212
rect 4927 2158 4983 2160
rect 4927 2026 4983 2028
rect 4927 1974 4929 2026
rect 4929 1974 4981 2026
rect 4981 1974 4983 2026
rect 4927 1972 4983 1974
rect 4609 1786 4665 1788
rect 4609 1734 4611 1786
rect 4611 1734 4663 1786
rect 4663 1734 4665 1786
rect 4609 1732 4665 1734
rect 4821 1786 4877 1788
rect 4821 1734 4823 1786
rect 4823 1734 4875 1786
rect 4875 1734 4877 1786
rect 4821 1732 4877 1734
rect 1981 1350 2037 1352
rect 1981 1298 1983 1350
rect 1983 1298 2035 1350
rect 2035 1298 2037 1350
rect 1981 1296 2037 1298
rect 2191 1350 2247 1352
rect 2191 1298 2193 1350
rect 2193 1298 2245 1350
rect 2245 1298 2247 1350
rect 2191 1296 2247 1298
rect 2402 1350 2458 1352
rect 2402 1298 2404 1350
rect 2404 1298 2456 1350
rect 2456 1298 2458 1350
rect 2402 1296 2458 1298
rect 2613 1350 2669 1352
rect 2613 1298 2615 1350
rect 2615 1298 2667 1350
rect 2667 1298 2669 1350
rect 2613 1296 2669 1298
rect 2824 1350 2880 1352
rect 2824 1298 2826 1350
rect 2826 1298 2878 1350
rect 2878 1298 2880 1350
rect 2824 1296 2880 1298
rect 3035 1350 3091 1352
rect 3035 1298 3037 1350
rect 3037 1298 3089 1350
rect 3089 1298 3091 1350
rect 3035 1296 3091 1298
rect 3246 1350 3302 1352
rect 3246 1298 3248 1350
rect 3248 1298 3300 1350
rect 3300 1298 3302 1350
rect 3246 1296 3302 1298
rect 3457 1350 3513 1352
rect 3457 1298 3459 1350
rect 3459 1298 3511 1350
rect 3511 1298 3513 1350
rect 3457 1296 3513 1298
rect 3668 1350 3724 1352
rect 3668 1298 3670 1350
rect 3670 1298 3722 1350
rect 3722 1298 3724 1350
rect 3668 1296 3724 1298
rect 3879 1350 3935 1352
rect 3879 1298 3881 1350
rect 3881 1298 3933 1350
rect 3933 1298 3935 1350
rect 3879 1296 3935 1298
rect 4089 1350 4145 1352
rect 4089 1298 4091 1350
rect 4091 1298 4143 1350
rect 4143 1298 4145 1350
rect 4089 1296 4145 1298
rect -338 1108 -282 1110
rect -338 1056 -336 1108
rect -336 1056 -284 1108
rect -284 1056 -282 1108
rect -338 1054 -282 1056
rect -338 922 -282 924
rect -338 870 -336 922
rect -336 870 -284 922
rect -284 870 -282 922
rect -338 868 -282 870
rect 90 1069 92 1112
rect 92 1069 144 1112
rect 144 1069 146 1112
rect 90 1056 146 1069
rect 90 883 92 926
rect 92 883 144 926
rect 144 883 146 926
rect 90 870 146 883
rect 510 1069 512 1112
rect 512 1069 564 1112
rect 564 1069 566 1112
rect 510 1056 566 1069
rect 510 883 512 926
rect 512 883 564 926
rect 564 883 566 926
rect 510 870 566 883
rect 982 1069 984 1112
rect 984 1069 1036 1112
rect 1036 1069 1038 1112
rect 982 1056 1038 1069
rect 982 883 984 926
rect 984 883 1036 926
rect 1036 883 1038 926
rect 982 870 1038 883
rect 1838 1069 1840 1112
rect 1840 1069 1892 1112
rect 1892 1069 1894 1112
rect 1838 1056 1894 1069
rect 1838 883 1840 926
rect 1840 883 1892 926
rect 1892 883 1894 926
rect 1838 870 1894 883
rect 2499 1069 2501 1112
rect 2501 1069 2553 1112
rect 2553 1069 2555 1112
rect 2499 1056 2555 1069
rect 2499 883 2501 926
rect 2501 883 2553 926
rect 2553 883 2555 926
rect 2499 870 2555 883
rect 3222 1069 3224 1112
rect 3224 1069 3276 1112
rect 3276 1069 3278 1112
rect 3222 1056 3278 1069
rect 3222 883 3224 926
rect 3224 883 3276 926
rect 3276 883 3278 926
rect 3222 870 3278 883
rect 3947 1069 3949 1112
rect 3949 1069 4001 1112
rect 4001 1069 4003 1112
rect 3947 1056 4003 1069
rect 3947 883 3949 926
rect 3949 883 4001 926
rect 4001 883 4003 926
rect 3947 870 4003 883
rect 4171 1069 4173 1112
rect 4173 1069 4225 1112
rect 4225 1069 4227 1112
rect 4171 1056 4227 1069
rect 4171 883 4173 926
rect 4173 883 4225 926
rect 4225 883 4227 926
rect 4171 870 4227 883
rect 4609 1568 4665 1570
rect 4609 1516 4611 1568
rect 4611 1516 4663 1568
rect 4663 1516 4665 1568
rect 4609 1514 4665 1516
rect 4821 1568 4877 1570
rect 4821 1516 4823 1568
rect 4823 1516 4875 1568
rect 4875 1516 4877 1568
rect 4821 1514 4877 1516
rect 4609 1350 4665 1352
rect 4609 1298 4611 1350
rect 4611 1298 4663 1350
rect 4663 1298 4665 1350
rect 4609 1296 4665 1298
rect 4821 1350 4877 1352
rect 4821 1298 4823 1350
rect 4823 1298 4875 1350
rect 4875 1298 4877 1350
rect 4821 1296 4877 1298
rect 4927 1108 4983 1110
rect 4927 1056 4929 1108
rect 4929 1056 4981 1108
rect 4981 1056 4983 1108
rect 4927 1054 4983 1056
rect 4927 922 4983 924
rect 4927 870 4929 922
rect 4929 870 4981 922
rect 4981 870 4983 922
rect 4927 868 4983 870
rect -338 515 -282 517
rect -338 463 -336 515
rect -336 463 -284 515
rect -284 463 -282 515
rect -338 461 -282 463
rect -338 329 -282 331
rect -338 277 -336 329
rect -336 277 -284 329
rect -284 277 -282 329
rect -338 275 -282 277
rect 90 472 146 474
rect 90 420 92 472
rect 92 420 144 472
rect 144 420 146 472
rect 90 418 146 420
rect 90 286 146 288
rect 90 234 92 286
rect 92 234 144 286
rect 144 234 146 286
rect 90 232 146 234
rect 539 470 595 472
rect 539 418 541 470
rect 541 418 593 470
rect 593 418 595 470
rect 539 416 595 418
rect 539 284 595 286
rect 539 232 541 284
rect 541 232 593 284
rect 593 232 595 284
rect 539 230 595 232
rect 986 468 1042 470
rect 986 416 988 468
rect 988 416 1040 468
rect 1040 416 1042 468
rect 986 414 1042 416
rect 986 282 1042 284
rect 986 230 988 282
rect 988 230 1040 282
rect 1040 230 1042 282
rect 986 228 1042 230
rect 1759 405 1815 407
rect 1759 353 1761 405
rect 1761 353 1813 405
rect 1813 353 1815 405
rect 1759 351 1815 353
rect 1759 219 1815 221
rect 1759 167 1761 219
rect 1761 167 1813 219
rect 1813 167 1815 219
rect 1759 165 1815 167
rect 2484 405 2540 407
rect 2484 353 2486 405
rect 2486 353 2538 405
rect 2538 353 2540 405
rect 2484 351 2540 353
rect 2484 219 2540 221
rect 2484 167 2486 219
rect 2486 167 2538 219
rect 2538 167 2540 219
rect 2484 165 2540 167
rect 3207 405 3263 407
rect 3207 353 3209 405
rect 3209 353 3261 405
rect 3261 353 3263 405
rect 3207 351 3263 353
rect 3207 219 3263 221
rect 3207 167 3209 219
rect 3209 167 3261 219
rect 3261 167 3263 219
rect 3207 165 3263 167
rect 3960 405 4016 407
rect 3960 353 3962 405
rect 3962 353 4014 405
rect 4014 353 4016 405
rect 3960 351 4016 353
rect 3960 219 4016 221
rect 3960 167 3962 219
rect 3962 167 4014 219
rect 4014 167 4016 219
rect 3960 165 4016 167
rect 4166 405 4222 407
rect 4166 353 4168 405
rect 4168 353 4220 405
rect 4220 353 4222 405
rect 4166 351 4222 353
rect 4166 219 4222 221
rect 4166 167 4168 219
rect 4168 167 4220 219
rect 4220 167 4222 219
rect 4166 165 4222 167
rect 4619 405 4675 407
rect 4619 353 4621 405
rect 4621 353 4673 405
rect 4673 353 4675 405
rect 4619 351 4675 353
rect 4619 219 4675 221
rect 4619 167 4621 219
rect 4621 167 4673 219
rect 4673 167 4675 219
rect 4619 165 4675 167
<< metal3 >>
rect -358 5512 5125 5655
rect -358 5456 -338 5512
rect -282 5493 5125 5512
rect -282 5456 31 5493
rect -358 5437 31 5456
rect 87 5437 527 5493
rect 583 5437 5125 5493
rect -358 5407 5125 5437
rect -358 5351 991 5407
rect 1047 5351 1430 5407
rect 1486 5351 1896 5407
rect 1952 5351 3813 5407
rect 3869 5351 4259 5407
rect 4315 5351 4711 5407
rect 4767 5351 5125 5407
rect -358 5326 5125 5351
rect -358 5270 -338 5326
rect -282 5307 5125 5326
rect -282 5270 31 5307
rect -358 5251 31 5270
rect 87 5251 527 5307
rect 583 5251 5125 5307
rect -358 5221 5125 5251
rect -358 5165 991 5221
rect 1047 5165 1430 5221
rect 1486 5165 1896 5221
rect 1952 5165 3813 5221
rect 3869 5165 4259 5221
rect 4315 5165 4711 5221
rect 4767 5165 5125 5221
rect -358 5127 5125 5165
rect -361 4414 5001 4467
rect -361 4371 993 4414
rect -361 4315 79 4371
rect 135 4315 527 4371
rect 583 4358 993 4371
rect 1049 4396 5001 4414
rect 1049 4371 2482 4396
rect 1049 4358 1430 4371
rect 583 4315 1430 4358
rect 1486 4315 1876 4371
rect 1932 4340 2482 4371
rect 2538 4340 2919 4396
rect 2975 4340 3361 4396
rect 3417 4340 3815 4396
rect 3871 4340 4261 4396
rect 4317 4340 4709 4396
rect 4765 4340 5001 4396
rect 1932 4315 5001 4340
rect -361 4228 5001 4315
rect -361 4185 993 4228
rect -361 4129 79 4185
rect 135 4129 527 4185
rect 583 4172 993 4185
rect 1049 4210 5001 4228
rect 1049 4185 2482 4210
rect 1049 4172 1430 4185
rect 583 4129 1430 4172
rect 1486 4129 1876 4185
rect 1932 4154 2482 4185
rect 2538 4154 2919 4210
rect 2975 4154 3361 4210
rect 3417 4154 3815 4210
rect 3871 4154 4261 4210
rect 4317 4154 4709 4210
rect 4765 4154 5001 4210
rect 1932 4129 5001 4154
rect -361 3964 5001 4129
rect -361 3908 -338 3964
rect -282 3908 5001 3964
rect -361 3881 5001 3908
rect -361 3853 5002 3881
rect -361 3797 4927 3853
rect 4983 3797 5002 3853
rect -361 3778 5002 3797
rect -361 3722 -338 3778
rect -282 3722 5002 3778
rect -361 3667 5002 3722
rect -361 3611 4927 3667
rect 4983 3611 5002 3667
rect -361 3598 5002 3611
rect -361 3542 31 3598
rect 87 3542 1430 3598
rect 1486 3572 5002 3598
rect 1486 3555 5001 3572
rect 1486 3542 2315 3555
rect -361 3499 2315 3542
rect 2371 3537 5001 3555
rect 2371 3499 2794 3537
rect -361 3481 2794 3499
rect 2850 3481 3224 3537
rect 3280 3481 3668 3537
rect 3724 3481 4118 3537
rect 4174 3481 5001 3537
rect -361 3414 5001 3481
rect -361 3412 5002 3414
rect -361 3386 31 3412
rect -361 3330 -338 3386
rect -282 3356 31 3386
rect 87 3356 1430 3412
rect 1486 3386 5002 3412
rect 1486 3369 4927 3386
rect 1486 3356 2315 3369
rect -282 3330 2315 3356
rect -361 3313 2315 3330
rect 2371 3351 4927 3369
rect 2371 3313 2794 3351
rect -361 3295 2794 3313
rect 2850 3295 3224 3351
rect 3280 3295 3668 3351
rect 3724 3295 4118 3351
rect 4174 3330 4927 3351
rect 4983 3330 5002 3386
rect 4174 3295 5002 3330
rect -361 3200 5002 3295
rect -361 3144 -338 3200
rect -282 3144 4927 3200
rect 4983 3144 5002 3200
rect -361 3105 5002 3144
rect 3875 2925 3968 2964
rect 3875 2869 3894 2925
rect 3950 2869 3968 2925
rect 3875 2742 3968 2869
rect 4325 2925 4418 2964
rect 4325 2869 4344 2925
rect 4400 2869 4418 2925
rect 4325 2742 4418 2869
rect 3875 2741 3970 2742
rect 4325 2741 4419 2742
rect 2189 2739 4419 2741
rect 2189 2720 3894 2739
rect 2189 2664 2217 2720
rect 2273 2664 2403 2720
rect 2459 2683 3894 2720
rect 3950 2683 4344 2739
rect 4400 2683 4419 2739
rect 2459 2664 4419 2683
rect 2189 2645 4419 2664
rect -361 2242 5001 2547
rect -361 2214 5002 2242
rect -361 2158 -338 2214
rect -282 2213 4927 2214
rect -282 2158 1432 2213
rect -361 2157 1432 2158
rect 1488 2157 2100 2213
rect 2156 2157 3448 2213
rect 3504 2157 3670 2213
rect 3726 2157 4116 2213
rect 4172 2158 4927 2213
rect 4983 2158 5002 2214
rect 4172 2157 5002 2158
rect -361 2028 5002 2157
rect -361 1972 -338 2028
rect -282 2027 4927 2028
rect -282 1972 1432 2027
rect -361 1971 1432 1972
rect 1488 1971 2100 2027
rect 2156 1971 3448 2027
rect 3504 1971 3670 2027
rect 3726 1971 4116 2027
rect 4172 1972 4927 2027
rect 4983 1972 5002 2028
rect 4172 1971 5002 1972
rect -361 1933 5002 1971
rect -374 1788 5025 1826
rect -374 1732 4609 1788
rect 4665 1732 4821 1788
rect 4877 1732 5025 1788
rect -374 1570 5025 1732
rect -374 1514 110 1570
rect 166 1514 322 1570
rect 378 1514 4609 1570
rect 4665 1514 4821 1570
rect 4877 1514 5025 1570
rect -374 1352 5025 1514
rect -374 1296 110 1352
rect 166 1296 322 1352
rect 378 1296 1981 1352
rect 2037 1296 2191 1352
rect 2247 1296 2402 1352
rect 2458 1296 2613 1352
rect 2669 1296 2824 1352
rect 2880 1296 3035 1352
rect 3091 1296 3246 1352
rect 3302 1296 3457 1352
rect 3513 1296 3668 1352
rect 3724 1296 3879 1352
rect 3935 1296 4089 1352
rect 4145 1296 4609 1352
rect 4665 1296 4821 1352
rect 4877 1296 5025 1352
rect -374 1257 5025 1296
rect -361 1138 5001 1150
rect -361 1112 5002 1138
rect -361 1110 90 1112
rect -361 1054 -338 1110
rect -282 1056 90 1110
rect 146 1056 510 1112
rect 566 1056 982 1112
rect 1038 1056 1838 1112
rect 1894 1056 2499 1112
rect 2555 1056 3222 1112
rect 3278 1056 3947 1112
rect 4003 1056 4171 1112
rect 4227 1110 5002 1112
rect 4227 1056 4927 1110
rect -282 1054 4927 1056
rect 4983 1054 5002 1110
rect -361 926 5002 1054
rect -361 924 90 926
rect -361 868 -338 924
rect -282 870 90 924
rect 146 870 510 926
rect 566 870 982 926
rect 1038 870 1838 926
rect 1894 870 2499 926
rect 2555 870 3222 926
rect 3278 870 3947 926
rect 4003 870 4171 926
rect 4227 924 5002 926
rect 4227 870 4927 924
rect -282 868 4927 870
rect 4983 868 5002 924
rect -361 829 5002 868
rect -361 718 5001 829
rect -361 517 5021 581
rect -361 461 -338 517
rect -282 474 5021 517
rect -282 461 90 474
rect -361 418 90 461
rect 146 472 5021 474
rect 146 418 539 472
rect -361 416 539 418
rect 595 470 5021 472
rect 595 416 986 470
rect -361 414 986 416
rect 1042 414 5021 470
rect -361 407 5021 414
rect -361 351 1759 407
rect 1815 351 2484 407
rect 2540 351 3207 407
rect 3263 351 3960 407
rect 4016 351 4166 407
rect 4222 351 4619 407
rect 4675 351 5021 407
rect -361 331 5021 351
rect -361 275 -338 331
rect -282 288 5021 331
rect -282 275 90 288
rect -361 232 90 275
rect 146 286 5021 288
rect 146 232 539 286
rect -361 230 539 232
rect 595 284 5021 286
rect 595 230 986 284
rect -361 228 986 230
rect 1042 228 5021 284
rect -361 221 5021 228
rect -361 165 1759 221
rect 1815 165 2484 221
rect 2540 165 3207 221
rect 3263 165 3960 221
rect 4016 165 4166 221
rect 4222 165 4619 221
rect 4675 165 5021 221
rect -361 126 5021 165
use M1_NWELL$$44998700_256x8m81  M1_NWELL$$44998700_256x8m81_0
timestamp 1698431365
transform 1 0 -310 0 -1 365
box 0 0 1 1
use M1_NWELL$$44999724_256x8m81  M1_NWELL$$44999724_256x8m81_0
timestamp 1698431365
transform 1 0 4876 0 1 3328
box 0 0 1 1
use M1_NWELL$$45000748_256x8m81  M1_NWELL$$45000748_256x8m81_0
timestamp 1698431365
transform 1 0 -310 0 1 3328
box 0 0 1 1
use M1_PACTIVE4310590878130_256x8m81  M1_PACTIVE4310590878130_256x8m81_0
timestamp 1698431365
transform 1 0 -310 0 1 5375
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_0
timestamp 1698431365
transform 1 0 984 0 1 1313
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_1
timestamp 1698431365
transform 1 0 343 0 1 1313
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_2
timestamp 1698431365
transform 1 0 321 0 1 4049
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_3
timestamp 1698431365
transform 1 0 758 0 1 4865
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_0
timestamp 1698431365
transform 1 0 2110 0 1 4502
box 0 0 1 1
use M1_POLY2$$45109292_256x8m81  M1_POLY2$$45109292_256x8m81_0
timestamp 1698431365
transform 1 0 2962 0 1 4765
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_0
timestamp 1698431365
transform 1 0 3610 0 1 2609
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_1
timestamp 1698431365
transform 1 0 2607 0 1 712
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_2
timestamp 1698431365
transform 1 0 2838 0 1 712
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_3
timestamp 1698431365
transform 1 0 3331 0 1 712
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_4
timestamp 1698431365
transform 1 0 3537 0 1 712
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_5
timestamp 1698431365
transform 1 0 4230 0 1 671
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_6
timestamp 1698431365
transform 1 0 3355 0 1 2426
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_7
timestamp 1698431365
transform 1 0 1882 0 1 773
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_8
timestamp 1698431365
transform 1 0 2071 0 1 773
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_9
timestamp 1698431365
transform 1 0 1347 0 1 714
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_10
timestamp 1698431365
transform 1 0 2240 0 1 2410
box 0 0 1 1
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_0
timestamp 1698431365
transform 1 0 2885 0 1 3765
box 0 0 1 1
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_1
timestamp 1698431365
transform 1 0 2388 0 1 2667
box 0 0 1 1
use M1_PSUB$$44997676_256x8m81  M1_PSUB$$44997676_256x8m81_0
timestamp 1698431365
transform 1 0 4797 0 -1 2086
box 0 0 1 1
use M1_PSUB$$44997676_256x8m81  M1_PSUB$$44997676_256x8m81_1
timestamp 1698431365
transform 1 0 -152 0 -1 2086
box 0 0 1 1
use M1_PSUB$$45110316_285_256x8m81  M1_PSUB$$45110316_285_256x8m81_0
timestamp 1698431365
transform 1 0 4876 0 -1 1065
box 0 0 1 1
use M1_PSUB$$45110316_285_256x8m81  M1_PSUB$$45110316_285_256x8m81_1
timestamp 1698431365
transform 1 0 -310 0 -1 1065
box 0 0 1 1
use M2_M1$$43374636_256x8m81  M2_M1$$43374636_256x8m81_0
timestamp 1698431365
transform 1 0 244 0 1 1433
box 0 0 1 1
use M2_M1$$45002796_256x8m81  M2_M1$$45002796_256x8m81_0
timestamp 1698431365
transform 1 0 3063 0 1 1324
box 0 0 1 1
use M2_M1$$45003820_256x8m81  M2_M1$$45003820_256x8m81_0
timestamp 1698431365
transform 1 0 4743 0 1 1542
box 0 0 1 1
use M2_M1c$$203396140_256x8m81  M2_M1c$$203396140_256x8m81_0
timestamp 1698431365
transform 1 0 997 0 1 3974
box 0 0 1 1
use M3_M2$$45005868_256x8m81  M3_M2$$45005868_256x8m81_0
timestamp 1698431365
transform 1 0 3063 0 1 1324
box 0 0 1 1
use M3_M2$$45006892_256x8m81  M3_M2$$45006892_256x8m81_0
timestamp 1698431365
transform 1 0 4743 0 1 1542
box 0 0 1 1
use M3_M2$$45008940_256x8m81  M3_M2$$45008940_256x8m81_0
timestamp 1698431365
transform 1 0 244 0 1 1433
box 0 0 1 1
use nmos_1p2$$45100076_256x8m81  nmos_1p2$$45100076_256x8m81_0
timestamp 1698431365
transform -1 0 4063 0 -1 2301
box -31 0 -30 1
use nmos_1p2$$45101100_256x8m81  nmos_1p2$$45101100_256x8m81_0
timestamp 1698431365
transform 1 0 202 0 1 855
box -31 0 -30 1
use nmos_1p2$$45102124_256x8m81  nmos_1p2$$45102124_256x8m81_0
timestamp 1698431365
transform -1 0 1823 0 -1 2301
box -31 0 -30 1
use nmos_1p2$$45103148_256x8m81  nmos_1p2$$45103148_256x8m81_0
timestamp 1698431365
transform -1 0 3391 0 -1 2301
box -31 0 -30 1
use nmos_5p04310590878112_256x8m81  nmos_5p04310590878112_256x8m81_0
timestamp 1698431365
transform -1 0 4684 0 1 5006
box 0 0 1 1
use nmos_5p04310590878123_256x8m81  nmos_5p04310590878123_256x8m81_0
timestamp 1698431365
transform 1 0 3065 0 1 884
box 0 0 1 1
use nmos_5p04310590878123_256x8m81  nmos_5p04310590878123_256x8m81_1
timestamp 1698431365
transform 1 0 1616 0 1 884
box 0 0 1 1
use nmos_5p04310590878123_256x8m81  nmos_5p04310590878123_256x8m81_2
timestamp 1698431365
transform 1 0 2341 0 1 884
box 0 0 1 1
use nmos_5p04310590878126_256x8m81  nmos_5p04310590878126_256x8m81_0
timestamp 1698431365
transform 1 0 1074 0 1 5006
box 0 0 1 1
use nmos_5p04310590878126_256x8m81  nmos_5p04310590878126_256x8m81_1
timestamp 1698431365
transform 1 0 2483 0 1 5006
box 0 0 1 1
use nmos_5p04310590878131_256x8m81  nmos_5p04310590878131_256x8m81_0
timestamp 1698431365
transform -1 0 503 0 1 5223
box 0 0 1 1
use nmos_5p04310590878132_256x8m81  nmos_5p04310590878132_256x8m81_0
timestamp 1698431365
transform 1 0 3790 0 1 884
box 0 0 1 1
use nmos_5p04310590878133_256x8m81  nmos_5p04310590878133_256x8m81_0
timestamp 1698431365
transform 1 0 4251 0 1 818
box 0 0 1 1
use pmos_1p2$$45095980_256x8m81  pmos_1p2$$45095980_256x8m81_0
timestamp 1698431365
transform -1 0 4653 0 1 4090
box -31 0 -30 1
use pmos_1p2$$46281772_256x8m81  pmos_1p2$$46281772_256x8m81_0
timestamp 1698431365
transform -1 0 4287 0 -1 3650
box -31 0 -30 1
use pmos_1p2$$46281772_256x8m81  pmos_1p2$$46281772_256x8m81_1
timestamp 1698431365
transform -1 0 3391 0 -1 3650
box -31 0 -30 1
use pmos_1p2$$46282796_256x8m81  pmos_1p2$$46282796_256x8m81_0
timestamp 1698431365
transform 1 0 202 0 1 118
box -31 0 -30 1
use pmos_1p2$$46283820_256x8m81  pmos_1p2$$46283820_256x8m81_0
timestamp 1698431365
transform -1 0 2271 0 -1 3629
box -31 0 -30 1
use pmos_1p2$$46284844_256x8m81  pmos_1p2$$46284844_256x8m81_0
timestamp 1698431365
transform 1 0 4282 0 1 197
box -31 0 -30 1
use pmos_1p2$$46285868_256x8m81  pmos_1p2$$46285868_256x8m81_0
timestamp 1698431365
transform 1 0 1777 0 1 4198
box -31 0 -30 1
use pmos_1p2$$46286892_256x8m81  pmos_1p2$$46286892_256x8m81_0
timestamp 1698431365
transform 1 0 1105 0 1 4198
box -31 0 -30 1
use pmos_1p2$$46287916_256x8m81  pmos_1p2$$46287916_256x8m81_0
timestamp 1698431365
transform -1 0 472 0 1 4189
box -31 0 -30 1
use pmos_5p04310590878125_256x8m81  pmos_5p04310590878125_256x8m81_0
timestamp 1698431365
transform 1 0 3065 0 1 296
box 0 0 1 1
use pmos_5p04310590878125_256x8m81  pmos_5p04310590878125_256x8m81_1
timestamp 1698431365
transform 1 0 1616 0 1 296
box 0 0 1 1
use pmos_5p04310590878125_256x8m81  pmos_5p04310590878125_256x8m81_2
timestamp 1698431365
transform 1 0 2341 0 1 296
box 0 0 1 1
use pmos_5p04310590878138_256x8m81  pmos_5p04310590878138_256x8m81_0
timestamp 1698431365
transform 1 0 3790 0 1 334
box 0 0 1 1
use po_m1_256x8m81  po_m1_256x8m81_0
timestamp 1698431365
transform 1 0 2743 0 1 1440
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_0
timestamp 1698431365
transform -1 0 3744 0 -1 2251
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_1
timestamp 1698431365
transform 1 0 3189 0 1 127
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_2
timestamp 1698431365
transform 1 0 2466 0 1 127
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_3
timestamp 1698431365
transform -1 0 3522 0 -1 2251
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_4
timestamp 1698431365
transform 1 0 4909 0 1 830
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_5
timestamp 1698431365
transform 1 0 4909 0 1 1934
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_6
timestamp 1698431365
transform 1 0 4601 0 1 127
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_7
timestamp 1698431365
transform 1 0 4148 0 1 127
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_8
timestamp 1698431365
transform 1 0 3942 0 1 127
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_9
timestamp 1698431365
transform -1 0 4190 0 -1 2251
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_10
timestamp 1698431365
transform 1 0 72 0 1 194
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_11
timestamp 1698431365
transform -1 0 -264 0 -1 555
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_12
timestamp 1698431365
transform -1 0 1506 0 -1 2251
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_13
timestamp 1698431365
transform 1 0 -356 0 1 830
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_14
timestamp 1698431365
transform 1 0 -356 0 1 1934
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_15
timestamp 1698431365
transform 1 0 1741 0 1 127
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_16
timestamp 1698431365
transform 1 0 968 0 1 190
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_17
timestamp 1698431365
transform 1 0 521 0 1 192
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_18
timestamp 1698431365
transform -1 0 2174 0 -1 2251
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_19
timestamp 1698431365
transform -1 0 1950 0 -1 4409
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_20
timestamp 1698431365
transform 1 0 -356 0 1 3106
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_21
timestamp 1698431365
transform -1 0 -264 0 -1 5550
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_22
timestamp 1698431365
transform -1 0 105 0 -1 5531
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_23
timestamp 1698431365
transform -1 0 153 0 -1 4409
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_24
timestamp 1698431365
transform -1 0 1065 0 -1 5445
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_25
timestamp 1698431365
transform -1 0 1504 0 -1 5445
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_26
timestamp 1698431365
transform -1 0 1970 0 -1 5445
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_27
timestamp 1698431365
transform -1 0 601 0 -1 5531
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_28
timestamp 1698431365
transform -1 0 601 0 -1 4409
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_29
timestamp 1698431365
transform -1 0 1067 0 -1 4452
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_30
timestamp 1698431365
transform -1 0 1504 0 -1 4409
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_31
timestamp 1698431365
transform -1 0 105 0 -1 3636
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_32
timestamp 1698431365
transform -1 0 1504 0 -1 3636
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_33
timestamp 1698431365
transform 1 0 -356 0 1 3684
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_34
timestamp 1698431365
transform 1 0 4909 0 1 3106
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_35
timestamp 1698431365
transform 1 0 4909 0 1 3573
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_36
timestamp 1698431365
transform -1 0 3742 0 -1 3575
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_37
timestamp 1698431365
transform -1 0 4192 0 -1 3575
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_38
timestamp 1698431365
transform -1 0 3298 0 -1 3575
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_39
timestamp 1698431365
transform -1 0 2868 0 -1 3575
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_40
timestamp 1698431365
transform -1 0 2556 0 -1 4434
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_41
timestamp 1698431365
transform -1 0 2993 0 -1 4434
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_42
timestamp 1698431365
transform -1 0 3435 0 -1 4434
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_43
timestamp 1698431365
transform -1 0 3889 0 -1 4434
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_44
timestamp 1698431365
transform -1 0 4335 0 -1 4434
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_45
timestamp 1698431365
transform -1 0 4783 0 -1 4434
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_46
timestamp 1698431365
transform -1 0 3887 0 -1 5445
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_47
timestamp 1698431365
transform -1 0 4333 0 -1 5445
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_48
timestamp 1698431365
transform -1 0 4785 0 -1 5445
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_49
timestamp 1698431365
transform -1 0 4418 0 -1 2963
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_50
timestamp 1698431365
transform -1 0 3968 0 -1 2963
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_51
timestamp 1698431365
transform -1 0 2389 0 -1 3593
box 0 0 1 1
use via1_R90_256x8m81  via1_R90_256x8m81_0
timestamp 1698431365
transform 0 -1 2422 1 0 2646
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_0
timestamp 1698431365
transform 1 0 4377 0 1 775
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_1
timestamp 1698431365
transform 1 0 2481 0 1 843
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_2
timestamp 1698431365
transform 1 0 3204 0 1 843
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_3
timestamp 1698431365
transform 1 0 3929 0 1 843
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_4
timestamp 1698431365
transform 1 0 4153 0 1 843
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_5
timestamp 1698431365
transform 1 0 1504 0 1 508
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_6
timestamp 1698431365
transform 1 0 1820 0 1 843
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_7
timestamp 1698431365
transform 1 0 72 0 1 843
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_8
timestamp 1698431365
transform 1 0 492 0 1 843
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_9
timestamp 1698431365
transform 1 0 964 0 1 843
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_10
timestamp 1698431365
transform -1 0 2145 0 -1 4616
box 0 0 1 1
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_0
timestamp 1698431365
transform 0 -1 4469 1 0 1512
box 0 0 1 1
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_1
timestamp 1698431365
transform 0 -1 4287 1 0 621
box 0 0 1 1
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_2
timestamp 1698431365
transform 0 -1 1168 1 0 1512
box 0 0 1 1
use via1_x2_R270_256x8m81  via1_x2_R270_256x8m81_0
timestamp 1698431365
transform 0 1 3083 -1 0 2471
box 0 0 1 1
use via1_x2_R270_256x8m81  via1_x2_R270_256x8m81_1
timestamp 1698431365
transform 0 1 1421 -1 0 1154
box 0 0 1 1
use via1_x2_R270_256x8m81  via1_x2_R270_256x8m81_2
timestamp 1698431365
transform 0 1 2778 -1 0 3818
box 0 0 1 1
use via1_x2_R270_256x8m81  via1_x2_R270_256x8m81_3
timestamp 1698431365
transform 0 1 2181 -1 0 2471
box 0 0 1 1
use via1_x2_R270_256x8m81  via1_x2_R270_256x8m81_4
timestamp 1698431365
transform 0 1 2275 -1 0 4833
box 0 0 1 1
use via2_x2_256x8m81  via2_x2_256x8m81_0
timestamp 1698431365
transform 1 0 3204 0 1 832
box 0 0 1 1
use via2_x2_256x8m81  via2_x2_256x8m81_1
timestamp 1698431365
transform 1 0 2481 0 1 832
box 0 0 1 1
use via2_x2_256x8m81  via2_x2_256x8m81_2
timestamp 1698431365
transform 1 0 3929 0 1 832
box 0 0 1 1
use via2_x2_256x8m81  via2_x2_256x8m81_3
timestamp 1698431365
transform 1 0 4153 0 1 832
box 0 0 1 1
use via2_x2_256x8m81  via2_x2_256x8m81_4
timestamp 1698431365
transform 1 0 964 0 1 832
box 0 0 1 1
use via2_x2_256x8m81  via2_x2_256x8m81_5
timestamp 1698431365
transform 1 0 492 0 1 832
box 0 0 1 1
use via2_x2_256x8m81  via2_x2_256x8m81_6
timestamp 1698431365
transform 1 0 72 0 1 832
box 0 0 1 1
use via2_x2_256x8m81  via2_x2_256x8m81_7
timestamp 1698431365
transform 1 0 1820 0 1 832
box 0 0 1 1
use via2_x2_R90_256x8m81  via2_x2_R90_256x8m81_0
timestamp 1698431365
transform 0 -1 2497 1 0 2646
box 0 0 1 1
<< labels >>
rlabel metal1 s 1456 2584 1456 2584 4 pcb
port 1 nsew
rlabel metal1 s 4066 5565 4066 5565 4 se
port 2 nsew
rlabel metal3 s 2398 3802 2398 3802 4 vdd
port 3 nsew
rlabel metal3 s 2163 5443 2163 5443 4 vss
port 4 nsew
rlabel metal3 s 2288 1061 2288 1061 4 vss
port 4 nsew
rlabel metal3 s 248 1437 248 1437 4 men
port 5 nsew
rlabel metal3 s 2288 2151 2288 2151 4 vss
port 4 nsew
rlabel metal3 s 1489 379 1489 379 4 vdd
port 3 nsew
<< properties >>
string GDS_END 495280
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 476310
string path 20.320 27.120 20.320 27.785 22.565 27.785 22.565 26.905 
<< end >>
