magic
tech gf180mcuB
timestamp 1698855177
<< properties >>
string gencell npn_00p54x10p00_0
string library gf180mcu
string parameter m=1
<< end >>
