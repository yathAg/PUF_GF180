magic
tech gf180mcuA
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 453 3558 1094
<< pwell >>
rect -86 -86 3558 453
<< mvnmos >>
rect 124 69 244 333
rect 308 69 428 333
rect 532 69 652 333
rect 716 69 836 333
rect 940 69 1060 333
rect 1124 69 1244 333
rect 1348 69 1468 333
rect 1542 69 1662 333
rect 1746 69 1866 333
rect 1940 69 2060 333
rect 2164 69 2284 333
rect 2348 69 2468 333
rect 2572 69 2692 333
rect 2756 69 2876 333
rect 2980 69 3100 333
rect 3164 69 3284 333
<< mvpmos >>
rect 124 683 224 939
rect 328 683 428 939
rect 532 683 632 939
rect 736 683 836 939
rect 940 683 1040 939
rect 1144 683 1244 939
rect 1348 683 1448 939
rect 1552 683 1652 939
rect 1756 683 1856 939
rect 1960 683 2060 939
rect 2164 683 2264 939
rect 2368 683 2468 939
rect 2572 683 2672 939
rect 2776 683 2876 939
rect 2980 683 3080 939
rect 3184 683 3284 939
<< mvndiff >>
rect 36 287 124 333
rect 36 147 49 287
rect 95 147 124 287
rect 36 69 124 147
rect 244 69 308 333
rect 428 193 532 333
rect 428 147 457 193
rect 503 147 532 193
rect 428 69 532 147
rect 652 69 716 333
rect 836 287 940 333
rect 836 147 865 287
rect 911 147 940 287
rect 836 69 940 147
rect 1060 69 1124 333
rect 1244 193 1348 333
rect 1244 147 1273 193
rect 1319 147 1348 193
rect 1244 69 1348 147
rect 1468 69 1542 333
rect 1662 69 1746 333
rect 1866 69 1940 333
rect 2060 285 2164 333
rect 2060 239 2089 285
rect 2135 239 2164 285
rect 2060 69 2164 239
rect 2284 69 2348 333
rect 2468 193 2572 333
rect 2468 147 2497 193
rect 2543 147 2572 193
rect 2468 69 2572 147
rect 2692 69 2756 333
rect 2876 285 2980 333
rect 2876 239 2905 285
rect 2951 239 2980 285
rect 2876 69 2980 239
rect 3100 69 3164 333
rect 3284 193 3372 333
rect 3284 147 3313 193
rect 3359 147 3372 193
rect 3284 69 3372 147
<< mvpdiff >>
rect 36 881 124 939
rect 36 741 49 881
rect 95 741 124 881
rect 36 683 124 741
rect 224 861 328 939
rect 224 721 253 861
rect 299 721 328 861
rect 224 683 328 721
rect 428 881 532 939
rect 428 741 457 881
rect 503 741 532 881
rect 428 683 532 741
rect 632 861 736 939
rect 632 721 661 861
rect 707 721 736 861
rect 632 683 736 721
rect 836 881 940 939
rect 836 741 865 881
rect 911 741 940 881
rect 836 683 940 741
rect 1040 861 1144 939
rect 1040 721 1069 861
rect 1115 721 1144 861
rect 1040 683 1144 721
rect 1244 881 1348 939
rect 1244 741 1273 881
rect 1319 741 1348 881
rect 1244 683 1348 741
rect 1448 861 1552 939
rect 1448 721 1477 861
rect 1523 721 1552 861
rect 1448 683 1552 721
rect 1652 881 1756 939
rect 1652 741 1681 881
rect 1727 741 1756 881
rect 1652 683 1756 741
rect 1856 861 1960 939
rect 1856 721 1885 861
rect 1931 721 1960 861
rect 1856 683 1960 721
rect 2060 881 2164 939
rect 2060 741 2089 881
rect 2135 741 2164 881
rect 2060 683 2164 741
rect 2264 861 2368 939
rect 2264 721 2293 861
rect 2339 721 2368 861
rect 2264 683 2368 721
rect 2468 881 2572 939
rect 2468 741 2497 881
rect 2543 741 2572 881
rect 2468 683 2572 741
rect 2672 861 2776 939
rect 2672 721 2701 861
rect 2747 721 2776 861
rect 2672 683 2776 721
rect 2876 881 2980 939
rect 2876 741 2905 881
rect 2951 741 2980 881
rect 2876 683 2980 741
rect 3080 861 3184 939
rect 3080 721 3109 861
rect 3155 721 3184 861
rect 3080 683 3184 721
rect 3284 881 3372 939
rect 3284 741 3313 881
rect 3359 741 3372 881
rect 3284 683 3372 741
<< mvndiffc >>
rect 49 147 95 287
rect 457 147 503 193
rect 865 147 911 287
rect 1273 147 1319 193
rect 2089 239 2135 285
rect 2497 147 2543 193
rect 2905 239 2951 285
rect 3313 147 3359 193
<< mvpdiffc >>
rect 49 741 95 881
rect 253 721 299 861
rect 457 741 503 881
rect 661 721 707 861
rect 865 741 911 881
rect 1069 721 1115 861
rect 1273 741 1319 881
rect 1477 721 1523 861
rect 1681 741 1727 881
rect 1885 721 1931 861
rect 2089 741 2135 881
rect 2293 721 2339 861
rect 2497 741 2543 881
rect 2701 721 2747 861
rect 2905 741 2951 881
rect 3109 721 3155 861
rect 3313 741 3359 881
<< polysilicon >>
rect 124 939 224 983
rect 328 939 428 983
rect 532 939 632 983
rect 736 939 836 983
rect 940 939 1040 983
rect 1144 939 1244 983
rect 1348 939 1448 983
rect 1552 939 1652 983
rect 1756 939 1856 983
rect 1960 939 2060 983
rect 2164 939 2264 983
rect 2368 939 2468 983
rect 2572 939 2672 983
rect 2776 939 2876 983
rect 2980 939 3080 983
rect 3184 939 3284 983
rect 124 500 224 683
rect 124 454 153 500
rect 199 454 224 500
rect 124 377 224 454
rect 328 513 428 683
rect 532 513 632 683
rect 328 500 632 513
rect 328 454 377 500
rect 423 454 632 500
rect 328 441 632 454
rect 328 377 428 441
rect 124 333 244 377
rect 308 333 428 377
rect 532 377 632 441
rect 736 513 836 683
rect 940 513 1040 683
rect 736 500 1040 513
rect 736 454 749 500
rect 795 454 1040 500
rect 736 441 1040 454
rect 736 377 836 441
rect 532 333 652 377
rect 716 333 836 377
rect 940 377 1040 441
rect 1144 513 1244 683
rect 1348 513 1448 683
rect 1144 500 1448 513
rect 1144 454 1157 500
rect 1203 454 1448 500
rect 1144 441 1448 454
rect 1144 377 1244 441
rect 940 333 1060 377
rect 1124 333 1244 377
rect 1348 377 1448 441
rect 1552 500 1652 683
rect 1552 454 1565 500
rect 1611 454 1652 500
rect 1552 377 1652 454
rect 1756 500 1856 683
rect 1756 454 1797 500
rect 1843 454 1856 500
rect 1756 377 1856 454
rect 1960 513 2060 683
rect 2164 513 2264 683
rect 1960 500 2264 513
rect 1960 454 1973 500
rect 2019 454 2264 500
rect 1960 441 2264 454
rect 1960 377 2060 441
rect 1348 333 1468 377
rect 1542 333 1662 377
rect 1746 333 1866 377
rect 1940 333 2060 377
rect 2164 377 2264 441
rect 2368 513 2468 683
rect 2572 513 2672 683
rect 2368 500 2672 513
rect 2368 454 2381 500
rect 2427 454 2672 500
rect 2368 441 2672 454
rect 2368 377 2468 441
rect 2164 333 2284 377
rect 2348 333 2468 377
rect 2572 377 2672 441
rect 2776 513 2876 683
rect 2980 513 3080 683
rect 3184 513 3284 683
rect 2776 500 3080 513
rect 2776 454 2789 500
rect 2835 454 3080 500
rect 2776 441 3080 454
rect 3128 500 3284 513
rect 3128 454 3141 500
rect 3187 454 3284 500
rect 3128 441 3284 454
rect 2776 377 2876 441
rect 2572 333 2692 377
rect 2756 333 2876 377
rect 2980 377 3080 441
rect 2980 333 3100 377
rect 3164 333 3284 441
rect 124 25 244 69
rect 308 25 428 69
rect 532 25 652 69
rect 716 25 836 69
rect 940 25 1060 69
rect 1124 25 1244 69
rect 1348 25 1468 69
rect 1542 25 1662 69
rect 1746 25 1866 69
rect 1940 25 2060 69
rect 2164 25 2284 69
rect 2348 25 2468 69
rect 2572 25 2692 69
rect 2756 25 2876 69
rect 2980 25 3100 69
rect 3164 25 3284 69
<< polycontact >>
rect 153 454 199 500
rect 377 454 423 500
rect 749 454 795 500
rect 1157 454 1203 500
rect 1565 454 1611 500
rect 1797 454 1843 500
rect 1973 454 2019 500
rect 2381 454 2427 500
rect 2789 454 2835 500
rect 3141 454 3187 500
<< metal1 >>
rect 0 918 3472 1098
rect 49 881 95 918
rect 457 881 503 918
rect 49 730 95 741
rect 253 861 299 872
rect 865 881 911 918
rect 457 730 503 741
rect 578 861 707 872
rect 253 684 299 721
rect 578 721 661 861
rect 1273 881 1319 918
rect 865 730 911 741
rect 1069 861 1115 872
rect 578 684 707 721
rect 1681 881 1727 918
rect 1273 730 1319 741
rect 1477 861 1523 872
rect 1069 684 1115 721
rect 2089 881 2135 918
rect 1681 730 1727 741
rect 1885 861 1931 872
rect 1477 684 1523 721
rect 2497 881 2543 918
rect 2089 730 2135 741
rect 2293 861 2339 872
rect 1885 684 1931 721
rect 2905 881 2951 918
rect 2497 730 2543 741
rect 2701 861 2747 872
rect 2293 684 2339 721
rect 3313 881 3359 918
rect 2905 730 2951 741
rect 3109 861 3155 872
rect 2701 684 2747 721
rect 3313 730 3359 741
rect 3109 684 3155 721
rect 253 638 3279 684
rect 142 546 1306 592
rect 142 500 210 546
rect 749 500 795 546
rect 1260 500 1306 546
rect 1786 546 3187 592
rect 1786 500 1854 546
rect 2270 500 2427 546
rect 3141 500 3187 546
rect 142 454 153 500
rect 199 454 210 500
rect 366 454 377 500
rect 423 454 434 500
rect 366 397 434 454
rect 749 443 795 454
rect 841 454 1157 500
rect 1203 454 1214 500
rect 1260 454 1565 500
rect 1611 454 1622 500
rect 1786 454 1797 500
rect 1843 454 1854 500
rect 1934 454 1973 500
rect 2019 454 2030 500
rect 841 397 887 454
rect 366 351 887 397
rect 1934 397 2030 454
rect 2270 454 2381 500
rect 2270 443 2427 454
rect 2473 454 2789 500
rect 2835 454 2846 500
rect 2473 397 2519 454
rect 3141 443 3187 454
rect 1934 351 2519 397
rect 49 287 2032 298
rect 95 252 865 287
rect 49 136 95 147
rect 457 193 503 204
rect 457 90 503 147
rect 911 252 2032 287
rect 3233 285 3279 638
rect 865 136 911 147
rect 1273 193 1319 204
rect 1986 193 2032 252
rect 2078 239 2089 285
rect 2135 239 2905 285
rect 2951 239 3279 285
rect 1986 147 2497 193
rect 2543 147 3313 193
rect 3359 147 3370 193
rect 1273 90 1319 147
rect 0 -90 3472 90
<< labels >>
flabel metal1 s 2473 454 2846 500 0 FreeSans 200 0 0 0 A1
port 1 nsew default input
flabel metal1 s 1786 546 3187 592 0 FreeSans 200 0 0 0 A2
port 2 nsew default input
flabel metal1 s 142 546 1306 592 0 FreeSans 200 0 0 0 A3
port 3 nsew default input
flabel metal1 s 841 454 1214 500 0 FreeSans 200 0 0 0 A4
port 4 nsew default input
flabel metal1 s 0 918 3472 1098 0 FreeSans 200 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 1273 90 1319 204 0 FreeSans 200 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel metal1 s 3109 684 3155 872 0 FreeSans 200 0 0 0 ZN
port 5 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 7 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 8 nsew ground bidirectional
rlabel metal1 s 1934 454 2030 500 1 A1
port 1 nsew default input
rlabel metal1 s 2473 397 2519 454 1 A1
port 1 nsew default input
rlabel metal1 s 1934 397 2030 454 1 A1
port 1 nsew default input
rlabel metal1 s 1934 351 2519 397 1 A1
port 1 nsew default input
rlabel metal1 s 3141 454 3187 546 1 A2
port 2 nsew default input
rlabel metal1 s 2270 454 2427 546 1 A2
port 2 nsew default input
rlabel metal1 s 1786 454 1854 546 1 A2
port 2 nsew default input
rlabel metal1 s 3141 443 3187 454 1 A2
port 2 nsew default input
rlabel metal1 s 2270 443 2427 454 1 A2
port 2 nsew default input
rlabel metal1 s 1260 500 1306 546 1 A3
port 3 nsew default input
rlabel metal1 s 749 500 795 546 1 A3
port 3 nsew default input
rlabel metal1 s 142 500 210 546 1 A3
port 3 nsew default input
rlabel metal1 s 1260 454 1622 500 1 A3
port 3 nsew default input
rlabel metal1 s 749 454 795 500 1 A3
port 3 nsew default input
rlabel metal1 s 142 454 210 500 1 A3
port 3 nsew default input
rlabel metal1 s 749 443 795 454 1 A3
port 3 nsew default input
rlabel metal1 s 366 454 434 500 1 A4
port 4 nsew default input
rlabel metal1 s 841 397 887 454 1 A4
port 4 nsew default input
rlabel metal1 s 366 397 434 454 1 A4
port 4 nsew default input
rlabel metal1 s 366 351 887 397 1 A4
port 4 nsew default input
rlabel metal1 s 2701 684 2747 872 1 ZN
port 5 nsew default output
rlabel metal1 s 2293 684 2339 872 1 ZN
port 5 nsew default output
rlabel metal1 s 1885 684 1931 872 1 ZN
port 5 nsew default output
rlabel metal1 s 1477 684 1523 872 1 ZN
port 5 nsew default output
rlabel metal1 s 1069 684 1115 872 1 ZN
port 5 nsew default output
rlabel metal1 s 578 684 707 872 1 ZN
port 5 nsew default output
rlabel metal1 s 253 684 299 872 1 ZN
port 5 nsew default output
rlabel metal1 s 253 638 3279 684 1 ZN
port 5 nsew default output
rlabel metal1 s 3233 285 3279 638 1 ZN
port 5 nsew default output
rlabel metal1 s 2078 239 3279 285 1 ZN
port 5 nsew default output
rlabel metal1 s 3313 730 3359 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2905 730 2951 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2497 730 2543 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2089 730 2135 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1681 730 1727 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1273 730 1319 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 865 730 911 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 457 730 503 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 49 730 95 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 457 90 503 204 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 3472 90 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3472 1008
string GDS_END 74330
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 66618
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
