magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 352 1654 870
<< pwell >>
rect -86 -86 1654 352
<< metal1 >>
rect 0 724 1568 844
rect 49 646 95 724
rect 477 632 523 724
rect 74 348 430 430
rect 757 536 803 678
rect 961 610 1007 724
rect 1185 536 1231 678
rect 1409 552 1455 724
rect 757 472 1231 536
rect 1026 289 1102 472
rect 38 60 106 208
rect 757 243 1251 289
rect 522 60 590 197
rect 757 138 803 243
rect 970 60 1038 197
rect 1205 138 1251 243
rect 1418 60 1486 197
rect 0 -60 1568 60
<< obsm1 >>
rect 253 552 299 676
rect 253 506 635 552
rect 589 405 635 506
rect 589 337 966 405
rect 589 300 635 337
rect 273 254 635 300
rect 1153 337 1387 405
rect 273 148 319 254
<< labels >>
rlabel metal1 s 74 348 430 430 6 I
port 1 nsew default input
rlabel metal1 s 1205 138 1251 243 6 Z
port 2 nsew default output
rlabel metal1 s 757 138 803 243 6 Z
port 2 nsew default output
rlabel metal1 s 757 243 1251 289 6 Z
port 2 nsew default output
rlabel metal1 s 1026 289 1102 472 6 Z
port 2 nsew default output
rlabel metal1 s 757 472 1231 536 6 Z
port 2 nsew default output
rlabel metal1 s 1185 536 1231 678 6 Z
port 2 nsew default output
rlabel metal1 s 757 536 803 678 6 Z
port 2 nsew default output
rlabel metal1 s 1409 552 1455 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 961 610 1007 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 477 632 523 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 646 95 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 724 1568 844 6 VDD
port 3 nsew power bidirectional abutment
rlabel nwell s -86 352 1654 870 6 VNW
port 4 nsew power bidirectional
rlabel pwell s -86 -86 1654 352 6 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 0 -60 1568 60 8 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1418 60 1486 197 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 970 60 1038 197 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 522 60 590 197 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 38 60 106 208 6 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1568 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 773314
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 768974
<< end >>
