magic
tech gf180mcuB
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 453 2886 1094
<< pwell >>
rect -86 -86 2886 453
<< mvnmos >>
rect 131 69 251 333
rect 315 69 435 333
rect 539 69 659 333
rect 723 69 843 333
rect 1071 69 1191 333
rect 1275 69 1395 333
rect 1499 69 1619 333
rect 1683 69 1803 333
rect 1910 69 2030 333
rect 2094 69 2214 333
rect 2318 69 2438 333
rect 2502 69 2622 333
<< mvpmos >>
rect 131 573 231 939
rect 335 573 435 939
rect 539 573 639 939
rect 743 573 843 939
rect 1091 573 1191 939
rect 1295 573 1395 939
rect 1499 573 1599 939
rect 1703 573 1803 939
rect 1910 573 2010 939
rect 2114 573 2214 939
rect 2318 573 2418 939
rect 2522 573 2622 939
<< mvndiff >>
rect 43 287 131 333
rect 43 147 56 287
rect 102 147 131 287
rect 43 69 131 147
rect 251 69 315 333
rect 435 128 539 333
rect 435 82 464 128
rect 510 82 539 128
rect 435 69 539 82
rect 659 69 723 333
rect 843 287 1071 333
rect 843 147 996 287
rect 1042 147 1071 287
rect 843 69 1071 147
rect 1191 69 1275 333
rect 1395 128 1499 333
rect 1395 82 1424 128
rect 1470 82 1499 128
rect 1395 69 1499 82
rect 1619 69 1683 333
rect 1803 320 1910 333
rect 1803 180 1832 320
rect 1878 180 1910 320
rect 1803 69 1910 180
rect 2030 69 2094 333
rect 2214 128 2318 333
rect 2214 82 2243 128
rect 2289 82 2318 128
rect 2214 69 2318 82
rect 2438 69 2502 333
rect 2622 320 2710 333
rect 2622 180 2651 320
rect 2697 180 2710 320
rect 2622 69 2710 180
<< mvpdiff >>
rect 43 926 131 939
rect 43 786 56 926
rect 102 786 131 926
rect 43 573 131 786
rect 231 726 335 939
rect 231 586 260 726
rect 306 586 335 726
rect 231 573 335 586
rect 435 926 539 939
rect 435 786 464 926
rect 510 786 539 926
rect 435 573 539 786
rect 639 726 743 939
rect 639 586 668 726
rect 714 586 743 726
rect 639 573 743 586
rect 843 926 931 939
rect 843 786 872 926
rect 918 786 931 926
rect 843 573 931 786
rect 1003 818 1091 939
rect 1003 678 1016 818
rect 1062 678 1091 818
rect 1003 573 1091 678
rect 1191 726 1295 939
rect 1191 586 1220 726
rect 1266 586 1295 726
rect 1191 573 1295 586
rect 1395 818 1499 939
rect 1395 678 1424 818
rect 1470 678 1499 818
rect 1395 573 1499 678
rect 1599 726 1703 939
rect 1599 586 1628 726
rect 1674 586 1703 726
rect 1599 573 1703 586
rect 1803 818 1910 939
rect 1803 678 1832 818
rect 1878 678 1910 818
rect 1803 573 1910 678
rect 2010 726 2114 939
rect 2010 586 2039 726
rect 2085 586 2114 726
rect 2010 573 2114 586
rect 2214 818 2318 939
rect 2214 678 2243 818
rect 2289 678 2318 818
rect 2214 573 2318 678
rect 2418 726 2522 939
rect 2418 586 2447 726
rect 2493 586 2522 726
rect 2418 573 2522 586
rect 2622 818 2710 939
rect 2622 678 2651 818
rect 2697 678 2710 818
rect 2622 573 2710 678
<< mvndiffc >>
rect 56 147 102 287
rect 464 82 510 128
rect 996 147 1042 287
rect 1424 82 1470 128
rect 1832 180 1878 320
rect 2243 82 2289 128
rect 2651 180 2697 320
<< mvpdiffc >>
rect 56 786 102 926
rect 260 586 306 726
rect 464 786 510 926
rect 668 586 714 726
rect 872 786 918 926
rect 1016 678 1062 818
rect 1220 586 1266 726
rect 1424 678 1470 818
rect 1628 586 1674 726
rect 1832 678 1878 818
rect 2039 586 2085 726
rect 2243 678 2289 818
rect 2447 586 2493 726
rect 2651 678 2697 818
<< polysilicon >>
rect 131 939 231 983
rect 335 939 435 983
rect 539 939 639 983
rect 743 939 843 983
rect 1091 939 1191 983
rect 1295 939 1395 983
rect 1499 939 1599 983
rect 1703 939 1803 983
rect 1910 939 2010 983
rect 2114 939 2214 983
rect 2318 939 2418 983
rect 2522 939 2622 983
rect 131 540 231 573
rect 131 494 144 540
rect 190 494 231 540
rect 131 377 231 494
rect 335 433 435 573
rect 539 433 639 573
rect 335 412 639 433
rect 335 377 366 412
rect 131 333 251 377
rect 315 366 366 377
rect 412 393 639 412
rect 412 366 435 393
rect 315 333 435 366
rect 539 377 639 393
rect 743 529 843 573
rect 743 483 756 529
rect 802 483 843 529
rect 743 377 843 483
rect 1091 522 1191 573
rect 1091 476 1132 522
rect 1178 476 1191 522
rect 1091 377 1191 476
rect 1295 433 1395 573
rect 1499 433 1599 573
rect 1295 412 1599 433
rect 1295 377 1308 412
rect 539 333 659 377
rect 723 333 843 377
rect 1071 333 1191 377
rect 1275 366 1308 377
rect 1354 393 1599 412
rect 1354 366 1395 393
rect 1275 333 1395 366
rect 1499 377 1599 393
rect 1703 412 1803 573
rect 1703 377 1716 412
rect 1499 333 1619 377
rect 1683 366 1716 377
rect 1762 366 1803 412
rect 1683 333 1803 366
rect 1910 515 2010 573
rect 1910 469 1951 515
rect 1997 469 2010 515
rect 1910 377 2010 469
rect 2114 433 2214 573
rect 2318 433 2418 573
rect 2114 412 2418 433
rect 2114 377 2155 412
rect 1910 333 2030 377
rect 2094 366 2155 377
rect 2201 393 2418 412
rect 2201 366 2214 393
rect 2094 333 2214 366
rect 2318 377 2418 393
rect 2522 515 2622 573
rect 2522 469 2535 515
rect 2581 469 2622 515
rect 2522 377 2622 469
rect 2318 333 2438 377
rect 2502 333 2622 377
rect 131 25 251 69
rect 315 25 435 69
rect 539 25 659 69
rect 723 25 843 69
rect 1071 25 1191 69
rect 1275 25 1395 69
rect 1499 25 1619 69
rect 1683 25 1803 69
rect 1910 25 2030 69
rect 2094 25 2214 69
rect 2318 25 2438 69
rect 2502 25 2622 69
<< polycontact >>
rect 144 494 190 540
rect 366 366 412 412
rect 756 483 802 529
rect 1132 476 1178 522
rect 1308 366 1354 412
rect 1716 366 1762 412
rect 1951 469 1997 515
rect 2155 366 2201 412
rect 2535 469 2581 515
<< metal1 >>
rect 0 926 2800 1098
rect 0 918 56 926
rect 102 918 464 926
rect 56 775 102 786
rect 510 918 872 926
rect 464 775 510 786
rect 918 918 2800 926
rect 872 775 918 786
rect 1016 818 2697 829
rect 260 726 306 737
rect 23 540 194 654
rect 668 726 714 737
rect 306 586 668 621
rect 1062 783 1424 818
rect 1016 667 1062 678
rect 1220 726 1266 737
rect 714 586 1220 621
rect 1470 783 1832 818
rect 1424 667 1470 678
rect 1628 726 1674 737
rect 1266 586 1628 621
rect 1878 783 2243 818
rect 1832 667 1878 678
rect 2039 726 2085 737
rect 260 575 1674 586
rect 1808 586 2039 621
rect 2289 783 2651 818
rect 2243 667 2289 678
rect 2447 726 2493 737
rect 2085 586 2447 621
rect 2651 667 2697 678
rect 2493 586 2697 621
rect 1808 575 2697 586
rect 23 494 144 540
rect 190 529 194 540
rect 190 494 756 529
rect 23 483 756 494
rect 802 483 813 529
rect 1121 476 1132 522
rect 1178 476 1762 522
rect 165 412 418 430
rect 165 366 366 412
rect 412 366 418 412
rect 165 354 418 366
rect 1051 412 1354 430
rect 1051 366 1308 412
rect 1051 354 1354 366
rect 1521 412 1762 476
rect 1521 366 1716 412
rect 1521 354 1762 366
rect 1808 320 1894 575
rect 1940 469 1951 515
rect 1997 469 2535 515
rect 2581 469 2592 515
rect 1808 298 1832 320
rect 56 287 1832 298
rect 102 185 996 287
rect 56 136 102 147
rect 1042 185 1832 287
rect 1878 180 1894 320
rect 1989 412 2210 423
rect 1989 366 2155 412
rect 2201 366 2210 412
rect 1989 242 2210 366
rect 2355 242 2592 469
rect 2651 320 2697 575
rect 1832 169 1894 180
rect 2651 169 2697 180
rect 464 128 510 139
rect 996 136 1042 147
rect 0 82 464 90
rect 1424 128 1470 139
rect 510 82 1424 90
rect 2243 128 2289 139
rect 1470 82 2243 90
rect 2289 82 2800 90
rect 0 -90 2800 82
<< labels >>
flabel metal1 s 1940 469 2592 515 0 FreeSans 200 0 0 0 A1
port 1 nsew default input
flabel metal1 s 1989 242 2210 423 0 FreeSans 200 0 0 0 A2
port 2 nsew default input
flabel metal1 s 1121 476 1762 522 0 FreeSans 200 0 0 0 B1
port 3 nsew default input
flabel metal1 s 1051 354 1354 430 0 FreeSans 200 0 0 0 B2
port 4 nsew default input
flabel metal1 s 23 529 194 654 0 FreeSans 200 0 0 0 C1
port 5 nsew default input
flabel metal1 s 165 354 418 430 0 FreeSans 200 0 0 0 C2
port 6 nsew default input
flabel metal1 s 0 918 2800 1098 0 FreeSans 200 0 0 0 VDD
port 8 nsew power bidirectional abutment
flabel metal1 s 2243 90 2289 139 0 FreeSans 200 0 0 0 VSS
port 11 nsew ground bidirectional abutment
flabel metal1 s 2447 621 2493 737 0 FreeSans 200 0 0 0 ZN
port 7 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 9 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 10 nsew ground bidirectional
rlabel metal1 s 2355 242 2592 469 1 A1
port 1 nsew default input
rlabel metal1 s 1521 354 1762 476 1 B1
port 3 nsew default input
rlabel metal1 s 23 483 813 529 1 C1
port 5 nsew default input
rlabel metal1 s 2039 621 2085 737 1 ZN
port 7 nsew default output
rlabel metal1 s 1808 575 2697 621 1 ZN
port 7 nsew default output
rlabel metal1 s 2651 298 2697 575 1 ZN
port 7 nsew default output
rlabel metal1 s 1808 298 1894 575 1 ZN
port 7 nsew default output
rlabel metal1 s 2651 202 2697 298 1 ZN
port 7 nsew default output
rlabel metal1 s 56 202 1894 298 1 ZN
port 7 nsew default output
rlabel metal1 s 2651 185 2697 202 1 ZN
port 7 nsew default output
rlabel metal1 s 56 185 1894 202 1 ZN
port 7 nsew default output
rlabel metal1 s 2651 169 2697 185 1 ZN
port 7 nsew default output
rlabel metal1 s 1832 169 1894 185 1 ZN
port 7 nsew default output
rlabel metal1 s 996 169 1042 185 1 ZN
port 7 nsew default output
rlabel metal1 s 56 169 102 185 1 ZN
port 7 nsew default output
rlabel metal1 s 996 136 1042 169 1 ZN
port 7 nsew default output
rlabel metal1 s 56 136 102 169 1 ZN
port 7 nsew default output
rlabel metal1 s 872 775 918 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 464 775 510 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 56 775 102 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1424 90 1470 139 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 464 90 510 139 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 2800 90 1 VSS
port 11 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2800 1008
string GDS_END 1247510
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1240474
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
