magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
use 5LM_METAL_RAIL  5LM_METAL_RAIL_0
timestamp 1698431365
transform 1 0 0 0 1 0
box -32 13097 15032 69968
use Bondpad_5LM  Bondpad_5LM_0
timestamp 1698431365
transform 1 0 1100 0 1 0
box -400 0 13200 13065
<< properties >>
string GDS_END 867940
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 867862
<< end >>
