magic
tech gf180mcuD
magscale 1 10
timestamp 1698431365
<< metal3 >>
rect 63 69625 139 69635
rect 63 69569 73 69625
rect 129 69569 139 69625
rect 63 69513 139 69569
rect 63 69457 73 69513
rect 129 69457 139 69513
rect 63 69401 139 69457
rect 63 69345 73 69401
rect 129 69345 139 69401
rect 63 69289 139 69345
rect 63 69233 73 69289
rect 129 69233 139 69289
rect 63 69177 139 69233
rect 63 69121 73 69177
rect 129 69121 139 69177
rect 63 69065 139 69121
rect 63 69009 73 69065
rect 129 69009 139 69065
rect 63 68953 139 69009
rect 63 68897 73 68953
rect 129 68897 139 68953
rect 63 68841 139 68897
rect 63 68785 73 68841
rect 129 68785 139 68841
rect 63 68729 139 68785
rect 63 68673 73 68729
rect 129 68673 139 68729
rect 63 68617 139 68673
rect 63 68561 73 68617
rect 129 68561 139 68617
rect 63 68505 139 68561
rect 63 68449 73 68505
rect 129 68449 139 68505
rect 63 68439 139 68449
rect 63 68153 139 68163
rect 63 68097 73 68153
rect 129 68097 139 68153
rect 63 68041 139 68097
rect 63 67985 73 68041
rect 129 67985 139 68041
rect 63 67929 139 67985
rect 63 67873 73 67929
rect 129 67873 139 67929
rect 63 67817 139 67873
rect 63 67761 73 67817
rect 129 67761 139 67817
rect 63 67705 139 67761
rect 63 67649 73 67705
rect 129 67649 139 67705
rect 63 67593 139 67649
rect 63 67537 73 67593
rect 129 67537 139 67593
rect 63 67481 139 67537
rect 63 67425 73 67481
rect 129 67425 139 67481
rect 63 67369 139 67425
rect 63 67313 73 67369
rect 129 67313 139 67369
rect 63 67257 139 67313
rect 63 67201 73 67257
rect 129 67201 139 67257
rect 63 67145 139 67201
rect 63 67089 73 67145
rect 129 67089 139 67145
rect 63 67033 139 67089
rect 63 66977 73 67033
rect 129 66977 139 67033
rect 63 66921 139 66977
rect 63 66865 73 66921
rect 129 66865 139 66921
rect 63 66855 139 66865
rect 63 66552 139 66562
rect 63 66496 73 66552
rect 129 66496 139 66552
rect 63 66440 139 66496
rect 63 66384 73 66440
rect 129 66384 139 66440
rect 63 66328 139 66384
rect 63 66272 73 66328
rect 129 66272 139 66328
rect 63 66216 139 66272
rect 63 66160 73 66216
rect 129 66160 139 66216
rect 63 66104 139 66160
rect 63 66048 73 66104
rect 129 66048 139 66104
rect 63 65992 139 66048
rect 63 65936 73 65992
rect 129 65936 139 65992
rect 63 65880 139 65936
rect 63 65824 73 65880
rect 129 65824 139 65880
rect 63 65768 139 65824
rect 63 65712 73 65768
rect 129 65712 139 65768
rect 63 65656 139 65712
rect 63 65600 73 65656
rect 129 65600 139 65656
rect 63 65544 139 65600
rect 63 65488 73 65544
rect 129 65488 139 65544
rect 63 65432 139 65488
rect 63 65376 73 65432
rect 129 65376 139 65432
rect 63 65320 139 65376
rect 63 65264 73 65320
rect 129 65264 139 65320
rect 63 65254 139 65264
rect 63 64944 139 64954
rect 63 64888 73 64944
rect 129 64888 139 64944
rect 63 64832 139 64888
rect 63 64776 73 64832
rect 129 64776 139 64832
rect 63 64720 139 64776
rect 63 64664 73 64720
rect 129 64664 139 64720
rect 63 64608 139 64664
rect 63 64552 73 64608
rect 129 64552 139 64608
rect 63 64496 139 64552
rect 63 64440 73 64496
rect 129 64440 139 64496
rect 63 64384 139 64440
rect 63 64328 73 64384
rect 129 64328 139 64384
rect 63 64272 139 64328
rect 63 64216 73 64272
rect 129 64216 139 64272
rect 63 64160 139 64216
rect 63 64104 73 64160
rect 129 64104 139 64160
rect 63 64048 139 64104
rect 63 63992 73 64048
rect 129 63992 139 64048
rect 63 63936 139 63992
rect 63 63880 73 63936
rect 129 63880 139 63936
rect 63 63824 139 63880
rect 63 63768 73 63824
rect 129 63768 139 63824
rect 63 63712 139 63768
rect 63 63656 73 63712
rect 129 63656 139 63712
rect 63 63646 139 63656
rect 63 63344 139 63354
rect 63 63288 73 63344
rect 129 63288 139 63344
rect 63 63232 139 63288
rect 63 63176 73 63232
rect 129 63176 139 63232
rect 63 63120 139 63176
rect 63 63064 73 63120
rect 129 63064 139 63120
rect 63 63008 139 63064
rect 63 62952 73 63008
rect 129 62952 139 63008
rect 63 62896 139 62952
rect 63 62840 73 62896
rect 129 62840 139 62896
rect 63 62784 139 62840
rect 63 62728 73 62784
rect 129 62728 139 62784
rect 63 62672 139 62728
rect 63 62616 73 62672
rect 129 62616 139 62672
rect 63 62560 139 62616
rect 63 62504 73 62560
rect 129 62504 139 62560
rect 63 62448 139 62504
rect 63 62392 73 62448
rect 129 62392 139 62448
rect 63 62336 139 62392
rect 63 62280 73 62336
rect 129 62280 139 62336
rect 63 62224 139 62280
rect 63 62168 73 62224
rect 129 62168 139 62224
rect 63 62112 139 62168
rect 63 62056 73 62112
rect 129 62056 139 62112
rect 63 62046 139 62056
rect 63 61745 139 61755
rect 63 61689 73 61745
rect 129 61689 139 61745
rect 63 61633 139 61689
rect 63 61577 73 61633
rect 129 61577 139 61633
rect 63 61521 139 61577
rect 63 61465 73 61521
rect 129 61465 139 61521
rect 63 61409 139 61465
rect 63 61353 73 61409
rect 129 61353 139 61409
rect 63 61297 139 61353
rect 63 61241 73 61297
rect 129 61241 139 61297
rect 63 61185 139 61241
rect 63 61129 73 61185
rect 129 61129 139 61185
rect 63 61073 139 61129
rect 63 61017 73 61073
rect 129 61017 139 61073
rect 63 60961 139 61017
rect 63 60905 73 60961
rect 129 60905 139 60961
rect 63 60849 139 60905
rect 63 60793 73 60849
rect 129 60793 139 60849
rect 63 60737 139 60793
rect 63 60681 73 60737
rect 129 60681 139 60737
rect 63 60625 139 60681
rect 63 60569 73 60625
rect 129 60569 139 60625
rect 63 60513 139 60569
rect 63 60457 73 60513
rect 129 60457 139 60513
rect 63 60447 139 60457
rect 63 60152 139 60162
rect 63 60096 73 60152
rect 129 60096 139 60152
rect 63 60040 139 60096
rect 63 59984 73 60040
rect 129 59984 139 60040
rect 63 59928 139 59984
rect 63 59872 73 59928
rect 129 59872 139 59928
rect 63 59816 139 59872
rect 63 59760 73 59816
rect 129 59760 139 59816
rect 63 59704 139 59760
rect 63 59648 73 59704
rect 129 59648 139 59704
rect 63 59592 139 59648
rect 63 59536 73 59592
rect 129 59536 139 59592
rect 63 59480 139 59536
rect 63 59424 73 59480
rect 129 59424 139 59480
rect 63 59368 139 59424
rect 63 59312 73 59368
rect 129 59312 139 59368
rect 63 59256 139 59312
rect 63 59200 73 59256
rect 129 59200 139 59256
rect 63 59144 139 59200
rect 63 59088 73 59144
rect 129 59088 139 59144
rect 63 59032 139 59088
rect 63 58976 73 59032
rect 129 58976 139 59032
rect 63 58920 139 58976
rect 63 58864 73 58920
rect 129 58864 139 58920
rect 63 58854 139 58864
rect 63 58547 139 58557
rect 63 58491 73 58547
rect 129 58491 139 58547
rect 63 58435 139 58491
rect 63 58379 73 58435
rect 129 58379 139 58435
rect 63 58323 139 58379
rect 63 58267 73 58323
rect 129 58267 139 58323
rect 63 58211 139 58267
rect 63 58155 73 58211
rect 129 58155 139 58211
rect 63 58099 139 58155
rect 63 58043 73 58099
rect 129 58043 139 58099
rect 63 57987 139 58043
rect 63 57931 73 57987
rect 129 57931 139 57987
rect 63 57875 139 57931
rect 63 57819 73 57875
rect 129 57819 139 57875
rect 63 57763 139 57819
rect 63 57707 73 57763
rect 129 57707 139 57763
rect 63 57651 139 57707
rect 63 57595 73 57651
rect 129 57595 139 57651
rect 63 57539 139 57595
rect 63 57483 73 57539
rect 129 57483 139 57539
rect 63 57427 139 57483
rect 63 57371 73 57427
rect 129 57371 139 57427
rect 63 57315 139 57371
rect 63 57259 73 57315
rect 129 57259 139 57315
rect 63 57249 139 57259
rect 63 56949 139 56959
rect 63 56893 73 56949
rect 129 56893 139 56949
rect 63 56837 139 56893
rect 63 56781 73 56837
rect 129 56781 139 56837
rect 63 56725 139 56781
rect 63 56669 73 56725
rect 129 56669 139 56725
rect 63 56613 139 56669
rect 63 56557 73 56613
rect 129 56557 139 56613
rect 63 56501 139 56557
rect 63 56445 73 56501
rect 129 56445 139 56501
rect 63 56389 139 56445
rect 63 56333 73 56389
rect 129 56333 139 56389
rect 63 56277 139 56333
rect 63 56221 73 56277
rect 129 56221 139 56277
rect 63 56165 139 56221
rect 63 56109 73 56165
rect 129 56109 139 56165
rect 63 56053 139 56109
rect 63 55997 73 56053
rect 129 55997 139 56053
rect 63 55941 139 55997
rect 63 55885 73 55941
rect 129 55885 139 55941
rect 63 55829 139 55885
rect 63 55773 73 55829
rect 129 55773 139 55829
rect 63 55717 139 55773
rect 63 55661 73 55717
rect 129 55661 139 55717
rect 63 55651 139 55661
rect 63 55348 139 55358
rect 63 55292 73 55348
rect 129 55292 139 55348
rect 63 55236 139 55292
rect 63 55180 73 55236
rect 129 55180 139 55236
rect 63 55124 139 55180
rect 63 55068 73 55124
rect 129 55068 139 55124
rect 63 55012 139 55068
rect 63 54956 73 55012
rect 129 54956 139 55012
rect 63 54900 139 54956
rect 63 54844 73 54900
rect 129 54844 139 54900
rect 63 54788 139 54844
rect 63 54732 73 54788
rect 129 54732 139 54788
rect 63 54676 139 54732
rect 63 54620 73 54676
rect 129 54620 139 54676
rect 63 54564 139 54620
rect 63 54508 73 54564
rect 129 54508 139 54564
rect 63 54452 139 54508
rect 63 54396 73 54452
rect 129 54396 139 54452
rect 63 54340 139 54396
rect 63 54284 73 54340
rect 129 54284 139 54340
rect 63 54228 139 54284
rect 63 54172 73 54228
rect 129 54172 139 54228
rect 63 54116 139 54172
rect 63 54060 73 54116
rect 129 54060 139 54116
rect 63 54050 139 54060
rect 63 53735 139 53745
rect 63 53679 73 53735
rect 129 53679 139 53735
rect 63 53623 139 53679
rect 63 53567 73 53623
rect 129 53567 139 53623
rect 63 53511 139 53567
rect 63 53455 73 53511
rect 129 53455 139 53511
rect 63 53399 139 53455
rect 63 53343 73 53399
rect 129 53343 139 53399
rect 63 53287 139 53343
rect 63 53231 73 53287
rect 129 53231 139 53287
rect 63 53175 139 53231
rect 63 53119 73 53175
rect 129 53119 139 53175
rect 63 53063 139 53119
rect 63 53007 73 53063
rect 129 53007 139 53063
rect 63 52951 139 53007
rect 63 52895 73 52951
rect 129 52895 139 52951
rect 63 52839 139 52895
rect 63 52783 73 52839
rect 129 52783 139 52839
rect 63 52727 139 52783
rect 63 52671 73 52727
rect 129 52671 139 52727
rect 63 52615 139 52671
rect 63 52559 73 52615
rect 129 52559 139 52615
rect 63 52503 139 52559
rect 63 52447 73 52503
rect 129 52447 139 52503
rect 63 52437 139 52447
rect 63 52149 139 52159
rect 63 52093 73 52149
rect 129 52093 139 52149
rect 63 52037 139 52093
rect 63 51981 73 52037
rect 129 51981 139 52037
rect 63 51925 139 51981
rect 63 51869 73 51925
rect 129 51869 139 51925
rect 63 51813 139 51869
rect 63 51757 73 51813
rect 129 51757 139 51813
rect 63 51701 139 51757
rect 63 51645 73 51701
rect 129 51645 139 51701
rect 63 51589 139 51645
rect 63 51533 73 51589
rect 129 51533 139 51589
rect 63 51477 139 51533
rect 63 51421 73 51477
rect 129 51421 139 51477
rect 63 51365 139 51421
rect 63 51309 73 51365
rect 129 51309 139 51365
rect 63 51253 139 51309
rect 63 51197 73 51253
rect 129 51197 139 51253
rect 63 51141 139 51197
rect 63 51085 73 51141
rect 129 51085 139 51141
rect 63 51029 139 51085
rect 63 50973 73 51029
rect 129 50973 139 51029
rect 63 50917 139 50973
rect 63 50861 73 50917
rect 129 50861 139 50917
rect 63 50851 139 50861
rect 64 50538 140 50548
rect 64 50482 74 50538
rect 130 50482 140 50538
rect 64 50426 140 50482
rect 64 50370 74 50426
rect 130 50370 140 50426
rect 64 50314 140 50370
rect 64 50258 74 50314
rect 130 50258 140 50314
rect 64 50202 140 50258
rect 64 50146 74 50202
rect 130 50146 140 50202
rect 64 50090 140 50146
rect 64 50034 74 50090
rect 130 50034 140 50090
rect 64 49978 140 50034
rect 64 49922 74 49978
rect 130 49922 140 49978
rect 64 49866 140 49922
rect 64 49810 74 49866
rect 130 49810 140 49866
rect 64 49754 140 49810
rect 64 49698 74 49754
rect 130 49698 140 49754
rect 64 49642 140 49698
rect 64 49586 74 49642
rect 130 49586 140 49642
rect 64 49530 140 49586
rect 64 49474 74 49530
rect 130 49474 140 49530
rect 64 49418 140 49474
rect 64 49362 74 49418
rect 130 49362 140 49418
rect 64 49306 140 49362
rect 64 49250 74 49306
rect 130 49250 140 49306
rect 64 49240 140 49250
rect 63 48884 139 48894
rect 63 48828 73 48884
rect 129 48828 139 48884
rect 63 48772 139 48828
rect 63 48716 73 48772
rect 129 48716 139 48772
rect 63 48660 139 48716
rect 63 48604 73 48660
rect 129 48604 139 48660
rect 63 48548 139 48604
rect 63 48492 73 48548
rect 129 48492 139 48548
rect 63 48436 139 48492
rect 63 48380 73 48436
rect 129 48380 139 48436
rect 63 48324 139 48380
rect 63 48268 73 48324
rect 129 48268 139 48324
rect 63 48212 139 48268
rect 63 48156 73 48212
rect 129 48156 139 48212
rect 63 48100 139 48156
rect 63 48044 73 48100
rect 129 48044 139 48100
rect 63 47988 139 48044
rect 63 47932 73 47988
rect 129 47932 139 47988
rect 63 47876 139 47932
rect 63 47820 73 47876
rect 129 47820 139 47876
rect 63 47764 139 47820
rect 63 47708 73 47764
rect 129 47708 139 47764
rect 63 47652 139 47708
rect 63 47596 73 47652
rect 129 47596 139 47652
rect 63 47540 139 47596
rect 63 47484 73 47540
rect 129 47484 139 47540
rect 63 47428 139 47484
rect 63 47372 73 47428
rect 129 47372 139 47428
rect 63 47316 139 47372
rect 63 47260 73 47316
rect 129 47260 139 47316
rect 63 47204 139 47260
rect 63 47148 73 47204
rect 129 47148 139 47204
rect 63 47092 139 47148
rect 63 47036 73 47092
rect 129 47036 139 47092
rect 63 46980 139 47036
rect 63 46924 73 46980
rect 129 46924 139 46980
rect 63 46868 139 46924
rect 63 46812 73 46868
rect 129 46812 139 46868
rect 63 46756 139 46812
rect 63 46700 73 46756
rect 129 46700 139 46756
rect 63 46644 139 46700
rect 63 46588 73 46644
rect 129 46588 139 46644
rect 63 46532 139 46588
rect 63 46476 73 46532
rect 129 46476 139 46532
rect 63 46420 139 46476
rect 63 46364 73 46420
rect 129 46364 139 46420
rect 63 46308 139 46364
rect 63 46252 73 46308
rect 129 46252 139 46308
rect 63 46196 139 46252
rect 63 46140 73 46196
rect 129 46140 139 46196
rect 63 46130 139 46140
rect 63 45670 139 45680
rect 63 45614 73 45670
rect 129 45614 139 45670
rect 63 45558 139 45614
rect 63 45502 73 45558
rect 129 45502 139 45558
rect 63 45446 139 45502
rect 63 45390 73 45446
rect 129 45390 139 45446
rect 63 45334 139 45390
rect 63 45278 73 45334
rect 129 45278 139 45334
rect 63 45222 139 45278
rect 63 45166 73 45222
rect 129 45166 139 45222
rect 63 45110 139 45166
rect 63 45054 73 45110
rect 129 45054 139 45110
rect 63 44998 139 45054
rect 63 44942 73 44998
rect 129 44942 139 44998
rect 63 44886 139 44942
rect 63 44830 73 44886
rect 129 44830 139 44886
rect 63 44774 139 44830
rect 63 44718 73 44774
rect 129 44718 139 44774
rect 63 44662 139 44718
rect 63 44606 73 44662
rect 129 44606 139 44662
rect 63 44550 139 44606
rect 63 44494 73 44550
rect 129 44494 139 44550
rect 63 44438 139 44494
rect 63 44382 73 44438
rect 129 44382 139 44438
rect 63 44326 139 44382
rect 63 44270 73 44326
rect 129 44270 139 44326
rect 63 44214 139 44270
rect 63 44158 73 44214
rect 129 44158 139 44214
rect 63 44102 139 44158
rect 63 44046 73 44102
rect 129 44046 139 44102
rect 63 43990 139 44046
rect 63 43934 73 43990
rect 129 43934 139 43990
rect 63 43878 139 43934
rect 63 43822 73 43878
rect 129 43822 139 43878
rect 63 43766 139 43822
rect 63 43710 73 43766
rect 129 43710 139 43766
rect 63 43654 139 43710
rect 63 43598 73 43654
rect 129 43598 139 43654
rect 63 43542 139 43598
rect 63 43486 73 43542
rect 129 43486 139 43542
rect 63 43430 139 43486
rect 63 43374 73 43430
rect 129 43374 139 43430
rect 63 43318 139 43374
rect 63 43262 73 43318
rect 129 43262 139 43318
rect 63 43206 139 43262
rect 63 43150 73 43206
rect 129 43150 139 43206
rect 63 43094 139 43150
rect 63 43038 73 43094
rect 129 43038 139 43094
rect 63 42982 139 43038
rect 63 42926 73 42982
rect 129 42926 139 42982
rect 63 42916 139 42926
rect 64 42549 140 42559
rect 64 42493 74 42549
rect 130 42493 140 42549
rect 64 42437 140 42493
rect 64 42381 74 42437
rect 130 42381 140 42437
rect 64 42325 140 42381
rect 64 42269 74 42325
rect 130 42269 140 42325
rect 64 42213 140 42269
rect 64 42157 74 42213
rect 130 42157 140 42213
rect 64 42101 140 42157
rect 64 42045 74 42101
rect 130 42045 140 42101
rect 64 41989 140 42045
rect 64 41933 74 41989
rect 130 41933 140 41989
rect 64 41877 140 41933
rect 64 41821 74 41877
rect 130 41821 140 41877
rect 64 41765 140 41821
rect 64 41709 74 41765
rect 130 41709 140 41765
rect 64 41653 140 41709
rect 64 41597 74 41653
rect 130 41597 140 41653
rect 64 41541 140 41597
rect 64 41485 74 41541
rect 130 41485 140 41541
rect 64 41429 140 41485
rect 64 41373 74 41429
rect 130 41373 140 41429
rect 64 41317 140 41373
rect 64 41261 74 41317
rect 130 41261 140 41317
rect 64 41251 140 41261
rect 64 40951 140 40961
rect 64 40895 74 40951
rect 130 40895 140 40951
rect 64 40839 140 40895
rect 64 40783 74 40839
rect 130 40783 140 40839
rect 64 40727 140 40783
rect 64 40671 74 40727
rect 130 40671 140 40727
rect 64 40615 140 40671
rect 64 40559 74 40615
rect 130 40559 140 40615
rect 64 40503 140 40559
rect 64 40447 74 40503
rect 130 40447 140 40503
rect 64 40391 140 40447
rect 64 40335 74 40391
rect 130 40335 140 40391
rect 64 40279 140 40335
rect 64 40223 74 40279
rect 130 40223 140 40279
rect 64 40167 140 40223
rect 64 40111 74 40167
rect 130 40111 140 40167
rect 64 40055 140 40111
rect 64 39999 74 40055
rect 130 39999 140 40055
rect 64 39943 140 39999
rect 64 39887 74 39943
rect 130 39887 140 39943
rect 64 39831 140 39887
rect 64 39775 74 39831
rect 130 39775 140 39831
rect 64 39719 140 39775
rect 64 39663 74 39719
rect 130 39663 140 39719
rect 64 39653 140 39663
rect 63 39276 139 39286
rect 63 39220 73 39276
rect 129 39220 139 39276
rect 63 39164 139 39220
rect 63 39108 73 39164
rect 129 39108 139 39164
rect 63 39052 139 39108
rect 63 38996 73 39052
rect 129 38996 139 39052
rect 63 38940 139 38996
rect 63 38884 73 38940
rect 129 38884 139 38940
rect 63 38828 139 38884
rect 63 38772 73 38828
rect 129 38772 139 38828
rect 63 38716 139 38772
rect 63 38660 73 38716
rect 129 38660 139 38716
rect 63 38604 139 38660
rect 63 38548 73 38604
rect 129 38548 139 38604
rect 63 38492 139 38548
rect 63 38436 73 38492
rect 129 38436 139 38492
rect 63 38380 139 38436
rect 63 38324 73 38380
rect 129 38324 139 38380
rect 63 38268 139 38324
rect 63 38212 73 38268
rect 129 38212 139 38268
rect 63 38156 139 38212
rect 63 38100 73 38156
rect 129 38100 139 38156
rect 63 38044 139 38100
rect 63 37988 73 38044
rect 129 37988 139 38044
rect 63 37932 139 37988
rect 63 37876 73 37932
rect 129 37876 139 37932
rect 63 37820 139 37876
rect 63 37764 73 37820
rect 129 37764 139 37820
rect 63 37708 139 37764
rect 63 37652 73 37708
rect 129 37652 139 37708
rect 63 37596 139 37652
rect 63 37540 73 37596
rect 129 37540 139 37596
rect 63 37484 139 37540
rect 63 37428 73 37484
rect 129 37428 139 37484
rect 63 37372 139 37428
rect 63 37316 73 37372
rect 129 37316 139 37372
rect 63 37260 139 37316
rect 63 37204 73 37260
rect 129 37204 139 37260
rect 63 37148 139 37204
rect 63 37092 73 37148
rect 129 37092 139 37148
rect 63 37036 139 37092
rect 63 36980 73 37036
rect 129 36980 139 37036
rect 63 36924 139 36980
rect 63 36868 73 36924
rect 129 36868 139 36924
rect 63 36812 139 36868
rect 63 36756 73 36812
rect 129 36756 139 36812
rect 63 36700 139 36756
rect 63 36644 73 36700
rect 129 36644 139 36700
rect 63 36588 139 36644
rect 63 36532 73 36588
rect 129 36532 139 36588
rect 63 36522 139 36532
rect 63 36075 139 36085
rect 63 36019 73 36075
rect 129 36019 139 36075
rect 63 35963 139 36019
rect 63 35907 73 35963
rect 129 35907 139 35963
rect 63 35851 139 35907
rect 63 35795 73 35851
rect 129 35795 139 35851
rect 63 35739 139 35795
rect 63 35683 73 35739
rect 129 35683 139 35739
rect 63 35627 139 35683
rect 63 35571 73 35627
rect 129 35571 139 35627
rect 63 35515 139 35571
rect 63 35459 73 35515
rect 129 35459 139 35515
rect 63 35403 139 35459
rect 63 35347 73 35403
rect 129 35347 139 35403
rect 63 35291 139 35347
rect 63 35235 73 35291
rect 129 35235 139 35291
rect 63 35179 139 35235
rect 63 35123 73 35179
rect 129 35123 139 35179
rect 63 35067 139 35123
rect 63 35011 73 35067
rect 129 35011 139 35067
rect 63 34955 139 35011
rect 63 34899 73 34955
rect 129 34899 139 34955
rect 63 34843 139 34899
rect 63 34787 73 34843
rect 129 34787 139 34843
rect 63 34731 139 34787
rect 63 34675 73 34731
rect 129 34675 139 34731
rect 63 34619 139 34675
rect 63 34563 73 34619
rect 129 34563 139 34619
rect 63 34507 139 34563
rect 63 34451 73 34507
rect 129 34451 139 34507
rect 63 34395 139 34451
rect 63 34339 73 34395
rect 129 34339 139 34395
rect 63 34283 139 34339
rect 63 34227 73 34283
rect 129 34227 139 34283
rect 63 34171 139 34227
rect 63 34115 73 34171
rect 129 34115 139 34171
rect 63 34059 139 34115
rect 63 34003 73 34059
rect 129 34003 139 34059
rect 63 33947 139 34003
rect 63 33891 73 33947
rect 129 33891 139 33947
rect 63 33835 139 33891
rect 63 33779 73 33835
rect 129 33779 139 33835
rect 63 33723 139 33779
rect 63 33667 73 33723
rect 129 33667 139 33723
rect 63 33611 139 33667
rect 63 33555 73 33611
rect 129 33555 139 33611
rect 63 33499 139 33555
rect 63 33443 73 33499
rect 129 33443 139 33499
rect 63 33387 139 33443
rect 63 33331 73 33387
rect 129 33331 139 33387
rect 63 33321 139 33331
rect 63 32879 139 32889
rect 63 32823 73 32879
rect 129 32823 139 32879
rect 63 32767 139 32823
rect 63 32711 73 32767
rect 129 32711 139 32767
rect 63 32655 139 32711
rect 63 32599 73 32655
rect 129 32599 139 32655
rect 63 32543 139 32599
rect 63 32487 73 32543
rect 129 32487 139 32543
rect 63 32431 139 32487
rect 63 32375 73 32431
rect 129 32375 139 32431
rect 63 32319 139 32375
rect 63 32263 73 32319
rect 129 32263 139 32319
rect 63 32207 139 32263
rect 63 32151 73 32207
rect 129 32151 139 32207
rect 63 32095 139 32151
rect 63 32039 73 32095
rect 129 32039 139 32095
rect 63 31983 139 32039
rect 63 31927 73 31983
rect 129 31927 139 31983
rect 63 31871 139 31927
rect 63 31815 73 31871
rect 129 31815 139 31871
rect 63 31759 139 31815
rect 63 31703 73 31759
rect 129 31703 139 31759
rect 63 31647 139 31703
rect 63 31591 73 31647
rect 129 31591 139 31647
rect 63 31535 139 31591
rect 63 31479 73 31535
rect 129 31479 139 31535
rect 63 31423 139 31479
rect 63 31367 73 31423
rect 129 31367 139 31423
rect 63 31311 139 31367
rect 63 31255 73 31311
rect 129 31255 139 31311
rect 63 31199 139 31255
rect 63 31143 73 31199
rect 129 31143 139 31199
rect 63 31087 139 31143
rect 63 31031 73 31087
rect 129 31031 139 31087
rect 63 30975 139 31031
rect 63 30919 73 30975
rect 129 30919 139 30975
rect 63 30863 139 30919
rect 63 30807 73 30863
rect 129 30807 139 30863
rect 63 30751 139 30807
rect 63 30695 73 30751
rect 129 30695 139 30751
rect 63 30639 139 30695
rect 63 30583 73 30639
rect 129 30583 139 30639
rect 63 30527 139 30583
rect 63 30471 73 30527
rect 129 30471 139 30527
rect 63 30415 139 30471
rect 63 30359 73 30415
rect 129 30359 139 30415
rect 63 30303 139 30359
rect 63 30247 73 30303
rect 129 30247 139 30303
rect 63 30191 139 30247
rect 63 30135 73 30191
rect 129 30135 139 30191
rect 63 30125 139 30135
rect 63 29685 139 29695
rect 63 29629 73 29685
rect 129 29629 139 29685
rect 63 29573 139 29629
rect 63 29517 73 29573
rect 129 29517 139 29573
rect 63 29461 139 29517
rect 63 29405 73 29461
rect 129 29405 139 29461
rect 63 29349 139 29405
rect 63 29293 73 29349
rect 129 29293 139 29349
rect 63 29237 139 29293
rect 63 29181 73 29237
rect 129 29181 139 29237
rect 63 29125 139 29181
rect 63 29069 73 29125
rect 129 29069 139 29125
rect 63 29013 139 29069
rect 63 28957 73 29013
rect 129 28957 139 29013
rect 63 28901 139 28957
rect 63 28845 73 28901
rect 129 28845 139 28901
rect 63 28789 139 28845
rect 63 28733 73 28789
rect 129 28733 139 28789
rect 63 28677 139 28733
rect 63 28621 73 28677
rect 129 28621 139 28677
rect 63 28565 139 28621
rect 63 28509 73 28565
rect 129 28509 139 28565
rect 63 28453 139 28509
rect 63 28397 73 28453
rect 129 28397 139 28453
rect 63 28341 139 28397
rect 63 28285 73 28341
rect 129 28285 139 28341
rect 63 28229 139 28285
rect 63 28173 73 28229
rect 129 28173 139 28229
rect 63 28117 139 28173
rect 63 28061 73 28117
rect 129 28061 139 28117
rect 63 28005 139 28061
rect 63 27949 73 28005
rect 129 27949 139 28005
rect 63 27893 139 27949
rect 63 27837 73 27893
rect 129 27837 139 27893
rect 63 27781 139 27837
rect 63 27725 73 27781
rect 129 27725 139 27781
rect 63 27669 139 27725
rect 63 27613 73 27669
rect 129 27613 139 27669
rect 63 27557 139 27613
rect 63 27501 73 27557
rect 129 27501 139 27557
rect 63 27445 139 27501
rect 63 27389 73 27445
rect 129 27389 139 27445
rect 63 27333 139 27389
rect 63 27277 73 27333
rect 129 27277 139 27333
rect 63 27221 139 27277
rect 63 27165 73 27221
rect 129 27165 139 27221
rect 63 27109 139 27165
rect 63 27053 73 27109
rect 129 27053 139 27109
rect 63 26997 139 27053
rect 63 26941 73 26997
rect 129 26941 139 26997
rect 63 26931 139 26941
rect 64 26550 140 26560
rect 64 26494 74 26550
rect 130 26494 140 26550
rect 64 26438 140 26494
rect 64 26382 74 26438
rect 130 26382 140 26438
rect 64 26326 140 26382
rect 64 26270 74 26326
rect 130 26270 140 26326
rect 64 26214 140 26270
rect 64 26158 74 26214
rect 130 26158 140 26214
rect 64 26102 140 26158
rect 64 26046 74 26102
rect 130 26046 140 26102
rect 64 25990 140 26046
rect 64 25934 74 25990
rect 130 25934 140 25990
rect 64 25878 140 25934
rect 64 25822 74 25878
rect 130 25822 140 25878
rect 64 25766 140 25822
rect 64 25710 74 25766
rect 130 25710 140 25766
rect 64 25654 140 25710
rect 64 25598 74 25654
rect 130 25598 140 25654
rect 64 25542 140 25598
rect 64 25486 74 25542
rect 130 25486 140 25542
rect 64 25430 140 25486
rect 64 25374 74 25430
rect 130 25374 140 25430
rect 64 25318 140 25374
rect 64 25262 74 25318
rect 130 25262 140 25318
rect 64 25252 140 25262
rect 64 24957 140 24967
rect 64 24901 74 24957
rect 130 24901 140 24957
rect 64 24845 140 24901
rect 64 24789 74 24845
rect 130 24789 140 24845
rect 64 24733 140 24789
rect 64 24677 74 24733
rect 130 24677 140 24733
rect 64 24621 140 24677
rect 64 24565 74 24621
rect 130 24565 140 24621
rect 64 24509 140 24565
rect 64 24453 74 24509
rect 130 24453 140 24509
rect 64 24397 140 24453
rect 64 24341 74 24397
rect 130 24341 140 24397
rect 64 24285 140 24341
rect 64 24229 74 24285
rect 130 24229 140 24285
rect 64 24173 140 24229
rect 64 24117 74 24173
rect 130 24117 140 24173
rect 64 24061 140 24117
rect 64 24005 74 24061
rect 130 24005 140 24061
rect 64 23949 140 24005
rect 64 23893 74 23949
rect 130 23893 140 23949
rect 64 23837 140 23893
rect 64 23781 74 23837
rect 130 23781 140 23837
rect 64 23725 140 23781
rect 64 23669 74 23725
rect 130 23669 140 23725
rect 64 23659 140 23669
rect 63 23323 139 23333
rect 63 23267 73 23323
rect 129 23267 139 23323
rect 63 23211 139 23267
rect 63 23155 73 23211
rect 129 23155 139 23211
rect 63 23099 139 23155
rect 63 23043 73 23099
rect 129 23043 139 23099
rect 63 22987 139 23043
rect 63 22931 73 22987
rect 129 22931 139 22987
rect 63 22875 139 22931
rect 63 22819 73 22875
rect 129 22819 139 22875
rect 63 22763 139 22819
rect 63 22707 73 22763
rect 129 22707 139 22763
rect 63 22651 139 22707
rect 63 22595 73 22651
rect 129 22595 139 22651
rect 63 22539 139 22595
rect 63 22483 73 22539
rect 129 22483 139 22539
rect 63 22427 139 22483
rect 63 22371 73 22427
rect 129 22371 139 22427
rect 63 22315 139 22371
rect 63 22259 73 22315
rect 129 22259 139 22315
rect 63 22203 139 22259
rect 63 22147 73 22203
rect 129 22147 139 22203
rect 63 22091 139 22147
rect 63 22035 73 22091
rect 129 22035 139 22091
rect 63 21979 139 22035
rect 63 21923 73 21979
rect 129 21923 139 21979
rect 63 21867 139 21923
rect 63 21811 73 21867
rect 129 21811 139 21867
rect 63 21755 139 21811
rect 63 21699 73 21755
rect 129 21699 139 21755
rect 63 21643 139 21699
rect 63 21587 73 21643
rect 129 21587 139 21643
rect 63 21531 139 21587
rect 63 21475 73 21531
rect 129 21475 139 21531
rect 63 21419 139 21475
rect 63 21363 73 21419
rect 129 21363 139 21419
rect 63 21307 139 21363
rect 63 21251 73 21307
rect 129 21251 139 21307
rect 63 21195 139 21251
rect 63 21139 73 21195
rect 129 21139 139 21195
rect 63 21083 139 21139
rect 63 21027 73 21083
rect 129 21027 139 21083
rect 63 20971 139 21027
rect 63 20915 73 20971
rect 129 20915 139 20971
rect 63 20859 139 20915
rect 63 20803 73 20859
rect 129 20803 139 20859
rect 63 20747 139 20803
rect 63 20691 73 20747
rect 129 20691 139 20747
rect 63 20635 139 20691
rect 63 20579 73 20635
rect 129 20579 139 20635
rect 63 20569 139 20579
rect 63 20073 139 20083
rect 63 20017 73 20073
rect 129 20017 139 20073
rect 63 19961 139 20017
rect 63 19905 73 19961
rect 129 19905 139 19961
rect 63 19849 139 19905
rect 63 19793 73 19849
rect 129 19793 139 19849
rect 63 19737 139 19793
rect 63 19681 73 19737
rect 129 19681 139 19737
rect 63 19625 139 19681
rect 63 19569 73 19625
rect 129 19569 139 19625
rect 63 19513 139 19569
rect 63 19457 73 19513
rect 129 19457 139 19513
rect 63 19401 139 19457
rect 63 19345 73 19401
rect 129 19345 139 19401
rect 63 19289 139 19345
rect 63 19233 73 19289
rect 129 19233 139 19289
rect 63 19177 139 19233
rect 63 19121 73 19177
rect 129 19121 139 19177
rect 63 19065 139 19121
rect 63 19009 73 19065
rect 129 19009 139 19065
rect 63 18953 139 19009
rect 63 18897 73 18953
rect 129 18897 139 18953
rect 63 18841 139 18897
rect 63 18785 73 18841
rect 129 18785 139 18841
rect 63 18729 139 18785
rect 63 18673 73 18729
rect 129 18673 139 18729
rect 63 18617 139 18673
rect 63 18561 73 18617
rect 129 18561 139 18617
rect 63 18505 139 18561
rect 63 18449 73 18505
rect 129 18449 139 18505
rect 63 18393 139 18449
rect 63 18337 73 18393
rect 129 18337 139 18393
rect 63 18281 139 18337
rect 63 18225 73 18281
rect 129 18225 139 18281
rect 63 18169 139 18225
rect 63 18113 73 18169
rect 129 18113 139 18169
rect 63 18057 139 18113
rect 63 18001 73 18057
rect 129 18001 139 18057
rect 63 17945 139 18001
rect 63 17889 73 17945
rect 129 17889 139 17945
rect 63 17833 139 17889
rect 63 17777 73 17833
rect 129 17777 139 17833
rect 63 17721 139 17777
rect 63 17665 73 17721
rect 129 17665 139 17721
rect 63 17609 139 17665
rect 63 17553 73 17609
rect 129 17553 139 17609
rect 63 17497 139 17553
rect 63 17441 73 17497
rect 129 17441 139 17497
rect 63 17385 139 17441
rect 63 17329 73 17385
rect 129 17329 139 17385
rect 63 17319 139 17329
rect 63 16872 139 16882
rect 63 16816 73 16872
rect 129 16816 139 16872
rect 63 16760 139 16816
rect 63 16704 73 16760
rect 129 16704 139 16760
rect 63 16648 139 16704
rect 63 16592 73 16648
rect 129 16592 139 16648
rect 63 16536 139 16592
rect 63 16480 73 16536
rect 129 16480 139 16536
rect 63 16424 139 16480
rect 63 16368 73 16424
rect 129 16368 139 16424
rect 63 16312 139 16368
rect 63 16256 73 16312
rect 129 16256 139 16312
rect 63 16200 139 16256
rect 63 16144 73 16200
rect 129 16144 139 16200
rect 63 16088 139 16144
rect 63 16032 73 16088
rect 129 16032 139 16088
rect 63 15976 139 16032
rect 63 15920 73 15976
rect 129 15920 139 15976
rect 63 15864 139 15920
rect 63 15808 73 15864
rect 129 15808 139 15864
rect 63 15752 139 15808
rect 63 15696 73 15752
rect 129 15696 139 15752
rect 63 15640 139 15696
rect 63 15584 73 15640
rect 129 15584 139 15640
rect 63 15528 139 15584
rect 63 15472 73 15528
rect 129 15472 139 15528
rect 63 15416 139 15472
rect 63 15360 73 15416
rect 129 15360 139 15416
rect 63 15304 139 15360
rect 63 15248 73 15304
rect 129 15248 139 15304
rect 63 15192 139 15248
rect 63 15136 73 15192
rect 129 15136 139 15192
rect 63 15080 139 15136
rect 63 15024 73 15080
rect 129 15024 139 15080
rect 63 14968 139 15024
rect 63 14912 73 14968
rect 129 14912 139 14968
rect 63 14856 139 14912
rect 63 14800 73 14856
rect 129 14800 139 14856
rect 63 14744 139 14800
rect 63 14688 73 14744
rect 129 14688 139 14744
rect 63 14632 139 14688
rect 63 14576 73 14632
rect 129 14576 139 14632
rect 63 14520 139 14576
rect 63 14464 73 14520
rect 129 14464 139 14520
rect 63 14408 139 14464
rect 63 14352 73 14408
rect 129 14352 139 14408
rect 63 14296 139 14352
rect 63 14240 73 14296
rect 129 14240 139 14296
rect 63 14184 139 14240
rect 63 14128 73 14184
rect 129 14128 139 14184
rect 63 14118 139 14128
<< via3 >>
rect 73 69569 129 69625
rect 73 69457 129 69513
rect 73 69345 129 69401
rect 73 69233 129 69289
rect 73 69121 129 69177
rect 73 69009 129 69065
rect 73 68897 129 68953
rect 73 68785 129 68841
rect 73 68673 129 68729
rect 73 68561 129 68617
rect 73 68449 129 68505
rect 73 68097 129 68153
rect 73 67985 129 68041
rect 73 67873 129 67929
rect 73 67761 129 67817
rect 73 67649 129 67705
rect 73 67537 129 67593
rect 73 67425 129 67481
rect 73 67313 129 67369
rect 73 67201 129 67257
rect 73 67089 129 67145
rect 73 66977 129 67033
rect 73 66865 129 66921
rect 73 66496 129 66552
rect 73 66384 129 66440
rect 73 66272 129 66328
rect 73 66160 129 66216
rect 73 66048 129 66104
rect 73 65936 129 65992
rect 73 65824 129 65880
rect 73 65712 129 65768
rect 73 65600 129 65656
rect 73 65488 129 65544
rect 73 65376 129 65432
rect 73 65264 129 65320
rect 73 64888 129 64944
rect 73 64776 129 64832
rect 73 64664 129 64720
rect 73 64552 129 64608
rect 73 64440 129 64496
rect 73 64328 129 64384
rect 73 64216 129 64272
rect 73 64104 129 64160
rect 73 63992 129 64048
rect 73 63880 129 63936
rect 73 63768 129 63824
rect 73 63656 129 63712
rect 73 63288 129 63344
rect 73 63176 129 63232
rect 73 63064 129 63120
rect 73 62952 129 63008
rect 73 62840 129 62896
rect 73 62728 129 62784
rect 73 62616 129 62672
rect 73 62504 129 62560
rect 73 62392 129 62448
rect 73 62280 129 62336
rect 73 62168 129 62224
rect 73 62056 129 62112
rect 73 61689 129 61745
rect 73 61577 129 61633
rect 73 61465 129 61521
rect 73 61353 129 61409
rect 73 61241 129 61297
rect 73 61129 129 61185
rect 73 61017 129 61073
rect 73 60905 129 60961
rect 73 60793 129 60849
rect 73 60681 129 60737
rect 73 60569 129 60625
rect 73 60457 129 60513
rect 73 60096 129 60152
rect 73 59984 129 60040
rect 73 59872 129 59928
rect 73 59760 129 59816
rect 73 59648 129 59704
rect 73 59536 129 59592
rect 73 59424 129 59480
rect 73 59312 129 59368
rect 73 59200 129 59256
rect 73 59088 129 59144
rect 73 58976 129 59032
rect 73 58864 129 58920
rect 73 58491 129 58547
rect 73 58379 129 58435
rect 73 58267 129 58323
rect 73 58155 129 58211
rect 73 58043 129 58099
rect 73 57931 129 57987
rect 73 57819 129 57875
rect 73 57707 129 57763
rect 73 57595 129 57651
rect 73 57483 129 57539
rect 73 57371 129 57427
rect 73 57259 129 57315
rect 73 56893 129 56949
rect 73 56781 129 56837
rect 73 56669 129 56725
rect 73 56557 129 56613
rect 73 56445 129 56501
rect 73 56333 129 56389
rect 73 56221 129 56277
rect 73 56109 129 56165
rect 73 55997 129 56053
rect 73 55885 129 55941
rect 73 55773 129 55829
rect 73 55661 129 55717
rect 73 55292 129 55348
rect 73 55180 129 55236
rect 73 55068 129 55124
rect 73 54956 129 55012
rect 73 54844 129 54900
rect 73 54732 129 54788
rect 73 54620 129 54676
rect 73 54508 129 54564
rect 73 54396 129 54452
rect 73 54284 129 54340
rect 73 54172 129 54228
rect 73 54060 129 54116
rect 73 53679 129 53735
rect 73 53567 129 53623
rect 73 53455 129 53511
rect 73 53343 129 53399
rect 73 53231 129 53287
rect 73 53119 129 53175
rect 73 53007 129 53063
rect 73 52895 129 52951
rect 73 52783 129 52839
rect 73 52671 129 52727
rect 73 52559 129 52615
rect 73 52447 129 52503
rect 73 52093 129 52149
rect 73 51981 129 52037
rect 73 51869 129 51925
rect 73 51757 129 51813
rect 73 51645 129 51701
rect 73 51533 129 51589
rect 73 51421 129 51477
rect 73 51309 129 51365
rect 73 51197 129 51253
rect 73 51085 129 51141
rect 73 50973 129 51029
rect 73 50861 129 50917
rect 74 50482 130 50538
rect 74 50370 130 50426
rect 74 50258 130 50314
rect 74 50146 130 50202
rect 74 50034 130 50090
rect 74 49922 130 49978
rect 74 49810 130 49866
rect 74 49698 130 49754
rect 74 49586 130 49642
rect 74 49474 130 49530
rect 74 49362 130 49418
rect 74 49250 130 49306
rect 73 48828 129 48884
rect 73 48716 129 48772
rect 73 48604 129 48660
rect 73 48492 129 48548
rect 73 48380 129 48436
rect 73 48268 129 48324
rect 73 48156 129 48212
rect 73 48044 129 48100
rect 73 47932 129 47988
rect 73 47820 129 47876
rect 73 47708 129 47764
rect 73 47596 129 47652
rect 73 47484 129 47540
rect 73 47372 129 47428
rect 73 47260 129 47316
rect 73 47148 129 47204
rect 73 47036 129 47092
rect 73 46924 129 46980
rect 73 46812 129 46868
rect 73 46700 129 46756
rect 73 46588 129 46644
rect 73 46476 129 46532
rect 73 46364 129 46420
rect 73 46252 129 46308
rect 73 46140 129 46196
rect 73 45614 129 45670
rect 73 45502 129 45558
rect 73 45390 129 45446
rect 73 45278 129 45334
rect 73 45166 129 45222
rect 73 45054 129 45110
rect 73 44942 129 44998
rect 73 44830 129 44886
rect 73 44718 129 44774
rect 73 44606 129 44662
rect 73 44494 129 44550
rect 73 44382 129 44438
rect 73 44270 129 44326
rect 73 44158 129 44214
rect 73 44046 129 44102
rect 73 43934 129 43990
rect 73 43822 129 43878
rect 73 43710 129 43766
rect 73 43598 129 43654
rect 73 43486 129 43542
rect 73 43374 129 43430
rect 73 43262 129 43318
rect 73 43150 129 43206
rect 73 43038 129 43094
rect 73 42926 129 42982
rect 74 42493 130 42549
rect 74 42381 130 42437
rect 74 42269 130 42325
rect 74 42157 130 42213
rect 74 42045 130 42101
rect 74 41933 130 41989
rect 74 41821 130 41877
rect 74 41709 130 41765
rect 74 41597 130 41653
rect 74 41485 130 41541
rect 74 41373 130 41429
rect 74 41261 130 41317
rect 74 40895 130 40951
rect 74 40783 130 40839
rect 74 40671 130 40727
rect 74 40559 130 40615
rect 74 40447 130 40503
rect 74 40335 130 40391
rect 74 40223 130 40279
rect 74 40111 130 40167
rect 74 39999 130 40055
rect 74 39887 130 39943
rect 74 39775 130 39831
rect 74 39663 130 39719
rect 73 39220 129 39276
rect 73 39108 129 39164
rect 73 38996 129 39052
rect 73 38884 129 38940
rect 73 38772 129 38828
rect 73 38660 129 38716
rect 73 38548 129 38604
rect 73 38436 129 38492
rect 73 38324 129 38380
rect 73 38212 129 38268
rect 73 38100 129 38156
rect 73 37988 129 38044
rect 73 37876 129 37932
rect 73 37764 129 37820
rect 73 37652 129 37708
rect 73 37540 129 37596
rect 73 37428 129 37484
rect 73 37316 129 37372
rect 73 37204 129 37260
rect 73 37092 129 37148
rect 73 36980 129 37036
rect 73 36868 129 36924
rect 73 36756 129 36812
rect 73 36644 129 36700
rect 73 36532 129 36588
rect 73 36019 129 36075
rect 73 35907 129 35963
rect 73 35795 129 35851
rect 73 35683 129 35739
rect 73 35571 129 35627
rect 73 35459 129 35515
rect 73 35347 129 35403
rect 73 35235 129 35291
rect 73 35123 129 35179
rect 73 35011 129 35067
rect 73 34899 129 34955
rect 73 34787 129 34843
rect 73 34675 129 34731
rect 73 34563 129 34619
rect 73 34451 129 34507
rect 73 34339 129 34395
rect 73 34227 129 34283
rect 73 34115 129 34171
rect 73 34003 129 34059
rect 73 33891 129 33947
rect 73 33779 129 33835
rect 73 33667 129 33723
rect 73 33555 129 33611
rect 73 33443 129 33499
rect 73 33331 129 33387
rect 73 32823 129 32879
rect 73 32711 129 32767
rect 73 32599 129 32655
rect 73 32487 129 32543
rect 73 32375 129 32431
rect 73 32263 129 32319
rect 73 32151 129 32207
rect 73 32039 129 32095
rect 73 31927 129 31983
rect 73 31815 129 31871
rect 73 31703 129 31759
rect 73 31591 129 31647
rect 73 31479 129 31535
rect 73 31367 129 31423
rect 73 31255 129 31311
rect 73 31143 129 31199
rect 73 31031 129 31087
rect 73 30919 129 30975
rect 73 30807 129 30863
rect 73 30695 129 30751
rect 73 30583 129 30639
rect 73 30471 129 30527
rect 73 30359 129 30415
rect 73 30247 129 30303
rect 73 30135 129 30191
rect 73 29629 129 29685
rect 73 29517 129 29573
rect 73 29405 129 29461
rect 73 29293 129 29349
rect 73 29181 129 29237
rect 73 29069 129 29125
rect 73 28957 129 29013
rect 73 28845 129 28901
rect 73 28733 129 28789
rect 73 28621 129 28677
rect 73 28509 129 28565
rect 73 28397 129 28453
rect 73 28285 129 28341
rect 73 28173 129 28229
rect 73 28061 129 28117
rect 73 27949 129 28005
rect 73 27837 129 27893
rect 73 27725 129 27781
rect 73 27613 129 27669
rect 73 27501 129 27557
rect 73 27389 129 27445
rect 73 27277 129 27333
rect 73 27165 129 27221
rect 73 27053 129 27109
rect 73 26941 129 26997
rect 74 26494 130 26550
rect 74 26382 130 26438
rect 74 26270 130 26326
rect 74 26158 130 26214
rect 74 26046 130 26102
rect 74 25934 130 25990
rect 74 25822 130 25878
rect 74 25710 130 25766
rect 74 25598 130 25654
rect 74 25486 130 25542
rect 74 25374 130 25430
rect 74 25262 130 25318
rect 74 24901 130 24957
rect 74 24789 130 24845
rect 74 24677 130 24733
rect 74 24565 130 24621
rect 74 24453 130 24509
rect 74 24341 130 24397
rect 74 24229 130 24285
rect 74 24117 130 24173
rect 74 24005 130 24061
rect 74 23893 130 23949
rect 74 23781 130 23837
rect 74 23669 130 23725
rect 73 23267 129 23323
rect 73 23155 129 23211
rect 73 23043 129 23099
rect 73 22931 129 22987
rect 73 22819 129 22875
rect 73 22707 129 22763
rect 73 22595 129 22651
rect 73 22483 129 22539
rect 73 22371 129 22427
rect 73 22259 129 22315
rect 73 22147 129 22203
rect 73 22035 129 22091
rect 73 21923 129 21979
rect 73 21811 129 21867
rect 73 21699 129 21755
rect 73 21587 129 21643
rect 73 21475 129 21531
rect 73 21363 129 21419
rect 73 21251 129 21307
rect 73 21139 129 21195
rect 73 21027 129 21083
rect 73 20915 129 20971
rect 73 20803 129 20859
rect 73 20691 129 20747
rect 73 20579 129 20635
rect 73 20017 129 20073
rect 73 19905 129 19961
rect 73 19793 129 19849
rect 73 19681 129 19737
rect 73 19569 129 19625
rect 73 19457 129 19513
rect 73 19345 129 19401
rect 73 19233 129 19289
rect 73 19121 129 19177
rect 73 19009 129 19065
rect 73 18897 129 18953
rect 73 18785 129 18841
rect 73 18673 129 18729
rect 73 18561 129 18617
rect 73 18449 129 18505
rect 73 18337 129 18393
rect 73 18225 129 18281
rect 73 18113 129 18169
rect 73 18001 129 18057
rect 73 17889 129 17945
rect 73 17777 129 17833
rect 73 17665 129 17721
rect 73 17553 129 17609
rect 73 17441 129 17497
rect 73 17329 129 17385
rect 73 16816 129 16872
rect 73 16704 129 16760
rect 73 16592 129 16648
rect 73 16480 129 16536
rect 73 16368 129 16424
rect 73 16256 129 16312
rect 73 16144 129 16200
rect 73 16032 129 16088
rect 73 15920 129 15976
rect 73 15808 129 15864
rect 73 15696 129 15752
rect 73 15584 129 15640
rect 73 15472 129 15528
rect 73 15360 129 15416
rect 73 15248 129 15304
rect 73 15136 129 15192
rect 73 15024 129 15080
rect 73 14912 129 14968
rect 73 14800 129 14856
rect 73 14688 129 14744
rect 73 14576 129 14632
rect 73 14464 129 14520
rect 73 14352 129 14408
rect 73 14240 129 14296
rect 73 14128 129 14184
<< metal4 >>
rect 0 69625 200 69678
rect 0 69569 73 69625
rect 129 69569 200 69625
rect 0 69513 200 69569
rect 0 69457 73 69513
rect 129 69457 200 69513
rect 0 69401 200 69457
rect 0 69345 73 69401
rect 129 69345 200 69401
rect 0 69289 200 69345
rect 0 69233 73 69289
rect 129 69233 200 69289
rect 0 69177 200 69233
rect 0 69121 73 69177
rect 129 69121 200 69177
rect 0 69065 200 69121
rect 0 69009 73 69065
rect 129 69009 200 69065
rect 0 68953 200 69009
rect 0 68897 73 68953
rect 129 68897 200 68953
rect 0 68841 200 68897
rect 0 68785 73 68841
rect 129 68785 200 68841
rect 0 68729 200 68785
rect 0 68673 73 68729
rect 129 68673 200 68729
rect 0 68617 200 68673
rect 0 68561 73 68617
rect 129 68561 200 68617
rect 0 68505 200 68561
rect 0 68449 73 68505
rect 129 68449 200 68505
rect 0 68400 200 68449
rect 0 68153 200 68200
rect 0 68097 73 68153
rect 129 68097 200 68153
rect 0 68041 200 68097
rect 0 67985 73 68041
rect 129 67985 200 68041
rect 0 67929 200 67985
rect 0 67873 73 67929
rect 129 67873 200 67929
rect 0 67817 200 67873
rect 0 67761 73 67817
rect 129 67761 200 67817
rect 0 67705 200 67761
rect 0 67649 73 67705
rect 129 67649 200 67705
rect 0 67593 200 67649
rect 0 67537 73 67593
rect 129 67537 200 67593
rect 0 67481 200 67537
rect 0 67425 73 67481
rect 129 67425 200 67481
rect 0 67369 200 67425
rect 0 67313 73 67369
rect 129 67313 200 67369
rect 0 67257 200 67313
rect 0 67201 73 67257
rect 129 67201 200 67257
rect 0 67145 200 67201
rect 0 67089 73 67145
rect 129 67089 200 67145
rect 0 67033 200 67089
rect 0 66977 73 67033
rect 129 66977 200 67033
rect 0 66921 200 66977
rect 0 66865 73 66921
rect 129 66865 200 66921
rect 0 66800 200 66865
rect 0 66552 200 66600
rect 0 66496 73 66552
rect 129 66496 200 66552
rect 0 66440 200 66496
rect 0 66384 73 66440
rect 129 66384 200 66440
rect 0 66328 200 66384
rect 0 66272 73 66328
rect 129 66272 200 66328
rect 0 66216 200 66272
rect 0 66160 73 66216
rect 129 66160 200 66216
rect 0 66104 200 66160
rect 0 66048 73 66104
rect 129 66048 200 66104
rect 0 65992 200 66048
rect 0 65936 73 65992
rect 129 65936 200 65992
rect 0 65880 200 65936
rect 0 65824 73 65880
rect 129 65824 200 65880
rect 0 65768 200 65824
rect 0 65712 73 65768
rect 129 65712 200 65768
rect 0 65656 200 65712
rect 0 65600 73 65656
rect 129 65600 200 65656
rect 0 65544 200 65600
rect 0 65488 73 65544
rect 129 65488 200 65544
rect 0 65432 200 65488
rect 0 65376 73 65432
rect 129 65376 200 65432
rect 0 65320 200 65376
rect 0 65264 73 65320
rect 129 65264 200 65320
rect 0 65200 200 65264
rect 0 64944 200 65000
rect 0 64888 73 64944
rect 129 64888 200 64944
rect 0 64832 200 64888
rect 0 64776 73 64832
rect 129 64776 200 64832
rect 0 64720 200 64776
rect 0 64664 73 64720
rect 129 64664 200 64720
rect 0 64608 200 64664
rect 0 64552 73 64608
rect 129 64552 200 64608
rect 0 64496 200 64552
rect 0 64440 73 64496
rect 129 64440 200 64496
rect 0 64384 200 64440
rect 0 64328 73 64384
rect 129 64328 200 64384
rect 0 64272 200 64328
rect 0 64216 73 64272
rect 129 64216 200 64272
rect 0 64160 200 64216
rect 0 64104 73 64160
rect 129 64104 200 64160
rect 0 64048 200 64104
rect 0 63992 73 64048
rect 129 63992 200 64048
rect 0 63936 200 63992
rect 0 63880 73 63936
rect 129 63880 200 63936
rect 0 63824 200 63880
rect 0 63768 73 63824
rect 129 63768 200 63824
rect 0 63712 200 63768
rect 0 63656 73 63712
rect 129 63656 200 63712
rect 0 63600 200 63656
rect 0 63344 200 63400
rect 0 63288 73 63344
rect 129 63288 200 63344
rect 0 63232 200 63288
rect 0 63176 73 63232
rect 129 63176 200 63232
rect 0 63120 200 63176
rect 0 63064 73 63120
rect 129 63064 200 63120
rect 0 63008 200 63064
rect 0 62952 73 63008
rect 129 62952 200 63008
rect 0 62896 200 62952
rect 0 62840 73 62896
rect 129 62840 200 62896
rect 0 62784 200 62840
rect 0 62728 73 62784
rect 129 62728 200 62784
rect 0 62672 200 62728
rect 0 62616 73 62672
rect 129 62616 200 62672
rect 0 62560 200 62616
rect 0 62504 73 62560
rect 129 62504 200 62560
rect 0 62448 200 62504
rect 0 62392 73 62448
rect 129 62392 200 62448
rect 0 62336 200 62392
rect 0 62280 73 62336
rect 129 62280 200 62336
rect 0 62224 200 62280
rect 0 62168 73 62224
rect 129 62168 200 62224
rect 0 62112 200 62168
rect 0 62056 73 62112
rect 129 62056 200 62112
rect 0 62000 200 62056
rect 0 61745 200 61800
rect 0 61689 73 61745
rect 129 61689 200 61745
rect 0 61633 200 61689
rect 0 61577 73 61633
rect 129 61577 200 61633
rect 0 61521 200 61577
rect 0 61465 73 61521
rect 129 61465 200 61521
rect 0 61409 200 61465
rect 0 61353 73 61409
rect 129 61353 200 61409
rect 0 61297 200 61353
rect 0 61241 73 61297
rect 129 61241 200 61297
rect 0 61185 200 61241
rect 0 61129 73 61185
rect 129 61129 200 61185
rect 0 61073 200 61129
rect 0 61017 73 61073
rect 129 61017 200 61073
rect 0 60961 200 61017
rect 0 60905 73 60961
rect 129 60905 200 60961
rect 0 60849 200 60905
rect 0 60793 73 60849
rect 129 60793 200 60849
rect 0 60737 200 60793
rect 0 60681 73 60737
rect 129 60681 200 60737
rect 0 60625 200 60681
rect 0 60569 73 60625
rect 129 60569 200 60625
rect 0 60513 200 60569
rect 0 60457 73 60513
rect 129 60457 200 60513
rect 0 60400 200 60457
rect 0 60152 200 60200
rect 0 60096 73 60152
rect 129 60096 200 60152
rect 0 60040 200 60096
rect 0 59984 73 60040
rect 129 59984 200 60040
rect 0 59928 200 59984
rect 0 59872 73 59928
rect 129 59872 200 59928
rect 0 59816 200 59872
rect 0 59760 73 59816
rect 129 59760 200 59816
rect 0 59704 200 59760
rect 0 59648 73 59704
rect 129 59648 200 59704
rect 0 59592 200 59648
rect 0 59536 73 59592
rect 129 59536 200 59592
rect 0 59480 200 59536
rect 0 59424 73 59480
rect 129 59424 200 59480
rect 0 59368 200 59424
rect 0 59312 73 59368
rect 129 59312 200 59368
rect 0 59256 200 59312
rect 0 59200 73 59256
rect 129 59200 200 59256
rect 0 59144 200 59200
rect 0 59088 73 59144
rect 129 59088 200 59144
rect 0 59032 200 59088
rect 0 58976 73 59032
rect 129 58976 200 59032
rect 0 58920 200 58976
rect 0 58864 73 58920
rect 129 58864 200 58920
rect 0 58800 200 58864
rect 0 58547 200 58600
rect 0 58491 73 58547
rect 129 58491 200 58547
rect 0 58435 200 58491
rect 0 58379 73 58435
rect 129 58379 200 58435
rect 0 58323 200 58379
rect 0 58267 73 58323
rect 129 58267 200 58323
rect 0 58211 200 58267
rect 0 58155 73 58211
rect 129 58155 200 58211
rect 0 58099 200 58155
rect 0 58043 73 58099
rect 129 58043 200 58099
rect 0 57987 200 58043
rect 0 57931 73 57987
rect 129 57931 200 57987
rect 0 57875 200 57931
rect 0 57819 73 57875
rect 129 57819 200 57875
rect 0 57763 200 57819
rect 0 57707 73 57763
rect 129 57707 200 57763
rect 0 57651 200 57707
rect 0 57595 73 57651
rect 129 57595 200 57651
rect 0 57539 200 57595
rect 0 57483 73 57539
rect 129 57483 200 57539
rect 0 57427 200 57483
rect 0 57371 73 57427
rect 129 57371 200 57427
rect 0 57315 200 57371
rect 0 57259 73 57315
rect 129 57259 200 57315
rect 0 57200 200 57259
rect 0 56949 200 57000
rect 0 56893 73 56949
rect 129 56893 200 56949
rect 0 56837 200 56893
rect 0 56781 73 56837
rect 129 56781 200 56837
rect 0 56725 200 56781
rect 0 56669 73 56725
rect 129 56669 200 56725
rect 0 56613 200 56669
rect 0 56557 73 56613
rect 129 56557 200 56613
rect 0 56501 200 56557
rect 0 56445 73 56501
rect 129 56445 200 56501
rect 0 56389 200 56445
rect 0 56333 73 56389
rect 129 56333 200 56389
rect 0 56277 200 56333
rect 0 56221 73 56277
rect 129 56221 200 56277
rect 0 56165 200 56221
rect 0 56109 73 56165
rect 129 56109 200 56165
rect 0 56053 200 56109
rect 0 55997 73 56053
rect 129 55997 200 56053
rect 0 55941 200 55997
rect 0 55885 73 55941
rect 129 55885 200 55941
rect 0 55829 200 55885
rect 0 55773 73 55829
rect 129 55773 200 55829
rect 0 55717 200 55773
rect 0 55661 73 55717
rect 129 55661 200 55717
rect 0 55600 200 55661
rect 0 55348 200 55400
rect 0 55292 73 55348
rect 129 55292 200 55348
rect 0 55236 200 55292
rect 0 55180 73 55236
rect 129 55180 200 55236
rect 0 55124 200 55180
rect 0 55068 73 55124
rect 129 55068 200 55124
rect 0 55012 200 55068
rect 0 54956 73 55012
rect 129 54956 200 55012
rect 0 54900 200 54956
rect 0 54844 73 54900
rect 129 54844 200 54900
rect 0 54788 200 54844
rect 0 54732 73 54788
rect 129 54732 200 54788
rect 0 54676 200 54732
rect 0 54620 73 54676
rect 129 54620 200 54676
rect 0 54564 200 54620
rect 0 54508 73 54564
rect 129 54508 200 54564
rect 0 54452 200 54508
rect 0 54396 73 54452
rect 129 54396 200 54452
rect 0 54340 200 54396
rect 0 54284 73 54340
rect 129 54284 200 54340
rect 0 54228 200 54284
rect 0 54172 73 54228
rect 129 54172 200 54228
rect 0 54116 200 54172
rect 0 54060 73 54116
rect 129 54060 200 54116
rect 0 54000 200 54060
rect 0 53735 200 53800
rect 0 53679 73 53735
rect 129 53679 200 53735
rect 0 53623 200 53679
rect 0 53567 73 53623
rect 129 53567 200 53623
rect 0 53511 200 53567
rect 0 53455 73 53511
rect 129 53455 200 53511
rect 0 53399 200 53455
rect 0 53343 73 53399
rect 129 53343 200 53399
rect 0 53287 200 53343
rect 0 53231 73 53287
rect 129 53231 200 53287
rect 0 53175 200 53231
rect 0 53119 73 53175
rect 129 53119 200 53175
rect 0 53063 200 53119
rect 0 53007 73 53063
rect 129 53007 200 53063
rect 0 52951 200 53007
rect 0 52895 73 52951
rect 129 52895 200 52951
rect 0 52839 200 52895
rect 0 52783 73 52839
rect 129 52783 200 52839
rect 0 52727 200 52783
rect 0 52671 73 52727
rect 129 52671 200 52727
rect 0 52615 200 52671
rect 0 52559 73 52615
rect 129 52559 200 52615
rect 0 52503 200 52559
rect 0 52447 73 52503
rect 129 52447 200 52503
rect 0 52400 200 52447
rect 0 52149 200 52200
rect 0 52093 73 52149
rect 129 52093 200 52149
rect 0 52037 200 52093
rect 0 51981 73 52037
rect 129 51981 200 52037
rect 0 51925 200 51981
rect 0 51869 73 51925
rect 129 51869 200 51925
rect 0 51813 200 51869
rect 0 51757 73 51813
rect 129 51757 200 51813
rect 0 51701 200 51757
rect 0 51645 73 51701
rect 129 51645 200 51701
rect 0 51589 200 51645
rect 0 51533 73 51589
rect 129 51533 200 51589
rect 0 51477 200 51533
rect 0 51421 73 51477
rect 129 51421 200 51477
rect 0 51365 200 51421
rect 0 51309 73 51365
rect 129 51309 200 51365
rect 0 51253 200 51309
rect 0 51197 73 51253
rect 129 51197 200 51253
rect 0 51141 200 51197
rect 0 51085 73 51141
rect 129 51085 200 51141
rect 0 51029 200 51085
rect 0 50973 73 51029
rect 129 50973 200 51029
rect 0 50917 200 50973
rect 0 50861 73 50917
rect 129 50861 200 50917
rect 0 50800 200 50861
rect 0 50538 200 50600
rect 0 50482 74 50538
rect 130 50482 200 50538
rect 0 50426 200 50482
rect 0 50370 74 50426
rect 130 50370 200 50426
rect 0 50314 200 50370
rect 0 50258 74 50314
rect 130 50258 200 50314
rect 0 50202 200 50258
rect 0 50146 74 50202
rect 130 50146 200 50202
rect 0 50090 200 50146
rect 0 50034 74 50090
rect 130 50034 200 50090
rect 0 49978 200 50034
rect 0 49922 74 49978
rect 130 49922 200 49978
rect 0 49866 200 49922
rect 0 49810 74 49866
rect 130 49810 200 49866
rect 0 49754 200 49810
rect 0 49698 74 49754
rect 130 49698 200 49754
rect 0 49642 200 49698
rect 0 49586 74 49642
rect 130 49586 200 49642
rect 0 49530 200 49586
rect 0 49474 74 49530
rect 130 49474 200 49530
rect 0 49418 200 49474
rect 0 49362 74 49418
rect 130 49362 200 49418
rect 0 49306 200 49362
rect 0 49250 74 49306
rect 130 49250 200 49306
rect 0 49200 200 49250
rect 0 48884 200 49000
rect 0 48828 73 48884
rect 129 48828 200 48884
rect 0 48772 200 48828
rect 0 48716 73 48772
rect 129 48716 200 48772
rect 0 48660 200 48716
rect 0 48604 73 48660
rect 129 48604 200 48660
rect 0 48548 200 48604
rect 0 48492 73 48548
rect 129 48492 200 48548
rect 0 48436 200 48492
rect 0 48380 73 48436
rect 129 48380 200 48436
rect 0 48324 200 48380
rect 0 48268 73 48324
rect 129 48268 200 48324
rect 0 48212 200 48268
rect 0 48156 73 48212
rect 129 48156 200 48212
rect 0 48100 200 48156
rect 0 48044 73 48100
rect 129 48044 200 48100
rect 0 47988 200 48044
rect 0 47932 73 47988
rect 129 47932 200 47988
rect 0 47876 200 47932
rect 0 47820 73 47876
rect 129 47820 200 47876
rect 0 47764 200 47820
rect 0 47708 73 47764
rect 129 47708 200 47764
rect 0 47652 200 47708
rect 0 47596 73 47652
rect 129 47596 200 47652
rect 0 47540 200 47596
rect 0 47484 73 47540
rect 129 47484 200 47540
rect 0 47428 200 47484
rect 0 47372 73 47428
rect 129 47372 200 47428
rect 0 47316 200 47372
rect 0 47260 73 47316
rect 129 47260 200 47316
rect 0 47204 200 47260
rect 0 47148 73 47204
rect 129 47148 200 47204
rect 0 47092 200 47148
rect 0 47036 73 47092
rect 129 47036 200 47092
rect 0 46980 200 47036
rect 0 46924 73 46980
rect 129 46924 200 46980
rect 0 46868 200 46924
rect 0 46812 73 46868
rect 129 46812 200 46868
rect 0 46756 200 46812
rect 0 46700 73 46756
rect 129 46700 200 46756
rect 0 46644 200 46700
rect 0 46588 73 46644
rect 129 46588 200 46644
rect 0 46532 200 46588
rect 0 46476 73 46532
rect 129 46476 200 46532
rect 0 46420 200 46476
rect 0 46364 73 46420
rect 129 46364 200 46420
rect 0 46308 200 46364
rect 0 46252 73 46308
rect 129 46252 200 46308
rect 0 46196 200 46252
rect 0 46140 73 46196
rect 129 46140 200 46196
rect 0 46000 200 46140
rect 0 45670 200 45800
rect 0 45614 73 45670
rect 129 45614 200 45670
rect 0 45558 200 45614
rect 0 45502 73 45558
rect 129 45502 200 45558
rect 0 45446 200 45502
rect 0 45390 73 45446
rect 129 45390 200 45446
rect 0 45334 200 45390
rect 0 45278 73 45334
rect 129 45278 200 45334
rect 0 45222 200 45278
rect 0 45166 73 45222
rect 129 45166 200 45222
rect 0 45110 200 45166
rect 0 45054 73 45110
rect 129 45054 200 45110
rect 0 44998 200 45054
rect 0 44942 73 44998
rect 129 44942 200 44998
rect 0 44886 200 44942
rect 0 44830 73 44886
rect 129 44830 200 44886
rect 0 44774 200 44830
rect 0 44718 73 44774
rect 129 44718 200 44774
rect 0 44662 200 44718
rect 0 44606 73 44662
rect 129 44606 200 44662
rect 0 44550 200 44606
rect 0 44494 73 44550
rect 129 44494 200 44550
rect 0 44438 200 44494
rect 0 44382 73 44438
rect 129 44382 200 44438
rect 0 44326 200 44382
rect 0 44270 73 44326
rect 129 44270 200 44326
rect 0 44214 200 44270
rect 0 44158 73 44214
rect 129 44158 200 44214
rect 0 44102 200 44158
rect 0 44046 73 44102
rect 129 44046 200 44102
rect 0 43990 200 44046
rect 0 43934 73 43990
rect 129 43934 200 43990
rect 0 43878 200 43934
rect 0 43822 73 43878
rect 129 43822 200 43878
rect 0 43766 200 43822
rect 0 43710 73 43766
rect 129 43710 200 43766
rect 0 43654 200 43710
rect 0 43598 73 43654
rect 129 43598 200 43654
rect 0 43542 200 43598
rect 0 43486 73 43542
rect 129 43486 200 43542
rect 0 43430 200 43486
rect 0 43374 73 43430
rect 129 43374 200 43430
rect 0 43318 200 43374
rect 0 43262 73 43318
rect 129 43262 200 43318
rect 0 43206 200 43262
rect 0 43150 73 43206
rect 129 43150 200 43206
rect 0 43094 200 43150
rect 0 43038 73 43094
rect 129 43038 200 43094
rect 0 42982 200 43038
rect 0 42926 73 42982
rect 129 42926 200 42982
rect 0 42800 200 42926
rect 0 42549 200 42600
rect 0 42493 74 42549
rect 130 42493 200 42549
rect 0 42437 200 42493
rect 0 42381 74 42437
rect 130 42381 200 42437
rect 0 42325 200 42381
rect 0 42269 74 42325
rect 130 42269 200 42325
rect 0 42213 200 42269
rect 0 42157 74 42213
rect 130 42157 200 42213
rect 0 42101 200 42157
rect 0 42045 74 42101
rect 130 42045 200 42101
rect 0 41989 200 42045
rect 0 41933 74 41989
rect 130 41933 200 41989
rect 0 41877 200 41933
rect 0 41821 74 41877
rect 130 41821 200 41877
rect 0 41765 200 41821
rect 0 41709 74 41765
rect 130 41709 200 41765
rect 0 41653 200 41709
rect 0 41597 74 41653
rect 130 41597 200 41653
rect 0 41541 200 41597
rect 0 41485 74 41541
rect 130 41485 200 41541
rect 0 41429 200 41485
rect 0 41373 74 41429
rect 130 41373 200 41429
rect 0 41317 200 41373
rect 0 41261 74 41317
rect 130 41261 200 41317
rect 0 41200 200 41261
rect 0 40951 200 41000
rect 0 40895 74 40951
rect 130 40895 200 40951
rect 0 40839 200 40895
rect 0 40783 74 40839
rect 130 40783 200 40839
rect 0 40727 200 40783
rect 0 40671 74 40727
rect 130 40671 200 40727
rect 0 40615 200 40671
rect 0 40559 74 40615
rect 130 40559 200 40615
rect 0 40503 200 40559
rect 0 40447 74 40503
rect 130 40447 200 40503
rect 0 40391 200 40447
rect 0 40335 74 40391
rect 130 40335 200 40391
rect 0 40279 200 40335
rect 0 40223 74 40279
rect 130 40223 200 40279
rect 0 40167 200 40223
rect 0 40111 74 40167
rect 130 40111 200 40167
rect 0 40055 200 40111
rect 0 39999 74 40055
rect 130 39999 200 40055
rect 0 39943 200 39999
rect 0 39887 74 39943
rect 130 39887 200 39943
rect 0 39831 200 39887
rect 0 39775 74 39831
rect 130 39775 200 39831
rect 0 39719 200 39775
rect 0 39663 74 39719
rect 130 39663 200 39719
rect 0 39600 200 39663
rect 0 39276 200 39400
rect 0 39220 73 39276
rect 129 39220 200 39276
rect 0 39164 200 39220
rect 0 39108 73 39164
rect 129 39108 200 39164
rect 0 39052 200 39108
rect 0 38996 73 39052
rect 129 38996 200 39052
rect 0 38940 200 38996
rect 0 38884 73 38940
rect 129 38884 200 38940
rect 0 38828 200 38884
rect 0 38772 73 38828
rect 129 38772 200 38828
rect 0 38716 200 38772
rect 0 38660 73 38716
rect 129 38660 200 38716
rect 0 38604 200 38660
rect 0 38548 73 38604
rect 129 38548 200 38604
rect 0 38492 200 38548
rect 0 38436 73 38492
rect 129 38436 200 38492
rect 0 38380 200 38436
rect 0 38324 73 38380
rect 129 38324 200 38380
rect 0 38268 200 38324
rect 0 38212 73 38268
rect 129 38212 200 38268
rect 0 38156 200 38212
rect 0 38100 73 38156
rect 129 38100 200 38156
rect 0 38044 200 38100
rect 0 37988 73 38044
rect 129 37988 200 38044
rect 0 37932 200 37988
rect 0 37876 73 37932
rect 129 37876 200 37932
rect 0 37820 200 37876
rect 0 37764 73 37820
rect 129 37764 200 37820
rect 0 37708 200 37764
rect 0 37652 73 37708
rect 129 37652 200 37708
rect 0 37596 200 37652
rect 0 37540 73 37596
rect 129 37540 200 37596
rect 0 37484 200 37540
rect 0 37428 73 37484
rect 129 37428 200 37484
rect 0 37372 200 37428
rect 0 37316 73 37372
rect 129 37316 200 37372
rect 0 37260 200 37316
rect 0 37204 73 37260
rect 129 37204 200 37260
rect 0 37148 200 37204
rect 0 37092 73 37148
rect 129 37092 200 37148
rect 0 37036 200 37092
rect 0 36980 73 37036
rect 129 36980 200 37036
rect 0 36924 200 36980
rect 0 36868 73 36924
rect 129 36868 200 36924
rect 0 36812 200 36868
rect 0 36756 73 36812
rect 129 36756 200 36812
rect 0 36700 200 36756
rect 0 36644 73 36700
rect 129 36644 200 36700
rect 0 36588 200 36644
rect 0 36532 73 36588
rect 129 36532 200 36588
rect 0 36400 200 36532
rect 0 36075 200 36200
rect 0 36019 73 36075
rect 129 36019 200 36075
rect 0 35963 200 36019
rect 0 35907 73 35963
rect 129 35907 200 35963
rect 0 35851 200 35907
rect 0 35795 73 35851
rect 129 35795 200 35851
rect 0 35739 200 35795
rect 0 35683 73 35739
rect 129 35683 200 35739
rect 0 35627 200 35683
rect 0 35571 73 35627
rect 129 35571 200 35627
rect 0 35515 200 35571
rect 0 35459 73 35515
rect 129 35459 200 35515
rect 0 35403 200 35459
rect 0 35347 73 35403
rect 129 35347 200 35403
rect 0 35291 200 35347
rect 0 35235 73 35291
rect 129 35235 200 35291
rect 0 35179 200 35235
rect 0 35123 73 35179
rect 129 35123 200 35179
rect 0 35067 200 35123
rect 0 35011 73 35067
rect 129 35011 200 35067
rect 0 34955 200 35011
rect 0 34899 73 34955
rect 129 34899 200 34955
rect 0 34843 200 34899
rect 0 34787 73 34843
rect 129 34787 200 34843
rect 0 34731 200 34787
rect 0 34675 73 34731
rect 129 34675 200 34731
rect 0 34619 200 34675
rect 0 34563 73 34619
rect 129 34563 200 34619
rect 0 34507 200 34563
rect 0 34451 73 34507
rect 129 34451 200 34507
rect 0 34395 200 34451
rect 0 34339 73 34395
rect 129 34339 200 34395
rect 0 34283 200 34339
rect 0 34227 73 34283
rect 129 34227 200 34283
rect 0 34171 200 34227
rect 0 34115 73 34171
rect 129 34115 200 34171
rect 0 34059 200 34115
rect 0 34003 73 34059
rect 129 34003 200 34059
rect 0 33947 200 34003
rect 0 33891 73 33947
rect 129 33891 200 33947
rect 0 33835 200 33891
rect 0 33779 73 33835
rect 129 33779 200 33835
rect 0 33723 200 33779
rect 0 33667 73 33723
rect 129 33667 200 33723
rect 0 33611 200 33667
rect 0 33555 73 33611
rect 129 33555 200 33611
rect 0 33499 200 33555
rect 0 33443 73 33499
rect 129 33443 200 33499
rect 0 33387 200 33443
rect 0 33331 73 33387
rect 129 33331 200 33387
rect 0 33200 200 33331
rect 0 32879 200 33000
rect 0 32823 73 32879
rect 129 32823 200 32879
rect 0 32767 200 32823
rect 0 32711 73 32767
rect 129 32711 200 32767
rect 0 32655 200 32711
rect 0 32599 73 32655
rect 129 32599 200 32655
rect 0 32543 200 32599
rect 0 32487 73 32543
rect 129 32487 200 32543
rect 0 32431 200 32487
rect 0 32375 73 32431
rect 129 32375 200 32431
rect 0 32319 200 32375
rect 0 32263 73 32319
rect 129 32263 200 32319
rect 0 32207 200 32263
rect 0 32151 73 32207
rect 129 32151 200 32207
rect 0 32095 200 32151
rect 0 32039 73 32095
rect 129 32039 200 32095
rect 0 31983 200 32039
rect 0 31927 73 31983
rect 129 31927 200 31983
rect 0 31871 200 31927
rect 0 31815 73 31871
rect 129 31815 200 31871
rect 0 31759 200 31815
rect 0 31703 73 31759
rect 129 31703 200 31759
rect 0 31647 200 31703
rect 0 31591 73 31647
rect 129 31591 200 31647
rect 0 31535 200 31591
rect 0 31479 73 31535
rect 129 31479 200 31535
rect 0 31423 200 31479
rect 0 31367 73 31423
rect 129 31367 200 31423
rect 0 31311 200 31367
rect 0 31255 73 31311
rect 129 31255 200 31311
rect 0 31199 200 31255
rect 0 31143 73 31199
rect 129 31143 200 31199
rect 0 31087 200 31143
rect 0 31031 73 31087
rect 129 31031 200 31087
rect 0 30975 200 31031
rect 0 30919 73 30975
rect 129 30919 200 30975
rect 0 30863 200 30919
rect 0 30807 73 30863
rect 129 30807 200 30863
rect 0 30751 200 30807
rect 0 30695 73 30751
rect 129 30695 200 30751
rect 0 30639 200 30695
rect 0 30583 73 30639
rect 129 30583 200 30639
rect 0 30527 200 30583
rect 0 30471 73 30527
rect 129 30471 200 30527
rect 0 30415 200 30471
rect 0 30359 73 30415
rect 129 30359 200 30415
rect 0 30303 200 30359
rect 0 30247 73 30303
rect 129 30247 200 30303
rect 0 30191 200 30247
rect 0 30135 73 30191
rect 129 30135 200 30191
rect 0 30000 200 30135
rect 0 29685 200 29800
rect 0 29629 73 29685
rect 129 29629 200 29685
rect 0 29573 200 29629
rect 0 29517 73 29573
rect 129 29517 200 29573
rect 0 29461 200 29517
rect 0 29405 73 29461
rect 129 29405 200 29461
rect 0 29349 200 29405
rect 0 29293 73 29349
rect 129 29293 200 29349
rect 0 29237 200 29293
rect 0 29181 73 29237
rect 129 29181 200 29237
rect 0 29125 200 29181
rect 0 29069 73 29125
rect 129 29069 200 29125
rect 0 29013 200 29069
rect 0 28957 73 29013
rect 129 28957 200 29013
rect 0 28901 200 28957
rect 0 28845 73 28901
rect 129 28845 200 28901
rect 0 28789 200 28845
rect 0 28733 73 28789
rect 129 28733 200 28789
rect 0 28677 200 28733
rect 0 28621 73 28677
rect 129 28621 200 28677
rect 0 28565 200 28621
rect 0 28509 73 28565
rect 129 28509 200 28565
rect 0 28453 200 28509
rect 0 28397 73 28453
rect 129 28397 200 28453
rect 0 28341 200 28397
rect 0 28285 73 28341
rect 129 28285 200 28341
rect 0 28229 200 28285
rect 0 28173 73 28229
rect 129 28173 200 28229
rect 0 28117 200 28173
rect 0 28061 73 28117
rect 129 28061 200 28117
rect 0 28005 200 28061
rect 0 27949 73 28005
rect 129 27949 200 28005
rect 0 27893 200 27949
rect 0 27837 73 27893
rect 129 27837 200 27893
rect 0 27781 200 27837
rect 0 27725 73 27781
rect 129 27725 200 27781
rect 0 27669 200 27725
rect 0 27613 73 27669
rect 129 27613 200 27669
rect 0 27557 200 27613
rect 0 27501 73 27557
rect 129 27501 200 27557
rect 0 27445 200 27501
rect 0 27389 73 27445
rect 129 27389 200 27445
rect 0 27333 200 27389
rect 0 27277 73 27333
rect 129 27277 200 27333
rect 0 27221 200 27277
rect 0 27165 73 27221
rect 129 27165 200 27221
rect 0 27109 200 27165
rect 0 27053 73 27109
rect 129 27053 200 27109
rect 0 26997 200 27053
rect 0 26941 73 26997
rect 129 26941 200 26997
rect 0 26800 200 26941
rect 0 26550 200 26600
rect 0 26494 74 26550
rect 130 26494 200 26550
rect 0 26438 200 26494
rect 0 26382 74 26438
rect 130 26382 200 26438
rect 0 26326 200 26382
rect 0 26270 74 26326
rect 130 26270 200 26326
rect 0 26214 200 26270
rect 0 26158 74 26214
rect 130 26158 200 26214
rect 0 26102 200 26158
rect 0 26046 74 26102
rect 130 26046 200 26102
rect 0 25990 200 26046
rect 0 25934 74 25990
rect 130 25934 200 25990
rect 0 25878 200 25934
rect 0 25822 74 25878
rect 130 25822 200 25878
rect 0 25766 200 25822
rect 0 25710 74 25766
rect 130 25710 200 25766
rect 0 25654 200 25710
rect 0 25598 74 25654
rect 130 25598 200 25654
rect 0 25542 200 25598
rect 0 25486 74 25542
rect 130 25486 200 25542
rect 0 25430 200 25486
rect 0 25374 74 25430
rect 130 25374 200 25430
rect 0 25318 200 25374
rect 0 25262 74 25318
rect 130 25262 200 25318
rect 0 25200 200 25262
rect 0 24957 200 25000
rect 0 24901 74 24957
rect 130 24901 200 24957
rect 0 24845 200 24901
rect 0 24789 74 24845
rect 130 24789 200 24845
rect 0 24733 200 24789
rect 0 24677 74 24733
rect 130 24677 200 24733
rect 0 24621 200 24677
rect 0 24565 74 24621
rect 130 24565 200 24621
rect 0 24509 200 24565
rect 0 24453 74 24509
rect 130 24453 200 24509
rect 0 24397 200 24453
rect 0 24341 74 24397
rect 130 24341 200 24397
rect 0 24285 200 24341
rect 0 24229 74 24285
rect 130 24229 200 24285
rect 0 24173 200 24229
rect 0 24117 74 24173
rect 130 24117 200 24173
rect 0 24061 200 24117
rect 0 24005 74 24061
rect 130 24005 200 24061
rect 0 23949 200 24005
rect 0 23893 74 23949
rect 130 23893 200 23949
rect 0 23837 200 23893
rect 0 23781 74 23837
rect 130 23781 200 23837
rect 0 23725 200 23781
rect 0 23669 74 23725
rect 130 23669 200 23725
rect 0 23600 200 23669
rect 0 23323 200 23400
rect 0 23267 73 23323
rect 129 23267 200 23323
rect 0 23211 200 23267
rect 0 23155 73 23211
rect 129 23155 200 23211
rect 0 23099 200 23155
rect 0 23043 73 23099
rect 129 23043 200 23099
rect 0 22987 200 23043
rect 0 22931 73 22987
rect 129 22931 200 22987
rect 0 22875 200 22931
rect 0 22819 73 22875
rect 129 22819 200 22875
rect 0 22763 200 22819
rect 0 22707 73 22763
rect 129 22707 200 22763
rect 0 22651 200 22707
rect 0 22595 73 22651
rect 129 22595 200 22651
rect 0 22539 200 22595
rect 0 22483 73 22539
rect 129 22483 200 22539
rect 0 22427 200 22483
rect 0 22371 73 22427
rect 129 22371 200 22427
rect 0 22315 200 22371
rect 0 22259 73 22315
rect 129 22259 200 22315
rect 0 22203 200 22259
rect 0 22147 73 22203
rect 129 22147 200 22203
rect 0 22091 200 22147
rect 0 22035 73 22091
rect 129 22035 200 22091
rect 0 21979 200 22035
rect 0 21923 73 21979
rect 129 21923 200 21979
rect 0 21867 200 21923
rect 0 21811 73 21867
rect 129 21811 200 21867
rect 0 21755 200 21811
rect 0 21699 73 21755
rect 129 21699 200 21755
rect 0 21643 200 21699
rect 0 21587 73 21643
rect 129 21587 200 21643
rect 0 21531 200 21587
rect 0 21475 73 21531
rect 129 21475 200 21531
rect 0 21419 200 21475
rect 0 21363 73 21419
rect 129 21363 200 21419
rect 0 21307 200 21363
rect 0 21251 73 21307
rect 129 21251 200 21307
rect 0 21195 200 21251
rect 0 21139 73 21195
rect 129 21139 200 21195
rect 0 21083 200 21139
rect 0 21027 73 21083
rect 129 21027 200 21083
rect 0 20971 200 21027
rect 0 20915 73 20971
rect 129 20915 200 20971
rect 0 20859 200 20915
rect 0 20803 73 20859
rect 129 20803 200 20859
rect 0 20747 200 20803
rect 0 20691 73 20747
rect 129 20691 200 20747
rect 0 20635 200 20691
rect 0 20579 73 20635
rect 129 20579 200 20635
rect 0 20400 200 20579
rect 0 20073 200 20200
rect 0 20017 73 20073
rect 129 20017 200 20073
rect 0 19961 200 20017
rect 0 19905 73 19961
rect 129 19905 200 19961
rect 0 19849 200 19905
rect 0 19793 73 19849
rect 129 19793 200 19849
rect 0 19737 200 19793
rect 0 19681 73 19737
rect 129 19681 200 19737
rect 0 19625 200 19681
rect 0 19569 73 19625
rect 129 19569 200 19625
rect 0 19513 200 19569
rect 0 19457 73 19513
rect 129 19457 200 19513
rect 0 19401 200 19457
rect 0 19345 73 19401
rect 129 19345 200 19401
rect 0 19289 200 19345
rect 0 19233 73 19289
rect 129 19233 200 19289
rect 0 19177 200 19233
rect 0 19121 73 19177
rect 129 19121 200 19177
rect 0 19065 200 19121
rect 0 19009 73 19065
rect 129 19009 200 19065
rect 0 18953 200 19009
rect 0 18897 73 18953
rect 129 18897 200 18953
rect 0 18841 200 18897
rect 0 18785 73 18841
rect 129 18785 200 18841
rect 0 18729 200 18785
rect 0 18673 73 18729
rect 129 18673 200 18729
rect 0 18617 200 18673
rect 0 18561 73 18617
rect 129 18561 200 18617
rect 0 18505 200 18561
rect 0 18449 73 18505
rect 129 18449 200 18505
rect 0 18393 200 18449
rect 0 18337 73 18393
rect 129 18337 200 18393
rect 0 18281 200 18337
rect 0 18225 73 18281
rect 129 18225 200 18281
rect 0 18169 200 18225
rect 0 18113 73 18169
rect 129 18113 200 18169
rect 0 18057 200 18113
rect 0 18001 73 18057
rect 129 18001 200 18057
rect 0 17945 200 18001
rect 0 17889 73 17945
rect 129 17889 200 17945
rect 0 17833 200 17889
rect 0 17777 73 17833
rect 129 17777 200 17833
rect 0 17721 200 17777
rect 0 17665 73 17721
rect 129 17665 200 17721
rect 0 17609 200 17665
rect 0 17553 73 17609
rect 129 17553 200 17609
rect 0 17497 200 17553
rect 0 17441 73 17497
rect 129 17441 200 17497
rect 0 17385 200 17441
rect 0 17329 73 17385
rect 129 17329 200 17385
rect 0 17200 200 17329
rect 0 16872 200 17000
rect 0 16816 73 16872
rect 129 16816 200 16872
rect 0 16760 200 16816
rect 0 16704 73 16760
rect 129 16704 200 16760
rect 0 16648 200 16704
rect 0 16592 73 16648
rect 129 16592 200 16648
rect 0 16536 200 16592
rect 0 16480 73 16536
rect 129 16480 200 16536
rect 0 16424 200 16480
rect 0 16368 73 16424
rect 129 16368 200 16424
rect 0 16312 200 16368
rect 0 16256 73 16312
rect 129 16256 200 16312
rect 0 16200 200 16256
rect 0 16144 73 16200
rect 129 16144 200 16200
rect 0 16088 200 16144
rect 0 16032 73 16088
rect 129 16032 200 16088
rect 0 15976 200 16032
rect 0 15920 73 15976
rect 129 15920 200 15976
rect 0 15864 200 15920
rect 0 15808 73 15864
rect 129 15808 200 15864
rect 0 15752 200 15808
rect 0 15696 73 15752
rect 129 15696 200 15752
rect 0 15640 200 15696
rect 0 15584 73 15640
rect 129 15584 200 15640
rect 0 15528 200 15584
rect 0 15472 73 15528
rect 129 15472 200 15528
rect 0 15416 200 15472
rect 0 15360 73 15416
rect 129 15360 200 15416
rect 0 15304 200 15360
rect 0 15248 73 15304
rect 129 15248 200 15304
rect 0 15192 200 15248
rect 0 15136 73 15192
rect 129 15136 200 15192
rect 0 15080 200 15136
rect 0 15024 73 15080
rect 129 15024 200 15080
rect 0 14968 200 15024
rect 0 14912 73 14968
rect 129 14912 200 14968
rect 0 14856 200 14912
rect 0 14800 73 14856
rect 129 14800 200 14856
rect 0 14744 200 14800
rect 0 14688 73 14744
rect 129 14688 200 14744
rect 0 14632 200 14688
rect 0 14576 73 14632
rect 129 14576 200 14632
rect 0 14520 200 14576
rect 0 14464 73 14520
rect 129 14464 200 14520
rect 0 14408 200 14464
rect 0 14352 73 14408
rect 129 14352 200 14408
rect 0 14296 200 14352
rect 0 14240 73 14296
rect 129 14240 200 14296
rect 0 14184 200 14240
rect 0 14128 73 14184
rect 129 14128 200 14184
rect 0 14000 200 14128
use GF_NI_FILL1_1  GF_NI_FILL1_1_0
timestamp 1698431365
transform 1 0 0 0 1 0
box -32 13097 232 69968
use M4_M3_CDNS_4066195314522  M4_M3_CDNS_4066195314522_0
timestamp 1698431365
transform 1 0 101 0 1 56305
box 0 0 1 1
use M4_M3_CDNS_4066195314522  M4_M3_CDNS_4066195314522_1
timestamp 1698431365
transform 1 0 101 0 1 64300
box 0 0 1 1
use M4_M3_CDNS_4066195314522  M4_M3_CDNS_4066195314522_2
timestamp 1698431365
transform 1 0 101 0 1 65908
box 0 0 1 1
use M4_M3_CDNS_4066195314522  M4_M3_CDNS_4066195314522_3
timestamp 1698431365
transform 1 0 101 0 1 67509
box 0 0 1 1
use M4_M3_CDNS_4066195314522  M4_M3_CDNS_4066195314522_4
timestamp 1698431365
transform 1 0 101 0 1 62700
box 0 0 1 1
use M4_M3_CDNS_4066195314522  M4_M3_CDNS_4066195314522_5
timestamp 1698431365
transform 1 0 101 0 1 61101
box 0 0 1 1
use M4_M3_CDNS_4066195314522  M4_M3_CDNS_4066195314522_6
timestamp 1698431365
transform 1 0 101 0 1 59508
box 0 0 1 1
use M4_M3_CDNS_4066195314522  M4_M3_CDNS_4066195314522_7
timestamp 1698431365
transform 1 0 101 0 1 57903
box 0 0 1 1
use M4_M3_CDNS_4066195314522  M4_M3_CDNS_4066195314522_8
timestamp 1698431365
transform 1 0 101 0 1 54704
box 0 0 1 1
use M4_M3_CDNS_4066195314522  M4_M3_CDNS_4066195314522_9
timestamp 1698431365
transform 1 0 101 0 1 53091
box 0 0 1 1
use M4_M3_CDNS_4066195314522  M4_M3_CDNS_4066195314522_10
timestamp 1698431365
transform 1 0 101 0 1 51505
box 0 0 1 1
use M4_M3_CDNS_4066195314522  M4_M3_CDNS_4066195314522_11
timestamp 1698431365
transform 1 0 102 0 1 41905
box 0 0 1 1
use M4_M3_CDNS_4066195314522  M4_M3_CDNS_4066195314522_12
timestamp 1698431365
transform 1 0 102 0 1 40307
box 0 0 1 1
use M4_M3_CDNS_4066195314522  M4_M3_CDNS_4066195314522_13
timestamp 1698431365
transform 1 0 102 0 1 25906
box 0 0 1 1
use M4_M3_CDNS_4066195314522  M4_M3_CDNS_4066195314522_14
timestamp 1698431365
transform 1 0 102 0 1 24313
box 0 0 1 1
use M4_M3_CDNS_4066195314522  M4_M3_CDNS_4066195314522_15
timestamp 1698431365
transform 1 0 102 0 1 49894
box 0 0 1 1
use M4_M3_CDNS_4066195314523  M4_M3_CDNS_4066195314523_0
timestamp 1698431365
transform 1 0 101 0 1 69037
box 0 0 1 1
use M4_M3_CDNS_4066195314524  M4_M3_CDNS_4066195314524_0
timestamp 1698431365
transform 1 0 101 0 1 44298
box 0 0 1 1
use M4_M3_CDNS_4066195314524  M4_M3_CDNS_4066195314524_1
timestamp 1698431365
transform 1 0 101 0 1 37904
box 0 0 1 1
use M4_M3_CDNS_4066195314524  M4_M3_CDNS_4066195314524_2
timestamp 1698431365
transform 1 0 101 0 1 34703
box 0 0 1 1
use M4_M3_CDNS_4066195314524  M4_M3_CDNS_4066195314524_3
timestamp 1698431365
transform 1 0 101 0 1 31507
box 0 0 1 1
use M4_M3_CDNS_4066195314524  M4_M3_CDNS_4066195314524_4
timestamp 1698431365
transform 1 0 101 0 1 28313
box 0 0 1 1
use M4_M3_CDNS_4066195314524  M4_M3_CDNS_4066195314524_5
timestamp 1698431365
transform 1 0 101 0 1 21951
box 0 0 1 1
use M4_M3_CDNS_4066195314524  M4_M3_CDNS_4066195314524_6
timestamp 1698431365
transform 1 0 101 0 1 18701
box 0 0 1 1
use M4_M3_CDNS_4066195314524  M4_M3_CDNS_4066195314524_7
timestamp 1698431365
transform 1 0 101 0 1 15500
box 0 0 1 1
use M4_M3_CDNS_4066195314524  M4_M3_CDNS_4066195314524_8
timestamp 1698431365
transform 1 0 101 0 1 47512
box 0 0 1 1
<< labels >>
rlabel metal3 s 94 37959 94 37959 4 DVDD
port 1 nsew
rlabel metal3 s 94 34723 94 34723 4 DVDD
port 1 nsew
rlabel metal3 s 94 44368 94 44368 4 DVDD
port 1 nsew
rlabel metal3 s 94 41977 94 41977 4 DVDD
port 1 nsew
rlabel metal3 s 94 61058 94 61058 4 DVSS
port 2 nsew
rlabel metal3 s 94 66023 94 66023 4 DVSS
port 2 nsew
rlabel metal3 s 94 69049 94 69049 4 DVSS
port 2 nsew
rlabel metal3 s 94 31609 94 31609 4 DVDD
port 1 nsew
rlabel metal3 s 94 28394 94 28394 4 DVDD
port 1 nsew
rlabel metal3 s 94 24284 94 24284 4 DVDD
port 1 nsew
rlabel metal3 s 94 59623 94 59623 4 DVDD
port 1 nsew
rlabel metal3 s 94 56423 94 56423 4 DVDD
port 1 nsew
rlabel metal3 s 94 54658 94 54658 4 DVDD
port 1 nsew
rlabel metal3 s 94 53223 94 53223 4 DVDD
port 1 nsew
rlabel metal3 s 94 64258 94 64258 4 VSS
port 3 nsew
rlabel metal3 s 94 50023 94 50023 4 VSS
port 3 nsew
rlabel metal3 s 94 51458 94 51458 4 VDD
port 4 nsew
rlabel metal3 s 94 62823 94 62823 4 VDD
port 4 nsew
rlabel metal3 s 94 18921 94 18921 4 DVSS
port 2 nsew
rlabel metal3 s 94 15750 94 15750 4 DVSS
port 2 nsew
rlabel metal3 s 94 21907 94 21907 4 DVSS
port 2 nsew
rlabel metal3 s 94 26100 94 26100 4 DVSS
port 2 nsew
rlabel metal3 s 94 40342 94 40342 4 DVSS
port 2 nsew
rlabel metal3 s 94 47595 94 47595 4 DVSS
port 2 nsew
rlabel metal3 s 94 57858 94 57858 4 DVSS
port 2 nsew
rlabel metal3 s 94 67458 94 67458 4 DVDD
port 1 nsew
rlabel metal4 s 94 67458 94 67458 4 DVDD
port 1 nsew
rlabel metal4 s 94 50023 94 50023 4 VSS
port 3 nsew
rlabel metal4 s 94 34723 94 34723 4 DVDD
port 1 nsew
rlabel metal4 s 94 37959 94 37959 4 DVDD
port 1 nsew
rlabel metal4 s 94 41977 94 41977 4 DVDD
port 1 nsew
rlabel metal4 s 94 44368 94 44368 4 DVDD
port 1 nsew
rlabel metal4 s 94 53223 94 53223 4 DVDD
port 1 nsew
rlabel metal4 s 94 54658 94 54658 4 DVDD
port 1 nsew
rlabel metal4 s 94 56423 94 56423 4 DVDD
port 1 nsew
rlabel metal4 s 94 59623 94 59623 4 DVDD
port 1 nsew
rlabel metal4 s 94 64258 94 64258 4 VSS
port 3 nsew
rlabel metal4 s 94 62823 94 62823 4 VDD
port 4 nsew
rlabel metal4 s 94 51458 94 51458 4 VDD
port 4 nsew
rlabel metal4 s 94 69049 94 69049 4 DVSS
port 2 nsew
rlabel metal4 s 94 66023 94 66023 4 DVSS
port 2 nsew
rlabel metal4 s 94 61058 94 61058 4 DVSS
port 2 nsew
rlabel metal4 s 94 57858 94 57858 4 DVSS
port 2 nsew
rlabel metal4 s 94 47595 94 47595 4 DVSS
port 2 nsew
rlabel metal4 s 94 40342 94 40342 4 DVSS
port 2 nsew
rlabel metal4 s 94 26100 94 26100 4 DVSS
port 2 nsew
rlabel metal4 s 94 21907 94 21907 4 DVSS
port 2 nsew
rlabel metal4 s 94 15750 94 15750 4 DVSS
port 2 nsew
rlabel metal4 s 94 18921 94 18921 4 DVSS
port 2 nsew
rlabel metal4 s 94 24284 94 24284 4 DVDD
port 1 nsew
rlabel metal4 s 94 28394 94 28394 4 DVDD
port 1 nsew
rlabel metal4 s 94 31609 94 31609 4 DVDD
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 200 70000
string GDS_END 5040828
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 5035730
<< end >>
