magic
tech gf180mcuB
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -83 1292 1139 2586
<< mvnmos >>
rect 336 281 476 881
rect 580 281 720 881
<< mvpmos >>
rect 336 1633 476 2233
rect 580 1633 720 2233
<< mvndiff >>
rect 248 868 336 881
rect 248 822 261 868
rect 307 822 336 868
rect 248 763 336 822
rect 248 717 261 763
rect 307 717 336 763
rect 248 658 336 717
rect 248 612 261 658
rect 307 612 336 658
rect 248 552 336 612
rect 248 506 261 552
rect 307 506 336 552
rect 248 446 336 506
rect 248 400 261 446
rect 307 400 336 446
rect 248 340 336 400
rect 248 294 261 340
rect 307 294 336 340
rect 248 281 336 294
rect 476 868 580 881
rect 476 822 505 868
rect 551 822 580 868
rect 476 763 580 822
rect 476 717 505 763
rect 551 717 580 763
rect 476 658 580 717
rect 476 612 505 658
rect 551 612 580 658
rect 476 552 580 612
rect 476 506 505 552
rect 551 506 580 552
rect 476 446 580 506
rect 476 400 505 446
rect 551 400 580 446
rect 476 340 580 400
rect 476 294 505 340
rect 551 294 580 340
rect 476 281 580 294
rect 720 868 808 881
rect 720 822 749 868
rect 795 822 808 868
rect 720 763 808 822
rect 720 717 749 763
rect 795 717 808 763
rect 720 658 808 717
rect 720 612 749 658
rect 795 612 808 658
rect 720 552 808 612
rect 720 506 749 552
rect 795 506 808 552
rect 720 446 808 506
rect 720 400 749 446
rect 795 400 808 446
rect 720 340 808 400
rect 720 294 749 340
rect 795 294 808 340
rect 720 281 808 294
<< mvpdiff >>
rect 248 2220 336 2233
rect 248 2174 261 2220
rect 307 2174 336 2220
rect 248 2115 336 2174
rect 248 2069 261 2115
rect 307 2069 336 2115
rect 248 2010 336 2069
rect 248 1964 261 2010
rect 307 1964 336 2010
rect 248 1904 336 1964
rect 248 1858 261 1904
rect 307 1858 336 1904
rect 248 1798 336 1858
rect 248 1752 261 1798
rect 307 1752 336 1798
rect 248 1692 336 1752
rect 248 1646 261 1692
rect 307 1646 336 1692
rect 248 1633 336 1646
rect 476 2220 580 2233
rect 476 2174 505 2220
rect 551 2174 580 2220
rect 476 2115 580 2174
rect 476 2069 505 2115
rect 551 2069 580 2115
rect 476 2010 580 2069
rect 476 1964 505 2010
rect 551 1964 580 2010
rect 476 1904 580 1964
rect 476 1858 505 1904
rect 551 1858 580 1904
rect 476 1798 580 1858
rect 476 1752 505 1798
rect 551 1752 580 1798
rect 476 1692 580 1752
rect 476 1646 505 1692
rect 551 1646 580 1692
rect 476 1633 580 1646
rect 720 2220 808 2233
rect 720 2174 749 2220
rect 795 2174 808 2220
rect 720 2115 808 2174
rect 720 2069 749 2115
rect 795 2069 808 2115
rect 720 2010 808 2069
rect 720 1964 749 2010
rect 795 1964 808 2010
rect 720 1904 808 1964
rect 720 1858 749 1904
rect 795 1858 808 1904
rect 720 1798 808 1858
rect 720 1752 749 1798
rect 795 1752 808 1798
rect 720 1692 808 1752
rect 720 1646 749 1692
rect 795 1646 808 1692
rect 720 1633 808 1646
<< mvndiffc >>
rect 261 822 307 868
rect 261 717 307 763
rect 261 612 307 658
rect 261 506 307 552
rect 261 400 307 446
rect 261 294 307 340
rect 505 822 551 868
rect 505 717 551 763
rect 505 612 551 658
rect 505 506 551 552
rect 505 400 551 446
rect 505 294 551 340
rect 749 822 795 868
rect 749 717 795 763
rect 749 612 795 658
rect 749 506 795 552
rect 749 400 795 446
rect 749 294 795 340
<< mvpdiffc >>
rect 261 2174 307 2220
rect 261 2069 307 2115
rect 261 1964 307 2010
rect 261 1858 307 1904
rect 261 1752 307 1798
rect 261 1646 307 1692
rect 505 2174 551 2220
rect 505 2069 551 2115
rect 505 1964 551 2010
rect 505 1858 551 1904
rect 505 1752 551 1798
rect 505 1646 551 1692
rect 749 2174 795 2220
rect 749 2069 795 2115
rect 749 1964 795 2010
rect 749 1858 795 1904
rect 749 1752 795 1798
rect 749 1646 795 1692
<< psubdiff >>
rect 0 1019 90 1041
rect 0 33 22 1019
rect 68 101 90 1019
rect 966 1019 1056 1041
rect 966 101 988 1019
rect 68 79 988 101
rect 68 33 176 79
rect 880 33 988 79
rect 1034 33 1056 1019
rect 0 11 1056 33
<< nsubdiff >>
rect 0 2481 1056 2503
rect 0 1495 22 2481
rect 68 2435 176 2481
rect 880 2435 988 2481
rect 68 2413 988 2435
rect 68 1495 90 2413
rect 0 1473 90 1495
rect 966 1495 988 2413
rect 1034 1495 1056 2481
rect 966 1473 1056 1495
<< psubdiffcont >>
rect 22 33 68 1019
rect 176 33 880 79
rect 988 33 1034 1019
<< nsubdiffcont >>
rect 22 1495 68 2481
rect 176 2435 880 2481
rect 988 1495 1034 2481
<< polysilicon >>
rect 336 2233 476 2277
rect 580 2233 720 2277
rect 336 1333 476 1633
rect 336 1193 383 1333
rect 429 1193 476 1333
rect 336 881 476 1193
rect 580 1333 720 1633
rect 580 1193 627 1333
rect 673 1193 720 1333
rect 580 881 720 1193
rect 336 237 476 281
rect 580 237 720 281
<< polycontact >>
rect 383 1193 429 1333
rect 627 1193 673 1333
<< metal1 >>
rect 11 2481 1045 2492
rect 11 1495 22 2481
rect 68 2435 176 2481
rect 880 2435 988 2481
rect 68 2424 988 2435
rect 68 1495 79 2424
rect 246 2220 322 2424
rect 246 2174 261 2220
rect 307 2174 322 2220
rect 246 2115 322 2174
rect 246 2069 261 2115
rect 307 2069 322 2115
rect 246 2010 322 2069
rect 246 1964 261 2010
rect 307 1964 322 2010
rect 246 1904 322 1964
rect 246 1858 261 1904
rect 307 1858 322 1904
rect 246 1798 322 1858
rect 246 1752 261 1798
rect 307 1752 322 1798
rect 246 1692 322 1752
rect 246 1646 261 1692
rect 307 1646 322 1692
rect 246 1633 322 1646
rect 490 2220 566 2233
rect 490 2174 505 2220
rect 551 2174 566 2220
rect 490 2115 566 2174
rect 490 2069 505 2115
rect 551 2069 566 2115
rect 490 2010 566 2069
rect 490 1964 505 2010
rect 551 1964 566 2010
rect 490 1904 566 1964
rect 490 1858 505 1904
rect 551 1858 566 1904
rect 490 1798 566 1858
rect 490 1752 505 1798
rect 551 1752 566 1798
rect 490 1692 566 1752
rect 490 1646 505 1692
rect 551 1646 566 1692
rect 11 1484 79 1495
rect 372 1333 440 1344
rect 372 1193 383 1333
rect 429 1193 440 1333
rect 372 1182 440 1193
rect 490 1088 566 1646
rect 734 2220 810 2424
rect 734 2174 749 2220
rect 795 2174 810 2220
rect 734 2115 810 2174
rect 734 2069 749 2115
rect 795 2069 810 2115
rect 734 2010 810 2069
rect 734 1964 749 2010
rect 795 1964 810 2010
rect 734 1904 810 1964
rect 734 1858 749 1904
rect 795 1858 810 1904
rect 734 1798 810 1858
rect 734 1752 749 1798
rect 795 1752 810 1798
rect 734 1692 810 1752
rect 734 1646 749 1692
rect 795 1646 810 1692
rect 734 1633 810 1646
rect 977 1495 988 2424
rect 1034 1495 1045 2481
rect 977 1484 1045 1495
rect 616 1333 684 1344
rect 616 1193 627 1333
rect 673 1193 684 1333
rect 616 1182 684 1193
rect 11 1019 79 1030
rect 11 33 22 1019
rect 68 90 79 1019
rect 490 1012 810 1088
rect 246 868 322 881
rect 246 822 261 868
rect 307 822 322 868
rect 246 763 322 822
rect 246 717 261 763
rect 307 717 322 763
rect 246 658 322 717
rect 246 612 261 658
rect 307 612 322 658
rect 246 552 322 612
rect 246 506 261 552
rect 307 506 322 552
rect 246 446 322 506
rect 246 400 261 446
rect 307 400 322 446
rect 246 340 322 400
rect 246 294 261 340
rect 307 294 322 340
rect 246 90 322 294
rect 505 868 551 881
rect 505 763 551 822
rect 505 658 551 717
rect 505 552 551 612
rect 505 446 551 506
rect 505 340 551 400
rect 505 281 551 294
rect 734 868 810 1012
rect 734 822 749 868
rect 795 822 810 868
rect 734 763 810 822
rect 734 717 749 763
rect 795 717 810 763
rect 734 658 810 717
rect 734 612 749 658
rect 795 612 810 658
rect 734 552 810 612
rect 734 506 749 552
rect 795 506 810 552
rect 734 446 810 506
rect 734 400 749 446
rect 795 400 810 446
rect 734 340 810 400
rect 734 294 749 340
rect 795 294 810 340
rect 734 281 810 294
rect 977 1019 1045 1030
rect 977 90 988 1019
rect 68 79 988 90
rect 68 33 176 79
rect 880 33 988 79
rect 1034 33 1045 1019
rect 11 22 1045 33
use M1_NWELL_CDNS_40661954729412  M1_NWELL_CDNS_40661954729412_0
timestamp 1698431365
transform 1 0 1011 0 1 1988
box 0 0 1 1
use M1_NWELL_CDNS_40661954729412  M1_NWELL_CDNS_40661954729412_1
timestamp 1698431365
transform 1 0 45 0 1 1988
box 0 0 1 1
use M1_NWELL_CDNS_40661954729426  M1_NWELL_CDNS_40661954729426_0
timestamp 1698431365
transform 1 0 528 0 1 2458
box 0 0 1 1
use M1_POLY2_CDNS_40661954729415  M1_POLY2_CDNS_40661954729415_0
timestamp 1698431365
transform 1 0 650 0 1 1263
box 0 0 1 1
use M1_POLY2_CDNS_40661954729415  M1_POLY2_CDNS_40661954729415_1
timestamp 1698431365
transform 1 0 406 0 1 1263
box 0 0 1 1
use M1_PSUB_CDNS_40661954729413  M1_PSUB_CDNS_40661954729413_0
timestamp 1698431365
transform 1 0 1011 0 -1 526
box 0 0 1 1
use M1_PSUB_CDNS_40661954729413  M1_PSUB_CDNS_40661954729413_1
timestamp 1698431365
transform 1 0 45 0 -1 526
box 0 0 1 1
use M1_PSUB_CDNS_40661954729427  M1_PSUB_CDNS_40661954729427_0
timestamp 1698431365
transform 1 0 528 0 -1 56
box 0 0 1 1
use nmos_6p0_CDNS_4066195472927  nmos_6p0_CDNS_4066195472927_0
timestamp 1698431365
transform 1 0 336 0 1 281
box 0 0 1 1
use nmos_6p0_CDNS_4066195472927  nmos_6p0_CDNS_4066195472927_1
timestamp 1698431365
transform 1 0 580 0 1 281
box 0 0 1 1
use pmos_6p0_CDNS_4066195472911  pmos_6p0_CDNS_4066195472911_0
timestamp 1698431365
transform -1 0 720 0 1 1633
box 0 0 1 1
use pmos_6p0_CDNS_4066195472911  pmos_6p0_CDNS_4066195472911_1
timestamp 1698431365
transform 1 0 336 0 1 1633
box 0 0 1 1
<< labels >>
rlabel metal1 s 75 2463 75 2463 4 VDD
port 1 nsew
rlabel metal1 s 244 56 244 56 4 VSS
port 2 nsew
rlabel metal1 s 407 1268 407 1268 4 A
port 3 nsew
rlabel metal1 s 652 1268 652 1268 4 B
port 4 nsew
rlabel metal1 s 528 1268 528 1268 4 Z
port 5 nsew
<< properties >>
string GDS_END 1419138
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 1417280
string path 19.300 40.825 19.300 61.900 
<< end >>
