magic
tech gf180mcuA
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 459 2550 1094
rect -86 453 86 459
rect 1863 453 2550 459
<< pwell >>
rect 86 453 1863 459
rect -86 -86 2550 453
<< mvnmos >>
rect 386 267 506 339
rect 124 123 244 195
rect 386 123 506 195
rect 818 212 938 284
rect 1186 212 1306 284
rect 818 68 938 140
rect 1186 68 1306 140
rect 1618 213 1738 285
rect 1618 69 1738 141
rect 1978 69 2098 333
rect 2202 69 2322 333
<< mvpmos >>
rect 124 781 224 853
rect 386 781 486 853
rect 386 637 486 709
rect 818 781 918 853
rect 1186 781 1286 853
rect 818 637 918 709
rect 1186 637 1286 709
rect 1618 781 1718 853
rect 1618 637 1718 709
rect 1978 574 2078 940
rect 2212 574 2312 940
<< mvndiff >>
rect 298 326 386 339
rect 298 280 311 326
rect 357 280 386 326
rect 298 267 386 280
rect 506 267 626 339
rect 566 195 626 267
rect 36 182 124 195
rect 36 136 49 182
rect 95 136 124 182
rect 36 123 124 136
rect 244 182 386 195
rect 244 136 273 182
rect 319 136 386 182
rect 244 123 386 136
rect 506 123 626 195
rect 698 212 818 284
rect 938 271 1026 284
rect 938 225 967 271
rect 1013 225 1026 271
rect 938 212 1026 225
rect 1098 271 1186 284
rect 1098 225 1111 271
rect 1157 225 1186 271
rect 1098 212 1186 225
rect 1306 212 1426 284
rect 698 140 758 212
rect 1366 140 1426 212
rect 698 68 818 140
rect 938 127 1186 140
rect 938 81 967 127
rect 1013 81 1186 127
rect 938 68 1186 81
rect 1306 68 1426 140
rect 1498 213 1618 285
rect 1738 272 1826 285
rect 1738 226 1767 272
rect 1813 226 1826 272
rect 1738 213 1826 226
rect 1498 141 1558 213
rect 1898 141 1978 333
rect 1498 69 1618 141
rect 1738 128 1978 141
rect 1738 82 1767 128
rect 1813 82 1978 128
rect 1738 69 1978 82
rect 2098 287 2202 333
rect 2098 147 2127 287
rect 2173 147 2202 287
rect 2098 69 2202 147
rect 2322 276 2410 333
rect 2322 136 2351 276
rect 2397 136 2410 276
rect 2322 69 2410 136
<< mvpdiff >>
rect 1898 853 1978 940
rect 36 840 124 853
rect 36 794 49 840
rect 95 794 124 840
rect 36 781 124 794
rect 224 840 386 853
rect 224 794 253 840
rect 299 794 386 840
rect 224 781 386 794
rect 486 781 606 853
rect 546 709 606 781
rect 298 696 386 709
rect 298 650 311 696
rect 357 650 386 696
rect 298 637 386 650
rect 486 637 606 709
rect 698 781 818 853
rect 918 840 1186 853
rect 918 794 947 840
rect 993 794 1186 840
rect 918 781 1186 794
rect 1286 781 1406 853
rect 698 709 758 781
rect 1346 709 1406 781
rect 698 637 818 709
rect 918 696 1006 709
rect 918 650 947 696
rect 993 650 1006 696
rect 918 637 1006 650
rect 1098 696 1186 709
rect 1098 650 1111 696
rect 1157 650 1186 696
rect 1098 637 1186 650
rect 1286 637 1406 709
rect 1498 781 1618 853
rect 1718 840 1978 853
rect 1718 794 1747 840
rect 1793 794 1978 840
rect 1718 781 1978 794
rect 1498 709 1558 781
rect 1498 637 1618 709
rect 1718 696 1806 709
rect 1718 650 1747 696
rect 1793 650 1806 696
rect 1718 637 1806 650
rect 1898 574 1978 781
rect 2078 861 2212 940
rect 2078 721 2127 861
rect 2173 721 2212 861
rect 2078 574 2212 721
rect 2312 927 2400 940
rect 2312 787 2341 927
rect 2387 787 2400 927
rect 2312 574 2400 787
<< mvndiffc >>
rect 311 280 357 326
rect 49 136 95 182
rect 273 136 319 182
rect 967 225 1013 271
rect 1111 225 1157 271
rect 967 81 1013 127
rect 1767 226 1813 272
rect 1767 82 1813 128
rect 2127 147 2173 287
rect 2351 136 2397 276
<< mvpdiffc >>
rect 49 794 95 840
rect 253 794 299 840
rect 311 650 357 696
rect 947 794 993 840
rect 947 650 993 696
rect 1111 650 1157 696
rect 1747 794 1793 840
rect 1747 650 1793 696
rect 2127 721 2173 861
rect 2341 787 2387 927
<< polysilicon >>
rect 1978 940 2078 984
rect 2212 940 2312 984
rect 124 853 224 897
rect 386 853 486 897
rect 818 853 918 897
rect 1186 853 1286 897
rect 1618 853 1718 897
rect 124 512 224 781
rect 386 709 486 781
rect 818 709 918 781
rect 1186 709 1286 781
rect 1618 709 1718 781
rect 124 372 141 512
rect 187 372 224 512
rect 124 239 224 372
rect 386 512 486 637
rect 386 372 399 512
rect 445 383 486 512
rect 818 512 918 637
rect 445 372 506 383
rect 386 339 506 372
rect 818 372 831 512
rect 877 372 918 512
rect 818 328 918 372
rect 1186 512 1286 637
rect 1186 372 1199 512
rect 1245 372 1286 512
rect 1186 328 1286 372
rect 1618 512 1718 637
rect 1618 372 1631 512
rect 1677 372 1718 512
rect 1978 478 2078 574
rect 1818 465 2078 478
rect 2212 465 2312 574
rect 1818 419 1831 465
rect 2065 419 2312 465
rect 1818 406 2312 419
rect 1618 329 1718 372
rect 1978 393 2312 406
rect 1978 333 2098 393
rect 2202 377 2312 393
rect 2202 333 2322 377
rect 818 284 938 328
rect 1186 284 1306 328
rect 1618 285 1738 329
rect 124 195 244 239
rect 386 195 506 267
rect 818 140 938 212
rect 1186 140 1306 212
rect 124 79 244 123
rect 386 79 506 123
rect 1618 141 1738 213
rect 818 24 938 68
rect 1186 24 1306 68
rect 1618 25 1738 69
rect 1978 25 2098 69
rect 2202 25 2322 69
<< polycontact >>
rect 141 372 187 512
rect 399 372 445 512
rect 831 372 877 512
rect 1199 372 1245 512
rect 1631 372 1677 512
rect 1831 419 2065 465
<< metal1 >>
rect 0 927 2464 1098
rect 0 918 2341 927
rect 38 840 95 851
rect 38 794 49 840
rect 38 604 95 794
rect 253 840 299 918
rect 253 783 299 794
rect 947 840 993 918
rect 947 783 993 794
rect 1747 840 1793 918
rect 1747 783 1793 794
rect 2127 861 2173 872
rect 2387 918 2464 927
rect 2341 776 2387 787
rect 947 696 993 707
rect 300 650 311 696
rect 357 650 548 696
rect 38 558 456 604
rect 38 182 84 558
rect 388 512 456 558
rect 130 372 141 512
rect 187 372 198 512
rect 388 372 399 512
rect 445 372 456 512
rect 130 354 198 372
rect 502 326 548 650
rect 831 512 877 523
rect 831 326 877 372
rect 300 280 311 326
rect 357 280 877 326
rect 947 418 993 650
rect 1111 696 1157 707
rect 1111 604 1157 650
rect 1747 696 1793 707
rect 1111 558 1348 604
rect 1188 418 1199 512
rect 947 372 1199 418
rect 1245 372 1256 512
rect 947 271 1013 372
rect 1302 326 1348 558
rect 1631 512 1677 523
rect 1631 326 1677 372
rect 947 225 967 271
rect 947 214 1013 225
rect 1111 280 1677 326
rect 1747 465 1793 650
rect 1747 419 1831 465
rect 2065 419 2076 465
rect 1111 271 1157 280
rect 1111 214 1157 225
rect 1747 272 1813 419
rect 2127 318 2173 721
rect 1747 226 1767 272
rect 2046 287 2173 318
rect 2046 242 2127 287
rect 1747 215 1813 226
rect 273 182 319 193
rect 38 136 49 182
rect 95 136 106 182
rect 273 90 319 136
rect 967 127 1013 138
rect 0 81 967 90
rect 1767 128 1813 139
rect 2127 136 2173 147
rect 2351 276 2397 287
rect 1013 82 1767 90
rect 2351 90 2397 136
rect 1813 82 2464 90
rect 1013 81 2464 82
rect 0 -90 2464 81
<< labels >>
flabel metal1 s 130 354 198 512 0 FreeSans 200 0 0 0 I
port 1 nsew default input
flabel metal1 s 0 918 2464 1098 0 FreeSans 200 0 0 0 VDD
port 3 nsew power bidirectional abutment
flabel metal1 s 2351 193 2397 287 0 FreeSans 200 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel metal1 s 2127 318 2173 872 0 FreeSans 200 0 0 0 Z
port 2 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 4 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 2046 242 2173 318 1 Z
port 2 nsew default output
rlabel metal1 s 2127 136 2173 242 1 Z
port 2 nsew default output
rlabel metal1 s 2341 783 2387 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1747 783 1793 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 947 783 993 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 253 783 299 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2341 776 2387 783 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2351 139 2397 193 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 273 139 319 193 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2351 138 2397 139 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1767 138 1813 139 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 273 138 319 139 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2351 90 2397 138 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1767 90 1813 138 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 967 90 1013 138 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 138 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 2464 90 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2464 1008
string GDS_END 733666
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 727644
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
