magic
tech gf180mcuA
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 377 6134 870
rect -86 352 688 377
rect 1688 352 6134 377
<< pwell >>
rect 688 352 1688 377
rect -86 -86 6134 352
<< mvnmos >>
rect 134 68 254 232
rect 358 68 478 232
rect 582 68 702 232
rect 1050 68 1170 232
rect 1362 68 1482 232
rect 1674 68 1794 232
rect 1986 68 2106 232
rect 2210 68 2330 232
rect 2434 68 2554 232
rect 2658 68 2778 232
rect 2882 68 3002 232
rect 3106 68 3226 232
rect 3330 68 3450 232
rect 3554 68 3674 232
rect 3778 68 3898 232
rect 4002 68 4122 232
rect 4226 68 4346 232
rect 4450 68 4570 232
rect 4674 68 4794 232
rect 4898 68 5018 232
rect 5122 68 5242 232
rect 5346 68 5466 232
rect 5570 68 5690 232
rect 5794 68 5914 232
<< mvpmos >>
rect 197 497 297 716
rect 401 497 501 716
rect 605 497 705 716
rect 1118 497 1218 716
rect 1410 497 1510 716
rect 1614 497 1714 716
rect 2082 480 2182 716
rect 2286 480 2386 716
rect 2490 480 2590 716
rect 2694 480 2794 716
rect 2898 480 2998 716
rect 3116 480 3216 716
rect 3340 480 3440 716
rect 3564 480 3664 716
rect 3788 480 3888 716
rect 4012 480 4112 716
rect 4236 480 4336 716
rect 4460 480 4560 716
rect 4664 480 4764 716
rect 4868 480 4968 716
rect 5072 480 5172 716
rect 5276 480 5376 716
rect 5480 480 5580 716
rect 5684 480 5784 716
<< mvndiff >>
rect 762 244 834 257
rect 762 232 775 244
rect 46 200 134 232
rect 46 154 59 200
rect 105 154 134 200
rect 46 68 134 154
rect 254 139 358 232
rect 254 93 283 139
rect 329 93 358 139
rect 254 68 358 93
rect 478 166 582 232
rect 478 120 507 166
rect 553 120 582 166
rect 478 68 582 120
rect 702 198 775 232
rect 821 198 834 244
rect 702 68 834 198
rect 918 244 990 257
rect 918 198 931 244
rect 977 232 990 244
rect 1542 244 1614 257
rect 1542 232 1555 244
rect 977 198 1050 232
rect 918 68 1050 198
rect 1170 95 1362 232
rect 1170 68 1243 95
rect 1230 49 1243 68
rect 1289 68 1362 95
rect 1482 198 1555 232
rect 1601 232 1614 244
rect 1601 198 1674 232
rect 1482 68 1674 198
rect 1794 95 1986 232
rect 1794 68 1867 95
rect 1289 49 1302 68
rect 1230 36 1302 49
rect 1854 49 1867 68
rect 1913 68 1986 95
rect 2106 187 2210 232
rect 2106 141 2135 187
rect 2181 141 2210 187
rect 2106 68 2210 141
rect 2330 175 2434 232
rect 2330 129 2359 175
rect 2405 129 2434 175
rect 2330 68 2434 129
rect 2554 175 2658 232
rect 2554 129 2583 175
rect 2629 129 2658 175
rect 2554 68 2658 129
rect 2778 175 2882 232
rect 2778 129 2807 175
rect 2853 129 2882 175
rect 2778 68 2882 129
rect 3002 175 3106 232
rect 3002 129 3031 175
rect 3077 129 3106 175
rect 3002 68 3106 129
rect 3226 175 3330 232
rect 3226 129 3255 175
rect 3301 129 3330 175
rect 3226 68 3330 129
rect 3450 219 3554 232
rect 3450 173 3479 219
rect 3525 173 3554 219
rect 3450 68 3554 173
rect 3674 127 3778 232
rect 3674 81 3703 127
rect 3749 81 3778 127
rect 3674 68 3778 81
rect 3898 219 4002 232
rect 3898 173 3927 219
rect 3973 173 4002 219
rect 3898 68 4002 173
rect 4122 127 4226 232
rect 4122 81 4151 127
rect 4197 81 4226 127
rect 4122 68 4226 81
rect 4346 219 4450 232
rect 4346 173 4375 219
rect 4421 173 4450 219
rect 4346 68 4450 173
rect 4570 127 4674 232
rect 4570 81 4599 127
rect 4645 81 4674 127
rect 4570 68 4674 81
rect 4794 219 4898 232
rect 4794 173 4823 219
rect 4869 173 4898 219
rect 4794 68 4898 173
rect 5018 127 5122 232
rect 5018 81 5047 127
rect 5093 81 5122 127
rect 5018 68 5122 81
rect 5242 219 5346 232
rect 5242 173 5271 219
rect 5317 173 5346 219
rect 5242 68 5346 173
rect 5466 127 5570 232
rect 5466 81 5495 127
rect 5541 81 5570 127
rect 5466 68 5570 81
rect 5690 219 5794 232
rect 5690 173 5719 219
rect 5765 173 5794 219
rect 5690 68 5794 173
rect 5914 172 6002 232
rect 5914 126 5943 172
rect 5989 126 6002 172
rect 5914 68 6002 126
rect 1913 49 1926 68
rect 1854 36 1926 49
<< mvpdiff >>
rect 1278 735 1350 748
rect 1278 716 1291 735
rect 109 665 197 716
rect 109 525 122 665
rect 168 525 197 665
rect 109 497 197 525
rect 297 683 401 716
rect 297 637 326 683
rect 372 637 401 683
rect 297 497 401 637
rect 501 671 605 716
rect 501 625 530 671
rect 576 625 605 671
rect 501 497 605 625
rect 705 556 793 716
rect 705 510 734 556
rect 780 510 793 556
rect 705 497 793 510
rect 1030 556 1118 716
rect 1030 510 1043 556
rect 1089 510 1118 556
rect 1030 497 1118 510
rect 1218 689 1291 716
rect 1337 716 1350 735
rect 1337 689 1410 716
rect 1218 497 1410 689
rect 1510 556 1614 716
rect 1510 510 1539 556
rect 1585 510 1614 556
rect 1510 497 1614 510
rect 1714 677 2082 716
rect 1714 631 1963 677
rect 2009 631 2082 677
rect 1714 497 2082 631
rect 1874 480 2082 497
rect 2182 665 2286 716
rect 2182 525 2211 665
rect 2257 525 2286 665
rect 2182 480 2286 525
rect 2386 665 2490 716
rect 2386 525 2415 665
rect 2461 525 2490 665
rect 2386 480 2490 525
rect 2590 665 2694 716
rect 2590 525 2619 665
rect 2665 525 2694 665
rect 2590 480 2694 525
rect 2794 665 2898 716
rect 2794 525 2823 665
rect 2869 525 2898 665
rect 2794 480 2898 525
rect 2998 665 3116 716
rect 2998 525 3027 665
rect 3073 525 3116 665
rect 2998 480 3116 525
rect 3216 665 3340 716
rect 3216 525 3245 665
rect 3291 525 3340 665
rect 3216 480 3340 525
rect 3440 665 3564 716
rect 3440 525 3489 665
rect 3535 525 3564 665
rect 3440 480 3564 525
rect 3664 703 3788 716
rect 3664 657 3693 703
rect 3739 657 3788 703
rect 3664 480 3788 657
rect 3888 665 4012 716
rect 3888 525 3917 665
rect 3963 525 4012 665
rect 3888 480 4012 525
rect 4112 703 4236 716
rect 4112 657 4141 703
rect 4187 657 4236 703
rect 4112 480 4236 657
rect 4336 665 4460 716
rect 4336 525 4365 665
rect 4411 525 4460 665
rect 4336 480 4460 525
rect 4560 703 4664 716
rect 4560 657 4589 703
rect 4635 657 4664 703
rect 4560 480 4664 657
rect 4764 665 4868 716
rect 4764 525 4793 665
rect 4839 525 4868 665
rect 4764 480 4868 525
rect 4968 703 5072 716
rect 4968 657 4997 703
rect 5043 657 5072 703
rect 4968 480 5072 657
rect 5172 665 5276 716
rect 5172 525 5201 665
rect 5247 525 5276 665
rect 5172 480 5276 525
rect 5376 703 5480 716
rect 5376 657 5405 703
rect 5451 657 5480 703
rect 5376 480 5480 657
rect 5580 665 5684 716
rect 5580 525 5609 665
rect 5655 525 5684 665
rect 5580 480 5684 525
rect 5784 665 5872 716
rect 5784 525 5813 665
rect 5859 525 5872 665
rect 5784 480 5872 525
<< mvndiffc >>
rect 59 154 105 200
rect 283 93 329 139
rect 507 120 553 166
rect 775 198 821 244
rect 931 198 977 244
rect 1243 49 1289 95
rect 1555 198 1601 244
rect 1867 49 1913 95
rect 2135 141 2181 187
rect 2359 129 2405 175
rect 2583 129 2629 175
rect 2807 129 2853 175
rect 3031 129 3077 175
rect 3255 129 3301 175
rect 3479 173 3525 219
rect 3703 81 3749 127
rect 3927 173 3973 219
rect 4151 81 4197 127
rect 4375 173 4421 219
rect 4599 81 4645 127
rect 4823 173 4869 219
rect 5047 81 5093 127
rect 5271 173 5317 219
rect 5495 81 5541 127
rect 5719 173 5765 219
rect 5943 126 5989 172
<< mvpdiffc >>
rect 122 525 168 665
rect 326 637 372 683
rect 530 625 576 671
rect 734 510 780 556
rect 1043 510 1089 556
rect 1291 689 1337 735
rect 1539 510 1585 556
rect 1963 631 2009 677
rect 2211 525 2257 665
rect 2415 525 2461 665
rect 2619 525 2665 665
rect 2823 525 2869 665
rect 3027 525 3073 665
rect 3245 525 3291 665
rect 3489 525 3535 665
rect 3693 657 3739 703
rect 3917 525 3963 665
rect 4141 657 4187 703
rect 4365 525 4411 665
rect 4589 657 4635 703
rect 4793 525 4839 665
rect 4997 657 5043 703
rect 5201 525 5247 665
rect 5405 657 5451 703
rect 5609 525 5655 665
rect 5813 525 5859 665
<< polysilicon >>
rect 197 716 297 760
rect 401 716 501 760
rect 605 716 705 760
rect 1118 716 1218 760
rect 1410 716 1510 760
rect 1614 716 1714 760
rect 2082 716 2182 760
rect 2286 716 2386 760
rect 2490 716 2590 760
rect 2694 716 2794 760
rect 2898 716 2998 760
rect 3116 716 3216 760
rect 3340 716 3440 760
rect 3564 716 3664 760
rect 3788 716 3888 760
rect 4012 716 4112 760
rect 4236 716 4336 760
rect 4460 716 4560 760
rect 4664 716 4764 760
rect 4868 716 4968 760
rect 5072 716 5172 760
rect 5276 716 5376 760
rect 5480 716 5580 760
rect 5684 716 5784 760
rect 197 437 297 497
rect 134 424 297 437
rect 134 378 158 424
rect 204 412 297 424
rect 401 412 501 497
rect 605 464 705 497
rect 605 418 618 464
rect 664 418 705 464
rect 1118 437 1218 497
rect 1410 437 1510 497
rect 1614 437 1714 497
rect 204 378 557 412
rect 605 405 705 418
rect 1050 424 1714 437
rect 134 372 557 378
rect 134 232 254 372
rect 517 345 557 372
rect 1050 378 1066 424
rect 1676 378 1714 424
rect 2082 391 2182 480
rect 2286 391 2386 480
rect 2490 391 2590 480
rect 2694 391 2794 480
rect 2898 391 2998 480
rect 3116 391 3216 480
rect 1050 365 1714 378
rect 358 311 457 324
rect 358 265 387 311
rect 433 276 457 311
rect 517 305 622 345
rect 582 288 622 305
rect 433 265 478 276
rect 358 232 478 265
rect 582 232 702 288
rect 1050 232 1170 365
rect 1362 232 1482 365
rect 1674 363 1714 365
rect 1986 378 3216 391
rect 3340 439 3440 480
rect 3340 393 3366 439
rect 3412 420 3440 439
rect 3564 439 3664 480
rect 3564 420 3591 439
rect 3412 393 3591 420
rect 3637 420 3664 439
rect 3788 439 3888 480
rect 3788 420 3817 439
rect 3637 393 3817 420
rect 3863 420 3888 439
rect 4012 439 4112 480
rect 4012 420 4039 439
rect 3863 393 4039 420
rect 4085 420 4112 439
rect 4236 439 4336 480
rect 4236 420 4251 439
rect 4085 393 4251 420
rect 4297 420 4336 439
rect 4460 439 4560 480
rect 4460 420 4473 439
rect 4297 393 4473 420
rect 4519 420 4560 439
rect 4664 420 4764 480
rect 4868 439 4968 480
rect 4868 420 4892 439
rect 4519 393 4892 420
rect 4938 420 4968 439
rect 5072 439 5172 480
rect 5072 420 5099 439
rect 4938 393 5099 420
rect 5145 420 5172 439
rect 5276 439 5376 480
rect 5276 420 5305 439
rect 5145 393 5305 420
rect 5351 420 5376 439
rect 5480 439 5580 480
rect 5480 420 5508 439
rect 5351 393 5508 420
rect 5554 420 5580 439
rect 5684 439 5784 480
rect 5684 420 5711 439
rect 5554 393 5711 420
rect 5757 393 5784 439
rect 3340 380 5784 393
rect 134 24 254 68
rect 358 24 478 68
rect 582 24 702 68
rect 1050 24 1170 68
rect 1674 232 1794 363
rect 1986 332 2004 378
rect 3178 332 3216 378
rect 1986 319 3216 332
rect 1986 232 2106 319
rect 2210 232 2330 319
rect 2434 232 2554 319
rect 2658 232 2778 319
rect 2882 232 3002 319
rect 3106 287 3216 319
rect 3330 319 5914 332
rect 3106 232 3226 287
rect 3330 273 3362 319
rect 3408 292 3591 319
rect 3408 273 3450 292
rect 3330 232 3450 273
rect 3554 273 3591 292
rect 3637 292 3819 319
rect 3637 273 3674 292
rect 3554 232 3674 273
rect 3778 273 3819 292
rect 3865 292 4038 319
rect 3865 273 3898 292
rect 3778 232 3898 273
rect 4002 273 4038 292
rect 4084 292 5383 319
rect 4084 273 4122 292
rect 4002 232 4122 273
rect 4226 232 4346 292
rect 4450 232 4570 292
rect 4674 232 4794 292
rect 4898 232 5018 292
rect 5122 232 5242 292
rect 5346 273 5383 292
rect 5429 292 5608 319
rect 5429 273 5466 292
rect 5346 232 5466 273
rect 5570 273 5608 292
rect 5654 292 5831 319
rect 5654 273 5690 292
rect 5570 232 5690 273
rect 5794 273 5831 292
rect 5877 273 5914 319
rect 5794 232 5914 273
rect 1362 24 1482 68
rect 1674 24 1794 68
rect 1986 24 2106 68
rect 2210 24 2330 68
rect 2434 24 2554 68
rect 2658 24 2778 68
rect 2882 24 3002 68
rect 3106 24 3226 68
rect 3330 24 3450 68
rect 3554 24 3674 68
rect 3778 24 3898 68
rect 4002 24 4122 68
rect 4226 24 4346 68
rect 4450 24 4570 68
rect 4674 24 4794 68
rect 4898 24 5018 68
rect 5122 24 5242 68
rect 5346 24 5466 68
rect 5570 24 5690 68
rect 5794 24 5914 68
<< polycontact >>
rect 158 378 204 424
rect 618 418 664 464
rect 1066 378 1676 424
rect 387 265 433 311
rect 3366 393 3412 439
rect 3591 393 3637 439
rect 3817 393 3863 439
rect 4039 393 4085 439
rect 4251 393 4297 439
rect 4473 393 4519 439
rect 4892 393 4938 439
rect 5099 393 5145 439
rect 5305 393 5351 439
rect 5508 393 5554 439
rect 5711 393 5757 439
rect 2004 332 3178 378
rect 3362 273 3408 319
rect 3591 273 3637 319
rect 3819 273 3865 319
rect 4038 273 4084 319
rect 5383 273 5429 319
rect 5608 273 5654 319
rect 5831 273 5877 319
<< metal1 >>
rect 0 735 6048 844
rect 0 724 1291 735
rect 326 683 372 724
rect 1280 689 1291 724
rect 1337 724 6048 735
rect 1337 689 1348 724
rect 122 665 168 676
rect 1963 677 2009 724
rect 326 626 372 637
rect 519 625 530 671
rect 576 643 1234 671
rect 1394 643 1898 671
rect 576 625 1898 643
rect 826 602 1898 625
rect 1963 620 2009 631
rect 2211 665 2257 676
rect 168 525 433 573
rect 122 514 433 525
rect 387 464 433 514
rect 734 556 780 578
rect 74 424 318 430
rect 74 378 158 424
rect 204 378 318 424
rect 74 354 318 378
rect 387 418 618 464
rect 664 418 675 464
rect 387 311 433 418
rect 734 372 780 510
rect 387 245 433 265
rect 59 200 433 245
rect 105 198 433 200
rect 605 326 780 372
rect 605 177 651 326
rect 826 280 872 602
rect 1188 597 1440 602
rect 1852 568 1898 602
rect 1030 510 1043 556
rect 1089 551 1133 556
rect 1486 551 1539 556
rect 1089 510 1539 551
rect 1585 510 1800 556
rect 1852 525 2211 568
rect 1852 522 2257 525
rect 1030 505 1800 510
rect 923 424 1695 430
rect 923 378 1066 424
rect 1676 378 1695 424
rect 923 354 1695 378
rect 1754 380 1800 505
rect 2211 472 2257 522
rect 2404 665 2472 724
rect 2404 525 2415 665
rect 2461 525 2472 665
rect 2404 518 2472 525
rect 2619 665 2665 676
rect 2619 472 2665 525
rect 2812 665 2880 724
rect 2812 525 2823 665
rect 2869 525 2880 665
rect 2812 518 2880 525
rect 3027 665 3073 676
rect 3027 472 3073 525
rect 3234 665 3302 724
rect 3693 703 3739 724
rect 3234 525 3245 665
rect 3291 525 3302 665
rect 3234 518 3302 525
rect 3489 665 3535 676
rect 4141 703 4187 724
rect 3693 646 3739 657
rect 3917 665 3963 676
rect 3535 525 3917 572
rect 4589 703 4635 724
rect 4141 646 4187 657
rect 4365 665 4411 676
rect 3963 525 4365 572
rect 4997 703 5043 724
rect 4589 646 4635 657
rect 4793 665 4839 676
rect 4411 525 4793 572
rect 5405 703 5451 724
rect 4997 646 5043 657
rect 5201 665 5247 676
rect 4839 525 5201 572
rect 5405 646 5451 657
rect 5609 665 5656 676
rect 5247 525 5609 572
rect 5655 525 5656 665
rect 3489 492 5656 525
rect 5813 665 5859 724
rect 5813 506 5859 525
rect 2211 439 3301 472
rect 2211 426 3366 439
rect 3255 393 3366 426
rect 3412 393 3591 439
rect 3637 393 3817 439
rect 3863 393 4039 439
rect 4085 393 4251 439
rect 4297 393 4473 439
rect 4519 393 4530 439
rect 3255 392 4530 393
rect 1754 378 3193 380
rect 762 244 872 280
rect 1754 332 2004 378
rect 3178 332 3193 378
rect 1754 330 3193 332
rect 1754 279 1800 330
rect 3255 284 3362 319
rect 762 198 775 244
rect 821 198 872 244
rect 918 244 1800 279
rect 918 198 931 244
rect 977 233 1555 244
rect 977 198 990 233
rect 1542 198 1555 233
rect 1601 233 1800 244
rect 2211 273 3362 284
rect 3408 273 3591 319
rect 3637 273 3819 319
rect 3865 273 4038 319
rect 4084 273 4095 319
rect 2211 238 3301 273
rect 4608 253 4688 492
rect 4881 393 4892 439
rect 4938 393 5099 439
rect 5145 393 5305 439
rect 5351 393 5508 439
rect 5554 393 5711 439
rect 5757 393 5768 439
rect 4881 392 5768 393
rect 5372 273 5383 319
rect 5429 273 5608 319
rect 5654 273 5831 319
rect 5877 273 5897 319
rect 1601 198 1614 233
rect 2211 187 2257 238
rect 59 143 105 154
rect 507 166 651 177
rect 283 139 329 152
rect 553 152 651 166
rect 1138 152 1431 187
rect 1711 152 2135 187
rect 553 141 2135 152
rect 2181 141 2257 187
rect 2359 175 2405 186
rect 553 120 1184 141
rect 507 106 1184 120
rect 1385 106 1757 141
rect 283 60 329 93
rect 1230 60 1243 95
rect 0 49 1243 60
rect 1289 60 1302 95
rect 1854 60 1867 95
rect 1289 49 1867 60
rect 1913 60 1926 95
rect 2359 60 2405 129
rect 2583 175 2629 238
rect 2583 116 2629 129
rect 2807 175 2853 186
rect 2807 60 2853 129
rect 3031 175 3077 238
rect 4150 227 5322 253
rect 3424 219 5776 227
rect 3031 116 3077 129
rect 3255 175 3301 186
rect 3424 173 3479 219
rect 3525 173 3927 219
rect 3973 173 4375 219
rect 4421 173 4823 219
rect 4869 173 5271 219
rect 5317 173 5719 219
rect 5765 173 5776 219
rect 3255 60 3301 129
rect 5943 172 5989 183
rect 3692 81 3703 127
rect 3749 81 3760 127
rect 3692 60 3760 81
rect 4140 81 4151 127
rect 4197 81 4208 127
rect 4140 60 4208 81
rect 4588 81 4599 127
rect 4645 81 4656 127
rect 4588 60 4656 81
rect 5036 81 5047 127
rect 5093 81 5104 127
rect 5036 60 5104 81
rect 5445 81 5495 127
rect 5541 81 5552 127
rect 5445 60 5552 81
rect 5943 60 5989 126
rect 1913 49 6048 60
rect 0 -60 6048 49
<< labels >>
flabel metal1 s 0 724 6048 844 0 FreeSans 400 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 3255 183 3301 186 0 FreeSans 400 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel metal1 s 5609 572 5656 676 0 FreeSans 400 0 0 0 ZN
port 3 nsew default output
flabel metal1 s 74 354 318 430 0 FreeSans 400 0 0 0 EN
port 1 nsew default input
flabel metal1 s 923 354 1695 430 0 FreeSans 400 0 0 0 I
port 2 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 5 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 6 nsew ground bidirectional
rlabel metal1 s 5201 572 5247 676 1 ZN
port 3 nsew default output
rlabel metal1 s 4793 572 4839 676 1 ZN
port 3 nsew default output
rlabel metal1 s 4365 572 4411 676 1 ZN
port 3 nsew default output
rlabel metal1 s 3917 572 3963 676 1 ZN
port 3 nsew default output
rlabel metal1 s 3489 572 3535 676 1 ZN
port 3 nsew default output
rlabel metal1 s 3489 492 5656 572 1 ZN
port 3 nsew default output
rlabel metal1 s 4608 253 4688 492 1 ZN
port 3 nsew default output
rlabel metal1 s 4150 227 5322 253 1 ZN
port 3 nsew default output
rlabel metal1 s 3424 173 5776 227 1 ZN
port 3 nsew default output
rlabel metal1 s 5813 689 5859 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5405 689 5451 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4997 689 5043 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4589 689 4635 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4141 689 4187 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3693 689 3739 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3234 689 3302 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2812 689 2880 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2404 689 2472 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1963 689 2009 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1280 689 1348 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 326 689 372 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5813 646 5859 689 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5405 646 5451 689 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4997 646 5043 689 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4589 646 4635 689 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4141 646 4187 689 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3693 646 3739 689 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3234 646 3302 689 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2812 646 2880 689 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2404 646 2472 689 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1963 646 2009 689 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 326 646 372 689 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5813 626 5859 646 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3234 626 3302 646 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2812 626 2880 646 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2404 626 2472 646 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1963 626 2009 646 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 326 626 372 646 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5813 620 5859 626 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3234 620 3302 626 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2812 620 2880 626 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2404 620 2472 626 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1963 620 2009 626 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5813 518 5859 620 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3234 518 3302 620 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2812 518 2880 620 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2404 518 2472 620 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5813 506 5859 518 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2807 183 2853 186 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2359 183 2405 186 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5943 152 5989 183 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3255 152 3301 183 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2807 152 2853 183 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2359 152 2405 183 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5943 127 5989 152 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3255 127 3301 152 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2807 127 2853 152 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2359 127 2405 152 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 283 127 329 152 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5943 95 5989 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5445 95 5552 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5036 95 5104 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4588 95 4656 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4140 95 4208 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3692 95 3760 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3255 95 3301 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2807 95 2853 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2359 95 2405 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 283 95 329 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5943 60 5989 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5445 60 5552 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5036 60 5104 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4588 60 4656 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4140 60 4208 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3692 60 3760 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3255 60 3301 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2807 60 2853 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2359 60 2405 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1854 60 1926 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1230 60 1302 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 283 60 329 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 6048 60 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 6048 784
string GDS_END 564332
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 551338
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
